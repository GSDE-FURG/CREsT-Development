//Converted to Combinational (Partial output: n55) , Module name: s1494_n55 , Timestamp: 2018-12-03T15:51:02.651861 
module s1494_n55 ( v1, CLR, v7, v2, v10, v8, v9, v11, v12, v3, v0, v5, v4, v6, n55 );
input v1, CLR, v7, v2, v10, v8, v9, v11, v12, v3, v0, v5, v4, v6;
output n55;
wire n267, n283, n291, n68, n271, n282, n290, n285, n93, n268, n270, n281, n45, n275, n289, n64, n148, n284, n184, n139, n67, n70_1, n269, n277, n280, n279, n272, n83, n274, n286, n287, n288, n94, n203, n62, n100, n276, n140, n57, n87, n278, n109, n273, n107, n86, n174, n131, n123;
AOI21X1  g246(.A0(n291), .A1(n283), .B0(n267), .Y(n55));
INVX1    g221(.A(CLR), .Y(n267));
OAI21X1  g237(.A0(n282), .A1(n271), .B0(n68), .Y(n283));
AOI21X1  g245(.A0(n285), .A1(v7), .B0(n290), .Y(n291));
INVX1    g023(.A(v7), .Y(n68));
AOI21X1  g225(.A0(n270), .A1(n268), .B0(n93), .Y(n271));
OAI21X1  g236(.A0(n275), .A1(n45), .B0(n281), .Y(n282));
OAI22X1  g244(.A0(n148), .A1(n64), .B0(v2), .B1(n289), .Y(n290));
OAI22X1  g239(.A0(n139), .A1(n184), .B0(v10), .B1(n284), .Y(n285));
INVX1    g048(.A(v8), .Y(n93));
NAND4X1  g222(.A(n45), .B(v11), .C(n67), .D(v9), .Y(n268));
OAI21X1  g224(.A0(n269), .A1(n70_1), .B0(v10), .Y(n270));
AOI22X1  g235(.A0(n279), .A1(n280), .B0(n277), .B1(n93), .Y(n281));
INVX1    g000(.A(v10), .Y(n45));
AOI21X1  g229(.A0(n274), .A1(n83), .B0(n272), .Y(n275));
AOI21X1  g243(.A0(n288), .A1(n287), .B0(n286), .Y(n289));
OR2X1    g019(.A(v9), .B(v12), .Y(n64));
NAND2X1  g102(.A(v8), .B(v10), .Y(n148));
AOI22X1  g238(.A0(n203), .A1(n93), .B0(n64), .B1(n94), .Y(n284));
NAND2X1  g138(.A(v9), .B(v10), .Y(n184));
NAND2X1  g093(.A(v11), .B(n67), .Y(n139));
INVX1    g022(.A(v12), .Y(n67));
INVX1    g025(.A(v9), .Y(n70_1));
AOI21X1  g223(.A0(n100), .A1(n62), .B0(n139), .Y(n269));
OAI21X1  g231(.A0(n140), .A1(n70_1), .B0(n276), .Y(n277));
AND2X1   g234(.A(v12), .B(v3), .Y(n280));
OAI22X1  g233(.A0(n109), .A1(n278), .B0(n87), .B1(n57), .Y(n279));
NOR3X1   g226(.A(v9), .B(v11), .C(v12), .Y(n272));
INVX1    g038(.A(v0), .Y(n83));
OAI22X1  g228(.A0(n100), .A1(n64), .B0(n107), .B1(n273), .Y(n274));
NOR3X1   g240(.A(n140), .B(n93), .C(v9), .Y(n286));
NOR3X1   g241(.A(n131), .B(n174), .C(n86), .Y(n287));
NOR3X1   g242(.A(n87), .B(v8), .C(n70_1), .Y(n288));
NOR2X1   g049(.A(n93), .B(v11), .Y(n94));
INVX1    g157(.A(n139), .Y(n203));
INVX1    g017(.A(v2), .Y(n62));
NAND2X1  g055(.A(v4), .B(v5), .Y(n100));
NAND4X1  g230(.A(n70_1), .B(v12), .C(v6), .D(n123), .Y(n276));
NAND2X1  g094(.A(v10), .B(v11), .Y(n140));
OR2X1    g012(.A(v8), .B(v9), .Y(n57));
OR2X1    g042(.A(v10), .B(v11), .Y(n87));
NAND4X1  g232(.A(v10), .B(v11), .C(v0), .D(v8), .Y(n278));
NOR2X1   g064(.A(v1), .B(n86), .Y(n109));
NAND4X1  g227(.A(n174), .B(v3), .C(v6), .D(v8), .Y(n273));
NAND2X1  g062(.A(v11), .B(v12), .Y(n107));
INVX1    g041(.A(v6), .Y(n86));
INVX1    g128(.A(v1), .Y(n174));
OR2X1    g085(.A(v7), .B(v12), .Y(n131));
NOR2X1   g077(.A(v10), .B(v11), .Y(n123));

endmodule
