//Converted to Combinational (Partial output: n90) , Module name: s832_n90
module s832_n90 ( G1, G3, G4, G18, G38, G0, G40, G41, G42, G39, G2, G15, G16, G9, G6, G7, G8, G13, G14, G5, n90 );
input G1, G3, G4, G18, G38, G0, G40, G41, G42, G39, G2, G15, G16, G9, G6, G7, G8, G13, G14, G5;
output n90;
wire n200, n218, n76, n191, n199, n217, n208, n212, n213, n190, n186, n187, n188, n193, n196, n198, n197, n214, n215, n216, n207, n202, n204, n205, n209, n211, n86, n73, n78, n189, n172, n62, n174, n185, n53, n114, n192, n194, n195, n80_1, n61, n147, n66, n57, n60, n206, n95_1, n96, n201, n203, n210, n102, n54, n52, n109;
AOI21X1  g165(.A0(n218), .A1(n200), .B0(G18), .Y(n90));
OAI21X1  g146(.A0(n199), .A1(n191), .B0(n76), .Y(n200));
NOR4X1   g164(.A(n213), .B(n212), .C(n208), .D(n217), .Y(n218));
INVX1    g024(.A(G38), .Y(n76));
NOR4X1   g137(.A(n188), .B(n187), .C(n186), .D(n190), .Y(n191));
OAI22X1  g145(.A0(n197), .A1(n198), .B0(n196), .B1(n193), .Y(n199));
NOR3X1   g163(.A(n216), .B(n215), .C(n214), .Y(n217));
NOR4X1   g154(.A(n205), .B(n204), .C(n202), .D(n207), .Y(n208));
NOR2X1   g158(.A(n211), .B(n209), .Y(n212));
NOR3X1   g159(.A(n209), .B(n86), .C(G0), .Y(n213));
OAI22X1  g136(.A0(n172), .A1(n189), .B0(n78), .B1(n73), .Y(n190));
NOR3X1   g132(.A(n185), .B(n174), .C(n62), .Y(n186));
NOR3X1   g133(.A(G42), .B(G41), .C(G40), .Y(n187));
OAI21X1  g134(.A0(n114), .A1(n73), .B0(n53), .Y(n188));
NOR2X1   g139(.A(n192), .B(G39), .Y(n193));
NAND2X1  g142(.A(n195), .B(n194), .Y(n196));
NAND4X1  g144(.A(n147), .B(G2), .C(n61), .D(n80_1), .Y(n198));
AOI22X1  g143(.A0(n57), .A1(G42), .B0(n62), .B1(n66), .Y(n197));
NAND4X1  g160(.A(n114), .B(G39), .C(n73), .D(n78), .Y(n214));
NOR2X1   g161(.A(n60), .B(n62), .Y(n215));
NOR3X1   g162(.A(G41), .B(n62), .C(G15), .Y(n216));
OAI21X1  g153(.A0(n95_1), .A1(G42), .B0(n206), .Y(n207));
NOR2X1   g148(.A(n201), .B(n96), .Y(n202));
OAI21X1  g150(.A0(G39), .A1(n76), .B0(n203), .Y(n204));
AOI21X1  g151(.A0(G42), .A1(G15), .B0(G41), .Y(n205));
NAND3X1  g155(.A(G42), .B(G41), .C(G40), .Y(n209));
NAND3X1  g157(.A(n210), .B(n53), .C(n73), .Y(n211));
NAND2X1  g034(.A(G39), .B(G38), .Y(n86));
INVX1    g021(.A(G4), .Y(n73));
NAND2X1  g026(.A(G42), .B(G41), .Y(n78));
OR2X1    g135(.A(G42), .B(G40), .Y(n189));
NAND2X1  g118(.A(G15), .B(n102), .Y(n172));
INVX1    g010(.A(G16), .Y(n62));
NOR2X1   g120(.A(G42), .B(G40), .Y(n174));
NOR4X1   g131(.A(G41), .B(n114), .C(n52), .D(n54), .Y(n185));
INVX1    g001(.A(G39), .Y(n53));
INVX1    g060(.A(G40), .Y(n114));
NOR3X1   g138(.A(G42), .B(n80_1), .C(G4), .Y(n192));
AOI21X1  g140(.A0(n80_1), .A1(n109), .B0(n114), .Y(n194));
OAI21X1  g141(.A0(n80_1), .A1(G16), .B0(G42), .Y(n195));
INVX1    g028(.A(G41), .Y(n80_1));
INVX1    g009(.A(G1), .Y(n61));
INVX1    g093(.A(G3), .Y(n147));
NOR2X1   g014(.A(G40), .B(G39), .Y(n66));
AND2X1   g005(.A(G40), .B(G39), .Y(n57));
OR2X1    g008(.A(G42), .B(G41), .Y(n60));
AOI21X1  g152(.A0(n53), .A1(G15), .B0(G4), .Y(n206));
NAND2X1  g043(.A(G38), .B(G15), .Y(n95_1));
NAND4X1  g044(.A(G8), .B(G7), .C(G6), .D(G9), .Y(n96));
AOI21X1  g147(.A0(G38), .A1(G15), .B0(n80_1), .Y(n201));
NOR2X1   g149(.A(G40), .B(n62), .Y(n203));
NAND3X1  g156(.A(G16), .B(G15), .C(G13), .Y(n210));
INVX1    g048(.A(G14), .Y(n102));
INVX1    g002(.A(G42), .Y(n54));
INVX1    g000(.A(G15), .Y(n52));
INVX1    g055(.A(G5), .Y(n109));

endmodule
