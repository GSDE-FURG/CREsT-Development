// Benchmark "b08_C" written by ABC on Wed Aug 05 14:39:06 2020

module b08_C ( 
    O_REG_0__SCAN_IN, START, I_7_, I_6_, I_5_, I_4_, I_3_, I_2_, I_1_,
    I_0_, STATO_REG_1__SCAN_IN, STATO_REG_0__SCAN_IN, MAR_REG_2__SCAN_IN,
    MAR_REG_1__SCAN_IN, MAR_REG_0__SCAN_IN, IN_R_REG_7__SCAN_IN,
    IN_R_REG_6__SCAN_IN, IN_R_REG_5__SCAN_IN, IN_R_REG_4__SCAN_IN,
    IN_R_REG_3__SCAN_IN, IN_R_REG_2__SCAN_IN, IN_R_REG_1__SCAN_IN,
    IN_R_REG_0__SCAN_IN, OUT_R_REG_3__SCAN_IN, OUT_R_REG_2__SCAN_IN,
    OUT_R_REG_1__SCAN_IN, OUT_R_REG_0__SCAN_IN, O_REG_3__SCAN_IN,
    O_REG_2__SCAN_IN, O_REG_1__SCAN_IN,
    U189, U188, U187, U206, U207, U208, U209, U210, U211, U212, U213, U214,
    U215, U186, U185, U184, U183, U216, U217, U218, U219  );
  input  O_REG_0__SCAN_IN, START, I_7_, I_6_, I_5_, I_4_, I_3_, I_2_,
    I_1_, I_0_, STATO_REG_1__SCAN_IN, STATO_REG_0__SCAN_IN,
    MAR_REG_2__SCAN_IN, MAR_REG_1__SCAN_IN, MAR_REG_0__SCAN_IN,
    IN_R_REG_7__SCAN_IN, IN_R_REG_6__SCAN_IN, IN_R_REG_5__SCAN_IN,
    IN_R_REG_4__SCAN_IN, IN_R_REG_3__SCAN_IN, IN_R_REG_2__SCAN_IN,
    IN_R_REG_1__SCAN_IN, IN_R_REG_0__SCAN_IN, OUT_R_REG_3__SCAN_IN,
    OUT_R_REG_2__SCAN_IN, OUT_R_REG_1__SCAN_IN, OUT_R_REG_0__SCAN_IN,
    O_REG_3__SCAN_IN, O_REG_2__SCAN_IN, O_REG_1__SCAN_IN;
  output U189, U188, U187, U206, U207, U208, U209, U210, U211, U212, U213,
    U214, U215, U186, U185, U184, U183, U216, U217, U218, U219;
  wire n55, n56, n57, n58, n59, n60, n62, n63, n65, n66, n67, n68, n69, n71,
    n72, n73, n74, n76, n78, n79, n81, n82, n84, n85, n87, n88, n90, n91,
    n93, n94, n96, n97, n99, n100, n102, n103, n104, n105, n106, n107,
    n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
    n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
    n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
    n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
    n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
    n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
    n181, n182, n183, n185, n186, n187, n189, n191, n192, n193, n195, n196,
    n198, n199, n201, n202;
  NAND3X1 g000(.A(MAR_REG_0__SCAN_IN), .B(MAR_REG_1__SCAN_IN), .C(MAR_REG_2__SCAN_IN), .Y(n55));
  OAI21X1 g001(.A0(n55), .A1(START), .B0(STATO_REG_0__SCAN_IN), .Y(n56));
  INVX1   g002(.A(STATO_REG_1__SCAN_IN), .Y(n57));
  NAND2X1 g003(.A(STATO_REG_0__SCAN_IN), .B(n57), .Y(n58));
  NOR2X1  g004(.A(STATO_REG_0__SCAN_IN), .B(n57), .Y(n59));
  INVX1   g005(.A(n59), .Y(n60));
  NAND3X1 g006(.A(n60), .B(n58), .C(n56), .Y(U189));
  OAI21X1 g007(.A0(n55), .A1(n57), .B0(STATO_REG_0__SCAN_IN), .Y(n62));
  NAND2X1 g008(.A(n62), .B(START), .Y(n63));
  NAND2X1 g009(.A(n63), .B(n60), .Y(U188));
  NAND2X1 g010(.A(STATO_REG_0__SCAN_IN), .B(STATO_REG_1__SCAN_IN), .Y(n65));
  INVX1   g011(.A(MAR_REG_2__SCAN_IN), .Y(n66));
  NAND3X1 g012(.A(MAR_REG_0__SCAN_IN), .B(MAR_REG_1__SCAN_IN), .C(n66), .Y(n67));
  INVX1   g013(.A(STATO_REG_0__SCAN_IN), .Y(n68));
  OAI21X1 g014(.A0(n68), .A1(STATO_REG_1__SCAN_IN), .B0(MAR_REG_2__SCAN_IN), .Y(n69));
  OAI21X1 g015(.A0(n67), .A1(n65), .B0(n69), .Y(U187));
  INVX1   g016(.A(MAR_REG_1__SCAN_IN), .Y(n71));
  NAND4X1 g017(.A(n71), .B(STATO_REG_0__SCAN_IN), .C(STATO_REG_1__SCAN_IN), .D(MAR_REG_0__SCAN_IN), .Y(n72));
  INVX1   g018(.A(MAR_REG_0__SCAN_IN), .Y(n73));
  AOI21X1 g019(.A0(n73), .A1(STATO_REG_1__SCAN_IN), .B0(n62), .Y(n74));
  OAI21X1 g020(.A0(n74), .A1(n71), .B0(n72), .Y(U206));
  NAND2X1 g021(.A(n62), .B(MAR_REG_0__SCAN_IN), .Y(n76));
  OAI21X1 g022(.A0(n65), .A1(MAR_REG_0__SCAN_IN), .B0(n76), .Y(U207));
  NAND3X1 g023(.A(STATO_REG_0__SCAN_IN), .B(n57), .C(I_7_), .Y(n78));
  OAI21X1 g024(.A0(n68), .A1(STATO_REG_1__SCAN_IN), .B0(IN_R_REG_7__SCAN_IN), .Y(n79));
  NAND2X1 g025(.A(n79), .B(n78), .Y(U208));
  NAND3X1 g026(.A(STATO_REG_0__SCAN_IN), .B(n57), .C(I_6_), .Y(n81));
  OAI21X1 g027(.A0(n68), .A1(STATO_REG_1__SCAN_IN), .B0(IN_R_REG_6__SCAN_IN), .Y(n82));
  NAND2X1 g028(.A(n82), .B(n81), .Y(U209));
  NAND3X1 g029(.A(STATO_REG_0__SCAN_IN), .B(n57), .C(I_5_), .Y(n84));
  OAI21X1 g030(.A0(n68), .A1(STATO_REG_1__SCAN_IN), .B0(IN_R_REG_5__SCAN_IN), .Y(n85));
  NAND2X1 g031(.A(n85), .B(n84), .Y(U210));
  NAND3X1 g032(.A(STATO_REG_0__SCAN_IN), .B(n57), .C(I_4_), .Y(n87));
  OAI21X1 g033(.A0(n68), .A1(STATO_REG_1__SCAN_IN), .B0(IN_R_REG_4__SCAN_IN), .Y(n88));
  NAND2X1 g034(.A(n88), .B(n87), .Y(U211));
  NAND3X1 g035(.A(STATO_REG_0__SCAN_IN), .B(n57), .C(I_3_), .Y(n90));
  OAI21X1 g036(.A0(n68), .A1(STATO_REG_1__SCAN_IN), .B0(IN_R_REG_3__SCAN_IN), .Y(n91));
  NAND2X1 g037(.A(n91), .B(n90), .Y(U212));
  NAND3X1 g038(.A(STATO_REG_0__SCAN_IN), .B(n57), .C(I_2_), .Y(n93));
  OAI21X1 g039(.A0(n68), .A1(STATO_REG_1__SCAN_IN), .B0(IN_R_REG_2__SCAN_IN), .Y(n94));
  NAND2X1 g040(.A(n94), .B(n93), .Y(U213));
  NAND3X1 g041(.A(STATO_REG_0__SCAN_IN), .B(n57), .C(I_1_), .Y(n96));
  OAI21X1 g042(.A0(n68), .A1(STATO_REG_1__SCAN_IN), .B0(IN_R_REG_1__SCAN_IN), .Y(n97));
  NAND2X1 g043(.A(n97), .B(n96), .Y(U214));
  NAND3X1 g044(.A(STATO_REG_0__SCAN_IN), .B(n57), .C(I_0_), .Y(n99));
  OAI21X1 g045(.A0(n68), .A1(STATO_REG_1__SCAN_IN), .B0(IN_R_REG_0__SCAN_IN), .Y(n100));
  NAND2X1 g046(.A(n100), .B(n99), .Y(U215));
  NAND3X1 g047(.A(n73), .B(n71), .C(n66), .Y(n102));
  NAND2X1 g048(.A(n71), .B(MAR_REG_2__SCAN_IN), .Y(n103));
  NAND3X1 g049(.A(n103), .B(n102), .C(n67), .Y(n104));
  NOR3X1  g050(.A(n73), .B(n71), .C(MAR_REG_2__SCAN_IN), .Y(n105));
  NOR2X1  g051(.A(MAR_REG_1__SCAN_IN), .B(n66), .Y(n106));
  AOI21X1 g052(.A0(MAR_REG_0__SCAN_IN), .A1(n66), .B0(n71), .Y(n107));
  NOR4X1  g053(.A(n106), .B(n105), .C(IN_R_REG_5__SCAN_IN), .D(n107), .Y(n108));
  NOR3X1  g054(.A(MAR_REG_0__SCAN_IN), .B(MAR_REG_1__SCAN_IN), .C(MAR_REG_2__SCAN_IN), .Y(n109));
  NOR3X1  g055(.A(n73), .B(MAR_REG_1__SCAN_IN), .C(n66), .Y(n110));
  NAND3X1 g056(.A(n73), .B(n71), .C(MAR_REG_2__SCAN_IN), .Y(n111));
  NAND3X1 g057(.A(n73), .B(MAR_REG_1__SCAN_IN), .C(n66), .Y(n112));
  NAND3X1 g058(.A(MAR_REG_0__SCAN_IN), .B(n71), .C(n66), .Y(n113));
  NAND4X1 g059(.A(n112), .B(n111), .C(n55), .D(n113), .Y(n114));
  NOR4X1  g060(.A(n110), .B(n109), .C(IN_R_REG_7__SCAN_IN), .D(n114), .Y(n115));
  INVX1   g061(.A(IN_R_REG_5__SCAN_IN), .Y(n116));
  NOR4X1  g062(.A(MAR_REG_0__SCAN_IN), .B(n71), .C(n66), .D(n116), .Y(n117));
  NOR3X1  g063(.A(n117), .B(n115), .C(n108), .Y(n118));
  INVX1   g064(.A(IN_R_REG_4__SCAN_IN), .Y(n119));
  OAI21X1 g065(.A0(n107), .A1(n106), .B0(n119), .Y(n120));
  OAI21X1 g066(.A0(n106), .A1(n105), .B0(IN_R_REG_4__SCAN_IN), .Y(n121));
  NAND4X1 g067(.A(n120), .B(n113), .C(n102), .D(n121), .Y(n122));
  NOR3X1  g068(.A(n110), .B(n105), .C(IN_R_REG_3__SCAN_IN), .Y(n123));
  NAND3X1 g069(.A(n123), .B(n112), .C(n55), .Y(n124));
  NOR2X1  g070(.A(n106), .B(n105), .Y(n125));
  INVX1   g071(.A(IN_R_REG_7__SCAN_IN), .Y(n126));
  NOR3X1  g072(.A(MAR_REG_0__SCAN_IN), .B(n71), .C(n66), .Y(n127));
  NOR3X1  g073(.A(MAR_REG_0__SCAN_IN), .B(n71), .C(MAR_REG_2__SCAN_IN), .Y(n128));
  NOR3X1  g074(.A(n128), .B(n127), .C(n126), .Y(n129));
  AOI21X1 g075(.A0(n129), .A1(n125), .B0(n60), .Y(n130));
  NAND4X1 g076(.A(n124), .B(n122), .C(n118), .D(n130), .Y(n131));
  INVX1   g077(.A(IN_R_REG_2__SCAN_IN), .Y(n132));
  OAI21X1 g078(.A0(n114), .A1(n127), .B0(n132), .Y(n133));
  NAND3X1 g079(.A(n103), .B(n67), .C(n55), .Y(n134));
  AOI21X1 g080(.A0(n134), .A1(IN_R_REG_2__SCAN_IN), .B0(n109), .Y(n135));
  INVX1   g081(.A(IN_R_REG_6__SCAN_IN), .Y(n136));
  OAI21X1 g082(.A0(n114), .A1(n105), .B0(n136), .Y(n137));
  AOI21X1 g083(.A0(n104), .A1(IN_R_REG_6__SCAN_IN), .B0(n127), .Y(n138));
  AOI22X1 g084(.A0(n137), .A1(n138), .B0(n135), .B1(n133), .Y(n139));
  OAI21X1 g085(.A0(n134), .A1(n127), .B0(IN_R_REG_1__SCAN_IN), .Y(n140));
  INVX1   g086(.A(IN_R_REG_1__SCAN_IN), .Y(n141));
  NAND2X1 g087(.A(n103), .B(n67), .Y(n142));
  NAND3X1 g088(.A(n113), .B(n112), .C(n55), .Y(n143));
  OAI21X1 g089(.A0(n143), .A1(n142), .B0(n141), .Y(n144));
  NAND3X1 g090(.A(n144), .B(n140), .C(n102), .Y(n145));
  NOR3X1  g091(.A(n73), .B(MAR_REG_1__SCAN_IN), .C(MAR_REG_2__SCAN_IN), .Y(n146));
  OAI21X1 g092(.A0(n134), .A1(n146), .B0(IN_R_REG_0__SCAN_IN), .Y(n147));
  OAI21X1 g093(.A0(n73), .A1(MAR_REG_2__SCAN_IN), .B0(MAR_REG_1__SCAN_IN), .Y(n148));
  AOI21X1 g094(.A0(n148), .A1(n67), .B0(IN_R_REG_0__SCAN_IN), .Y(n149));
  NOR2X1  g095(.A(n149), .B(n109), .Y(n150));
  NAND2X1 g096(.A(n150), .B(n147), .Y(n151));
  NAND3X1 g097(.A(n151), .B(n145), .C(n139), .Y(n152));
  OAI21X1 g098(.A0(n152), .A1(n131), .B0(n58), .Y(n153));
  NAND3X1 g099(.A(n153), .B(n104), .C(STATO_REG_1__SCAN_IN), .Y(n154));
  NAND3X1 g100(.A(n130), .B(n124), .C(n122), .Y(n155));
  NOR4X1  g101(.A(n117), .B(n115), .C(n108), .D(n155), .Y(n156));
  NAND3X1 g102(.A(n73), .B(MAR_REG_1__SCAN_IN), .C(MAR_REG_2__SCAN_IN), .Y(n157));
  NOR3X1  g103(.A(n73), .B(n71), .C(n66), .Y(n158));
  NOR3X1  g104(.A(MAR_REG_0__SCAN_IN), .B(MAR_REG_1__SCAN_IN), .C(n66), .Y(n159));
  NOR4X1  g105(.A(n128), .B(n159), .C(n158), .D(n146), .Y(n160));
  AOI21X1 g106(.A0(n160), .A1(n157), .B0(IN_R_REG_2__SCAN_IN), .Y(n161));
  NOR3X1  g107(.A(n106), .B(n105), .C(n158), .Y(n162));
  OAI21X1 g108(.A0(n162), .A1(n132), .B0(n102), .Y(n163));
  AOI21X1 g109(.A0(n160), .A1(n67), .B0(IN_R_REG_6__SCAN_IN), .Y(n164));
  NOR3X1  g110(.A(n106), .B(n109), .C(n105), .Y(n165));
  OAI21X1 g111(.A0(n165), .A1(n136), .B0(n157), .Y(n166));
  OAI22X1 g112(.A0(n164), .A1(n166), .B0(n163), .B1(n161), .Y(n167));
  AOI21X1 g113(.A0(n162), .A1(n157), .B0(n141), .Y(n168));
  NOR3X1  g114(.A(n146), .B(n128), .C(n158), .Y(n169));
  AOI21X1 g115(.A0(n169), .A1(n125), .B0(IN_R_REG_1__SCAN_IN), .Y(n170));
  NOR3X1  g116(.A(n170), .B(n168), .C(n109), .Y(n171));
  INVX1   g117(.A(IN_R_REG_0__SCAN_IN), .Y(n172));
  AOI21X1 g118(.A0(n162), .A1(n113), .B0(n172), .Y(n173));
  NOR3X1  g119(.A(n149), .B(n173), .C(n109), .Y(n174));
  NOR3X1  g120(.A(n174), .B(n171), .C(n167), .Y(n175));
  AOI22X1 g121(.A0(n156), .A1(n175), .B0(STATO_REG_0__SCAN_IN), .B1(n57), .Y(n176));
  OAI21X1 g122(.A0(n176), .A1(STATO_REG_1__SCAN_IN), .B0(OUT_R_REG_3__SCAN_IN), .Y(n177));
  NAND2X1 g123(.A(n112), .B(n157), .Y(n178));
  NAND3X1 g124(.A(n153), .B(n178), .C(STATO_REG_1__SCAN_IN), .Y(n179));
  NAND3X1 g125(.A(n179), .B(n177), .C(n154), .Y(U186));
  OAI21X1 g126(.A0(n176), .A1(STATO_REG_1__SCAN_IN), .B0(OUT_R_REG_2__SCAN_IN), .Y(n181));
  NAND3X1 g127(.A(n112), .B(n111), .C(n55), .Y(n182));
  NAND3X1 g128(.A(n153), .B(n182), .C(STATO_REG_1__SCAN_IN), .Y(n183));
  NAND2X1 g129(.A(n183), .B(n181), .Y(U185));
  OAI21X1 g130(.A0(n176), .A1(STATO_REG_1__SCAN_IN), .B0(OUT_R_REG_1__SCAN_IN), .Y(n185));
  NAND4X1 g131(.A(n111), .B(n102), .C(n67), .D(n113), .Y(n186));
  NAND3X1 g132(.A(n186), .B(n153), .C(STATO_REG_1__SCAN_IN), .Y(n187));
  NAND3X1 g133(.A(n187), .B(n185), .C(n179), .Y(U184));
  OAI21X1 g134(.A0(n176), .A1(STATO_REG_1__SCAN_IN), .B0(OUT_R_REG_0__SCAN_IN), .Y(n189));
  NAND2X1 g135(.A(n189), .B(n179), .Y(U183));
  INVX1   g136(.A(O_REG_3__SCAN_IN), .Y(n191));
  NOR3X1  g137(.A(n65), .B(n55), .C(START), .Y(n192));
  NAND2X1 g138(.A(n192), .B(OUT_R_REG_3__SCAN_IN), .Y(n193));
  OAI21X1 g139(.A0(n192), .A1(n191), .B0(n193), .Y(U216));
  INVX1   g140(.A(O_REG_2__SCAN_IN), .Y(n195));
  NAND2X1 g141(.A(n192), .B(OUT_R_REG_2__SCAN_IN), .Y(n196));
  OAI21X1 g142(.A0(n192), .A1(n195), .B0(n196), .Y(U217));
  INVX1   g143(.A(O_REG_1__SCAN_IN), .Y(n198));
  NAND2X1 g144(.A(n192), .B(OUT_R_REG_1__SCAN_IN), .Y(n199));
  OAI21X1 g145(.A0(n192), .A1(n198), .B0(n199), .Y(U218));
  INVX1   g146(.A(O_REG_0__SCAN_IN), .Y(n201));
  NAND2X1 g147(.A(n192), .B(OUT_R_REG_0__SCAN_IN), .Y(n202));
  OAI21X1 g148(.A0(n192), .A1(n201), .B0(n202), .Y(U219));
endmodule


