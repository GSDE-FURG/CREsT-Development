//Converted to Combinational (Partial output: n8450) , Module name: s35932_n8450 , Timestamp: 2018-12-03T15:51:10.543058 
module s35932_n8450 ( RESET, TM1, DATA_0_0, TM0, WX10891, WX11115, WX11243, WX11051, WX11179, WX11181, WX11183, WX11185, WX11187, WX11189, WX11191, WX11193, WX11195, WX11197, WX11199, WX11201, WX11203, WX11205, WX11207, WX11209, WX11211, WX11213, WX11215, WX11217, WX11219, WX11221, WX11223, WX11225, WX11227, WX11229, WX11231, WX11233, WX11235, WX11237, WX11239, WX11241, n8450 );
input RESET, TM1, DATA_0_0, TM0, WX10891, WX11115, WX11243, WX11051, WX11179, WX11181, WX11183, WX11185, WX11187, WX11189, WX11191, WX11193, WX11195, WX11197, WX11199, WX11201, WX11203, WX11205, WX11207, WX11209, WX11211, WX11213, WX11215, WX11217, WX11219, WX11221, WX11223, WX11225, WX11227, WX11229, WX11231, WX11233, WX11235, WX11237, WX11239, WX11241;
output n8450;
wire n5827, n10651, n10650, n10648, n5539, n10259, n10649, n10647, n10256, n10258, CRC_OUT_1_0, n10255, n10257, n10749, CRC_OUT_1_31, n10814, CRC_OUT_1_30, n10812, CRC_OUT_1_29, n10810, CRC_OUT_1_28, n10808, CRC_OUT_1_27, n10806, CRC_OUT_1_26, n10804, CRC_OUT_1_25, n10802, CRC_OUT_1_24, n10800, CRC_OUT_1_23, n10798, CRC_OUT_1_22, n10796, CRC_OUT_1_21, n10794, CRC_OUT_1_20, n10792, CRC_OUT_1_19, n10790, CRC_OUT_1_18, n10788, CRC_OUT_1_17, n10786, CRC_OUT_1_16, n10784, CRC_OUT_1_15, n10783, n10781, CRC_OUT_1_14, n10779, CRC_OUT_1_13, n10777, CRC_OUT_1_12, n10775, CRC_OUT_1_11, n10773, CRC_OUT_1_10, n10772, n10770, CRC_OUT_1_9, n10768, CRC_OUT_1_8, n10766, CRC_OUT_1_7, n10764, CRC_OUT_1_6, n10762, CRC_OUT_1_5, n10760, CRC_OUT_1_4, n10758, CRC_OUT_1_3, n10757, n10755, CRC_OUT_1_2, n10753, CRC_OUT_1_1, n10751;
NOR2X1   g4857(.A(n10651), .B(n5827), .Y(n8450));
INVX1    g0288(.A(RESET), .Y(n5827));
MX2X1    g4856(.A(n10648), .B(n10650), .S0(TM1), .Y(n10651));
MX2X1    g4855(.A(n10649), .B(n10259), .S0(n5539), .Y(n10650));
AOI21X1  g4853(.A0(n5539), .A1(DATA_0_0), .B0(n10647), .Y(n10648));
INVX1    g0000(.A(TM0), .Y(n5539));
XOR2X1   g4465(.A(n10258), .B(n10256), .Y(n10259));
INVX1    g4854(.A(WX10891), .Y(n10649));
AND2X1   g4852(.A(CRC_OUT_1_0), .B(TM0), .Y(n10647));
XOR2X1   g4462(.A(n10255), .B(WX11115), .Y(n10256));
XOR2X1   g4464(.A(WX11243), .B(n10257), .Y(n10258));
NOR2X1   g4955(.A(n10749), .B(n5827), .Y(CRC_OUT_1_0));
XOR2X1   g4461(.A(WX11051), .B(TM0), .Y(n10255));
INVX1    g4463(.A(WX11179), .Y(n10257));
XOR2X1   g4954(.A(CRC_OUT_1_31), .B(WX11243), .Y(n10749));
NOR2X1   g5020(.A(n10814), .B(n5827), .Y(CRC_OUT_1_31));
XOR2X1   g5019(.A(CRC_OUT_1_30), .B(WX11181), .Y(n10814));
NOR2X1   g5018(.A(n10812), .B(n5827), .Y(CRC_OUT_1_30));
XOR2X1   g5017(.A(CRC_OUT_1_29), .B(WX11183), .Y(n10812));
NOR2X1   g5016(.A(n10810), .B(n5827), .Y(CRC_OUT_1_29));
XOR2X1   g5015(.A(CRC_OUT_1_28), .B(WX11185), .Y(n10810));
NOR2X1   g5014(.A(n10808), .B(n5827), .Y(CRC_OUT_1_28));
XOR2X1   g5013(.A(CRC_OUT_1_27), .B(WX11187), .Y(n10808));
NOR2X1   g5012(.A(n10806), .B(n5827), .Y(CRC_OUT_1_27));
XOR2X1   g5011(.A(CRC_OUT_1_26), .B(WX11189), .Y(n10806));
NOR2X1   g5010(.A(n10804), .B(n5827), .Y(CRC_OUT_1_26));
XOR2X1   g5009(.A(CRC_OUT_1_25), .B(WX11191), .Y(n10804));
NOR2X1   g5008(.A(n10802), .B(n5827), .Y(CRC_OUT_1_25));
XOR2X1   g5007(.A(CRC_OUT_1_24), .B(WX11193), .Y(n10802));
NOR2X1   g5006(.A(n10800), .B(n5827), .Y(CRC_OUT_1_24));
XOR2X1   g5005(.A(CRC_OUT_1_23), .B(WX11195), .Y(n10800));
NOR2X1   g5004(.A(n10798), .B(n5827), .Y(CRC_OUT_1_23));
XOR2X1   g5003(.A(CRC_OUT_1_22), .B(WX11197), .Y(n10798));
NOR2X1   g5002(.A(n10796), .B(n5827), .Y(CRC_OUT_1_22));
XOR2X1   g5001(.A(CRC_OUT_1_21), .B(WX11199), .Y(n10796));
NOR2X1   g5000(.A(n10794), .B(n5827), .Y(CRC_OUT_1_21));
XOR2X1   g4999(.A(CRC_OUT_1_20), .B(WX11201), .Y(n10794));
NOR2X1   g4998(.A(n10792), .B(n5827), .Y(CRC_OUT_1_20));
XOR2X1   g4997(.A(CRC_OUT_1_19), .B(WX11203), .Y(n10792));
NOR2X1   g4996(.A(n10790), .B(n5827), .Y(CRC_OUT_1_19));
XOR2X1   g4995(.A(CRC_OUT_1_18), .B(WX11205), .Y(n10790));
NOR2X1   g4994(.A(n10788), .B(n5827), .Y(CRC_OUT_1_18));
XOR2X1   g4993(.A(CRC_OUT_1_17), .B(WX11207), .Y(n10788));
NOR2X1   g4992(.A(n10786), .B(n5827), .Y(CRC_OUT_1_17));
XOR2X1   g4991(.A(CRC_OUT_1_16), .B(WX11209), .Y(n10786));
NOR2X1   g4990(.A(n10784), .B(n5827), .Y(CRC_OUT_1_16));
XOR2X1   g4989(.A(n10783), .B(CRC_OUT_1_15), .Y(n10784));
NOR2X1   g4987(.A(n10781), .B(n5827), .Y(CRC_OUT_1_15));
XOR2X1   g4988(.A(CRC_OUT_1_31), .B(WX11211), .Y(n10783));
XOR2X1   g4986(.A(CRC_OUT_1_14), .B(WX11213), .Y(n10781));
NOR2X1   g4985(.A(n10779), .B(n5827), .Y(CRC_OUT_1_14));
XOR2X1   g4984(.A(CRC_OUT_1_13), .B(WX11215), .Y(n10779));
NOR2X1   g4983(.A(n10777), .B(n5827), .Y(CRC_OUT_1_13));
XOR2X1   g4982(.A(CRC_OUT_1_12), .B(WX11217), .Y(n10777));
NOR2X1   g4981(.A(n10775), .B(n5827), .Y(CRC_OUT_1_12));
XOR2X1   g4980(.A(CRC_OUT_1_11), .B(WX11219), .Y(n10775));
NOR2X1   g4979(.A(n10773), .B(n5827), .Y(CRC_OUT_1_11));
XOR2X1   g4978(.A(n10772), .B(CRC_OUT_1_10), .Y(n10773));
NOR2X1   g4976(.A(n10770), .B(n5827), .Y(CRC_OUT_1_10));
XOR2X1   g4977(.A(CRC_OUT_1_31), .B(WX11221), .Y(n10772));
XOR2X1   g4975(.A(CRC_OUT_1_9), .B(WX11223), .Y(n10770));
NOR2X1   g4974(.A(n10768), .B(n5827), .Y(CRC_OUT_1_9));
XOR2X1   g4973(.A(CRC_OUT_1_8), .B(WX11225), .Y(n10768));
NOR2X1   g4972(.A(n10766), .B(n5827), .Y(CRC_OUT_1_8));
XOR2X1   g4971(.A(CRC_OUT_1_7), .B(WX11227), .Y(n10766));
NOR2X1   g4970(.A(n10764), .B(n5827), .Y(CRC_OUT_1_7));
XOR2X1   g4969(.A(CRC_OUT_1_6), .B(WX11229), .Y(n10764));
NOR2X1   g4968(.A(n10762), .B(n5827), .Y(CRC_OUT_1_6));
XOR2X1   g4967(.A(CRC_OUT_1_5), .B(WX11231), .Y(n10762));
NOR2X1   g4966(.A(n10760), .B(n5827), .Y(CRC_OUT_1_5));
XOR2X1   g4965(.A(CRC_OUT_1_4), .B(WX11233), .Y(n10760));
NOR2X1   g4964(.A(n10758), .B(n5827), .Y(CRC_OUT_1_4));
XOR2X1   g4963(.A(n10757), .B(CRC_OUT_1_3), .Y(n10758));
NOR2X1   g4961(.A(n10755), .B(n5827), .Y(CRC_OUT_1_3));
XOR2X1   g4962(.A(CRC_OUT_1_31), .B(WX11235), .Y(n10757));
XOR2X1   g4960(.A(CRC_OUT_1_2), .B(WX11237), .Y(n10755));
NOR2X1   g4959(.A(n10753), .B(n5827), .Y(CRC_OUT_1_2));
XOR2X1   g4958(.A(CRC_OUT_1_1), .B(WX11239), .Y(n10753));
NOR2X1   g4957(.A(n10751), .B(n5827), .Y(CRC_OUT_1_1));
XOR2X1   g4956(.A(CRC_OUT_1_0), .B(WX11241), .Y(n10751));

endmodule
