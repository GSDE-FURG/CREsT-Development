//Converted to Combinational (Partial output: g34237) , Module name: s38584_g34237 , Timestamp: 2018-12-03T15:51:18.317834 
module s38584_g34237 ( g53, g56, g57, g28, g19, g34, g54, g7, g31, g6, g8, g16, g9, g34237 );
input g53, g56, g57, g28, g19, g34, g54, g7, g31, g6, g8, g16, g9;
output g34237;
wire n5035, n5100, n5106_1, n5110, n5033, n5034, n5093, n5096_1, n5099, n5040, n5103, n5105, n5091_1, n5066_1, n5092, n4987, n5004, n5024, n4383, n5055, n5095, n5087, n5094, n5097, n5098, n5029, n5043, n5102, n5104, n4991, n5041, n5090, n5017_1, n5089, n4977, n4976, n4983, n4979_1, n5005, n5047_1, n5049, n5085, n5086_1, n5010, n5030, n5088, n5025, n5026, n5028, n5020, n5046, n4990, n4988_1, n5048, n5050, n4984_1, n5016, n5019, n5006, n5002_1, n4998, n4999, n5000, n5007_1, n5012_1, n5013, n5009, n5008, n5023, n5021, n5027_1, n4989, n4980, n4982, n4995, n5001, n4997_1, n5011, n5022_1, n4994, n4992_1, n4993, n4996;
NAND4X1  g0481(.A(n5110), .B(n5106_1), .C(n5100), .D(n5035), .Y(g34237));
NOR2X1   g0415(.A(n5034), .B(n5033), .Y(n5035));
NOR3X1   g0473(.A(n5099), .B(n5096_1), .C(n5093), .Y(n5100));
NOR3X1   g0478(.A(n5105), .B(n5103), .C(n5040), .Y(n5106_1));
AOI21X1  g0480(.A0(n5092), .A1(n5066_1), .B0(n5091_1), .Y(n5110));
NOR3X1   g0413(.A(n5024), .B(n5004), .C(n4987), .Y(n5033));
NOR2X1   g0414(.A(n4383), .B(g53), .Y(n5034));
AND2X1   g0466(.A(n5092), .B(n5055), .Y(n5093));
NOR4X1   g0469(.A(n5094), .B(n5091_1), .C(n5087), .D(n5095), .Y(n5096_1));
NOR3X1   g0472(.A(n5098), .B(n5097), .C(n5095), .Y(n5099));
NOR2X1   g0420(.A(n5029), .B(n4987), .Y(n5040));
NOR2X1   g0475(.A(n5102), .B(n5043), .Y(n5103));
NOR4X1   g0477(.A(n5041), .B(n5040), .C(n4991), .D(n5104), .Y(n5105));
INVX1    g0464(.A(n5090), .Y(n5091_1));
NOR3X1   g0443(.A(n5041), .B(n5040), .C(n5017_1), .Y(n5066_1));
NOR3X1   g0465(.A(n5091_1), .B(n5089), .C(n5087), .Y(n5092));
OR4X1    g0367(.A(n4976), .B(g57), .C(g56), .D(n4977), .Y(n4987));
NAND2X1  g0384(.A(n4983), .B(g28), .Y(n5004));
NAND3X1  g0404(.A(g19), .B(n5005), .C(n4979_1), .Y(n5024));
NOR4X1   g0358(.A(n4976), .B(g57), .C(g56), .D(n4977), .Y(n4383));
NOR4X1   g0435(.A(n5033), .B(n5040), .C(n5047_1), .D(n5034), .Y(n5055));
NAND3X1  g0468(.A(n5049), .B(n5017_1), .C(n4991), .Y(n5095));
AOI21X1  g0460(.A0(n5086_1), .A1(n5085), .B0(n4987), .Y(n5087));
NAND4X1  g0467(.A(n5029), .B(n5010), .C(n4383), .D(n5035), .Y(n5094));
NAND3X1  g0470(.A(n5087), .B(n5035), .C(n5030), .Y(n5097));
NAND2X1  g0471(.A(n5090), .B(n5088), .Y(n5098));
NOR3X1   g0409(.A(n5028), .B(n5026), .C(n5025), .Y(n5029));
NAND3X1  g0423(.A(n5035), .B(n5030), .C(n5020), .Y(n5043));
OR4X1    g0474(.A(n5087), .B(n5047_1), .C(n5046), .D(n5098), .Y(n5102));
OR4X1    g0476(.A(n5087), .B(n5020), .C(n5047_1), .D(n5098), .Y(n5104));
OR4X1    g0371(.A(n4988_1), .B(n4987), .C(g28), .D(n4990), .Y(n4991));
INVX1    g0421(.A(n5035), .Y(n5041));
NAND3X1  g0463(.A(n5050), .B(n5048), .C(n4383), .Y(n5090));
NAND3X1  g0397(.A(n5016), .B(n4984_1), .C(n4383), .Y(n5017_1));
NAND3X1  g0462(.A(n5088), .B(n5049), .C(n4991), .Y(n5089));
OR2X1    g0357(.A(g34), .B(g53), .Y(n4977));
INVX1    g0356(.A(g54), .Y(n4976));
NOR4X1   g0363(.A(g8), .B(g6), .C(g31), .D(g7), .Y(n4983));
INVX1    g0359(.A(g16), .Y(n4979_1));
INVX1    g0385(.A(g9), .Y(n5005));
NOR3X1   g0427(.A(n5006), .B(n5019), .C(n4987), .Y(n5047_1));
NAND3X1  g0429(.A(n5048), .B(n4984_1), .C(n4383), .Y(n5049));
NOR4X1   g0458(.A(n5000), .B(n4999), .C(n4998), .D(n5002_1), .Y(n5085));
NOR3X1   g0459(.A(n5013), .B(n5012_1), .C(n5007_1), .Y(n5086_1));
NOR4X1   g0390(.A(n5008), .B(g28), .C(n5005), .D(n5009), .Y(n5010));
OR2X1    g0410(.A(n5029), .B(n4987), .Y(n5030));
NAND2X1  g0461(.A(n5010), .B(n4383), .Y(n5088));
OAI21X1  g0405(.A0(n5024), .A1(n5021), .B0(n5023), .Y(n5025));
NOR4X1   g0406(.A(n5008), .B(g28), .C(g9), .D(n5009), .Y(n5026));
OAI21X1  g0408(.A0(n5024), .A1(n5019), .B0(n5027_1), .Y(n5028));
NOR3X1   g0400(.A(n4988_1), .B(n5019), .C(n4987), .Y(n5020));
NOR3X1   g0426(.A(n5021), .B(n4988_1), .C(n4987), .Y(n5046));
NAND2X1  g0370(.A(n4989), .B(g31), .Y(n4990));
NAND3X1  g0368(.A(g19), .B(g9), .C(n4979_1), .Y(n4988_1));
NOR3X1   g0428(.A(n4980), .B(n5005), .C(g16), .Y(n5048));
AND2X1   g0430(.A(n4983), .B(g28), .Y(n5050));
AND2X1   g0364(.A(n4983), .B(n4982), .Y(n4984_1));
NOR3X1   g0396(.A(g19), .B(g9), .C(n4979_1), .Y(n5016));
NAND2X1  g0399(.A(n4983), .B(n4982), .Y(n5019));
NAND3X1  g0386(.A(n4980), .B(n5005), .C(g16), .Y(n5006));
NOR3X1   g0382(.A(n5001), .B(n4995), .C(g28), .Y(n5002_1));
NOR3X1   g0378(.A(n4997_1), .B(n4995), .C(g28), .Y(n4998));
NOR3X1   g0379(.A(n4995), .B(n4988_1), .C(n4982), .Y(n4999));
NOR3X1   g0380(.A(n4997_1), .B(n4995), .C(n4982), .Y(n5000));
NOR2X1   g0387(.A(n5006), .B(n5004), .Y(n5007_1));
NOR2X1   g0392(.A(n5011), .B(n5006), .Y(n5012_1));
NOR4X1   g0393(.A(n5008), .B(n4982), .C(n5005), .D(n5009), .Y(n5013));
OR2X1    g0389(.A(g19), .B(g16), .Y(n5009));
OR4X1    g0388(.A(g8), .B(g6), .C(g31), .D(g7), .Y(n5008));
NAND4X1  g0403(.A(n4989), .B(g28), .C(g31), .D(n5022_1), .Y(n5023));
NAND3X1  g0401(.A(n4989), .B(n4982), .C(g31), .Y(n5021));
NAND3X1  g0407(.A(n5022_1), .B(n4983), .C(g28), .Y(n5027_1));
NOR3X1   g0369(.A(g7), .B(g8), .C(g6), .Y(n4989));
INVX1    g0360(.A(g19), .Y(n4980));
INVX1    g0362(.A(g28), .Y(n4982));
OR4X1    g0375(.A(n4993), .B(n4992_1), .C(g31), .D(n4994), .Y(n4995));
NAND3X1  g0381(.A(n4980), .B(g9), .C(g16), .Y(n5001));
NAND2X1  g0377(.A(n4996), .B(g9), .Y(n4997_1));
NAND3X1  g0391(.A(n4989), .B(g28), .C(g31), .Y(n5011));
NOR3X1   g0402(.A(g19), .B(g9), .C(g16), .Y(n5022_1));
INVX1    g0374(.A(g7), .Y(n4994));
INVX1    g0372(.A(g6), .Y(n4992_1));
INVX1    g0373(.A(g8), .Y(n4993));
NOR2X1   g0376(.A(g19), .B(g16), .Y(n4996));

endmodule
