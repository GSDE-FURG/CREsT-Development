//Converted to Combinational , Module name: s13207 , Timestamp: 2018-12-03T15:51:03.711215 
module s13207 ( g43, g49, g633, g634, g635, g645, g647, g648, g690, g694, g698, g702, g722, g723, g751, g752, g753, g754, g755, g756, g757, g781, g941, g962, g1000, g1008, g1016, g1080, g1234, g1553, g1554, g786, g1206, g929, g955, g795, g1194, g1198, g1202, g24, g1203, g1196, g29, g22, g28, g23, g37, g26, g27, g42, g32, g41, g31, g45, g44, g21, g30, g25, g397, g1271, g312, g273, g452, g948, g629, g207, g1541, g1153, g940, g976, g498, g314, g1092, g454, g196, g535, g292, g772, g1375, g689, g183, g359, g1384, g1339, g1424, g767, g393, g1077, g1231, g294, g1477, g608, g465, g774, g921, g1304, g243, g1499, g80, g1444, g1269, g600, g423, g771, g803, g843, g315, g455, g906, g622, g891, g1014, g984, g117, g527, g1513, g278, g1378, g718, g598, g1182, g1288, g1382, g179, g624, g48, g362, g878, g270, g763, g710, g730, g295, g1037, g1102, g483, g775, g621, g1364, g1454, g1296, g1532, g587, g741, g606, g1012, g646, g1412, g327, g1189, g1389, g1029, g1371, g1429, g398, g985, g354, g619, g113, g180, g1138, g1309, g889, g390, g625, g417, g681, g437, g351, g1049, g1098, g200, g240, g479, g596, g1268, g222, g420, g172, g387, g840, g365, g1486, g1504, g1185, g1385, g583, g822, g1025, g969, g768, g174, g685, g1087, g355, g911, g1226, g99, g1045, g1173, g1373, g186, g760, g959, g1369, g1007, g1459, g758, g480, g396, g612, g632, g1415, g1227, g246, g449, g517, g16, g284, g219, g426, g1388, g806, g846, g1428, g579, g1030, g614, g1430, g1247, g669, g225, g281, g819, g1308, g611, g631, g1217, g1365, g825, g1333, g474, g1396, g1509, g766, g1018, g588, g1467, g317, g457, g486, g471, g1381, g513, g1397, g533, g1021, g1421, g952, g1263, g580, g615, g1257, g402, g998, g1041, g297, g954, g105, g212, g1368, g232, g990, g475, g33, g951, g799, g812, g567, g313, g333, g168, g214, g234, g652, g1126, g1400, g1326, g309, g211, g834, g231, g557, g1383, g1220, g158, g627, g661, g831, g1327, g293, g1146, g773, g859, g1240, g518, g1472, g1443, g436, g405, g1034, g1147, g374, g563, g510, g530, g215, g235, g1013, g1317, g504, g665, g544, g371, g792, g468, g815, g1460, g553, g623, g501, g1190, g1390, g1156, g318, g458, g342, g1250, g1163, g1363, g1432, g1053, g252, g330, g264, g1157, g1357, g375, g852, g261, g516, g536, g979, g778, g199, g1292, g290, g1084, g1439, g770, g1276, g890, g1004, g1404, g93, g287, g560, g1224, g1320, g617, g316, g336, g933, g456, g345, g628, g887, g789, g173, g550, g255, g949, g1244, g620, g1435, g477, g926, g368, g855, g1214, g1110, g1310, g296, g972, g1402, g1236, g896, g613, g566, g1394, g1489, g883, g971, g609, g1254, g556, g1409, g626, g1229, g782, g237, g942, g228, g706, g746, g1462, g963, g837, g599, g1192, g828, g1392, g492, g944, g195, g1431, g1252, g356, g953, g1176, g1376, g1005, g1405, g901, g1270, g1225, g1073, g1324, g1069, g443, g1377, g377, g618, g602, g213, g233, g1199, g1399, g888, g573, g399, g1245, g507, g547, g610, g630, g1207, g249, g916, g936, g478, g604, g945, g1114, g429, g809, g849, g1408, g1336, g601, g1065, g1122, g1228, g495, g1322, g1230, g1033, g267, g1395, g373, g274, g1266, g714, g734, g1142, g1342, g769, g1081, g1481, g1097, g543, g1154, g1354, g489, g874, g591, g616, g1267, g1312, g605, g182, g1401, g950, g1329, g408, g871, g759, g202, g440, g476, g184, g1149, g1398, g210, g394, g86, g570, g275, g303, g181, g1524, g595, g1319, g863, g1211, g966, g1186, g1386, g875, g1170, g1370, g201, g1325, g1280, g1106, g1061, g1387, g762, g1461, g378, g1200, g1514, g1403, g1345, g1191, g1391, g185, g1307, g1159, g1223, g446, g1416, g395, g764, g1251, g216, g236, g205, g540, g576, g1537, g727, g999, g761, g1272, g1243, g1328, g1130, g1330, g1166, g524, g1366, g348, g1148, g1348, g1155, g1260, g258, g521, g300, g765, g1118, g1167, g1318, g1367, g677, g376, g1057, g973, g1393, g1549, g1321, g1253, g1519, g584, g539, g324, g432, g1158, g321, g1311, g414, g1374, g1284, g1545, g1380, g673, g607, g306, g943, g162, g411, g866, g1204, g1300, g384, g339, g459, g1323, g381, g1528, g1351, g597, g1372, g435, g970, g1134, g995, g190, g1313, g603, g1494, g462, g1160, g1360, g1450, g187, g1179, g1379, g206, g291, g372, g453, g534, g594, g785, g1006, g1015, g1017, g1246, g1724, g1783, g1798, g1804, g1810, g1817, g1824, g1829, g1870, g1871, g1894, g1911, g1944, g2662, g2844, g2888, g3077, g3096, g3130, g3159, g3191, g3829, g3859, g3860, g4267, g4316, g4370, g4371, g4372, g4373, g4655, g4657, g4660, g4661, g4663, g4664, g5143, g5164, g5571, g5669, g5678, g5682, g5684, g5687, g5729, g6207, g6212, g6223, g6236, g6269, g6425, g6648, g6653, g6675, g6849, g6850, g6895, g6909, g7048, g7063, g7103, g7283, g7284, g7285, g7286, g7287, g7288, g7289, g7290, g7291, g7292, g7293, g7294, g7295, g7298, g7423, g7424, g7425, g7474, g7504, g7505, g7506, g7507, g7508, g7514, g7729, g7730, g7731, g7732, g8216, g8217, g8218, g8219, g8234, g8661, g8663, g8872, g8958, g9128, g9132, g9204, g9280, g9297, g9299, g9305, g9308, g9310, g9312, g9314, g9378, g7763, g1205, g3856, g3857, g3854, g1193, g1197, g1201, g6294, g6376, g1195, g6300, g6292, g6298, g6291, g6293, g6304, g6296, g6289, g6297, g6306, g6290, g6303, g6305, g6302, g6308, g6288, g6307, g6299, g6301, g6295, n429, n434, n439, n444, n449, n454, n459, n464, n469, n474, n479, n484, n489, n494, n499, n504, n509, n514, n519, n524, n529, n534, n539, n544, n549, n554, n559, n564, n569, n574, n579, n584, n589, n594, n599, n604, n613, n618, n623, n628, n633, n638, n643, n648, n653, n658, n663, n668, n673, n678, n683, n688, n693, n698, n703, n708, n713, n718, n723, n728, n733, n738, n743, n748, n753, n758, n763, n768, n773, n778, n783, n788, n793, n798, n803, n808, n813, n818, n823, n828, n833, n838, n843, n848, n853, n858, n863, n868, n873, n878, n883, n888, n893, n897, n902, n907, n912, n917, n922, n927, n932, n937, n942, n947, n952, n957, n962, n967, n972, n977, n982, n987, n992, n997, n1002, n1007, n1012, n1017, n1026, n1031, n1036, n1041, n1046, n1051, n1056, n1061, n1066, n1071, n1076, n1081, n1086, n1091, n1096, n1101, n1106, n1111, n1116, n1121, n1126, n1131, n1136, n1141, n1146, n1151, n1156, n1161, n1166, n1171, n1175, n1180, n1185, n1190, n1195, n1200, n1205, n1210, n1215, n1220, n1225, n1230, n1235, n1240, n1245, n1250, n1255, n1260, n1265, n1270, n1275, n1280, n1284, n1289, n1294, n1299, n1304, n1309, n1314, n1319, n1324, n1329, n1334, n1339, n1344, n1349, n1354, n1359, n1364, n1369, n1373, n1378, n1383, n1388, n1393, n1398, n1402, n1407, n1412, n1417, n1422, n1427, n1432, n1437, n1442, n1447, n1452, n1457, n1462, n1467, n1472, n1477, n1482, n1487, n1492, n1497, n1505, n1510, n1515, n1520, n1525, n1530, n1535, n1540, n1545, n1550, n1555, n1560, n1565, n1570, n1575, n1580, n1584, n1589, n1594, n1599, n1604, n1609, n1614, n1619, n1624, n1629, n1634, n1639, n1644, n1649, n1654, n1659, n1664, n1668, n1673, n1678, n1683, n1688, n1693, n1698, n1703, n1708, n1713, n1718, n1723, n1728, n1733, n1738, n1743, n1748, n1753, n1758, n1763, n1767, n1772, n1777, n1782, n1787, n1792, n1797, n1802, n1807, n1812, n1817, n1821, n1826, n1831, n1836, n1841, n1846, n1850, n1855, n1859, n1864, n1869, n1874, n1879, n1884, n1889, n1894, n1899, n1904, n1909, n1914, n1919, n1924, n1929, n1934, n1939, n1944, n1949, n1954, n1959, n1964, n1969, n1974, n1979, n1984, n1989, n1994, n1999, n2004, n2009, n2013, n2018, n2023, n2028, n2033, n2038, n2043, n2048, n2053, n2058, n2063, n2067, n2072, n2077, n2082, n2087, n2092, n2097, n2101, n2106, n2110, n2115, n2120, n2124, n2129, n2134, n2139, n2144, n2149, n2154, n2159, n2164, n2169, n2174, n2179, n2184, n2189, n2194, n2199, n2204, n2209, n2214, n2219, n2224, n2228, n2233, n2237, n2242, n2247, n2251, n2256, n2261, n2266, n2270, n2273, n2278, n2283, n2288, n2293, n2297, n2302, n2307, n2312, n2317, n2322, n2327, n2332, n2337, n2342, n2347, n2352, n2357, n2362, n2367, n2372, n2377, n2382, n2387, n2392, n2397, n2402, n2407, n2412, n2417, n2422, n2427, n2432, n2437, n2442, n2447, n2452, n2457, n2462, n2466, n2470, n2474, n2477, n2481, n2486, n2491, n2496, n2501, n2506, n2511, n2516, n2521, n2526, n2531, n2536, n2541, n2546, n2551, n2556, n2561, n2565, n2570, n2575, n2580, n2585, n2590, n2595, n2600, n2605, n2609, n2613, n2618, n2623, n2628, n2633, n2637, n2642, n2647, n2652, n2657, n2662, n2667, n2672, n2677, n2682, n2687, n2692, n2697, n2702, n2707, n2712, n2721, n2726, n2731, n2736, n2741, n2746, n2751, n2756, n2761, n2766, n2770, n2774, n2779, n2783, n2788, n2793, n2798, n2803, n2808, n2813, n2818, n2823, n2827, n2832, n2836, n2841, n2846, n2851, n2856, n2861, n2866, n2871, n2876, n2881, n2886, n2891, n2895, n2900, n2905, n2910, n2915, n2920, n2925, n2930, n2935, n2940, n2944, n2949, n2954, n2959, n2964, n2967, n2972, n2977, n2981, n2986, n2990, n2995, n3000, n3005, n3010, n3015, n3020, n3025, n3030, n3034, n3038, n3042, n3046, n3051, n3054, n3059, n3064, n3068, n3073, n3078, n3083, n3088, n3093, n3098, n3103, n3108, n3113, n3118, n3123, n3127, n3132, n3137, n3142, n3147, n3152, n3157, n3162, n3167, n3172, n3177, n3182, n3187, n3192, n3197, n3201, n3206, n3210, n3214, n3219, n3224, n3229, n3234, n3239, n3244, n3248, n3252, n3257, n3262, n3267, n3272, n3277, n3285, n3289, n3294, n3299, n3304, n3309, n3314, n3319, n3324, n3328, n3333, n3337, n3341, n3346, n3351, n3355, n3360, n3365, n3370, n3375, n3380, n3385, n3390, n3395, n3400, n3404, n3408, n3413, n3418, n3423, n3428, n3433, n3438, n3443, n3448, n3453, n3458, n3463, n3467, n3472, n3477, n3481, n3486, n3491, n3496, n3501, n3505, n3509, n3514, n3519, n3523, n3528, n3533, n3538 );
input g94, g92, g104, g109, g9, g20, g145, g125, g137, g108, g133, g121, g129, g12, g11, g141, g98, g103, g38, g46, g13, g47, g146, g114, g118, g150, g122, g126, g89, g154, g130, g95, g134, g100, g138, g142, g110, g55, g10, g62, g65, g8, g3, g2, g4, g5, g6, g58, g7, g71, g77, g74, g68, g52, g83, g1, g43, g49, g633, g634, g635, g645, g647, g648, g690, g694, g698, g702, g722, g723, g751, g752, g753, g754, g755, g756, g757, g781, g941, g962, g1000, g1008, g1016, g1080, g1234, g1553, g1554, g786, g1206, g929, g955, g795, g1194, g1198, g1202, g24, g1203, g1196, g29, g22, g28, g23, g37, g26, g27, g42, g32, g41, g31, g45, g44, g21, g30, g25, g397, g1271, g312, g273, g452, g948, g629, g207, g1541, g1153, g940, g976, g498, g314, g1092, g454, g196, g535, g292, g772, g1375, g689, g183, g359, g1384, g1339, g1424, g767, g393, g1077, g1231, g294, g1477, g608, g465, g774, g921, g1304, g243, g1499, g80, g1444, g1269, g600, g423, g771, g803, g843, g315, g455, g906, g622, g891, g1014, g984, g117, g527, g1513, g278, g1378, g718, g598, g1182, g1288, g1382, g179, g624, g48, g362, g878, g270, g763, g710, g730, g295, g1037, g1102, g483, g775, g621, g1364, g1454, g1296, g1532, g587, g741, g606, g1012, g646, g1412, g327, g1189, g1389, g1029, g1371, g1429, g398, g985, g354, g619, g113, g180, g1138, g1309, g889, g390, g625, g417, g681, g437, g351, g1049, g1098, g200, g240, g479, g596, g1268, g222, g420, g172, g387, g840, g365, g1486, g1504, g1185, g1385, g583, g822, g1025, g969, g768, g174, g685, g1087, g355, g911, g1226, g99, g1045, g1173, g1373, g186, g760, g959, g1369, g1007, g1459, g758, g480, g396, g612, g632, g1415, g1227, g246, g449, g517, g16, g284, g219, g426, g1388, g806, g846, g1428, g579, g1030, g614, g1430, g1247, g669, g225, g281, g819, g1308, g611, g631, g1217, g1365, g825, g1333, g474, g1396, g1509, g766, g1018, g588, g1467, g317, g457, g486, g471, g1381, g513, g1397, g533, g1021, g1421, g952, g1263, g580, g615, g1257, g402, g998, g1041, g297, g954, g105, g212, g1368, g232, g990, g475, g33, g951, g799, g812, g567, g313, g333, g168, g214, g234, g652, g1126, g1400, g1326, g309, g211, g834, g231, g557, g1383, g1220, g158, g627, g661, g831, g1327, g293, g1146, g773, g859, g1240, g518, g1472, g1443, g436, g405, g1034, g1147, g374, g563, g510, g530, g215, g235, g1013, g1317, g504, g665, g544, g371, g792, g468, g815, g1460, g553, g623, g501, g1190, g1390, g1156, g318, g458, g342, g1250, g1163, g1363, g1432, g1053, g252, g330, g264, g1157, g1357, g375, g852, g261, g516, g536, g979, g778, g199, g1292, g290, g1084, g1439, g770, g1276, g890, g1004, g1404, g93, g287, g560, g1224, g1320, g617, g316, g336, g933, g456, g345, g628, g887, g789, g173, g550, g255, g949, g1244, g620, g1435, g477, g926, g368, g855, g1214, g1110, g1310, g296, g972, g1402, g1236, g896, g613, g566, g1394, g1489, g883, g971, g609, g1254, g556, g1409, g626, g1229, g782, g237, g942, g228, g706, g746, g1462, g963, g837, g599, g1192, g828, g1392, g492, g944, g195, g1431, g1252, g356, g953, g1176, g1376, g1005, g1405, g901, g1270, g1225, g1073, g1324, g1069, g443, g1377, g377, g618, g602, g213, g233, g1199, g1399, g888, g573, g399, g1245, g507, g547, g610, g630, g1207, g249, g916, g936, g478, g604, g945, g1114, g429, g809, g849, g1408, g1336, g601, g1065, g1122, g1228, g495, g1322, g1230, g1033, g267, g1395, g373, g274, g1266, g714, g734, g1142, g1342, g769, g1081, g1481, g1097, g543, g1154, g1354, g489, g874, g591, g616, g1267, g1312, g605, g182, g1401, g950, g1329, g408, g871, g759, g202, g440, g476, g184, g1149, g1398, g210, g394, g86, g570, g275, g303, g181, g1524, g595, g1319, g863, g1211, g966, g1186, g1386, g875, g1170, g1370, g201, g1325, g1280, g1106, g1061, g1387, g762, g1461, g378, g1200, g1514, g1403, g1345, g1191, g1391, g185, g1307, g1159, g1223, g446, g1416, g395, g764, g1251, g216, g236, g205, g540, g576, g1537, g727, g999, g761, g1272, g1243, g1328, g1130, g1330, g1166, g524, g1366, g348, g1148, g1348, g1155, g1260, g258, g521, g300, g765, g1118, g1167, g1318, g1367, g677, g376, g1057, g973, g1393, g1549, g1321, g1253, g1519, g584, g539, g324, g432, g1158, g321, g1311, g414, g1374, g1284, g1545, g1380, g673, g607, g306, g943, g162, g411, g866, g1204, g1300, g384, g339, g459, g1323, g381, g1528, g1351, g597, g1372, g435, g970, g1134, g995, g190, g1313, g603, g1494, g462, g1160, g1360, g1450, g187, g1179, g1379;
output g206, g291, g372, g453, g534, g594, g785, g1006, g1015, g1017, g1246, g1724, g1783, g1798, g1804, g1810, g1817, g1824, g1829, g1870, g1871, g1894, g1911, g1944, g2662, g2844, g2888, g3077, g3096, g3130, g3159, g3191, g3829, g3859, g3860, g4267, g4316, g4370, g4371, g4372, g4373, g4655, g4657, g4660, g4661, g4663, g4664, g5143, g5164, g5571, g5669, g5678, g5682, g5684, g5687, g5729, g6207, g6212, g6223, g6236, g6269, g6425, g6648, g6653, g6675, g6849, g6850, g6895, g6909, g7048, g7063, g7103, g7283, g7284, g7285, g7286, g7287, g7288, g7289, g7290, g7291, g7292, g7293, g7294, g7295, g7298, g7423, g7424, g7425, g7474, g7504, g7505, g7506, g7507, g7508, g7514, g7729, g7730, g7731, g7732, g8216, g8217, g8218, g8219, g8234, g8661, g8663, g8872, g8958, g9128, g9132, g9204, g9280, g9297, g9299, g9305, g9308, g9310, g9312, g9314, g9378, g7763, g1205, g3856, g3857, g3854, g1193, g1197, g1201, g6294, g6376, g1195, g6300, g6292, g6298, g6291, g6293, g6304, g6296, g6289, g6297, g6306, g6290, g6303, g6305, g6302, g6308, g6288, g6307, g6299, g6301, g6295, n429, n434, n439, n444, n449, n454, n459, n464, n469, n474, n479, n484, n489, n494, n499, n504, n509, n514, n519, n524, n529, n534, n539, n544, n549, n554, n559, n564, n569, n574, n579, n584, n589, n594, n599, n604, n613, n618, n623, n628, n633, n638, n643, n648, n653, n658, n663, n668, n673, n678, n683, n688, n693, n698, n703, n708, n713, n718, n723, n728, n733, n738, n743, n748, n753, n758, n763, n768, n773, n778, n783, n788, n793, n798, n803, n808, n813, n818, n823, n828, n833, n838, n843, n848, n853, n858, n863, n868, n873, n878, n883, n888, n893, n897, n902, n907, n912, n917, n922, n927, n932, n937, n942, n947, n952, n957, n962, n967, n972, n977, n982, n987, n992, n997, n1002, n1007, n1012, n1017, n1026, n1031, n1036, n1041, n1046, n1051, n1056, n1061, n1066, n1071, n1076, n1081, n1086, n1091, n1096, n1101, n1106, n1111, n1116, n1121, n1126, n1131, n1136, n1141, n1146, n1151, n1156, n1161, n1166, n1171, n1175, n1180, n1185, n1190, n1195, n1200, n1205, n1210, n1215, n1220, n1225, n1230, n1235, n1240, n1245, n1250, n1255, n1260, n1265, n1270, n1275, n1280, n1284, n1289, n1294, n1299, n1304, n1309, n1314, n1319, n1324, n1329, n1334, n1339, n1344, n1349, n1354, n1359, n1364, n1369, n1373, n1378, n1383, n1388, n1393, n1398, n1402, n1407, n1412, n1417, n1422, n1427, n1432, n1437, n1442, n1447, n1452, n1457, n1462, n1467, n1472, n1477, n1482, n1487, n1492, n1497, n1505, n1510, n1515, n1520, n1525, n1530, n1535, n1540, n1545, n1550, n1555, n1560, n1565, n1570, n1575, n1580, n1584, n1589, n1594, n1599, n1604, n1609, n1614, n1619, n1624, n1629, n1634, n1639, n1644, n1649, n1654, n1659, n1664, n1668, n1673, n1678, n1683, n1688, n1693, n1698, n1703, n1708, n1713, n1718, n1723, n1728, n1733, n1738, n1743, n1748, n1753, n1758, n1763, n1767, n1772, n1777, n1782, n1787, n1792, n1797, n1802, n1807, n1812, n1817, n1821, n1826, n1831, n1836, n1841, n1846, n1850, n1855, n1859, n1864, n1869, n1874, n1879, n1884, n1889, n1894, n1899, n1904, n1909, n1914, n1919, n1924, n1929, n1934, n1939, n1944, n1949, n1954, n1959, n1964, n1969, n1974, n1979, n1984, n1989, n1994, n1999, n2004, n2009, n2013, n2018, n2023, n2028, n2033, n2038, n2043, n2048, n2053, n2058, n2063, n2067, n2072, n2077, n2082, n2087, n2092, n2097, n2101, n2106, n2110, n2115, n2120, n2124, n2129, n2134, n2139, n2144, n2149, n2154, n2159, n2164, n2169, n2174, n2179, n2184, n2189, n2194, n2199, n2204, n2209, n2214, n2219, n2224, n2228, n2233, n2237, n2242, n2247, n2251, n2256, n2261, n2266, n2270, n2273, n2278, n2283, n2288, n2293, n2297, n2302, n2307, n2312, n2317, n2322, n2327, n2332, n2337, n2342, n2347, n2352, n2357, n2362, n2367, n2372, n2377, n2382, n2387, n2392, n2397, n2402, n2407, n2412, n2417, n2422, n2427, n2432, n2437, n2442, n2447, n2452, n2457, n2462, n2466, n2470, n2474, n2477, n2481, n2486, n2491, n2496, n2501, n2506, n2511, n2516, n2521, n2526, n2531, n2536, n2541, n2546, n2551, n2556, n2561, n2565, n2570, n2575, n2580, n2585, n2590, n2595, n2600, n2605, n2609, n2613, n2618, n2623, n2628, n2633, n2637, n2642, n2647, n2652, n2657, n2662, n2667, n2672, n2677, n2682, n2687, n2692, n2697, n2702, n2707, n2712, n2721, n2726, n2731, n2736, n2741, n2746, n2751, n2756, n2761, n2766, n2770, n2774, n2779, n2783, n2788, n2793, n2798, n2803, n2808, n2813, n2818, n2823, n2827, n2832, n2836, n2841, n2846, n2851, n2856, n2861, n2866, n2871, n2876, n2881, n2886, n2891, n2895, n2900, n2905, n2910, n2915, n2920, n2925, n2930, n2935, n2940, n2944, n2949, n2954, n2959, n2964, n2967, n2972, n2977, n2981, n2986, n2990, n2995, n3000, n3005, n3010, n3015, n3020, n3025, n3030, n3034, n3038, n3042, n3046, n3051, n3054, n3059, n3064, n3068, n3073, n3078, n3083, n3088, n3093, n3098, n3103, n3108, n3113, n3118, n3123, n3127, n3132, n3137, n3142, n3147, n3152, n3157, n3162, n3167, n3172, n3177, n3182, n3187, n3192, n3197, n3201, n3206, n3210, n3214, n3219, n3224, n3229, n3234, n3239, n3244, n3248, n3252, n3257, n3262, n3267, n3272, n3277, n3285, n3289, n3294, n3299, n3304, n3309, n3314, n3319, n3324, n3328, n3333, n3337, n3341, n3346, n3351, n3355, n3360, n3365, n3370, n3375, n3380, n3385, n3390, n3395, n3400, n3404, n3408, n3413, n3418, n3423, n3428, n3433, n3438, n3443, n3448, n3453, n3458, n3463, n3467, n3472, n3477, n3481, n3486, n3491, n3496, n3501, n3505, n3509, n3514, n3519, n3523, n3528, n3533, n3538;
wire n2129_1, n2130, n2131, n2132, n2133, n2134_1, n2135, n2139_1, n2142, n2143, n2144_1, n2145, n2147, n2148, n2150, n2151, n2153, n2154_1, n2155, n2157, n2159_1, n2161, n2163, n2165, n2166, n2167, n2172, n2173, n2174_1, n2175, n2176, n2177, n2178, n2179_1, n2180, n2181, n2182, n2185, n2188, n2189_1, n2190, n2191, n2200, n2204_1, n2205, n2206, n2208, n2211, n2212, n2215, n2216, n2217, n2218, n2219_1, n2220, n2222, n2223, n2226, n2227, n2229, n2230, n2231, n2232, n2233_1, n2234, n2235, n2236, n2237_1, n2238, n2239, n2240, n2241, n2242_1, n2243, n2244, n2245, n2246, n2247_1, n2248, n2249, n2250, n2251_1, n2252, n2253, n2254, n2255, n2256_1, n2257, n2258, n2259, n2260, n2261_1, n2262, n2263, n2264, n2265, n2266_1, n2267, n2268, n2269, n2270_1, n2271, n2272, n2273_1, n2274, n2275, n2276, n2277, n2278_1, n2279, n2280, n2281, n2282, n2283_1, n2284, n2285, n2286, n2287, n2288_1, n2289, n2290, n2291, n2292, n2293_1, n2294, n2295, n2296, n2297_1, n2298, n2299, n2300, n2301, n2302_1, n2303, n2304, n2305, n2306, n2307_1, n2308, n2309, n2310, n2311, n2312_1, n2313, n2314, n2315, n2316, n2317_1, n2318, n2319, n2320, n2321, n2322_1, n2323, n2324, n2325, n2326, n2327_1, n2328, n2329, n2330, n2331, n2332_1, n2333, n2334, n2335, n2336, n2337_1, n2338, n2339, n2340, n2341, n2342_1, n2343, n2344, n2345, n2346, n2347_1, n2348, n2349, n2350, n2351, n2352_1, n2353, n2354, n2355, n2356, n2357_1, n2358, n2359, n2360, n2361, n2362_1, n2363, n2364, n2365, n2366, n2367_1, n2368, n2369, n2370, n2371, n2372_1, n2373, n2374, n2375, n2376, n2377_1, n2378, n2379, n2380, n2381, n2382_1, n2384, n2385, n2386, n2387_1, n2388, n2389, n2390, n2391, n2392_1, n2393, n2394, n2395, n2398, n2399, n2400, n2401, n2402_1, n2403, n2404, n2405, n2406, n2407_1, n2408, n2409, n2410, n2411, n2412_1, n2413, n2414, n2415, n2416, n2417_1, n2418, n2419, n2420, n2421, n2422_1, n2423, n2424, n2425, n2426, n2427_1, n2428, n2429, n2430, n2431, n2432_1, n2434, n2435, n2436, n2437_1, n2438, n2439, n2440, n2441, n2442_1, n2443, n2444, n2445, n2446, n2447_1, n2448, n2449, n2450, n2451, n2452_1, n2453, n2454, n2455, n2456, n2457_1, n2458, n2459, n2460, n2461, n2462_1, n2463, n2464, n2466_1, n2467, n2468, n2469, n2470_1, n2471, n2472, n2473, n2474_1, n2475, n2476, n2477_1, n2478, n2479, n2480, n2481_1, n2482, n2483, n2484, n2485, n2486_1, n2487, n2488, n2489, n2490, n2491_1, n2492, n2493, n2494, n2496_1, n2497, n2498, n2499, n2500, n2501_1, n2502, n2503, n2504, n2505, n2506_1, n2507, n2508, n2509, n2510, n2511_1, n2512, n2513, n2514, n2515, n2516_1, n2517, n2518, n2519, n2520, n2521_1, n2522, n2523, n2524, n2525, n2526_1, n2527, n2529, n2530, n2531_1, n2532, n2533, n2534, n2535, n2536_1, n2537, n2538, n2539, n2540, n2541_1, n2542, n2543, n2544, n2545, n2546_1, n2547, n2548, n2549, n2550, n2551_1, n2552, n2553, n2555, n2556_1, n2557, n2558, n2559, n2560, n2561_1, n2562, n2563, n2564, n2565_1, n2566, n2567, n2568, n2569, n2570_1, n2571, n2572, n2573, n2574, n2575_1, n2576, n2577, n2578, n2579, n2580_1, n2582, n2583, n2584, n2585_1, n2586, n2587, n2588, n2589, n2590_1, n2591, n2592, n2593, n2594, n2595_1, n2596, n2597, n2598, n2599, n2600_1, n2601, n2602, n2603, n2604, n2606, n2607, n2608, n2609_1, n2610, n2611, n2612, n2613_1, n2615, n2616, n2617, n2618_1, n2619, n2620, n2621, n2622, n2623_1, n2625, n2626, n2627, n2632, n2634, n2635, n2636, n2638, n2639, n2640, n2641, n2643, n2644, n2645, n2646, n2647_1, n2648, n2649, n2650, n2651, n2652_1, n2654, n2655, n2658, n2662_1, n2664, n2665, n2667_1, n2668, n2669, n2672_1, n2673, n2674, n2675, n2676, n2677_1, n2678, n2679, n2680, n2682_1, n2683, n2686, n2687_1, n2688, n2690, n2691, n2692_1, n2693, n2694, n2695, n2696, n2697_1, n2698, n2699, n2700, n2701, n2702_1, n2703, n2706, n2707_1, n2708, n2709, n2710, n2711, n2712_1, n2714, n2716, n2717_1, n2718, n2719, n2720, n2721_1, n2722, n2723, n2724, n2725, n2726_1, n2727, n2728, n2729, n2730, n2731_1, n2732, n2733, n2734, n2735, n2736_1, n2737, n2738, n2739, n2740, n2741_1, n2742, n2743, n2744, n2745, n2746_1, n2748, n2749, n2751_1, n2752, n2754, n2755, n2757, n2758, n2759, n2761_1, n2763, n2764, n2767, n2768, n2769, n2770_1, n2771, n2772, n2778, n2780, n2781, n2782, n2783_1, n2784, n2785, n2786, n2789, n2790, n2796, n2797, n2798_1, n2799, n2800, n2801, n2803_1, n2804, n2805, n2806, n2809, n2812, n2813_1, n2815, n2816, n2817, n2818_1, n2820, n2821, n2822, n2824, n2825, n2827_1, n2829, n2830, n2831, n2832_1, n2834, n2835, n2836_1, n2837, n2838, n2839, n2840, n2841_1, n2842, n2843, n2845, n2848, n2849, n2850, n2851_1, n2852, n2853, n2854, n2855, n2856_1, n2857, n2859, n2860, n2861_1, n2864, n2865, n2866_1, n2868, n2869, n2870, n2871_1, n2873, n2874, n2875, n2876_1, n2878, n2879, n2880, n2881_1, n2882, n2883, n2884, n2885, n2886_1, n2887, n2888, n2890, n2891_1, n2894, n2898, n2899, n2900_1, n2901, n2902, n2903, n2905_1, n2906, n2909, n2910_1, n2914, n2915_1, n2917, n2918, n2921, n2923, n2925_1, n2926, n2929, n2930_1, n2931, n2933, n2934, n2935_1, n2936, n2937, n2938, n2940_1, n2943, n2945, n2946, n2947, n2948, n2949_1, n2950, n2952, n2953, n2954_1, n2959_1, n2962, n2963, n2964_1, n2965, n2966, n2967_1, n2970, n2971, n2972_1, n2975, n2980, n2981_1, n2985, n2986_1, n2987, n2988, n2993, n2994, n2997, n2998, n2999, n3000_1, n3003, n3004, n3006, n3008, n3009, n3010_1, n3012, n3013, n3014, n3017, n3018, n3019, n3025_1, n3027, n3030_1, n3032, n3033, n3035, n3037, n3038_1, n3041, n3042_1, n3043, n3048, n3050, n3053, n3055, n3060, n3061, n3063, n3064_1, n3065, n3066, n3071, n3072, n3073_1, n3077, n3078_1, n3079, n3080, n3083_1, n3086, n3087, n3088_1, n3091, n3092, n3093_1, n3097, n3098_1, n3100, n3108_1, n3112, n3113_1, n3114, n3115, n3116, n3117, n3118_1, n3119, n3120, n3124, n3125, n3129, n3130, n3132_1, n3133, n3134, n3135, n3140, n3141, n3148, n3149, n3150, n3152_1, n3153, n3155, n3157_1, n3158, n3162_1, n3163, n3166, n3167_1, n3168, n3169, n3171, n3172_1, n3173, n3178, n3179, n3181, n3182_1, n3183, n3184, n3185, n3186, n3187_1, n3188, n3197_1, n3198, n3199, n3201_1, n3202, n3204, n3205, n3206_1, n3207, n3208, n3209, n3210_1, n3211, n3212, n3213, n3214_1, n3215, n3216, n3217, n3218, n3219_1, n3220, n3221, n3222, n3224_1, n3225, n3227, n3228, n3232, n3233, n3234_1, n3236, n3241, n3242, n3243, n3245, n3246, n3248_1, n3254, n3255, n3258, n3260, n3261, n3262_1, n3263, n3264, n3266, n3267_1, n3268, n3269, n3270, n3271, n3272_1, n3274, n3275, n3277_1, n3278, n3279, n3280, n3284, n3285_1, n3286, n3287, n3296, n3299_1, n3300, n3301, n3304_1, n3305, n3308, n3309_1, n3311, n3312, n3314_1, n3315, n3317, n3318, n3321, n3322, n3323, n3324_1, n3325, n3327, n3328_1, n3329, n3331, n3337_1, n3338, n3340, n3342, n3344, n3346_1, n3355_1, n3356, n3357, n3360_1, n3361, n3366, n3367, n3369, n3371, n3376, n3377, n3378, n3380_1, n3381, n3382, n3384, n3385_1, n3386, n3387, n3389, n3390_1, n3393, n3394, n3397, n3398, n3399, n3401, n3402, n3404_1, n3405, n3408_1, n3412, n3413_1, n3414, n3418_1, n3420, n3421, n3422, n3424, n3425, n3426, n3432, n3433_1, n3434, n3437, n3438_1, n3443_1, n3444, n3445, n3447, n3448_1, n3452, n3453_1, n3454, n3457, n3458_1, n3459, n3461, n3462, n3465, n3466, n3474, n3475, n3476, n3477_1, n3479, n3480, n3489, n3490, n3491_1, n3496_1, n3497, n3500, n3501_1, n3503, n3504, n3507, n3509_1, n3510, n3511, n3513, n3514_1, n3515, n3518, n3519_1, n3522, n3523_1, n3525, n3527, n3528_1, n3529;
INVX1    g0000(.A(g43), .Y(g6850));
INVX1    g0001(.A(g162), .Y(n2129_1));
NOR4X1   g0002(.A(g971), .B(g972), .C(g962), .D(g963), .Y(n2130));
INVX1    g0003(.A(n2130), .Y(n2131));
NOR4X1   g0004(.A(g970), .B(g966), .C(g969), .D(n2131), .Y(n2132));
INVX1    g0005(.A(n2132), .Y(n2133));
INVX1    g0006(.A(g973), .Y(n2134_1));
INVX1    g0007(.A(g1), .Y(n2135));
NOR2X1   g0008(.A(n2132), .B(n2135), .Y(g7298));
NOR2X1   g0009(.A(n2132), .B(g1), .Y(g7103));
NOR4X1   g0010(.A(g7298), .B(n2134_1), .C(g6850), .D(g7103), .Y(n2964));
OAI21X1  g0011(.A0(n2132), .A1(n2135), .B0(g976), .Y(n2139_1));
NOR3X1   g0012(.A(n2139_1), .B(g7103), .C(g6850), .Y(n2382));
INVX1    g0013(.A(g1034), .Y(n2307));
INVX1    g0014(.A(g979), .Y(n2142));
NAND3X1  g0015(.A(n2142), .B(g984), .C(g43), .Y(n2143));
NAND3X1  g0016(.A(n2143), .B(n2142), .C(n2307), .Y(n2144_1));
OR4X1    g0017(.A(n2382), .B(n2964), .C(n2133), .D(n2144_1), .Y(n2145));
NOR4X1   g0018(.A(n2129_1), .B(g1000), .C(g6850), .D(n2145), .Y(g1006));
NAND3X1  g0019(.A(n2143), .B(n2142), .C(g1013), .Y(n2147));
OR4X1    g0020(.A(n2382), .B(n2964), .C(n2133), .D(n2147), .Y(n2148));
NOR4X1   g0021(.A(n2129_1), .B(g1034), .C(n2135), .D(n2148), .Y(g1015));
INVX1    g0022(.A(g940), .Y(n2150));
XOR2X1   g0023(.A(g936), .B(n2150), .Y(n2151));
INVX1    g0024(.A(n2151), .Y(g4655));
OR4X1    g0025(.A(g1367), .B(g1373), .C(g1375), .D(g1374), .Y(n2153));
OR4X1    g0026(.A(g1363), .B(g1368), .C(g1369), .D(g1370), .Y(n2154_1));
OR4X1    g0027(.A(g1366), .B(g1365), .C(g1364), .D(n2154_1), .Y(n2155));
NOR4X1   g0028(.A(n2153), .B(g1372), .C(g1371), .D(n2155), .Y(g4657));
INVX1    g0029(.A(g1392), .Y(n2157));
NOR2X1   g0030(.A(g1391), .B(n2157), .Y(g4660));
INVX1    g0031(.A(g1394), .Y(n2159_1));
NOR2X1   g0032(.A(g1395), .B(n2159_1), .Y(g4661));
INVX1    g0033(.A(g1397), .Y(n2161));
NOR2X1   g0034(.A(g1398), .B(n2161), .Y(g4663));
INVX1    g0035(.A(g1400), .Y(n2163));
NOR2X1   g0036(.A(g1401), .B(n2163), .Y(g4664));
INVX1    g0037(.A(g889), .Y(n2165));
INVX1    g0038(.A(g887), .Y(n2166));
INVX1    g0039(.A(g888), .Y(n2167));
NOR3X1   g0040(.A(n2167), .B(n2166), .C(n2165), .Y(g5164));
INVX1    g0041(.A(g1486), .Y(g6223));
OR2X1    g0042(.A(g16), .B(g1189), .Y(g6236));
INVX1    g0043(.A(g1432), .Y(g6675));
XOR2X1   g0044(.A(g883), .B(g852), .Y(n2172));
XOR2X1   g0045(.A(g840), .B(g906), .Y(n2173));
XOR2X1   g0046(.A(g901), .B(g837), .Y(n2174_1));
XOR2X1   g0047(.A(g849), .B(g921), .Y(n2175));
NOR4X1   g0048(.A(n2174_1), .B(n2173), .C(n2172), .D(n2175), .Y(n2176));
XOR2X1   g0049(.A(g896), .B(g834), .Y(n2177));
XOR2X1   g0050(.A(g916), .B(g846), .Y(n2178));
XOR2X1   g0051(.A(g911), .B(g843), .Y(n2179_1));
XOR2X1   g0052(.A(g831), .B(g891), .Y(n2180));
NOR4X1   g0053(.A(n2179_1), .B(n2178), .C(n2177), .D(n2180), .Y(n2181));
OR4X1    g0054(.A(g887), .B(g778), .C(g889), .D(g888), .Y(n2182));
AOI21X1  g0055(.A0(n2181), .A1(n2176), .B0(n2182), .Y(g6849));
INVX1    g0056(.A(g689), .Y(g6895));
INVX1    g0057(.A(g855), .Y(n2185));
NAND2X1  g0058(.A(g944), .B(n2185), .Y(g7048));
NAND2X1  g0059(.A(g1405), .B(g1412), .Y(g7063));
NAND4X1  g0060(.A(g83), .B(g52), .C(g80), .D(g86), .Y(n2188));
INVX1    g0061(.A(n2188), .Y(n2189_1));
INVX1    g0062(.A(g68), .Y(n2190));
NOR4X1   g0063(.A(n2190), .B(g74), .C(g77), .D(g71), .Y(n2191));
NAND4X1  g0064(.A(n2189_1), .B(g7), .C(g58), .D(n2191), .Y(g7283));
NAND4X1  g0065(.A(n2189_1), .B(g6), .C(g58), .D(n2191), .Y(g7284));
NAND4X1  g0066(.A(n2189_1), .B(g58), .C(g5), .D(n2191), .Y(g7285));
NAND4X1  g0067(.A(n2189_1), .B(g58), .C(g4), .D(n2191), .Y(g7286));
NAND4X1  g0068(.A(n2189_1), .B(g2), .C(g58), .D(n2191), .Y(g7287));
NAND4X1  g0069(.A(n2189_1), .B(g58), .C(g3), .D(n2191), .Y(g7288));
NAND4X1  g0070(.A(n2189_1), .B(g58), .C(g48), .D(n2191), .Y(g7289));
NAND4X1  g0071(.A(n2189_1), .B(g8), .C(g58), .D(n2191), .Y(g7290));
NOR4X1   g0072(.A(g68), .B(g74), .C(g77), .D(g71), .Y(n2200));
NAND4X1  g0073(.A(n2189_1), .B(g58), .C(g48), .D(n2200), .Y(g7291));
NAND4X1  g0074(.A(n2189_1), .B(g58), .C(g3), .D(n2200), .Y(g7292));
NAND4X1  g0075(.A(n2189_1), .B(g2), .C(g58), .D(n2200), .Y(g7293));
INVX1    g0076(.A(g4), .Y(n2204_1));
INVX1    g0077(.A(g58), .Y(n2205));
OR4X1    g0078(.A(g68), .B(g74), .C(g77), .D(g71), .Y(n2206));
OR4X1    g0079(.A(n2188), .B(n2205), .C(n2204_1), .D(n2206), .Y(g7294));
NOR2X1   g0080(.A(g65), .B(g62), .Y(n2208));
OR2X1    g0081(.A(n2208), .B(g45), .Y(g7474));
AND2X1   g0082(.A(n2143), .B(g1034), .Y(g7514));
INVX1    g0083(.A(g1033), .Y(n2211));
NOR3X1   g0084(.A(n2211), .B(g1029), .C(g6850), .Y(n2212));
INVX1    g0085(.A(n2212), .Y(g8234));
ZERO     g0086(.Y(g8661));
INVX1    g0087(.A(g998), .Y(n2215));
INVX1    g0088(.A(g999), .Y(n2216));
NOR4X1   g0089(.A(n2215), .B(g1), .C(g1000), .D(n2216), .Y(n2217));
INVX1    g0090(.A(g1030), .Y(n2218));
INVX1    g0091(.A(n2964), .Y(n2219_1));
NAND3X1  g0092(.A(n2143), .B(n2219_1), .C(n2218), .Y(n2220));
OAI21X1  g0093(.A0(n2220), .A1(n2217), .B0(g1), .Y(g8872));
NOR2X1   g0094(.A(n2212), .B(g10), .Y(n2222));
OR2X1    g0095(.A(n2222), .B(n2217), .Y(n2223));
OAI21X1  g0096(.A0(n2223), .A1(n2220), .B0(g1), .Y(g8958));
MX2X1    g0097(.A(g31), .B(g30), .S0(g32), .Y(g9128));
INVX1    g0098(.A(g44), .Y(n2226));
OR2X1    g0099(.A(g55), .B(g42), .Y(n2227));
NOR4X1   g0100(.A(n2226), .B(g45), .C(g41), .D(n2227), .Y(n1899));
INVX1    g0101(.A(g77), .Y(n2229));
NOR4X1   g0102(.A(n2190), .B(g74), .C(n2229), .D(g71), .Y(n2230));
NAND3X1  g0103(.A(n2230), .B(n1899), .C(n2189_1), .Y(n2231));
INVX1    g0104(.A(g71), .Y(n2232));
NOR4X1   g0105(.A(g68), .B(g74), .C(g77), .D(n2232), .Y(n2233_1));
NAND3X1  g0106(.A(n2233_1), .B(n1899), .C(n2189_1), .Y(n2234));
NOR4X1   g0107(.A(g68), .B(g74), .C(n2229), .D(g71), .Y(n2235));
NAND3X1  g0108(.A(n2235), .B(n1899), .C(n2189_1), .Y(n2236));
NAND3X1  g0109(.A(n2236), .B(n2234), .C(n2231), .Y(n2237_1));
OR4X1    g0110(.A(n2226), .B(g45), .C(g41), .D(n2227), .Y(n2238));
INVX1    g0111(.A(g80), .Y(n2239));
OR4X1    g0112(.A(g83), .B(g52), .C(n2239), .D(g86), .Y(n2240));
AND2X1   g0113(.A(g74), .B(g77), .Y(n2241));
NAND3X1  g0114(.A(n2241), .B(n2232), .C(n2190), .Y(n2242_1));
NOR3X1   g0115(.A(n2242_1), .B(n2240), .C(n2238), .Y(n2243));
NAND3X1  g0116(.A(n2241), .B(n2232), .C(g68), .Y(n2244));
NOR3X1   g0117(.A(n2244), .B(n2240), .C(n2238), .Y(n2245));
NOR3X1   g0118(.A(n2238), .B(n2206), .C(n2188), .Y(n2246));
INVX1    g0119(.A(g74), .Y(n2247_1));
NAND4X1  g0120(.A(g68), .B(n2247_1), .C(n2229), .D(n2232), .Y(n2248));
NOR3X1   g0121(.A(n2238), .B(n2248), .C(n2188), .Y(n2249));
NAND4X1  g0122(.A(n2190), .B(g74), .C(n2229), .D(g71), .Y(n2250));
NOR3X1   g0123(.A(n2250), .B(n2238), .C(n2188), .Y(n2251_1));
NAND4X1  g0124(.A(g68), .B(n2247_1), .C(n2229), .D(g71), .Y(n2252));
NOR3X1   g0125(.A(n2252), .B(n2238), .C(n2188), .Y(n2253));
OR4X1    g0126(.A(n2251_1), .B(n2249), .C(n2246), .D(n2253), .Y(n2254));
NOR4X1   g0127(.A(n2245), .B(n2243), .C(n2237_1), .D(n2254), .Y(n2255));
NOR4X1   g0128(.A(g68), .B(n2247_1), .C(g77), .D(n2232), .Y(n2256_1));
NAND4X1  g0129(.A(n1899), .B(n2189_1), .C(g49), .D(n2256_1), .Y(n2257));
NAND4X1  g0130(.A(n1899), .B(n2189_1), .C(g710), .D(n2233_1), .Y(n2258));
NAND2X1  g0131(.A(n2258), .B(n2257), .Y(n2259));
INVX1    g0132(.A(g746), .Y(n2260));
NAND4X1  g0133(.A(n2200), .B(n2189_1), .C(g694), .D(n1899), .Y(n2261_1));
OAI21X1  g0134(.A0(n2231), .A1(n2260), .B0(n2261_1), .Y(n2262));
NOR4X1   g0135(.A(g83), .B(g52), .C(n2239), .D(g86), .Y(n2263));
NOR4X1   g0136(.A(g68), .B(n2247_1), .C(n2229), .D(g71), .Y(n2264));
NAND4X1  g0137(.A(n2263), .B(n1899), .C(g471), .D(n2264), .Y(n2265));
NOR4X1   g0138(.A(n2190), .B(n2247_1), .C(n2229), .D(g71), .Y(n2266_1));
NAND4X1  g0139(.A(n2263), .B(n1899), .C(g527), .D(n2266_1), .Y(n2267));
NOR4X1   g0140(.A(n2190), .B(g74), .C(g77), .D(n2232), .Y(n2268));
NAND4X1  g0141(.A(n1899), .B(n2189_1), .C(g685), .D(n2268), .Y(n2269));
NAND4X1  g0142(.A(n2191), .B(n2189_1), .C(g648), .D(n1899), .Y(n2270_1));
NAND4X1  g0143(.A(n2269), .B(n2267), .C(n2265), .D(n2270_1), .Y(n2271));
OR4X1    g0144(.A(n2262), .B(n2259), .C(n2255), .D(n2271), .Y(n2272));
NAND4X1  g0145(.A(n2190), .B(n2247_1), .C(g77), .D(g71), .Y(n2273_1));
INVX1    g0146(.A(n2273_1), .Y(n2274));
OAI21X1  g0147(.A0(n2274), .A1(n2235), .B0(n2263), .Y(n2275));
NOR4X1   g0148(.A(n2190), .B(g74), .C(n2229), .D(n2232), .Y(n2276));
OAI21X1  g0149(.A0(n2276), .A1(n2230), .B0(n2263), .Y(n2277));
NAND4X1  g0150(.A(n2190), .B(n2247_1), .C(n2229), .D(g71), .Y(n2278_1));
AOI21X1  g0151(.A0(n2252), .A1(n2278_1), .B0(n2240), .Y(n2279));
NAND4X1  g0152(.A(g68), .B(g74), .C(n2229), .D(n2232), .Y(n2280));
AOI21X1  g0153(.A0(n2280), .A1(n2250), .B0(n2240), .Y(n2281));
NAND4X1  g0154(.A(g68), .B(g74), .C(n2229), .D(g71), .Y(n2282));
NAND4X1  g0155(.A(n2190), .B(g74), .C(n2229), .D(n2232), .Y(n2283_1));
AOI21X1  g0156(.A0(n2283_1), .A1(n2282), .B0(n2240), .Y(n2284));
NOR3X1   g0157(.A(n2284), .B(n2281), .C(n2279), .Y(n2285));
NAND3X1  g0158(.A(n2285), .B(n2277), .C(n2275), .Y(n2286));
NOR3X1   g0159(.A(n2273_1), .B(n2240), .C(n2238), .Y(n2287));
NOR3X1   g0160(.A(n2250), .B(n2240), .C(n2238), .Y(n2288_1));
NAND4X1  g0161(.A(n2190), .B(n2247_1), .C(g77), .D(n2232), .Y(n2289));
NOR3X1   g0162(.A(n2240), .B(n2289), .C(n2238), .Y(n2290));
NAND3X1  g0163(.A(n2276), .B(n2263), .C(n1899), .Y(n2291));
NAND3X1  g0164(.A(n2263), .B(n2230), .C(n1899), .Y(n2292));
NOR4X1   g0165(.A(n2190), .B(n2247_1), .C(g77), .D(n2232), .Y(n2293_1));
NAND3X1  g0166(.A(n2293_1), .B(n2263), .C(n1899), .Y(n2294));
NAND3X1  g0167(.A(n2294), .B(n2292), .C(n2291), .Y(n2295));
NOR4X1   g0168(.A(n2290), .B(n2288_1), .C(n2287), .D(n2295), .Y(n2296));
NAND4X1  g0169(.A(n2263), .B(n1899), .C(g852), .D(n2276), .Y(n2297_1));
NAND4X1  g0170(.A(g68), .B(n2247_1), .C(g77), .D(n2232), .Y(n2298));
NOR3X1   g0171(.A(n2240), .B(n2298), .C(n2238), .Y(n2299));
NOR3X1   g0172(.A(n2282), .B(n2240), .C(n2238), .Y(n2300));
AOI22X1  g0173(.A0(n2299), .A1(g48), .B0(g855), .B1(n2300), .Y(n2301));
NAND2X1  g0174(.A(n2301), .B(n2297_1), .Y(n2302_1));
NAND4X1  g0175(.A(g68), .B(n2247_1), .C(g77), .D(g71), .Y(n2303));
NOR3X1   g0176(.A(n2303), .B(n2240), .C(n2238), .Y(n2304));
OR2X1    g0177(.A(n2304), .B(n2290), .Y(n2305));
OR4X1    g0178(.A(n2299), .B(n2288_1), .C(n2287), .D(n2300), .Y(n2306));
OR2X1    g0179(.A(n2306), .B(n2305), .Y(n2307_1));
OAI21X1  g0180(.A0(n2302_1), .A1(n2296), .B0(n2307_1), .Y(n2308));
NOR3X1   g0181(.A(n2280), .B(n2240), .C(n2238), .Y(n2309));
NOR3X1   g0182(.A(n2283_1), .B(n2240), .C(n2238), .Y(n2310));
NOR3X1   g0183(.A(n2252), .B(n2240), .C(n2238), .Y(n2311));
NOR3X1   g0184(.A(n2240), .B(n2278_1), .C(n2238), .Y(n2312_1));
OR4X1    g0185(.A(n2311), .B(n2310), .C(n2309), .D(n2312_1), .Y(n2313));
OR4X1    g0186(.A(n2306), .B(n2304), .C(n2290), .D(n2313), .Y(n2314));
NAND4X1  g0187(.A(n2233_1), .B(n1899), .C(g758), .D(n2263), .Y(n2315));
AOI22X1  g0188(.A0(n2309), .A1(g774), .B0(g766), .B1(n2311), .Y(n2316));
NAND4X1  g0189(.A(n2315), .B(n2314), .C(n2308), .D(n2316), .Y(n2317_1));
MX2X1    g0190(.A(n2272), .B(n2317_1), .S0(n2286), .Y(n2318));
NOR4X1   g0191(.A(g83), .B(g52), .C(g80), .D(g86), .Y(n2319));
OAI21X1  g0192(.A0(n2274), .A1(n2230), .B0(n2319), .Y(n2320));
OAI21X1  g0193(.A0(n2264), .A1(n2235), .B0(n2319), .Y(n2321));
OAI21X1  g0194(.A0(n2276), .A1(n2266_1), .B0(n2319), .Y(n2322_1));
NAND3X1  g0195(.A(n2322_1), .B(n2321), .C(n2320), .Y(n2323));
NOR4X1   g0196(.A(g68), .B(n2247_1), .C(g77), .D(g71), .Y(n2324));
OAI21X1  g0197(.A0(n2324), .A1(n2200), .B0(n2319), .Y(n2325));
NOR4X1   g0198(.A(n2190), .B(n2247_1), .C(g77), .D(g71), .Y(n2326));
OAI21X1  g0199(.A0(n2326), .A1(n2268), .B0(n2319), .Y(n2327_1));
NAND2X1  g0200(.A(n2327_1), .B(n2325), .Y(n2328));
AOI22X1  g0201(.A0(n2293_1), .A1(n2319), .B0(n2263), .B1(n2191), .Y(n2329));
OAI21X1  g0202(.A0(n2233_1), .A1(n2191), .B0(n2319), .Y(n2330));
NAND2X1  g0203(.A(n2330), .B(n2329), .Y(n2331));
NAND4X1  g0204(.A(n2241), .B(g71), .C(g68), .D(n2319), .Y(n2332_1));
OAI21X1  g0205(.A0(n2240), .A1(n2206), .B0(n2332_1), .Y(n2333));
OR4X1    g0206(.A(g83), .B(g52), .C(g80), .D(g86), .Y(n2334));
NAND4X1  g0207(.A(n2241), .B(g71), .C(n2190), .D(n2319), .Y(n2335));
OAI21X1  g0208(.A0(n2334), .A1(n2250), .B0(n2335), .Y(n2336));
OR2X1    g0209(.A(n2336), .B(n2333), .Y(n2337_1));
NOR4X1   g0210(.A(n2331), .B(n2328), .C(n2323), .D(n2337_1), .Y(n2338));
NOR3X1   g0211(.A(n2240), .B(n2238), .C(n2248), .Y(n2339));
NOR3X1   g0212(.A(n2240), .B(n2238), .C(n2206), .Y(n2340));
NOR3X1   g0213(.A(n2334), .B(n2283_1), .C(n2238), .Y(n2341));
NOR3X1   g0214(.A(n2334), .B(n2280), .C(n2238), .Y(n2342_1));
NOR3X1   g0215(.A(n2334), .B(n2282), .C(n2238), .Y(n2343));
NOR3X1   g0216(.A(n2334), .B(n2250), .C(n2238), .Y(n2344));
OR4X1    g0217(.A(n2343), .B(n2342_1), .C(n2341), .D(n2344), .Y(n2345));
NOR3X1   g0218(.A(n2334), .B(n2242_1), .C(n2238), .Y(n2346));
NOR3X1   g0219(.A(n2334), .B(n2244), .C(n2238), .Y(n2347_1));
NOR2X1   g0220(.A(n2335), .B(n2238), .Y(n2348));
NOR2X1   g0221(.A(n2332_1), .B(n2238), .Y(n2349));
NOR4X1   g0222(.A(n2348), .B(n2347_1), .C(n2346), .D(n2349), .Y(n2350));
NOR3X1   g0223(.A(n2334), .B(n2289), .C(n2238), .Y(n2351));
NOR3X1   g0224(.A(n2334), .B(n2298), .C(n2238), .Y(n2352_1));
NOR3X1   g0225(.A(n2334), .B(n2303), .C(n2238), .Y(n2353));
NOR3X1   g0226(.A(n2334), .B(n2273_1), .C(n2238), .Y(n2354));
NOR4X1   g0227(.A(n2353), .B(n2352_1), .C(n2351), .D(n2354), .Y(n2355));
NOR3X1   g0228(.A(n2334), .B(n2278_1), .C(n2238), .Y(n2356));
NOR3X1   g0229(.A(n2334), .B(n2252), .C(n2238), .Y(n2357_1));
NOR3X1   g0230(.A(n2334), .B(n2238), .C(n2248), .Y(n2358));
NOR3X1   g0231(.A(n2334), .B(n2238), .C(n2206), .Y(n2359));
NOR4X1   g0232(.A(n2358), .B(n2357_1), .C(n2356), .D(n2359), .Y(n2360));
NAND3X1  g0233(.A(n2360), .B(n2355), .C(n2350), .Y(n2361));
OR4X1    g0234(.A(n2345), .B(n2340), .C(n2339), .D(n2361), .Y(n2362_1));
AOI22X1  g0235(.A0(n2339), .A1(g632), .B0(g624), .B1(n2340), .Y(n2363));
AOI22X1  g0236(.A0(n2341), .A1(g228), .B0(g284), .B1(n2342_1), .Y(n2364));
AOI22X1  g0237(.A0(n2343), .A1(g365), .B0(g309), .B1(n2344), .Y(n2365));
NAND3X1  g0238(.A(n2365), .B(n2364), .C(n2363), .Y(n2366));
NAND2X1  g0239(.A(n2348), .B(g613), .Y(n2367_1));
AOI22X1  g0240(.A0(n2346), .A1(g600), .B0(g621), .B1(n2349), .Y(n2368));
NAND2X1  g0241(.A(n2368), .B(n2367_1), .Y(n2369));
NAND4X1  g0242(.A(n2235), .B(n1899), .C(g390), .D(n2319), .Y(n2370));
NAND4X1  g0243(.A(n2230), .B(n1899), .C(g446), .D(n2319), .Y(n2371));
NAND4X1  g0244(.A(n2266_1), .B(n1899), .C(g608), .D(n2319), .Y(n2372_1));
NAND4X1  g0245(.A(n2276), .B(n1899), .C(g553), .D(n2319), .Y(n2373));
NAND4X1  g0246(.A(n2372_1), .B(n2371), .C(n2370), .D(n2373), .Y(n2374));
NAND4X1  g0247(.A(n2233_1), .B(n1899), .C(g110), .D(n2319), .Y(n2375));
NAND4X1  g0248(.A(n2268), .B(n1899), .C(g142), .D(n2319), .Y(n2376));
NAND4X1  g0249(.A(n1899), .B(n2191), .C(g185), .D(n2319), .Y(n2377_1));
NAND4X1  g0250(.A(n1899), .B(n2200), .C(g168), .D(n2319), .Y(n2378));
NAND4X1  g0251(.A(n2377_1), .B(n2376), .C(n2375), .D(n2378), .Y(n2379));
NOR4X1   g0252(.A(n2374), .B(n2369), .C(n2366), .D(n2379), .Y(n2380));
AOI21X1  g0253(.A0(n2380), .A1(n2362_1), .B0(n2338), .Y(n2381));
AOI21X1  g0254(.A0(n2338), .A1(n2318), .B0(n2381), .Y(n2382_1));
NAND2X1  g0255(.A(n2382_1), .B(g62), .Y(g9280));
INVX1    g0256(.A(g62), .Y(n2384));
OR4X1    g0257(.A(n2331), .B(n2328), .C(n2323), .D(n2337_1), .Y(n2385));
NOR3X1   g0258(.A(n2278_1), .B(n2238), .C(n2188), .Y(n2386));
AOI22X1  g0259(.A0(n2386), .A1(g714), .B0(g757), .B1(n2251_1), .Y(n2387_1));
INVX1    g0260(.A(g741), .Y(n2388));
NOR4X1   g0261(.A(n2238), .B(n2188), .C(n2388), .D(n2298), .Y(n2389));
AOI21X1  g0262(.A0(n2246), .A1(g698), .B0(n2389), .Y(n2390));
AOI22X1  g0263(.A0(n2243), .A1(g468), .B0(g524), .B1(n2245), .Y(n2391));
AOI22X1  g0264(.A0(n2249), .A1(g647), .B0(g681), .B1(n2253), .Y(n2392_1));
NAND4X1  g0265(.A(n2391), .B(n2390), .C(n2387_1), .D(n2392_1), .Y(n2393));
NOR2X1   g0266(.A(n2393), .B(n2255), .Y(n2394));
NOR3X1   g0267(.A(n2313), .B(n2306), .C(n2305), .Y(n2395));
NAND4X1  g0268(.A(n2263), .B(n1899), .C(g849), .D(n2276), .Y(n2398));
AOI22X1  g0269(.A0(n2299), .A1(g3), .B0(g859), .B1(n2300), .Y(n2399));
AND2X1   g0270(.A(n2399), .B(n2398), .Y(n2400));
AOI21X1  g0271(.A0(n2400), .A1(n2307_1), .B0(n2296), .Y(n2401));
NAND4X1  g0272(.A(n2263), .B(n1899), .C(g765), .D(n2268), .Y(n2402_1));
NAND4X1  g0273(.A(n2263), .B(n1899), .C(g773), .D(n2326), .Y(n2403));
NAND2X1  g0274(.A(n2403), .B(n2402_1), .Y(n2404));
NOR3X1   g0275(.A(n2404), .B(n2401), .C(n2395), .Y(n2405));
MX2X1    g0276(.A(n2394), .B(n2405), .S0(n2286), .Y(n2406));
NOR4X1   g0277(.A(n2345), .B(n2340), .C(n2339), .D(n2361), .Y(n2407_1));
NAND4X1  g0278(.A(n1899), .B(n2200), .C(g623), .D(n2263), .Y(n2408));
NAND4X1  g0279(.A(n1899), .B(n2191), .C(g631), .D(n2263), .Y(n2409));
NAND2X1  g0280(.A(n2409), .B(n2408), .Y(n2410));
NAND4X1  g0281(.A(n2324), .B(n1899), .C(g225), .D(n2319), .Y(n2411));
NAND4X1  g0282(.A(n2326), .B(n1899), .C(g281), .D(n2319), .Y(n2412_1));
NAND4X1  g0283(.A(n2293_1), .B(n1899), .C(g362), .D(n2319), .Y(n2413));
NAND4X1  g0284(.A(n2256_1), .B(n1899), .C(g306), .D(n2319), .Y(n2414));
NAND4X1  g0285(.A(n2413), .B(n2412_1), .C(n2411), .D(n2414), .Y(n2415));
NOR2X1   g0286(.A(n2415), .B(n2410), .Y(n2416));
NAND2X1  g0287(.A(n2349), .B(g620), .Y(n2417_1));
AOI22X1  g0288(.A0(n2347_1), .A1(g607), .B0(g612), .B1(n2348), .Y(n2418));
NAND4X1  g0289(.A(n2235), .B(n1899), .C(g387), .D(n2319), .Y(n2419));
NAND4X1  g0290(.A(n2230), .B(n1899), .C(g443), .D(n2319), .Y(n2420));
NAND4X1  g0291(.A(n2264), .B(n1899), .C(g599), .D(n2319), .Y(n2421));
NAND4X1  g0292(.A(n2276), .B(n1899), .C(g550), .D(n2319), .Y(n2422_1));
NAND4X1  g0293(.A(n2421), .B(n2420), .C(n2419), .D(n2422_1), .Y(n2423));
NAND4X1  g0294(.A(n2233_1), .B(n1899), .C(g105), .D(n2319), .Y(n2424));
NAND4X1  g0295(.A(n2268), .B(n1899), .C(g138), .D(n2319), .Y(n2425));
NAND4X1  g0296(.A(n1899), .B(n2191), .C(g182), .D(n2319), .Y(n2426));
NAND4X1  g0297(.A(n1899), .B(n2200), .C(g162), .D(n2319), .Y(n2427_1));
NAND4X1  g0298(.A(n2426), .B(n2425), .C(n2424), .D(n2427_1), .Y(n2428));
NOR2X1   g0299(.A(n2428), .B(n2423), .Y(n2429));
NAND4X1  g0300(.A(n2418), .B(n2417_1), .C(n2416), .D(n2429), .Y(n2430));
OAI21X1  g0301(.A0(n2430), .A1(n2407_1), .B0(n2385), .Y(n2431));
OAI21X1  g0302(.A0(n2406), .A1(n2385), .B0(n2431), .Y(n2432_1));
OR2X1    g0303(.A(n2432_1), .B(n2384), .Y(g9297));
OR4X1    g0304(.A(n2245), .B(n2243), .C(n2237_1), .D(n2254), .Y(n2434));
NAND4X1  g0305(.A(n2191), .B(n2189_1), .C(g652), .D(n1899), .Y(n2435));
NAND4X1  g0306(.A(n2263), .B(n1899), .C(g513), .D(n2266_1), .Y(n2436));
NAND2X1  g0307(.A(n2436), .B(n2435), .Y(n2437_1));
AOI21X1  g0308(.A0(n2243), .A1(g465), .B0(n2437_1), .Y(n2438));
AOI22X1  g0309(.A0(n2386), .A1(g718), .B0(g677), .B1(n2253), .Y(n2439));
AOI22X1  g0310(.A0(n2246), .A1(g702), .B0(g756), .B1(n2251_1), .Y(n2440));
NAND4X1  g0311(.A(n2439), .B(n2438), .C(n2434), .D(n2440), .Y(n2441));
NAND4X1  g0312(.A(n2263), .B(n1899), .C(g846), .D(n2276), .Y(n2442_1));
AOI22X1  g0313(.A0(n2299), .A1(g2), .B0(g863), .B1(n2300), .Y(n2443));
NAND2X1  g0314(.A(n2443), .B(n2442_1), .Y(n2444));
OAI21X1  g0315(.A0(n2444), .A1(n2296), .B0(n2307_1), .Y(n2445));
AOI22X1  g0316(.A0(n2309), .A1(g772), .B0(g764), .B1(n2311), .Y(n2446));
NAND3X1  g0317(.A(n2446), .B(n2445), .C(n2314), .Y(n2447_1));
MX2X1    g0318(.A(n2441), .B(n2447_1), .S0(n2286), .Y(n2448));
AOI22X1  g0319(.A0(n2339), .A1(g630), .B0(g622), .B1(n2340), .Y(n2449));
AOI22X1  g0320(.A0(n2341), .A1(g222), .B0(g270), .B1(n2342_1), .Y(n2450));
AOI22X1  g0321(.A0(n2343), .A1(g351), .B0(g303), .B1(n2344), .Y(n2451));
NAND3X1  g0322(.A(n2451), .B(n2450), .C(n2449), .Y(n2452_1));
AND2X1   g0323(.A(n2349), .B(g619), .Y(n2453));
NAND4X1  g0324(.A(n2266_1), .B(n1899), .C(g606), .D(n2319), .Y(n2454));
NAND2X1  g0325(.A(n2348), .B(g611), .Y(n2455));
NAND2X1  g0326(.A(n2455), .B(n2454), .Y(n2456));
AOI22X1  g0327(.A0(n2351), .A1(g384), .B0(g432), .B1(n2352_1), .Y(n2457_1));
AOI22X1  g0328(.A0(n2346), .A1(g598), .B0(g547), .B1(n2353), .Y(n2458));
AOI22X1  g0329(.A0(n2356), .A1(g100), .B0(g134), .B1(n2357_1), .Y(n2459));
AOI22X1  g0330(.A0(n2358), .A1(g181), .B0(g158), .B1(n2359), .Y(n2460));
NAND4X1  g0331(.A(n2459), .B(n2458), .C(n2457_1), .D(n2460), .Y(n2461));
NOR4X1   g0332(.A(n2456), .B(n2453), .C(n2452_1), .D(n2461), .Y(n2462_1));
AOI21X1  g0333(.A0(n2462_1), .A1(n2362_1), .B0(n2338), .Y(n2463));
AOI21X1  g0334(.A0(n2448), .A1(n2338), .B0(n2463), .Y(n2464));
NAND2X1  g0335(.A(n2464), .B(g62), .Y(g9299));
NAND4X1  g0336(.A(n2191), .B(n2189_1), .C(g645), .D(n1899), .Y(n2466_1));
NAND4X1  g0337(.A(n2263), .B(n1899), .C(g510), .D(n2266_1), .Y(n2467));
NAND2X1  g0338(.A(n2467), .B(n2466_1), .Y(n2468));
AOI21X1  g0339(.A0(n2243), .A1(g462), .B0(n2468), .Y(n2469));
AOI22X1  g0340(.A0(n2246), .A1(g722), .B0(g673), .B1(n2253), .Y(n2470_1));
AOI22X1  g0341(.A0(n2386), .A1(g734), .B0(g753), .B1(n2251_1), .Y(n2471));
NAND4X1  g0342(.A(n2470_1), .B(n2469), .C(n2434), .D(n2471), .Y(n2472));
AOI22X1  g0343(.A0(n2304), .A1(g843), .B0(g4), .B1(n2299), .Y(n2473));
AOI21X1  g0344(.A0(n2473), .A1(n2307_1), .B0(n2296), .Y(n2474_1));
AOI22X1  g0345(.A0(n2309), .A1(g771), .B0(g763), .B1(n2311), .Y(n2475));
NAND2X1  g0346(.A(n2475), .B(n2314), .Y(n2476));
OR2X1    g0347(.A(n2476), .B(n2474_1), .Y(n2477_1));
MX2X1    g0348(.A(n2472), .B(n2477_1), .S0(n2286), .Y(n2478));
AOI22X1  g0349(.A0(n2356), .A1(g95), .B0(g130), .B1(n2357_1), .Y(n2479));
AOI22X1  g0350(.A0(n2358), .A1(g180), .B0(g154), .B1(n2359), .Y(n2480));
NAND2X1  g0351(.A(n2480), .B(n2479), .Y(n2481_1));
NAND4X1  g0352(.A(n2324), .B(n1899), .C(g219), .D(n2319), .Y(n2482));
NAND4X1  g0353(.A(n2326), .B(n1899), .C(g267), .D(n2319), .Y(n2483));
NAND4X1  g0354(.A(n2293_1), .B(n1899), .C(g348), .D(n2319), .Y(n2484));
NAND4X1  g0355(.A(n2256_1), .B(n1899), .C(g300), .D(n2319), .Y(n2485));
NAND4X1  g0356(.A(n2484), .B(n2483), .C(n2482), .D(n2485), .Y(n2486_1));
AOI22X1  g0357(.A0(n2347_1), .A1(g605), .B0(g610), .B1(n2348), .Y(n2487));
AOI22X1  g0358(.A0(n2339), .A1(g629), .B0(g618), .B1(n2349), .Y(n2488));
AOI22X1  g0359(.A0(n2351), .A1(g381), .B0(g429), .B1(n2352_1), .Y(n2489));
AOI22X1  g0360(.A0(n2346), .A1(g597), .B0(g573), .B1(n2353), .Y(n2490));
NAND4X1  g0361(.A(n2489), .B(n2488), .C(n2487), .D(n2490), .Y(n2491_1));
NOR3X1   g0362(.A(n2491_1), .B(n2486_1), .C(n2481_1), .Y(n2492));
AOI21X1  g0363(.A0(n2492), .A1(n2362_1), .B0(n2338), .Y(n2493));
AOI21X1  g0364(.A0(n2478), .A1(n2338), .B0(n2493), .Y(n2494));
NAND2X1  g0365(.A(n2494), .B(g62), .Y(g9305));
NAND4X1  g0366(.A(n2263), .B(n1899), .C(g459), .D(n2264), .Y(n2496_1));
AOI22X1  g0367(.A0(n2245), .A1(g507), .B0(g635), .B1(n2249), .Y(n2497));
AOI22X1  g0368(.A0(n2386), .A1(g730), .B0(g669), .B1(n2253), .Y(n2498));
AOI22X1  g0369(.A0(n2246), .A1(g723), .B0(g752), .B1(n2251_1), .Y(n2499));
NAND4X1  g0370(.A(n2498), .B(n2497), .C(n2496_1), .D(n2499), .Y(n2500));
NOR2X1   g0371(.A(n2500), .B(n2255), .Y(n2501_1));
AOI22X1  g0372(.A0(n2304), .A1(g840), .B0(g5), .B1(n2299), .Y(n2502));
AOI21X1  g0373(.A0(n2502), .A1(n2307_1), .B0(n2296), .Y(n2503));
NAND4X1  g0374(.A(n2263), .B(n1899), .C(g762), .D(n2268), .Y(n2504));
NAND4X1  g0375(.A(n2263), .B(n1899), .C(g770), .D(n2326), .Y(n2505));
NAND2X1  g0376(.A(n2505), .B(n2504), .Y(n2506_1));
NOR3X1   g0377(.A(n2506_1), .B(n2503), .C(n2395), .Y(n2507));
MX2X1    g0378(.A(n2501_1), .B(n2507), .S0(n2286), .Y(n2508));
AOI22X1  g0379(.A0(n2356), .A1(g89), .B0(g126), .B1(n2357_1), .Y(n2509));
AOI22X1  g0380(.A0(n2358), .A1(g179), .B0(g174), .B1(n2359), .Y(n2510));
NAND2X1  g0381(.A(n2510), .B(n2509), .Y(n2511_1));
NAND4X1  g0382(.A(n2324), .B(n1899), .C(g216), .D(n2319), .Y(n2512));
NAND4X1  g0383(.A(n2326), .B(n1899), .C(g264), .D(n2319), .Y(n2513));
NAND4X1  g0384(.A(n2293_1), .B(n1899), .C(g345), .D(n2319), .Y(n2514));
NAND4X1  g0385(.A(n2256_1), .B(n1899), .C(g297), .D(n2319), .Y(n2515));
NAND4X1  g0386(.A(n2514), .B(n2513), .C(n2512), .D(n2515), .Y(n2516_1));
AOI22X1  g0387(.A0(n2347_1), .A1(g604), .B0(g609), .B1(n2348), .Y(n2517));
AOI22X1  g0388(.A0(n2339), .A1(g628), .B0(g617), .B1(n2349), .Y(n2518));
NAND2X1  g0389(.A(n2518), .B(n2517), .Y(n2519));
NAND4X1  g0390(.A(n2235), .B(n1899), .C(g378), .D(n2319), .Y(n2520));
NAND4X1  g0391(.A(n2230), .B(n1899), .C(g426), .D(n2319), .Y(n2521_1));
NAND4X1  g0392(.A(n2264), .B(n1899), .C(g596), .D(n2319), .Y(n2522));
NAND4X1  g0393(.A(n2276), .B(n1899), .C(g591), .D(n2319), .Y(n2523));
NAND4X1  g0394(.A(n2522), .B(n2521_1), .C(n2520), .D(n2523), .Y(n2524));
OR4X1    g0395(.A(n2519), .B(n2516_1), .C(n2511_1), .D(n2524), .Y(n2525));
OAI21X1  g0396(.A0(n2525), .A1(n2407_1), .B0(n2385), .Y(n2526_1));
OAI21X1  g0397(.A0(n2508), .A1(n2385), .B0(n2526_1), .Y(n2527));
OR2X1    g0398(.A(n2527), .B(n2384), .Y(g9308));
AOI22X1  g0399(.A0(n2251_1), .A1(g754), .B0(g665), .B1(n2253), .Y(n2529));
AOI22X1  g0400(.A0(n2245), .A1(g504), .B0(g634), .B1(n2249), .Y(n2530));
NAND3X1  g0401(.A(n2530), .B(n2529), .C(n2434), .Y(n2531_1));
NAND4X1  g0402(.A(n2263), .B(n1899), .C(g837), .D(n2276), .Y(n2532));
NAND4X1  g0403(.A(n2230), .B(n1899), .C(g6), .D(n2263), .Y(n2533));
NAND2X1  g0404(.A(n2533), .B(n2532), .Y(n2534));
OAI21X1  g0405(.A0(n2534), .A1(n2296), .B0(n2307_1), .Y(n2535));
AOI22X1  g0406(.A0(n2309), .A1(g769), .B0(g761), .B1(n2311), .Y(n2536_1));
NAND3X1  g0407(.A(n2536_1), .B(n2535), .C(n2314), .Y(n2537));
MX2X1    g0408(.A(n2531_1), .B(n2537), .S0(n2286), .Y(n2538));
NAND4X1  g0409(.A(n2326), .B(n1899), .C(g261), .D(n2319), .Y(n2539));
NAND4X1  g0410(.A(n1899), .B(n2191), .C(g184), .D(n2319), .Y(n2540));
NAND2X1  g0411(.A(n2540), .B(n2539), .Y(n2541_1));
INVX1    g0412(.A(g616), .Y(n2542));
OR2X1    g0413(.A(n2332_1), .B(n2238), .Y(n2543));
NAND4X1  g0414(.A(n1899), .B(n2191), .C(g627), .D(n2263), .Y(n2544));
OAI21X1  g0415(.A0(n2543), .A1(n2542), .B0(n2544), .Y(n2545));
NAND4X1  g0416(.A(n2293_1), .B(n1899), .C(g342), .D(n2319), .Y(n2546_1));
NAND4X1  g0417(.A(n2230), .B(n1899), .C(g423), .D(n2319), .Y(n2547));
AOI22X1  g0418(.A0(n2347_1), .A1(g603), .B0(g588), .B1(n2353), .Y(n2548));
AOI22X1  g0419(.A0(n2357_1), .A1(g122), .B0(g150), .B1(n2359), .Y(n2549));
NAND4X1  g0420(.A(n2548), .B(n2547), .C(n2546_1), .D(n2549), .Y(n2550));
NOR3X1   g0421(.A(n2550), .B(n2545), .C(n2541_1), .Y(n2551_1));
AOI21X1  g0422(.A0(n2551_1), .A1(n2362_1), .B0(n2338), .Y(n2552));
AOI21X1  g0423(.A0(n2538), .A1(n2338), .B0(n2552), .Y(n2553));
NAND2X1  g0424(.A(n2553), .B(g62), .Y(g9310));
NAND4X1  g0425(.A(n1899), .B(n2189_1), .C(g661), .D(n2268), .Y(n2555));
NAND4X1  g0426(.A(n1899), .B(n2189_1), .C(g755), .D(n2256_1), .Y(n2556_1));
NAND4X1  g0427(.A(n2263), .B(n1899), .C(g501), .D(n2266_1), .Y(n2557));
NAND4X1  g0428(.A(n2191), .B(n2189_1), .C(g633), .D(n1899), .Y(n2558));
NAND4X1  g0429(.A(n2557), .B(n2556_1), .C(n2555), .D(n2558), .Y(n2559));
NOR2X1   g0430(.A(n2559), .B(n2255), .Y(n2560));
AOI22X1  g0431(.A0(n2304), .A1(g834), .B0(g7), .B1(n2299), .Y(n2561_1));
AOI21X1  g0432(.A0(n2561_1), .A1(n2307_1), .B0(n2296), .Y(n2562));
NAND4X1  g0433(.A(n2263), .B(n1899), .C(g760), .D(n2268), .Y(n2563));
NAND4X1  g0434(.A(n2263), .B(n1899), .C(g768), .D(n2326), .Y(n2564));
NAND3X1  g0435(.A(n2564), .B(n2563), .C(n2314), .Y(n2565_1));
OAI21X1  g0436(.A0(n2565_1), .A1(n2562), .B0(n2286), .Y(n2566));
OAI21X1  g0437(.A0(n2560), .A1(n2286), .B0(n2566), .Y(n2567));
NAND4X1  g0438(.A(n2326), .B(n1899), .C(g258), .D(n2319), .Y(n2568));
NAND4X1  g0439(.A(n1899), .B(n2191), .C(g183), .D(n2319), .Y(n2569));
AND2X1   g0440(.A(n2569), .B(n2568), .Y(n2570_1));
AOI22X1  g0441(.A0(n2339), .A1(g626), .B0(g615), .B1(n2349), .Y(n2571));
NAND4X1  g0442(.A(n2293_1), .B(n1899), .C(g339), .D(n2319), .Y(n2572));
NAND4X1  g0443(.A(n2230), .B(n1899), .C(g420), .D(n2319), .Y(n2573));
AND2X1   g0444(.A(n2573), .B(n2572), .Y(n2574));
AOI22X1  g0445(.A0(n2347_1), .A1(g602), .B0(g570), .B1(n2353), .Y(n2575_1));
AOI22X1  g0446(.A0(n2357_1), .A1(g118), .B0(g173), .B1(n2359), .Y(n2576));
AND2X1   g0447(.A(n2576), .B(n2575_1), .Y(n2577));
NAND4X1  g0448(.A(n2574), .B(n2571), .C(n2570_1), .D(n2577), .Y(n2578));
OR2X1    g0449(.A(n2578), .B(n2407_1), .Y(n2579));
MX2X1    g0450(.A(n2567), .B(n2579), .S0(n2385), .Y(n2580_1));
OR2X1    g0451(.A(n2580_1), .B(n2384), .Y(g9312));
AOI22X1  g0452(.A0(n2251_1), .A1(g751), .B0(g706), .B1(n2253), .Y(n2582));
AOI22X1  g0453(.A0(n2245), .A1(g498), .B0(g690), .B1(n2249), .Y(n2583));
NAND3X1  g0454(.A(n2583), .B(n2582), .C(n2434), .Y(n2584));
AOI22X1  g0455(.A0(n2304), .A1(g831), .B0(g8), .B1(n2299), .Y(n2585_1));
AOI21X1  g0456(.A0(n2585_1), .A1(n2307_1), .B0(n2296), .Y(n2586));
AOI22X1  g0457(.A0(n2309), .A1(g767), .B0(g759), .B1(n2311), .Y(n2587));
NAND2X1  g0458(.A(n2587), .B(n2314), .Y(n2588));
OR2X1    g0459(.A(n2588), .B(n2586), .Y(n2589));
MX2X1    g0460(.A(n2584), .B(n2589), .S0(n2286), .Y(n2590_1));
NAND4X1  g0461(.A(n2266_1), .B(n1899), .C(g601), .D(n2319), .Y(n2591));
AOI22X1  g0462(.A0(n2352_1), .A1(g417), .B0(g563), .B1(n2353), .Y(n2592));
NAND2X1  g0463(.A(n2592), .B(n2591), .Y(n2593));
INVX1    g0464(.A(g614), .Y(n2594));
NAND4X1  g0465(.A(n1899), .B(n2191), .C(g625), .D(n2263), .Y(n2595_1));
OAI21X1  g0466(.A0(n2543), .A1(n2594), .B0(n2595_1), .Y(n2596));
NAND4X1  g0467(.A(n2268), .B(n1899), .C(g114), .D(n2319), .Y(n2597));
NAND4X1  g0468(.A(n1899), .B(n2200), .C(g146), .D(n2319), .Y(n2598));
NAND4X1  g0469(.A(n2293_1), .B(n1899), .C(g336), .D(n2319), .Y(n2599));
NAND4X1  g0470(.A(n2326), .B(n1899), .C(g255), .D(n2319), .Y(n2600_1));
NAND4X1  g0471(.A(n2599), .B(n2598), .C(n2597), .D(n2600_1), .Y(n2601));
NOR3X1   g0472(.A(n2601), .B(n2596), .C(n2593), .Y(n2602));
AOI21X1  g0473(.A0(n2602), .A1(n2362_1), .B0(n2338), .Y(n2603));
AOI21X1  g0474(.A0(n2590_1), .A1(n2338), .B0(n2603), .Y(n2604));
NAND2X1  g0475(.A(n2604), .B(g62), .Y(g9314));
XOR2X1   g0476(.A(g7), .B(g8), .Y(n2606));
XOR2X1   g0477(.A(g6), .B(g5), .Y(n2607));
XOR2X1   g0478(.A(n2607), .B(n2606), .Y(n2608));
XOR2X1   g0479(.A(g2), .B(g4), .Y(n2609_1));
XOR2X1   g0480(.A(g3), .B(g48), .Y(n2610));
XOR2X1   g0481(.A(n2610), .B(n2609_1), .Y(n2611));
XOR2X1   g0482(.A(n2611), .B(n2608), .Y(n2612));
OAI21X1  g0483(.A0(n2226), .A1(g45), .B0(g47), .Y(n2613_1));
XOR2X1   g0484(.A(n2613_1), .B(n2612), .Y(n1869));
XOR2X1   g0485(.A(n2494), .B(n2464), .Y(n2615));
XOR2X1   g0486(.A(n2432_1), .B(n2382_1), .Y(n2616));
XOR2X1   g0487(.A(n2616), .B(n2615), .Y(n2617));
XOR2X1   g0488(.A(n2604), .B(n2580_1), .Y(n2618_1));
XOR2X1   g0489(.A(n2553), .B(n2527), .Y(n2619));
XOR2X1   g0490(.A(n2619), .B(n2618_1), .Y(n2620));
OR2X1    g0491(.A(n2620), .B(n2617), .Y(n2621));
AOI21X1  g0492(.A0(n2620), .A1(n2617), .B0(n2226), .Y(n2622));
AOI22X1  g0493(.A0(n2621), .A1(n2622), .B0(n1869), .B1(n2226), .Y(n2623_1));
NAND2X1  g0494(.A(n2623_1), .B(g62), .Y(g9378));
INVX1    g0495(.A(g828), .Y(n2625));
NAND4X1  g0496(.A(g825), .B(g819), .C(g822), .D(g815), .Y(n2626));
NOR2X1   g0497(.A(n2626), .B(n2625), .Y(n2627));
XOR2X1   g0498(.A(n2627), .B(g786), .Y(g7763));
INVX1    g0499(.A(g929), .Y(g3856));
INVX1    g0500(.A(g955), .Y(g3857));
INVX1    g0501(.A(g795), .Y(g3854));
INVX1    g0502(.A(g154), .Y(n2632));
NOR2X1   g0503(.A(n2632), .B(g1034), .Y(n434));
INVX1    g0504(.A(g936), .Y(n2634));
NOR2X1   g0505(.A(n2634), .B(g940), .Y(n2635));
INVX1    g0506(.A(n2635), .Y(n2636));
OR2X1    g0507(.A(n2636), .B(g8), .Y(n454));
INVX1    g0508(.A(g190), .Y(n2638));
INVX1    g0509(.A(g210), .Y(n2639));
OR2X1    g0510(.A(n2639), .B(g1206), .Y(n2640));
AOI21X1  g0511(.A0(n2639), .A1(g1206), .B0(g207), .Y(n2641));
AOI21X1  g0512(.A0(n2641), .A1(n2640), .B0(n2638), .Y(n464));
INVX1    g0513(.A(g1549), .Y(n2643));
INVX1    g0514(.A(g1545), .Y(n2644));
NAND4X1  g0515(.A(g1537), .B(g1532), .C(g1541), .D(g1528), .Y(n2645));
NOR4X1   g0516(.A(n2644), .B(n2643), .C(g1251), .D(n2645), .Y(n2646));
NOR2X1   g0517(.A(n2646), .B(g1553), .Y(n2647_1));
INVX1    g0518(.A(g1541), .Y(n2648));
INVX1    g0519(.A(g1251), .Y(n2649));
NAND3X1  g0520(.A(g1528), .B(g1537), .C(g1532), .Y(n2650));
XOR2X1   g0521(.A(n2650), .B(g1541), .Y(n2651));
MX2X1    g0522(.A(n2648), .B(n2651), .S0(n2649), .Y(n2652_1));
NAND2X1  g0523(.A(n2652_1), .B(n2647_1), .Y(n469));
NAND2X1  g0524(.A(g1084), .B(g1077), .Y(n2654));
NAND3X1  g0525(.A(g1158), .B(g1176), .C(g652), .Y(n2655));
NAND2X1  g0526(.A(n2655), .B(n2654), .Y(n474));
AND2X1   g0527(.A(g959), .B(g955), .Y(n2658));
AOI21X1  g0528(.A0(n2658), .A1(g945), .B0(n2151), .Y(n479));
NOR3X1   g0529(.A(n2132), .B(n2135), .C(g6850), .Y(n484));
MX2X1    g0530(.A(g498), .B(g480), .S0(n2243), .Y(n489));
INVX1    g0531(.A(g1092), .Y(n2662_1));
INVX1    g0532(.A(g1158), .Y(n902));
NOR2X1   g0533(.A(n902), .B(g1251), .Y(n2664));
XOR2X1   g0534(.A(n2664), .B(n2662_1), .Y(n2665));
AOI21X1  g0535(.A0(g1158), .A1(g1073), .B0(n2665), .Y(n499));
INVX1    g0536(.A(g195), .Y(n2667_1));
OR2X1    g0537(.A(n2667_1), .B(g1194), .Y(n2668));
AOI21X1  g0538(.A0(n2667_1), .A1(g1194), .B0(g196), .Y(n2669));
AOI21X1  g0539(.A0(n2669), .A1(n2668), .B0(n2638), .Y(n509));
XOR2X1   g0540(.A(g1207), .B(g608), .Y(n529));
AOI22X1  g0541(.A0(g661), .A1(g633), .B0(g634), .B1(g665), .Y(n2672_1));
AOI22X1  g0542(.A0(g734), .A1(g722), .B0(g645), .B1(g673), .Y(n2673));
AOI22X1  g0543(.A0(g652), .A1(g677), .B0(g669), .B1(g635), .Y(n2674));
NAND3X1  g0544(.A(n2674), .B(n2673), .C(n2672_1), .Y(n2675));
NAND2X1  g0545(.A(g710), .B(g694), .Y(n2676));
AOI22X1  g0546(.A0(g730), .A1(g723), .B0(g698), .B1(g714), .Y(n2677_1));
AOI22X1  g0547(.A0(g685), .A1(g648), .B0(g690), .B1(g706), .Y(n2678));
AOI22X1  g0548(.A0(g718), .A1(g702), .B0(g647), .B1(g681), .Y(n2679));
NAND4X1  g0549(.A(n2678), .B(n2677_1), .C(n2676), .D(n2679), .Y(n2680));
OR2X1    g0550(.A(n2680), .B(n2675), .Y(n534));
INVX1    g0551(.A(g371), .Y(n2682_1));
NOR2X1   g0552(.A(g368), .B(n2682_1), .Y(n2683));
MX2X1    g0553(.A(g359), .B(g355), .S0(n2683), .Y(n544));
XOR2X1   g0554(.A(g1211), .B(g620), .Y(n549));
INVX1    g0555(.A(g1247), .Y(n2686));
NAND3X1  g0556(.A(g1330), .B(g1336), .C(g1333), .Y(n2687_1));
XOR2X1   g0557(.A(n2687_1), .B(g1339), .Y(n2688));
NOR2X1   g0558(.A(n2688), .B(n2686), .Y(n554));
XOR2X1   g0559(.A(g1342), .B(g628), .Y(n2690));
XOR2X1   g0560(.A(g1339), .B(g629), .Y(n2691));
XOR2X1   g0561(.A(g1345), .B(g627), .Y(n2692_1));
NOR3X1   g0562(.A(n2692_1), .B(n2691), .C(n2690), .Y(n2693));
XOR2X1   g0563(.A(g1330), .B(g632), .Y(n2694));
XOR2X1   g0564(.A(g1336), .B(g630), .Y(n2695));
XOR2X1   g0565(.A(g1348), .B(g626), .Y(n2696));
XOR2X1   g0566(.A(g1333), .B(g631), .Y(n2697_1));
NOR4X1   g0567(.A(n2696), .B(n2695), .C(n2694), .D(n2697_1), .Y(n2698));
XOR2X1   g0568(.A(g1357), .B(g623), .Y(n2699));
XOR2X1   g0569(.A(g1360), .B(g622), .Y(n2700));
XOR2X1   g0570(.A(g1354), .B(g624), .Y(n2701));
XOR2X1   g0571(.A(g1351), .B(g625), .Y(n2702_1));
NOR4X1   g0572(.A(n2701), .B(n2700), .C(n2699), .D(n2702_1), .Y(n2703));
NAND3X1  g0573(.A(n2703), .B(n2698), .C(n2693), .Y(n559));
INVX1    g0574(.A(g1260), .Y(n564));
INVX1    g0575(.A(g1110), .Y(n2706));
INVX1    g0576(.A(g1114), .Y(n2707_1));
INVX1    g0577(.A(g1118), .Y(n2708));
NAND4X1  g0578(.A(g1087), .B(g1098), .C(g1102), .D(g1106), .Y(n2709));
NOR4X1   g0579(.A(n2708), .B(n2707_1), .C(n2706), .D(n2709), .Y(n2710));
AND2X1   g0580(.A(n2710), .B(g1122), .Y(n2711));
AND2X1   g0581(.A(n2711), .B(g1126), .Y(n2712_1));
AND2X1   g0582(.A(n2712_1), .B(g1142), .Y(n1195));
OR4X1    g0583(.A(g1166), .B(g1170), .C(g1173), .D(g1167), .Y(n2714));
OR2X1    g0584(.A(n2714), .B(n1195), .Y(n579));
INVX1    g0585(.A(g1477), .Y(n2716));
INVX1    g0586(.A(g1504), .Y(n2717_1));
INVX1    g0587(.A(g1509), .Y(n2718));
INVX1    g0588(.A(g1514), .Y(n2719));
NAND4X1  g0589(.A(g1481), .B(g1489), .C(g1499), .D(g1494), .Y(n2720));
NOR4X1   g0590(.A(n2719), .B(n2718), .C(n2717_1), .D(n2720), .Y(n2721_1));
AND2X1   g0591(.A(n2721_1), .B(g1519), .Y(n2722));
NAND4X1  g0592(.A(g1462), .B(g1472), .C(g1467), .D(n2722), .Y(n2723));
XOR2X1   g0593(.A(n2723), .B(g1477), .Y(n2724));
MX2X1    g0594(.A(n2716), .B(n2724), .S0(n2649), .Y(n2725));
AND2X1   g0595(.A(n2307), .B(g150), .Y(n2726_1));
INVX1    g0596(.A(n2726_1), .Y(n2727));
AND2X1   g0597(.A(g1481), .B(g1489), .Y(n2728));
AND2X1   g0598(.A(n2728), .B(g1494), .Y(n2729));
NAND4X1  g0599(.A(g174), .B(g1504), .C(g1499), .D(g1467), .Y(n2730));
NAND4X1  g0600(.A(g1462), .B(g1472), .C(g1477), .D(g1519), .Y(n2731_1));
NOR2X1   g0601(.A(n2731_1), .B(n2730), .Y(n2732));
AND2X1   g0602(.A(n2732), .B(n2729), .Y(n2733));
INVX1    g0603(.A(g1462), .Y(n2734));
INVX1    g0604(.A(g1519), .Y(n2735));
INVX1    g0605(.A(g1467), .Y(n2736_1));
INVX1    g0606(.A(g1472), .Y(n2737));
OR4X1    g0607(.A(n2737), .B(n2736_1), .C(g174), .D(n2719), .Y(n2738));
NOR4X1   g0608(.A(n2720), .B(n2735), .C(n2734), .D(n2738), .Y(n2739));
OR2X1    g0609(.A(n2739), .B(n2733), .Y(n2740));
AOI21X1  g0610(.A0(n2307), .A1(g150), .B0(g1251), .Y(n2741_1));
AND2X1   g0611(.A(n2741_1), .B(n2740), .Y(n2742));
INVX1    g0612(.A(n2742), .Y(n2743));
INVX1    g0613(.A(g1524), .Y(n2744));
XOR2X1   g0614(.A(n2744), .B(g1513), .Y(n2745));
OAI21X1  g0615(.A0(n2745), .A1(n2727), .B0(n2743), .Y(n2746_1));
NOR2X1   g0616(.A(n2746_1), .B(n2725), .Y(n594));
OR2X1    g0617(.A(n2494), .B(g62), .Y(n2748));
OR2X1    g0618(.A(n2494), .B(n2384), .Y(n2749));
NAND2X1  g0619(.A(n2749), .B(n2748), .Y(n599));
INVX1    g0620(.A(g533), .Y(n2751_1));
NOR2X1   g0621(.A(g530), .B(n2751_1), .Y(n2752));
MX2X1    g0622(.A(g465), .B(g456), .S0(n2752), .Y(n613));
INVX1    g0623(.A(g290), .Y(n2754));
NOR2X1   g0624(.A(g287), .B(n2754), .Y(n2755));
MX2X1    g0625(.A(g243), .B(g233), .S0(n2755), .Y(n633));
INVX1    g0626(.A(n2746_1), .Y(n2757));
XOR2X1   g0627(.A(n2729), .B(g1499), .Y(n2758));
MX2X1    g0628(.A(g1499), .B(n2758), .S0(n2649), .Y(n2759));
AND2X1   g0629(.A(n2759), .B(n2757), .Y(n638));
AOI21X1  g0630(.A0(g1450), .A1(g1454), .B0(g1459), .Y(n2761_1));
NAND2X1  g0631(.A(n2761_1), .B(g1444), .Y(n648));
INVX1    g0632(.A(g1217), .Y(n2763));
INVX1    g0633(.A(g1220), .Y(n2764));
NAND4X1  g0634(.A(g1214), .B(n2764), .C(n2763), .D(g1211), .Y(n653));
MX2X1    g0635(.A(g423), .B(g405), .S0(n2351), .Y(n663));
INVX1    g0636(.A(g781), .Y(n2767));
INVX1    g0637(.A(g812), .Y(n2768));
NAND4X1  g0638(.A(g799), .B(g806), .C(g803), .D(g809), .Y(n2769));
NOR2X1   g0639(.A(n2769), .B(n2768), .Y(n2770_1));
AOI21X1  g0640(.A0(n2770_1), .A1(g775), .B0(n2767), .Y(n2771));
XOR2X1   g0641(.A(g799), .B(g803), .Y(n2772));
AND2X1   g0642(.A(n2772), .B(n2771), .Y(n673));
NOR3X1   g0643(.A(n2219_1), .B(g979), .C(g6850), .Y(n713));
MX2X1    g0644(.A(g527), .B(g521), .S0(n2243), .Y(n728));
MX2X1    g0645(.A(g278), .B(g274), .S0(n2755), .Y(n738));
XOR2X1   g0646(.A(g610), .B(g1229), .Y(n743));
NOR3X1   g0647(.A(n2278_1), .B(n2188), .C(n2205), .Y(n2778));
MX2X1    g0648(.A(g718), .B(g2), .S0(n2778), .Y(n748));
INVX1    g0649(.A(g1307), .Y(n2780));
NAND4X1  g0650(.A(g1272), .B(g1280), .C(g1276), .D(g1284), .Y(n2781));
NAND4X1  g0651(.A(g1280), .B(g1276), .C(g1296), .D(g1300), .Y(n2782));
NAND4X1  g0652(.A(g1272), .B(g1292), .C(g1288), .D(g1284), .Y(n2783_1));
OAI22X1  g0653(.A0(n2782), .A1(n2783_1), .B0(n2781), .B1(g1288), .Y(n2784));
AOI21X1  g0654(.A0(n2781), .A1(g1288), .B0(n2784), .Y(n2785));
AOI21X1  g0655(.A0(n2780), .A1(g1288), .B0(g1304), .Y(n2786));
OAI21X1  g0656(.A0(n2785), .A1(n2780), .B0(n2786), .Y(n763));
XOR2X1   g0657(.A(g1225), .B(g614), .Y(n768));
OR2X1    g0658(.A(n2382_1), .B(g62), .Y(n2789));
OR2X1    g0659(.A(n2382_1), .B(n2384), .Y(n2790));
NAND2X1  g0660(.A(n2790), .B(n2789), .Y(n783));
MX2X1    g0661(.A(g362), .B(g356), .S0(n2344), .Y(n788));
MX2X1    g0662(.A(g270), .B(g252), .S0(n2341), .Y(n798));
MX2X1    g0663(.A(g710), .B(g48), .S0(n2778), .Y(n808));
MX2X1    g0664(.A(g730), .B(g5), .S0(n2778), .Y(n813));
INVX1    g0665(.A(g1037), .Y(n2796));
INVX1    g0666(.A(g1149), .Y(n2797));
NAND4X1  g0667(.A(g1130), .B(g1138), .C(g1092), .D(g1134), .Y(n2798_1));
NOR2X1   g0668(.A(n2798_1), .B(n2797), .Y(n2799));
XOR2X1   g0669(.A(n2799), .B(n2796), .Y(n2800));
MX2X1    g0670(.A(n2796), .B(n2800), .S0(n2664), .Y(n2801));
AOI21X1  g0671(.A0(g1158), .A1(g1073), .B0(n2801), .Y(n823));
INVX1    g0672(.A(g1097), .Y(n2803_1));
AND2X1   g0673(.A(g1087), .B(g1098), .Y(n2804));
XOR2X1   g0674(.A(n2804), .B(g1102), .Y(n2805));
MX2X1    g0675(.A(g1102), .B(n2805), .S0(g1148), .Y(n2806));
AND2X1   g0676(.A(n2806), .B(n2803_1), .Y(n828));
MX2X1    g0677(.A(g483), .B(g475), .S0(n2752), .Y(n833));
XOR2X1   g0678(.A(n2770_1), .B(g775), .Y(n2809));
AND2X1   g0679(.A(n2809), .B(n2771), .Y(n838));
XOR2X1   g0680(.A(g1228), .B(g598), .Y(n848));
AND2X1   g0681(.A(g1450), .B(g1444), .Y(n2812));
XOR2X1   g0682(.A(n2812), .B(g1454), .Y(n2813_1));
AND2X1   g0683(.A(n2813_1), .B(n2761_1), .Y(n853));
INVX1    g0684(.A(g1304), .Y(n2815));
INVX1    g0685(.A(g1288), .Y(n2816));
INVX1    g0686(.A(g1292), .Y(n2817));
INVX1    g0687(.A(g1300), .Y(n2818_1));
NOR4X1   g0688(.A(n2818_1), .B(n2817), .C(n2816), .D(n2781), .Y(n2820));
XOR2X1   g0689(.A(n2820), .B(g1296), .Y(n2821));
MX2X1    g0690(.A(g1296), .B(n2821), .S0(g1307), .Y(n2822));
AND2X1   g0691(.A(n2822), .B(n2815), .Y(n858));
NAND2X1  g0692(.A(n2527), .B(n2384), .Y(n2824));
NAND2X1  g0693(.A(n2527), .B(g62), .Y(n2825));
NAND2X1  g0694(.A(n2825), .B(n2824), .Y(n863));
XOR2X1   g0695(.A(g1251), .B(g1532), .Y(n2827_1));
NOR3X1   g0696(.A(n2827_1), .B(n2646), .C(g1553), .Y(n868));
NOR3X1   g0697(.A(g45), .B(g41), .C(g42), .Y(n2829));
NAND3X1  g0698(.A(n2829), .B(n2388), .C(n2226), .Y(n2830));
OAI21X1  g0699(.A0(n2830), .A1(n2623_1), .B0(n2388), .Y(n2831));
NAND3X1  g0700(.A(n2230), .B(n2189_1), .C(g58), .Y(n2832_1));
MX2X1    g0701(.A(g3), .B(n2831), .S0(n2832_1), .Y(n878));
INVX1    g0702(.A(g13), .Y(n2834));
INVX1    g0703(.A(g1322), .Y(n2835));
INVX1    g0704(.A(g1321), .Y(n2836_1));
INVX1    g0705(.A(g1323), .Y(n2837));
NAND4X1  g0706(.A(g1319), .B(g1320), .C(g1317), .D(g1318), .Y(n2838));
NOR4X1   g0707(.A(n2837), .B(n2836_1), .C(n2835), .D(n2838), .Y(n2839));
NAND2X1  g0708(.A(g1327), .B(g1326), .Y(n2840));
NAND2X1  g0709(.A(g1325), .B(g1324), .Y(n2841_1));
NOR2X1   g0710(.A(n2841_1), .B(n2840), .Y(n2842));
NAND4X1  g0711(.A(n2839), .B(g1313), .C(g1328), .D(n2842), .Y(n2843));
AOI21X1  g0712(.A0(n2843), .A1(n2834), .B0(g1329), .Y(n883));
OR2X1    g0713(.A(g1431), .B(g1430), .Y(n2845));
AOI21X1  g0714(.A0(g1415), .A1(g1412), .B0(n2845), .Y(n907));
MX2X1    g0715(.A(g327), .B(g315), .S0(n2683), .Y(n912));
XOR2X1   g0716(.A(g1276), .B(g773), .Y(n2848));
XOR2X1   g0717(.A(g1272), .B(g774), .Y(n2849));
XOR2X1   g0718(.A(g1280), .B(g772), .Y(n2850));
XOR2X1   g0719(.A(g1284), .B(g771), .Y(n2851_1));
NOR4X1   g0720(.A(n2850), .B(n2849), .C(n2848), .D(n2851_1), .Y(n2852));
XOR2X1   g0721(.A(g769), .B(g1292), .Y(n2853));
XOR2X1   g0722(.A(g770), .B(g1288), .Y(n2854));
XOR2X1   g0723(.A(g1300), .B(g768), .Y(n2855));
XOR2X1   g0724(.A(g1296), .B(g767), .Y(n2856_1));
NOR4X1   g0725(.A(n2855), .B(n2854), .C(n2853), .D(n2856_1), .Y(n2857));
NAND2X1  g0726(.A(n2857), .B(n2852), .Y(n917));
OR4X1    g0727(.A(g1387), .B(g1386), .C(g1388), .D(g1380), .Y(n2859));
OR4X1    g0728(.A(g1383), .B(g1381), .C(g1382), .D(g1377), .Y(n2860));
OR4X1    g0729(.A(g1379), .B(g1376), .C(g1378), .D(n2860), .Y(n2861_1));
NOR4X1   g0730(.A(n2859), .B(g1385), .C(g1384), .D(n2861_1), .Y(n922));
XOR2X1   g0731(.A(g607), .B(g1211), .Y(n932));
NOR2X1   g0732(.A(g990), .B(g985), .Y(n2864));
AND2X1   g0733(.A(n2864), .B(g995), .Y(n2865));
XOR2X1   g0734(.A(n2865), .B(g985), .Y(n2866_1));
NOR2X1   g0735(.A(n2866_1), .B(g43), .Y(n947));
INVX1    g0736(.A(g1138), .Y(n2868));
NAND3X1  g0737(.A(g1134), .B(g1130), .C(g1092), .Y(n2869));
XOR2X1   g0738(.A(n2869), .B(g1138), .Y(n2870));
MX2X1    g0739(.A(n2868), .B(n2870), .S0(n2664), .Y(n2871_1));
AOI21X1  g0740(.A0(g1158), .A1(g1073), .B0(n2871_1), .Y(n977));
NOR4X1   g0741(.A(g883), .B(g896), .C(g891), .D(g901), .Y(n2873));
NOR4X1   g0742(.A(g911), .B(g906), .C(g921), .D(g916), .Y(n2874));
AOI21X1  g0743(.A0(n2874), .A1(n2873), .B0(g866), .Y(n2875));
AND2X1   g0744(.A(g933), .B(g929), .Y(n2876_1));
AND2X1   g0745(.A(n2876_1), .B(g871), .Y(n2798));
OR4X1    g0746(.A(g926), .B(g887), .C(g889), .D(g888), .Y(n2878));
NOR3X1   g0747(.A(n2878), .B(n2798), .C(n2875), .Y(n2879));
INVX1    g0748(.A(g874), .Y(n2880));
NOR4X1   g0749(.A(g888), .B(n2166), .C(n2165), .D(n2880), .Y(n2881_1));
NOR4X1   g0750(.A(g926), .B(g887), .C(n2165), .D(g888), .Y(n2882));
NAND3X1  g0751(.A(g888), .B(g887), .C(n2165), .Y(n2883));
INVX1    g0752(.A(g875), .Y(n2884));
NOR2X1   g0753(.A(g866), .B(g926), .Y(n2885));
NAND2X1  g0754(.A(n2885), .B(n2884), .Y(n2886_1));
OR4X1    g0755(.A(n2167), .B(n2166), .C(n2165), .D(n2798), .Y(n2887));
OAI21X1  g0756(.A0(n2886_1), .A1(n2883), .B0(n2887), .Y(n2888));
OR4X1    g0757(.A(n2882), .B(n2881_1), .C(n2879), .D(n2888), .Y(n987));
INVX1    g0758(.A(g452), .Y(n2890));
NOR2X1   g0759(.A(g449), .B(n2890), .Y(n2891_1));
MX2X1    g0760(.A(g390), .B(g377), .S0(n2891_1), .Y(n992));
MX2X1    g0761(.A(g417), .B(g399), .S0(n2351), .Y(n1002));
NOR3X1   g0762(.A(n2252), .B(n2188), .C(n2205), .Y(n2894));
MX2X1    g0763(.A(g681), .B(g3), .S0(n2894), .Y(n1007));
MX2X1    g0764(.A(g437), .B(g435), .S0(n2891_1), .Y(n1012));
MX2X1    g0765(.A(g351), .B(g333), .S0(n2344), .Y(n1017));
INVX1    g0766(.A(g1049), .Y(n2898));
INVX1    g0767(.A(g1041), .Y(n2899));
NOR4X1   g0768(.A(n2797), .B(n2899), .C(n2796), .D(n2798_1), .Y(n2900_1));
AND2X1   g0769(.A(n2900_1), .B(g1045), .Y(n2901));
XOR2X1   g0770(.A(n2901), .B(n2898), .Y(n2902));
MX2X1    g0771(.A(n2898), .B(n2902), .S0(n2664), .Y(n2903));
AOI21X1  g0772(.A0(g1158), .A1(g1073), .B0(n2903), .Y(n1031));
XOR2X1   g0773(.A(g1087), .B(g1098), .Y(n2905_1));
MX2X1    g0774(.A(g1098), .B(n2905_1), .S0(g1148), .Y(n2906));
AND2X1   g0775(.A(n2906), .B(n2803_1), .Y(n1036));
MX2X1    g0776(.A(g240), .B(g232), .S0(n2755), .Y(n1046));
NOR4X1   g0777(.A(g1230), .B(g1225), .C(g1224), .D(g1223), .Y(n2909));
NOR4X1   g0778(.A(g1229), .B(g1227), .C(g1226), .D(g1228), .Y(n2910_1));
NAND2X1  g0779(.A(n2910_1), .B(n2909), .Y(n1066));
MX2X1    g0780(.A(g222), .B(g213), .S0(n2755), .Y(n1071));
MX2X1    g0781(.A(g420), .B(g402), .S0(n2351), .Y(n1076));
NAND2X1  g0782(.A(n2432_1), .B(n2384), .Y(n2914));
NAND2X1  g0783(.A(n2432_1), .B(g62), .Y(n2915_1));
NAND2X1  g0784(.A(n2915_1), .B(n2914), .Y(n1081));
INVX1    g0785(.A(g45), .Y(n2917));
NAND4X1  g0786(.A(n2205), .B(n2226), .C(n2917), .D(g46), .Y(n2918));
NOR4X1   g0787(.A(n2227), .B(n2226), .C(g41), .D(n2918), .Y(n1086));
MX2X1    g0788(.A(g387), .B(g376), .S0(n2891_1), .Y(n1096));
NAND3X1  g0789(.A(n2319), .B(n2256_1), .C(n1899), .Y(n2921));
MX2X1    g0790(.A(g359), .B(g365), .S0(n2921), .Y(n1106));
XOR2X1   g0791(.A(n2742), .B(g1486), .Y(n2923));
MX2X1    g0792(.A(n2744), .B(n2923), .S0(n2727), .Y(n1111));
XOR2X1   g0793(.A(n2720), .B(g1504), .Y(n2925_1));
MX2X1    g0794(.A(n2717_1), .B(n2925_1), .S0(n2649), .Y(n2926));
NOR2X1   g0795(.A(n2926), .B(n2746_1), .Y(n1116));
XOR2X1   g0796(.A(g1214), .B(g619), .Y(n1126));
AND2X1   g0797(.A(n2627), .B(g786), .Y(n2929));
AND2X1   g0798(.A(g815), .B(g819), .Y(n2930_1));
XOR2X1   g0799(.A(n2930_1), .B(g822), .Y(n2931));
OR2X1    g0800(.A(n2931), .B(n2929), .Y(n1136));
NOR2X1   g0801(.A(g1021), .B(g1018), .Y(n2933));
XOR2X1   g0802(.A(n2933), .B(g1025), .Y(n2934));
NOR3X1   g0803(.A(g1021), .B(g1018), .C(g1025), .Y(n2935_1));
INVX1    g0804(.A(n2935_1), .Y(n2936));
AOI21X1  g0805(.A0(n2936), .A1(n2934), .B0(g1029), .Y(n2937));
OAI21X1  g0806(.A0(n2212), .A1(g1034), .B0(g43), .Y(n2938));
NOR2X1   g0807(.A(n2938), .B(n2937), .Y(n1141));
NOR3X1   g0808(.A(n2334), .B(n2206), .C(n2205), .Y(n2940_1));
MX2X1    g0809(.A(g174), .B(g5), .S0(n2940_1), .Y(n1156));
MX2X1    g0810(.A(g685), .B(g48), .S0(n2894), .Y(n1161));
XOR2X1   g0811(.A(g1148), .B(g1087), .Y(n2943));
AND2X1   g0812(.A(n2943), .B(n2803_1), .Y(n1166));
INVX1    g0813(.A(g1226), .Y(n2945));
INVX1    g0814(.A(g1207), .Y(n2946));
NAND4X1  g0815(.A(g1214), .B(g1220), .C(g1217), .D(g1211), .Y(n2947));
NAND3X1  g0816(.A(g1223), .B(g1225), .C(g1224), .Y(n2948));
NOR3X1   g0817(.A(n2948), .B(n2947), .C(n2946), .Y(n2949_1));
AOI21X1  g0818(.A0(n2949_1), .A1(n2945), .B0(g1231), .Y(n2950));
OAI21X1  g0819(.A0(n2949_1), .A1(n2945), .B0(n2950), .Y(n1180));
INVX1    g0820(.A(g1045), .Y(n2952));
XOR2X1   g0821(.A(n2900_1), .B(n2952), .Y(n2953));
MX2X1    g0822(.A(n2952), .B(n2953), .S0(n2664), .Y(n2954_1));
AOI21X1  g0823(.A0(g1158), .A1(g1073), .B0(n2954_1), .Y(n1190));
XOR2X1   g0824(.A(g605), .B(g1217), .Y(n1200));
XOR2X1   g0825(.A(g959), .B(g955), .Y(n1215));
XOR2X1   g0826(.A(g601), .B(g1225), .Y(n1220));
NAND3X1  g0827(.A(g1), .B(g10), .C(g43), .Y(n2959_1));
NOR4X1   g0828(.A(n2148), .B(g162), .C(g1034), .D(n2959_1), .Y(n1225));
MX2X1    g0829(.A(g480), .B(g474), .S0(n2752), .Y(n1240));
INVX1    g0830(.A(g1443), .Y(n2962));
INVX1    g0831(.A(g1439), .Y(n2963));
OR4X1    g0832(.A(g6675), .B(g33), .C(g38), .D(n2963), .Y(n2964_1));
AND2X1   g0833(.A(g1439), .B(g1432), .Y(n2965));
INVX1    g0834(.A(n2965), .Y(n2966));
OAI21X1  g0835(.A0(n2966), .A1(g33), .B0(g38), .Y(n2967_1));
NAND3X1  g0836(.A(n2967_1), .B(n2964_1), .C(n2962), .Y(n1255));
OR2X1    g0837(.A(n2845), .B(g1412), .Y(n1265));
INVX1    g0838(.A(g1227), .Y(n2970));
NOR4X1   g0839(.A(n2947), .B(n2946), .C(n2945), .D(n2948), .Y(n2971));
AOI21X1  g0840(.A0(n2971), .A1(n2970), .B0(g1231), .Y(n2972_1));
OAI21X1  g0841(.A0(n2971), .A1(n2970), .B0(n2972_1), .Y(n1270));
MX2X1    g0842(.A(g246), .B(g234), .S0(n2755), .Y(n1275));
NAND3X1  g0843(.A(n2319), .B(n2324), .C(n1899), .Y(n2975));
MX2X1    g0844(.A(g278), .B(g284), .S0(n2975), .Y(n1304));
MX2X1    g0845(.A(g219), .B(g212), .S0(n2755), .Y(n1314));
MX2X1    g0846(.A(g426), .B(g408), .S0(n2351), .Y(n1319));
XOR2X1   g0847(.A(g1207), .B(g621), .Y(n1324));
NAND2X1  g0848(.A(g799), .B(g803), .Y(n2980));
XOR2X1   g0849(.A(n2980), .B(g806), .Y(n2981_1));
NAND2X1  g0850(.A(n2981_1), .B(n2771), .Y(n1329));
NOR3X1   g0851(.A(g8234), .B(g146), .C(n2307), .Y(n1349));
INVX1    g0852(.A(g1252), .Y(n1359));
INVX1    g0853(.A(g1228), .Y(n2985));
INVX1    g0854(.A(g1229), .Y(n2986_1));
NAND3X1  g0855(.A(g1230), .B(n2986_1), .C(g1227), .Y(n2987));
NOR4X1   g0856(.A(n2948), .B(n2985), .C(n2945), .D(n2987), .Y(n2988));
NAND2X1  g0857(.A(n2988), .B(g1263), .Y(n1364));
MX2X1    g0858(.A(g669), .B(g5), .S0(n2894), .Y(n1369));
MX2X1    g0859(.A(g225), .B(g214), .S0(n2755), .Y(n1383));
MX2X1    g0860(.A(g281), .B(g275), .S0(n2341), .Y(n1388));
INVX1    g0861(.A(n2929), .Y(n2993));
XOR2X1   g0862(.A(g815), .B(g819), .Y(n2994));
AND2X1   g0863(.A(n2994), .B(n2993), .Y(n1393));
OR2X1    g0864(.A(n434), .B(g1236), .Y(n1398));
INVX1    g0865(.A(g1231), .Y(n2997));
NAND2X1  g0866(.A(g1211), .B(g1214), .Y(n2998));
OAI21X1  g0867(.A0(n2998), .A1(n2946), .B0(g1217), .Y(n2999));
NAND4X1  g0868(.A(g1207), .B(g1214), .C(n2763), .D(g1211), .Y(n3000_1));
NAND3X1  g0869(.A(n3000_1), .B(n2999), .C(n2997), .Y(n1412));
XOR2X1   g0870(.A(g597), .B(g1229), .Y(n1422));
NAND3X1  g0871(.A(g815), .B(g819), .C(g822), .Y(n3003));
XOR2X1   g0872(.A(n3003), .B(g825), .Y(n3004));
NAND2X1  g0873(.A(n3004), .B(n2993), .Y(n1427));
XOR2X1   g0874(.A(g1330), .B(g1333), .Y(n3006));
AND2X1   g0875(.A(n3006), .B(g1247), .Y(n1432));
NOR2X1   g0876(.A(n2720), .B(n2717_1), .Y(n3008));
XOR2X1   g0877(.A(n3008), .B(n2718), .Y(n3009));
MX2X1    g0878(.A(n2718), .B(n3009), .S0(n2649), .Y(n3010_1));
NOR2X1   g0879(.A(n3010_1), .B(n2746_1), .Y(n1452));
NOR2X1   g0880(.A(g1021), .B(g1025), .Y(n3012));
NOR3X1   g0881(.A(n3012), .B(g1018), .C(g1029), .Y(n3013));
NOR2X1   g0882(.A(n3013), .B(g1029), .Y(n3014));
NOR2X1   g0883(.A(n3014), .B(n2938), .Y(n1462));
MX2X1    g0884(.A(g588), .B(g580), .S0(n2351), .Y(n1467));
AND2X1   g0885(.A(n2722), .B(g1462), .Y(n3017));
XOR2X1   g0886(.A(n3017), .B(n2736_1), .Y(n3018));
MX2X1    g0887(.A(n2736_1), .B(n3018), .S0(n2649), .Y(n3019));
NOR2X1   g0888(.A(n3019), .B(n2746_1), .Y(n1472));
MX2X1    g0889(.A(g486), .B(g476), .S0(n2752), .Y(n1487));
MX2X1    g0890(.A(g471), .B(g458), .S0(n2752), .Y(n1492));
XOR2X1   g0891(.A(g1224), .B(g615), .Y(n1497));
MX2X1    g0892(.A(g513), .B(g495), .S0(n2243), .Y(n1505));
XOR2X1   g0893(.A(g1021), .B(g1018), .Y(n3025_1));
NOR4X1   g0894(.A(n2938), .B(n2935_1), .C(g1029), .D(n3025_1), .Y(n1520));
INVX1    g0895(.A(g1416), .Y(n3027));
NOR3X1   g0896(.A(n3027), .B(g1421), .C(g1424), .Y(n1525));
MX2X1    g0897(.A(g951), .B(g4), .S0(n2635), .Y(n1530));
NAND2X1  g0898(.A(g1220), .B(g1217), .Y(n3030_1));
NOR3X1   g0899(.A(n3030_1), .B(n2998), .C(g1207), .Y(n1535));
INVX1    g0900(.A(g595), .Y(n3032));
NOR2X1   g0901(.A(g576), .B(n3032), .Y(n3033));
MX2X1    g0902(.A(g580), .B(g579), .S0(n3033), .Y(n1540));
INVX1    g0903(.A(g1214), .Y(n3035));
NOR4X1   g0904(.A(g1211), .B(n2946), .C(n3035), .D(n3030_1), .Y(n1550));
NAND2X1  g0905(.A(n2208), .B(g45), .Y(n3037));
OAI21X1  g0906(.A0(g65), .A1(g62), .B0(g45), .Y(n3038_1));
NAND2X1  g0907(.A(n3038_1), .B(n3037), .Y(n1555));
MX2X1    g0908(.A(g402), .B(g394), .S0(n2891_1), .Y(n1560));
NOR3X1   g0909(.A(n2798_1), .B(n2797), .C(n2796), .Y(n3041));
XOR2X1   g0910(.A(n3041), .B(n2899), .Y(n3042_1));
MX2X1    g0911(.A(n2899), .B(n3042_1), .S0(n2664), .Y(n3043));
AOI21X1  g0912(.A0(g1158), .A1(g1073), .B0(n3043), .Y(n1570));
MX2X1    g0913(.A(g297), .B(g292), .S0(n2683), .Y(n1575));
MX2X1    g0914(.A(g953), .B(g3), .S0(n2635), .Y(n1580));
XOR2X1   g0915(.A(g602), .B(g1224), .Y(n1599));
XOR2X1   g0916(.A(g990), .B(g985), .Y(n3048));
AND2X1   g0917(.A(n3048), .B(g6850), .Y(n1609));
AOI21X1  g0918(.A0(n2966), .A1(g33), .B0(g1443), .Y(n3050));
OAI21X1  g0919(.A0(n2966), .A1(g33), .B0(n3050), .Y(n1619));
MX2X1    g0920(.A(g950), .B(g5), .S0(n2635), .Y(n1624));
AND2X1   g0921(.A(n2770_1), .B(g775), .Y(n3053));
NOR3X1   g0922(.A(n3053), .B(g799), .C(n2767), .Y(n1629));
XOR2X1   g0923(.A(n2769), .B(n2768), .Y(n3055));
AND2X1   g0924(.A(n3055), .B(n2771), .Y(n1634));
MX2X1    g0925(.A(g567), .B(g566), .S0(n3033), .Y(n1639));
MX2X1    g0926(.A(g333), .B(g317), .S0(n2683), .Y(n1649));
MX2X1    g0927(.A(g168), .B(g48), .S0(n2940_1), .Y(n1654));
XOR2X1   g0928(.A(n2711), .B(g1126), .Y(n3060));
MX2X1    g0929(.A(g1126), .B(n3060), .S0(g1148), .Y(n3061));
OR2X1    g0930(.A(n3061), .B(g1097), .Y(n1673));
INVX1    g0931(.A(g1329), .Y(n3063));
INVX1    g0932(.A(g1326), .Y(n3064_1));
NAND4X1  g0933(.A(g1313), .B(g1325), .C(g1324), .D(n2839), .Y(n3065));
XOR2X1   g0934(.A(n3065), .B(n3064_1), .Y(n3066));
MX2X1    g0935(.A(g103), .B(n3066), .S0(n3063), .Y(n1683));
MX2X1    g0936(.A(g309), .B(g296), .S0(n2683), .Y(n1693));
MX2X1    g0937(.A(g557), .B(g556), .S0(n3033), .Y(n1713));
XOR2X1   g0938(.A(g613), .B(g1226), .Y(n1718));
INVX1    g0939(.A(g1211), .Y(n3071));
NOR4X1   g0940(.A(n2946), .B(n3035), .C(n2763), .D(n3071), .Y(n3072));
AOI21X1  g0941(.A0(n3072), .A1(n2764), .B0(g1231), .Y(n3073_1));
OAI21X1  g0942(.A0(n3072), .A1(n2764), .B0(n3073_1), .Y(n1723));
MX2X1    g0943(.A(g158), .B(g2), .S0(n2940_1), .Y(n1728));
MX2X1    g0944(.A(g661), .B(g7), .S0(n2894), .Y(n1738));
INVX1    g0945(.A(g1313), .Y(n3077));
INVX1    g0946(.A(n2839), .Y(n3078_1));
NOR4X1   g0947(.A(n3078_1), .B(n3077), .C(n3064_1), .D(n2841_1), .Y(n3079));
XOR2X1   g0948(.A(n3079), .B(g1327), .Y(n3080));
MX2X1    g0949(.A(g98), .B(n3080), .S0(n3063), .Y(n1753));
MX2X1    g0950(.A(g150), .B(g6), .S0(n2940_1), .Y(n1772));
NAND3X1  g0951(.A(n2293_1), .B(n2263), .C(g58), .Y(n3083_1));
MX2X1    g0952(.A(g3), .B(g859), .S0(n3083_1), .Y(n1782));
MX2X1    g0953(.A(g518), .B(g516), .S0(n2752), .Y(n1792));
AND2X1   g0954(.A(n3017), .B(g1467), .Y(n3086));
XOR2X1   g0955(.A(n3086), .B(n2737), .Y(n3087));
MX2X1    g0956(.A(n2737), .B(n3087), .S0(n2649), .Y(n3088_1));
NOR2X1   g0957(.A(n3088_1), .B(n2746_1), .Y(n1797));
MX2X1    g0958(.A(g405), .B(g395), .S0(n2891_1), .Y(n1812));
INVX1    g0959(.A(g1007), .Y(n3091));
NOR4X1   g0960(.A(n3091), .B(g1016), .C(g1008), .D(n2959_1), .Y(n3092));
NOR3X1   g0961(.A(n3092), .B(n2217), .C(n2964), .Y(n3093_1));
AOI21X1  g0962(.A0(n3093_1), .A1(n2307), .B0(n2865), .Y(n1817));
MX2X1    g0963(.A(g563), .B(g557), .S0(n2351), .Y(n1836));
MX2X1    g0964(.A(g510), .B(g492), .S0(n2243), .Y(n1841));
OR2X1    g0965(.A(n2553), .B(g62), .Y(n3097));
OR2X1    g0966(.A(n2553), .B(n2384), .Y(n3098_1));
NAND2X1  g0967(.A(n3098_1), .B(n3097), .Y(n1864));
XOR2X1   g0968(.A(g1313), .B(g1317), .Y(n3100));
MX2X1    g0969(.A(g141), .B(n3100), .S0(n3063), .Y(n1874));
MX2X1    g0970(.A(g504), .B(g486), .S0(n2243), .Y(n1879));
MX2X1    g0971(.A(g665), .B(g6), .S0(n2894), .Y(n1884));
MX2X1    g0972(.A(g544), .B(g543), .S0(n3033), .Y(n1889));
XOR2X1   g0973(.A(g792), .B(g795), .Y(n1904));
MX2X1    g0974(.A(g468), .B(g457), .S0(n2752), .Y(n1909));
AOI21X1  g0975(.A0(n2627), .A1(g786), .B0(g815), .Y(n1914));
INVX1    g0976(.A(g1450), .Y(n3108_1));
NOR3X1   g0977(.A(n3108_1), .B(g1454), .C(g1444), .Y(n1919));
MX2X1    g0978(.A(g553), .B(g544), .S0(n2351), .Y(n1924));
MX2X1    g0979(.A(g501), .B(g483), .S0(n2243), .Y(n1934));
INVX1    g0980(.A(g1357), .Y(n3112));
INVX1    g0981(.A(g1354), .Y(n3113_1));
INVX1    g0982(.A(g1360), .Y(n3114));
INVX1    g0983(.A(g1342), .Y(n3115));
NAND4X1  g0984(.A(g1336), .B(g1333), .C(g1339), .D(g1330), .Y(n3116));
NOR2X1   g0985(.A(n3116), .B(n3115), .Y(n3117));
NAND4X1  g0986(.A(g1351), .B(g1348), .C(g1345), .D(n3117), .Y(n3118_1));
OR4X1    g0987(.A(n3114), .B(n3113_1), .C(n3112), .D(n3118_1), .Y(n3119));
XOR2X1   g0988(.A(n3119), .B(g1190), .Y(n3120));
NOR2X1   g0989(.A(n3120), .B(n2686), .Y(n1939));
MX2X1    g0990(.A(g318), .B(g312), .S0(n2683), .Y(n1959));
MX2X1    g0991(.A(g342), .B(g324), .S0(n2344), .Y(n1969));
INVX1    g0992(.A(g1253), .Y(n3124));
OR2X1    g0993(.A(g1257), .B(g1263), .Y(n3125));
AOI21X1  g0994(.A0(n3125), .A1(n2988), .B0(n2686), .Y(n3098));
OR2X1    g0995(.A(n3098), .B(n3124), .Y(n1974));
XOR2X1   g0996(.A(g599), .B(g1227), .Y(n1984));
AND2X1   g0997(.A(g1435), .B(g1439), .Y(n3129));
XOR2X1   g0998(.A(n3129), .B(g6675), .Y(n3130));
NOR3X1   g0999(.A(n3130), .B(n2965), .C(g1443), .Y(n1989));
NAND2X1  g1000(.A(g1158), .B(g1073), .Y(n3132_1));
AND2X1   g1001(.A(n2901), .B(g1049), .Y(n3133));
XOR2X1   g1002(.A(n3133), .B(g1053), .Y(n3134));
MX2X1    g1003(.A(g1053), .B(n3134), .S0(n2664), .Y(n3135));
AND2X1   g1004(.A(n3135), .B(n3132_1), .Y(n1994));
MX2X1    g1005(.A(g252), .B(g236), .S0(n2755), .Y(n1999));
MX2X1    g1006(.A(g330), .B(g316), .S0(n2683), .Y(n2004));
MX2X1    g1007(.A(g246), .B(g264), .S0(n2975), .Y(n2009));
NOR2X1   g1008(.A(n3118_1), .B(n3113_1), .Y(n3140));
XOR2X1   g1009(.A(n3140), .B(n3112), .Y(n3141));
NOR2X1   g1010(.A(n3141), .B(n2686), .Y(n2018));
MX2X1    g1011(.A(g243), .B(g261), .S0(n2975), .Y(n2038));
MX2X1    g1012(.A(g536), .B(g535), .S0(n3033), .Y(n2048));
INVX1    g1013(.A(n2143), .Y(n2053));
XOR2X1   g1014(.A(n3053), .B(g778), .Y(n2058));
INVX1    g1015(.A(g158), .Y(n2063));
NOR2X1   g1016(.A(n2781), .B(n2816), .Y(n3148));
XOR2X1   g1017(.A(n3148), .B(n2817), .Y(n3149));
MX2X1    g1018(.A(n2817), .B(n3149), .S0(g1307), .Y(n3150));
NOR2X1   g1019(.A(n3150), .B(g1304), .Y(n2067));
NAND3X1  g1020(.A(g1179), .B(g1158), .C(g652), .Y(n3152_1));
NAND2X1  g1021(.A(n3152_1), .B(n2654), .Y(n3153));
XOR2X1   g1022(.A(n3153), .B(g1084), .Y(n2077));
XOR2X1   g1023(.A(g1435), .B(n2963), .Y(n3155));
NOR3X1   g1024(.A(n3155), .B(n2965), .C(g1443), .Y(n2082));
XOR2X1   g1025(.A(g1272), .B(g1276), .Y(n3157_1));
MX2X1    g1026(.A(g1276), .B(n3157_1), .S0(g1307), .Y(n3158));
AND2X1   g1027(.A(n3158), .B(n2815), .Y(n2092));
MX2X1    g1028(.A(g11), .B(g12), .S0(g859), .Y(n2097));
NOR2X1   g1029(.A(g162), .B(g6850), .Y(n2101));
OR2X1    g1030(.A(n2464), .B(g62), .Y(n3162_1));
OR2X1    g1031(.A(n2464), .B(n2384), .Y(n3163));
NAND2X1  g1032(.A(n3163), .B(n3162_1), .Y(n2115));
MX2X1    g1033(.A(g560), .B(g587), .S0(n3033), .Y(n2124));
NAND3X1  g1034(.A(g1211), .B(g1214), .C(g1217), .Y(n3166));
NAND3X1  g1035(.A(g1223), .B(g1207), .C(g1220), .Y(n3167_1));
OAI21X1  g1036(.A0(n3167_1), .A1(n3166), .B0(g1224), .Y(n3168));
OR4X1    g1037(.A(n2998), .B(g1224), .C(n2763), .D(n3167_1), .Y(n3169));
NAND3X1  g1038(.A(n3169), .B(n3168), .C(n2997), .Y(n2129));
INVX1    g1039(.A(g1320), .Y(n3171));
NAND4X1  g1040(.A(g1318), .B(g1319), .C(g1317), .D(g1313), .Y(n3172_1));
XOR2X1   g1041(.A(n3172_1), .B(n3171), .Y(n3173));
MX2X1    g1042(.A(g129), .B(n3173), .S0(n3063), .Y(n2134));
MX2X1    g1043(.A(g318), .B(g336), .S0(n2921), .Y(n2149));
XOR2X1   g1044(.A(g933), .B(g929), .Y(n2154));
MX2X1    g1045(.A(g327), .B(g345), .S0(n2921), .Y(n2164));
OR2X1    g1046(.A(n2604), .B(g62), .Y(n3178));
OR2X1    g1047(.A(n2604), .B(n2384), .Y(n3179));
NAND2X1  g1048(.A(n3179), .B(n3178), .Y(n2174));
NAND2X1  g1049(.A(n2874), .B(n2873), .Y(n3181));
AOI21X1  g1050(.A0(n3181), .A1(g866), .B0(g926), .Y(n3182_1));
OR4X1    g1051(.A(g888), .B(g887), .C(g889), .D(n2798), .Y(n3183));
NOR2X1   g1052(.A(n3183), .B(n3182_1), .Y(n3184));
AND2X1   g1053(.A(g888), .B(g889), .Y(n3185));
AND2X1   g1054(.A(n2798), .B(n3185), .Y(n3186));
NAND4X1  g1055(.A(g926), .B(n2166), .C(g889), .D(n2167), .Y(n3187_1));
OAI21X1  g1056(.A0(n3186), .A1(n2166), .B0(n3187_1), .Y(n3188));
OR2X1    g1057(.A(n3188), .B(n3184), .Y(n2179));
XOR2X1   g1058(.A(n2929), .B(g789), .Y(n2184));
MX2X1    g1059(.A(g173), .B(g7), .S0(n2940_1), .Y(n2189));
MX2X1    g1060(.A(g550), .B(g540), .S0(n2351), .Y(n2194));
MX2X1    g1061(.A(g255), .B(g237), .S0(n2341), .Y(n2199));
MX2X1    g1062(.A(g948), .B(g7), .S0(n2635), .Y(n2204));
NAND3X1  g1063(.A(n2966), .B(g1435), .C(n2962), .Y(n2219));
MX2X1    g1064(.A(g48), .B(g855), .S0(n3083_1), .Y(n2237));
INVX1    g1065(.A(g1254), .Y(n3197_1));
AND2X1   g1066(.A(g1211), .B(g1207), .Y(n3198));
XOR2X1   g1067(.A(n3198), .B(n3035), .Y(n3199));
NOR3X1   g1068(.A(n3199), .B(n3197_1), .C(g1231), .Y(n2242));
XOR2X1   g1069(.A(n2709), .B(g1110), .Y(n3201_1));
MX2X1    g1070(.A(n2706), .B(n3201_1), .S0(g1148), .Y(n3202));
NAND2X1  g1071(.A(n3202), .B(n2803_1), .Y(n2247));
XOR2X1   g1072(.A(g1345), .B(g763), .Y(n3204));
XOR2X1   g1073(.A(g1348), .B(g762), .Y(n3205));
INVX1    g1074(.A(g764), .Y(n3206_1));
NOR2X1   g1075(.A(g1330), .B(g1333), .Y(n3207));
OAI21X1  g1076(.A0(n3206_1), .A1(g1342), .B0(n3207), .Y(n3208));
XOR2X1   g1077(.A(g765), .B(g1339), .Y(n3209));
NOR4X1   g1078(.A(n3208), .B(n3205), .C(n3204), .D(n3209), .Y(n3210_1));
INVX1    g1079(.A(g758), .Y(n3211));
OAI22X1  g1080(.A0(g759), .A1(n3112), .B0(n3211), .B1(g1360), .Y(n3212));
AOI21X1  g1081(.A0(g1360), .A1(n3211), .B0(n3212), .Y(n3213));
INVX1    g1082(.A(g761), .Y(n3214_1));
OAI22X1  g1083(.A0(n3214_1), .A1(g1351), .B0(n3113_1), .B1(g760), .Y(n3215));
INVX1    g1084(.A(g759), .Y(n3216));
INVX1    g1085(.A(g1351), .Y(n3217));
OAI22X1  g1086(.A0(g761), .A1(n3217), .B0(n3216), .B1(g1357), .Y(n3218));
XOR2X1   g1087(.A(g1336), .B(g766), .Y(n3219_1));
INVX1    g1088(.A(g760), .Y(n3220));
OAI22X1  g1089(.A0(g1354), .A1(n3220), .B0(n3115), .B1(g764), .Y(n3221));
NOR4X1   g1090(.A(n3219_1), .B(n3218), .C(n3215), .D(n3221), .Y(n3222));
NAND3X1  g1091(.A(n3222), .B(n3213), .C(n3210_1), .Y(n2266));
XOR2X1   g1092(.A(g1481), .B(g1489), .Y(n3224_1));
MX2X1    g1093(.A(g1489), .B(n3224_1), .S0(n2649), .Y(n3225));
AND2X1   g1094(.A(n3225), .B(n2757), .Y(n2293));
OR2X1    g1095(.A(n2623_1), .B(g62), .Y(n3227));
OR2X1    g1096(.A(n2623_1), .B(n2384), .Y(n3228));
NAND2X1  g1097(.A(n3228), .B(n3227), .Y(n2302));
NAND2X1  g1098(.A(n2988), .B(g1257), .Y(n2322));
MX2X1    g1099(.A(g1409), .B(g7063), .S0(n3027), .Y(n2332));
OR4X1    g1100(.A(n2947), .B(n2970), .C(n2945), .D(n2948), .Y(n3232));
NOR3X1   g1101(.A(n3232), .B(n2985), .C(n2946), .Y(n3233));
XOR2X1   g1102(.A(n3233), .B(n2986_1), .Y(n3234_1));
NOR3X1   g1103(.A(n3234_1), .B(n3197_1), .C(g1231), .Y(n2342));
AND2X1   g1104(.A(g792), .B(g795), .Y(n3236));
XOR2X1   g1105(.A(n3236), .B(g782), .Y(n2347));
MX2X1    g1106(.A(g237), .B(g231), .S0(n2755), .Y(n2352));
MX2X1    g1107(.A(g228), .B(g215), .S0(n2755), .Y(n2362));
MX2X1    g1108(.A(g706), .B(g8), .S0(n2894), .Y(n2367));
NOR2X1   g1109(.A(g41), .B(g42), .Y(n3241));
NAND4X1  g1110(.A(n2260), .B(g55), .C(n2917), .D(n3241), .Y(n3242));
NAND2X1  g1111(.A(n3242), .B(n2260), .Y(n3243));
MX2X1    g1112(.A(g48), .B(n3243), .S0(n2832_1), .Y(n2372));
XOR2X1   g1113(.A(n2722), .B(n2734), .Y(n3245));
MX2X1    g1114(.A(n2734), .B(n3245), .S0(n2649), .Y(n3246));
NOR2X1   g1115(.A(n3246), .B(n2746_1), .Y(n2377));
XOR2X1   g1116(.A(n2626), .B(g828), .Y(n3248_1));
AOI21X1  g1117(.A0(n2627), .A1(g786), .B0(n3248_1), .Y(n2407));
MX2X1    g1118(.A(g492), .B(g478), .S0(n2752), .Y(n2417));
OAI21X1  g1119(.A0(n2151), .A1(g943), .B0(n2636), .Y(n2427));
MX2X1    g1120(.A(g356), .B(g354), .S0(n2683), .Y(n2447));
MX2X1    g1121(.A(g952), .B(g2), .S0(n2635), .Y(n2452));
NOR2X1   g1122(.A(g1160), .B(g1186), .Y(n3254));
NOR4X1   g1123(.A(g1073), .B(g1163), .C(g1182), .D(g1179), .Y(n3255));
NAND2X1  g1124(.A(n3255), .B(n3254), .Y(n2457));
XOR2X1   g1125(.A(g1227), .B(g612), .Y(n2462));
OR2X1    g1126(.A(g1428), .B(g1429), .Y(n3258));
AOI21X1  g1127(.A0(g1408), .A1(g1405), .B0(n3258), .Y(n2470));
INVX1    g1128(.A(g1225), .Y(n3260));
NAND3X1  g1129(.A(g1224), .B(g1220), .C(g1217), .Y(n3261));
NAND4X1  g1130(.A(g1211), .B(g1207), .C(g1214), .D(g1223), .Y(n3262_1));
NOR2X1   g1131(.A(n3262_1), .B(n3261), .Y(n3263));
AOI21X1  g1132(.A0(n3263), .A1(n3260), .B0(g1231), .Y(n3264));
OAI21X1  g1133(.A0(n3263), .A1(n3260), .B0(n3264), .Y(n2481));
INVX1    g1134(.A(g1069), .Y(n3266));
INVX1    g1135(.A(g1065), .Y(n3267_1));
INVX1    g1136(.A(g1061), .Y(n3268));
NAND4X1  g1137(.A(g1057), .B(g1053), .C(g1049), .D(n2901), .Y(n3269));
NOR4X1   g1138(.A(n3268), .B(n3267_1), .C(n3266), .D(n3269), .Y(n3270));
XOR2X1   g1139(.A(n3270), .B(g1073), .Y(n3271));
MX2X1    g1140(.A(g1073), .B(n3271), .S0(n2664), .Y(n3272_1));
AND2X1   g1141(.A(n3272_1), .B(n3132_1), .Y(n2486));
AND2X1   g1142(.A(n2839), .B(g1313), .Y(n3274));
XOR2X1   g1143(.A(n3274), .B(g1324), .Y(n3275));
MX2X1    g1144(.A(g113), .B(n3275), .S0(n3063), .Y(n2491));
OR2X1    g1145(.A(n3269), .B(n3268), .Y(n3277_1));
OR2X1    g1146(.A(n3277_1), .B(n3267_1), .Y(n3278));
XOR2X1   g1147(.A(n3278), .B(g1069), .Y(n3279));
MX2X1    g1148(.A(n3266), .B(n3279), .S0(n2664), .Y(n3280));
AOI21X1  g1149(.A0(g1158), .A1(g1073), .B0(n3280), .Y(n2496));
MX2X1    g1150(.A(g443), .B(g437), .S0(n2351), .Y(n2501));
XOR2X1   g1151(.A(g1228), .B(g611), .Y(n2506));
INVX1    g1152(.A(g878), .Y(n3284));
NAND4X1  g1153(.A(g887), .B(n2165), .C(n3284), .D(n2167), .Y(n3285_1));
NAND4X1  g1154(.A(g888), .B(g887), .C(n2165), .D(n2884), .Y(n3286));
NAND4X1  g1155(.A(n2167), .B(n2166), .C(g889), .D(g866), .Y(n3287));
NAND4X1  g1156(.A(n3286), .B(n3285_1), .C(n2887), .D(n3287), .Y(n2551));
MX2X1    g1157(.A(g573), .B(g560), .S0(n2351), .Y(n2556));
MX2X1    g1158(.A(g399), .B(g393), .S0(n2891_1), .Y(n2561));
MX2X1    g1159(.A(g507), .B(g489), .S0(n2243), .Y(n2570));
MX2X1    g1160(.A(g547), .B(g536), .S0(n2351), .Y(n2575));
NAND2X1  g1161(.A(g1207), .B(n2997), .Y(n2595));
MX2X1    g1162(.A(g249), .B(g235), .S0(n2755), .Y(n2600));
OR2X1    g1163(.A(g65), .B(g58), .Y(n2605));
INVX1    g1164(.A(g942), .Y(n3296));
AOI21X1  g1165(.A0(n2634), .A1(g940), .B0(n3296), .Y(n2613));
XOR2X1   g1166(.A(n2658), .B(g945), .Y(n2628));
NOR2X1   g1167(.A(n2709), .B(n2706), .Y(n3299_1));
XOR2X1   g1168(.A(n3299_1), .B(n2707_1), .Y(n3300));
MX2X1    g1169(.A(n2707_1), .B(n3300), .S0(g1148), .Y(n3301));
NAND2X1  g1170(.A(n3301), .B(n2803_1), .Y(n2633));
MX2X1    g1171(.A(g429), .B(g411), .S0(n2351), .Y(n2642));
NAND3X1  g1172(.A(g799), .B(g806), .C(g803), .Y(n3304_1));
XOR2X1   g1173(.A(n3304_1), .B(g809), .Y(n3305));
NAND2X1  g1174(.A(n3305), .B(n2771), .Y(n2647));
OR2X1    g1175(.A(n3258), .B(g1405), .Y(n2657));
NAND2X1  g1176(.A(g1330), .B(g1333), .Y(n3308));
XOR2X1   g1177(.A(n3308), .B(g1336), .Y(n3309_1));
NOR2X1   g1178(.A(n3309_1), .B(n2686), .Y(n2662));
XOR2X1   g1179(.A(n3277_1), .B(n3267_1), .Y(n3311));
MX2X1    g1180(.A(g1065), .B(n3311), .S0(n2664), .Y(n3312));
AND2X1   g1181(.A(n3312), .B(n3132_1), .Y(n2677));
XOR2X1   g1182(.A(n2710), .B(g1122), .Y(n3314_1));
MX2X1    g1183(.A(g1122), .B(n3314_1), .S0(g1148), .Y(n3315));
OR2X1    g1184(.A(n3315), .B(g1097), .Y(n2682));
NOR2X1   g1185(.A(n3232), .B(n2946), .Y(n3317));
AOI21X1  g1186(.A0(n3317), .A1(n2985), .B0(g1231), .Y(n3318));
OAI21X1  g1187(.A0(n3317), .A1(n2985), .B0(n3318), .Y(n2687));
MX2X1    g1188(.A(g495), .B(g479), .S0(n2752), .Y(n2692));
INVX1    g1189(.A(g1319), .Y(n3321));
NAND2X1  g1190(.A(g1318), .B(g1317), .Y(n3322));
NAND3X1  g1191(.A(g1313), .B(g1321), .C(g1320), .Y(n3323));
NOR3X1   g1192(.A(n3323), .B(n3322), .C(n3321), .Y(n3324_1));
XOR2X1   g1193(.A(n3324_1), .B(g1322), .Y(n3325));
MX2X1    g1194(.A(g121), .B(n3325), .S0(n3063), .Y(n2697));
NAND4X1  g1195(.A(g1207), .B(g1229), .C(g1227), .D(g1228), .Y(n3327));
OR4X1    g1196(.A(n2948), .B(n2947), .C(n2945), .D(n3327), .Y(n3328_1));
XOR2X1   g1197(.A(n3328_1), .B(g1230), .Y(n3329));
OAI21X1  g1198(.A0(n3329), .A1(n3197_1), .B0(n2997), .Y(n2702));
AOI21X1  g1199(.A0(n3012), .A1(g1018), .B0(n2212), .Y(n3331));
AOI21X1  g1200(.A0(n3331), .A1(n3093_1), .B0(n2382), .Y(n2707));
MX2X1    g1201(.A(g249), .B(g267), .S0(n2975), .Y(n2712));
NOR4X1   g1202(.A(g1211), .B(g1207), .C(n3035), .D(n3030_1), .Y(n2736));
MX2X1    g1203(.A(g714), .B(g3), .S0(n2778), .Y(n2741));
MX2X1    g1204(.A(g734), .B(g4), .S0(n2778), .Y(n2746));
XOR2X1   g1205(.A(n2712_1), .B(g1142), .Y(n3337_1));
MX2X1    g1206(.A(g1142), .B(n3337_1), .S0(g1148), .Y(n3338));
AND2X1   g1207(.A(n3338), .B(n2803_1), .Y(n2751));
XOR2X1   g1208(.A(n3116), .B(g1342), .Y(n3340));
NOR2X1   g1209(.A(n3340), .B(n2686), .Y(n2756));
INVX1    g1210(.A(g1176), .Y(n3342));
MX2X1    g1211(.A(g1080), .B(n3342), .S0(g1081), .Y(n2766));
XOR2X1   g1212(.A(g1251), .B(g1481), .Y(n3344));
NOR2X1   g1213(.A(n3344), .B(n2746_1), .Y(n2770));
XOR2X1   g1214(.A(n3118_1), .B(g1354), .Y(n3346_1));
NOR2X1   g1215(.A(n3346_1), .B(n2686), .Y(n2788));
MX2X1    g1216(.A(g489), .B(g477), .S0(n2752), .Y(n2793));
MX2X1    g1217(.A(g591), .B(g584), .S0(n2351), .Y(n2808));
NOR2X1   g1218(.A(g1268), .B(g1269), .Y(n2818));
MX2X1    g1219(.A(g949), .B(g6), .S0(n2635), .Y(n2841));
MX2X1    g1220(.A(g408), .B(g396), .S0(n2891_1), .Y(n2851));
XOR2X1   g1221(.A(n2876_1), .B(g871), .Y(n2856));
MX2X1    g1222(.A(g146), .B(g8), .S0(n2940_1), .Y(n2866));
INVX1    g1223(.A(g205), .Y(n3355_1));
OR2X1    g1224(.A(n3355_1), .B(g1202), .Y(n3356));
AOI21X1  g1225(.A0(n3355_1), .A1(g1202), .B0(g202), .Y(n3357));
AOI21X1  g1226(.A0(n3357), .A1(n3356), .B0(n2638), .Y(n2871));
MX2X1    g1227(.A(g440), .B(g436), .S0(n2891_1), .Y(n2876));
XOR2X1   g1228(.A(n2798_1), .B(n2797), .Y(n3360_1));
MX2X1    g1229(.A(g1149), .B(n3360_1), .S0(n2664), .Y(n3361));
AND2X1   g1230(.A(n3361), .B(n3132_1), .Y(n2891));
MX2X1    g1231(.A(g570), .B(g567), .S0(n2351), .Y(n2915));
MX2X1    g1232(.A(g275), .B(g273), .S0(n2755), .Y(n2920));
MX2X1    g1233(.A(g303), .B(g294), .S0(n2683), .Y(n2925));
NAND3X1  g1234(.A(g1313), .B(g1318), .C(g1317), .Y(n3366));
XOR2X1   g1235(.A(n3366), .B(n3321), .Y(n3367));
MX2X1    g1236(.A(g133), .B(n3367), .S0(n3063), .Y(n2949));
OR2X1    g1237(.A(g866), .B(g863), .Y(n3369));
MX2X1    g1238(.A(g2), .B(n3369), .S0(n3083_1), .Y(n2954));
AOI21X1  g1239(.A0(n3071), .A1(g1207), .B0(g1231), .Y(n3371));
OAI21X1  g1240(.A0(n3071), .A1(g1207), .B0(n3371), .Y(n2959));
XOR2X1   g1241(.A(g618), .B(g1217), .Y(n2972));
NOR4X1   g1242(.A(n2166), .B(g889), .C(n3284), .D(n2167), .Y(n2977));
XOR2X1   g1243(.A(g1226), .B(g600), .Y(n2986));
INVX1    g1244(.A(g1324), .Y(n3376));
NOR3X1   g1245(.A(n3078_1), .B(n3077), .C(n3376), .Y(n3377));
XOR2X1   g1246(.A(n3377), .B(g1325), .Y(n3378));
MX2X1    g1247(.A(g108), .B(n3378), .S0(n3063), .Y(n2995));
AND2X1   g1248(.A(g1272), .B(g1276), .Y(n3380_1));
XOR2X1   g1249(.A(n3380_1), .B(g1280), .Y(n3381));
MX2X1    g1250(.A(g1280), .B(n3381), .S0(g1307), .Y(n3382));
AND2X1   g1251(.A(n3382), .B(n2815), .Y(n3000));
INVX1    g1252(.A(g1106), .Y(n3384));
NAND3X1  g1253(.A(g1087), .B(g1098), .C(g1102), .Y(n3385_1));
XOR2X1   g1254(.A(n3385_1), .B(g1106), .Y(n3386));
MX2X1    g1255(.A(n3384), .B(n3386), .S0(g1148), .Y(n3387));
NAND2X1  g1256(.A(n3387), .B(n2803_1), .Y(n3005));
XOR2X1   g1257(.A(n3269), .B(n3268), .Y(n3389));
MX2X1    g1258(.A(g1061), .B(n3389), .S0(n2664), .Y(n3390_1));
AND2X1   g1259(.A(n3390_1), .B(n3132_1), .Y(n3010));
XOR2X1   g1260(.A(g617), .B(g1220), .Y(n3015));
INVX1    g1261(.A(g1444), .Y(n3393));
INVX1    g1262(.A(g1454), .Y(n3394));
NOR3X1   g1263(.A(g1450), .B(n3394), .C(n3393), .Y(n3025));
MX2X1    g1264(.A(g378), .B(g373), .S0(n2891_1), .Y(n3030));
NOR3X1   g1265(.A(n2720), .B(n2718), .C(n2717_1), .Y(n3397));
XOR2X1   g1266(.A(n3397), .B(n2719), .Y(n3398));
MX2X1    g1267(.A(n2719), .B(n3398), .S0(n2649), .Y(n3399));
NOR2X1   g1268(.A(n3399), .B(n2746_1), .Y(n3038));
INVX1    g1269(.A(g1345), .Y(n3401));
XOR2X1   g1270(.A(n3117), .B(n3401), .Y(n3402));
NOR2X1   g1271(.A(n3402), .B(n2686), .Y(n3046));
OAI21X1  g1272(.A0(n2947), .A1(n2946), .B0(g1223), .Y(n3404_1));
OR4X1    g1273(.A(g1223), .B(n2946), .C(n2764), .D(n3166), .Y(n3405));
NAND3X1  g1274(.A(n3405), .B(n3404_1), .C(n2997), .Y(n3073));
MX2X1    g1275(.A(g446), .B(g440), .S0(n2351), .Y(n3078));
NOR2X1   g1276(.A(g1416), .B(g1421), .Y(n3408_1));
OR2X1    g1277(.A(n3408_1), .B(g1424), .Y(n3083));
MX2X1    g1278(.A(g216), .B(g211), .S0(n2755), .Y(n3103));
MX2X1    g1279(.A(g540), .B(g539), .S0(n3033), .Y(n3118));
AND2X1   g1280(.A(g1528), .B(g1532), .Y(n3412));
XOR2X1   g1281(.A(n3412), .B(g1537), .Y(n3413_1));
MX2X1    g1282(.A(g1537), .B(n3413_1), .S0(n2649), .Y(n3414));
AND2X1   g1283(.A(n3414), .B(n2647_1), .Y(n3127));
XOR2X1   g1284(.A(n2646), .B(g727), .Y(n3132));
NOR4X1   g1285(.A(n2215), .B(g1), .C(g1000), .D(n2145), .Y(n3137));
XOR2X1   g1286(.A(g1272), .B(g1307), .Y(n3418_1));
AND2X1   g1287(.A(n3418_1), .B(n2815), .Y(n3147));
NAND4X1  g1288(.A(g1325), .B(g1327), .C(g1326), .D(g1313), .Y(n3420));
NOR3X1   g1289(.A(n3420), .B(n3078_1), .C(n3376), .Y(n3421));
XOR2X1   g1290(.A(n3421), .B(g1328), .Y(n3422));
MX2X1    g1291(.A(g93), .B(n3422), .S0(n3063), .Y(n3157));
OAI21X1  g1292(.A0(n902), .A1(g1251), .B0(g1130), .Y(n3424));
XOR2X1   g1293(.A(g1130), .B(g1092), .Y(n3425));
NAND3X1  g1294(.A(n3425), .B(g1158), .C(n2649), .Y(n3426));
AOI22X1  g1295(.A0(n3424), .A1(n3426), .B0(g1158), .B1(g1073), .Y(n3162));
NOR2X1   g1296(.A(g1330), .B(n2686), .Y(n3167));
MX2X1    g1297(.A(g524), .B(g518), .S0(n2243), .Y(n3187));
XOR2X1   g1298(.A(g1230), .B(g596), .Y(n3192));
MX2X1    g1299(.A(g330), .B(g348), .S0(n2921), .Y(n3197));
INVX1    g1300(.A(g1348), .Y(n3432));
NOR3X1   g1301(.A(n3116), .B(n3401), .C(n3115), .Y(n3433_1));
XOR2X1   g1302(.A(n3433_1), .B(n3432), .Y(n3434));
NOR2X1   g1303(.A(n3434), .B(n2686), .Y(n3206));
NAND2X1  g1304(.A(n2988), .B(g1266), .Y(n3214));
NAND2X1  g1305(.A(n2580_1), .B(n2384), .Y(n3437));
NAND2X1  g1306(.A(n2580_1), .B(g62), .Y(n3438_1));
NAND2X1  g1307(.A(n3438_1), .B(n3437), .Y(n3219));
MX2X1    g1308(.A(g240), .B(g258), .S0(n2975), .Y(n3224));
MX2X1    g1309(.A(g521), .B(g517), .S0(n2752), .Y(n3229));
MX2X1    g1310(.A(g300), .B(g293), .S0(n2683), .Y(n3234));
NOR3X1   g1311(.A(n2709), .B(n2707_1), .C(n2706), .Y(n3443_1));
XOR2X1   g1312(.A(n3443_1), .B(n2708), .Y(n3444));
MX2X1    g1313(.A(n2708), .B(n3444), .S0(g1148), .Y(n3445));
NAND2X1  g1314(.A(n3445), .B(n2803_1), .Y(n3244));
AND2X1   g1315(.A(g1313), .B(g1317), .Y(n3447));
XOR2X1   g1316(.A(n3447), .B(g1318), .Y(n3448_1));
MX2X1    g1317(.A(g137), .B(n3448_1), .S0(n3063), .Y(n3252));
XOR2X1   g1318(.A(g603), .B(g1223), .Y(n3257));
MX2X1    g1319(.A(g677), .B(g2), .S0(n2894), .Y(n3262));
AND2X1   g1320(.A(n3133), .B(g1053), .Y(n3452));
XOR2X1   g1321(.A(n3452), .B(g1057), .Y(n3453_1));
MX2X1    g1322(.A(g1057), .B(n3453_1), .S0(n2664), .Y(n3454));
AND2X1   g1323(.A(n3454), .B(n3132_1), .Y(n3272));
NOR3X1   g1324(.A(n2132), .B(g1), .C(g6850), .Y(n3277));
NOR2X1   g1325(.A(n2645), .B(n2644), .Y(n3457));
XOR2X1   g1326(.A(n3457), .B(g1549), .Y(n3458_1));
MX2X1    g1327(.A(g1549), .B(n3458_1), .S0(n2649), .Y(n3459));
AND2X1   g1328(.A(n3459), .B(n2647_1), .Y(n3289));
NOR2X1   g1329(.A(n2838), .B(n3077), .Y(n3461));
XOR2X1   g1330(.A(n3461), .B(g1321), .Y(n3462));
MX2X1    g1331(.A(g125), .B(n3462), .S0(n3063), .Y(n3294));
NOR2X1   g1332(.A(n2783_1), .B(n2782), .Y(n3299));
XOR2X1   g1333(.A(n2721_1), .B(n2735), .Y(n3465));
MX2X1    g1334(.A(n2735), .B(n3465), .S0(n2649), .Y(n3466));
NOR2X1   g1335(.A(n3466), .B(n2746_1), .Y(n3304));
MX2X1    g1336(.A(g584), .B(g583), .S0(n3033), .Y(n3309));
MX2X1    g1337(.A(g324), .B(g314), .S0(n2683), .Y(n3319));
MX2X1    g1338(.A(g432), .B(g414), .S0(n2351), .Y(n3324));
MX2X1    g1339(.A(g321), .B(g313), .S0(n2683), .Y(n3333));
MX2X1    g1340(.A(g414), .B(g398), .S0(n2891_1), .Y(n3341));
XOR2X1   g1341(.A(g604), .B(g1220), .Y(n3346));
INVX1    g1342(.A(g1284), .Y(n3474));
NAND3X1  g1343(.A(g1272), .B(g1280), .C(g1276), .Y(n3475));
XOR2X1   g1344(.A(n3475), .B(g1284), .Y(n3476));
MX2X1    g1345(.A(n3474), .B(n3476), .S0(g1307), .Y(n3477_1));
NOR2X1   g1346(.A(n3477_1), .B(g1304), .Y(n3355));
XOR2X1   g1347(.A(n2645), .B(g1545), .Y(n3479));
MX2X1    g1348(.A(n2644), .B(n3479), .S0(n2649), .Y(n3480));
NAND2X1  g1349(.A(n3480), .B(n2647_1), .Y(n3360));
XOR2X1   g1350(.A(g1223), .B(g616), .Y(n3365));
MX2X1    g1351(.A(g673), .B(g4), .S0(n2894), .Y(n3370));
MX2X1    g1352(.A(g306), .B(g295), .S0(n2683), .Y(n3380));
MX2X1    g1353(.A(g954), .B(g48), .S0(n2635), .Y(n3385));
MX2X1    g1354(.A(g162), .B(g3), .S0(n2940_1), .Y(n3390));
MX2X1    g1355(.A(g411), .B(g397), .S0(n2891_1), .Y(n3395));
NOR2X1   g1356(.A(n2880), .B(g878), .Y(n3400));
NOR3X1   g1357(.A(n2781), .B(n2817), .C(n2816), .Y(n3489));
XOR2X1   g1358(.A(n3489), .B(n2818_1), .Y(n3490));
MX2X1    g1359(.A(n2818_1), .B(n3490), .S0(g1307), .Y(n3491_1));
NOR2X1   g1360(.A(n3491_1), .B(g1304), .Y(n3408));
MX2X1    g1361(.A(g384), .B(g375), .S0(n2891_1), .Y(n3413));
MX2X1    g1362(.A(g321), .B(g339), .S0(n2921), .Y(n3418));
MX2X1    g1363(.A(g459), .B(g454), .S0(n2752), .Y(n3423));
NOR4X1   g1364(.A(n3322), .B(n3321), .C(n2835), .D(n3323), .Y(n3496_1));
XOR2X1   g1365(.A(n3496_1), .B(g1323), .Y(n3497));
MX2X1    g1366(.A(g117), .B(n3497), .S0(n3063), .Y(n3428));
MX2X1    g1367(.A(g381), .B(g374), .S0(n2891_1), .Y(n3433));
XOR2X1   g1368(.A(g1528), .B(g1532), .Y(n3500));
MX2X1    g1369(.A(g1528), .B(n3500), .S0(n2649), .Y(n3501_1));
AND2X1   g1370(.A(n3501_1), .B(n2647_1), .Y(n3438));
NOR4X1   g1371(.A(n3432), .B(n3401), .C(n3115), .D(n3116), .Y(n3503));
XOR2X1   g1372(.A(n3503), .B(n3217), .Y(n3504));
NOR2X1   g1373(.A(n3504), .B(n2686), .Y(n3443));
XOR2X1   g1374(.A(g1214), .B(g606), .Y(n3453));
MX2X1    g1375(.A(n2632), .B(n2204_1), .S0(n2940_1), .Y(n3507));
NOR2X1   g1376(.A(n3507), .B(g172), .Y(n3458));
AND2X1   g1377(.A(g1130), .B(g1092), .Y(n3509_1));
XOR2X1   g1378(.A(n3509_1), .B(g1134), .Y(n3510));
MX2X1    g1379(.A(g1134), .B(n3510), .S0(n2664), .Y(n3511));
AND2X1   g1380(.A(n3511), .B(n3132_1), .Y(n3472));
AND2X1   g1381(.A(g990), .B(g985), .Y(n3513));
XOR2X1   g1382(.A(n3513), .B(g995), .Y(n3514_1));
AOI21X1  g1383(.A0(n2864), .A1(g995), .B0(n3514_1), .Y(n3515));
NOR2X1   g1384(.A(n3515), .B(g43), .Y(n3477));
MX2X1    g1385(.A(g145), .B(n3077), .S0(n3063), .Y(n3486));
XOR2X1   g1386(.A(n2728), .B(g1494), .Y(n3518));
MX2X1    g1387(.A(g1494), .B(n3518), .S0(n2649), .Y(n3519_1));
AND2X1   g1388(.A(n3519_1), .B(n2757), .Y(n3496));
MX2X1    g1389(.A(g462), .B(g455), .S0(n2752), .Y(n3501));
NOR3X1   g1390(.A(n3118_1), .B(n3113_1), .C(n3112), .Y(n3522));
XOR2X1   g1391(.A(n3522), .B(n3114), .Y(n3523_1));
NOR2X1   g1392(.A(n3523_1), .B(n2686), .Y(n3509));
XOR2X1   g1393(.A(g1450), .B(g1444), .Y(n3525));
AND2X1   g1394(.A(n3525), .B(n2761_1), .Y(n3514));
INVX1    g1395(.A(g186), .Y(n3527));
OR2X1    g1396(.A(n3527), .B(g1198), .Y(n3528_1));
AOI21X1  g1397(.A0(n3527), .A1(g1198), .B0(g187), .Y(n3529));
AOI21X1  g1398(.A0(n3529), .A1(n3528_1), .B0(n2638), .Y(n3519));
XOR2X1   g1399(.A(g1230), .B(g609), .Y(n3528));
BUFX1    g1400(.A(g1460), .Y(g206));
BUFX1    g1401(.A(g1460), .Y(g291));
BUFX1    g1402(.A(g1460), .Y(g372));
BUFX1    g1403(.A(g1460), .Y(g453));
BUFX1    g1404(.A(g1460), .Y(g534));
BUFX1    g1405(.A(g1460), .Y(g594));
BUFX1    g1406(.A(g888), .Y(g785));
BUFX1    g1407(.A(g1029), .Y(g1017));
BUFX1    g1408(.A(g1245), .Y(g1246));
BUFX1    g1409(.A(g1409), .Y(g1724));
BUFX1    g1410(.A(g891), .Y(g1783));
BUFX1    g1411(.A(g921), .Y(g1798));
BUFX1    g1412(.A(g916), .Y(g1804));
BUFX1    g1413(.A(g911), .Y(g1810));
BUFX1    g1414(.A(g906), .Y(g1817));
BUFX1    g1415(.A(g901), .Y(g1824));
BUFX1    g1416(.A(g896), .Y(g1829));
BUFX1    g1417(.A(g963), .Y(g1870));
BUFX1    g1418(.A(g966), .Y(g1871));
BUFX1    g1419(.A(g1240), .Y(g1894));
BUFX1    g1420(.A(g1524), .Y(g1911));
BUFX1    g1421(.A(g1081), .Y(g1944));
BUFX1    g1422(.A(g1254), .Y(g2662));
BUFX1    g1423(.A(g576), .Y(g2844));
BUFX1    g1424(.A(g1084), .Y(g2888));
BUFX1    g1425(.A(g1029), .Y(g3077));
BUFX1    g1426(.A(g287), .Y(g3096));
BUFX1    g1427(.A(g368), .Y(g3130));
BUFX1    g1428(.A(g449), .Y(g3159));
BUFX1    g1429(.A(g530), .Y(g3191));
BUFX1    g1430(.A(g1461), .Y(g3829));
BUFX1    g1431(.A(g1461), .Y(g3859));
BUFX1    g1432(.A(g1461), .Y(g3860));
BUFX1    g1433(.A(g1073), .Y(g4267));
BUFX1    g1434(.A(g878), .Y(g4316));
BUFX1    g1435(.A(g1160), .Y(g4370));
BUFX1    g1436(.A(g1163), .Y(g4371));
BUFX1    g1437(.A(g1182), .Y(g4372));
BUFX1    g1438(.A(g1186), .Y(g4373));
BUFX1    g1439(.A(g1554), .Y(g5143));
BUFX1    g1440(.A(g1236), .Y(g5571));
BUFX1    g1441(.A(g13), .Y(g5669));
BUFX1    g1442(.A(g16), .Y(g5678));
BUFX1    g1443(.A(g20), .Y(g5682));
BUFX1    g1444(.A(g33), .Y(g5684));
BUFX1    g1445(.A(g38), .Y(g5687));
BUFX1    g1446(.A(g49), .Y(g5729));
BUFX1    g1447(.A(g173), .Y(g6207));
BUFX1    g1448(.A(g1389), .Y(g6212));
BUFX1    g1449(.A(g1000), .Y(g6269));
BUFX1    g1450(.A(g1034), .Y(g6425));
BUFX1    g1451(.A(g1251), .Y(g6648));
BUFX1    g1452(.A(g1250), .Y(g6653));
BUFX1    g1453(.A(g1008), .Y(g6909));
OR4X1    g1454(.A(n2188), .B(n2205), .C(n2204_1), .D(n2206), .Y(g7295));
BUFX1    g1455(.A(g1167), .Y(g7423));
BUFX1    g1456(.A(g1170), .Y(g7424));
BUFX1    g1457(.A(g1173), .Y(g7425));
BUFX1    g1458(.A(g13), .Y(g7504));
BUFX1    g1459(.A(g16), .Y(g7505));
BUFX1    g1460(.A(g20), .Y(g7506));
BUFX1    g1461(.A(g33), .Y(g7507));
BUFX1    g1462(.A(g38), .Y(g7508));
BUFX1    g1463(.A(g173), .Y(g7729));
BUFX1    g1464(.A(g1389), .Y(g7730));
OR2X1    g1465(.A(g16), .B(g1189), .Y(g7731));
INVX1    g1466(.A(g1486), .Y(g7732));
BUFX1    g1467(.A(g1251), .Y(g8216));
BUFX1    g1468(.A(g1250), .Y(g8217));
BUFX1    g1469(.A(g1034), .Y(g8218));
INVX1    g1470(.A(g1432), .Y(g8219));
NAND2X1  g1471(.A(g1405), .B(g1412), .Y(g8663));
INVX1    g1472(.A(n2212), .Y(g9132));
MX2X1    g1473(.A(g31), .B(g30), .S0(g32), .Y(g9204));
BUFX1    g1474(.A(g24), .Y(g6294));
BUFX1    g1475(.A(g25), .Y(g6376));
BUFX1    g1476(.A(g29), .Y(g6300));
BUFX1    g1477(.A(g22), .Y(g6292));
BUFX1    g1478(.A(g28), .Y(g6298));
BUFX1    g1479(.A(g10), .Y(g6291));
BUFX1    g1480(.A(g23), .Y(g6293));
BUFX1    g1481(.A(g37), .Y(g6304));
BUFX1    g1482(.A(g26), .Y(g6296));
BUFX1    g1483(.A(g1), .Y(g6289));
BUFX1    g1484(.A(g27), .Y(g6297));
BUFX1    g1485(.A(g42), .Y(g6306));
BUFX1    g1486(.A(g11), .Y(g6290));
BUFX1    g1487(.A(g32), .Y(g6303));
BUFX1    g1488(.A(g41), .Y(g6305));
BUFX1    g1489(.A(g31), .Y(g6302));
BUFX1    g1490(.A(g45), .Y(g6308));
BUFX1    g1491(.A(g9), .Y(g6288));
BUFX1    g1492(.A(g44), .Y(g6307));
BUFX1    g1493(.A(g21), .Y(g6299));
BUFX1    g1494(.A(g30), .Y(g6301));
BUFX1    g1495(.A(g25), .Y(g6295));
BUFX1    g1496(.A(g1217), .Y(n429));
BUFX1    g1497(.A(g1225), .Y(n439));
BUFX1    g1498(.A(g1211), .Y(n444));
BUFX1    g1499(.A(g449), .Y(n449));
BUFX1    g1500(.A(g4), .Y(n459));
BUFX1    g1501(.A(g1223), .Y(n494));
BUFX1    g1502(.A(g1230), .Y(n504));
BUFX1    g1503(.A(g1280), .Y(n514));
BUFX1    g1504(.A(g1230), .Y(n519));
BUFX1    g1505(.A(g2), .Y(n524));
BUFX1    g1506(.A(g10), .Y(n539));
BUFX1    g1507(.A(g8), .Y(n569));
BUFX1    g1508(.A(g1225), .Y(n574));
BUFX1    g1509(.A(g1236), .Y(n584));
BUFX1    g1510(.A(g1228), .Y(n589));
BUFX1    g1511(.A(g48), .Y(n604));
BUFX1    g1512(.A(g1204), .Y(g1205));
BUFX1    g1513(.A(g48), .Y(n618));
BUFX1    g1514(.A(g916), .Y(n623));
BUFX1    g1515(.A(g1312), .Y(n628));
BUFX1    g1516(.A(g5), .Y(n643));
BUFX1    g1517(.A(g48), .Y(n658));
BUFX1    g1518(.A(g4), .Y(n668));
BUFX1    g1519(.A(g911), .Y(n678));
BUFX1    g1520(.A(g1220), .Y(n683));
BUFX1    g1521(.A(g1229), .Y(n688));
BUFX1    g1522(.A(g901), .Y(n693));
BUFX1    g1523(.A(g2), .Y(n698));
BUFX1    g1524(.A(g926), .Y(n703));
BUFX1    g1525(.A(g1012), .Y(n708));
BUFX1    g1526(.A(g114), .Y(n718));
BUFX1    g1527(.A(g134), .Y(n723));
BUFX1    g1528(.A(g1524), .Y(n733));
BUFX1    g1529(.A(g2), .Y(n753));
BUFX1    g1530(.A(g1160), .Y(n758));
BUFX1    g1531(.A(g196), .Y(n773));
BUFX1    g1532(.A(g48), .Y(n778));
BUFX1    g1533(.A(g890), .Y(n793));
BUFX1    g1534(.A(g4), .Y(n803));
BUFX1    g1535(.A(g1227), .Y(n818));
BUFX1    g1536(.A(g48), .Y(n843));
BUFX1    g1537(.A(g1284), .Y(n873));
BUFX1    g1538(.A(g2), .Y(n888));
BUFX1    g1539(.A(g43), .Y(n893));
BUFX1    g1540(.A(g8), .Y(n897));
BUFX1    g1541(.A(g168), .Y(n927));
BUFX1    g1542(.A(g1236), .Y(n937));
BUFX1    g1543(.A(g1214), .Y(n942));
BUFX1    g1544(.A(g1211), .Y(n952));
BUFX1    g1545(.A(g2), .Y(n957));
BUFX1    g1546(.A(g110), .Y(n962));
BUFX1    g1547(.A(g130), .Y(n967));
BUFX1    g1548(.A(g187), .Y(n972));
BUFX1    g1549(.A(g1308), .Y(n982));
BUFX1    g1550(.A(g8), .Y(n997));
BUFX1    g1551(.A(g1200), .Y(g1201));
BUFX1    g1552(.A(g48), .Y(n1026));
BUFX1    g1553(.A(g199), .Y(n1041));
BUFX1    g1554(.A(g1214), .Y(n1051));
BUFX1    g1555(.A(g5), .Y(n1056));
BUFX1    g1556(.A(g5), .Y(n1061));
BUFX1    g1557(.A(g1270), .Y(n1091));
BUFX1    g1558(.A(g906), .Y(n1101));
BUFX1    g1559(.A(g1155), .Y(n1121));
BUFX1    g1560(.A(g1288), .Y(n1131));
BUFX1    g1561(.A(g966), .Y(n1146));
BUFX1    g1562(.A(g7), .Y(n1151));
BUFX1    g1563(.A(g1207), .Y(n1171));
BUFX1    g1564(.A(g906), .Y(n1175));
BUFX1    g1565(.A(g2), .Y(n1185));
BUFX1    g1566(.A(g1198), .Y(n1205));
BUFX1    g1567(.A(g7), .Y(n1210));
INVX1    g1568(.A(g1260), .Y(n1230));
BUFX1    g1569(.A(g48), .Y(n1235));
BUFX1    g1570(.A(g1220), .Y(n1245));
BUFX1    g1571(.A(g3), .Y(n1250));
BUFX1    g1572(.A(g48), .Y(n1260));
BUFX1    g1573(.A(g1206), .Y(n1280));
BUFX1    g1574(.A(g1207), .Y(n1284));
BUFX1    g1575(.A(g7), .Y(n1289));
BUFX1    g1576(.A(g3), .Y(n1294));
BUFX1    g1577(.A(g1404), .Y(n1299));
BUFX1    g1578(.A(g48), .Y(n1309));
BUFX1    g1579(.A(g916), .Y(n1334));
BUFX1    g1580(.A(g1424), .Y(n1339));
BUFX1    g1581(.A(g1292), .Y(n1344));
BUFX1    g1582(.A(g8), .Y(n1354));
BUFX1    g1583(.A(g109), .Y(n1373));
BUFX1    g1584(.A(g4), .Y(n1378));
BUFX1    g1585(.A(g2), .Y(n1402));
BUFX1    g1586(.A(g3), .Y(n1407));
BUFX1    g1587(.A(g3), .Y(n1417));
BUFX1    g1588(.A(g1225), .Y(n1437));
BUFX1    g1589(.A(g1250), .Y(n1442));
BUFX1    g1590(.A(g138), .Y(n1447));
BUFX1    g1591(.A(g48), .Y(n1457));
BUFX1    g1592(.A(g1214), .Y(n1477));
BUFX1    g1593(.A(g1227), .Y(n1482));
BUFX1    g1594(.A(g1196), .Y(g1197));
BUFX1    g1595(.A(g28), .Y(n1510));
BUFX1    g1596(.A(g530), .Y(n1515));
BUFX1    g1597(.A(g7), .Y(n1545));
BUFX1    g1598(.A(g1005), .Y(n1565));
BUFX1    g1599(.A(g104), .Y(n1584));
BUFX1    g1600(.A(g142), .Y(n1589));
BUFX1    g1601(.A(g1229), .Y(n1594));
BUFX1    g1602(.A(g1224), .Y(n1604));
BUFX1    g1603(.A(g1224), .Y(n1614));
BUFX1    g1604(.A(g1224), .Y(n1644));
BUFX1    g1605(.A(g1227), .Y(n1659));
BUFX1    g1606(.A(g1220), .Y(n1664));
BUFX1    g1607(.A(g646), .Y(n1668));
BUFX1    g1608(.A(g29), .Y(n1678));
BUFX1    g1609(.A(g5), .Y(n1688));
BUFX1    g1610(.A(g1230), .Y(n1698));
BUFX1    g1611(.A(g896), .Y(n1703));
BUFX1    g1612(.A(g1225), .Y(n1708));
BUFX1    g1613(.A(g6), .Y(n1733));
BUFX1    g1614(.A(g4), .Y(n1743));
BUFX1    g1615(.A(g891), .Y(n1748));
BUFX1    g1616(.A(g1229), .Y(n1758));
BUFX1    g1617(.A(g1084), .Y(n1763));
BUFX1    g1618(.A(g92), .Y(n1767));
BUFX1    g1619(.A(g3), .Y(n1777));
BUFX1    g1620(.A(g1234), .Y(n1787));
INVX1    g1621(.A(g1252), .Y(n1802));
BUFX1    g1622(.A(g1207), .Y(n1807));
BUFX1    g1623(.A(g1146), .Y(n1821));
BUFX1    g1624(.A(g1229), .Y(n1826));
BUFX1    g1625(.A(g95), .Y(n1831));
BUFX1    g1626(.A(g1202), .Y(n1846));
BUFX1    g1627(.A(g1226), .Y(n1850));
BUFX1    g1628(.A(g1217), .Y(n1855));
BUFX1    g1629(.A(g1014), .Y(n1859));
BUFX1    g1630(.A(g368), .Y(n1894));
BUFX1    g1631(.A(g3), .Y(n1929));
BUFX1    g1632(.A(g1251), .Y(n1944));
BUFX1    g1633(.A(g2), .Y(n1949));
BUFX1    g1634(.A(g1081), .Y(n1954));
BUFX1    g1635(.A(g1226), .Y(n1964));
BUFX1    g1636(.A(g1073), .Y(n1979));
BUFX1    g1637(.A(g1156), .Y(n2013));
BUFX1    g1638(.A(g1228), .Y(n2023));
BUFX1    g1639(.A(g48), .Y(n2028));
BUFX1    g1640(.A(g883), .Y(n2033));
BUFX1    g1641(.A(g1211), .Y(n2043));
BUFX1    g1642(.A(g287), .Y(n2072));
BUFX1    g1643(.A(g5), .Y(n2087));
BUFX1    g1644(.A(g1403), .Y(n2106));
BUFX1    g1645(.A(g89), .Y(n2110));
BUFX1    g1646(.A(g1194), .Y(n2120));
BUFX1    g1647(.A(g5), .Y(n2139));
BUFX1    g1648(.A(g1217), .Y(n2144));
BUFX1    g1649(.A(g1228), .Y(n2159));
BUFX1    g1650(.A(g5), .Y(n2169));
BUFX1    g1651(.A(g1231), .Y(n2209));
BUFX1    g1652(.A(g3), .Y(n2214));
BUFX1    g1653(.A(g1220), .Y(n2224));
BUFX1    g1654(.A(g878), .Y(n2228));
BUFX1    g1655(.A(g1198), .Y(n2233));
BUFX1    g1656(.A(g1309), .Y(n2251));
BUFX1    g1657(.A(g1226), .Y(n2256));
BUFX1    g1658(.A(g979), .Y(n2261));
BUFX1    g1659(.A(g1240), .Y(n2270));
BUFX1    g1660(.A(g891), .Y(n2273));
BUFX1    g1661(.A(g48), .Y(n2278));
BUFX1    g1662(.A(g1300), .Y(n2283));
BUFX1    g1663(.A(g27), .Y(n2288));
BUFX1    g1664(.A(g921), .Y(n2297));
BUFX1    g1665(.A(g5), .Y(n2312));
BUFX1    g1666(.A(g100), .Y(n2317));
BUFX1    g1667(.A(g1296), .Y(n2327));
BUFX1    g1668(.A(g7), .Y(n2337));
BUFX1    g1669(.A(g941), .Y(n2357));
BUFX1    g1670(.A(g126), .Y(n2387));
BUFX1    g1671(.A(g901), .Y(n2392));
BUFX1    g1672(.A(g3), .Y(n2397));
BUFX1    g1673(.A(g1191), .Y(n2402));
BUFX1    g1674(.A(g26), .Y(n2412));
BUFX1    g1675(.A(g94), .Y(n2422));
BUFX1    g1676(.A(g1194), .Y(n2432));
BUFX1    g1677(.A(g1243), .Y(n2437));
BUFX1    g1678(.A(g1260), .Y(n2442));
BUFX1    g1679(.A(g1004), .Y(n2466));
BUFX1    g1680(.A(g896), .Y(n2474));
BUFX1    g1681(.A(g1271), .Y(n2477));
BUFX1    g1682(.A(g1226), .Y(n2511));
BUFX1    g1683(.A(g4), .Y(n2516));
BUFX1    g1684(.A(g7), .Y(n2521));
BUFX1    g1685(.A(g1228), .Y(n2526));
BUFX1    g1686(.A(g1223), .Y(n2531));
BUFX1    g1687(.A(g24), .Y(n2536));
OR2X1    g1688(.A(g16), .B(g1189), .Y(n2541));
BUFX1    g1689(.A(g6), .Y(n2546));
BUFX1    g1690(.A(g1244), .Y(n2565));
BUFX1    g1691(.A(g105), .Y(n2580));
BUFX1    g1692(.A(g4), .Y(n2585));
BUFX1    g1693(.A(g2), .Y(n2590));
BUFX1    g1694(.A(g911), .Y(n2609));
BUFX1    g1695(.A(g1217), .Y(n2618));
BUFX1    g1696(.A(g5), .Y(n2623));
BUFX1    g1697(.A(g99), .Y(n2637));
BUFX1    g1698(.A(g921), .Y(n2652));
BUFX1    g1699(.A(g8), .Y(n2667));
BUFX1    g1700(.A(g6), .Y(n2672));
BUFX1    g1701(.A(g23), .Y(g1195));
BUFX1    g1702(.A(g1393), .Y(n2721));
BUFX1    g1703(.A(g1230), .Y(n2726));
BUFX1    g1704(.A(g1207), .Y(n2731));
BUFX1    g1705(.A(g6), .Y(n2761));
BUFX1    g1706(.A(g1185), .Y(n2774));
BUFX1    g1707(.A(g1272), .Y(n2779));
BUFX1    g1708(.A(g1153), .Y(n2783));
BUFX1    g1709(.A(g118), .Y(n2803));
BUFX1    g1710(.A(g6), .Y(n2813));
BUFX1    g1711(.A(g1311), .Y(n2823));
BUFX1    g1712(.A(g4), .Y(n2827));
BUFX1    g1713(.A(g207), .Y(n2832));
BUFX1    g1714(.A(g1399), .Y(n2836));
BUFX1    g1715(.A(g1267), .Y(n2846));
BUFX1    g1716(.A(g8), .Y(n2861));
BUFX1    g1717(.A(g1223), .Y(n2881));
BUFX1    g1718(.A(g1), .Y(n2886));
BUFX1    g1719(.A(g1396), .Y(n2895));
BUFX1    g1720(.A(g1206), .Y(n2900));
BUFX1    g1721(.A(g1224), .Y(n2905));
BUFX1    g1722(.A(g7), .Y(n2910));
BUFX1    g1723(.A(g122), .Y(n2930));
BUFX1    g1724(.A(g202), .Y(n2935));
BUFX1    g1725(.A(g37), .Y(n2940));
BUFX1    g1726(.A(g576), .Y(n2944));
BUFX1    g1727(.A(g1182), .Y(n2967));
BUFX1    g1728(.A(g1173), .Y(n2981));
BUFX1    g1729(.A(g200), .Y(n2990));
BUFX1    g1730(.A(g5), .Y(n3020));
BUFX1    g1731(.A(g1199), .Y(n3034));
BUFX1    g1732(.A(g1402), .Y(n3042));
BUFX1    g1733(.A(g22), .Y(n3051));
BUFX1    g1734(.A(g1390), .Y(n3054));
BUFX1    g1735(.A(g1034), .Y(n3059));
INVX1    g1736(.A(g1260), .Y(n3064));
BUFX1    g1737(.A(g1157), .Y(n3068));
BUFX1    g1738(.A(g1223), .Y(n3088));
BUFX1    g1739(.A(g2), .Y(n3093));
BUFX1    g1740(.A(g1214), .Y(n3108));
BUFX1    g1741(.A(g1202), .Y(n3113));
BUFX1    g1742(.A(g1206), .Y(n3123));
BUFX1    g1743(.A(g6), .Y(n3142));
BUFX1    g1744(.A(g1240), .Y(n3152));
BUFX1    g1745(.A(g8), .Y(n3172));
BUFX1    g1746(.A(g2), .Y(n3177));
BUFX1    g1747(.A(g1167), .Y(n3182));
BUFX1    g1748(.A(g1147), .Y(n3201));
BUFX1    g1749(.A(g1154), .Y(n3210));
BUFX1    g1750(.A(g3), .Y(n3239));
BUFX1    g1751(.A(g1170), .Y(n3248));
BUFX1    g1752(.A(g1227), .Y(n3267));
BUFX1    g1753(.A(g1192), .Y(g1193));
BUFX1    g1754(.A(g16), .Y(n3285));
BUFX1    g1755(.A(g1276), .Y(n3314));
BUFX1    g1756(.A(g1159), .Y(n3328));
BUFX1    g1757(.A(g1310), .Y(n3337));
BUFX1    g1758(.A(g4), .Y(n3351));
BUFX1    g1759(.A(g3), .Y(n3375));
BUFX1    g1760(.A(g1203), .Y(n3404));
BUFX1    g1761(.A(g4), .Y(n3448));
BUFX1    g1762(.A(g1211), .Y(n3463));
BUFX1    g1763(.A(g963), .Y(n3467));
BUFX1    g1764(.A(g201), .Y(n3481));
BUFX1    g1765(.A(g6), .Y(n3491));
BUFX1    g1766(.A(g1163), .Y(n3505));
BUFX1    g1767(.A(g1186), .Y(n3523));
NAND2X1  g1768(.A(g944), .B(n2185), .Y(n3533));
BUFX1    g1769(.A(g3), .Y(n3538));
endmodule
