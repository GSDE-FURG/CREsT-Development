// Benchmark "b12_C" written by ABC on Wed Aug 05 14:40:08 2020

module b12_C ( 
    GAMMA_REG_0__SCAN_IN, START, K_3_, K_2_, K_1_, K_0_,
    COUNT_REG_0__SCAN_IN, MEMORY_REG_31__1__SCAN_IN,
    MEMORY_REG_31__0__SCAN_IN, MEMORY_REG_30__1__SCAN_IN,
    MEMORY_REG_30__0__SCAN_IN, MEMORY_REG_29__1__SCAN_IN,
    MEMORY_REG_29__0__SCAN_IN, MEMORY_REG_28__1__SCAN_IN,
    MEMORY_REG_28__0__SCAN_IN, MEMORY_REG_27__1__SCAN_IN,
    MEMORY_REG_27__0__SCAN_IN, MEMORY_REG_26__1__SCAN_IN,
    MEMORY_REG_26__0__SCAN_IN, MEMORY_REG_25__1__SCAN_IN,
    MEMORY_REG_25__0__SCAN_IN, MEMORY_REG_24__1__SCAN_IN,
    MEMORY_REG_24__0__SCAN_IN, MEMORY_REG_23__1__SCAN_IN,
    MEMORY_REG_23__0__SCAN_IN, MEMORY_REG_22__1__SCAN_IN,
    MEMORY_REG_22__0__SCAN_IN, MEMORY_REG_21__1__SCAN_IN,
    MEMORY_REG_21__0__SCAN_IN, MEMORY_REG_20__1__SCAN_IN,
    MEMORY_REG_20__0__SCAN_IN, MEMORY_REG_19__1__SCAN_IN,
    MEMORY_REG_19__0__SCAN_IN, MEMORY_REG_18__1__SCAN_IN,
    MEMORY_REG_18__0__SCAN_IN, MEMORY_REG_17__1__SCAN_IN,
    MEMORY_REG_17__0__SCAN_IN, MEMORY_REG_16__1__SCAN_IN,
    MEMORY_REG_16__0__SCAN_IN, MEMORY_REG_15__1__SCAN_IN,
    MEMORY_REG_15__0__SCAN_IN, MEMORY_REG_14__1__SCAN_IN,
    MEMORY_REG_14__0__SCAN_IN, MEMORY_REG_13__1__SCAN_IN,
    MEMORY_REG_13__0__SCAN_IN, MEMORY_REG_12__1__SCAN_IN,
    MEMORY_REG_12__0__SCAN_IN, MEMORY_REG_11__1__SCAN_IN,
    MEMORY_REG_11__0__SCAN_IN, MEMORY_REG_10__1__SCAN_IN,
    MEMORY_REG_10__0__SCAN_IN, MEMORY_REG_9__1__SCAN_IN,
    MEMORY_REG_9__0__SCAN_IN, MEMORY_REG_8__1__SCAN_IN,
    MEMORY_REG_8__0__SCAN_IN, MEMORY_REG_7__1__SCAN_IN,
    MEMORY_REG_7__0__SCAN_IN, MEMORY_REG_6__1__SCAN_IN,
    MEMORY_REG_6__0__SCAN_IN, MEMORY_REG_5__1__SCAN_IN,
    MEMORY_REG_5__0__SCAN_IN, MEMORY_REG_4__1__SCAN_IN,
    MEMORY_REG_4__0__SCAN_IN, MEMORY_REG_3__1__SCAN_IN,
    MEMORY_REG_3__0__SCAN_IN, MEMORY_REG_2__1__SCAN_IN,
    MEMORY_REG_2__0__SCAN_IN, MEMORY_REG_1__1__SCAN_IN,
    MEMORY_REG_1__0__SCAN_IN, MEMORY_REG_0__1__SCAN_IN,
    MEMORY_REG_0__0__SCAN_IN, NL_REG_3__SCAN_IN, NL_REG_2__SCAN_IN,
    NL_REG_1__SCAN_IN, NL_REG_0__SCAN_IN, SCAN_REG_4__SCAN_IN,
    SCAN_REG_3__SCAN_IN, SCAN_REG_2__SCAN_IN, SCAN_REG_1__SCAN_IN,
    SCAN_REG_0__SCAN_IN, MAX_REG_4__SCAN_IN, MAX_REG_3__SCAN_IN,
    MAX_REG_2__SCAN_IN, MAX_REG_1__SCAN_IN, MAX_REG_0__SCAN_IN,
    IND_REG_1__SCAN_IN, IND_REG_0__SCAN_IN, TIMEBASE_REG_5__SCAN_IN,
    TIMEBASE_REG_4__SCAN_IN, TIMEBASE_REG_3__SCAN_IN,
    TIMEBASE_REG_2__SCAN_IN, TIMEBASE_REG_1__SCAN_IN,
    TIMEBASE_REG_0__SCAN_IN, COUNT_REG2_5__SCAN_IN, COUNT_REG2_4__SCAN_IN,
    COUNT_REG2_3__SCAN_IN, COUNT_REG2_2__SCAN_IN, COUNT_REG2_1__SCAN_IN,
    COUNT_REG2_0__SCAN_IN, SOUND_REG_2__SCAN_IN, SOUND_REG_1__SCAN_IN,
    SOUND_REG_0__SCAN_IN, ADDRESS_REG_4__SCAN_IN, ADDRESS_REG_3__SCAN_IN,
    ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN,
    DATA_IN_REG_1__SCAN_IN, DATA_IN_REG_0__SCAN_IN, S_REG_SCAN_IN,
    PLAY_REG_SCAN_IN, NLOSS_REG_SCAN_IN, SPEAKER_REG_SCAN_IN,
    WR_REG_SCAN_IN, COUNTER_REG_2__SCAN_IN, COUNTER_REG_1__SCAN_IN,
    COUNTER_REG_0__SCAN_IN, COUNT_REG_1__SCAN_IN, NUM_REG_1__SCAN_IN,
    NUM_REG_0__SCAN_IN, DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN,
    GAMMA_REG_4__SCAN_IN, GAMMA_REG_3__SCAN_IN, GAMMA_REG_2__SCAN_IN,
    GAMMA_REG_1__SCAN_IN,
    U1391, U1486, U1485, U1484, U1483, U1482, U1481, U1480, U1479, U1478,
    U1477, U1476, U1475, U1474, U1473, U1472, U1471, U1470, U1469, U1468,
    U1467, U1466, U1465, U1464, U1463, U1462, U1461, U1460, U1459, U1458,
    U1457, U1456, U1455, U1454, U1453, U1452, U1451, U1450, U1449, U1448,
    U1447, U1446, U1445, U1444, U1443, U1442, U1441, U1440, U1439, U1438,
    U1437, U1436, U1435, U1434, U1433, U1432, U1431, U1430, U1429, U1428,
    U1427, U1426, U1425, U1424, U1423, U1422, U1421, U1420, U1419, U1418,
    U1417, U1416, U1415, U1414, U1413, U1412, U1411, U1410, U1409, U1564,
    U1565, U1566, U1408, U1407, U1406, U1405, U1567, U1404, U1403, U1568,
    U1402, U1401, U1400, U1569, U1570, U1571, U1399, U1398, U1397, U1396,
    U1395, U1572, U1573, U1394, U1574, U1575, U1393, U1392, U1381, U1382,
    U1383, U1563, U1563, U1391, U1390, U1389, U1384, U1385, U1386, U1387,
    U1388  );
  input  GAMMA_REG_0__SCAN_IN, START, K_3_, K_2_, K_1_, K_0_,
    COUNT_REG_0__SCAN_IN, MEMORY_REG_31__1__SCAN_IN,
    MEMORY_REG_31__0__SCAN_IN, MEMORY_REG_30__1__SCAN_IN,
    MEMORY_REG_30__0__SCAN_IN, MEMORY_REG_29__1__SCAN_IN,
    MEMORY_REG_29__0__SCAN_IN, MEMORY_REG_28__1__SCAN_IN,
    MEMORY_REG_28__0__SCAN_IN, MEMORY_REG_27__1__SCAN_IN,
    MEMORY_REG_27__0__SCAN_IN, MEMORY_REG_26__1__SCAN_IN,
    MEMORY_REG_26__0__SCAN_IN, MEMORY_REG_25__1__SCAN_IN,
    MEMORY_REG_25__0__SCAN_IN, MEMORY_REG_24__1__SCAN_IN,
    MEMORY_REG_24__0__SCAN_IN, MEMORY_REG_23__1__SCAN_IN,
    MEMORY_REG_23__0__SCAN_IN, MEMORY_REG_22__1__SCAN_IN,
    MEMORY_REG_22__0__SCAN_IN, MEMORY_REG_21__1__SCAN_IN,
    MEMORY_REG_21__0__SCAN_IN, MEMORY_REG_20__1__SCAN_IN,
    MEMORY_REG_20__0__SCAN_IN, MEMORY_REG_19__1__SCAN_IN,
    MEMORY_REG_19__0__SCAN_IN, MEMORY_REG_18__1__SCAN_IN,
    MEMORY_REG_18__0__SCAN_IN, MEMORY_REG_17__1__SCAN_IN,
    MEMORY_REG_17__0__SCAN_IN, MEMORY_REG_16__1__SCAN_IN,
    MEMORY_REG_16__0__SCAN_IN, MEMORY_REG_15__1__SCAN_IN,
    MEMORY_REG_15__0__SCAN_IN, MEMORY_REG_14__1__SCAN_IN,
    MEMORY_REG_14__0__SCAN_IN, MEMORY_REG_13__1__SCAN_IN,
    MEMORY_REG_13__0__SCAN_IN, MEMORY_REG_12__1__SCAN_IN,
    MEMORY_REG_12__0__SCAN_IN, MEMORY_REG_11__1__SCAN_IN,
    MEMORY_REG_11__0__SCAN_IN, MEMORY_REG_10__1__SCAN_IN,
    MEMORY_REG_10__0__SCAN_IN, MEMORY_REG_9__1__SCAN_IN,
    MEMORY_REG_9__0__SCAN_IN, MEMORY_REG_8__1__SCAN_IN,
    MEMORY_REG_8__0__SCAN_IN, MEMORY_REG_7__1__SCAN_IN,
    MEMORY_REG_7__0__SCAN_IN, MEMORY_REG_6__1__SCAN_IN,
    MEMORY_REG_6__0__SCAN_IN, MEMORY_REG_5__1__SCAN_IN,
    MEMORY_REG_5__0__SCAN_IN, MEMORY_REG_4__1__SCAN_IN,
    MEMORY_REG_4__0__SCAN_IN, MEMORY_REG_3__1__SCAN_IN,
    MEMORY_REG_3__0__SCAN_IN, MEMORY_REG_2__1__SCAN_IN,
    MEMORY_REG_2__0__SCAN_IN, MEMORY_REG_1__1__SCAN_IN,
    MEMORY_REG_1__0__SCAN_IN, MEMORY_REG_0__1__SCAN_IN,
    MEMORY_REG_0__0__SCAN_IN, NL_REG_3__SCAN_IN, NL_REG_2__SCAN_IN,
    NL_REG_1__SCAN_IN, NL_REG_0__SCAN_IN, SCAN_REG_4__SCAN_IN,
    SCAN_REG_3__SCAN_IN, SCAN_REG_2__SCAN_IN, SCAN_REG_1__SCAN_IN,
    SCAN_REG_0__SCAN_IN, MAX_REG_4__SCAN_IN, MAX_REG_3__SCAN_IN,
    MAX_REG_2__SCAN_IN, MAX_REG_1__SCAN_IN, MAX_REG_0__SCAN_IN,
    IND_REG_1__SCAN_IN, IND_REG_0__SCAN_IN, TIMEBASE_REG_5__SCAN_IN,
    TIMEBASE_REG_4__SCAN_IN, TIMEBASE_REG_3__SCAN_IN,
    TIMEBASE_REG_2__SCAN_IN, TIMEBASE_REG_1__SCAN_IN,
    TIMEBASE_REG_0__SCAN_IN, COUNT_REG2_5__SCAN_IN, COUNT_REG2_4__SCAN_IN,
    COUNT_REG2_3__SCAN_IN, COUNT_REG2_2__SCAN_IN, COUNT_REG2_1__SCAN_IN,
    COUNT_REG2_0__SCAN_IN, SOUND_REG_2__SCAN_IN, SOUND_REG_1__SCAN_IN,
    SOUND_REG_0__SCAN_IN, ADDRESS_REG_4__SCAN_IN, ADDRESS_REG_3__SCAN_IN,
    ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN,
    DATA_IN_REG_1__SCAN_IN, DATA_IN_REG_0__SCAN_IN, S_REG_SCAN_IN,
    PLAY_REG_SCAN_IN, NLOSS_REG_SCAN_IN, SPEAKER_REG_SCAN_IN,
    WR_REG_SCAN_IN, COUNTER_REG_2__SCAN_IN, COUNTER_REG_1__SCAN_IN,
    COUNTER_REG_0__SCAN_IN, COUNT_REG_1__SCAN_IN, NUM_REG_1__SCAN_IN,
    NUM_REG_0__SCAN_IN, DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN,
    GAMMA_REG_4__SCAN_IN, GAMMA_REG_3__SCAN_IN, GAMMA_REG_2__SCAN_IN,
    GAMMA_REG_1__SCAN_IN;
  output U1391, U1486, U1485, U1484, U1483, U1482, U1481, U1480, U1479, U1478,
    U1477, U1476, U1475, U1474, U1473, U1472, U1471, U1470, U1469, U1468,
    U1467, U1466, U1465, U1464, U1463, U1462, U1461, U1460, U1459, U1458,
    U1457, U1456, U1455, U1454, U1453, U1452, U1451, U1450, U1449, U1448,
    U1447, U1446, U1445, U1444, U1443, U1442, U1441, U1440, U1439, U1438,
    U1437, U1436, U1435, U1434, U1433, U1432, U1431, U1430, U1429, U1428,
    U1427, U1426, U1425, U1424, U1423, U1422, U1421, U1420, U1419, U1418,
    U1417, U1416, U1415, U1414, U1413, U1412, U1411, U1410, U1409, U1564,
    U1565, U1566, U1408, U1407, U1406, U1405, U1567, U1404, U1403, U1568,
    U1402, U1401, U1400, U1569, U1570, U1571, U1399, U1398, U1397, U1396,
    U1395, U1572, U1573, U1394, U1574, U1575, U1393, U1392, U1381, U1382,
    U1383, U1563, U1563, U1391, U1390, U1389, U1384, U1385, U1386, U1387,
    U1388;
  wire n254, n255, n256, n257, n258, n259, n260, n261, n263, n264, n266,
    n267, n268, n269, n271, n273, n274, n275, n276, n278, n280, n281, n282,
    n284, n286, n287, n288, n289, n291, n293, n294, n295, n296, n298, n300,
    n301, n302, n304, n306, n307, n308, n310, n312, n313, n314, n315, n317,
    n319, n320, n321, n323, n325, n326, n327, n329, n331, n332, n333, n335,
    n337, n338, n339, n341, n343, n344, n345, n347, n349, n350, n351, n353,
    n355, n356, n357, n359, n361, n362, n363, n364, n366, n368, n369, n370,
    n372, n374, n375, n376, n378, n380, n381, n382, n384, n386, n387, n388,
    n390, n392, n393, n394, n396, n398, n399, n400, n402, n404, n405, n406,
    n408, n410, n411, n412, n414, n416, n417, n418, n420, n422, n423, n424,
    n426, n428, n429, n430, n432, n434, n435, n436, n438, n440, n441, n442,
    n444, n446, n447, n448, n450, n452, n453, n454, n456, n458, n459, n460,
    n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
    n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
    n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
    n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
    n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
    n521, n522, n523, n524, n525, n526, n528, n529, n530, n531, n533, n534,
    n535, n536, n537, n539, n540, n541, n542, n543, n545, n546, n547, n548,
    n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
    n562, n563, n564, n565, n566, n567, n568, n570, n571, n572, n574, n575,
    n576, n578, n579, n581, n583, n584, n585, n586, n587, n588, n589, n590,
    n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
    n603, n604, n605, n606, n608, n609, n610, n611, n613, n614, n616, n618,
    n620, n621, n622, n623, n624, n625, n627, n628, n629, n631, n632, n633,
    n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
    n646, n648, n649, n650, n652, n653, n654, n655, n657, n658, n659, n661,
    n662, n663, n664, n665, n666, n668, n669, n671, n672, n673, n674, n675,
    n676, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
    n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
    n701, n702, n703, n704, n705, n706, n707, n708, n710, n711, n712, n713,
    n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n726,
    n727, n728, n729, n730, n731, n732, n734, n735, n736, n738, n739, n740,
    n742, n743, n744, n746, n747, n748, n749, n750, n751, n752, n753, n755,
    n756, n758, n759, n760, n762, n763, n764, n765, n766, n767, n768, n770,
    n772, n774, n776, n777, n779, n780, n782, n783, n785, n786, n787, n788,
    n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
    n801, n802, n803, n804, n806, n807, n808, n809, n810, n811, n812, n813,
    n814, n815, n816, n817, n818, n819, n820, n822, n823, n824, n825, n826,
    n827, n828, n829, n830, n831, n832, n833, n834, n836, n838, n840, n841,
    n843, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
    n858, n859, n860, n861, n862, n863, n864, n865, n866, n868, n869, n870,
    n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
    n883, n884, n885, n886, n887, n889, n890, n892, n893, n894, n895, n896,
    n897, n898, n899, n900, n901, n902, n904, n905, n906, n907, n908, n909,
    n910, n911, n913, n914, n915, n916, n917, n918, n919, n920, n922, n923,
    n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934;
  INVX1   g000(.A(COUNT_REG_0__SCAN_IN), .Y(U1391));
  INVX1   g001(.A(MEMORY_REG_31__1__SCAN_IN), .Y(n254));
  NAND2X1 g002(.A(WR_REG_SCAN_IN), .B(DATA_IN_REG_1__SCAN_IN), .Y(n255));
  INVX1   g003(.A(ADDRESS_REG_2__SCAN_IN), .Y(n256));
  INVX1   g004(.A(ADDRESS_REG_0__SCAN_IN), .Y(n257));
  NOR2X1  g005(.A(n257), .B(n256), .Y(n258));
  NAND4X1 g006(.A(ADDRESS_REG_1__SCAN_IN), .B(ADDRESS_REG_3__SCAN_IN), .C(ADDRESS_REG_4__SCAN_IN), .D(n258), .Y(n259));
  INVX1   g007(.A(WR_REG_SCAN_IN), .Y(n260));
  NOR2X1  g008(.A(n259), .B(n260), .Y(n261));
  OAI22X1 g009(.A0(n259), .A1(n255), .B0(n254), .B1(n261), .Y(U1486));
  INVX1   g010(.A(MEMORY_REG_31__0__SCAN_IN), .Y(n263));
  NAND2X1 g011(.A(WR_REG_SCAN_IN), .B(DATA_IN_REG_0__SCAN_IN), .Y(n264));
  OAI22X1 g012(.A0(n261), .A1(n263), .B0(n259), .B1(n264), .Y(U1485));
  INVX1   g013(.A(MEMORY_REG_30__1__SCAN_IN), .Y(n266));
  NOR2X1  g014(.A(ADDRESS_REG_0__SCAN_IN), .B(n256), .Y(n267));
  NAND4X1 g015(.A(ADDRESS_REG_1__SCAN_IN), .B(ADDRESS_REG_3__SCAN_IN), .C(ADDRESS_REG_4__SCAN_IN), .D(n267), .Y(n268));
  NOR2X1  g016(.A(n268), .B(n260), .Y(n269));
  OAI22X1 g017(.A0(n268), .A1(n255), .B0(n266), .B1(n269), .Y(U1484));
  INVX1   g018(.A(MEMORY_REG_30__0__SCAN_IN), .Y(n271));
  OAI22X1 g019(.A0(n268), .A1(n264), .B0(n271), .B1(n269), .Y(U1483));
  INVX1   g020(.A(MEMORY_REG_29__1__SCAN_IN), .Y(n273));
  INVX1   g021(.A(ADDRESS_REG_1__SCAN_IN), .Y(n274));
  NAND4X1 g022(.A(n274), .B(ADDRESS_REG_3__SCAN_IN), .C(ADDRESS_REG_4__SCAN_IN), .D(n258), .Y(n275));
  NOR2X1  g023(.A(n275), .B(n260), .Y(n276));
  OAI22X1 g024(.A0(n275), .A1(n255), .B0(n273), .B1(n276), .Y(U1482));
  INVX1   g025(.A(MEMORY_REG_29__0__SCAN_IN), .Y(n278));
  OAI22X1 g026(.A0(n275), .A1(n264), .B0(n278), .B1(n276), .Y(U1481));
  INVX1   g027(.A(MEMORY_REG_28__1__SCAN_IN), .Y(n280));
  NAND4X1 g028(.A(n274), .B(ADDRESS_REG_3__SCAN_IN), .C(ADDRESS_REG_4__SCAN_IN), .D(n267), .Y(n281));
  NOR2X1  g029(.A(n281), .B(n260), .Y(n282));
  OAI22X1 g030(.A0(n281), .A1(n255), .B0(n280), .B1(n282), .Y(U1480));
  INVX1   g031(.A(MEMORY_REG_28__0__SCAN_IN), .Y(n284));
  OAI22X1 g032(.A0(n281), .A1(n264), .B0(n284), .B1(n282), .Y(U1479));
  INVX1   g033(.A(MEMORY_REG_27__1__SCAN_IN), .Y(n286));
  NOR2X1  g034(.A(n257), .B(ADDRESS_REG_2__SCAN_IN), .Y(n287));
  NAND4X1 g035(.A(ADDRESS_REG_1__SCAN_IN), .B(ADDRESS_REG_3__SCAN_IN), .C(ADDRESS_REG_4__SCAN_IN), .D(n287), .Y(n288));
  NOR2X1  g036(.A(n288), .B(n260), .Y(n289));
  OAI22X1 g037(.A0(n288), .A1(n255), .B0(n286), .B1(n289), .Y(U1478));
  INVX1   g038(.A(MEMORY_REG_27__0__SCAN_IN), .Y(n291));
  OAI22X1 g039(.A0(n288), .A1(n264), .B0(n291), .B1(n289), .Y(U1477));
  INVX1   g040(.A(MEMORY_REG_26__1__SCAN_IN), .Y(n293));
  NOR2X1  g041(.A(ADDRESS_REG_0__SCAN_IN), .B(ADDRESS_REG_2__SCAN_IN), .Y(n294));
  NAND4X1 g042(.A(ADDRESS_REG_1__SCAN_IN), .B(ADDRESS_REG_3__SCAN_IN), .C(ADDRESS_REG_4__SCAN_IN), .D(n294), .Y(n295));
  NOR2X1  g043(.A(n295), .B(n260), .Y(n296));
  OAI22X1 g044(.A0(n295), .A1(n255), .B0(n293), .B1(n296), .Y(U1476));
  INVX1   g045(.A(MEMORY_REG_26__0__SCAN_IN), .Y(n298));
  OAI22X1 g046(.A0(n295), .A1(n264), .B0(n298), .B1(n296), .Y(U1475));
  INVX1   g047(.A(MEMORY_REG_25__1__SCAN_IN), .Y(n300));
  NAND4X1 g048(.A(n274), .B(ADDRESS_REG_3__SCAN_IN), .C(ADDRESS_REG_4__SCAN_IN), .D(n287), .Y(n301));
  NOR2X1  g049(.A(n301), .B(n260), .Y(n302));
  OAI22X1 g050(.A0(n301), .A1(n255), .B0(n300), .B1(n302), .Y(U1474));
  INVX1   g051(.A(MEMORY_REG_25__0__SCAN_IN), .Y(n304));
  OAI22X1 g052(.A0(n301), .A1(n264), .B0(n304), .B1(n302), .Y(U1473));
  INVX1   g053(.A(MEMORY_REG_24__1__SCAN_IN), .Y(n306));
  NAND4X1 g054(.A(n274), .B(ADDRESS_REG_3__SCAN_IN), .C(ADDRESS_REG_4__SCAN_IN), .D(n294), .Y(n307));
  NOR2X1  g055(.A(n307), .B(n260), .Y(n308));
  OAI22X1 g056(.A0(n307), .A1(n255), .B0(n306), .B1(n308), .Y(U1472));
  INVX1   g057(.A(MEMORY_REG_24__0__SCAN_IN), .Y(n310));
  OAI22X1 g058(.A0(n307), .A1(n264), .B0(n310), .B1(n308), .Y(U1471));
  INVX1   g059(.A(MEMORY_REG_23__1__SCAN_IN), .Y(n312));
  INVX1   g060(.A(ADDRESS_REG_3__SCAN_IN), .Y(n313));
  NAND4X1 g061(.A(ADDRESS_REG_1__SCAN_IN), .B(n313), .C(ADDRESS_REG_4__SCAN_IN), .D(n258), .Y(n314));
  NOR2X1  g062(.A(n314), .B(n260), .Y(n315));
  OAI22X1 g063(.A0(n314), .A1(n255), .B0(n312), .B1(n315), .Y(U1470));
  INVX1   g064(.A(MEMORY_REG_23__0__SCAN_IN), .Y(n317));
  OAI22X1 g065(.A0(n314), .A1(n264), .B0(n317), .B1(n315), .Y(U1469));
  INVX1   g066(.A(MEMORY_REG_22__1__SCAN_IN), .Y(n319));
  NAND4X1 g067(.A(ADDRESS_REG_1__SCAN_IN), .B(n313), .C(ADDRESS_REG_4__SCAN_IN), .D(n267), .Y(n320));
  NOR2X1  g068(.A(n320), .B(n260), .Y(n321));
  OAI22X1 g069(.A0(n320), .A1(n255), .B0(n319), .B1(n321), .Y(U1468));
  INVX1   g070(.A(MEMORY_REG_22__0__SCAN_IN), .Y(n323));
  OAI22X1 g071(.A0(n320), .A1(n264), .B0(n323), .B1(n321), .Y(U1467));
  INVX1   g072(.A(MEMORY_REG_21__1__SCAN_IN), .Y(n325));
  NAND4X1 g073(.A(n274), .B(n313), .C(ADDRESS_REG_4__SCAN_IN), .D(n258), .Y(n326));
  NOR2X1  g074(.A(n326), .B(n260), .Y(n327));
  OAI22X1 g075(.A0(n326), .A1(n255), .B0(n325), .B1(n327), .Y(U1466));
  INVX1   g076(.A(MEMORY_REG_21__0__SCAN_IN), .Y(n329));
  OAI22X1 g077(.A0(n326), .A1(n264), .B0(n329), .B1(n327), .Y(U1465));
  INVX1   g078(.A(MEMORY_REG_20__1__SCAN_IN), .Y(n331));
  NAND4X1 g079(.A(n274), .B(n313), .C(ADDRESS_REG_4__SCAN_IN), .D(n267), .Y(n332));
  NOR2X1  g080(.A(n332), .B(n260), .Y(n333));
  OAI22X1 g081(.A0(n332), .A1(n255), .B0(n331), .B1(n333), .Y(U1464));
  INVX1   g082(.A(MEMORY_REG_20__0__SCAN_IN), .Y(n335));
  OAI22X1 g083(.A0(n332), .A1(n264), .B0(n335), .B1(n333), .Y(U1463));
  INVX1   g084(.A(MEMORY_REG_19__1__SCAN_IN), .Y(n337));
  NAND4X1 g085(.A(ADDRESS_REG_1__SCAN_IN), .B(n313), .C(ADDRESS_REG_4__SCAN_IN), .D(n287), .Y(n338));
  NOR2X1  g086(.A(n338), .B(n260), .Y(n339));
  OAI22X1 g087(.A0(n338), .A1(n255), .B0(n337), .B1(n339), .Y(U1462));
  INVX1   g088(.A(MEMORY_REG_19__0__SCAN_IN), .Y(n341));
  OAI22X1 g089(.A0(n338), .A1(n264), .B0(n341), .B1(n339), .Y(U1461));
  INVX1   g090(.A(MEMORY_REG_18__1__SCAN_IN), .Y(n343));
  NAND4X1 g091(.A(ADDRESS_REG_1__SCAN_IN), .B(n313), .C(ADDRESS_REG_4__SCAN_IN), .D(n294), .Y(n344));
  NOR2X1  g092(.A(n344), .B(n260), .Y(n345));
  OAI22X1 g093(.A0(n344), .A1(n255), .B0(n343), .B1(n345), .Y(U1460));
  INVX1   g094(.A(MEMORY_REG_18__0__SCAN_IN), .Y(n347));
  OAI22X1 g095(.A0(n344), .A1(n264), .B0(n347), .B1(n345), .Y(U1459));
  INVX1   g096(.A(MEMORY_REG_17__1__SCAN_IN), .Y(n349));
  NAND4X1 g097(.A(n274), .B(n313), .C(ADDRESS_REG_4__SCAN_IN), .D(n287), .Y(n350));
  NOR2X1  g098(.A(n350), .B(n260), .Y(n351));
  OAI22X1 g099(.A0(n350), .A1(n255), .B0(n349), .B1(n351), .Y(U1458));
  INVX1   g100(.A(MEMORY_REG_17__0__SCAN_IN), .Y(n353));
  OAI22X1 g101(.A0(n350), .A1(n264), .B0(n353), .B1(n351), .Y(U1457));
  INVX1   g102(.A(MEMORY_REG_16__1__SCAN_IN), .Y(n355));
  NAND4X1 g103(.A(n274), .B(n313), .C(ADDRESS_REG_4__SCAN_IN), .D(n294), .Y(n356));
  NOR2X1  g104(.A(n356), .B(n260), .Y(n357));
  OAI22X1 g105(.A0(n356), .A1(n255), .B0(n355), .B1(n357), .Y(U1456));
  INVX1   g106(.A(MEMORY_REG_16__0__SCAN_IN), .Y(n359));
  OAI22X1 g107(.A0(n356), .A1(n264), .B0(n359), .B1(n357), .Y(U1455));
  INVX1   g108(.A(MEMORY_REG_15__1__SCAN_IN), .Y(n361));
  INVX1   g109(.A(ADDRESS_REG_4__SCAN_IN), .Y(n362));
  NAND4X1 g110(.A(ADDRESS_REG_1__SCAN_IN), .B(ADDRESS_REG_3__SCAN_IN), .C(n362), .D(n258), .Y(n363));
  NOR2X1  g111(.A(n363), .B(n260), .Y(n364));
  OAI22X1 g112(.A0(n363), .A1(n255), .B0(n361), .B1(n364), .Y(U1454));
  INVX1   g113(.A(MEMORY_REG_15__0__SCAN_IN), .Y(n366));
  OAI22X1 g114(.A0(n363), .A1(n264), .B0(n366), .B1(n364), .Y(U1453));
  INVX1   g115(.A(MEMORY_REG_14__1__SCAN_IN), .Y(n368));
  NAND4X1 g116(.A(ADDRESS_REG_1__SCAN_IN), .B(ADDRESS_REG_3__SCAN_IN), .C(n362), .D(n267), .Y(n369));
  NOR2X1  g117(.A(n369), .B(n260), .Y(n370));
  OAI22X1 g118(.A0(n369), .A1(n255), .B0(n368), .B1(n370), .Y(U1452));
  INVX1   g119(.A(MEMORY_REG_14__0__SCAN_IN), .Y(n372));
  OAI22X1 g120(.A0(n369), .A1(n264), .B0(n372), .B1(n370), .Y(U1451));
  INVX1   g121(.A(MEMORY_REG_13__1__SCAN_IN), .Y(n374));
  NAND4X1 g122(.A(n274), .B(ADDRESS_REG_3__SCAN_IN), .C(n362), .D(n258), .Y(n375));
  NOR2X1  g123(.A(n375), .B(n260), .Y(n376));
  OAI22X1 g124(.A0(n375), .A1(n255), .B0(n374), .B1(n376), .Y(U1450));
  INVX1   g125(.A(MEMORY_REG_13__0__SCAN_IN), .Y(n378));
  OAI22X1 g126(.A0(n375), .A1(n264), .B0(n378), .B1(n376), .Y(U1449));
  INVX1   g127(.A(MEMORY_REG_12__1__SCAN_IN), .Y(n380));
  NAND4X1 g128(.A(n274), .B(ADDRESS_REG_3__SCAN_IN), .C(n362), .D(n267), .Y(n381));
  NOR2X1  g129(.A(n381), .B(n260), .Y(n382));
  OAI22X1 g130(.A0(n381), .A1(n255), .B0(n380), .B1(n382), .Y(U1448));
  INVX1   g131(.A(MEMORY_REG_12__0__SCAN_IN), .Y(n384));
  OAI22X1 g132(.A0(n381), .A1(n264), .B0(n384), .B1(n382), .Y(U1447));
  INVX1   g133(.A(MEMORY_REG_11__1__SCAN_IN), .Y(n386));
  NAND4X1 g134(.A(ADDRESS_REG_1__SCAN_IN), .B(ADDRESS_REG_3__SCAN_IN), .C(n362), .D(n287), .Y(n387));
  NOR2X1  g135(.A(n387), .B(n260), .Y(n388));
  OAI22X1 g136(.A0(n387), .A1(n255), .B0(n386), .B1(n388), .Y(U1446));
  INVX1   g137(.A(MEMORY_REG_11__0__SCAN_IN), .Y(n390));
  OAI22X1 g138(.A0(n387), .A1(n264), .B0(n390), .B1(n388), .Y(U1445));
  INVX1   g139(.A(MEMORY_REG_10__1__SCAN_IN), .Y(n392));
  NAND4X1 g140(.A(ADDRESS_REG_1__SCAN_IN), .B(ADDRESS_REG_3__SCAN_IN), .C(n362), .D(n294), .Y(n393));
  NOR2X1  g141(.A(n393), .B(n260), .Y(n394));
  OAI22X1 g142(.A0(n393), .A1(n255), .B0(n392), .B1(n394), .Y(U1444));
  INVX1   g143(.A(MEMORY_REG_10__0__SCAN_IN), .Y(n396));
  OAI22X1 g144(.A0(n393), .A1(n264), .B0(n396), .B1(n394), .Y(U1443));
  INVX1   g145(.A(MEMORY_REG_9__1__SCAN_IN), .Y(n398));
  NAND4X1 g146(.A(n274), .B(ADDRESS_REG_3__SCAN_IN), .C(n362), .D(n287), .Y(n399));
  NOR2X1  g147(.A(n399), .B(n260), .Y(n400));
  OAI22X1 g148(.A0(n399), .A1(n255), .B0(n398), .B1(n400), .Y(U1442));
  INVX1   g149(.A(MEMORY_REG_9__0__SCAN_IN), .Y(n402));
  OAI22X1 g150(.A0(n399), .A1(n264), .B0(n402), .B1(n400), .Y(U1441));
  INVX1   g151(.A(MEMORY_REG_8__1__SCAN_IN), .Y(n404));
  NAND4X1 g152(.A(n274), .B(ADDRESS_REG_3__SCAN_IN), .C(n362), .D(n294), .Y(n405));
  NOR2X1  g153(.A(n405), .B(n260), .Y(n406));
  OAI22X1 g154(.A0(n405), .A1(n255), .B0(n404), .B1(n406), .Y(U1440));
  INVX1   g155(.A(MEMORY_REG_8__0__SCAN_IN), .Y(n408));
  OAI22X1 g156(.A0(n405), .A1(n264), .B0(n408), .B1(n406), .Y(U1439));
  INVX1   g157(.A(MEMORY_REG_7__1__SCAN_IN), .Y(n410));
  NAND4X1 g158(.A(ADDRESS_REG_1__SCAN_IN), .B(n313), .C(n362), .D(n258), .Y(n411));
  NOR2X1  g159(.A(n411), .B(n260), .Y(n412));
  OAI22X1 g160(.A0(n411), .A1(n255), .B0(n410), .B1(n412), .Y(U1438));
  INVX1   g161(.A(MEMORY_REG_7__0__SCAN_IN), .Y(n414));
  OAI22X1 g162(.A0(n411), .A1(n264), .B0(n414), .B1(n412), .Y(U1437));
  INVX1   g163(.A(MEMORY_REG_6__1__SCAN_IN), .Y(n416));
  NAND4X1 g164(.A(ADDRESS_REG_1__SCAN_IN), .B(n313), .C(n362), .D(n267), .Y(n417));
  NOR2X1  g165(.A(n417), .B(n260), .Y(n418));
  OAI22X1 g166(.A0(n417), .A1(n255), .B0(n416), .B1(n418), .Y(U1436));
  INVX1   g167(.A(MEMORY_REG_6__0__SCAN_IN), .Y(n420));
  OAI22X1 g168(.A0(n417), .A1(n264), .B0(n420), .B1(n418), .Y(U1435));
  INVX1   g169(.A(MEMORY_REG_5__1__SCAN_IN), .Y(n422));
  NAND4X1 g170(.A(n274), .B(n313), .C(n362), .D(n258), .Y(n423));
  NOR2X1  g171(.A(n423), .B(n260), .Y(n424));
  OAI22X1 g172(.A0(n423), .A1(n255), .B0(n422), .B1(n424), .Y(U1434));
  INVX1   g173(.A(MEMORY_REG_5__0__SCAN_IN), .Y(n426));
  OAI22X1 g174(.A0(n423), .A1(n264), .B0(n426), .B1(n424), .Y(U1433));
  INVX1   g175(.A(MEMORY_REG_4__1__SCAN_IN), .Y(n428));
  NAND4X1 g176(.A(n274), .B(n313), .C(n362), .D(n267), .Y(n429));
  NOR2X1  g177(.A(n429), .B(n260), .Y(n430));
  OAI22X1 g178(.A0(n429), .A1(n255), .B0(n428), .B1(n430), .Y(U1432));
  INVX1   g179(.A(MEMORY_REG_4__0__SCAN_IN), .Y(n432));
  OAI22X1 g180(.A0(n429), .A1(n264), .B0(n432), .B1(n430), .Y(U1431));
  INVX1   g181(.A(MEMORY_REG_3__1__SCAN_IN), .Y(n434));
  NAND4X1 g182(.A(ADDRESS_REG_1__SCAN_IN), .B(n313), .C(n362), .D(n287), .Y(n435));
  NOR2X1  g183(.A(n435), .B(n260), .Y(n436));
  OAI22X1 g184(.A0(n435), .A1(n255), .B0(n434), .B1(n436), .Y(U1430));
  INVX1   g185(.A(MEMORY_REG_3__0__SCAN_IN), .Y(n438));
  OAI22X1 g186(.A0(n435), .A1(n264), .B0(n438), .B1(n436), .Y(U1429));
  INVX1   g187(.A(MEMORY_REG_2__1__SCAN_IN), .Y(n440));
  NAND4X1 g188(.A(ADDRESS_REG_1__SCAN_IN), .B(n313), .C(n362), .D(n294), .Y(n441));
  NOR2X1  g189(.A(n441), .B(n260), .Y(n442));
  OAI22X1 g190(.A0(n441), .A1(n255), .B0(n440), .B1(n442), .Y(U1428));
  INVX1   g191(.A(MEMORY_REG_2__0__SCAN_IN), .Y(n444));
  OAI22X1 g192(.A0(n441), .A1(n264), .B0(n444), .B1(n442), .Y(U1427));
  INVX1   g193(.A(MEMORY_REG_1__1__SCAN_IN), .Y(n446));
  NAND4X1 g194(.A(n274), .B(n313), .C(n362), .D(n287), .Y(n447));
  NOR2X1  g195(.A(n447), .B(n260), .Y(n448));
  OAI22X1 g196(.A0(n447), .A1(n255), .B0(n446), .B1(n448), .Y(U1426));
  INVX1   g197(.A(MEMORY_REG_1__0__SCAN_IN), .Y(n450));
  OAI22X1 g198(.A0(n447), .A1(n264), .B0(n450), .B1(n448), .Y(U1425));
  INVX1   g199(.A(MEMORY_REG_0__1__SCAN_IN), .Y(n452));
  NAND4X1 g200(.A(n274), .B(n313), .C(n362), .D(n294), .Y(n453));
  NOR2X1  g201(.A(n453), .B(n260), .Y(n454));
  OAI22X1 g202(.A0(n453), .A1(n255), .B0(n452), .B1(n454), .Y(U1424));
  INVX1   g203(.A(MEMORY_REG_0__0__SCAN_IN), .Y(n456));
  OAI22X1 g204(.A0(n453), .A1(n264), .B0(n456), .B1(n454), .Y(U1423));
  INVX1   g205(.A(GAMMA_REG_0__SCAN_IN), .Y(n458));
  INVX1   g206(.A(START), .Y(n459));
  NAND2X1 g207(.A(n459), .B(n458), .Y(n460));
  NAND2X1 g208(.A(GAMMA_REG_3__SCAN_IN), .B(n459), .Y(n461));
  OAI21X1 g209(.A0(GAMMA_REG_1__SCAN_IN), .A1(n458), .B0(n459), .Y(n462));
  XOR2X1  g210(.A(MAX_REG_4__SCAN_IN), .B(SCAN_REG_4__SCAN_IN), .Y(n463));
  XOR2X1  g211(.A(MAX_REG_3__SCAN_IN), .B(SCAN_REG_3__SCAN_IN), .Y(n464));
  NOR2X1  g212(.A(n464), .B(n463), .Y(n465));
  XOR2X1  g213(.A(MAX_REG_2__SCAN_IN), .B(SCAN_REG_2__SCAN_IN), .Y(n466));
  XOR2X1  g214(.A(MAX_REG_1__SCAN_IN), .B(SCAN_REG_1__SCAN_IN), .Y(n467));
  XOR2X1  g215(.A(MAX_REG_0__SCAN_IN), .B(SCAN_REG_0__SCAN_IN), .Y(n468));
  NOR3X1  g216(.A(n468), .B(n467), .C(n466), .Y(n469));
  NAND4X1 g217(.A(n465), .B(n462), .C(n461), .D(n469), .Y(n470));
  INVX1   g218(.A(GAMMA_REG_3__SCAN_IN), .Y(n471));
  NOR2X1  g219(.A(n471), .B(START), .Y(n472));
  INVX1   g220(.A(GAMMA_REG_1__SCAN_IN), .Y(n473));
  AOI21X1 g221(.A0(n473), .A1(GAMMA_REG_0__SCAN_IN), .B0(START), .Y(n474));
  NOR3X1  g222(.A(n473), .B(START), .C(GAMMA_REG_0__SCAN_IN), .Y(n475));
  AOI21X1 g223(.A0(n474), .A1(n472), .B0(n475), .Y(n476));
  INVX1   g224(.A(COUNT_REG2_3__SCAN_IN), .Y(n477));
  INVX1   g225(.A(COUNT_REG2_1__SCAN_IN), .Y(n478));
  INVX1   g226(.A(GAMMA_REG_2__SCAN_IN), .Y(n479));
  NOR2X1  g227(.A(n479), .B(START), .Y(n480));
  NOR4X1  g228(.A(COUNT_REG2_2__SCAN_IN), .B(COUNT_REG2_4__SCAN_IN), .C(COUNT_REG2_5__SCAN_IN), .D(COUNT_REG2_0__SCAN_IN), .Y(n481));
  NAND4X1 g229(.A(n480), .B(n478), .C(n477), .D(n481), .Y(n482));
  AOI21X1 g230(.A0(n476), .A1(n470), .B0(n482), .Y(n483));
  NAND2X1 g231(.A(GAMMA_REG_4__SCAN_IN), .B(n459), .Y(n484));
  NAND3X1 g232(.A(n484), .B(n462), .C(n461), .Y(n485));
  AOI21X1 g233(.A0(n480), .A1(n474), .B0(n472), .Y(n486));
  INVX1   g234(.A(GAMMA_REG_4__SCAN_IN), .Y(n487));
  NOR2X1  g235(.A(n487), .B(START), .Y(n488));
  NAND4X1 g236(.A(n481), .B(n478), .C(n477), .D(n488), .Y(n489));
  OAI21X1 g237(.A0(n489), .A1(n486), .B0(n485), .Y(n490));
  NOR3X1  g238(.A(n473), .B(START), .C(n458), .Y(n491));
  OAI21X1 g239(.A0(GAMMA_REG_2__SCAN_IN), .A1(GAMMA_REG_4__SCAN_IN), .B0(n459), .Y(n492));
  NAND3X1 g240(.A(n492), .B(n491), .C(n472), .Y(n493));
  NOR2X1  g241(.A(START), .B(GAMMA_REG_0__SCAN_IN), .Y(n494));
  NOR2X1  g242(.A(n473), .B(START), .Y(n495));
  NOR3X1  g243(.A(n479), .B(n471), .C(START), .Y(n496));
  NAND4X1 g244(.A(n484), .B(n495), .C(n494), .D(n496), .Y(n497));
  OAI21X1 g245(.A0(GAMMA_REG_2__SCAN_IN), .A1(GAMMA_REG_3__SCAN_IN), .B0(n459), .Y(n498));
  NOR4X1  g246(.A(n487), .B(START), .C(n458), .D(n473), .Y(n499));
  NAND2X1 g247(.A(n499), .B(n498), .Y(n500));
  NAND3X1 g248(.A(n500), .B(n497), .C(n493), .Y(n501));
  NOR3X1  g249(.A(n501), .B(n490), .C(n483), .Y(n502));
  NAND3X1 g250(.A(GAMMA_REG_3__SCAN_IN), .B(GAMMA_REG_4__SCAN_IN), .C(n459), .Y(n503));
  NOR3X1  g251(.A(n503), .B(n502), .C(n460), .Y(n504));
  NOR2X1  g252(.A(n474), .B(n472), .Y(n505));
  OAI21X1 g253(.A0(n498), .A1(n505), .B0(n488), .Y(n506));
  OAI21X1 g254(.A0(GAMMA_REG_3__SCAN_IN), .A1(GAMMA_REG_4__SCAN_IN), .B0(n459), .Y(n507));
  NOR3X1  g255(.A(GAMMA_REG_1__SCAN_IN), .B(n479), .C(START), .Y(n508));
  AOI22X1 g256(.A0(n507), .A1(n508), .B0(n499), .B1(n480), .Y(n509));
  AOI21X1 g257(.A0(n509), .A1(n506), .B0(n502), .Y(n510));
  NAND2X1 g258(.A(DATA_OUT_REG_0__SCAN_IN), .B(DATA_OUT_REG_1__SCAN_IN), .Y(n511));
  INVX1   g259(.A(n511), .Y(n512));
  AOI21X1 g260(.A0(n512), .A1(n510), .B0(n504), .Y(n513));
  INVX1   g261(.A(IND_REG_1__SCAN_IN), .Y(n514));
  INVX1   g262(.A(IND_REG_0__SCAN_IN), .Y(n515));
  NAND3X1 g263(.A(GAMMA_REG_1__SCAN_IN), .B(n459), .C(n458), .Y(n516));
  AOI21X1 g264(.A0(n479), .A1(n487), .B0(START), .Y(n517));
  AOI21X1 g265(.A0(n517), .A1(n516), .B0(n461), .Y(n518));
  INVX1   g266(.A(n518), .Y(n519));
  NOR4X1  g267(.A(n502), .B(n515), .C(n514), .D(n519), .Y(n520));
  NAND2X1 g268(.A(GAMMA_REG_2__SCAN_IN), .B(n459), .Y(n521));
  OAI21X1 g269(.A0(n521), .A1(n462), .B0(n461), .Y(n522));
  NAND3X1 g270(.A(n481), .B(n478), .C(n477), .Y(n523));
  NOR2X1  g271(.A(n484), .B(n523), .Y(n524));
  AOI22X1 g272(.A0(n522), .A1(n524), .B0(n484), .B1(n505), .Y(n525));
  NAND4X1 g273(.A(n497), .B(n493), .C(n525), .D(n500), .Y(n526));
  OAI21X1 g274(.A0(n522), .A1(n484), .B0(n509), .Y(n528));
  NOR2X1  g275(.A(n518), .B(n528), .Y(n529));
  OAI21X1 g276(.A0(n526), .A1(n483), .B0(n529), .Y(n530));
  AOI21X1 g277(.A0(n530), .A1(NL_REG_3__SCAN_IN), .B0(n520), .Y(n531));
  NAND2X1 g278(.A(n531), .B(n513), .Y(U1422));
  NOR4X1  g279(.A(n502), .B(IND_REG_0__SCAN_IN), .C(n514), .D(n519), .Y(n533));
  NOR2X1  g280(.A(n533), .B(n504), .Y(n534));
  INVX1   g281(.A(DATA_OUT_REG_1__SCAN_IN), .Y(n535));
  NOR2X1  g282(.A(DATA_OUT_REG_0__SCAN_IN), .B(n535), .Y(n536));
  AOI22X1 g283(.A0(n530), .A1(NL_REG_2__SCAN_IN), .B0(n510), .B1(n536), .Y(n537));
  NAND2X1 g284(.A(n537), .B(n534), .Y(U1421));
  INVX1   g285(.A(DATA_OUT_REG_0__SCAN_IN), .Y(n539));
  NOR2X1  g286(.A(n539), .B(DATA_OUT_REG_1__SCAN_IN), .Y(n540));
  AOI21X1 g287(.A0(n540), .A1(n510), .B0(n504), .Y(n541));
  NOR4X1  g288(.A(n502), .B(n515), .C(IND_REG_1__SCAN_IN), .D(n519), .Y(n542));
  AOI21X1 g289(.A0(n530), .A1(NL_REG_1__SCAN_IN), .B0(n542), .Y(n543));
  NAND2X1 g290(.A(n543), .B(n541), .Y(U1420));
  NOR4X1  g291(.A(n502), .B(IND_REG_0__SCAN_IN), .C(IND_REG_1__SCAN_IN), .D(n519), .Y(n545));
  NOR2X1  g292(.A(n545), .B(n504), .Y(n546));
  NOR2X1  g293(.A(DATA_OUT_REG_0__SCAN_IN), .B(DATA_OUT_REG_1__SCAN_IN), .Y(n547));
  AOI22X1 g294(.A0(n530), .A1(NL_REG_0__SCAN_IN), .B0(n510), .B1(n547), .Y(n548));
  NAND2X1 g295(.A(n548), .B(n546), .Y(U1419));
  INVX1   g296(.A(SCAN_REG_4__SCAN_IN), .Y(n550));
  NAND2X1 g297(.A(n469), .B(n465), .Y(n551));
  INVX1   g298(.A(COUNT_REG2_2__SCAN_IN), .Y(n552));
  INVX1   g299(.A(COUNT_REG2_0__SCAN_IN), .Y(n553));
  NOR2X1  g300(.A(COUNT_REG2_4__SCAN_IN), .B(COUNT_REG2_5__SCAN_IN), .Y(n554));
  NAND3X1 g301(.A(n554), .B(n553), .C(n552), .Y(n555));
  NOR3X1  g302(.A(n555), .B(COUNT_REG2_1__SCAN_IN), .C(COUNT_REG2_3__SCAN_IN), .Y(n556));
  NAND3X1 g303(.A(GAMMA_REG_2__SCAN_IN), .B(GAMMA_REG_3__SCAN_IN), .C(n459), .Y(n557));
  NOR2X1  g304(.A(n557), .B(n474), .Y(n558));
  NAND3X1 g305(.A(n558), .B(n556), .C(n551), .Y(n559));
  NAND4X1 g306(.A(n521), .B(n495), .C(n494), .D(n507), .Y(n560));
  NAND2X1 g307(.A(GAMMA_REG_1__SCAN_IN), .B(n459), .Y(n561));
  AOI21X1 g308(.A0(n471), .A1(n487), .B0(START), .Y(n562));
  NOR4X1  g309(.A(n521), .B(n561), .C(n494), .D(n562), .Y(n563));
  NAND2X1 g310(.A(n563), .B(n556), .Y(n564));
  NAND3X1 g311(.A(n564), .B(n560), .C(n559), .Y(n565));
  NAND4X1 g312(.A(SCAN_REG_1__SCAN_IN), .B(SCAN_REG_2__SCAN_IN), .C(SCAN_REG_3__SCAN_IN), .D(SCAN_REG_0__SCAN_IN), .Y(n566));
  XOR2X1  g313(.A(n566), .B(SCAN_REG_4__SCAN_IN), .Y(n567));
  NAND3X1 g314(.A(n565), .B(n480), .C(n551), .Y(n568));
  OAI22X1 g315(.A0(n567), .A1(n568), .B0(n565), .B1(n550), .Y(U1418));
  INVX1   g316(.A(SCAN_REG_3__SCAN_IN), .Y(n570));
  NAND3X1 g317(.A(SCAN_REG_0__SCAN_IN), .B(SCAN_REG_1__SCAN_IN), .C(SCAN_REG_2__SCAN_IN), .Y(n571));
  XOR2X1  g318(.A(n571), .B(SCAN_REG_3__SCAN_IN), .Y(n572));
  OAI22X1 g319(.A0(n568), .A1(n572), .B0(n565), .B1(n570), .Y(U1417));
  INVX1   g320(.A(SCAN_REG_2__SCAN_IN), .Y(n574));
  NAND2X1 g321(.A(SCAN_REG_0__SCAN_IN), .B(SCAN_REG_1__SCAN_IN), .Y(n575));
  XOR2X1  g322(.A(n575), .B(SCAN_REG_2__SCAN_IN), .Y(n576));
  OAI22X1 g323(.A0(n568), .A1(n576), .B0(n565), .B1(n574), .Y(U1416));
  INVX1   g324(.A(SCAN_REG_1__SCAN_IN), .Y(n578));
  XOR2X1  g325(.A(SCAN_REG_0__SCAN_IN), .B(n578), .Y(n579));
  OAI22X1 g326(.A0(n568), .A1(n579), .B0(n565), .B1(n578), .Y(U1415));
  NAND4X1 g327(.A(n560), .B(n559), .C(SCAN_REG_0__SCAN_IN), .D(n564), .Y(n581));
  OAI21X1 g328(.A0(n568), .A1(SCAN_REG_0__SCAN_IN), .B0(n581), .Y(U1414));
  INVX1   g329(.A(MAX_REG_4__SCAN_IN), .Y(n583));
  NAND3X1 g330(.A(n556), .B(n469), .C(n465), .Y(n584));
  INVX1   g331(.A(MAX_REG_2__SCAN_IN), .Y(n585));
  INVX1   g332(.A(MAX_REG_1__SCAN_IN), .Y(n586));
  NOR3X1  g333(.A(n586), .B(n585), .C(n583), .Y(n587));
  NAND3X1 g334(.A(n587), .B(MAX_REG_0__SCAN_IN), .C(MAX_REG_3__SCAN_IN), .Y(n588));
  NAND2X1 g335(.A(n588), .B(n558), .Y(n589));
  NOR2X1  g336(.A(n589), .B(n584), .Y(n590));
  AOI21X1 g337(.A0(n492), .A1(n505), .B0(n590), .Y(n591));
  NOR3X1  g338(.A(n480), .B(n516), .C(n461), .Y(n592));
  NAND4X1 g339(.A(GAMMA_REG_4__SCAN_IN), .B(n459), .C(GAMMA_REG_0__SCAN_IN), .D(n473), .Y(n593));
  NOR2X1  g340(.A(n593), .B(n521), .Y(n594));
  AOI21X1 g341(.A0(n594), .A1(n551), .B0(n592), .Y(n595));
  NOR3X1  g342(.A(GAMMA_REG_1__SCAN_IN), .B(START), .C(GAMMA_REG_0__SCAN_IN), .Y(n596));
  NAND3X1 g343(.A(n596), .B(n498), .C(n488), .Y(n597));
  NAND2X1 g344(.A(n597), .B(n595), .Y(n598));
  NAND2X1 g345(.A(n598), .B(n556), .Y(n599));
  NAND2X1 g346(.A(n599), .B(n591), .Y(n600));
  NAND4X1 g347(.A(MAX_REG_1__SCAN_IN), .B(MAX_REG_2__SCAN_IN), .C(MAX_REG_3__SCAN_IN), .D(MAX_REG_0__SCAN_IN), .Y(n601));
  XOR2X1  g348(.A(n601), .B(MAX_REG_4__SCAN_IN), .Y(n602));
  NAND3X1 g349(.A(n492), .B(n462), .C(n461), .Y(n603));
  OAI21X1 g350(.A0(n589), .A1(n584), .B0(n603), .Y(n604));
  AOI21X1 g351(.A0(n597), .A1(n595), .B0(n523), .Y(n605));
  OAI21X1 g352(.A0(n605), .A1(n604), .B0(n480), .Y(n606));
  OAI22X1 g353(.A0(n602), .A1(n606), .B0(n600), .B1(n583), .Y(U1413));
  NOR2X1  g354(.A(n605), .B(n604), .Y(n608));
  NAND2X1 g355(.A(n608), .B(MAX_REG_3__SCAN_IN), .Y(n609));
  NAND3X1 g356(.A(MAX_REG_0__SCAN_IN), .B(MAX_REG_1__SCAN_IN), .C(MAX_REG_2__SCAN_IN), .Y(n610));
  XOR2X1  g357(.A(n610), .B(MAX_REG_3__SCAN_IN), .Y(n611));
  OAI21X1 g358(.A0(n611), .A1(n606), .B0(n609), .Y(U1412));
  NAND2X1 g359(.A(MAX_REG_0__SCAN_IN), .B(MAX_REG_1__SCAN_IN), .Y(n613));
  XOR2X1  g360(.A(n613), .B(MAX_REG_2__SCAN_IN), .Y(n614));
  OAI22X1 g361(.A0(n606), .A1(n614), .B0(n600), .B1(n585), .Y(U1411));
  XOR2X1  g362(.A(MAX_REG_0__SCAN_IN), .B(n586), .Y(n616));
  OAI22X1 g363(.A0(n606), .A1(n616), .B0(n600), .B1(n586), .Y(U1410));
  NAND2X1 g364(.A(n608), .B(MAX_REG_0__SCAN_IN), .Y(n618));
  OAI21X1 g365(.A0(n606), .A1(MAX_REG_0__SCAN_IN), .B0(n618), .Y(U1409));
  NOR4X1  g366(.A(K_1_), .B(K_2_), .C(K_3_), .D(K_0_), .Y(n620));
  INVX1   g367(.A(n620), .Y(n621));
  NAND3X1 g368(.A(n621), .B(n592), .C(n523), .Y(n622));
  INVX1   g369(.A(n622), .Y(n623));
  NOR2X1  g370(.A(K_0_), .B(K_1_), .Y(n624));
  NAND4X1 g371(.A(n624), .B(n592), .C(n523), .D(n621), .Y(n625));
  OAI21X1 g372(.A0(n623), .A1(n514), .B0(n625), .Y(U1564));
  INVX1   g373(.A(K_1_), .Y(n627));
  AOI21X1 g374(.A0(n627), .A1(K_2_), .B0(K_0_), .Y(n628));
  NAND4X1 g375(.A(n621), .B(n592), .C(n523), .D(n628), .Y(n629));
  OAI21X1 g376(.A0(n623), .A1(n515), .B0(n629), .Y(U1565));
  INVX1   g377(.A(TIMEBASE_REG_5__SCAN_IN), .Y(n631));
  NAND4X1 g378(.A(n478), .B(n477), .C(TIMEBASE_REG_0__SCAN_IN), .D(n481), .Y(n632));
  NAND4X1 g379(.A(n478), .B(n477), .C(TIMEBASE_REG_1__SCAN_IN), .D(n481), .Y(n633));
  NAND4X1 g380(.A(n632), .B(n553), .C(n478), .D(n633), .Y(n634));
  INVX1   g381(.A(TIMEBASE_REG_2__SCAN_IN), .Y(n635));
  OAI21X1 g382(.A0(n523), .A1(n635), .B0(n552), .Y(n636));
  INVX1   g383(.A(TIMEBASE_REG_3__SCAN_IN), .Y(n637));
  OAI21X1 g384(.A0(n523), .A1(n637), .B0(n477), .Y(n638));
  INVX1   g385(.A(TIMEBASE_REG_4__SCAN_IN), .Y(n639));
  INVX1   g386(.A(COUNT_REG2_4__SCAN_IN), .Y(n640));
  OAI21X1 g387(.A0(n523), .A1(n639), .B0(n640), .Y(n641));
  NOR4X1  g388(.A(n638), .B(n636), .C(n634), .D(n641), .Y(n642));
  AOI21X1 g389(.A0(n556), .A1(TIMEBASE_REG_5__SCAN_IN), .B0(COUNT_REG2_5__SCAN_IN), .Y(n643));
  XOR2X1  g390(.A(n643), .B(n642), .Y(n644));
  NAND2X1 g391(.A(n644), .B(n472), .Y(n645));
  NAND2X1 g392(.A(n645), .B(n604), .Y(n646));
  OAI21X1 g393(.A0(n604), .A1(n631), .B0(n646), .Y(U1566));
  NOR3X1  g394(.A(n638), .B(n636), .C(n634), .Y(n648));
  XOR2X1  g395(.A(n641), .B(n648), .Y(n649));
  NAND3X1 g396(.A(n649), .B(n604), .C(n472), .Y(n650));
  OAI21X1 g397(.A0(n604), .A1(n639), .B0(n650), .Y(U1408));
  NAND2X1 g398(.A(n604), .B(n472), .Y(n652));
  NOR2X1  g399(.A(n636), .B(n634), .Y(n653));
  AOI21X1 g400(.A0(n556), .A1(TIMEBASE_REG_3__SCAN_IN), .B0(COUNT_REG2_3__SCAN_IN), .Y(n654));
  XOR2X1  g401(.A(n654), .B(n653), .Y(n655));
  OAI22X1 g402(.A0(n652), .A1(n655), .B0(n604), .B1(n637), .Y(U1407));
  INVX1   g403(.A(n634), .Y(n657));
  XOR2X1  g404(.A(n636), .B(n657), .Y(n658));
  NAND3X1 g405(.A(n658), .B(n604), .C(n472), .Y(n659));
  OAI21X1 g406(.A0(n604), .A1(n635), .B0(n659), .Y(U1406));
  INVX1   g407(.A(TIMEBASE_REG_1__SCAN_IN), .Y(n661));
  NAND2X1 g408(.A(n632), .B(n553), .Y(n662));
  INVX1   g409(.A(n662), .Y(n663));
  NAND2X1 g410(.A(n633), .B(n478), .Y(n664));
  XOR2X1  g411(.A(n664), .B(n663), .Y(n665));
  NAND3X1 g412(.A(n665), .B(n604), .C(n472), .Y(n666));
  OAI21X1 g413(.A0(n604), .A1(n661), .B0(n666), .Y(U1405));
  INVX1   g414(.A(TIMEBASE_REG_0__SCAN_IN), .Y(n668));
  OAI21X1 g415(.A0(n663), .A1(n461), .B0(n604), .Y(n669));
  OAI21X1 g416(.A0(n604), .A1(n668), .B0(n669), .Y(U1567));
  NOR4X1  g417(.A(n523), .B(n521), .C(n551), .D(n593), .Y(n671));
  OAI22X1 g418(.A0(n557), .A1(n474), .B0(n521), .B1(n593), .Y(n672));
  AOI21X1 g419(.A0(n672), .A1(n523), .B0(n671), .Y(n673));
  NAND3X1 g420(.A(n491), .B(n484), .C(n523), .Y(n674));
  NAND3X1 g421(.A(n488), .B(n474), .C(n461), .Y(n675));
  NAND3X1 g422(.A(n507), .B(n495), .C(n494), .Y(n676));
  NAND4X1 g423(.A(n676), .B(n675), .C(n674), .D(n485), .Y(n678));
  NAND2X1 g424(.A(n678), .B(n480), .Y(n679));
  NAND2X1 g425(.A(n496), .B(n462), .Y(n680));
  NOR4X1  g426(.A(n680), .B(n523), .C(n551), .D(n588), .Y(n681));
  NAND3X1 g427(.A(n523), .B(n521), .C(n494), .Y(n682));
  NOR3X1  g428(.A(GAMMA_REG_2__SCAN_IN), .B(n487), .C(START), .Y(n683));
  AOI22X1 g429(.A0(n596), .A1(n484), .B0(n561), .B1(n683), .Y(n684));
  AOI21X1 g430(.A0(n684), .A1(n682), .B0(n461), .Y(n685));
  NAND3X1 g431(.A(n496), .B(n495), .C(n460), .Y(n686));
  AOI22X1 g432(.A0(n596), .A1(n683), .B0(n499), .B1(n498), .Y(n687));
  OAI21X1 g433(.A0(n686), .A1(n488), .B0(n687), .Y(n688));
  NOR3X1  g434(.A(n688), .B(n685), .C(n681), .Y(n689));
  NAND3X1 g435(.A(n689), .B(n679), .C(n673), .Y(n690));
  NAND4X1 g436(.A(n487), .B(n459), .C(n458), .D(n471), .Y(n691));
  NAND4X1 g437(.A(GAMMA_REG_2__SCAN_IN), .B(GAMMA_REG_3__SCAN_IN), .C(n459), .D(GAMMA_REG_1__SCAN_IN), .Y(n692));
  AOI21X1 g438(.A0(n692), .A1(n691), .B0(n523), .Y(n693));
  INVX1   g439(.A(n596), .Y(n694));
  NOR3X1  g440(.A(n694), .B(n523), .C(n521), .Y(n695));
  NOR4X1  g441(.A(GAMMA_REG_2__SCAN_IN), .B(GAMMA_REG_3__SCAN_IN), .C(START), .D(n473), .Y(n696));
  OAI22X1 g442(.A0(n562), .A1(n495), .B0(n517), .B1(n620), .Y(n697));
  NOR4X1  g443(.A(n696), .B(n695), .C(n693), .D(n697), .Y(n698));
  NAND4X1 g444(.A(GAMMA_REG_3__SCAN_IN), .B(n459), .C(GAMMA_REG_0__SCAN_IN), .D(n473), .Y(n699));
  NAND3X1 g445(.A(n471), .B(n459), .C(n458), .Y(n700));
  NAND4X1 g446(.A(n699), .B(n593), .C(n503), .D(n700), .Y(n701));
  AOI21X1 g447(.A0(n480), .A1(n495), .B0(n596), .Y(n702));
  OAI22X1 g448(.A0(n621), .A1(n517), .B0(n556), .B1(n702), .Y(n703));
  AOI21X1 g449(.A0(n701), .A1(n523), .B0(n703), .Y(n704));
  OAI22X1 g450(.A0(n698), .A1(n631), .B0(n644), .B1(n704), .Y(n705));
  NAND2X1 g451(.A(n705), .B(n690), .Y(n706));
  NAND3X1 g452(.A(n690), .B(n492), .C(n561), .Y(n707));
  NAND4X1 g453(.A(n679), .B(n673), .C(COUNT_REG2_5__SCAN_IN), .D(n689), .Y(n708));
  NAND3X1 g454(.A(n708), .B(n707), .C(n706), .Y(U1404));
  NAND2X1 g455(.A(n701), .B(n523), .Y(n710));
  NOR2X1  g456(.A(n521), .B(n462), .Y(n711));
  NOR3X1  g457(.A(n621), .B(n517), .C(n561), .Y(n712));
  AOI21X1 g458(.A0(n711), .A1(n523), .B0(n712), .Y(n713));
  NAND2X1 g459(.A(n713), .B(n710), .Y(n714));
  NAND3X1 g460(.A(n714), .B(n690), .C(n649), .Y(n715));
  NAND4X1 g461(.A(n679), .B(n673), .C(COUNT_REG2_4__SCAN_IN), .D(n689), .Y(n716));
  INVX1   g462(.A(n695), .Y(n717));
  AOI21X1 g463(.A0(n479), .A1(n471), .B0(START), .Y(n718));
  NAND3X1 g464(.A(n473), .B(GAMMA_REG_2__SCAN_IN), .C(n459), .Y(n719));
  OAI22X1 g465(.A0(n562), .A1(n719), .B0(n718), .B1(n561), .Y(n720));
  NOR3X1  g466(.A(n620), .B(n517), .C(n561), .Y(n721));
  NOR3X1  g467(.A(n721), .B(n720), .C(n693), .Y(n722));
  NAND2X1 g468(.A(n722), .B(n717), .Y(n723));
  NAND3X1 g469(.A(n723), .B(n690), .C(TIMEBASE_REG_4__SCAN_IN), .Y(n724));
  NAND3X1 g470(.A(n724), .B(n716), .C(n715), .Y(U1403));
  AOI21X1 g471(.A0(n713), .A1(n710), .B0(n655), .Y(n726));
  NAND3X1 g472(.A(n699), .B(n593), .C(n503), .Y(n727));
  NAND3X1 g473(.A(GAMMA_REG_2__SCAN_IN), .B(GAMMA_REG_4__SCAN_IN), .C(n459), .Y(n728));
  OAI22X1 g474(.A0(n521), .A1(n637), .B0(n561), .B1(n728), .Y(n729));
  OAI21X1 g475(.A0(n729), .A1(n727), .B0(n556), .Y(n730));
  OAI21X1 g476(.A0(n722), .A1(n637), .B0(n730), .Y(n731));
  OAI21X1 g477(.A0(n731), .A1(n726), .B0(n690), .Y(n732));
  OAI21X1 g478(.A0(n690), .A1(n477), .B0(n732), .Y(U1568));
  NAND3X1 g479(.A(n714), .B(n690), .C(n658), .Y(n734));
  NAND4X1 g480(.A(n679), .B(n673), .C(COUNT_REG2_2__SCAN_IN), .D(n689), .Y(n735));
  NAND3X1 g481(.A(n723), .B(n690), .C(TIMEBASE_REG_2__SCAN_IN), .Y(n736));
  NAND3X1 g482(.A(n736), .B(n735), .C(n734), .Y(U1402));
  NAND3X1 g483(.A(n714), .B(n690), .C(n665), .Y(n738));
  NAND4X1 g484(.A(n679), .B(n673), .C(COUNT_REG2_1__SCAN_IN), .D(n689), .Y(n739));
  NAND3X1 g485(.A(n723), .B(n690), .C(TIMEBASE_REG_1__SCAN_IN), .Y(n740));
  NAND3X1 g486(.A(n740), .B(n739), .C(n738), .Y(U1401));
  OAI22X1 g487(.A0(n698), .A1(n668), .B0(n662), .B1(n704), .Y(n742));
  NAND2X1 g488(.A(n742), .B(n690), .Y(n743));
  NAND4X1 g489(.A(n679), .B(n673), .C(COUNT_REG2_0__SCAN_IN), .D(n689), .Y(n744));
  NAND3X1 g490(.A(n744), .B(n743), .C(n707), .Y(U1400));
  AOI21X1 g491(.A0(n718), .A1(n488), .B0(n496), .Y(n746));
  NOR4X1  g492(.A(n584), .B(n521), .C(n474), .D(n588), .Y(n747));
  NAND2X1 g493(.A(n622), .B(n500), .Y(n748));
  NOR4X1  g494(.A(n487), .B(START), .C(n458), .D(n471), .Y(n749));
  NOR2X1  g495(.A(n749), .B(n499), .Y(n750));
  OAI22X1 g496(.A0(n485), .A1(n521), .B0(n523), .B1(n750), .Y(n751));
  NOR4X1  g497(.A(n748), .B(n747), .C(n671), .D(n751), .Y(n752));
  NAND2X1 g498(.A(n752), .B(SOUND_REG_2__SCAN_IN), .Y(n753));
  OAI21X1 g499(.A0(n752), .A1(n746), .B0(n753), .Y(U1569));
  AOI22X1 g500(.A0(n624), .A1(n492), .B0(DATA_OUT_REG_1__SCAN_IN), .B1(n720), .Y(n755));
  NAND2X1 g501(.A(n752), .B(SOUND_REG_1__SCAN_IN), .Y(n756));
  OAI21X1 g502(.A0(n755), .A1(n752), .B0(n756), .Y(U1570));
  OAI21X1 g503(.A0(n472), .A1(n539), .B0(n728), .Y(n758));
  AOI21X1 g504(.A0(n628), .A1(n492), .B0(n758), .Y(n759));
  NAND2X1 g505(.A(n752), .B(SOUND_REG_0__SCAN_IN), .Y(n760));
  OAI21X1 g506(.A0(n759), .A1(n752), .B0(n760), .Y(U1571));
  NOR3X1  g507(.A(n694), .B(n517), .C(n461), .Y(n762));
  NAND3X1 g508(.A(GAMMA_REG_1__SCAN_IN), .B(n487), .C(n459), .Y(n763));
  AOI21X1 g509(.A0(n593), .A1(n763), .B0(n718), .Y(n764));
  OAI22X1 g510(.A0(n762), .A1(n764), .B0(n491), .B1(n472), .Y(n765));
  NOR2X1  g511(.A(n764), .B(n762), .Y(n766));
  AOI21X1 g512(.A0(n593), .A1(n516), .B0(n766), .Y(n767));
  AOI22X1 g513(.A0(n766), .A1(ADDRESS_REG_4__SCAN_IN), .B0(MAX_REG_4__SCAN_IN), .B1(n767), .Y(n768));
  OAI21X1 g514(.A0(n765), .A1(n550), .B0(n768), .Y(U1399));
  AOI22X1 g515(.A0(n766), .A1(ADDRESS_REG_3__SCAN_IN), .B0(MAX_REG_3__SCAN_IN), .B1(n767), .Y(n770));
  OAI21X1 g516(.A0(n765), .A1(n570), .B0(n770), .Y(U1398));
  AOI22X1 g517(.A0(n766), .A1(ADDRESS_REG_2__SCAN_IN), .B0(MAX_REG_2__SCAN_IN), .B1(n767), .Y(n772));
  OAI21X1 g518(.A0(n765), .A1(n574), .B0(n772), .Y(U1397));
  AOI22X1 g519(.A0(n766), .A1(ADDRESS_REG_1__SCAN_IN), .B0(MAX_REG_1__SCAN_IN), .B1(n767), .Y(n774));
  OAI21X1 g520(.A0(n765), .A1(n578), .B0(n774), .Y(U1396));
  INVX1   g521(.A(SCAN_REG_0__SCAN_IN), .Y(n776));
  AOI22X1 g522(.A0(n766), .A1(ADDRESS_REG_0__SCAN_IN), .B0(MAX_REG_0__SCAN_IN), .B1(n767), .Y(n777));
  OAI21X1 g523(.A0(n765), .A1(n776), .B0(n777), .Y(U1395));
  INVX1   g524(.A(NUM_REG_1__SCAN_IN), .Y(n779));
  NAND2X1 g525(.A(n560), .B(DATA_IN_REG_1__SCAN_IN), .Y(n780));
  OAI21X1 g526(.A0(n560), .A1(n779), .B0(n780), .Y(U1572));
  INVX1   g527(.A(NUM_REG_0__SCAN_IN), .Y(n782));
  NAND2X1 g528(.A(n560), .B(DATA_IN_REG_0__SCAN_IN), .Y(n783));
  OAI21X1 g529(.A0(n560), .A1(n782), .B0(n783), .Y(U1573));
  INVX1   g530(.A(COUNTER_REG_2__SCAN_IN), .Y(n785));
  INVX1   g531(.A(SOUND_REG_2__SCAN_IN), .Y(n786));
  INVX1   g532(.A(SOUND_REG_0__SCAN_IN), .Y(n787));
  NOR2X1  g533(.A(n787), .B(n786), .Y(n788));
  INVX1   g534(.A(SOUND_REG_1__SCAN_IN), .Y(n789));
  INVX1   g535(.A(COUNTER_REG_0__SCAN_IN), .Y(n790));
  OAI21X1 g536(.A0(n790), .A1(SOUND_REG_0__SCAN_IN), .B0(n789), .Y(n791));
  OAI21X1 g537(.A0(n791), .A1(n788), .B0(COUNTER_REG_1__SCAN_IN), .Y(n792));
  NAND3X1 g538(.A(COUNTER_REG_0__SCAN_IN), .B(n787), .C(SOUND_REG_1__SCAN_IN), .Y(n793));
  OAI21X1 g539(.A0(SOUND_REG_0__SCAN_IN), .A1(n786), .B0(n789), .Y(n794));
  AOI22X1 g540(.A0(n793), .A1(n792), .B0(n785), .B1(n794), .Y(n795));
  NOR2X1  g541(.A(n794), .B(n785), .Y(n796));
  NOR2X1  g542(.A(n796), .B(n795), .Y(n797));
  AOI21X1 g543(.A0(SOUND_REG_1__SCAN_IN), .A1(SOUND_REG_2__SCAN_IN), .B0(n797), .Y(n798));
  INVX1   g544(.A(PLAY_REG_SCAN_IN), .Y(n799));
  NOR2X1  g545(.A(n799), .B(S_REG_SCAN_IN), .Y(n800));
  NAND2X1 g546(.A(n800), .B(n798), .Y(n801));
  NAND2X1 g547(.A(SOUND_REG_1__SCAN_IN), .B(SOUND_REG_2__SCAN_IN), .Y(n802));
  OAI21X1 g548(.A0(n796), .A1(n795), .B0(n802), .Y(n803));
  OAI21X1 g549(.A0(n803), .A1(n799), .B0(S_REG_SCAN_IN), .Y(n804));
  NAND2X1 g550(.A(n804), .B(n801), .Y(U1394));
  NAND4X1 g551(.A(GAMMA_REG_4__SCAN_IN), .B(n459), .C(GAMMA_REG_0__SCAN_IN), .D(GAMMA_REG_1__SCAN_IN), .Y(n806));
  OAI21X1 g552(.A0(n728), .A1(n494), .B0(n806), .Y(n807));
  NAND3X1 g553(.A(n521), .B(n475), .C(n472), .Y(n808));
  AOI21X1 g554(.A0(n488), .A1(n472), .B0(n480), .Y(n809));
  NAND2X1 g555(.A(n728), .B(n462), .Y(n810));
  OAI22X1 g556(.A0(n809), .A1(n810), .B0(n808), .B1(n488), .Y(n811));
  AOI21X1 g557(.A0(n807), .A1(n461), .B0(n811), .Y(n812));
  NOR2X1  g558(.A(n692), .B(n494), .Y(n813));
  NAND4X1 g559(.A(GAMMA_REG_3__SCAN_IN), .B(n459), .C(n458), .D(GAMMA_REG_2__SCAN_IN), .Y(n814));
  NAND3X1 g560(.A(GAMMA_REG_2__SCAN_IN), .B(n471), .C(n459), .Y(n815));
  OAI22X1 g561(.A0(n814), .A1(n495), .B0(n516), .B1(n815), .Y(n816));
  OAI21X1 g562(.A0(n816), .A1(n813), .B0(n556), .Y(n817));
  NAND2X1 g563(.A(n817), .B(n525), .Y(n818));
  NOR4X1  g564(.A(n748), .B(n747), .C(n671), .D(n818), .Y(n819));
  NAND2X1 g565(.A(n819), .B(PLAY_REG_SCAN_IN), .Y(n820));
  OAI21X1 g566(.A0(n819), .A1(n812), .B0(n820), .Y(U1574));
  AOI21X1 g567(.A0(n511), .A1(K_3_), .B0(K_2_), .Y(n822));
  INVX1   g568(.A(K_2_), .Y(n823));
  NOR3X1  g569(.A(DATA_OUT_REG_0__SCAN_IN), .B(n535), .C(n823), .Y(n824));
  NOR4X1  g570(.A(n822), .B(K_0_), .C(K_1_), .D(n824), .Y(n825));
  INVX1   g571(.A(K_0_), .Y(n826));
  NAND2X1 g572(.A(n826), .B(K_1_), .Y(n827));
  OAI22X1 g573(.A0(n547), .A1(n826), .B0(n540), .B1(n827), .Y(n828));
  NOR2X1  g574(.A(n808), .B(n556), .Y(n829));
  OAI21X1 g575(.A0(n828), .A1(n825), .B0(n829), .Y(n830));
  AOI22X1 g576(.A0(n492), .A1(n505), .B0(n556), .B1(n592), .Y(n831));
  NAND2X1 g577(.A(n831), .B(n830), .Y(n832));
  NAND2X1 g578(.A(n832), .B(n472), .Y(n833));
  NAND3X1 g579(.A(n831), .B(n830), .C(NLOSS_REG_SCAN_IN), .Y(n834));
  NAND2X1 g580(.A(n834), .B(n833), .Y(U1575));
  NAND3X1 g581(.A(n803), .B(SPEAKER_REG_SCAN_IN), .C(PLAY_REG_SCAN_IN), .Y(n836));
  NAND2X1 g582(.A(n836), .B(n801), .Y(U1393));
  NOR3X1  g583(.A(n562), .B(n480), .C(n494), .Y(n838));
  OAI21X1 g584(.A0(n838), .A1(n260), .B0(n560), .Y(U1392));
  NAND3X1 g585(.A(n802), .B(n797), .C(PLAY_REG_SCAN_IN), .Y(n840));
  AOI21X1 g586(.A0(COUNTER_REG_0__SCAN_IN), .A1(COUNTER_REG_1__SCAN_IN), .B0(COUNTER_REG_2__SCAN_IN), .Y(n841));
  NOR2X1  g587(.A(n841), .B(n840), .Y(U1381));
  XOR2X1  g588(.A(n790), .B(COUNTER_REG_1__SCAN_IN), .Y(n843));
  NOR2X1  g589(.A(n843), .B(n840), .Y(U1382));
  NOR2X1  g590(.A(n840), .B(COUNTER_REG_0__SCAN_IN), .Y(U1383));
  XOR2X1  g591(.A(COUNT_REG_1__SCAN_IN), .B(COUNT_REG_0__SCAN_IN), .Y(U1563));
  OAI22X1 g592(.A0(n387), .A1(n386), .B0(n392), .B1(n393), .Y(n847));
  OAI22X1 g593(.A0(n399), .A1(n398), .B0(n404), .B1(n405), .Y(n848));
  OAI22X1 g594(.A0(n363), .A1(n361), .B0(n368), .B1(n369), .Y(n849));
  OAI22X1 g595(.A0(n375), .A1(n374), .B0(n380), .B1(n381), .Y(n850));
  NOR4X1  g596(.A(n849), .B(n848), .C(n847), .D(n850), .Y(n851));
  OAI22X1 g597(.A0(n435), .A1(n434), .B0(n440), .B1(n441), .Y(n852));
  OAI22X1 g598(.A0(n447), .A1(n446), .B0(n452), .B1(n453), .Y(n853));
  OAI22X1 g599(.A0(n411), .A1(n410), .B0(n416), .B1(n417), .Y(n854));
  OAI22X1 g600(.A0(n423), .A1(n422), .B0(n428), .B1(n429), .Y(n855));
  NOR4X1  g601(.A(n854), .B(n853), .C(n852), .D(n855), .Y(n856));
  OAI22X1 g602(.A0(n338), .A1(n337), .B0(n343), .B1(n344), .Y(n857));
  OAI22X1 g603(.A0(n350), .A1(n349), .B0(n355), .B1(n356), .Y(n858));
  OAI22X1 g604(.A0(n314), .A1(n312), .B0(n319), .B1(n320), .Y(n859));
  OAI22X1 g605(.A0(n326), .A1(n325), .B0(n331), .B1(n332), .Y(n860));
  NOR4X1  g606(.A(n859), .B(n858), .C(n857), .D(n860), .Y(n861));
  OAI22X1 g607(.A0(n288), .A1(n286), .B0(n293), .B1(n295), .Y(n862));
  OAI22X1 g608(.A0(n301), .A1(n300), .B0(n306), .B1(n307), .Y(n863));
  OAI22X1 g609(.A0(n259), .A1(n254), .B0(n266), .B1(n268), .Y(n864));
  OAI22X1 g610(.A0(n275), .A1(n273), .B0(n280), .B1(n281), .Y(n865));
  NOR4X1  g611(.A(n864), .B(n863), .C(n862), .D(n865), .Y(n866));
  NAND4X1 g612(.A(n861), .B(n856), .C(n851), .D(n866), .Y(U1390));
  OAI22X1 g613(.A0(n387), .A1(n390), .B0(n396), .B1(n393), .Y(n868));
  OAI22X1 g614(.A0(n399), .A1(n402), .B0(n408), .B1(n405), .Y(n869));
  OAI22X1 g615(.A0(n363), .A1(n366), .B0(n372), .B1(n369), .Y(n870));
  OAI22X1 g616(.A0(n375), .A1(n378), .B0(n384), .B1(n381), .Y(n871));
  NOR4X1  g617(.A(n870), .B(n869), .C(n868), .D(n871), .Y(n872));
  OAI22X1 g618(.A0(n435), .A1(n438), .B0(n444), .B1(n441), .Y(n873));
  OAI22X1 g619(.A0(n447), .A1(n450), .B0(n456), .B1(n453), .Y(n874));
  OAI22X1 g620(.A0(n411), .A1(n414), .B0(n420), .B1(n417), .Y(n875));
  OAI22X1 g621(.A0(n423), .A1(n426), .B0(n432), .B1(n429), .Y(n876));
  NOR4X1  g622(.A(n875), .B(n874), .C(n873), .D(n876), .Y(n877));
  OAI22X1 g623(.A0(n338), .A1(n341), .B0(n347), .B1(n344), .Y(n878));
  OAI22X1 g624(.A0(n350), .A1(n353), .B0(n359), .B1(n356), .Y(n879));
  OAI22X1 g625(.A0(n314), .A1(n317), .B0(n323), .B1(n320), .Y(n880));
  OAI22X1 g626(.A0(n326), .A1(n329), .B0(n335), .B1(n332), .Y(n881));
  NOR4X1  g627(.A(n880), .B(n879), .C(n878), .D(n881), .Y(n882));
  OAI22X1 g628(.A0(n288), .A1(n291), .B0(n298), .B1(n295), .Y(n883));
  OAI22X1 g629(.A0(n301), .A1(n304), .B0(n310), .B1(n307), .Y(n884));
  OAI22X1 g630(.A0(n259), .A1(n263), .B0(n271), .B1(n268), .Y(n885));
  OAI22X1 g631(.A0(n275), .A1(n278), .B0(n284), .B1(n281), .Y(n886));
  NOR4X1  g632(.A(n885), .B(n884), .C(n883), .D(n886), .Y(n887));
  NAND4X1 g633(.A(n882), .B(n877), .C(n872), .D(n887), .Y(U1389));
  INVX1   g634(.A(n681), .Y(n889));
  OAI21X1 g635(.A0(n813), .A1(n592), .B0(n556), .Y(n890));
  NAND3X1 g636(.A(n890), .B(n889), .C(n484), .Y(U1384));
  OAI21X1 g637(.A0(GAMMA_REG_1__SCAN_IN), .A1(GAMMA_REG_2__SCAN_IN), .B0(n459), .Y(n892));
  NOR4X1  g638(.A(GAMMA_REG_2__SCAN_IN), .B(START), .C(n458), .D(n473), .Y(n893));
  OAI21X1 g639(.A0(n893), .A1(n892), .B0(n472), .Y(n894));
  NOR3X1  g640(.A(n557), .B(n495), .C(n460), .Y(n895));
  AOI22X1 g641(.A0(n488), .A1(n472), .B0(n475), .B1(n496), .Y(n896));
  OAI21X1 g642(.A0(n588), .A1(n680), .B0(n896), .Y(n897));
  NOR2X1  g643(.A(n897), .B(n895), .Y(n898));
  NAND3X1 g644(.A(n686), .B(n808), .C(n680), .Y(n899));
  INVX1   g645(.A(n563), .Y(n900));
  NOR2X1  g646(.A(n584), .B(n900), .Y(n901));
  AOI21X1 g647(.A0(n899), .A1(n523), .B0(n901), .Y(n902));
  NAND4X1 g648(.A(n898), .B(n894), .C(n559), .D(n902), .Y(U1385));
  AOI21X1 g649(.A0(n686), .A1(n900), .B0(n556), .Y(n904));
  AOI21X1 g650(.A0(n496), .A1(n475), .B0(n904), .Y(n905));
  NOR2X1  g651(.A(n806), .B(n521), .Y(n906));
  NOR2X1  g652(.A(n691), .B(n719), .Y(n907));
  OAI22X1 g653(.A0(n694), .A1(n728), .B0(n521), .B1(n516), .Y(n908));
  NOR2X1  g654(.A(n908), .B(n895), .Y(n909));
  OAI21X1 g655(.A0(n485), .A1(n521), .B0(n909), .Y(n910));
  NOR4X1  g656(.A(n907), .B(n893), .C(n906), .D(n910), .Y(n911));
  NAND4X1 g657(.A(n905), .B(n830), .C(n673), .D(n911), .Y(U1386));
  INVX1   g658(.A(n683), .Y(n913));
  AOI21X1 g659(.A0(n913), .A1(n718), .B0(n516), .Y(n914));
  AOI21X1 g660(.A0(n563), .A1(n551), .B0(n914), .Y(n915));
  OAI22X1 g661(.A0(n521), .A1(n516), .B0(n474), .B1(n517), .Y(n916));
  AOI21X1 g662(.A0(n521), .A1(n505), .B0(n916), .Y(n917));
  AOI21X1 g663(.A0(n592), .A1(n523), .B0(n906), .Y(n918));
  NAND3X1 g664(.A(n918), .B(n917), .C(n485), .Y(n919));
  NOR3X1  g665(.A(n919), .B(n671), .C(n590), .Y(n920));
  NAND3X1 g666(.A(n920), .B(n915), .C(n905), .Y(U1387));
  NAND4X1 g667(.A(n479), .B(GAMMA_REG_4__SCAN_IN), .C(n459), .D(n596), .Y(n922));
  NAND3X1 g668(.A(n909), .B(n922), .C(n595), .Y(n923));
  NAND2X1 g669(.A(n923), .B(n556), .Y(n924));
  AOI21X1 g670(.A0(n826), .A1(K_1_), .B0(n539), .Y(n925));
  NOR2X1  g671(.A(DATA_OUT_REG_0__SCAN_IN), .B(K_0_), .Y(n926));
  OAI21X1 g672(.A0(n926), .A1(n925), .B0(n535), .Y(n927));
  AOI21X1 g673(.A0(n823), .A1(K_3_), .B0(n539), .Y(n928));
  OAI21X1 g674(.A0(DATA_OUT_REG_0__SCAN_IN), .A1(K_2_), .B0(n624), .Y(n929));
  OAI21X1 g675(.A0(n929), .A1(n928), .B0(DATA_OUT_REG_1__SCAN_IN), .Y(n930));
  NAND3X1 g676(.A(n930), .B(n927), .C(n592), .Y(n931));
  NOR3X1  g677(.A(n749), .B(n672), .C(n906), .Y(n932));
  AOI21X1 g678(.A0(n932), .A1(n931), .B0(n556), .Y(n933));
  NOR3X1  g679(.A(n933), .B(n907), .C(n762), .Y(n934));
  NAND4X1 g680(.A(n924), .B(n915), .C(n905), .D(n934), .Y(U1388));
endmodule


