//Converted to Combinational (Partial output: n3795) , Module name: s35932_n3795 , Timestamp: 2018-12-03T15:51:09.266841 
module s35932_n3795 ( RESET, TM1, TM0, WX4420, WX4644, WX4772, WX5937, WX6065, WX4580, WX4708, WX5873, WX6001, WX4774, WX4776, WX4778, WX4716, WX4718, WX4720, WX4722, WX4724, WX4726, WX4728, WX4730, WX4732, WX4734, WX4736, WX4738, WX4740, WX4742, WX4744, WX4746, WX4748, WX4750, WX4752, WX4754, WX4756, WX4758, WX4760, WX4762, WX4764, WX4766, WX4768, WX4770, n3795 );
input RESET, TM1, TM0, WX4420, WX4644, WX4772, WX5937, WX6065, WX4580, WX4708, WX5873, WX6001, WX4774, WX4776, WX4778, WX4716, WX4718, WX4720, WX4722, WX4724, WX4726, WX4728, WX4730, WX4732, WX4734, WX4736, WX4738, WX4740, WX4742, WX4744, WX4746, WX4748, WX4750, WX4752, WX4754, WX4756, WX4758, WX4760, WX4762, WX4764, WX4766, WX4768, WX4770;
output n3795;
wire n5827, n7912_1, n7911, n7909, n5539, n7328, n7910, n7907_1, n7902_1, n7325, n7327_1, n7904, n7906, CRC_OUT_6_3, n7324, n7326, n7903, n7905, n8052, CRC_OUT_6_2, n8050, CRC_OUT_6_1, n8048, CRC_OUT_6_0, n8046, CRC_OUT_6_31, n8111_1, CRC_OUT_6_30, n8109, CRC_OUT_6_29, n8107_1, CRC_OUT_6_28, n8105, CRC_OUT_6_27, n8103_1, CRC_OUT_6_26, n8101, CRC_OUT_6_25, n8099_1, CRC_OUT_6_24, n8097, CRC_OUT_6_23, n8095_1, CRC_OUT_6_22, n8093, CRC_OUT_6_21, n8091_1, CRC_OUT_6_20, n8089, CRC_OUT_6_19, n8087_1, CRC_OUT_6_18, n8085, CRC_OUT_6_17, n8083_1, CRC_OUT_6_16, n8081, CRC_OUT_6_15, n8080, n8078, CRC_OUT_6_14, n8076, CRC_OUT_6_13, n8074, CRC_OUT_6_12, n8072, CRC_OUT_6_11, n8070, CRC_OUT_6_10, n8069, n8067_1, CRC_OUT_6_9, n8065, CRC_OUT_6_8, n8063_1, CRC_OUT_6_7, n8061, CRC_OUT_6_6, n8059_1, CRC_OUT_6_5, n8057, CRC_OUT_6_4, n8055_1, n8054;
NOR2X1   g2249(.A(n7912_1), .B(n5827), .Y(n3795));
INVX1    g0288(.A(RESET), .Y(n5827));
MX2X1    g2248(.A(n7909), .B(n7911), .S0(TM1), .Y(n7912_1));
MX2X1    g2247(.A(n7910), .B(n7328), .S0(n5539), .Y(n7911));
MX2X1    g2245(.A(n7902_1), .B(n7907_1), .S0(n5539), .Y(n7909));
INVX1    g0000(.A(TM0), .Y(n5539));
XOR2X1   g1697(.A(n7327_1), .B(n7325), .Y(n7328));
INVX1    g2246(.A(WX4420), .Y(n7910));
XOR2X1   g2244(.A(n7906), .B(n7904), .Y(n7907_1));
INVX1    g2239(.A(CRC_OUT_6_3), .Y(n7902_1));
XOR2X1   g1694(.A(n7324), .B(WX4644), .Y(n7325));
XOR2X1   g1696(.A(WX4772), .B(n7326), .Y(n7327_1));
XOR2X1   g2241(.A(n7903), .B(WX5937), .Y(n7904));
XOR2X1   g2243(.A(WX6065), .B(n7905), .Y(n7906));
NOR2X1   g2386(.A(n8052), .B(n5827), .Y(CRC_OUT_6_3));
XOR2X1   g1693(.A(WX4580), .B(TM0), .Y(n7324));
INVX1    g1695(.A(WX4708), .Y(n7326));
XOR2X1   g2240(.A(WX5873), .B(TM0), .Y(n7903));
INVX1    g2242(.A(WX6001), .Y(n7905));
XOR2X1   g2385(.A(CRC_OUT_6_2), .B(WX4772), .Y(n8052));
NOR2X1   g2384(.A(n8050), .B(n5827), .Y(CRC_OUT_6_2));
XOR2X1   g2383(.A(CRC_OUT_6_1), .B(WX4774), .Y(n8050));
NOR2X1   g2382(.A(n8048), .B(n5827), .Y(CRC_OUT_6_1));
XOR2X1   g2381(.A(CRC_OUT_6_0), .B(WX4776), .Y(n8048));
NOR2X1   g2380(.A(n8046), .B(n5827), .Y(CRC_OUT_6_0));
XOR2X1   g2379(.A(CRC_OUT_6_31), .B(WX4778), .Y(n8046));
NOR2X1   g2445(.A(n8111_1), .B(n5827), .Y(CRC_OUT_6_31));
XOR2X1   g2444(.A(CRC_OUT_6_30), .B(WX4716), .Y(n8111_1));
NOR2X1   g2443(.A(n8109), .B(n5827), .Y(CRC_OUT_6_30));
XOR2X1   g2442(.A(CRC_OUT_6_29), .B(WX4718), .Y(n8109));
NOR2X1   g2441(.A(n8107_1), .B(n5827), .Y(CRC_OUT_6_29));
XOR2X1   g2440(.A(CRC_OUT_6_28), .B(WX4720), .Y(n8107_1));
NOR2X1   g2439(.A(n8105), .B(n5827), .Y(CRC_OUT_6_28));
XOR2X1   g2438(.A(CRC_OUT_6_27), .B(WX4722), .Y(n8105));
NOR2X1   g2437(.A(n8103_1), .B(n5827), .Y(CRC_OUT_6_27));
XOR2X1   g2436(.A(CRC_OUT_6_26), .B(WX4724), .Y(n8103_1));
NOR2X1   g2435(.A(n8101), .B(n5827), .Y(CRC_OUT_6_26));
XOR2X1   g2434(.A(CRC_OUT_6_25), .B(WX4726), .Y(n8101));
NOR2X1   g2433(.A(n8099_1), .B(n5827), .Y(CRC_OUT_6_25));
XOR2X1   g2432(.A(CRC_OUT_6_24), .B(WX4728), .Y(n8099_1));
NOR2X1   g2431(.A(n8097), .B(n5827), .Y(CRC_OUT_6_24));
XOR2X1   g2430(.A(CRC_OUT_6_23), .B(WX4730), .Y(n8097));
NOR2X1   g2429(.A(n8095_1), .B(n5827), .Y(CRC_OUT_6_23));
XOR2X1   g2428(.A(CRC_OUT_6_22), .B(WX4732), .Y(n8095_1));
NOR2X1   g2427(.A(n8093), .B(n5827), .Y(CRC_OUT_6_22));
XOR2X1   g2426(.A(CRC_OUT_6_21), .B(WX4734), .Y(n8093));
NOR2X1   g2425(.A(n8091_1), .B(n5827), .Y(CRC_OUT_6_21));
XOR2X1   g2424(.A(CRC_OUT_6_20), .B(WX4736), .Y(n8091_1));
NOR2X1   g2423(.A(n8089), .B(n5827), .Y(CRC_OUT_6_20));
XOR2X1   g2422(.A(CRC_OUT_6_19), .B(WX4738), .Y(n8089));
NOR2X1   g2421(.A(n8087_1), .B(n5827), .Y(CRC_OUT_6_19));
XOR2X1   g2420(.A(CRC_OUT_6_18), .B(WX4740), .Y(n8087_1));
NOR2X1   g2419(.A(n8085), .B(n5827), .Y(CRC_OUT_6_18));
XOR2X1   g2418(.A(CRC_OUT_6_17), .B(WX4742), .Y(n8085));
NOR2X1   g2417(.A(n8083_1), .B(n5827), .Y(CRC_OUT_6_17));
XOR2X1   g2416(.A(CRC_OUT_6_16), .B(WX4744), .Y(n8083_1));
NOR2X1   g2415(.A(n8081), .B(n5827), .Y(CRC_OUT_6_16));
XOR2X1   g2414(.A(n8080), .B(CRC_OUT_6_15), .Y(n8081));
NOR2X1   g2412(.A(n8078), .B(n5827), .Y(CRC_OUT_6_15));
XOR2X1   g2413(.A(CRC_OUT_6_31), .B(WX4746), .Y(n8080));
XOR2X1   g2411(.A(CRC_OUT_6_14), .B(WX4748), .Y(n8078));
NOR2X1   g2410(.A(n8076), .B(n5827), .Y(CRC_OUT_6_14));
XOR2X1   g2409(.A(CRC_OUT_6_13), .B(WX4750), .Y(n8076));
NOR2X1   g2408(.A(n8074), .B(n5827), .Y(CRC_OUT_6_13));
XOR2X1   g2407(.A(CRC_OUT_6_12), .B(WX4752), .Y(n8074));
NOR2X1   g2406(.A(n8072), .B(n5827), .Y(CRC_OUT_6_12));
XOR2X1   g2405(.A(CRC_OUT_6_11), .B(WX4754), .Y(n8072));
NOR2X1   g2404(.A(n8070), .B(n5827), .Y(CRC_OUT_6_11));
XOR2X1   g2403(.A(n8069), .B(CRC_OUT_6_10), .Y(n8070));
NOR2X1   g2401(.A(n8067_1), .B(n5827), .Y(CRC_OUT_6_10));
XOR2X1   g2402(.A(CRC_OUT_6_31), .B(WX4756), .Y(n8069));
XOR2X1   g2400(.A(CRC_OUT_6_9), .B(WX4758), .Y(n8067_1));
NOR2X1   g2399(.A(n8065), .B(n5827), .Y(CRC_OUT_6_9));
XOR2X1   g2398(.A(CRC_OUT_6_8), .B(WX4760), .Y(n8065));
NOR2X1   g2397(.A(n8063_1), .B(n5827), .Y(CRC_OUT_6_8));
XOR2X1   g2396(.A(CRC_OUT_6_7), .B(WX4762), .Y(n8063_1));
NOR2X1   g2395(.A(n8061), .B(n5827), .Y(CRC_OUT_6_7));
XOR2X1   g2394(.A(CRC_OUT_6_6), .B(WX4764), .Y(n8061));
NOR2X1   g2393(.A(n8059_1), .B(n5827), .Y(CRC_OUT_6_6));
XOR2X1   g2392(.A(CRC_OUT_6_5), .B(WX4766), .Y(n8059_1));
NOR2X1   g2391(.A(n8057), .B(n5827), .Y(CRC_OUT_6_5));
XOR2X1   g2390(.A(CRC_OUT_6_4), .B(WX4768), .Y(n8057));
NOR2X1   g2389(.A(n8055_1), .B(n5827), .Y(CRC_OUT_6_4));
XOR2X1   g2388(.A(n8054), .B(CRC_OUT_6_3), .Y(n8055_1));
XOR2X1   g2387(.A(CRC_OUT_6_31), .B(WX4770), .Y(n8054));

endmodule
