// Benchmark "b03_C" written by ABC on Wed Aug 05 14:36:09 2020

module b03_C ( 
    STATO_REG_0__SCAN_IN, REQUEST1, REQUEST2, REQUEST3, REQUEST4,
    CODA0_REG_2__SCAN_IN, CODA0_REG_1__SCAN_IN, CODA0_REG_0__SCAN_IN,
    CODA1_REG_2__SCAN_IN, CODA1_REG_1__SCAN_IN, CODA1_REG_0__SCAN_IN,
    CODA2_REG_2__SCAN_IN, CODA2_REG_1__SCAN_IN, CODA2_REG_0__SCAN_IN,
    CODA3_REG_2__SCAN_IN, CODA3_REG_1__SCAN_IN, CODA3_REG_0__SCAN_IN,
    GRANT_REG_3__SCAN_IN, GRANT_REG_2__SCAN_IN, GRANT_REG_1__SCAN_IN,
    GRANT_REG_0__SCAN_IN, GRANT_O_REG_3__SCAN_IN, GRANT_O_REG_2__SCAN_IN,
    GRANT_O_REG_1__SCAN_IN, GRANT_O_REG_0__SCAN_IN, RU3_REG_SCAN_IN,
    FU1_REG_SCAN_IN, FU3_REG_SCAN_IN, RU1_REG_SCAN_IN, RU4_REG_SCAN_IN,
    FU2_REG_SCAN_IN, FU4_REG_SCAN_IN, RU2_REG_SCAN_IN,
    STATO_REG_1__SCAN_IN,
    U217, U216, U215, U214, U213, U212, U211, U210, U209, U208, U207, U206,
    U229, U230, U231, U232, U233, U234, U235, U236, U237, U205, U238, U204,
    U239, U240, U241, U242, U203  );
  input  STATO_REG_0__SCAN_IN, REQUEST1, REQUEST2, REQUEST3, REQUEST4,
    CODA0_REG_2__SCAN_IN, CODA0_REG_1__SCAN_IN, CODA0_REG_0__SCAN_IN,
    CODA1_REG_2__SCAN_IN, CODA1_REG_1__SCAN_IN, CODA1_REG_0__SCAN_IN,
    CODA2_REG_2__SCAN_IN, CODA2_REG_1__SCAN_IN, CODA2_REG_0__SCAN_IN,
    CODA3_REG_2__SCAN_IN, CODA3_REG_1__SCAN_IN, CODA3_REG_0__SCAN_IN,
    GRANT_REG_3__SCAN_IN, GRANT_REG_2__SCAN_IN, GRANT_REG_1__SCAN_IN,
    GRANT_REG_0__SCAN_IN, GRANT_O_REG_3__SCAN_IN, GRANT_O_REG_2__SCAN_IN,
    GRANT_O_REG_1__SCAN_IN, GRANT_O_REG_0__SCAN_IN, RU3_REG_SCAN_IN,
    FU1_REG_SCAN_IN, FU3_REG_SCAN_IN, RU1_REG_SCAN_IN, RU4_REG_SCAN_IN,
    FU2_REG_SCAN_IN, FU4_REG_SCAN_IN, RU2_REG_SCAN_IN,
    STATO_REG_1__SCAN_IN;
  output U217, U216, U215, U214, U213, U212, U211, U210, U209, U208, U207,
    U206, U229, U230, U231, U232, U233, U234, U235, U236, U237, U205, U238,
    U204, U239, U240, U241, U242, U203;
  wire n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
    n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n93, n94, n95, n96,
    n97, n98, n100, n101, n102, n103, n105, n106, n107, n109, n110, n111,
    n113, n114, n115, n117, n118, n119, n121, n122, n123, n125, n126, n127,
    n129, n130, n131, n133, n134, n136, n137, n139, n140, n142, n143, n144,
    n145, n147, n148, n149, n151, n152, n154, n155, n157, n158, n160, n161,
    n163, n164, n166, n167, n169, n170, n172, n175, n177, n178, n180, n183;
  INVX1   g000(.A(RU4_REG_SCAN_IN), .Y(n68));
  NOR4X1  g001(.A(FU4_REG_SCAN_IN), .B(n68), .C(RU3_REG_SCAN_IN), .D(RU2_REG_SCAN_IN), .Y(n69));
  INVX1   g002(.A(RU3_REG_SCAN_IN), .Y(n70));
  NOR3X1  g003(.A(RU2_REG_SCAN_IN), .B(FU3_REG_SCAN_IN), .C(n70), .Y(n71));
  INVX1   g004(.A(RU2_REG_SCAN_IN), .Y(n72));
  NOR2X1  g005(.A(n72), .B(FU2_REG_SCAN_IN), .Y(n73));
  NOR3X1  g006(.A(n73), .B(n71), .C(n69), .Y(n74));
  INVX1   g007(.A(RU1_REG_SCAN_IN), .Y(n75));
  NAND2X1 g008(.A(n75), .B(STATO_REG_0__SCAN_IN), .Y(n76));
  NAND2X1 g009(.A(RU1_REG_SCAN_IN), .B(STATO_REG_0__SCAN_IN), .Y(n77));
  NOR2X1  g010(.A(n77), .B(FU1_REG_SCAN_IN), .Y(n78));
  INVX1   g011(.A(STATO_REG_1__SCAN_IN), .Y(n79));
  NOR4X1  g012(.A(FU2_REG_SCAN_IN), .B(FU3_REG_SCAN_IN), .C(FU1_REG_SCAN_IN), .D(FU4_REG_SCAN_IN), .Y(n80));
  NOR2X1  g013(.A(n80), .B(n79), .Y(n81));
  NOR2X1  g014(.A(n81), .B(n78), .Y(n82));
  OAI21X1 g015(.A0(n76), .A1(n74), .B0(n82), .Y(n83));
  NAND3X1 g016(.A(n83), .B(STATO_REG_1__SCAN_IN), .C(CODA1_REG_2__SCAN_IN), .Y(n84));
  INVX1   g017(.A(FU4_REG_SCAN_IN), .Y(n85));
  NAND4X1 g018(.A(n85), .B(RU4_REG_SCAN_IN), .C(n70), .D(n72), .Y(n86));
  INVX1   g019(.A(FU3_REG_SCAN_IN), .Y(n87));
  NAND3X1 g020(.A(n72), .B(n87), .C(RU3_REG_SCAN_IN), .Y(n88));
  INVX1   g021(.A(FU2_REG_SCAN_IN), .Y(n89));
  NAND2X1 g022(.A(RU2_REG_SCAN_IN), .B(n89), .Y(n90));
  NAND3X1 g023(.A(n90), .B(n88), .C(n86), .Y(n91));
  INVX1   g024(.A(STATO_REG_0__SCAN_IN), .Y(U203));
  NOR2X1  g025(.A(RU1_REG_SCAN_IN), .B(U203), .Y(n93));
  OAI22X1 g026(.A0(n77), .A1(FU1_REG_SCAN_IN), .B0(n79), .B1(n80), .Y(n94));
  AOI21X1 g027(.A0(n93), .A1(n91), .B0(n94), .Y(n95));
  NAND2X1 g028(.A(n95), .B(CODA0_REG_2__SCAN_IN), .Y(n96));
  OAI21X1 g029(.A0(RU2_REG_SCAN_IN), .A1(RU3_REG_SCAN_IN), .B0(n75), .Y(n97));
  NAND3X1 g030(.A(n97), .B(n83), .C(n79), .Y(n98));
  NAND3X1 g031(.A(n98), .B(n96), .C(n84), .Y(U217));
  NAND3X1 g032(.A(n83), .B(STATO_REG_1__SCAN_IN), .C(CODA1_REG_1__SCAN_IN), .Y(n100));
  NAND2X1 g033(.A(n95), .B(CODA0_REG_1__SCAN_IN), .Y(n101));
  AOI21X1 g034(.A0(n72), .A1(RU3_REG_SCAN_IN), .B0(RU1_REG_SCAN_IN), .Y(n102));
  NAND3X1 g035(.A(n102), .B(n83), .C(n79), .Y(n103));
  NAND3X1 g036(.A(n103), .B(n101), .C(n100), .Y(U216));
  NAND3X1 g037(.A(n83), .B(STATO_REG_1__SCAN_IN), .C(CODA1_REG_0__SCAN_IN), .Y(n105));
  NAND2X1 g038(.A(n95), .B(CODA0_REG_0__SCAN_IN), .Y(n106));
  NAND4X1 g039(.A(n79), .B(n72), .C(n75), .D(n83), .Y(n107));
  NAND3X1 g040(.A(n107), .B(n106), .C(n105), .Y(U215));
  NAND3X1 g041(.A(n83), .B(n79), .C(CODA0_REG_2__SCAN_IN), .Y(n109));
  NAND2X1 g042(.A(n95), .B(CODA1_REG_2__SCAN_IN), .Y(n110));
  NAND3X1 g043(.A(n83), .B(STATO_REG_1__SCAN_IN), .C(CODA2_REG_2__SCAN_IN), .Y(n111));
  NAND3X1 g044(.A(n111), .B(n110), .C(n109), .Y(U214));
  NAND3X1 g045(.A(n83), .B(n79), .C(CODA0_REG_1__SCAN_IN), .Y(n113));
  NAND2X1 g046(.A(n95), .B(CODA1_REG_1__SCAN_IN), .Y(n114));
  NAND3X1 g047(.A(n83), .B(STATO_REG_1__SCAN_IN), .C(CODA2_REG_1__SCAN_IN), .Y(n115));
  NAND3X1 g048(.A(n115), .B(n114), .C(n113), .Y(U213));
  NAND3X1 g049(.A(n83), .B(n79), .C(CODA0_REG_0__SCAN_IN), .Y(n117));
  NAND2X1 g050(.A(n95), .B(CODA1_REG_0__SCAN_IN), .Y(n118));
  NAND3X1 g051(.A(n83), .B(STATO_REG_1__SCAN_IN), .C(CODA2_REG_0__SCAN_IN), .Y(n119));
  NAND3X1 g052(.A(n119), .B(n118), .C(n117), .Y(U212));
  NAND3X1 g053(.A(n83), .B(n79), .C(CODA1_REG_2__SCAN_IN), .Y(n121));
  NAND2X1 g054(.A(n95), .B(CODA2_REG_2__SCAN_IN), .Y(n122));
  NAND3X1 g055(.A(n83), .B(STATO_REG_1__SCAN_IN), .C(CODA3_REG_2__SCAN_IN), .Y(n123));
  NAND3X1 g056(.A(n123), .B(n122), .C(n121), .Y(U211));
  NAND3X1 g057(.A(n83), .B(n79), .C(CODA1_REG_1__SCAN_IN), .Y(n125));
  NAND2X1 g058(.A(n95), .B(CODA2_REG_1__SCAN_IN), .Y(n126));
  NAND3X1 g059(.A(n83), .B(STATO_REG_1__SCAN_IN), .C(CODA3_REG_1__SCAN_IN), .Y(n127));
  NAND3X1 g060(.A(n127), .B(n126), .C(n125), .Y(U210));
  NAND3X1 g061(.A(n83), .B(n79), .C(CODA1_REG_0__SCAN_IN), .Y(n129));
  NAND2X1 g062(.A(n95), .B(CODA2_REG_0__SCAN_IN), .Y(n130));
  NAND3X1 g063(.A(n83), .B(STATO_REG_1__SCAN_IN), .C(CODA3_REG_0__SCAN_IN), .Y(n131));
  NAND3X1 g064(.A(n131), .B(n130), .C(n129), .Y(U209));
  NAND2X1 g065(.A(n95), .B(CODA3_REG_2__SCAN_IN), .Y(n133));
  NAND3X1 g066(.A(n83), .B(n79), .C(CODA2_REG_2__SCAN_IN), .Y(n134));
  NAND2X1 g067(.A(n134), .B(n133), .Y(U208));
  NAND2X1 g068(.A(n95), .B(CODA3_REG_1__SCAN_IN), .Y(n136));
  NAND3X1 g069(.A(n83), .B(n79), .C(CODA2_REG_1__SCAN_IN), .Y(n137));
  NAND2X1 g070(.A(n137), .B(n136), .Y(U207));
  NAND2X1 g071(.A(n95), .B(CODA3_REG_0__SCAN_IN), .Y(n139));
  NAND3X1 g072(.A(n83), .B(n79), .C(CODA2_REG_0__SCAN_IN), .Y(n140));
  NAND2X1 g073(.A(n140), .B(n139), .Y(U206));
  INVX1   g074(.A(CODA0_REG_1__SCAN_IN), .Y(n142));
  INVX1   g075(.A(CODA0_REG_0__SCAN_IN), .Y(n143));
  NAND4X1 g076(.A(n143), .B(n142), .C(CODA0_REG_2__SCAN_IN), .D(n81), .Y(n144));
  OAI21X1 g077(.A0(n80), .A1(n79), .B0(GRANT_REG_3__SCAN_IN), .Y(n145));
  NAND2X1 g078(.A(n145), .B(n144), .Y(U229));
  INVX1   g079(.A(CODA0_REG_2__SCAN_IN), .Y(n147));
  NAND4X1 g080(.A(n143), .B(CODA0_REG_1__SCAN_IN), .C(n147), .D(n81), .Y(n148));
  OAI21X1 g081(.A0(n80), .A1(n79), .B0(GRANT_REG_2__SCAN_IN), .Y(n149));
  NAND2X1 g082(.A(n149), .B(n148), .Y(U230));
  NAND4X1 g083(.A(CODA0_REG_0__SCAN_IN), .B(n142), .C(n147), .D(n81), .Y(n151));
  OAI21X1 g084(.A0(n80), .A1(n79), .B0(GRANT_REG_1__SCAN_IN), .Y(n152));
  NAND2X1 g085(.A(n152), .B(n151), .Y(U231));
  NAND4X1 g086(.A(CODA0_REG_0__SCAN_IN), .B(CODA0_REG_1__SCAN_IN), .C(CODA0_REG_2__SCAN_IN), .D(n81), .Y(n154));
  OAI21X1 g087(.A0(n80), .A1(n79), .B0(GRANT_REG_0__SCAN_IN), .Y(n155));
  NAND2X1 g088(.A(n155), .B(n154), .Y(U232));
  INVX1   g089(.A(GRANT_O_REG_3__SCAN_IN), .Y(n157));
  NAND2X1 g090(.A(GRANT_REG_3__SCAN_IN), .B(STATO_REG_0__SCAN_IN), .Y(n158));
  OAI21X1 g091(.A0(n157), .A1(STATO_REG_0__SCAN_IN), .B0(n158), .Y(U233));
  INVX1   g092(.A(GRANT_O_REG_2__SCAN_IN), .Y(n160));
  NAND2X1 g093(.A(GRANT_REG_2__SCAN_IN), .B(STATO_REG_0__SCAN_IN), .Y(n161));
  OAI21X1 g094(.A0(n160), .A1(STATO_REG_0__SCAN_IN), .B0(n161), .Y(U234));
  INVX1   g095(.A(GRANT_O_REG_1__SCAN_IN), .Y(n163));
  NAND2X1 g096(.A(GRANT_REG_1__SCAN_IN), .B(STATO_REG_0__SCAN_IN), .Y(n164));
  OAI21X1 g097(.A0(n163), .A1(STATO_REG_0__SCAN_IN), .B0(n164), .Y(U235));
  INVX1   g098(.A(GRANT_O_REG_0__SCAN_IN), .Y(n166));
  NAND2X1 g099(.A(GRANT_REG_0__SCAN_IN), .B(STATO_REG_0__SCAN_IN), .Y(n167));
  OAI21X1 g100(.A0(n166), .A1(STATO_REG_0__SCAN_IN), .B0(n167), .Y(U236));
  INVX1   g101(.A(REQUEST3), .Y(n169));
  NAND2X1 g102(.A(RU3_REG_SCAN_IN), .B(STATO_REG_0__SCAN_IN), .Y(n170));
  OAI21X1 g103(.A0(n169), .A1(STATO_REG_0__SCAN_IN), .B0(n170), .Y(U237));
  INVX1   g104(.A(FU1_REG_SCAN_IN), .Y(n172));
  OAI21X1 g105(.A0(n172), .A1(STATO_REG_0__SCAN_IN), .B0(n77), .Y(U205));
  OAI21X1 g106(.A0(n87), .A1(STATO_REG_0__SCAN_IN), .B0(n170), .Y(U238));
  INVX1   g107(.A(REQUEST1), .Y(n175));
  OAI21X1 g108(.A0(n175), .A1(STATO_REG_0__SCAN_IN), .B0(n77), .Y(U204));
  INVX1   g109(.A(REQUEST4), .Y(n177));
  NAND2X1 g110(.A(RU4_REG_SCAN_IN), .B(STATO_REG_0__SCAN_IN), .Y(n178));
  OAI21X1 g111(.A0(n177), .A1(STATO_REG_0__SCAN_IN), .B0(n178), .Y(U239));
  NAND2X1 g112(.A(RU2_REG_SCAN_IN), .B(STATO_REG_0__SCAN_IN), .Y(n180));
  OAI21X1 g113(.A0(n89), .A1(STATO_REG_0__SCAN_IN), .B0(n180), .Y(U240));
  OAI21X1 g114(.A0(n85), .A1(STATO_REG_0__SCAN_IN), .B0(n178), .Y(U241));
  INVX1   g115(.A(REQUEST2), .Y(n183));
  OAI21X1 g116(.A0(n183), .A1(STATO_REG_0__SCAN_IN), .B0(n180), .Y(U242));
endmodule


