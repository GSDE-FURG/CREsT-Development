//Benchmark atmr_5xp11

module atmr_5xp11(i0, i1, i2, i3, i4, i5, i6, z0, z1, z2, z3, z4, z5, z6, z7, z8, z9);
 input i0, i1, i2, i3, i4, i5, i6;
 output z0, z1, z2, z3, z4, z5, z6, z7, z8, z9;
 wire ori_n18_, ori_n19_, ori_n20_, ori_n21_, ori_n22_, ori_n23_, ori_n24_, ori_n25_, ori_n26_, ori_n27_, ori_n28_, ori_n29_, ori_n30_, ori_n31_, ori_n32_, ori_n34_, ori_n35_, ori_n36_, ori_n37_, ori_n38_, ori_n39_, ori_n40_, ori_n41_, ori_n42_, ori_n43_, ori_n44_, ori_n45_, ori_n46_, ori_n47_, ori_n48_, ori_n49_, ori_n50_, ori_n51_, ori_n52_, ori_n53_, ori_n54_, ori_n55_, ori_n56_, ori_n58_, ori_n59_, ori_n61_, ori_n63_, ori_n66_, ori_n67_, ori_n68_, ori_n70_, ori_n71_, ori_n73_, ori_n74_, ori_n75_, ori_n76_, ori_n77_, ori_n78_, ori_n79_, ori_n80_, ori_n81_, ori_n82_, ori_n83_, ori_n85_, ori_n86_, ori_n87_, ori_n88_, ori_n89_, mai_n18_, mai_n19_, mai_n20_, mai_n21_, mai_n22_, mai_n23_, mai_n24_, mai_n25_, mai_n26_, mai_n27_, mai_n28_, mai_n30_, mai_n31_, mai_n32_, mai_n33_, mai_n34_, mai_n35_, mai_n36_, mai_n37_, mai_n38_, mai_n39_, mai_n40_, mai_n41_, mai_n43_, mai_n45_, mai_n46_, mai_n50_, mai_n52_, mai_n53_, mai_n54_, mai_n55_, mai_n57_, mai_n58_, mai_n59_, mai_n60_, mai_n61_, mai_n62_, mai_n63_, mai_n64_, men_n18_, men_n19_, men_n20_, men_n21_, men_n22_, men_n23_, men_n24_, men_n25_, men_n26_, men_n27_, men_n28_, men_n29_, men_n31_, men_n32_, men_n33_, men_n34_, men_n35_, men_n36_, men_n37_, men_n38_, men_n39_, men_n40_, men_n42_, men_n45_, men_n46_, men_n49_, men_n51_, men_n53_, men_n54_, men_n55_, men_n56_, men_n57_, men_n59_, men_n60_, zori10, zmaior0, zmenor0, zori11, zmaior1, zmenor1, zori12, zmaior2, zmenor2, zori13, zmaior3, zmenor3, zori14, zmaior4, zmenor4, zori15, zmaior5, zmenor5, zori16, zmaior6, zmenor6, zori17, zmaior7, zmenor7, zori18, zmaior8, zmenor8, zori19, zmaior9, zmenor9;
  INV        o00(.A(i1), .Y(ori_n18_));
  INV        o01(.A(i3), .Y(ori_n19_));
  NA2        o02(.A(ori_n19_), .B(ori_n18_), .Y(ori_n20_));
  NO2        o03(.A(i4), .B(i1), .Y(ori_n21_));
  NA2        o04(.A(i5), .B(i2), .Y(ori_n22_));
  NO2        o05(.A(ori_n22_), .B(ori_n21_), .Y(ori_n23_));
  INV        o06(.A(i6), .Y(ori_n24_));
  OAI210     o07(.A0(i4), .A1(i3), .B0(i1), .Y(ori_n25_));
  NA2        o08(.A(ori_n25_), .B(ori_n24_), .Y(ori_n26_));
  OAI210     o09(.A0(ori_n26_), .A1(ori_n23_), .B0(ori_n20_), .Y(ori_n27_));
  NO2        o10(.A(i5), .B(i4), .Y(ori_n28_));
  OAI210     o11(.A0(i5), .A1(i2), .B0(i4), .Y(ori_n29_));
  OA220      o12(.A0(ori_n29_), .A1(ori_n19_), .B0(ori_n28_), .B1(ori_n18_), .Y(ori_n30_));
  NA2        o13(.A(i3), .B(i1), .Y(ori_n31_));
  OAI210     o14(.A0(ori_n30_), .A1(ori_n24_), .B0(ori_n31_), .Y(ori_n32_));
  MUX2       o15(.S(i0), .A(ori_n32_), .B(ori_n27_), .Y(zori10));
  INV        o16(.A(i0), .Y(ori_n34_));
  OAI210     o17(.A0(ori_n28_), .A1(ori_n24_), .B0(ori_n34_), .Y(ori_n35_));
  INV        o18(.A(i4), .Y(ori_n36_));
  AOI210     o19(.A0(i5), .A1(i2), .B0(i6), .Y(ori_n37_));
  NA2        o20(.A(ori_n37_), .B(ori_n36_), .Y(ori_n38_));
  AOI210     o21(.A0(ori_n38_), .A1(ori_n35_), .B0(ori_n18_), .Y(ori_n39_));
  NA2        o22(.A(i4), .B(i2), .Y(ori_n40_));
  NA2        o23(.A(i6), .B(ori_n18_), .Y(ori_n41_));
  AOI210     o24(.A0(ori_n40_), .A1(ori_n34_), .B0(ori_n41_), .Y(ori_n42_));
  OAI210     o25(.A0(ori_n42_), .A1(ori_n39_), .B0(ori_n19_), .Y(ori_n43_));
  AOI210     o26(.A0(i4), .A1(i0), .B0(ori_n18_), .Y(ori_n44_));
  NA2        o27(.A(i2), .B(i0), .Y(ori_n45_));
  NA2        o28(.A(i5), .B(i4), .Y(ori_n46_));
  OAI210     o29(.A0(ori_n46_), .A1(ori_n45_), .B0(ori_n24_), .Y(ori_n47_));
  OR2        o30(.A(i4), .B(i0), .Y(ori_n48_));
  AN2        o31(.A(i6), .B(i1), .Y(ori_n49_));
  NO2        o32(.A(i1), .B(i0), .Y(ori_n50_));
  AOI220     o33(.A0(ori_n50_), .A1(ori_n29_), .B0(ori_n49_), .B1(ori_n48_), .Y(ori_n51_));
  OAI210     o34(.A0(ori_n47_), .A1(ori_n44_), .B0(ori_n51_), .Y(ori_n52_));
  OAI210     o35(.A0(ori_n20_), .A1(ori_n36_), .B0(ori_n31_), .Y(ori_n53_));
  INV        o36(.A(i5), .Y(ori_n54_));
  AOI210     o37(.A0(ori_n45_), .A1(ori_n24_), .B0(ori_n54_), .Y(ori_n55_));
  AOI220     o38(.A0(ori_n55_), .A1(ori_n53_), .B0(ori_n52_), .B1(i3), .Y(ori_n56_));
  NA2        o39(.A(ori_n56_), .B(ori_n43_), .Y(zori11));
  NO2        o40(.A(i6), .B(i1), .Y(ori_n58_));
  OAI210     o41(.A0(ori_n40_), .A1(ori_n54_), .B0(ori_n58_), .Y(ori_n59_));
  NOi31      o42(.An(ori_n59_), .B(ori_n19_), .C(ori_n34_), .Y(zori13));
  NA3        o43(.A(ori_n38_), .B(i1), .C(i0), .Y(ori_n61_));
  AOI210     o44(.A0(ori_n61_), .A1(ori_n19_), .B0(zori13), .Y(zori12));
  NO2        o45(.A(i5), .B(i2), .Y(ori_n63_));
  NOi21      o46(.An(ori_n22_), .B(ori_n63_), .Y(zori14));
  INV        o47(.A(i2), .Y(zori15));
  NA2        o48(.A(ori_n28_), .B(i2), .Y(ori_n66_));
  XO2        o49(.A(zori14), .B(i6), .Y(ori_n67_));
  NA2        o50(.A(ori_n67_), .B(ori_n66_), .Y(ori_n68_));
  OAI210     o51(.A0(ori_n66_), .A1(ori_n24_), .B0(ori_n68_), .Y(zori16));
  NA2        o52(.A(ori_n54_), .B(i2), .Y(ori_n70_));
  NA2        o53(.A(ori_n70_), .B(i4), .Y(ori_n71_));
  NA2        o54(.A(ori_n71_), .B(ori_n66_), .Y(zori17));
  NO2        o55(.A(i6), .B(ori_n34_), .Y(ori_n73_));
  NO2        o56(.A(ori_n24_), .B(i0), .Y(ori_n74_));
  AOI220     o57(.A0(ori_n74_), .A1(ori_n29_), .B0(ori_n73_), .B1(ori_n40_), .Y(ori_n75_));
  NO2        o58(.A(ori_n75_), .B(i1), .Y(ori_n76_));
  AOI220     o59(.A0(ori_n74_), .A1(ori_n54_), .B0(ori_n37_), .B1(i0), .Y(ori_n77_));
  NO2        o60(.A(ori_n77_), .B(i4), .Y(ori_n78_));
  NO3        o61(.A(i5), .B(zori15), .C(i1), .Y(ori_n79_));
  NO3        o62(.A(ori_n79_), .B(ori_n49_), .C(ori_n34_), .Y(ori_n80_));
  NO4        o63(.A(ori_n80_), .B(ori_n74_), .C(ori_n50_), .D(ori_n36_), .Y(ori_n81_));
  OAI210     o64(.A0(i6), .A1(i2), .B0(i5), .Y(ori_n82_));
  NO4        o65(.A(ori_n82_), .B(ori_n74_), .C(ori_n73_), .D(ori_n21_), .Y(ori_n83_));
  OR4        o66(.A(ori_n83_), .B(ori_n81_), .C(ori_n78_), .D(ori_n76_), .Y(zori18));
  NA2        o67(.A(ori_n82_), .B(ori_n36_), .Y(ori_n85_));
  AOI210     o68(.A0(ori_n70_), .A1(ori_n46_), .B0(ori_n37_), .Y(ori_n86_));
  NOi21      o69(.An(ori_n85_), .B(ori_n86_), .Y(ori_n87_));
  NO2        o70(.A(ori_n37_), .B(ori_n29_), .Y(ori_n88_));
  NA2        o71(.A(ori_n85_), .B(ori_n18_), .Y(ori_n89_));
  OAI220     o72(.A0(ori_n89_), .A1(ori_n88_), .B0(ori_n87_), .B1(ori_n18_), .Y(zori19));
  INV        m00(.A(i5), .Y(mai_n18_));
  INV        m01(.A(i0), .Y(mai_n19_));
  INV        m02(.A(i1), .Y(mai_n20_));
  AOI210     m03(.A0(i6), .A1(i4), .B0(i3), .Y(mai_n21_));
  NA2        m04(.A(i6), .B(i3), .Y(mai_n22_));
  NA2        m05(.A(i4), .B(i2), .Y(mai_n23_));
  OAI220     m06(.A0(mai_n23_), .A1(mai_n22_), .B0(mai_n21_), .B1(mai_n20_), .Y(mai_n24_));
  NA2        m07(.A(mai_n24_), .B(mai_n19_), .Y(mai_n25_));
  NO3        m08(.A(i6), .B(i4), .C(i3), .Y(mai_n26_));
  NOi21      m09(.An(mai_n22_), .B(mai_n19_), .Y(mai_n27_));
  OAI210     m10(.A0(mai_n26_), .A1(mai_n20_), .B0(mai_n27_), .Y(mai_n28_));
  NA3        m11(.A(mai_n28_), .B(mai_n25_), .C(mai_n18_), .Y(zmaior0));
  INV        m12(.A(i3), .Y(mai_n30_));
  INV        m13(.A(i6), .Y(mai_n31_));
  NA3        m14(.A(i5), .B(i4), .C(i2), .Y(mai_n32_));
  AOI210     m15(.A0(mai_n32_), .A1(mai_n31_), .B0(mai_n19_), .Y(mai_n33_));
  OAI210     m16(.A0(i5), .A1(i2), .B0(i4), .Y(mai_n34_));
  NO2        m17(.A(mai_n34_), .B(mai_n31_), .Y(mai_n35_));
  OAI210     m18(.A0(mai_n35_), .A1(mai_n33_), .B0(mai_n20_), .Y(mai_n36_));
  OR2        m19(.A(i5), .B(i4), .Y(mai_n37_));
  AOI210     m20(.A0(mai_n37_), .A1(i6), .B0(i0), .Y(mai_n38_));
  AOI210     m21(.A0(i5), .A1(i2), .B0(i4), .Y(mai_n39_));
  NOi21      m22(.An(mai_n39_), .B(i6), .Y(mai_n40_));
  OAI210     m23(.A0(mai_n40_), .A1(mai_n38_), .B0(i1), .Y(mai_n41_));
  NA3        m24(.A(mai_n41_), .B(mai_n36_), .C(mai_n30_), .Y(zmaior1));
  NA2        m25(.A(i1), .B(i0), .Y(mai_n43_));
  OAI210     m26(.A0(mai_n43_), .A1(mai_n40_), .B0(mai_n30_), .Y(zmaior2));
  INV        m27(.A(i2), .Y(mai_n45_));
  AOI210     m28(.A0(i5), .A1(mai_n45_), .B0(i6), .Y(mai_n46_));
  OAI210     m29(.A0(i5), .A1(mai_n45_), .B0(mai_n46_), .Y(zmaior4));
  NA2        m30(.A(mai_n31_), .B(i2), .Y(zmaior5));
  OAI210     m31(.A0(mai_n23_), .A1(i5), .B0(mai_n46_), .Y(zmaior6));
  INV        m32(.A(i4), .Y(mai_n50_));
  OAI210     m33(.A0(i5), .A1(mai_n45_), .B0(mai_n50_), .Y(zmaior7));
  OAI210     m34(.A0(mai_n39_), .A1(mai_n20_), .B0(mai_n32_), .Y(mai_n52_));
  NA2        m35(.A(mai_n52_), .B(mai_n31_), .Y(mai_n53_));
  NA2        m36(.A(mai_n37_), .B(i1), .Y(mai_n54_));
  NA3        m37(.A(mai_n54_), .B(mai_n34_), .C(i6), .Y(mai_n55_));
  NA3        m38(.A(mai_n55_), .B(mai_n53_), .C(mai_n19_), .Y(zmaior8));
  NA2        m39(.A(i5), .B(i2), .Y(mai_n57_));
  OAI210     m40(.A0(i5), .A1(i2), .B0(i6), .Y(mai_n58_));
  NA3        m41(.A(mai_n58_), .B(mai_n57_), .C(i4), .Y(mai_n59_));
  NA2        m42(.A(mai_n31_), .B(mai_n45_), .Y(mai_n60_));
  NA3        m43(.A(mai_n60_), .B(i5), .C(mai_n50_), .Y(mai_n61_));
  NO2        m44(.A(i5), .B(i2), .Y(mai_n62_));
  NO2        m45(.A(i3), .B(i0), .Y(mai_n63_));
  AOI210     m46(.A0(mai_n63_), .A1(mai_n62_), .B0(i1), .Y(mai_n64_));
  NA3        m47(.A(mai_n64_), .B(mai_n61_), .C(mai_n59_), .Y(zmaior9));
  BUFFER     m48(.A(i3), .Y(zmaior3));
  INV        u00(.A(i1), .Y(men_n18_));
  INV        u01(.A(i3), .Y(men_n19_));
  NO3        u02(.A(i6), .B(i4), .C(i2), .Y(men_n20_));
  OAI210     u03(.A0(men_n20_), .A1(men_n18_), .B0(men_n19_), .Y(men_n21_));
  INV        u04(.A(i0), .Y(men_n22_));
  NA2        u05(.A(i4), .B(i2), .Y(men_n23_));
  NO2        u06(.A(i6), .B(i1), .Y(men_n24_));
  AOI210     u07(.A0(men_n24_), .A1(men_n23_), .B0(men_n22_), .Y(men_n25_));
  AOI210     u08(.A0(i6), .A1(i4), .B0(i1), .Y(men_n26_));
  AOI210     u09(.A0(i6), .A1(i1), .B0(i0), .Y(men_n27_));
  OAI210     u10(.A0(men_n26_), .A1(men_n19_), .B0(men_n27_), .Y(men_n28_));
  NA2        u11(.A(men_n28_), .B(i5), .Y(men_n29_));
  AOI210     u12(.A0(men_n25_), .A1(men_n21_), .B0(men_n29_), .Y(zmenor0));
  INV        u13(.A(i6), .Y(men_n31_));
  NA3        u14(.A(i5), .B(i4), .C(i2), .Y(men_n32_));
  NOi21      u15(.An(men_n32_), .B(i6), .Y(men_n33_));
  OAI210     u16(.A0(i5), .A1(i2), .B0(i4), .Y(men_n34_));
  OAI220     u17(.A0(men_n34_), .A1(men_n31_), .B0(men_n33_), .B1(men_n22_), .Y(men_n35_));
  AOI210     u18(.A0(i5), .A1(i2), .B0(i4), .Y(men_n36_));
  NO2        u19(.A(men_n36_), .B(men_n22_), .Y(men_n37_));
  NO3        u20(.A(i5), .B(i4), .C(i0), .Y(men_n38_));
  OAI210     u21(.A0(men_n38_), .A1(men_n31_), .B0(i1), .Y(men_n39_));
  OAI210     u22(.A0(men_n39_), .A1(men_n37_), .B0(i3), .Y(men_n40_));
  AOI210     u23(.A0(men_n35_), .A1(men_n18_), .B0(men_n40_), .Y(zmenor1));
  AO210      u24(.A0(men_n33_), .A1(men_n18_), .B0(men_n22_), .Y(men_n42_));
  NOi21      u25(.An(men_n42_), .B(men_n19_), .Y(zmenor2));
  NO2        u26(.A(men_n42_), .B(men_n19_), .Y(zmenor3));
  NOi21      u27(.An(i5), .B(i2), .Y(men_n45_));
  NOi21      u28(.An(i2), .B(i5), .Y(men_n46_));
  OA210      u29(.A0(men_n46_), .A1(men_n45_), .B0(i6), .Y(zmenor4));
  NO2        u30(.A(men_n31_), .B(i2), .Y(zmenor5));
  NO2        u31(.A(men_n23_), .B(i5), .Y(men_n49_));
  NO3        u32(.A(men_n49_), .B(men_n45_), .C(men_n31_), .Y(zmenor6));
  INV        u33(.A(i4), .Y(men_n51_));
  NO2        u34(.A(men_n46_), .B(men_n51_), .Y(zmenor7));
  OAI210     u35(.A0(men_n36_), .A1(men_n18_), .B0(men_n32_), .Y(men_n53_));
  NO2        u36(.A(i5), .B(i4), .Y(men_n54_));
  NO2        u37(.A(men_n54_), .B(men_n18_), .Y(men_n55_));
  NA2        u38(.A(men_n34_), .B(i6), .Y(men_n56_));
  OAI210     u39(.A0(men_n56_), .A1(men_n55_), .B0(i0), .Y(men_n57_));
  AOI210     u40(.A0(men_n53_), .A1(men_n31_), .B0(men_n57_), .Y(zmenor8));
  OR2        u41(.A(men_n34_), .B(men_n33_), .Y(men_n59_));
  NO2        u42(.A(men_n54_), .B(men_n20_), .Y(men_n60_));
  AOI210     u43(.A0(men_n60_), .A1(men_n59_), .B0(men_n18_), .Y(zmenor9));
  VOTADOR g0(.A(zori10), .B(zmaior0), .C(zmenor0), .Y(z0));
  VOTADOR g1(.A(zori11), .B(zmaior1), .C(zmenor1), .Y(z1));
  VOTADOR g2(.A(zori12), .B(zmaior2), .C(zmenor2), .Y(z2));
  VOTADOR g3(.A(zori13), .B(zmaior3), .C(zmenor3), .Y(z3));
  VOTADOR g4(.A(zori14), .B(zmaior4), .C(zmenor4), .Y(z4));
  VOTADOR g5(.A(zori15), .B(zmaior5), .C(zmenor5), .Y(z5));
  VOTADOR g6(.A(zori16), .B(zmaior6), .C(zmenor6), .Y(z6));
  VOTADOR g7(.A(zori17), .B(zmaior7), .C(zmenor7), .Y(z7));
  VOTADOR g8(.A(zori18), .B(zmaior8), .C(zmenor8), .Y(z8));
  VOTADOR g9(.A(zori19), .B(zmaior9), .C(zmenor9), .Y(z9));
endmodule