//Converted to Combinational , Module name: s15850 , Timestamp: 2018-12-03T15:51:04.781284 
module s15850 ( g18, g27, g109, g741, g742, g743, g744, g872, g873, g877, g881, g1712, g1960, g1961, g1696, g750, g85, g42, g1700, g102, g104, g101, g29, g28, g103, g83, g23, g922, g892, g84, g919, g1182, g925, g48, g895, g889, g1185, g41, g43, g99, g1173, g1203, g1188, g1197, g46, g31, g45, g898, g93, g913, g82, g1194, g47, g96, g910, g95, g904, g1176, g901, g44, g916, g100, g886, g30, g86, g1170, g1200, g1191, g907, g94, g1179, g1289, g1882, g312, g452, g123, g207, g713, g1153, g1209, g1744, g1558, g695, g461, g940, g976, g709, g1092, g1574, g1864, g369, g1580, g1736, g39, g1651, g1424, g1737, g1672, g1077, g1231, g774, g1104, g1304, g243, g1499, g1044, g1444, g757, g786, g1543, g552, g315, g1534, g622, g1927, g1660, g278, g1436, g718, g76, g554, g496, g981, g878, g590, g829, g1095, g704, g1265, g1786, g682, g1296, g587, g52, g646, g327, g1389, g1371, g1956, g1675, g354, g113, g639, g1684, g1639, g1791, g248, g1707, g1759, g351, g1604, g1098, g932, g1896, g736, g1019, g1362, g745, g1419, g876, g1086, g1486, g1730, g1504, g1470, g822, g583, g1678, g1766, g1801, g959, g1169, g1007, g1407, g1059, g1868, g758, g1718, g396, g1015, g38, g632, g1415, g1227, g1721, g882, g284, g426, g219, g1216, g806, g1428, g579, g1564, g1741, g225, g281, g1308, g611, g631, g1217, g1589, g1466, g1571, g1861, g1365, g1448, g1711, g1133, g1333, g962, g766, g588, g486, g471, g1397, g580, g1950, g756, g635, g1101, g549, g1041, g1669, g1368, g1531, g1458, g572, g1011, g33, g1411, g1074, g444, g1474, g1080, g1713, g333, g269, g401, g1857, g664, g965, g1400, g309, g814, g231, g557, g586, g869, g1383, g627, g1023, g259, g1361, g1327, g654, g293, g1346, g1633, g1753, g1508, g1240, g538, g416, g542, g1681, g374, g563, g1914, g530, g575, g1936, g1117, g1317, g357, g386, g1601, g553, g501, g262, g1840, g318, g1356, g794, g302, g342, g1250, g1163, g1810, g1032, g1432, g1053, g1453, g363, g330, g1157, g1357, g928, g261, g516, g254, g778, g861, g1627, g1292, g290, g1850, g770, g1583, g466, g1561, g1527, g1546, g287, g560, g617, g336, g456, g305, g345, g1771, g865, g255, g1945, g1738, g1478, g1035, g1959, g1690, g1482, g1110, g296, g1663, g700, g1762, g360, g1657, g722, g566, g1394, g1089, g883, g1071, g986, g971, g1955, g1814, g1038, g1212, g1918, g782, g1822, g237, g746, g1062, g1462, g366, g837, g599, g1854, g944, g1941, g1520, g686, g953, g1958, g1765, g1733, g1270, g1610, g1796, g1324, g1540, g1377, g1206, g491, g1849, g213, g1781, g1900, g1245, g630, g833, g1923, g936, g1215, g1314, g849, g1336, g272, g1806, g826, g1065, g1887, g968, g1845, g1137, g1891, g1255, g257, g874, g591, g731, g636, g1218, g605, g950, g1129, g857, g448, g1828, g1727, g1592, g1703, g1932, g1624, g1068, g578, g440, g476, g668, g1149, g1848, g263, g818, g1747, g802, g275, g1524, g1577, g810, g391, g658, g1386, g253, g875, g1125, g201, g1280, g1083, g650, g1636, g853, g421, g762, g956, g378, g1756, g589, g841, g1027, g1003, g1403, g1145, g1107, g1223, g406, g1811, g1642, g1047, g1654, g197, g1595, g1537, g727, g999, g798, g481, g754, g1330, g845, g790, g1512, g1490, g1166, g1056, g348, g868, g1260, g260, g258, g521, g1318, g1872, g677, g582, g1393, g1549, g947, g1834, g1598, g1121, g1321, g506, g546, g1909, g755, g1552, g584, g1687, g1586, g324, g1141, g1570, g1341, g1710, g1645, g525, g581, g1607, g321, g1275, g1311, g1615, g382, g1374, g266, g1284, g1380, g673, g1853, g411, g431, g1905, g1515, g1630, g991, g1300, g339, g256, g1750, g585, g1440, g1666, g1528, g1351, g1648, g1618, g1235, g299, g435, g1555, g995, g1621, g1113, g643, g1494, g1567, g691, g534, g1776, g569, g1160, g1360, g1050, g511, g1724, g1878, g2355, g2601, g2602, g2603, g2604, g2605, g2606, g2607, g2608, g2609, g2610, g2611, g2612, g2648, g2986, g3007, g3069, g4172, g4173, g4174, g4175, g4176, g4177, g4178, g4179, g4180, g4181, g4887, g4888, g5101, g5105, g5658, g5659, g5816, g6920, g6926, g6932, g6942, g6949, g6955, g7744, g8061, g8062, g8271, g8313, g8316, g8318, g8323, g8328, g8331, g8335, g8340, g8347, g8349, g8352, g8561, g8562, g8563, g8564, g8565, g8566, g8976, g8977, g8978, g8979, g8980, g8981, g8982, g8983, g8984, g8985, g8986, g9451, g9961, g10377, g10379, g10455, g10457, g10459, g10461, g10463, g10465, g10628, g10801, g11163, g11206, g11489, g6842, g4171, g6267, g6257, g1957, g6282, g6284, g6281, g6253, g6285, g6283, g6265, g3327, g6269, g4204, g4193, g6266, g4203, g4212, g4196, g6263, g4194, g4192, g4213, g6256, g6258, g6279, g4209, g4208, g4214, g4206, g6261, g6255, g6260, g6274, g6271, g4195, g6273, g6275, g4201, g6264, g6270, g4216, g6262, g6278, g4200, g6277, g4198, g4210, g4197, g6259, g4202, g6280, g4191, g6254, g6268, g4205, g4207, g4215, g4199, g6272, g6276, g4211, n455, n460, n465, n470, n475, n480, n485, n490, n495, n500, n505, n510, n515, n520, n525, n530, n535, n540, n545, n550, n555, n560, n565, n570, n575, n579, n584, n589, n594, n599, n604, n609, n614, n619, n624, n629, n634, n639, n644, n649, n654, n659, n664, n669, n674, n679, n684, n689, n694, n699, n704, n709, n714, n719, n724, n729, n734, n739, n744, n749, n754, n759, n764, n769, n774, n779, n784, n789, n794, n799, n804, n809, n814, n819, n824, n829, n834, n839, n844, n849, n857, n862, n867, n872, n877, n882, n887, n892, n897, n902, n907, n912, n916, n921, n926, n931, n936, n941, n946, n951, n956, n961, n966, n971, n976, n981, n986, n991, n996, n1001, n1006, n1011, n1016, n1021, n1026, n1031, n1036, n1041, n1046, n1051, n1056, n1061, n1066, n1071, n1076, n1081, n1086, n1091, n1096, n1101, n1106, n1111, n1116, n1121, n1126, n1131, n1136, n1141, n1146, n1151, n1156, n1161, n1166, n1171, n1176, n1181, n1186, n1191, n1196, n1201, n1206, n1211, n1216, n1221, n1226, n1231, n1236, n1241, n1246, n1251, n1256, n1261, n1266, n1271, n1276, n1281, n1286, n1291, n1296, n1301, n1306, n1311, n1316, n1321, n1326, n1331, n1336, n1341, n1346, n1351, n1356, n1361, n1366, n1371, n1376, n1381, n1386, n1391, n1396, n1401, n1406, n1411, n1416, n1421, n1426, n1431, n1436, n1441, n1446, n1451, n1456, n1461, n1466, n1471, n1476, n1481, n1486, n1491, n1496, n1501, n1506, n1511, n1516, n1521, n1526, n1531, n1536, n1541, n1546, n1551, n1556, n1561, n1566, n1571, n1576, n1581, n1585, n1590, n1595, n1600, n1605, n1610, n1615, n1620, n1625, n1630, n1635, n1640, n1645, n1650, n1655, n1660, n1665, n1670, n1675, n1680, n1685, n1690, n1695, n1700, n1705, n1710, n1715, n1720, n1725, n1730, n1735, n1740, n1745, n1750, n1755, n1760, n1765, n1770, n1775, n1780, n1785, n1790, n1795, n1800, n1805, n1810, n1815, n1820, n1825, n1830, n1835, n1840, n1845, n1850, n1855, n1860, n1865, n1870, n1875, n1880, n1885, n1890, n1895, n1900, n1905, n1909, n1914, n1919, n1924, n1928, n1933, n1938, n1942, n1947, n1952, n1957, n1962, n1967, n1972, n1977, n1982, n1987, n1992, n1997, n2002, n2007, n2012, n2017, n2022, n2027, n2032, n2037, n2042, n2047, n2052, n2057, n2062, n2067, n2072, n2077, n2082, n2087, n2091, n2096, n2101, n2106, n2111, n2116, n2121, n2126, n2131, n2136, n2141, n2146, n2151, n2156, n2161, n2166, n2171, n2176, n2181, n2186, n2191, n2196, n2201, n2206, n2211, n2216, n2221, n2226, n2231, n2236, n2241, n2246, n2251, n2256, n2261, n2266, n2271, n2276, n2281, n2286, n2291, n2296, n2301, n2306, n2311, n2316, n2321, n2326, n2331, n2336, n2341, n2346, n2351, n2356, n2361, n2366, n2371, n2376, n2381, n2386, n2391, n2396, n2401, n2406, n2411, n2416, n2421, n2426, n2431, n2436, n2440, n2445, n2450, n2455, n2460, n2465, n2470, n2475, n2480, n2485, n2490, n2495, n2500, n2505, n2510, n2515, n2520, n2525, n2530, n2535, n2540, n2545, n2550, n2555, n2560, n2565, n2570, n2575, n2580, n2585, n2590, n2595, n2600, n2605, n2610, n2615, n2620, n2624, n2629, n2634, n2639, n2644, n2648, n2653, n2658, n2663, n2668, n2673, n2678, n2683, n2688, n2693, n2698, n2703, n2708, n2713, n2718, n2723, n2728, n2733, n2738, n2743, n2748, n2753, n2757, n2762, n2767, n2772, n2777, n2782, n2787, n2792, n2797, n2802, n2807, n2812, n2817, n2822, n2827, n2832, n2837, n2842, n2847, n2852, n2857, n2862, n2867, n2872, n2877, n2882, n2887, n2892, n2897, n2902, n2907, n2912, n2917, n2922, n2927, n2932, n2937, n2942, n2947, n2952, n2957, n2962, n2967, n2972, n2977, n2982, n2987, n2992, n2997, n3002, n3007, n3012, n3017, n3022, n3027, n3032, n3037, n3042, n3047, n3052, n3057, n3062, n3067, n3072, n3076, n3081, n3086, n3091, n3096, n3101, n3106 );
input g88, g90, g87, g26, g92, g89, g192, g91, g126, g186, g114, g135, g148, g139, g166, g127, g143, g170, g174, g178, g182, g131, g162, g153, g158, g115, g105, g108, g32, g37, g7, g16, g36, g8, g17, g35, g9, g1, g34, g12, g4, g119, g40, g79, g49, g73, g70, g67, g64, g61, g58, g55, g18, g27, g109, g741, g742, g743, g744, g872, g873, g877, g881, g1712, g1960, g1961, g1696, g750, g85, g42, g1700, g102, g104, g101, g29, g28, g103, g83, g23, g922, g892, g84, g919, g1182, g925, g48, g895, g889, g1185, g41, g43, g99, g1173, g1203, g1188, g1197, g46, g31, g45, g898, g93, g913, g82, g1194, g47, g96, g910, g95, g904, g1176, g901, g44, g916, g100, g886, g30, g86, g1170, g1200, g1191, g907, g94, g1179, g1289, g1882, g312, g452, g123, g207, g713, g1153, g1209, g1744, g1558, g695, g461, g940, g976, g709, g1092, g1574, g1864, g369, g1580, g1736, g39, g1651, g1424, g1737, g1672, g1077, g1231, g774, g1104, g1304, g243, g1499, g1044, g1444, g757, g786, g1543, g552, g315, g1534, g622, g1927, g1660, g278, g1436, g718, g76, g554, g496, g981, g878, g590, g829, g1095, g704, g1265, g1786, g682, g1296, g587, g52, g646, g327, g1389, g1371, g1956, g1675, g354, g113, g639, g1684, g1639, g1791, g248, g1707, g1759, g351, g1604, g1098, g932, g1896, g736, g1019, g1362, g745, g1419, g876, g1086, g1486, g1730, g1504, g1470, g822, g583, g1678, g1766, g1801, g959, g1169, g1007, g1407, g1059, g1868, g758, g1718, g396, g1015, g38, g632, g1415, g1227, g1721, g882, g284, g426, g219, g1216, g806, g1428, g579, g1564, g1741, g225, g281, g1308, g611, g631, g1217, g1589, g1466, g1571, g1861, g1365, g1448, g1711, g1133, g1333, g962, g766, g588, g486, g471, g1397, g580, g1950, g756, g635, g1101, g549, g1041, g1669, g1368, g1531, g1458, g572, g1011, g33, g1411, g1074, g444, g1474, g1080, g1713, g333, g269, g401, g1857, g664, g965, g1400, g309, g814, g231, g557, g586, g869, g1383, g627, g1023, g259, g1361, g1327, g654, g293, g1346, g1633, g1753, g1508, g1240, g538, g416, g542, g1681, g374, g563, g1914, g530, g575, g1936, g1117, g1317, g357, g386, g1601, g553, g501, g262, g1840, g318, g1356, g794, g302, g342, g1250, g1163, g1810, g1032, g1432, g1053, g1453, g363, g330, g1157, g1357, g928, g261, g516, g254, g778, g861, g1627, g1292, g290, g1850, g770, g1583, g466, g1561, g1527, g1546, g287, g560, g617, g336, g456, g305, g345, g1771, g865, g255, g1945, g1738, g1478, g1035, g1959, g1690, g1482, g1110, g296, g1663, g700, g1762, g360, g1657, g722, g566, g1394, g1089, g883, g1071, g986, g971, g1955, g1814, g1038, g1212, g1918, g782, g1822, g237, g746, g1062, g1462, g366, g837, g599, g1854, g944, g1941, g1520, g686, g953, g1958, g1765, g1733, g1270, g1610, g1796, g1324, g1540, g1377, g1206, g491, g1849, g213, g1781, g1900, g1245, g630, g833, g1923, g936, g1215, g1314, g849, g1336, g272, g1806, g826, g1065, g1887, g968, g1845, g1137, g1891, g1255, g257, g874, g591, g731, g636, g1218, g605, g950, g1129, g857, g448, g1828, g1727, g1592, g1703, g1932, g1624, g1068, g578, g440, g476, g668, g1149, g1848, g263, g818, g1747, g802, g275, g1524, g1577, g810, g391, g658, g1386, g253, g875, g1125, g201, g1280, g1083, g650, g1636, g853, g421, g762, g956, g378, g1756, g589, g841, g1027, g1003, g1403, g1145, g1107, g1223, g406, g1811, g1642, g1047, g1654, g197, g1595, g1537, g727, g999, g798, g481, g754, g1330, g845, g790, g1512, g1490, g1166, g1056, g348, g868, g1260, g260, g258, g521, g1318, g1872, g677, g582, g1393, g1549, g947, g1834, g1598, g1121, g1321, g506, g546, g1909, g755, g1552, g584, g1687, g1586, g324, g1141, g1570, g1341, g1710, g1645, g525, g581, g1607, g321, g1275, g1311, g1615, g382, g1374, g266, g1284, g1380, g673, g1853, g411, g431, g1905, g1515, g1630, g991, g1300, g339, g256, g1750, g585, g1440, g1666, g1528, g1351, g1648, g1618, g1235, g299, g435, g1555, g995, g1621, g1113, g643, g1494, g1567, g691, g534, g1776, g569, g1160, g1360, g1050, g511, g1724, g1878;
output g2355, g2601, g2602, g2603, g2604, g2605, g2606, g2607, g2608, g2609, g2610, g2611, g2612, g2648, g2986, g3007, g3069, g4172, g4173, g4174, g4175, g4176, g4177, g4178, g4179, g4180, g4181, g4887, g4888, g5101, g5105, g5658, g5659, g5816, g6920, g6926, g6932, g6942, g6949, g6955, g7744, g8061, g8062, g8271, g8313, g8316, g8318, g8323, g8328, g8331, g8335, g8340, g8347, g8349, g8352, g8561, g8562, g8563, g8564, g8565, g8566, g8976, g8977, g8978, g8979, g8980, g8981, g8982, g8983, g8984, g8985, g8986, g9451, g9961, g10377, g10379, g10455, g10457, g10459, g10461, g10463, g10465, g10628, g10801, g11163, g11206, g11489, g6842, g4171, g6267, g6257, g1957, g6282, g6284, g6281, g6253, g6285, g6283, g6265, g3327, g6269, g4204, g4193, g6266, g4203, g4212, g4196, g6263, g4194, g4192, g4213, g6256, g6258, g6279, g4209, g4208, g4214, g4206, g6261, g6255, g6260, g6274, g6271, g4195, g6273, g6275, g4201, g6264, g6270, g4216, g6262, g6278, g4200, g6277, g4198, g4210, g4197, g6259, g4202, g6280, g4191, g6254, g6268, g4205, g4207, g4215, g4199, g6272, g6276, g4211, n455, n460, n465, n470, n475, n480, n485, n490, n495, n500, n505, n510, n515, n520, n525, n530, n535, n540, n545, n550, n555, n560, n565, n570, n575, n579, n584, n589, n594, n599, n604, n609, n614, n619, n624, n629, n634, n639, n644, n649, n654, n659, n664, n669, n674, n679, n684, n689, n694, n699, n704, n709, n714, n719, n724, n729, n734, n739, n744, n749, n754, n759, n764, n769, n774, n779, n784, n789, n794, n799, n804, n809, n814, n819, n824, n829, n834, n839, n844, n849, n857, n862, n867, n872, n877, n882, n887, n892, n897, n902, n907, n912, n916, n921, n926, n931, n936, n941, n946, n951, n956, n961, n966, n971, n976, n981, n986, n991, n996, n1001, n1006, n1011, n1016, n1021, n1026, n1031, n1036, n1041, n1046, n1051, n1056, n1061, n1066, n1071, n1076, n1081, n1086, n1091, n1096, n1101, n1106, n1111, n1116, n1121, n1126, n1131, n1136, n1141, n1146, n1151, n1156, n1161, n1166, n1171, n1176, n1181, n1186, n1191, n1196, n1201, n1206, n1211, n1216, n1221, n1226, n1231, n1236, n1241, n1246, n1251, n1256, n1261, n1266, n1271, n1276, n1281, n1286, n1291, n1296, n1301, n1306, n1311, n1316, n1321, n1326, n1331, n1336, n1341, n1346, n1351, n1356, n1361, n1366, n1371, n1376, n1381, n1386, n1391, n1396, n1401, n1406, n1411, n1416, n1421, n1426, n1431, n1436, n1441, n1446, n1451, n1456, n1461, n1466, n1471, n1476, n1481, n1486, n1491, n1496, n1501, n1506, n1511, n1516, n1521, n1526, n1531, n1536, n1541, n1546, n1551, n1556, n1561, n1566, n1571, n1576, n1581, n1585, n1590, n1595, n1600, n1605, n1610, n1615, n1620, n1625, n1630, n1635, n1640, n1645, n1650, n1655, n1660, n1665, n1670, n1675, n1680, n1685, n1690, n1695, n1700, n1705, n1710, n1715, n1720, n1725, n1730, n1735, n1740, n1745, n1750, n1755, n1760, n1765, n1770, n1775, n1780, n1785, n1790, n1795, n1800, n1805, n1810, n1815, n1820, n1825, n1830, n1835, n1840, n1845, n1850, n1855, n1860, n1865, n1870, n1875, n1880, n1885, n1890, n1895, n1900, n1905, n1909, n1914, n1919, n1924, n1928, n1933, n1938, n1942, n1947, n1952, n1957, n1962, n1967, n1972, n1977, n1982, n1987, n1992, n1997, n2002, n2007, n2012, n2017, n2022, n2027, n2032, n2037, n2042, n2047, n2052, n2057, n2062, n2067, n2072, n2077, n2082, n2087, n2091, n2096, n2101, n2106, n2111, n2116, n2121, n2126, n2131, n2136, n2141, n2146, n2151, n2156, n2161, n2166, n2171, n2176, n2181, n2186, n2191, n2196, n2201, n2206, n2211, n2216, n2221, n2226, n2231, n2236, n2241, n2246, n2251, n2256, n2261, n2266, n2271, n2276, n2281, n2286, n2291, n2296, n2301, n2306, n2311, n2316, n2321, n2326, n2331, n2336, n2341, n2346, n2351, n2356, n2361, n2366, n2371, n2376, n2381, n2386, n2391, n2396, n2401, n2406, n2411, n2416, n2421, n2426, n2431, n2436, n2440, n2445, n2450, n2455, n2460, n2465, n2470, n2475, n2480, n2485, n2490, n2495, n2500, n2505, n2510, n2515, n2520, n2525, n2530, n2535, n2540, n2545, n2550, n2555, n2560, n2565, n2570, n2575, n2580, n2585, n2590, n2595, n2600, n2605, n2610, n2615, n2620, n2624, n2629, n2634, n2639, n2644, n2648, n2653, n2658, n2663, n2668, n2673, n2678, n2683, n2688, n2693, n2698, n2703, n2708, n2713, n2718, n2723, n2728, n2733, n2738, n2743, n2748, n2753, n2757, n2762, n2767, n2772, n2777, n2782, n2787, n2792, n2797, n2802, n2807, n2812, n2817, n2822, n2827, n2832, n2837, n2842, n2847, n2852, n2857, n2862, n2867, n2872, n2877, n2882, n2887, n2892, n2897, n2902, n2907, n2912, n2917, n2922, n2927, n2932, n2937, n2942, n2947, n2952, n2957, n2962, n2967, n2972, n2977, n2982, n2987, n2992, n2997, n3002, n3007, n3012, n3017, n3022, n3027, n3032, n3037, n3042, n3047, n3052, n3057, n3062, n3067, n3072, n3076, n3081, n3086, n3091, n3096, n3101, n3106;
wire n1829, n1831, n1840_1, n1842, n1844, n1846, n1848, n1850_1, n1852, n1854, n1856, n1858, n1860_1, n1862, n1864, n1866, n1868, n1870_1, n1872, n1874, n1876, n1878, n1880_1, n1882, n1884, n1885_1, n1886, n1887, n1888, n1889, n1892, n1893, n1894, n1895_1, n1896, n1897, n1898, n1899, n1900_1, n1901, n1902, n1903, n1904, n1905_1, n1906, n1907, n1908, n1909_1, n1910, n1911, n1912, n1913, n1914_1, n1915, n1916, n1917, n1918, n1919_1, n1920, n1921, n1922, n1923, n1924_1, n1925, n1926, n1927, n1928_1, n1929, n1930, n1931, n1932, n1933_1, n1934, n1935, n1936, n1937, n1938_1, n1939, n1940, n1941, n1942_1, n1943, n1944, n1945, n1946, n1947_1, n1948, n1949, n1950, n1951, n1952_1, n1953, n1954, n1955, n1956, n1957_1, n1958, n1959, n1961, n1962_1, n1963, n1964, n1965, n1966, n1967_1, n1968, n1969, n1970, n1971, n1972_1, n1973, n1974, n1975, n1976, n1977_1, n1978, n1979, n1980, n1981, n1982_1, n1983, n1984, n1986, n1987_1, n1989, n1990, n1991, n1992_1, n1993, n1994, n1995, n1996, n1997_1, n1998, n1999, n2000, n2001, n2002_1, n2003, n2004, n2006, n2007_1, n2008, n2009, n2010, n2011, n2012_1, n2013, n2014, n2015, n2016, n2017_1, n2018, n2019, n2020, n2021, n2022_1, n2023, n2024, n2025, n2026, n2027_1, n2028, n2029, n2030, n2031, n2032_1, n2033, n2034, n2035, n2036, n2037_1, n2038, n2039, n2040, n2041, n2042_1, n2043, n2044, n2045, n2046, n2047_1, n2048, n2049, n2050, n2051, n2052_1, n2053, n2054, n2055, n2056, n2057_1, n2058, n2059, n2060, n2061, n2063, n2066, n2067_1, n2068, n2069, n2070, n2071, n2072_1, n2073, n2074, n2075, n2076, n2077_1, n2078, n2079, n2080, n2081, n2082_1, n2083, n2084, n2085, n2086, n2087_1, n2088, n2089, n2091_1, n2092, n2093, n2094, n2095, n2096_1, n2097, n2098, n2099, n2100, n2101_1, n2102, n2103, n2104, n2105, n2106_1, n2107, n2108, n2109, n2110, n2111_1, n2112, n2114, n2115, n2116_1, n2117, n2118, n2119, n2120, n2121_1, n2122, n2123, n2124, n2125, n2126_1, n2127, n2128, n2129, n2130, n2131_1, n2132, n2133, n2134, n2135, n2136_1, n2137, n2138, n2139, n2140, n2141_1, n2142, n2143, n2144, n2145, n2146_1, n2147, n2148, n2149, n2150, n2151_1, n2152, n2153, n2155, n2156_1, n2157, n2158, n2159, n2160, n2161_1, n2162, n2163, n2164, n2165, n2166_1, n2167, n2168, n2169, n2170, n2171_1, n2172, n2173, n2174, n2175, n2177, n2178, n2179, n2180, n2181_1, n2182, n2183, n2184, n2185, n2186_1, n2187, n2188, n2189, n2190, n2191_1, n2192, n2193, n2195, n2196_1, n2197, n2198, n2199, n2200, n2201_1, n2202, n2203, n2204, n2205, n2206_1, n2207, n2208, n2209, n2210, n2211_1, n2212, n2213, n2214, n2215, n2216_1, n2217, n2218, n2219, n2220, n2221_1, n2222, n2223, n2224, n2226_1, n2227, n2228, n2229, n2230, n2231_1, n2232, n2233, n2234, n2235, n2236_1, n2237, n2238, n2239, n2240, n2241_1, n2242, n2243, n2244, n2245, n2246_1, n2247, n2249, n2250, n2251_1, n2252, n2253, n2254, n2255, n2256_1, n2257, n2258, n2259, n2260, n2261_1, n2262, n2263, n2264, n2265, n2267, n2268, n2269, n2270, n2271_1, n2272, n2273, n2274, n2275, n2276_1, n2277, n2278, n2279, n2283, n2284, n2285, n2286_1, n2287, n2288, n2289, n2290, n2291_1, n2292, n2294, n2295, n2296_1, n2302, n2306_1, n2307, n2308, n2309, n2310, n2311_1, n2312, n2313, n2314, n2315, n2316_1, n2317, n2318, n2319, n2320, n2321_1, n2322, n2323, n2324, n2325, n2326_1, n2327, n2328, n2329, n2330, n2331_1, n2332, n2333, n2334, n2335, n2336_1, n2337, n2338, n2339, n2340, n2341_1, n2342, n2343, n2344, n2345, n2346_1, n2347, n2348, n2350, n2351_1, n2352, n2353, n2354, n2355, n2356_1, n2357, n2358, n2359, n2360, n2362, n2364, n2365, n2366_1, n2367, n2368, n2369, n2370, n2371_1, n2372, n2373, n2374, n2375, n2376_1, n2377, n2378, n2379, n2380, n2381_1, n2382, n2383, n2384, n2385, n2386_1, n2387, n2388, n2389, n2390, n2391_1, n2392, n2393, n2394, n2395, n2396_1, n2397, n2399, n2400, n2401_1, n2402, n2403, n2404, n2405, n2406_1, n2407, n2408, n2409, n2410, n2411_1, n2412, n2413, n2414, n2416_1, n2417, n2418, n2419, n2420, n2421_1, n2422, n2423, n2424, n2425, n2426_1, n2427, n2430, n2431_1, n2432, n2433, n2434, n2435, n2436_1, n2437, n2438, n2439, n2440_1, n2441, n2442, n2443, n2444, n2445_1, n2446, n2447, n2448, n2449, n2450_1, n2451, n2452, n2453, n2454, n2455_1, n2456, n2457, n2458, n2459, n2460_1, n2461, n2462, n2463, n2464, n2465_1, n2466, n2467, n2468, n2469, n2470_1, n2471, n2472, n2473, n2474, n2475_1, n2476, n2477, n2478, n2481, n2482, n2483, n2484, n2485_1, n2486, n2487, n2488, n2489, n2490_1, n2491, n2492, n2493, n2494, n2495_1, n2496, n2497, n2498, n2499, n2500_1, n2501, n2502, n2503, n2504, n2505_1, n2508, n2509, n2511, n2512, n2513, n2514, n2515_1, n2516, n2518, n2519, n2520_1, n2521, n2522, n2523, n2525_1, n2527, n2528, n2530_1, n2531, n2532, n2533, n2534, n2535_1, n2536, n2537, n2538, n2539, n2540_1, n2541, n2542, n2543, n2544, n2545_1, n2546, n2547, n2548, n2549, n2550_1, n2551, n2552, n2553, n2554, n2555_1, n2556, n2557, n2558, n2560_1, n2561, n2562, n2563, n2564, n2566, n2567, n2568, n2569, n2571, n2572, n2574, n2576, n2577, n2578, n2580_1, n2581, n2582, n2585_1, n2587, n2590_1, n2591, n2592, n2593, n2594, n2595_1, n2598, n2599, n2600_1, n2601, n2602, n2603, n2605_1, n2606, n2607, n2608, n2609, n2610_1, n2611, n2612, n2613, n2614, n2615_1, n2617, n2618, n2620_1, n2622, n2625, n2626, n2629_1, n2630, n2631, n2632, n2633, n2634_1, n2635, n2636, n2638, n2639_1, n2640, n2641, n2642, n2643, n2646, n2647, n2650, n2651, n2652, n2654, n2655, n2656, n2657, n2658_1, n2659, n2660, n2661, n2662, n2664, n2665, n2666, n2667, n2669, n2670, n2672, n2673_1, n2674, n2675, n2676, n2678_1, n2680, n2681, n2682, n2684, n2685, n2686, n2688_1, n2690, n2691, n2692, n2693_1, n2695, n2698_1, n2699, n2700, n2701, n2702, n2703_1, n2705, n2707, n2708_1, n2709, n2710, n2711, n2713_1, n2714, n2716, n2719, n2720, n2721, n2726, n2727, n2728_1, n2729, n2730, n2731, n2732, n2734, n2735, n2736, n2737, n2738_1, n2740, n2741, n2742, n2743_1, n2745, n2746, n2748_1, n2749, n2750, n2755, n2756, n2757_1, n2758, n2759, n2765, n2766, n2767_1, n2768, n2770, n2771, n2773, n2778, n2779, n2782_1, n2783, n2785, n2788, n2789, n2791, n2792_1, n2793, n2794, n2795, n2796, n2797_1, n2798, n2800, n2801, n2802_1, n2803, n2804, n2807_1, n2809, n2811, n2812_1, n2813, n2816, n2819, n2821, n2822_1, n2823, n2824, n2825, n2828, n2829, n2830, n2831, n2835, n2837_1, n2839, n2841, n2844, n2845, n2846, n2847_1, n2848, n2851, n2852_1, n2855, n2858, n2859, n2861, n2862_1, n2863, n2864, n2870, n2871, n2872_1, n2873, n2874, n2875, n2876, n2877_1, n2878, n2879, n2880, n2881, n2882_1, n2883, n2884, n2885, n2886, n2887_1, n2888, n2889, n2890, n2891, n2892_1, n2893, n2894, n2895, n2896, n2897_1, n2898, n2899, n2900, n2901, n2902_1, n2903, n2904, n2905, n2906, n2907_1, n2909, n2910, n2911, n2912_1, n2917_1, n2920, n2923, n2924, n2925, n2926, n2927_1, n2928, n2929, n2930, n2931, n2932_1, n2933, n2934, n2935, n2941, n2944, n2945, n2947_1, n2949, n2950, n2953, n2954, n2958, n2959, n2960, n2963, n2964, n2965, n2966, n2967_1, n2968, n2969, n2970, n2971, n2972_1, n2974, n2979, n2980, n2982_1, n2984, n2988, n2990, n2991, n2996, n2998, n2999, n3000, n3001, n3002_1, n3003, n3004, n3005, n3006, n3007_1, n3008, n3009, n3010, n3011, n3012_1, n3013, n3014, n3015, n3016, n3017_1, n3018, n3019, n3021, n3023, n3027_1, n3028, n3031, n3035, n3038, n3041, n3042_1, n3045, n3047_1, n3048, n3049, n3051, n3052_1, n3054, n3055, n3056, n3060, n3062_1, n3064, n3066, n3068, n3069, n3071, n3072_1, n3075, n3076_1, n3078, n3081_1, n3082, n3083, n3084, n3085, n3086_1, n3087, n3091_1, n3092, n3093, n3094, n3095, n3096_1, n3098, n3103, n3106_1, n3107, n3111, n3114, n3115, n3116, n3117, n3119, n3122, n3124, n3125, n3126, n3127, n3130, n3131, n3132, n3134, n3135, n3136, n3140, n3144, n3147, n3148, n3151, n3155, n3156, n3159, n3160, n3167, n3168, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3215, n3217, n3219, n3220, n3222, n3223, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3235, n3236, n3239, n3241, n3246, n3249, n3253, n3254, n3255, n3256, n3257, n3260, n3261, n3262, n3263, n3265, n3270, n3271, n3273, n3275, n3276, n3277, n3278, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3297, n3298, n3300, n3301, n3302, n3303, n3307, n3310, n3312, n3313, n3314, n3315, n3316, n3317, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3331, n3334, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3346, n3347, n3348, n3349, n3351, n3352, n3355, n3357, n3359, n3361, n3362, n3363, n3368, n3370, n3374, n3375, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3385, n3387, n3390, n3392, n3397, n3400, n3401, n3402, n3404, n3405, n3408, n3410, n3415, n3416, n3417, n3418, n3419, n3420, n3422, n3424, n3426, n3427, n3428, n3429, n3430, n3432, n3433, n3434, n3435, n3436, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3455, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3469, n3471, n3472, n3473, n3474, n3475, n3480, n3482, n3484, n3485, n3486, n3490, n3492, n3494, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3504, n3507, n3511, n3512, n3515, n3516, n3521, n3523, n3525, n3526, n3527, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3548, n3551, n3552, n3553, n3554, n3557, n3559, n3560, n3563, n3564, n3567, n3569, n3571, n3572, n3576, n3577, n3579, n3581, n3582, n3584, n3587, n3588, n3589, n3594, n3596, n3598, n3600, n3601, n3603, n3606, n3608, n3609, n3611, n3615, n3617, n3619, n3622, n3625, n3626, n3627, n3628, n3630, n3631, n3632, n3633, n3634, n3635, n3637, n3638, n3639, n3643, n3644, n3649, n3652, n3653, n3654, n3655, n3656, n3659, n3664, n3665, n3667, n3669, n3671, n3673, n3677, n3681, n3685, n3688, n3691, n3693, n3695, n3697, n3702, n3704, n3706, n3709, n3710, n3714, n3715, n3717, n3719, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3734, n3737, n3741, n3745, n3747, n3750, n3752, n3754, n3755, n3756, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3770, n3773, n3775;
AND2X1   g0000(.A(g742), .B(g109), .Y(n1829));
AND2X1   g0001(.A(n1829), .B(g741), .Y(g5658));
AND2X1   g0002(.A(g744), .B(g109), .Y(n1831));
AND2X1   g0003(.A(n1831), .B(g743), .Y(g5659));
INVX1    g0004(.A(g1810), .Y(g5816));
MX2X1    g0005(.A(g1654), .B(g1672), .S0(g1690), .Y(g6920));
MX2X1    g0006(.A(g1657), .B(g1675), .S0(g1690), .Y(g6926));
MX2X1    g0007(.A(g1660), .B(g1678), .S0(g1690), .Y(g6932));
MX2X1    g0008(.A(g1663), .B(g1681), .S0(g1690), .Y(g6942));
MX2X1    g0009(.A(g1666), .B(g1684), .S0(g1690), .Y(g6949));
MX2X1    g0010(.A(g1669), .B(g1687), .S0(g1690), .Y(g6955));
NOR2X1   g0011(.A(g52), .B(g82), .Y(n1840_1));
INVX1    g0012(.A(n1840_1), .Y(g8313));
NOR2X1   g0013(.A(g55), .B(g82), .Y(n1842));
INVX1    g0014(.A(n1842), .Y(g8316));
NOR2X1   g0015(.A(g58), .B(g82), .Y(n1844));
INVX1    g0016(.A(n1844), .Y(g8318));
NOR2X1   g0017(.A(g61), .B(g82), .Y(n1846));
INVX1    g0018(.A(n1846), .Y(g8323));
NOR2X1   g0019(.A(g64), .B(g82), .Y(n1848));
INVX1    g0020(.A(n1848), .Y(g8328));
NOR2X1   g0021(.A(g67), .B(g82), .Y(n1850_1));
INVX1    g0022(.A(n1850_1), .Y(g8331));
NOR2X1   g0023(.A(g70), .B(g82), .Y(n1852));
INVX1    g0024(.A(n1852), .Y(g8335));
NOR2X1   g0025(.A(g73), .B(g82), .Y(n1854));
INVX1    g0026(.A(n1854), .Y(g8340));
NOR2X1   g0027(.A(g49), .B(g82), .Y(n1856));
INVX1    g0028(.A(n1856), .Y(g8347));
NOR2X1   g0029(.A(g76), .B(g82), .Y(n1858));
INVX1    g0030(.A(n1858), .Y(g8349));
NOR2X1   g0031(.A(g79), .B(g82), .Y(n1860_1));
INVX1    g0032(.A(n1860_1), .Y(g8352));
NAND2X1  g0033(.A(g49), .B(g82), .Y(n1862));
OAI21X1  g0034(.A0(n1856), .A1(g82), .B0(n1862), .Y(g8976));
NAND2X1  g0035(.A(g52), .B(g82), .Y(n1864));
OAI21X1  g0036(.A0(n1840_1), .A1(g82), .B0(n1864), .Y(g8977));
NAND2X1  g0037(.A(g55), .B(g82), .Y(n1866));
OAI21X1  g0038(.A0(n1842), .A1(g82), .B0(n1866), .Y(g8978));
NAND2X1  g0039(.A(g58), .B(g82), .Y(n1868));
OAI21X1  g0040(.A0(n1844), .A1(g82), .B0(n1868), .Y(g8979));
NAND2X1  g0041(.A(g61), .B(g82), .Y(n1870_1));
OAI21X1  g0042(.A0(n1846), .A1(g82), .B0(n1870_1), .Y(g8980));
NAND2X1  g0043(.A(g64), .B(g82), .Y(n1872));
OAI21X1  g0044(.A0(n1848), .A1(g82), .B0(n1872), .Y(g8981));
NAND2X1  g0045(.A(g67), .B(g82), .Y(n1874));
OAI21X1  g0046(.A0(n1850_1), .A1(g82), .B0(n1874), .Y(g8982));
NAND2X1  g0047(.A(g70), .B(g82), .Y(n1876));
OAI21X1  g0048(.A0(n1852), .A1(g82), .B0(n1876), .Y(g8983));
NAND2X1  g0049(.A(g73), .B(g82), .Y(n1878));
OAI21X1  g0050(.A0(n1854), .A1(g82), .B0(n1878), .Y(g8984));
NAND2X1  g0051(.A(g76), .B(g82), .Y(n1880_1));
OAI21X1  g0052(.A0(n1858), .A1(g82), .B0(n1880_1), .Y(g8985));
NAND2X1  g0053(.A(g79), .B(g82), .Y(n1882));
OAI21X1  g0054(.A0(n1860_1), .A1(g82), .B0(n1882), .Y(g8986));
INVX1    g0055(.A(g41), .Y(n1884));
AND2X1   g0056(.A(g31), .B(g48), .Y(n1885_1));
INVX1    g0057(.A(n1885_1), .Y(n1886));
INVX1    g0058(.A(g48), .Y(n1887));
NAND2X1  g0059(.A(g30), .B(n1887), .Y(n1888));
NOR2X1   g0060(.A(g30), .B(g31), .Y(n1889));
NAND4X1  g0061(.A(n1888), .B(n1886), .C(n1884), .D(n1889), .Y(g9451));
NAND4X1  g0062(.A(n1888), .B(n1886), .C(n1884), .D(n1889), .Y(g9961));
NOR4X1   g0063(.A(g31), .B(g41), .C(n1887), .D(g30), .Y(n1892));
OR2X1    g0064(.A(g41), .B(g42), .Y(n1893));
INVX1    g0065(.A(g43), .Y(n1894));
INVX1    g0066(.A(g44), .Y(n1895_1));
NAND3X1  g0067(.A(n1895_1), .B(g45), .C(n1894), .Y(n1896));
NOR3X1   g0068(.A(n1896), .B(n1893), .C(n1887), .Y(n1897));
INVX1    g0069(.A(g30), .Y(n1898));
OAI21X1  g0070(.A0(n1898), .A1(g48), .B0(n1884), .Y(n1899));
NOR4X1   g0071(.A(n1885_1), .B(g47), .C(g46), .D(n1899), .Y(n1900_1));
INVX1    g0072(.A(g42), .Y(n1901));
NOR4X1   g0073(.A(g41), .B(n1887), .C(n1901), .D(n1896), .Y(n1902));
OAI21X1  g0074(.A0(n1902), .A1(n1897), .B0(n1900_1), .Y(n1903));
NOR4X1   g0075(.A(n1895_1), .B(g45), .C(n1894), .D(n1893), .Y(n1904));
AND2X1   g0076(.A(n1904), .B(g48), .Y(n1905_1));
INVX1    g0077(.A(g45), .Y(n1906));
NAND3X1  g0078(.A(g44), .B(n1906), .C(g43), .Y(n1907));
NOR4X1   g0079(.A(g41), .B(n1887), .C(n1901), .D(n1907), .Y(n1908));
OAI21X1  g0080(.A0(n1908), .A1(n1905_1), .B0(n1900_1), .Y(n1909_1));
OR4X1    g0081(.A(n1885_1), .B(g47), .C(g46), .D(n1899), .Y(n1910));
NAND2X1  g0082(.A(n1904), .B(g48), .Y(n1911));
OAI21X1  g0083(.A0(n1911), .A1(n1910), .B0(g1543), .Y(n1912));
NOR2X1   g0084(.A(g41), .B(g42), .Y(n1913));
NOR3X1   g0085(.A(g44), .B(n1906), .C(g43), .Y(n1914_1));
NAND3X1  g0086(.A(n1914_1), .B(n1913), .C(g48), .Y(n1915));
OAI21X1  g0087(.A0(n1910), .A1(n1915), .B0(g1586), .Y(n1916));
OAI22X1  g0088(.A0(n1912), .A1(n1909_1), .B0(n1903), .B1(n1916), .Y(n1917));
INVX1    g0089(.A(g46), .Y(n1918));
OR4X1    g0090(.A(n1885_1), .B(g47), .C(n1918), .D(n1899), .Y(n1919_1));
NAND2X1  g0091(.A(g44), .B(g45), .Y(n1920));
NAND4X1  g0092(.A(n1884), .B(g48), .C(g42), .D(n1894), .Y(n1921));
OR2X1    g0093(.A(n1921), .B(n1920), .Y(n1922));
AOI21X1  g0094(.A0(n1922), .A1(n1911), .B0(n1919_1), .Y(n1923));
NAND4X1  g0095(.A(n1884), .B(g48), .C(g42), .D(n1914_1), .Y(n1924_1));
AOI21X1  g0096(.A0(n1924_1), .A1(n1915), .B0(n1919_1), .Y(n1925));
OR4X1    g0097(.A(g41), .B(n1887), .C(n1901), .D(n1907), .Y(n1926));
NOR2X1   g0098(.A(n1919_1), .B(n1926), .Y(n1927));
NAND2X1  g0099(.A(n1895_1), .B(g45), .Y(n1928_1));
NAND4X1  g0100(.A(n1884), .B(g48), .C(g42), .D(g43), .Y(n1929));
NOR3X1   g0101(.A(n1929), .B(n1919_1), .C(n1928_1), .Y(n1930));
OR4X1    g0102(.A(n1927), .B(n1925), .C(n1923), .D(n1930), .Y(n1931));
INVX1    g0103(.A(g31), .Y(n1932));
NAND2X1  g0104(.A(n1932), .B(g48), .Y(n1933_1));
INVX1    g0105(.A(n1933_1), .Y(n1934));
NAND3X1  g0106(.A(n1884), .B(g48), .C(n1901), .Y(n1935));
NOR4X1   g0107(.A(n1895_1), .B(g45), .C(g43), .D(n1935), .Y(n1936));
NAND3X1  g0108(.A(n1884), .B(g48), .C(g42), .Y(n1937));
NOR4X1   g0109(.A(n1895_1), .B(g45), .C(g43), .D(n1937), .Y(n1938_1));
OAI21X1  g0110(.A0(n1938_1), .A1(n1936), .B0(n1900_1), .Y(n1939));
INVX1    g0111(.A(g47), .Y(n1940));
NAND3X1  g0112(.A(n1904), .B(g46), .C(g48), .Y(n1941));
OR4X1    g0113(.A(n1899), .B(n1885_1), .C(n1940), .D(n1941), .Y(n1942_1));
NAND3X1  g0114(.A(n1942_1), .B(n1939), .C(n1934), .Y(n1943));
NOR4X1   g0115(.A(n1885_1), .B(n1940), .C(g46), .D(n1899), .Y(n1944));
NAND2X1  g0116(.A(n1944), .B(n1908), .Y(n1945));
NAND2X1  g0117(.A(n1944), .B(n1897), .Y(n1946));
NAND2X1  g0118(.A(n1944), .B(n1902), .Y(n1947_1));
NAND3X1  g0119(.A(n1947_1), .B(n1946), .C(n1945), .Y(n1948));
NAND3X1  g0120(.A(g44), .B(g45), .C(g43), .Y(n1949));
NOR4X1   g0121(.A(g41), .B(n1887), .C(n1901), .D(n1949), .Y(n1950));
NOR4X1   g0122(.A(g41), .B(n1887), .C(g42), .D(n1949), .Y(n1951));
OAI21X1  g0123(.A0(n1951), .A1(n1950), .B0(n1944), .Y(n1952_1));
NAND3X1  g0124(.A(n1952_1), .B(n1909_1), .C(n1903), .Y(n1953));
NOR4X1   g0125(.A(n1948), .B(n1943), .C(n1931), .D(n1953), .Y(n1954));
NAND3X1  g0126(.A(n1950), .B(n1944), .C(g1738), .Y(n1955));
NAND3X1  g0127(.A(n1951), .B(n1944), .C(g1762), .Y(n1956));
AOI21X1  g0128(.A0(n1956), .A1(n1955), .B0(n1952_1), .Y(n1957_1));
NOR3X1   g0129(.A(n1957_1), .B(n1954), .C(n1917), .Y(n1958));
OAI21X1  g0130(.A0(n1908), .A1(n1902), .B0(n1944), .Y(n1959));
NAND3X1  g0131(.A(n1944), .B(n1908), .C(g1188), .Y(n1961));
OR4X1    g0132(.A(n1885_1), .B(n1940), .C(g46), .D(n1899), .Y(n1962_1));
NOR2X1   g0133(.A(n1962_1), .B(n1915), .Y(n1963));
NOR2X1   g0134(.A(n1962_1), .B(n1924_1), .Y(n1964));
AOI22X1  g0135(.A0(n1963), .A1(g1333), .B0(g1308), .B1(n1964), .Y(n1965));
NAND3X1  g0136(.A(n1965), .B(n1961), .C(n1948), .Y(n1966));
NOR4X1   g0137(.A(n1927), .B(n1925), .C(n1923), .D(n1930), .Y(n1967_1));
INVX1    g0138(.A(g916), .Y(n1968));
NOR3X1   g0139(.A(n1919_1), .B(n1926), .C(n1968), .Y(n1969));
INVX1    g0140(.A(g968), .Y(n1970));
NOR3X1   g0141(.A(n1919_1), .B(n1915), .C(n1970), .Y(n1971));
INVX1    g0142(.A(g944), .Y(n1972_1));
NOR3X1   g0143(.A(n1919_1), .B(n1924_1), .C(n1972_1), .Y(n1973));
NOR3X1   g0144(.A(n1973), .B(n1971), .C(n1969), .Y(n1974));
NOR4X1   g0145(.A(n1899), .B(n1885_1), .C(n1940), .D(n1941), .Y(n1975));
INVX1    g0146(.A(g281), .Y(n1976));
OR4X1    g0147(.A(n1895_1), .B(g45), .C(g43), .D(n1937), .Y(n1977_1));
NOR4X1   g0148(.A(n1936), .B(n1910), .C(n1976), .D(n1977_1), .Y(n1978));
AND2X1   g0149(.A(n1933_1), .B(g39), .Y(n1979));
NOR3X1   g0150(.A(n1979), .B(n1978), .C(n1975), .Y(n1980));
OAI21X1  g0151(.A0(n1974), .A1(n1967_1), .B0(n1980), .Y(n1981));
AOI21X1  g0152(.A0(n1966), .A1(n1948), .B0(n1981), .Y(n1982_1));
AND2X1   g0153(.A(n1982_1), .B(n1958), .Y(n1983));
AND2X1   g0154(.A(n1983), .B(n1892), .Y(n1984));
INVX1    g0155(.A(n1984), .Y(g10377));
NOR2X1   g0156(.A(n1919_1), .B(n1924_1), .Y(n1986));
AOI22X1  g0157(.A0(n1986), .A1(g947), .B0(g919), .B1(n1927), .Y(n1987_1));
NAND3X1  g0158(.A(n1950), .B(n1944), .C(g1741), .Y(n1989));
OAI21X1  g0159(.A0(g31), .A1(n1887), .B0(g40), .Y(n1990));
NOR3X1   g0160(.A(g41), .B(n1887), .C(g42), .Y(n1991));
NAND4X1  g0161(.A(g44), .B(n1906), .C(n1894), .D(n1991), .Y(n1992_1));
NAND4X1  g0162(.A(n1992_1), .B(n1900_1), .C(g284), .D(n1938_1), .Y(n1993));
NAND4X1  g0163(.A(n1990), .B(n1989), .C(n1987_1), .D(n1993), .Y(n1994));
OAI21X1  g0164(.A0(n1911), .A1(n1910), .B0(g1546), .Y(n1995));
OAI21X1  g0165(.A0(n1910), .A1(n1915), .B0(g1589), .Y(n1996));
OAI22X1  g0166(.A0(n1995), .A1(n1909_1), .B0(n1903), .B1(n1996), .Y(n1997_1));
NAND2X1  g0167(.A(n1950), .B(n1944), .Y(n1998));
NAND4X1  g0168(.A(n1998), .B(n1909_1), .C(n1903), .D(n1959), .Y(n1999));
NOR3X1   g0169(.A(n1999), .B(n1943), .C(n1931), .Y(n2000));
NAND3X1  g0170(.A(n1944), .B(n1908), .C(g1191), .Y(n2001));
NAND3X1  g0171(.A(n1944), .B(n1902), .C(g1311), .Y(n2002_1));
AOI21X1  g0172(.A0(n2002_1), .A1(n2001), .B0(n1959), .Y(n2003));
NOR4X1   g0173(.A(n2000), .B(n1997_1), .C(n1994), .D(n2003), .Y(n2004));
NAND2X1  g0174(.A(n2004), .B(n1892), .Y(g10379));
INVX1    g0175(.A(n1892), .Y(n2006));
NAND3X1  g0176(.A(n1895_1), .B(n1906), .C(g43), .Y(n2007_1));
NOR2X1   g0177(.A(n2007_1), .B(n1937), .Y(n2008));
NOR2X1   g0178(.A(n2007_1), .B(n1935), .Y(n2009));
OAI21X1  g0179(.A0(n2009), .A1(n2008), .B0(n1900_1), .Y(n2010));
AND2X1   g0180(.A(n2010), .B(n1942_1), .Y(n2011));
NAND3X1  g0181(.A(n2009), .B(n1900_1), .C(g119), .Y(n2012_1));
AND2X1   g0182(.A(n2008), .B(n1900_1), .Y(n2013));
AOI21X1  g0183(.A0(n2013), .A1(g123), .B0(n1975), .Y(n2014));
AOI21X1  g0184(.A0(n2014), .A1(n2012_1), .B0(n2011), .Y(n2015));
NAND3X1  g0185(.A(n1936), .B(n1900_1), .C(g287), .Y(n2016));
OAI21X1  g0186(.A0(n1992_1), .A1(n1910), .B0(g263), .Y(n2017_1));
AND2X1   g0187(.A(n2017_1), .B(n2016), .Y(n2018));
OAI21X1  g0188(.A0(g31), .A1(n1887), .B0(g33), .Y(n2019));
OAI21X1  g0189(.A0(n2018), .A1(n1939), .B0(n2019), .Y(n2020));
NAND4X1  g0190(.A(n1942_1), .B(n1939), .C(n1934), .D(n2010), .Y(n2021));
NAND2X1  g0191(.A(n1944), .B(n1905_1), .Y(n2022_1));
NAND4X1  g0192(.A(n1947_1), .B(n1946), .C(n1945), .D(n2022_1), .Y(n2023));
NOR4X1   g0193(.A(n2021), .B(n1953), .C(n1931), .D(n2023), .Y(n2024));
NAND3X1  g0194(.A(n1950), .B(n1944), .C(g1721), .Y(n2025));
NAND3X1  g0195(.A(n1951), .B(n1944), .C(g1744), .Y(n2026));
AOI21X1  g0196(.A0(n2026), .A1(n2025), .B0(n1952_1), .Y(n2027_1));
OR4X1    g0197(.A(n2024), .B(n2020), .C(n2015), .D(n2027_1), .Y(n2028));
INVX1    g0198(.A(g1336), .Y(n2029));
NAND3X1  g0199(.A(n1944), .B(n1908), .C(g1170), .Y(n2030));
OAI21X1  g0200(.A0(n1947_1), .A1(n2029), .B0(n2030), .Y(n2031));
NAND3X1  g0201(.A(n1944), .B(n1905_1), .C(g1194), .Y(n2032_1));
NAND3X1  g0202(.A(n1944), .B(n1897), .C(g1314), .Y(n2033));
NAND2X1  g0203(.A(n2033), .B(n2032_1), .Y(n2034));
OAI21X1  g0204(.A0(n2034), .A1(n2031), .B0(n2023), .Y(n2035));
INVX1    g0205(.A(g928), .Y(n2036));
OR2X1    g0206(.A(n1922), .B(n1919_1), .Y(n2037_1));
NOR4X1   g0207(.A(n1885_1), .B(g47), .C(n1918), .D(n1899), .Y(n2038));
NAND3X1  g0208(.A(n2038), .B(n1897), .C(g950), .Y(n2039));
OAI21X1  g0209(.A0(n2037_1), .A1(n2036), .B0(n2039), .Y(n2040));
INVX1    g0210(.A(g922), .Y(n2041));
NOR3X1   g0211(.A(n1919_1), .B(n1911), .C(n2041), .Y(n2042_1));
INVX1    g0212(.A(g971), .Y(n2043));
NOR3X1   g0213(.A(n1919_1), .B(n1924_1), .C(n2043), .Y(n2044));
INVX1    g0214(.A(g886), .Y(n2045));
NOR4X1   g0215(.A(n1919_1), .B(n1928_1), .C(n2045), .D(n1929), .Y(n2046));
INVX1    g0216(.A(g898), .Y(n2047_1));
NOR3X1   g0217(.A(n1919_1), .B(n1926), .C(n2047_1), .Y(n2048));
OR4X1    g0218(.A(n2046), .B(n2044), .C(n2042_1), .D(n2048), .Y(n2049));
OAI21X1  g0219(.A0(n2049), .A1(n2040), .B0(n1931), .Y(n2050));
AOI21X1  g0220(.A0(n1924_1), .A1(n1915), .B0(n1910), .Y(n2051));
AOI21X1  g0221(.A0(n1926), .A1(n1911), .B0(n1910), .Y(n2052_1));
NAND3X1  g0222(.A(n1905_1), .B(n1900_1), .C(g1549), .Y(n2053));
OAI21X1  g0223(.A0(n1911), .A1(n1910), .B0(g1524), .Y(n2054));
NAND2X1  g0224(.A(n2054), .B(n2053), .Y(n2055));
NAND3X1  g0225(.A(n1900_1), .B(n1897), .C(g1592), .Y(n2056));
OAI21X1  g0226(.A0(n1910), .A1(n1915), .B0(g1567), .Y(n2057_1));
NAND2X1  g0227(.A(n2057_1), .B(n2056), .Y(n2058));
AOI22X1  g0228(.A0(n2055), .A1(n2052_1), .B0(n2051), .B1(n2058), .Y(n2059));
NAND3X1  g0229(.A(n2059), .B(n2050), .C(n2035), .Y(n2060));
NOR3X1   g0230(.A(n2060), .B(n2028), .C(n2006), .Y(n2061));
INVX1    g0231(.A(n2061), .Y(g10455));
OAI21X1  g0232(.A0(n1908), .A1(n1897), .B0(n1944), .Y(n2063));
NAND3X1  g0233(.A(n1950), .B(n1944), .C(g1724), .Y(n2066));
NAND3X1  g0234(.A(n1951), .B(n1944), .C(g1747), .Y(n2067_1));
AOI21X1  g0235(.A0(n2067_1), .A1(n2066), .B0(n1952_1), .Y(n2068));
AND2X1   g0236(.A(n2009), .B(n1900_1), .Y(n2069));
AOI22X1  g0237(.A0(n2013), .A1(g4), .B0(g12), .B1(n2069), .Y(n2070));
NOR2X1   g0238(.A(n2070), .B(n2011), .Y(n2071));
NAND3X1  g0239(.A(n1936), .B(n1900_1), .C(g290), .Y(n2072_1));
OAI21X1  g0240(.A0(n1992_1), .A1(n1910), .B0(g266), .Y(n2073));
AND2X1   g0241(.A(n2073), .B(n2072_1), .Y(n2074));
OAI21X1  g0242(.A0(g31), .A1(n1887), .B0(g34), .Y(n2075));
OAI21X1  g0243(.A0(n2074), .A1(n1939), .B0(n2075), .Y(n2076));
OR4X1    g0244(.A(n2071), .B(n2068), .C(n2024), .D(n2076), .Y(n2077_1));
NOR2X1   g0245(.A(n1962_1), .B(n1926), .Y(n2078));
NOR2X1   g0246(.A(n1962_1), .B(n1911), .Y(n2079));
NOR4X1   g0247(.A(n1964), .B(n1963), .C(n2078), .D(n2079), .Y(n2080));
INVX1    g0248(.A(g1341), .Y(n2081));
NOR3X1   g0249(.A(n1962_1), .B(n1924_1), .C(n2081), .Y(n2082_1));
INVX1    g0250(.A(g1318), .Y(n2083));
NOR3X1   g0251(.A(n1962_1), .B(n1915), .C(n2083), .Y(n2084));
INVX1    g0252(.A(g1173), .Y(n2085));
NOR3X1   g0253(.A(n1962_1), .B(n1926), .C(n2085), .Y(n2086));
INVX1    g0254(.A(g1197), .Y(n2087_1));
NOR3X1   g0255(.A(n1962_1), .B(n1911), .C(n2087_1), .Y(n2088));
OR4X1    g0256(.A(n2086), .B(n2084), .C(n2082_1), .D(n2088), .Y(n2089));
INVX1    g0257(.A(g932), .Y(n2091_1));
NAND3X1  g0258(.A(n2038), .B(n1897), .C(g953), .Y(n2092));
OAI21X1  g0259(.A0(n2037_1), .A1(n2091_1), .B0(n2092), .Y(n2093));
INVX1    g0260(.A(g925), .Y(n2094));
NOR3X1   g0261(.A(n1919_1), .B(n1911), .C(n2094), .Y(n2095));
INVX1    g0262(.A(g976), .Y(n2096_1));
NOR3X1   g0263(.A(n1919_1), .B(n1924_1), .C(n2096_1), .Y(n2097));
INVX1    g0264(.A(g889), .Y(n2098));
NOR4X1   g0265(.A(n1919_1), .B(n1928_1), .C(n2098), .D(n1929), .Y(n2099));
INVX1    g0266(.A(g901), .Y(n2100));
NOR3X1   g0267(.A(n1919_1), .B(n1926), .C(n2100), .Y(n2101_1));
OR4X1    g0268(.A(n2099), .B(n2097), .C(n2095), .D(n2101_1), .Y(n2102));
OAI21X1  g0269(.A0(n2102), .A1(n2093), .B0(n1931), .Y(n2103));
NAND3X1  g0270(.A(n1905_1), .B(n1900_1), .C(g1552), .Y(n2104));
OAI21X1  g0271(.A0(n1911), .A1(n1910), .B0(g1528), .Y(n2105));
NAND2X1  g0272(.A(n2105), .B(n2104), .Y(n2106_1));
NAND3X1  g0273(.A(n1900_1), .B(n1897), .C(g1595), .Y(n2107));
OAI21X1  g0274(.A0(n1910), .A1(n1915), .B0(g1571), .Y(n2108));
NAND2X1  g0275(.A(n2108), .B(n2107), .Y(n2109));
AOI22X1  g0276(.A0(n2106_1), .A1(n2052_1), .B0(n2051), .B1(n2109), .Y(n2110));
NAND3X1  g0277(.A(n2110), .B(n2103), .C(n2397), .Y(n2111_1));
NOR3X1   g0278(.A(n2111_1), .B(n2077_1), .C(n2006), .Y(n2112));
INVX1    g0279(.A(n2112), .Y(g10457));
NAND3X1  g0280(.A(n1950), .B(n1944), .C(g1727), .Y(n2114));
NAND3X1  g0281(.A(n1951), .B(n1944), .C(g1750), .Y(n2115));
AOI21X1  g0282(.A0(n2115), .A1(n2114), .B0(n1952_1), .Y(n2116_1));
AOI22X1  g0283(.A0(n2013), .A1(g1), .B0(g9), .B1(n2069), .Y(n2117));
NOR2X1   g0284(.A(n2117), .B(n2011), .Y(n2118));
NAND3X1  g0285(.A(n1936), .B(n1900_1), .C(g293), .Y(n2119));
OAI21X1  g0286(.A0(n1992_1), .A1(n1910), .B0(g269), .Y(n2120));
AND2X1   g0287(.A(n2120), .B(n2119), .Y(n2121_1));
OAI21X1  g0288(.A0(g31), .A1(n1887), .B0(g35), .Y(n2122));
OAI21X1  g0289(.A0(n2121_1), .A1(n1939), .B0(n2122), .Y(n2123));
OR4X1    g0290(.A(n2118), .B(n2116_1), .C(n2024), .D(n2123), .Y(n2124));
INVX1    g0291(.A(g1346), .Y(n2125));
NOR3X1   g0292(.A(n1962_1), .B(n1924_1), .C(n2125), .Y(n2126_1));
INVX1    g0293(.A(g1321), .Y(n2127));
NOR3X1   g0294(.A(n1962_1), .B(n1915), .C(n2127), .Y(n2128));
INVX1    g0295(.A(g1176), .Y(n2129));
NOR3X1   g0296(.A(n1962_1), .B(n1926), .C(n2129), .Y(n2130));
INVX1    g0297(.A(g1200), .Y(n2131_1));
NOR3X1   g0298(.A(n1962_1), .B(n1911), .C(n2131_1), .Y(n2132));
OR4X1    g0299(.A(n2130), .B(n2128), .C(n2126_1), .D(n2132), .Y(n2133));
OAI21X1  g0300(.A0(n2133), .A1(n2080), .B0(n2023), .Y(n2134));
INVX1    g0301(.A(g936), .Y(n2135));
NAND3X1  g0302(.A(n2038), .B(n1897), .C(g956), .Y(n2136_1));
OAI21X1  g0303(.A0(n2037_1), .A1(n2135), .B0(n2136_1), .Y(n2137));
NAND3X1  g0304(.A(n2038), .B(n1908), .C(g904), .Y(n2138));
NOR2X1   g0305(.A(g44), .B(n1906), .Y(n2139));
NOR4X1   g0306(.A(g41), .B(n1887), .C(n1901), .D(n1894), .Y(n2140));
NAND4X1  g0307(.A(n2038), .B(n2139), .C(g892), .D(n2140), .Y(n2141_1));
NAND3X1  g0308(.A(n2038), .B(n1902), .C(g981), .Y(n2142));
NAND3X1  g0309(.A(n2142), .B(n2141_1), .C(n2138), .Y(n2143));
OAI21X1  g0310(.A0(n2143), .A1(n2137), .B0(n1931), .Y(n2144));
NAND3X1  g0311(.A(n1905_1), .B(n1900_1), .C(g1555), .Y(n2145));
OAI21X1  g0312(.A0(n1911), .A1(n1910), .B0(g1531), .Y(n2146_1));
NAND2X1  g0313(.A(n2146_1), .B(n2145), .Y(n2147));
NAND3X1  g0314(.A(n1900_1), .B(n1897), .C(g1598), .Y(n2148));
OAI21X1  g0315(.A0(n1910), .A1(n1915), .B0(g1574), .Y(n2149));
NAND2X1  g0316(.A(n2149), .B(n2148), .Y(n2150));
AOI22X1  g0317(.A0(n2147), .A1(n2052_1), .B0(n2051), .B1(n2150), .Y(n2151_1));
NAND3X1  g0318(.A(n2151_1), .B(n2144), .C(n2134), .Y(n2152));
NOR3X1   g0319(.A(n2152), .B(n2124), .C(n2006), .Y(n2153));
INVX1    g0320(.A(n2153), .Y(g10459));
NAND3X1  g0321(.A(n1950), .B(n1944), .C(g1730), .Y(n2155));
NAND3X1  g0322(.A(n1951), .B(n1944), .C(g1753), .Y(n2156_1));
AOI21X1  g0323(.A0(n2156_1), .A1(n2155), .B0(n1952_1), .Y(n2157));
NAND3X1  g0324(.A(n2009), .B(n1900_1), .C(g17), .Y(n2158));
NAND3X1  g0325(.A(n2008), .B(n1900_1), .C(g8), .Y(n2159));
AOI22X1  g0326(.A0(n2158), .A1(n2159), .B0(n2010), .B1(n1942_1), .Y(n2160));
NAND3X1  g0327(.A(n1936), .B(n1900_1), .C(g296), .Y(n2161_1));
OAI21X1  g0328(.A0(n1992_1), .A1(n1910), .B0(g272), .Y(n2162));
AND2X1   g0329(.A(n2162), .B(n2161_1), .Y(n2163));
OAI21X1  g0330(.A0(g31), .A1(n1887), .B0(g36), .Y(n2164));
OAI21X1  g0331(.A0(n2163), .A1(n1939), .B0(n2164), .Y(n2165));
OR4X1    g0332(.A(n2160), .B(n2157), .C(n2024), .D(n2165), .Y(n2166_1));
INVX1    g0333(.A(g1351), .Y(n2167));
NOR3X1   g0334(.A(n1962_1), .B(n1924_1), .C(n2167), .Y(n2168));
INVX1    g0335(.A(g1324), .Y(n2169));
NOR3X1   g0336(.A(n1962_1), .B(n1915), .C(n2169), .Y(n2170));
INVX1    g0337(.A(g1179), .Y(n2171_1));
NOR3X1   g0338(.A(n1962_1), .B(n1926), .C(n2171_1), .Y(n2172));
INVX1    g0339(.A(g1203), .Y(n2173));
NOR3X1   g0340(.A(n1962_1), .B(n1911), .C(n2173), .Y(n2174));
OR4X1    g0341(.A(n2172), .B(n2170), .C(n2168), .D(n2174), .Y(n2175));
INVX1    g0342(.A(g940), .Y(n2177));
NAND3X1  g0343(.A(n2038), .B(n1897), .C(g959), .Y(n2178));
OAI21X1  g0344(.A0(n2037_1), .A1(n2177), .B0(n2178), .Y(n2179));
NAND3X1  g0345(.A(n2038), .B(n1908), .C(g907), .Y(n2180));
NAND4X1  g0346(.A(n2038), .B(n2139), .C(g895), .D(n2140), .Y(n2181_1));
NAND3X1  g0347(.A(n2038), .B(n1902), .C(g986), .Y(n2182));
NAND3X1  g0348(.A(n2182), .B(n2181_1), .C(n2180), .Y(n2183));
OAI21X1  g0349(.A0(n2183), .A1(n2179), .B0(n1931), .Y(n2184));
NAND3X1  g0350(.A(n1905_1), .B(n1900_1), .C(g1558), .Y(n2185));
OAI21X1  g0351(.A0(n1911), .A1(n1910), .B0(g1534), .Y(n2186_1));
NAND2X1  g0352(.A(n2186_1), .B(n2185), .Y(n2187));
NAND3X1  g0353(.A(n1900_1), .B(n1897), .C(g1601), .Y(n2188));
OAI21X1  g0354(.A0(n1910), .A1(n1915), .B0(g1577), .Y(n2189));
NAND2X1  g0355(.A(n2189), .B(n2188), .Y(n2190));
AOI22X1  g0356(.A0(n2187), .A1(n2052_1), .B0(n2051), .B1(n2190), .Y(n2191_1));
NAND3X1  g0357(.A(n2191_1), .B(n2184), .C(n2362), .Y(n2192));
NOR3X1   g0358(.A(n2192), .B(n2166_1), .C(n2006), .Y(n2193));
INVX1    g0359(.A(n2193), .Y(g10461));
NAND3X1  g0360(.A(n1944), .B(n1908), .C(g1182), .Y(n2195));
NAND3X1  g0361(.A(n1944), .B(n1897), .C(g1327), .Y(n2196_1));
AOI21X1  g0362(.A0(n2196_1), .A1(n2195), .B0(n2063), .Y(n2197));
AOI21X1  g0363(.A0(n1926), .A1(n1915), .B0(n1962_1), .Y(n2198));
NOR4X1   g0364(.A(n2021), .B(n1953), .C(n1931), .D(n2198), .Y(n2199));
NAND3X1  g0365(.A(n1950), .B(n1944), .C(g1733), .Y(n2200));
NAND3X1  g0366(.A(n1951), .B(n1944), .C(g1756), .Y(n2201_1));
AOI21X1  g0367(.A0(n2201_1), .A1(n2200), .B0(n1952_1), .Y(n2202));
NOR3X1   g0368(.A(n2202), .B(n2199), .C(n2197), .Y(n2203));
NAND3X1  g0369(.A(n1905_1), .B(n1900_1), .C(g1561), .Y(n2204));
OAI21X1  g0370(.A0(n1911), .A1(n1910), .B0(g1537), .Y(n2205));
AND2X1   g0371(.A(n2205), .B(n2204), .Y(n2206_1));
NAND3X1  g0372(.A(n1900_1), .B(n1897), .C(g1604), .Y(n2207));
OAI21X1  g0373(.A0(n1910), .A1(n1915), .B0(g1580), .Y(n2208));
AND2X1   g0374(.A(n2208), .B(n2207), .Y(n2209));
OAI22X1  g0375(.A0(n2206_1), .A1(n1909_1), .B0(n1903), .B1(n2209), .Y(n2210));
NOR2X1   g0376(.A(n1919_1), .B(n1915), .Y(n2211_1));
AOI22X1  g0377(.A0(n2211_1), .A1(g962), .B0(g910), .B1(n1927), .Y(n2212));
NOR2X1   g0378(.A(n2212), .B(n1967_1), .Y(n2213));
NAND3X1  g0379(.A(n2009), .B(n1900_1), .C(g16), .Y(n2214));
NAND3X1  g0380(.A(n2008), .B(n1900_1), .C(g7), .Y(n2215));
AOI22X1  g0381(.A0(n2214), .A1(n2215), .B0(n2010), .B1(n1942_1), .Y(n2216_1));
NAND3X1  g0382(.A(n1936), .B(n1900_1), .C(g299), .Y(n2217));
OAI21X1  g0383(.A0(n1992_1), .A1(n1910), .B0(g275), .Y(n2218));
AND2X1   g0384(.A(n2218), .B(n2217), .Y(n2219));
OAI21X1  g0385(.A0(g31), .A1(n1887), .B0(g37), .Y(n2220));
OAI21X1  g0386(.A0(n2219), .A1(n1939), .B0(n2220), .Y(n2221_1));
NOR4X1   g0387(.A(n2216_1), .B(n2213), .C(n2210), .D(n2221_1), .Y(n2222));
NAND2X1  g0388(.A(n2222), .B(n2203), .Y(n2223));
NOR2X1   g0389(.A(n2223), .B(n2006), .Y(n2224));
INVX1    g0390(.A(n2224), .Y(g10463));
NAND2X1  g0391(.A(n1905_1), .B(n1900_1), .Y(n2226_1));
MX2X1    g0392(.A(g1564), .B(g1540), .S0(n2226_1), .Y(n2227));
NOR2X1   g0393(.A(n1910), .B(n1915), .Y(n2228));
MX2X1    g0394(.A(g1583), .B(g1607), .S0(n2228), .Y(n2229));
AOI22X1  g0395(.A0(n2227), .A1(n2052_1), .B0(n2051), .B1(n2229), .Y(n2230));
NAND3X1  g0396(.A(n2038), .B(n1908), .C(g913), .Y(n2231_1));
NAND3X1  g0397(.A(n2038), .B(n1897), .C(g965), .Y(n2232));
NAND2X1  g0398(.A(n2232), .B(n2231_1), .Y(n2233));
NAND2X1  g0399(.A(n2233), .B(n1931), .Y(n2234));
INVX1    g0400(.A(n1949), .Y(n2235));
NAND4X1  g0401(.A(n1944), .B(n1991), .C(g1759), .D(n2235), .Y(n2236_1));
AOI21X1  g0402(.A0(n1977_1), .A1(n1992_1), .B0(n1910), .Y(n2237));
NOR2X1   g0403(.A(n1992_1), .B(n1910), .Y(n2238));
MX2X1    g0404(.A(g278), .B(g302), .S0(n2238), .Y(n2239));
AOI22X1  g0405(.A0(n2237), .A1(n2239), .B0(n1933_1), .B1(g38), .Y(n2240));
NAND3X1  g0406(.A(n2240), .B(n2236_1), .C(n2234), .Y(n2241_1));
OR4X1    g0407(.A(n1953), .B(n1943), .C(n1931), .D(n2198), .Y(n2242));
AOI22X1  g0408(.A0(n2078), .A1(g1185), .B0(g1330), .B1(n1963), .Y(n2243));
NAND2X1  g0409(.A(n2243), .B(n2242), .Y(n2244));
NOR2X1   g0410(.A(n2244), .B(n2241_1), .Y(n2245));
AND2X1   g0411(.A(n2245), .B(n2230), .Y(n2246_1));
AND2X1   g0412(.A(n2246_1), .B(n1892), .Y(n2247));
INVX1    g0413(.A(n2247), .Y(g10465));
INVX1    g0414(.A(g109), .Y(n2249));
INVX1    g0415(.A(g883), .Y(n2250));
NOR2X1   g0416(.A(n2152), .B(n2124), .Y(n2251_1));
NOR4X1   g0417(.A(n2250), .B(g882), .C(n2249), .D(n2251_1), .Y(n2252));
AOI21X1  g0418(.A0(n2222), .A1(n2203), .B0(n2249), .Y(n2253));
INVX1    g0419(.A(g878), .Y(n2254));
NOR3X1   g0420(.A(g876), .B(n2254), .C(n2249), .Y(n2255));
AND2X1   g0421(.A(n2255), .B(n2253), .Y(n2256_1));
OAI21X1  g0422(.A0(n2060), .A1(n2028), .B0(g109), .Y(n2257));
NAND2X1  g0423(.A(g877), .B(g109), .Y(n2258));
NOR2X1   g0424(.A(n2258), .B(n2257), .Y(n2259));
OAI21X1  g0425(.A0(n2192), .A1(n2166_1), .B0(g109), .Y(n2260));
AND2X1   g0426(.A(g757), .B(g109), .Y(n2261_1));
INVX1    g0427(.A(n2261_1), .Y(n2262));
OAI21X1  g0428(.A0(n2111_1), .A1(n2077_1), .B0(g109), .Y(n2263));
NAND2X1  g0429(.A(g881), .B(g109), .Y(n2264));
OAI22X1  g0430(.A0(n2263), .A1(n2264), .B0(n2262), .B1(n2260), .Y(n2265));
NOR4X1   g0431(.A(n2259), .B(n2256_1), .C(n2252), .D(n2265), .Y(g10628));
AOI21X1  g0432(.A0(n1932), .A1(g48), .B0(g32), .Y(n2267));
INVX1    g0433(.A(n1983), .Y(n2268));
XOR2X1   g0434(.A(n2004), .B(n2268), .Y(n2269));
XOR2X1   g0435(.A(n2246_1), .B(n2223), .Y(n2270));
XOR2X1   g0436(.A(n2270), .B(n2269), .Y(n2271_1));
NOR2X1   g0437(.A(n2192), .B(n2166_1), .Y(n2272));
XOR2X1   g0438(.A(n2272), .B(n2251_1), .Y(n2273));
OR2X1    g0439(.A(n2060), .B(n2028), .Y(n2274));
NOR2X1   g0440(.A(n2111_1), .B(n2077_1), .Y(n2275));
XOR2X1   g0441(.A(n2275), .B(n2274), .Y(n2276_1));
XOR2X1   g0442(.A(n2276_1), .B(n2273), .Y(n2277));
XOR2X1   g0443(.A(n2277), .B(n2271_1), .Y(n2278));
XOR2X1   g0444(.A(n2278), .B(n2267), .Y(n2279));
OR2X1    g0445(.A(n2279), .B(n2006), .Y(g10801));
NAND2X1  g0446(.A(g108), .B(g109), .Y(n2283));
NOR2X1   g0447(.A(n2283), .B(n2260), .Y(n2284));
NAND2X1  g0448(.A(g1206), .B(g109), .Y(n2285));
NOR2X1   g0449(.A(n2285), .B(g1361), .Y(n2286_1));
NAND2X1  g0450(.A(n2286_1), .B(n2253), .Y(n2287));
NOR2X1   g0451(.A(n2004), .B(n2249), .Y(n2288));
NAND3X1  g0452(.A(n2288), .B(g865), .C(g109), .Y(n2289));
NAND2X1  g0453(.A(n2289), .B(n2287), .Y(n2290));
AOI21X1  g0454(.A0(n1982_1), .A1(n1958), .B0(n2249), .Y(n2291_1));
AND2X1   g0455(.A(g1610), .B(g1765), .Y(n2292));
AND2X1   g0456(.A(n2292), .B(g109), .Y(n560));
AND2X1   g0457(.A(n560), .B(n2291_1), .Y(n2294));
NOR3X1   g0458(.A(n2246_1), .B(g105), .C(n2249), .Y(n2295));
NOR4X1   g0459(.A(n2294), .B(n2290), .C(n2284), .D(n2295), .Y(n2296_1));
XOR2X1   g0460(.A(n2296_1), .B(n2279), .Y(g11163));
AND2X1   g0461(.A(n2296_1), .B(g10628), .Y(g11206));
ZERO     g0462(.Y(g11489));
INVX1    g0463(.A(g1700), .Y(n1825));
NOR3X1   g0464(.A(g1959), .B(n1825), .C(g1696), .Y(g6842));
INVX1    g0465(.A(g746), .Y(n2302));
NOR2X1   g0466(.A(n2302), .B(g750), .Y(g4171));
INVX1    g0467(.A(g23), .Y(g3327));
OR2X1    g0468(.A(g1212), .B(g1289), .Y(n455));
INVX1    g0469(.A(g1882), .Y(n2306_1));
INVX1    g0470(.A(g1845), .Y(n2307));
NOR4X1   g0471(.A(g1861), .B(g1868), .C(g1864), .D(n2307), .Y(n2308));
INVX1    g0472(.A(g1857), .Y(n2309));
NOR2X1   g0473(.A(g1828), .B(g1822), .Y(n2310));
NOR2X1   g0474(.A(n2310), .B(n2309), .Y(n2311_1));
NAND2X1  g0475(.A(g1834), .B(g1814), .Y(n2312));
NOR2X1   g0476(.A(n2312), .B(g1840), .Y(n2313));
OAI21X1  g0477(.A0(n2313), .A1(n2311_1), .B0(n2308), .Y(n2314));
INVX1    g0478(.A(g1840), .Y(n2315));
INVX1    g0479(.A(g1834), .Y(n2316_1));
NAND4X1  g0480(.A(n2316_1), .B(g1814), .C(n2315), .D(n2310), .Y(n2317));
INVX1    g0481(.A(n2317), .Y(n2318));
OAI21X1  g0482(.A0(n2318), .A1(g1840), .B0(n2308), .Y(n2319));
NAND2X1  g0483(.A(n2319), .B(n2314), .Y(n2320));
INVX1    g0484(.A(g1887), .Y(n2321_1));
INVX1    g0485(.A(g1822), .Y(n2322));
NOR2X1   g0486(.A(n2322), .B(g1814), .Y(n2323));
INVX1    g0487(.A(n2323), .Y(n2324));
OAI21X1  g0488(.A0(g1828), .A1(g1814), .B0(n2322), .Y(n2325));
OAI21X1  g0489(.A0(n2324), .A1(g1828), .B0(n2325), .Y(n2326_1));
XOR2X1   g0490(.A(n2326_1), .B(g1872), .Y(n2327));
MX2X1    g0491(.A(n2321_1), .B(n2327), .S0(n2319), .Y(n2328));
XOR2X1   g0492(.A(n2328), .B(g1882), .Y(n2329));
MX2X1    g0493(.A(n2306_1), .B(n2329), .S0(n2320), .Y(n2330));
NOR4X1   g0494(.A(g1828), .B(g1822), .C(g1814), .D(g1834), .Y(n2331_1));
INVX1    g0495(.A(g1927), .Y(n2332));
INVX1    g0496(.A(g1918), .Y(n2333));
INVX1    g0497(.A(g1909), .Y(n2334));
NOR4X1   g0498(.A(g1891), .B(g1900), .C(g1882), .D(g1872), .Y(n2335));
NAND4X1  g0499(.A(n2334), .B(n2333), .C(n2332), .D(n2335), .Y(n2336_1));
OR4X1    g0500(.A(n2326_1), .B(g1945), .C(g1936), .D(n2336_1), .Y(n2337));
NAND4X1  g0501(.A(g1891), .B(g1900), .C(g1882), .D(g1872), .Y(n2338));
NOR4X1   g0502(.A(n2334), .B(n2333), .C(n2332), .D(n2338), .Y(n2339));
NAND4X1  g0503(.A(n2326_1), .B(g1945), .C(g1936), .D(n2339), .Y(n2340));
AOI21X1  g0504(.A0(n2340), .A1(n2337), .B0(n2314), .Y(n2341_1));
OR2X1    g0505(.A(n2341_1), .B(n2331_1), .Y(n2342));
INVX1    g0506(.A(g1828), .Y(n2343));
NOR3X1   g0507(.A(n2343), .B(g1822), .C(g1814), .Y(n2344));
INVX1    g0508(.A(n2344), .Y(n2345));
INVX1    g0509(.A(n2331_1), .Y(n2346_1));
AOI21X1  g0510(.A0(n2343), .A1(g1822), .B0(n2313), .Y(n2347));
NAND4X1  g0511(.A(n2341_1), .B(n2346_1), .C(n2345), .D(n2347), .Y(n2348));
OAI21X1  g0512(.A0(n2342), .A1(n2330), .B0(n2348), .Y(n460));
AOI21X1  g0513(.A0(n2245), .A1(n2230), .B0(n2249), .Y(n2350));
XOR2X1   g0514(.A(n2350), .B(g849), .Y(n2351_1));
XOR2X1   g0515(.A(n2288), .B(g857), .Y(n2352));
XOR2X1   g0516(.A(n2291_1), .B(g853), .Y(n2353));
XOR2X1   g0517(.A(n2253), .B(g845), .Y(n2354));
AND2X1   g0518(.A(n2257), .B(g829), .Y(n2355));
OAI21X1  g0519(.A0(n2152), .A1(n2124), .B0(g109), .Y(n2356_1));
NOR2X1   g0520(.A(n2356_1), .B(g837), .Y(n2357));
OR4X1    g0521(.A(n2355), .B(n2354), .C(n2353), .D(n2357), .Y(n2358));
INVX1    g0522(.A(g841), .Y(n2359));
NOR4X1   g0523(.A(n2160), .B(n2157), .C(n2024), .D(n2165), .Y(n2360));
NOR4X1   g0524(.A(n2172), .B(n2170), .C(n2168), .D(n2174), .Y(n2362));
NOR2X1   g0525(.A(n1922), .B(n1919_1), .Y(n2364));
AOI22X1  g0526(.A0(n2364), .A1(g940), .B0(g959), .B1(n2211_1), .Y(n2365));
INVX1    g0527(.A(g907), .Y(n2366_1));
NOR3X1   g0528(.A(n1919_1), .B(n1926), .C(n2366_1), .Y(n2367));
INVX1    g0529(.A(g895), .Y(n2368));
NOR4X1   g0530(.A(n1919_1), .B(n1928_1), .C(n2368), .D(n1929), .Y(n2369));
INVX1    g0531(.A(g986), .Y(n2370));
NOR3X1   g0532(.A(n1919_1), .B(n1924_1), .C(n2370), .Y(n2371_1));
NOR3X1   g0533(.A(n2371_1), .B(n2369), .C(n2367), .Y(n2372));
AOI21X1  g0534(.A0(n2372), .A1(n2365), .B0(n1967_1), .Y(n2373));
AND2X1   g0535(.A(n2186_1), .B(n2185), .Y(n2374));
AND2X1   g0536(.A(n2189), .B(n2188), .Y(n2375));
OAI22X1  g0537(.A0(n2374), .A1(n1909_1), .B0(n1903), .B1(n2375), .Y(n2376_1));
NOR3X1   g0538(.A(n2376_1), .B(n2373), .C(n2175), .Y(n2377));
AOI21X1  g0539(.A0(n2377), .A1(n2360), .B0(n2249), .Y(n2378));
AOI22X1  g0540(.A0(n2356_1), .A1(g837), .B0(n2359), .B1(n2378), .Y(n2379));
XOR2X1   g0541(.A(n2257), .B(g861), .Y(n2380));
INVX1    g0542(.A(g829), .Y(n2381_1));
NOR4X1   g0543(.A(n2024), .B(n2020), .C(n2015), .D(n2027_1), .Y(n2382));
AOI22X1  g0544(.A0(n2078), .A1(g1170), .B0(g1336), .B1(n1964), .Y(n2383));
AND2X1   g0545(.A(n2033), .B(n2032_1), .Y(n2384));
AOI21X1  g0546(.A0(n2384), .A1(n2383), .B0(n2080), .Y(n2385));
AOI22X1  g0547(.A0(n2364), .A1(g928), .B0(g950), .B1(n2211_1), .Y(n2386_1));
NOR4X1   g0548(.A(n2046), .B(n2044), .C(n2042_1), .D(n2048), .Y(n2387));
AOI21X1  g0549(.A0(n2387), .A1(n2386_1), .B0(n1967_1), .Y(n2388));
AND2X1   g0550(.A(n2054), .B(n2053), .Y(n2389));
AND2X1   g0551(.A(n2057_1), .B(n2056), .Y(n2390));
OAI22X1  g0552(.A0(n2389), .A1(n1909_1), .B0(n1903), .B1(n2390), .Y(n2391_1));
NOR3X1   g0553(.A(n2391_1), .B(n2388), .C(n2385), .Y(n2392));
AOI21X1  g0554(.A0(n2392), .A1(n2382), .B0(n2249), .Y(n2393));
AOI22X1  g0555(.A0(n2393), .A1(n2381_1), .B0(g833), .B1(n2263), .Y(n2394));
INVX1    g0556(.A(g833), .Y(n2395));
NOR4X1   g0557(.A(n2071), .B(n2068), .C(n2024), .D(n2076), .Y(n2396_1));
NOR4X1   g0558(.A(n2086), .B(n2084), .C(n2082_1), .D(n2088), .Y(n2397));
AOI22X1  g0559(.A0(n2364), .A1(g932), .B0(g953), .B1(n2211_1), .Y(n2399));
NOR4X1   g0560(.A(n2099), .B(n2097), .C(n2095), .D(n2101_1), .Y(n2400));
AOI21X1  g0561(.A0(n2400), .A1(n2399), .B0(n1967_1), .Y(n2401_1));
AND2X1   g0562(.A(n2105), .B(n2104), .Y(n2402));
AND2X1   g0563(.A(n2108), .B(n2107), .Y(n2403));
OAI22X1  g0564(.A0(n2402), .A1(n1909_1), .B0(n1903), .B1(n2403), .Y(n2404));
NOR3X1   g0565(.A(n2404), .B(n2401_1), .C(n2089), .Y(n2405));
AOI21X1  g0566(.A0(n2405), .A1(n2396_1), .B0(n2249), .Y(n2406_1));
AOI22X1  g0567(.A0(n2260), .A1(g841), .B0(n2395), .B1(n2406_1), .Y(n2407));
NAND4X1  g0568(.A(n2394), .B(n2380), .C(n2379), .D(n2407), .Y(n2408));
NOR4X1   g0569(.A(n2358), .B(n2352), .C(n2351_1), .D(n2408), .Y(n2409));
NOR3X1   g0570(.A(g853), .B(g849), .C(g861), .Y(n2410));
NOR4X1   g0571(.A(g841), .B(g857), .C(g837), .D(g845), .Y(n2411_1));
NAND4X1  g0572(.A(n2410), .B(n2395), .C(n2381_1), .D(n2411_1), .Y(n2412));
NOR2X1   g0573(.A(n2412), .B(n2409), .Y(n2413));
AND2X1   g0574(.A(g452), .B(g109), .Y(n2414));
MX2X1    g0575(.A(g421), .B(n2414), .S0(n2413), .Y(n470));
INVX1    g0576(.A(g123), .Y(n2416_1));
NAND2X1  g0577(.A(g115), .B(g18), .Y(n2417));
OR4X1    g0578(.A(g119), .B(g158), .C(g153), .D(g162), .Y(n2418));
OR2X1    g0579(.A(n2418), .B(n2417), .Y(n2419));
INVX1    g0580(.A(g131), .Y(n2420));
NAND3X1  g0581(.A(n2420), .B(g182), .C(g178), .Y(n2421_1));
INVX1    g0582(.A(g174), .Y(n2422));
INVX1    g0583(.A(g170), .Y(n2423));
OR4X1    g0584(.A(n2423), .B(g143), .C(n2422), .D(g127), .Y(n2424));
INVX1    g0585(.A(g166), .Y(n2425));
OR4X1    g0586(.A(g139), .B(g148), .C(n2425), .D(g135), .Y(n2426_1));
OR4X1    g0587(.A(n2424), .B(n2421_1), .C(n2419), .D(n2426_1), .Y(n2427));
AOI21X1  g0588(.A0(n2427), .A1(n2416_1), .B0(n2249), .Y(n475));
AND2X1   g0589(.A(g1380), .B(g109), .Y(n480));
INVX1    g0590(.A(g713), .Y(n2430));
INVX1    g0591(.A(g654), .Y(n2431_1));
NOR3X1   g0592(.A(g643), .B(g650), .C(g646), .Y(n2432));
NAND3X1  g0593(.A(n2432), .B(n2431_1), .C(g627), .Y(n2433));
INVX1    g0594(.A(n2433), .Y(n2434));
INVX1    g0595(.A(g639), .Y(n2435));
INVX1    g0596(.A(g599), .Y(n2436_1));
INVX1    g0597(.A(g605), .Y(n2437));
AOI21X1  g0598(.A0(n2437), .A1(n2436_1), .B0(n2435), .Y(n2438));
INVX1    g0599(.A(g611), .Y(n2439));
INVX1    g0600(.A(g591), .Y(n2440_1));
NOR3X1   g0601(.A(n2440_1), .B(g617), .C(n2439), .Y(n2441));
OAI21X1  g0602(.A0(n2441), .A1(n2438), .B0(n2434), .Y(n2442));
OR2X1    g0603(.A(g605), .B(g611), .Y(n2443));
NOR4X1   g0604(.A(n2440_1), .B(g599), .C(g617), .D(n2443), .Y(n2444));
OAI21X1  g0605(.A0(n2444), .A1(g617), .B0(n2434), .Y(n2445_1));
NAND2X1  g0606(.A(n2445_1), .B(n2442), .Y(n2446));
INVX1    g0607(.A(g718), .Y(n2447));
INVX1    g0608(.A(g695), .Y(n2448));
INVX1    g0609(.A(g704), .Y(n2449));
NOR4X1   g0610(.A(g658), .B(g668), .C(g686), .D(g677), .Y(n2450_1));
NAND3X1  g0611(.A(n2450_1), .B(n2449), .C(n2448), .Y(n2451));
NOR3X1   g0612(.A(g605), .B(g591), .C(n2436_1), .Y(n2452));
AOI21X1  g0613(.A0(n2437), .A1(n2440_1), .B0(g599), .Y(n2453));
NOR2X1   g0614(.A(n2453), .B(n2452), .Y(n2454));
INVX1    g0615(.A(g686), .Y(n2455_1));
NAND3X1  g0616(.A(g677), .B(g658), .C(g668), .Y(n2456));
OR4X1    g0617(.A(n2455_1), .B(n2449), .C(n2448), .D(n2456), .Y(n2457));
MX2X1    g0618(.A(n2457), .B(n2451), .S0(n2454), .Y(n2458));
MX2X1    g0619(.A(n2447), .B(n2458), .S0(n2445_1), .Y(n2459));
XOR2X1   g0620(.A(n2459), .B(g713), .Y(n2460_1));
MX2X1    g0621(.A(n2430), .B(n2460_1), .S0(n2446), .Y(n2461));
NOR4X1   g0622(.A(g591), .B(g599), .C(g611), .D(g605), .Y(n2462));
NAND4X1  g0623(.A(n2449), .B(n2448), .C(n2430), .D(n2450_1), .Y(n2463));
OR2X1    g0624(.A(n2463), .B(g722), .Y(n2464));
OR4X1    g0625(.A(n2453), .B(n2452), .C(g731), .D(n2464), .Y(n2465_1));
INVX1    g0626(.A(g722), .Y(n2466));
INVX1    g0627(.A(g731), .Y(n2467));
NAND4X1  g0628(.A(g658), .B(g668), .C(g686), .D(g677), .Y(n2468));
NOR4X1   g0629(.A(n2449), .B(n2448), .C(n2430), .D(n2468), .Y(n2469));
INVX1    g0630(.A(n2469), .Y(n2470_1));
OR4X1    g0631(.A(n2454), .B(n2467), .C(n2466), .D(n2470_1), .Y(n2471));
AOI21X1  g0632(.A0(n2471), .A1(n2465_1), .B0(n2442), .Y(n2472));
OR2X1    g0633(.A(n2472), .B(n2462), .Y(n2473));
NOR3X1   g0634(.A(n2437), .B(g591), .C(g599), .Y(n2474));
INVX1    g0635(.A(n2472), .Y(n2475_1));
AOI21X1  g0636(.A0(n2437), .A1(g599), .B0(n2441), .Y(n2476));
INVX1    g0637(.A(n2476), .Y(n2477));
OR4X1    g0638(.A(n2475_1), .B(n2462), .C(n2474), .D(n2477), .Y(n2478));
OAI21X1  g0639(.A0(n2473), .A1(n2461), .B0(n2478), .Y(n485));
AND2X1   g0640(.A(g1153), .B(g109), .Y(n490));
OAI21X1  g0641(.A0(g1703), .A1(g1696), .B0(g1209), .Y(n2481));
INVX1    g0642(.A(g1776), .Y(n2482));
INVX1    g0643(.A(n2356_1), .Y(n2483));
INVX1    g0644(.A(g1796), .Y(n2484));
NOR2X1   g0645(.A(g1703), .B(g1696), .Y(n2485_1));
OAI21X1  g0646(.A0(n2291_1), .A1(n2484), .B0(n2485_1), .Y(n2486));
AOI21X1  g0647(.A0(n2483), .A1(n2482), .B0(n2486), .Y(n2487));
XOR2X1   g0648(.A(n2257), .B(g1766), .Y(n2488));
AND2X1   g0649(.A(n2488), .B(n2487), .Y(n2489));
OAI21X1  g0650(.A0(n2004), .A1(n2249), .B0(g1801), .Y(n2490_1));
INVX1    g0651(.A(g1801), .Y(n2491));
INVX1    g0652(.A(n2350), .Y(n2492));
AOI22X1  g0653(.A0(n2288), .A1(n2491), .B0(g1791), .B1(n2492), .Y(n2493));
INVX1    g0654(.A(g1786), .Y(n2494));
AOI22X1  g0655(.A0(n2253), .A1(n2494), .B0(n2484), .B1(n2291_1), .Y(n2495_1));
INVX1    g0656(.A(g1791), .Y(n2496));
NOR2X1   g0657(.A(n2253), .B(n2494), .Y(n2497));
AOI21X1  g0658(.A0(n2350), .A1(n2496), .B0(n2497), .Y(n2498));
AND2X1   g0659(.A(n2498), .B(n2495_1), .Y(n2499));
NAND4X1  g0660(.A(n2493), .B(n2490_1), .C(n2489), .D(n2499), .Y(n2500_1));
NAND2X1  g0661(.A(n2356_1), .B(g1776), .Y(n2501));
XOR2X1   g0662(.A(n2257), .B(g1806), .Y(n2502));
XOR2X1   g0663(.A(n2263), .B(g1771), .Y(n2503));
XOR2X1   g0664(.A(n2260), .B(g1781), .Y(n2504));
NAND4X1  g0665(.A(n2503), .B(n2502), .C(n2501), .D(n2504), .Y(n2505_1));
OAI21X1  g0666(.A0(n2505_1), .A1(n2500_1), .B0(n2481), .Y(n495));
MX2X1    g0667(.A(g1744), .B(g1776), .S0(n2292), .Y(n500));
NOR2X1   g0668(.A(n2417), .B(g12), .Y(n2508));
NOR3X1   g0669(.A(n2508), .B(g1527), .C(n2249), .Y(n2509));
MX2X1    g0670(.A(g1462), .B(g1558), .S0(n2509), .Y(n505));
INVX1    g0671(.A(g700), .Y(n2511));
INVX1    g0672(.A(n2450_1), .Y(n2512));
MX2X1    g0673(.A(n2468), .B(n2512), .S0(n2454), .Y(n2513));
MX2X1    g0674(.A(n2511), .B(n2513), .S0(n2445_1), .Y(n2514));
XOR2X1   g0675(.A(n2514), .B(g695), .Y(n2515_1));
MX2X1    g0676(.A(n2448), .B(n2515_1), .S0(n2446), .Y(n2516));
OAI21X1  g0677(.A0(n2516), .A1(n2473), .B0(n2478), .Y(n510));
AND2X1   g0678(.A(g456), .B(g461), .Y(n2518));
AND2X1   g0679(.A(n2518), .B(g466), .Y(n2519));
AOI21X1  g0680(.A0(n2519), .A1(g471), .B0(n2413), .Y(n2520_1));
XOR2X1   g0681(.A(g456), .B(g461), .Y(n2521));
MX2X1    g0682(.A(g461), .B(n2521), .S0(n2520_1), .Y(n2522));
NOR2X1   g0683(.A(g868), .B(n2249), .Y(n2523));
AND2X1   g0684(.A(n2523), .B(n2522), .Y(n515));
NOR3X1   g0685(.A(n2250), .B(g882), .C(n2249), .Y(n2525_1));
AOI21X1  g0686(.A0(g881), .A1(g109), .B0(n2525_1), .Y(n809));
INVX1    g0687(.A(n809), .Y(n2527));
OAI21X1  g0688(.A0(n2527), .A1(g114), .B0(g109), .Y(n2528));
NOR2X1   g0689(.A(n2528), .B(n2177), .Y(n520));
AND2X1   g0690(.A(g374), .B(g369), .Y(n2530_1));
AND2X1   g0691(.A(n2530_1), .B(g378), .Y(n2531));
AND2X1   g0692(.A(n2531), .B(g382), .Y(n2532));
INVX1    g0693(.A(g305), .Y(n2533));
NOR4X1   g0694(.A(g406), .B(g416), .C(g401), .D(g411), .Y(n2534));
NOR4X1   g0695(.A(g386), .B(g426), .C(g396), .D(g391), .Y(n2535_1));
NOR3X1   g0696(.A(g431), .B(g440), .C(g444), .Y(n2536));
NOR4X1   g0697(.A(g421), .B(g448), .C(g452), .D(g435), .Y(n2537));
NAND4X1  g0698(.A(n2536), .B(n2535_1), .C(n2534), .D(n2537), .Y(n2538));
INVX1    g0699(.A(g431), .Y(n2539));
XOR2X1   g0700(.A(g435), .B(n2539), .Y(n2540_1));
NAND2X1  g0701(.A(n2540_1), .B(n2538), .Y(n2541));
MX2X1    g0702(.A(g305), .B(n2541), .S0(n2532), .Y(n2542));
AND2X1   g0703(.A(n2542), .B(n2533), .Y(n2543));
NAND4X1  g0704(.A(n2538), .B(n2532), .C(g305), .D(n2540_1), .Y(n2544));
XOR2X1   g0705(.A(g426), .B(g315), .Y(n2545_1));
XOR2X1   g0706(.A(g324), .B(g396), .Y(n2546));
XOR2X1   g0707(.A(g401), .B(g327), .Y(n2547));
NOR3X1   g0708(.A(n2547), .B(n2546), .C(n2545_1), .Y(n2548));
XOR2X1   g0709(.A(g411), .B(g333), .Y(n2549));
XOR2X1   g0710(.A(g406), .B(g330), .Y(n2550_1));
XOR2X1   g0711(.A(g416), .B(g309), .Y(n2551));
XOR2X1   g0712(.A(g421), .B(g312), .Y(n2552));
XOR2X1   g0713(.A(g321), .B(g391), .Y(n2553));
XOR2X1   g0714(.A(g318), .B(g386), .Y(n2554));
OR4X1    g0715(.A(n2553), .B(n2552), .C(n2551), .D(n2554), .Y(n2555_1));
NOR3X1   g0716(.A(n2555_1), .B(n2550_1), .C(n2549), .Y(n2556));
NAND3X1  g0717(.A(n2556), .B(n2548), .C(n2544), .Y(n2557));
OAI21X1  g0718(.A0(n2557), .A1(n2543), .B0(n2532), .Y(n2558));
NOR2X1   g0719(.A(n2558), .B(n2413), .Y(n639));
XOR2X1   g0720(.A(g971), .B(n2096_1), .Y(n2560_1));
MX2X1    g0721(.A(n2096_1), .B(n2560_1), .S0(n639), .Y(n2561));
NOR2X1   g0722(.A(n2261_1), .B(n2255), .Y(n2562));
NAND2X1  g0723(.A(n2562), .B(g869), .Y(n2563));
NAND2X1  g0724(.A(n2563), .B(g109), .Y(n2564));
NOR2X1   g0725(.A(n2564), .B(n2561), .Y(n525));
NAND4X1  g0726(.A(g617), .B(n2431_1), .C(g627), .D(n2432), .Y(n2566));
NOR2X1   g0727(.A(n2566), .B(g611), .Y(n2567));
INVX1    g0728(.A(g709), .Y(n2568));
NOR2X1   g0729(.A(n2462), .B(n2568), .Y(n2569));
MX2X1    g0730(.A(n2569), .B(g700), .S0(n2567), .Y(n530));
INVX1    g0731(.A(g1703), .Y(n2571));
NOR2X1   g0732(.A(n2571), .B(g1696), .Y(n2572));
MX2X1    g0733(.A(g1092), .B(g360), .S0(n2572), .Y(n535));
NOR3X1   g0734(.A(n2508), .B(g1570), .C(n2249), .Y(n2574));
MX2X1    g0735(.A(g1515), .B(g1574), .S0(n2574), .Y(n540));
INVX1    g0736(.A(g1864), .Y(n2576));
XOR2X1   g0737(.A(g1861), .B(g1864), .Y(n2577));
MX2X1    g0738(.A(n2576), .B(n2577), .S0(g1845), .Y(n2578));
NOR3X1   g0739(.A(n2578), .B(n2331_1), .C(n2308), .Y(n545));
NOR2X1   g0740(.A(n2532), .B(n2413), .Y(n2580_1));
XOR2X1   g0741(.A(n2580_1), .B(g369), .Y(n2581));
NOR2X1   g0742(.A(g869), .B(n2249), .Y(n2582));
AND2X1   g0743(.A(n2582), .B(n2581), .Y(n550));
MX2X1    g0744(.A(g1411), .B(g1580), .S0(n2574), .Y(n555));
OR2X1    g0745(.A(n1983), .B(n1892), .Y(n2585_1));
OAI21X1  g0746(.A0(n1984), .A1(n2006), .B0(n2585_1), .Y(n565));
INVX1    g0747(.A(g1651), .Y(n2587));
AOI21X1  g0748(.A0(n2571), .A1(g1696), .B0(n2587), .Y(n570));
AND2X1   g0749(.A(g1407), .B(g109), .Y(n575));
INVX1    g0750(.A(g1718), .Y(n2590_1));
NAND2X1  g0751(.A(g1357), .B(n2590_1), .Y(n2591));
NOR2X1   g0752(.A(g1357), .B(g1718), .Y(n2592));
MX2X1    g0753(.A(g1618), .B(g186), .S0(g18), .Y(n2593));
NAND2X1  g0754(.A(n2593), .B(n2592), .Y(n2594));
OAI21X1  g0755(.A0(n2591), .A1(n2257), .B0(n2594), .Y(n2595_1));
MX2X1    g0756(.A(g1672), .B(n2595_1), .S0(n2485_1), .Y(n584));
MX2X1    g0757(.A(g1077), .B(g345), .S0(n2572), .Y(n589));
AND2X1   g0758(.A(g1223), .B(g1218), .Y(n2598));
AND2X1   g0759(.A(n2598), .B(g1227), .Y(n2599));
INVX1    g0760(.A(g1713), .Y(n2600_1));
NAND3X1  g0761(.A(n2485_1), .B(n2600_1), .C(g1289), .Y(n2601));
INVX1    g0762(.A(n2601), .Y(n2602));
AOI21X1  g0763(.A0(n2602), .A1(n2599), .B0(g1231), .Y(n2603));
NOR3X1   g0764(.A(n2603), .B(g1212), .C(n2249), .Y(n594));
INVX1    g0765(.A(g4), .Y(n2605_1));
NAND4X1  g0766(.A(g1490), .B(g1508), .C(g1504), .D(g1494), .Y(n2606));
NOR3X1   g0767(.A(n2606), .B(g1482), .C(g1499), .Y(n2607));
INVX1    g0768(.A(g1453), .Y(n2608));
NOR4X1   g0769(.A(g1458), .B(g1466), .C(g1486), .D(n2608), .Y(n2609));
INVX1    g0770(.A(g1470), .Y(n2610_1));
INVX1    g0771(.A(g1474), .Y(n2611));
INVX1    g0772(.A(g1478), .Y(n2612));
INVX1    g0773(.A(g1462), .Y(n2613));
NOR4X1   g0774(.A(n2612), .B(n2611), .C(n2610_1), .D(n2613), .Y(n2614));
NAND4X1  g0775(.A(n2609), .B(n2607), .C(n2508), .D(n2614), .Y(n2615_1));
AOI21X1  g0776(.A0(n2615_1), .A1(n2605_1), .B0(n2249), .Y(n599));
NAND4X1  g0777(.A(g770), .B(g766), .C(g758), .D(g762), .Y(n2617));
XOR2X1   g0778(.A(n2617), .B(g774), .Y(n2618));
NOR3X1   g0779(.A(n2618), .B(g590), .C(n2249), .Y(n604));
INVX1    g0780(.A(g1104), .Y(n2620_1));
NOR3X1   g0781(.A(g1216), .B(n2620_1), .C(n2249), .Y(n609));
AND2X1   g0782(.A(g1304), .B(g109), .Y(n2622));
MX2X1    g0783(.A(g1270), .B(n2622), .S0(n2601), .Y(n614));
AND2X1   g0784(.A(g1400), .B(g109), .Y(n619));
INVX1    g0785(.A(g1494), .Y(n2625));
XOR2X1   g0786(.A(n2593), .B(n2625), .Y(n2626));
NOR2X1   g0787(.A(n2626), .B(n2249), .Y(n624));
MX2X1    g0788(.A(g96), .B(g1044), .S0(g85), .Y(n629));
INVX1    g0789(.A(g1448), .Y(n2629_1));
INVX1    g0790(.A(g18), .Y(n2630));
INVX1    g0791(.A(g1101), .Y(n2631));
INVX1    g0792(.A(g1110), .Y(n2632));
NOR4X1   g0793(.A(n2632), .B(n2631), .C(g1104), .D(g1107), .Y(n2633));
XOR2X1   g0794(.A(n2633), .B(g1145), .Y(n2634_1));
MX2X1    g0795(.A(g237), .B(n2634_1), .S0(n2630), .Y(n2635));
XOR2X1   g0796(.A(n2635), .B(n2629_1), .Y(n2636));
NOR2X1   g0797(.A(n2636), .B(n2249), .Y(n634));
INVX1    g0798(.A(g786), .Y(n2638));
INVX1    g0799(.A(g774), .Y(n2639_1));
INVX1    g0800(.A(g778), .Y(n2640));
INVX1    g0801(.A(g782), .Y(n2641));
NOR4X1   g0802(.A(n2641), .B(n2640), .C(n2639_1), .D(n2617), .Y(n2642));
XOR2X1   g0803(.A(n2642), .B(n2638), .Y(n2643));
NOR3X1   g0804(.A(n2643), .B(g590), .C(n2249), .Y(n644));
MX2X1    g0805(.A(g1482), .B(g1543), .S0(n2509), .Y(n649));
INVX1    g0806(.A(g1357), .Y(n2646));
OAI21X1  g0807(.A0(n2356_1), .A1(n2646), .B0(n2590_1), .Y(n2647));
MX2X1    g0808(.A(g552), .B(n2647), .S0(n2485_1), .Y(n654));
MX2X1    g0809(.A(g1494), .B(g1534), .S0(n2509), .Y(n664));
INVX1    g0810(.A(g622), .Y(n2650));
AND2X1   g0811(.A(n2472), .B(n2441), .Y(n2651));
XOR2X1   g0812(.A(n2651), .B(n2650), .Y(n2652));
NOR2X1   g0813(.A(n2652), .B(n2462), .Y(n669));
INVX1    g0814(.A(g1932), .Y(n2654));
NAND3X1  g0815(.A(n2335), .B(n2334), .C(n2333), .Y(n2655));
INVX1    g0816(.A(g1900), .Y(n2656));
NAND3X1  g0817(.A(g1872), .B(g1891), .C(g1882), .Y(n2657));
OR4X1    g0818(.A(n2334), .B(n2656), .C(n2333), .D(n2657), .Y(n2658_1));
MX2X1    g0819(.A(n2655), .B(n2658_1), .S0(n2326_1), .Y(n2659));
MX2X1    g0820(.A(n2654), .B(n2659), .S0(n2319), .Y(n2660));
XOR2X1   g0821(.A(n2660), .B(g1927), .Y(n2661));
MX2X1    g0822(.A(n2332), .B(n2661), .S0(n2320), .Y(n2662));
OAI21X1  g0823(.A0(n2662), .A1(n2342), .B0(n2348), .Y(n674));
INVX1    g0824(.A(n2592), .Y(n2664));
NAND4X1  g0825(.A(n2382), .B(n2590_1), .C(g109), .D(n2392), .Y(n2665));
MX2X1    g0826(.A(g1636), .B(g248), .S0(g18), .Y(n2666));
MX2X1    g0827(.A(n2666), .B(n2665), .S0(n2664), .Y(n2667));
MX2X1    g0828(.A(g1660), .B(n2667), .S0(n2572), .Y(n679));
NOR2X1   g0829(.A(n2417), .B(g119), .Y(n2669));
NOR3X1   g0830(.A(n2669), .B(g126), .C(n2249), .Y(n2670));
MX2X1    g0831(.A(g162), .B(g278), .S0(n2670), .Y(n684));
INVX1    g0832(.A(g1107), .Y(n2672));
NOR4X1   g0833(.A(g1110), .B(n2631), .C(n2620_1), .D(n2672), .Y(n2673_1));
XOR2X1   g0834(.A(n2673_1), .B(g1137), .Y(n2674));
MX2X1    g0835(.A(g225), .B(n2674), .S0(n2630), .Y(n2675));
XOR2X1   g0836(.A(n2675), .B(g1440), .Y(n2676));
AND2X1   g0837(.A(n2676), .B(g109), .Y(n689));
NOR2X1   g0838(.A(n2462), .B(n2447), .Y(n2678_1));
MX2X1    g0839(.A(n2678_1), .B(g709), .S0(n2567), .Y(n694));
INVX1    g0840(.A(g750), .Y(n2680));
NOR2X1   g0841(.A(g754), .B(n2680), .Y(n2681));
INVX1    g0842(.A(n2681), .Y(n2682));
AND2X1   g0843(.A(n2682), .B(g76), .Y(n699));
NAND4X1  g0844(.A(n2396_1), .B(n2590_1), .C(g109), .D(n2405), .Y(n2684));
MX2X1    g0845(.A(g1639), .B(g207), .S0(g18), .Y(n2685));
MX2X1    g0846(.A(n2685), .B(n2684), .S0(n2664), .Y(n2686));
MX2X1    g0847(.A(g554), .B(n2686), .S0(n2485_1), .Y(n704));
AND2X1   g0848(.A(g496), .B(g109), .Y(n2688_1));
MX2X1    g0849(.A(g491), .B(n2688_1), .S0(n2413), .Y(n709));
INVX1    g0850(.A(g981), .Y(n2690));
AND2X1   g0851(.A(g971), .B(g976), .Y(n2691));
XOR2X1   g0852(.A(n2691), .B(n2690), .Y(n2692));
MX2X1    g0853(.A(n2690), .B(n2692), .S0(n639), .Y(n2693_1));
NOR2X1   g0854(.A(n2693_1), .B(n2564), .Y(n714));
NAND3X1  g0855(.A(g971), .B(g981), .C(g976), .Y(n2695));
NOR2X1   g0856(.A(n2695), .B(n2370), .Y(n719));
MX2X1    g0857(.A(g1095), .B(g363), .S0(n2572), .Y(n734));
NAND2X1  g0858(.A(n2450_1), .B(n2448), .Y(n2698_1));
OR2X1    g0859(.A(n2468), .B(n2448), .Y(n2699));
MX2X1    g0860(.A(n2699), .B(n2698_1), .S0(n2454), .Y(n2700));
MX2X1    g0861(.A(n2568), .B(n2700), .S0(n2445_1), .Y(n2701));
XOR2X1   g0862(.A(n2701), .B(g704), .Y(n2702));
MX2X1    g0863(.A(n2449), .B(n2702), .S0(n2446), .Y(n2703_1));
OAI21X1  g0864(.A0(n2703_1), .A1(n2473), .B0(n2478), .Y(n739));
AND2X1   g0865(.A(g1265), .B(g109), .Y(n2705));
MX2X1    g0866(.A(g1260), .B(n2705), .S0(n2601), .Y(n744));
INVX1    g0867(.A(g1696), .Y(n2707));
NOR2X1   g0868(.A(g1703), .B(n2707), .Y(n2708_1));
NAND4X1  g0869(.A(g1781), .B(g1771), .C(g1766), .D(g1776), .Y(n2709));
XOR2X1   g0870(.A(n2709), .B(g1786), .Y(n2710));
MX2X1    g0871(.A(n2494), .B(n2710), .S0(n2708_1), .Y(n2711));
NOR2X1   g0872(.A(n2711), .B(g1713), .Y(n749));
INVX1    g0873(.A(g682), .Y(n2713_1));
NOR2X1   g0874(.A(n2462), .B(n2713_1), .Y(n2714));
MX2X1    g0875(.A(n2714), .B(g673), .S0(n2567), .Y(n754));
AND2X1   g0876(.A(g1296), .B(g109), .Y(n2716));
MX2X1    g0877(.A(g1300), .B(n2716), .S0(n2601), .Y(n759));
AND2X1   g0878(.A(n2682), .B(g52), .Y(n769));
INVX1    g0879(.A(g646), .Y(n2719));
XOR2X1   g0880(.A(g643), .B(g646), .Y(n2720));
MX2X1    g0881(.A(n2719), .B(n2720), .S0(g627), .Y(n2721));
NOR3X1   g0882(.A(n2721), .B(n2462), .C(n2434), .Y(n774));
AND2X1   g0883(.A(g197), .B(g109), .Y(n784));
AND2X1   g0884(.A(g225), .B(g109), .Y(n789));
MX2X1    g0885(.A(g1675), .B(n2686), .S0(n2485_1), .Y(n799));
OAI21X1  g0886(.A0(g754), .A1(n2680), .B0(g354), .Y(n2726));
INVX1    g0887(.A(g321), .Y(n2727));
INVX1    g0888(.A(g466), .Y(n2728_1));
NOR4X1   g0889(.A(n2728_1), .B(g471), .C(g461), .D(g456), .Y(n2729));
XOR2X1   g0890(.A(n2729), .B(g491), .Y(n2730));
INVX1    g0891(.A(n2730), .Y(n2731));
MX2X1    g0892(.A(n2731), .B(n2727), .S0(n2413), .Y(n2732));
OAI21X1  g0893(.A0(n2732), .A1(n2682), .B0(n2726), .Y(n804));
INVX1    g0894(.A(n2462), .Y(n2734));
OAI21X1  g0895(.A0(n2437), .A1(n2440_1), .B0(n2436_1), .Y(n2735));
OR2X1    g0896(.A(n2735), .B(n2474), .Y(n2736));
NAND3X1  g0897(.A(n2736), .B(n2434), .C(n2435), .Y(n2737));
NAND2X1  g0898(.A(n2433), .B(g639), .Y(n2738_1));
NAND3X1  g0899(.A(n2738_1), .B(n2737), .C(n2734), .Y(n814));
NOR2X1   g0900(.A(n2223), .B(n2249), .Y(n2740));
MX2X1    g0901(.A(g1624), .B(g225), .S0(g18), .Y(n2741));
NAND2X1  g0902(.A(n2741), .B(n2592), .Y(n2742));
OAI21X1  g0903(.A0(n2740), .A1(n2591), .B0(n2742), .Y(n2743_1));
MX2X1    g0904(.A(g1684), .B(n2743_1), .S0(n2485_1), .Y(n819));
NOR4X1   g0905(.A(g1110), .B(g1101), .C(n2620_1), .D(g1107), .Y(n2745));
XOR2X1   g0906(.A(n2745), .B(g1117), .Y(n2746));
MX2X1    g0907(.A(g1639), .B(n2746), .S0(n2485_1), .Y(n824));
NOR2X1   g0908(.A(n2709), .B(n2494), .Y(n2748_1));
XOR2X1   g0909(.A(n2748_1), .B(n2496), .Y(n2749));
MX2X1    g0910(.A(n2496), .B(n2749), .S0(n2708_1), .Y(n2750));
NOR2X1   g0911(.A(n2750), .B(g1713), .Y(n829));
AND2X1   g0912(.A(g1397), .B(g109), .Y(n834));
NOR2X1   g0913(.A(g1707), .B(n1825), .Y(n839));
MX2X1    g0914(.A(g1759), .B(g1801), .S0(n2292), .Y(n844));
INVX1    g0915(.A(g461), .Y(n2755));
INVX1    g0916(.A(g456), .Y(n2756));
NOR4X1   g0917(.A(g466), .B(g471), .C(n2755), .D(n2756), .Y(n2757_1));
XOR2X1   g0918(.A(n2757_1), .B(g486), .Y(n2758));
MX2X1    g0919(.A(n2758), .B(g318), .S0(n2413), .Y(n2759));
MX2X1    g0920(.A(g351), .B(n2759), .S0(n2681), .Y(n849));
MX2X1    g0921(.A(g1444), .B(g1604), .S0(n2574), .Y(n857));
MX2X1    g0922(.A(g1098), .B(g366), .S0(n2572), .Y(n862));
NOR2X1   g0923(.A(n2528), .B(n2091_1), .Y(n867));
ZERO     g0924(.Y(n872));
INVX1    g0925(.A(n2308), .Y(n2765));
NOR3X1   g0926(.A(n2765), .B(g1834), .C(n2315), .Y(n2766));
INVX1    g0927(.A(g1896), .Y(n2767_1));
NOR2X1   g0928(.A(n2331_1), .B(n2767_1), .Y(n2768));
MX2X1    g0929(.A(n2768), .B(g1887), .S0(n2766), .Y(n877));
INVX1    g0930(.A(g736), .Y(n2770));
NOR2X1   g0931(.A(n2462), .B(n2770), .Y(n2771));
MX2X1    g0932(.A(n2771), .B(g727), .S0(n2567), .Y(n882));
MX2X1    g0933(.A(g1065), .B(g1098), .S0(n2485_1), .Y(n2773));
MX2X1    g0934(.A(g1019), .B(n2773), .S0(n2485_1), .Y(n887));
AND2X1   g0935(.A(g243), .B(g109), .Y(n892));
AND2X1   g0936(.A(g1411), .B(g109), .Y(n902));
AND2X1   g0937(.A(n2682), .B(g58), .Y(n907));
NAND2X1  g0938(.A(n2279), .B(n2006), .Y(n2778));
NAND2X1  g0939(.A(n2279), .B(n1892), .Y(n2779));
NAND2X1  g0940(.A(n2779), .B(n2778), .Y(n912));
MX2X1    g0941(.A(g1086), .B(g354), .S0(n2572), .Y(n921));
MX2X1    g0942(.A(g1621), .B(g219), .S0(g18), .Y(n2782_1));
XOR2X1   g0943(.A(n2782_1), .B(g1482), .Y(n2783));
AND2X1   g0944(.A(n2783), .B(g109), .Y(n926));
AND2X1   g0945(.A(g1703), .B(g1696), .Y(n2785));
MX2X1    g0946(.A(g1730), .B(n2378), .S0(n2785), .Y(n931));
AND2X1   g0947(.A(g1499), .B(g109), .Y(n936));
MX2X1    g0948(.A(g1633), .B(g243), .S0(g18), .Y(n2788));
XOR2X1   g0949(.A(n2788), .B(g1466), .Y(n2789));
AND2X1   g0950(.A(n2789), .B(g109), .Y(n941));
INVX1    g0951(.A(g745), .Y(n2791));
INVX1    g0952(.A(g822), .Y(n2792_1));
INVX1    g0953(.A(g814), .Y(n2793));
INVX1    g0954(.A(g818), .Y(n2794));
INVX1    g0955(.A(g810), .Y(n2795));
NAND4X1  g0956(.A(g802), .B(g794), .C(g806), .D(g798), .Y(n2796));
NOR4X1   g0957(.A(n2795), .B(n2794), .C(n2793), .D(n2796), .Y(n2797_1));
XOR2X1   g0958(.A(n2797_1), .B(n2792_1), .Y(n2798));
NOR4X1   g0959(.A(n2302), .B(n2791), .C(n2249), .D(n2798), .Y(n946));
OAI21X1  g0960(.A0(g1703), .A1(g1696), .B0(g1678), .Y(n2800));
NOR3X1   g0961(.A(n2356_1), .B(n2646), .C(g1718), .Y(n2801));
MX2X1    g0962(.A(g1615), .B(g213), .S0(g18), .Y(n2802_1));
AND2X1   g0963(.A(n2802_1), .B(n2592), .Y(n2803));
OAI21X1  g0964(.A0(n2803), .A1(n2801), .B0(n2485_1), .Y(n2804));
NAND2X1  g0965(.A(n2804), .B(n2800), .Y(n956));
MX2X1    g0966(.A(g563), .B(g225), .S0(g18), .Y(n1416));
XOR2X1   g0967(.A(n1416), .B(n2423), .Y(n2807_1));
NOR2X1   g0968(.A(n2807_1), .B(n2249), .Y(n961));
XOR2X1   g0969(.A(n2708_1), .B(g1766), .Y(n2809));
OR2X1    g0970(.A(n2809), .B(g1713), .Y(n966));
NOR4X1   g0971(.A(n2484), .B(n2496), .C(n2494), .D(n2709), .Y(n2811));
XOR2X1   g0972(.A(n2811), .B(n2491), .Y(n2812_1));
MX2X1    g0973(.A(n2491), .B(n2812_1), .S0(n2708_1), .Y(n2813));
NOR2X1   g0974(.A(n2813), .B(g1713), .Y(n971));
AND2X1   g0975(.A(g1383), .B(g109), .Y(n976));
NOR4X1   g0976(.A(n2413), .B(n2261_1), .C(n2255), .D(n2558), .Y(n2816));
MX2X1    g0977(.A(g959), .B(g849), .S0(n2816), .Y(n981));
OR2X1    g0978(.A(n2485_1), .B(g1169), .Y(n986));
MX2X1    g0979(.A(g1062), .B(g1095), .S0(n2485_1), .Y(n2819));
MX2X1    g0980(.A(g1007), .B(n2819), .S0(n2485_1), .Y(n991));
INVX1    g0981(.A(g1428), .Y(n2821));
NOR4X1   g0982(.A(g1110), .B(n2631), .C(n2620_1), .D(g1107), .Y(n2822_1));
XOR2X1   g0983(.A(n2822_1), .B(g1121), .Y(n2823));
MX2X1    g0984(.A(g186), .B(n2823), .S0(n2630), .Y(n2824));
XOR2X1   g0985(.A(n2824), .B(n2821), .Y(n2825));
NOR2X1   g0986(.A(n2825), .B(n2249), .Y(n996));
MX2X1    g0987(.A(g91), .B(g1059), .S0(g85), .Y(n1001));
OR2X1    g0988(.A(n2331_1), .B(n2308), .Y(n2828));
NOR2X1   g0989(.A(g1861), .B(g1864), .Y(n2829));
XOR2X1   g0990(.A(n2829), .B(g1868), .Y(n2830));
MX2X1    g0991(.A(g1868), .B(n2830), .S0(g1845), .Y(n2831));
OR2X1    g0992(.A(n2831), .B(n2828), .Y(n1006));
NOR3X1   g0993(.A(g758), .B(g590), .C(n2249), .Y(n1011));
MX2X1    g0994(.A(g1718), .B(g1713), .S0(n2485_1), .Y(n1016));
AND2X1   g0995(.A(g396), .B(g109), .Y(n2835));
MX2X1    g0996(.A(g391), .B(n2835), .S0(n2413), .Y(n1021));
MX2X1    g0997(.A(g1038), .B(g1074), .S0(n2485_1), .Y(n2837_1));
MX2X1    g0998(.A(g1015), .B(n2837_1), .S0(n2485_1), .Y(n1026));
OR2X1    g0999(.A(n2246_1), .B(n1892), .Y(n2839));
OAI21X1  g1000(.A0(n2247), .A1(n2006), .B0(n2839), .Y(n1031));
AOI21X1  g1001(.A0(n2440_1), .A1(g611), .B0(n2462), .Y(n2841));
AND2X1   g1002(.A(n2841), .B(g631), .Y(n1036));
AND2X1   g1003(.A(g1520), .B(g109), .Y(n1041));
NOR2X1   g1004(.A(g1212), .B(n2249), .Y(n2844));
NAND4X1  g1005(.A(g1218), .B(g1227), .C(g1231), .D(g1223), .Y(n2845));
NAND4X1  g1006(.A(n2485_1), .B(n2600_1), .C(g1289), .D(n2845), .Y(n2846));
XOR2X1   g1007(.A(n2598), .B(g1227), .Y(n2847_1));
MX2X1    g1008(.A(n2847_1), .B(g1227), .S0(n2846), .Y(n2848));
AND2X1   g1009(.A(n2848), .B(n2844), .Y(n1046));
MX2X1    g1010(.A(g1721), .B(n2393), .S0(n2785), .Y(n1051));
INVX1    g1011(.A(g1814), .Y(n2851));
AOI21X1  g1012(.A0(g1834), .A1(n2851), .B0(n2331_1), .Y(n2852_1));
INVX1    g1013(.A(n2852_1), .Y(n1061));
MX2X1    g1014(.A(g170), .B(g284), .S0(n2670), .Y(n1066));
AND2X1   g1015(.A(g426), .B(g109), .Y(n2855));
MX2X1    g1016(.A(n2542), .B(n2855), .S0(n2413), .Y(n1071));
AND2X1   g1017(.A(g1371), .B(g109), .Y(n1076));
NAND3X1  g1018(.A(g798), .B(g802), .C(g794), .Y(n2858));
XOR2X1   g1019(.A(n2858), .B(g806), .Y(n2859));
NOR4X1   g1020(.A(n2302), .B(n2791), .C(n2249), .D(n2859), .Y(n1086));
NOR4X1   g1021(.A(g1110), .B(g1101), .C(g1104), .D(n2672), .Y(n2861));
XOR2X1   g1022(.A(n2861), .B(g1125), .Y(n2862_1));
MX2X1    g1023(.A(g207), .B(n2862_1), .S0(n2630), .Y(n2863));
XOR2X1   g1024(.A(n2863), .B(g1403), .Y(n2864));
AND2X1   g1025(.A(n2864), .B(g109), .Y(n1091));
MX2X1    g1026(.A(g1453), .B(g1564), .S0(n2509), .Y(n1101));
MX2X1    g1027(.A(g1741), .B(g1771), .S0(n2292), .Y(n1106));
AND2X1   g1028(.A(g1368), .B(g109), .Y(n1111));
MX2X1    g1029(.A(g174), .B(g281), .S0(n2670), .Y(n1116));
NOR3X1   g1030(.A(g44), .B(g45), .C(g43), .Y(n2870));
NAND4X1  g1031(.A(n1884), .B(n1887), .C(g42), .D(n2870), .Y(n2871));
OR2X1    g1032(.A(n2871), .B(n1910), .Y(n2872_1));
AND2X1   g1033(.A(n2872_1), .B(n2268), .Y(n2873));
OAI21X1  g1034(.A0(n1983), .A1(n2249), .B0(n2872_1), .Y(n2874));
OR2X1    g1035(.A(n2874), .B(n2873), .Y(n2875));
INVX1    g1036(.A(g1027), .Y(n2876));
XOR2X1   g1037(.A(n2876), .B(g1032), .Y(n2877_1));
INVX1    g1038(.A(n2877_1), .Y(n2878));
MX2X1    g1039(.A(g1027), .B(n2878), .S0(n2875), .Y(n2879));
INVX1    g1040(.A(n2879), .Y(n2880));
NOR4X1   g1041(.A(g1255), .B(g1250), .C(g1265), .D(g1260), .Y(n2881));
NOR4X1   g1042(.A(g1275), .B(g1245), .C(g1240), .D(g1235), .Y(n2882_1));
NOR3X1   g1043(.A(g1280), .B(g1292), .C(g1296), .Y(n2883));
NOR4X1   g1044(.A(g1284), .B(g1270), .C(g1304), .D(g1300), .Y(n2884));
NAND4X1  g1045(.A(n2883), .B(n2882_1), .C(n2881), .D(n2884), .Y(n2885));
INVX1    g1046(.A(g1280), .Y(n2886));
XOR2X1   g1047(.A(g1284), .B(n2886), .Y(n2887_1));
NAND2X1  g1048(.A(n2887_1), .B(n2885), .Y(n2888));
MX2X1    g1049(.A(n2888), .B(n2879), .S0(n2845), .Y(n2889));
AND2X1   g1050(.A(n2889), .B(n2880), .Y(n2890));
NOR2X1   g1051(.A(n2889), .B(n2880), .Y(n2891));
XOR2X1   g1052(.A(g995), .B(g1275), .Y(n2892_1));
XOR2X1   g1053(.A(g999), .B(g1245), .Y(n2893));
XOR2X1   g1054(.A(g1250), .B(g1011), .Y(n2894));
NOR3X1   g1055(.A(n2894), .B(n2893), .C(n2892_1), .Y(n2895));
XOR2X1   g1056(.A(g1260), .B(g1019), .Y(n2896));
XOR2X1   g1057(.A(g1255), .B(g1007), .Y(n2897_1));
NOR2X1   g1058(.A(n2897_1), .B(n2896), .Y(n2898));
XOR2X1   g1059(.A(g1015), .B(g1265), .Y(n2899));
XOR2X1   g1060(.A(g1270), .B(g1023), .Y(n2900));
XOR2X1   g1061(.A(g1003), .B(g1240), .Y(n2901));
XOR2X1   g1062(.A(g1235), .B(g991), .Y(n2902_1));
NOR4X1   g1063(.A(n2901), .B(n2900), .C(n2899), .D(n2902_1), .Y(n2903));
NAND3X1  g1064(.A(n2903), .B(n2898), .C(n2895), .Y(n2904));
NOR3X1   g1065(.A(n2904), .B(n2891), .C(n2890), .Y(n2905));
NAND2X1  g1066(.A(n2485_1), .B(g1317), .Y(n2906));
OR4X1    g1067(.A(n2905), .B(n2601), .C(n2845), .D(n2906), .Y(n2907_1));
MX2X1    g1068(.A(g1766), .B(g1308), .S0(n2907_1), .Y(n1121));
INVX1    g1069(.A(n2441), .Y(n2909));
AOI21X1  g1070(.A0(n2472), .A1(g622), .B0(n2909), .Y(n2910));
OAI21X1  g1071(.A0(n2910), .A1(g617), .B0(n2434), .Y(n2911));
XOR2X1   g1072(.A(n2911), .B(g611), .Y(n2912_1));
NOR2X1   g1073(.A(n2912_1), .B(n2630), .Y(n1126));
AND2X1   g1074(.A(n2841), .B(g630), .Y(n1131));
OR2X1    g1075(.A(n2871), .B(n1962_1), .Y(n1136));
MX2X1    g1076(.A(g1428), .B(g1589), .S0(n2574), .Y(n1141));
XOR2X1   g1077(.A(n2666), .B(n2613), .Y(n2917_1));
NOR2X1   g1078(.A(n2917_1), .B(n2249), .Y(n1146));
MX2X1    g1079(.A(g1520), .B(g1571), .S0(n2574), .Y(n1151));
XOR2X1   g1080(.A(n2307), .B(g1861), .Y(n2920));
NOR3X1   g1081(.A(n2920), .B(n2331_1), .C(n2308), .Y(n1156));
AND2X1   g1082(.A(g237), .B(g109), .Y(n1161));
INVX1    g1083(.A(g201), .Y(n2923));
INVX1    g1084(.A(g1811), .Y(n2924));
NAND3X1  g1085(.A(n2872_1), .B(n2492), .C(n2246_1), .Y(n2925));
OR4X1    g1086(.A(g1645), .B(g1642), .C(g1651), .D(g1648), .Y(n2926));
AOI21X1  g1087(.A0(n2926), .A1(n2925), .B0(n2924), .Y(n2927_1));
NAND2X1  g1088(.A(n2926), .B(n2924), .Y(n2928));
AOI21X1  g1089(.A0(n2926), .A1(n2925), .B0(n2928), .Y(n2929));
OR2X1    g1090(.A(n2929), .B(g18), .Y(n2930));
OAI22X1  g1091(.A0(n2927_1), .A1(n2930), .B0(n2923), .B1(n2630), .Y(n2931));
XOR2X1   g1092(.A(g1515), .B(g1415), .Y(n2932_1));
XOR2X1   g1093(.A(n2932_1), .B(g1419), .Y(n2933));
XOR2X1   g1094(.A(n2933), .B(n2629_1), .Y(n2934));
XOR2X1   g1095(.A(n2934), .B(n2931), .Y(n2935));
NOR2X1   g1096(.A(n2935), .B(n2249), .Y(n1166));
MX2X1    g1097(.A(g1711), .B(g1712), .S0(n2485_1), .Y(n1171));
AND2X1   g1098(.A(g1133), .B(g109), .Y(n1176));
MX2X1    g1099(.A(g1806), .B(g1333), .S0(n2907_1), .Y(n1181));
MX2X1    g1100(.A(g554), .B(g207), .S0(g18), .Y(n2942));
XOR2X1   g1101(.A(n2942), .B(g158), .Y(n2941));
AND2X1   g1102(.A(n2941), .B(g109), .Y(n1186));
MX2X1    g1103(.A(g962), .B(g853), .S0(n2816), .Y(n1191));
NAND2X1  g1104(.A(g762), .B(g758), .Y(n2944));
XOR2X1   g1105(.A(n2944), .B(g766), .Y(n2945));
NOR3X1   g1106(.A(n2945), .B(g590), .C(n2249), .Y(n1196));
AND2X1   g1107(.A(g486), .B(g109), .Y(n2947_1));
MX2X1    g1108(.A(g481), .B(n2947_1), .S0(n2413), .Y(n1206));
INVX1    g1109(.A(n2413), .Y(n2949));
AOI21X1  g1110(.A0(n2519), .A1(n2949), .B0(g471), .Y(n2950));
NOR3X1   g1111(.A(n2950), .B(g868), .C(n2249), .Y(n1211));
AND2X1   g1112(.A(g192), .B(g109), .Y(n1216));
INVX1    g1113(.A(g1950), .Y(n2953));
NOR2X1   g1114(.A(n2331_1), .B(n2953), .Y(n2954));
MX2X1    g1115(.A(n2954), .B(g1941), .S0(n2766), .Y(n1226));
AND2X1   g1116(.A(n2841), .B(g632), .Y(n1236));
NOR3X1   g1117(.A(n2631), .B(g1216), .C(n2249), .Y(n1241));
NAND2X1  g1118(.A(n2263), .B(n2590_1), .Y(n2958));
MX2X1    g1119(.A(g1512), .B(g192), .S0(g18), .Y(n2959));
MX2X1    g1120(.A(n2959), .B(n2958), .S0(n2664), .Y(n2960));
MX2X1    g1121(.A(g549), .B(n2960), .S0(n2485_1), .Y(n1246));
MX2X1    g1122(.A(g95), .B(g1041), .S0(g85), .Y(n1251));
XOR2X1   g1123(.A(g1015), .B(g1019), .Y(n2963));
XOR2X1   g1124(.A(g1011), .B(g1007), .Y(n2964));
XOR2X1   g1125(.A(n2964), .B(n2963), .Y(n2965));
XOR2X1   g1126(.A(g999), .B(g1003), .Y(n2966));
XOR2X1   g1127(.A(g995), .B(g991), .Y(n2967_1));
XOR2X1   g1128(.A(n2967_1), .B(n2966), .Y(n2968));
XOR2X1   g1129(.A(n2968), .B(n2965), .Y(n2969));
XOR2X1   g1130(.A(n2969), .B(g1023), .Y(n2970));
XOR2X1   g1131(.A(n2970), .B(n2876), .Y(n2971));
OAI21X1  g1132(.A0(n2874), .A1(n2873), .B0(n2971), .Y(n2972_1));
MX2X1    g1133(.A(g105), .B(n2972_1), .S0(n2485_1), .Y(n1256));
AOI21X1  g1134(.A0(n2272), .A1(g109), .B0(n2591), .Y(n2974));
MX2X1    g1135(.A(g1669), .B(n2974), .S0(n2572), .Y(n1261));
AND2X1   g1136(.A(g231), .B(g109), .Y(n1266));
MX2X1    g1137(.A(g1499), .B(g1531), .S0(n2509), .Y(n1271));
AND2X1   g1138(.A(g1453), .B(g109), .Y(n1276));
OAI21X1  g1139(.A0(n2004), .A1(n2249), .B0(n2590_1), .Y(n2979));
MX2X1    g1140(.A(n2788), .B(n2979), .S0(n2664), .Y(n2980));
MX2X1    g1141(.A(g572), .B(n2980), .S0(n2485_1), .Y(n1281));
MX2X1    g1142(.A(g1059), .B(g1092), .S0(n2485_1), .Y(n2982_1));
MX2X1    g1143(.A(g1011), .B(n2982_1), .S0(n2485_1), .Y(n1286));
OAI21X1  g1144(.A0(n2060), .A1(n2028), .B0(n2006), .Y(n2984));
OAI21X1  g1145(.A0(n2061), .A1(n2006), .B0(n2984), .Y(n1291));
AND2X1   g1146(.A(g1424), .B(g109), .Y(n1296));
MX2X1    g1147(.A(g1074), .B(g342), .S0(n2572), .Y(n1301));
AND2X1   g1148(.A(g444), .B(g109), .Y(n2988));
MX2X1    g1149(.A(g448), .B(n2988), .S0(n2413), .Y(n1306));
MX2X1    g1150(.A(g1630), .B(g237), .S0(g18), .Y(n2990));
XOR2X1   g1151(.A(n2990), .B(n2610_1), .Y(n2991));
NOR2X1   g1152(.A(n2991), .B(n2249), .Y(n1311));
MX2X1    g1153(.A(g1080), .B(g348), .S0(n2572), .Y(n1316));
MX2X1    g1154(.A(g1713), .B(g1710), .S0(n2485_1), .Y(n1321));
MX2X1    g1155(.A(g148), .B(g269), .S0(n2670), .Y(n1331));
AND2X1   g1156(.A(g401), .B(g109), .Y(n2996));
MX2X1    g1157(.A(g396), .B(n2996), .S0(n2413), .Y(n1336));
OAI21X1  g1158(.A0(n2343), .A1(n2851), .B0(n2322), .Y(n2998));
AND2X1   g1159(.A(n2308), .B(n2309), .Y(n2999));
OAI21X1  g1160(.A0(n2998), .A1(n2344), .B0(n2999), .Y(n3000));
OAI21X1  g1161(.A0(n2308), .A1(n2309), .B0(n3000), .Y(n3001));
MX2X1    g1162(.A(n2491), .B(n2004), .S0(g1690), .Y(n3002_1));
MX2X1    g1163(.A(n2484), .B(n1983), .S0(g1690), .Y(n3003));
MX2X1    g1164(.A(n2496), .B(n2246_1), .S0(g1690), .Y(n3004));
INVX1    g1165(.A(n2223), .Y(n3005));
MX2X1    g1166(.A(n2494), .B(n3005), .S0(g1690), .Y(n3006));
OAI22X1  g1167(.A0(n3004), .A1(n3006), .B0(n3003), .B1(n3002_1), .Y(n3007_1));
INVX1    g1168(.A(g1690), .Y(n3008));
NAND2X1  g1169(.A(g1781), .B(n3008), .Y(n3009));
OAI21X1  g1170(.A0(n2192), .A1(n2166_1), .B0(g1690), .Y(n3010));
NAND2X1  g1171(.A(g1776), .B(n3008), .Y(n3011));
OAI21X1  g1172(.A0(n2152), .A1(n2124), .B0(g1690), .Y(n3012_1));
AOI22X1  g1173(.A0(n3011), .A1(n3012_1), .B0(n3010), .B1(n3009), .Y(n3013));
NAND2X1  g1174(.A(n3008), .B(g1771), .Y(n3014));
OAI21X1  g1175(.A0(n2111_1), .A1(n2077_1), .B0(g1690), .Y(n3015));
AOI21X1  g1176(.A0(n2392), .A1(n2382), .B0(n3008), .Y(n3016));
AOI21X1  g1177(.A0(n3008), .A1(g1766), .B0(n3016), .Y(n3017_1));
AOI21X1  g1178(.A0(n3015), .A1(n3014), .B0(n3017_1), .Y(n3018));
OAI21X1  g1179(.A0(n3018), .A1(n3013), .B0(n3007_1), .Y(n3019));
MX2X1    g1180(.A(n3001), .B(n3019), .S0(n2331_1), .Y(n1341));
AOI21X1  g1181(.A0(g115), .A1(g18), .B0(g9), .Y(n3021));
NOR2X1   g1182(.A(n3021), .B(n2249), .Y(n1346));
MX2X1    g1183(.A(g664), .B(g736), .S0(n2567), .Y(n3023));
OR2X1    g1184(.A(n3023), .B(n2462), .Y(n1351));
MX2X1    g1185(.A(g965), .B(g857), .S0(n2816), .Y(n1356));
AND2X1   g1186(.A(g248), .B(g109), .Y(n1361));
NOR2X1   g1187(.A(n2796), .B(n2795), .Y(n3027_1));
XOR2X1   g1188(.A(n3027_1), .B(n2793), .Y(n3028));
NOR4X1   g1189(.A(n2302), .B(n2791), .C(n2249), .D(n3028), .Y(n1371));
AND2X1   g1190(.A(g1365), .B(g109), .Y(n1376));
OAI21X1  g1191(.A0(g1703), .A1(g1696), .B0(g557), .Y(n3031));
NAND2X1  g1192(.A(n3031), .B(n2804), .Y(n1381));
AND2X1   g1193(.A(g207), .B(g109), .Y(n1396));
MX2X1    g1194(.A(g557), .B(g213), .S0(g18), .Y(n2226));
XOR2X1   g1195(.A(n2226), .B(g162), .Y(n3035));
AND2X1   g1196(.A(n3035), .B(g109), .Y(n1401));
AND2X1   g1197(.A(n2841), .B(g635), .Y(n1406));
MX2X1    g1198(.A(g1041), .B(g1071), .S0(n2485_1), .Y(n3038));
MX2X1    g1199(.A(g1023), .B(n3038), .S0(n2485_1), .Y(n1411));
MX2X1    g1200(.A(g1796), .B(g1327), .S0(n2907_1), .Y(n1426));
XOR2X1   g1201(.A(n2432), .B(n2431_1), .Y(n3041));
MX2X1    g1202(.A(n2431_1), .B(n3041), .S0(g627), .Y(n3042_1));
NAND3X1  g1203(.A(n3042_1), .B(n2734), .C(n2433), .Y(n1431));
MX2X1    g1204(.A(g135), .B(g293), .S0(n2670), .Y(n1436));
INVX1    g1205(.A(n2485_1), .Y(n3045));
NOR4X1   g1206(.A(n2601), .B(n2845), .C(n3045), .D(n2905), .Y(n2121));
AND2X1   g1207(.A(g1341), .B(g1336), .Y(n3047_1));
XOR2X1   g1208(.A(n3047_1), .B(n2125), .Y(n3048));
MX2X1    g1209(.A(n2125), .B(n3048), .S0(n2121), .Y(n3049));
AOI21X1  g1210(.A0(g108), .A1(g109), .B0(n2286_1), .Y(n1581));
NAND2X1  g1211(.A(n1581), .B(g1212), .Y(n3051));
NAND2X1  g1212(.A(n3051), .B(g109), .Y(n3052_1));
NOR2X1   g1213(.A(n3052_1), .B(n3049), .Y(n1441));
NOR4X1   g1214(.A(n2632), .B(g1101), .C(g1104), .D(g1107), .Y(n3054));
XOR2X1   g1215(.A(n3054), .B(g1141), .Y(n3055));
MX2X1    g1216(.A(g231), .B(n3055), .S0(n2630), .Y(n3056));
MX2X1    g1217(.A(g1633), .B(n3056), .S0(n2485_1), .Y(n1446));
MX2X1    g1218(.A(g1753), .B(g1791), .S0(n2292), .Y(n1451));
AND2X1   g1219(.A(g1504), .B(g109), .Y(n1456));
AND2X1   g1220(.A(g1240), .B(g109), .Y(n3060));
MX2X1    g1221(.A(g1235), .B(n3060), .S0(n2601), .Y(n1461));
AND2X1   g1222(.A(g538), .B(g109), .Y(n3062_1));
MX2X1    g1223(.A(g542), .B(n3062_1), .S0(n2413), .Y(n1466));
AND2X1   g1224(.A(g416), .B(g109), .Y(n3064));
MX2X1    g1225(.A(g411), .B(n3064), .S0(n2413), .Y(n1471));
AND2X1   g1226(.A(g542), .B(g109), .Y(n3066));
MX2X1    g1227(.A(g476), .B(n3066), .S0(n2413), .Y(n1476));
NAND2X1  g1228(.A(n2782_1), .B(n2592), .Y(n3068));
OAI21X1  g1229(.A0(n2591), .A1(n2260), .B0(n3068), .Y(n3069));
MX2X1    g1230(.A(g1681), .B(n3069), .S0(n2485_1), .Y(n1481));
XOR2X1   g1231(.A(g374), .B(g369), .Y(n3071));
MX2X1    g1232(.A(g374), .B(n3071), .S0(n2580_1), .Y(n3072_1));
AND2X1   g1233(.A(n3072_1), .B(n2582), .Y(n1486));
MX2X1    g1234(.A(g563), .B(n2743_1), .S0(n2485_1), .Y(n1491));
INVX1    g1235(.A(g1914), .Y(n3075));
NOR2X1   g1236(.A(n2331_1), .B(n3075), .Y(n3076_1));
MX2X1    g1237(.A(n3076_1), .B(g1905), .S0(n2766), .Y(n1496));
AND2X1   g1238(.A(g530), .B(g109), .Y(n3078));
MX2X1    g1239(.A(g534), .B(n3078), .S0(n2413), .Y(n1501));
MX2X1    g1240(.A(g575), .B(n2667), .S0(n2485_1), .Y(n1506));
INVX1    g1241(.A(g1936), .Y(n3081_1));
INVX1    g1242(.A(g1941), .Y(n3082));
INVX1    g1243(.A(n2339), .Y(n3083));
MX2X1    g1244(.A(n2336_1), .B(n3083), .S0(n2326_1), .Y(n3084));
MX2X1    g1245(.A(n3082), .B(n3084), .S0(n2319), .Y(n3085));
XOR2X1   g1246(.A(n3085), .B(g1936), .Y(n3086_1));
MX2X1    g1247(.A(n3081_1), .B(n3086_1), .S0(n2320), .Y(n3087));
OAI21X1  g1248(.A0(n3087), .A1(n2342), .B0(n2348), .Y(n1511));
OR2X1    g1249(.A(n2681), .B(g55), .Y(n1516));
AND2X1   g1250(.A(g1117), .B(g109), .Y(n1521));
OAI21X1  g1251(.A0(g754), .A1(n2680), .B0(g357), .Y(n3091_1));
INVX1    g1252(.A(g324), .Y(n3092));
NOR4X1   g1253(.A(n2728_1), .B(g471), .C(g461), .D(n2756), .Y(n3093));
XOR2X1   g1254(.A(n3093), .B(g496), .Y(n3094));
INVX1    g1255(.A(n3094), .Y(n3095));
MX2X1    g1256(.A(n3095), .B(n3092), .S0(n2413), .Y(n3096_1));
OAI21X1  g1257(.A0(n3096_1), .A1(n2682), .B0(n3091_1), .Y(n1531));
AND2X1   g1258(.A(g386), .B(g109), .Y(n3098));
MX2X1    g1259(.A(g426), .B(n3098), .S0(n2413), .Y(n1536));
MX2X1    g1260(.A(g1440), .B(g1601), .S0(n2574), .Y(n1541));
MX2X1    g1261(.A(g553), .B(n2974), .S0(n2485_1), .Y(n1546));
AND2X1   g1262(.A(g143), .B(g109), .Y(n1551));
AND2X1   g1263(.A(g501), .B(g109), .Y(n3103));
MX2X1    g1264(.A(g496), .B(n3103), .S0(n2413), .Y(n1556));
MX2X1    g1265(.A(g572), .B(g243), .S0(g18), .Y(n1561));
AOI22X1  g1266(.A0(n2318), .A1(n2308), .B0(g1950), .B1(n2766), .Y(n3106_1));
XOR2X1   g1267(.A(n3106_1), .B(g1840), .Y(n3107));
NOR2X1   g1268(.A(n3107), .B(n2630), .Y(n1566));
AND2X1   g1269(.A(n2682), .B(g70), .Y(n1571));
NAND4X1  g1270(.A(g794), .B(g745), .C(g109), .D(g746), .Y(n1585));
OAI21X1  g1271(.A0(n2192), .A1(n2166_1), .B0(n2006), .Y(n3111));
OAI21X1  g1272(.A0(n2193), .A1(n2006), .B0(n3111), .Y(n1590));
MX2X1    g1273(.A(g143), .B(g302), .S0(n2670), .Y(n1595));
INVX1    g1274(.A(g471), .Y(n3114));
NOR4X1   g1275(.A(g466), .B(n3114), .C(g461), .D(n2756), .Y(n3115));
XOR2X1   g1276(.A(n3115), .B(g516), .Y(n3116));
MX2X1    g1277(.A(n3116), .B(g309), .S0(n2413), .Y(n3117));
MX2X1    g1278(.A(g342), .B(n3117), .S0(n2681), .Y(n1600));
AND2X1   g1279(.A(g1250), .B(g109), .Y(n3119));
MX2X1    g1280(.A(g1245), .B(n3119), .S0(n2601), .Y(n1605));
AND2X1   g1281(.A(g1163), .B(g109), .Y(n1610));
MX2X1    g1282(.A(g1044), .B(g1077), .S0(n2485_1), .Y(n3122));
MX2X1    g1283(.A(g1032), .B(n3122), .S0(n2485_1), .Y(n1620));
NOR4X1   g1284(.A(g1110), .B(g1101), .C(n2620_1), .D(n2672), .Y(n3124));
XOR2X1   g1285(.A(n3124), .B(g1133), .Y(n3125));
MX2X1    g1286(.A(g219), .B(n3125), .S0(n2630), .Y(n3126));
XOR2X1   g1287(.A(n3126), .B(g1436), .Y(n3127));
AND2X1   g1288(.A(n3127), .B(g109), .Y(n1625));
MX2X1    g1289(.A(g89), .B(g1053), .S0(g85), .Y(n1630));
XOR2X1   g1290(.A(g1508), .B(g1499), .Y(n3130));
XOR2X1   g1291(.A(n3130), .B(n2625), .Y(n3131));
XOR2X1   g1292(.A(n3131), .B(g1453), .Y(n3132));
NOR2X1   g1293(.A(n3132), .B(n2249), .Y(n1635));
NOR4X1   g1294(.A(n2728_1), .B(g471), .C(n2755), .D(n2756), .Y(n3134));
XOR2X1   g1295(.A(n3134), .B(g506), .Y(n3135));
MX2X1    g1296(.A(n3135), .B(g330), .S0(n2413), .Y(n3136));
MX2X1    g1297(.A(g363), .B(n3136), .S0(n2681), .Y(n1640));
AND2X1   g1298(.A(g1157), .B(g109), .Y(n1650));
NOR2X1   g1299(.A(n2485_1), .B(n2646), .Y(n1655));
OAI21X1  g1300(.A0(n2152), .A1(n2124), .B0(n2006), .Y(n3140));
OAI21X1  g1301(.A0(n2153), .A1(n2006), .B0(n3140), .Y(n1660));
NOR2X1   g1302(.A(n2528), .B(n2036), .Y(n1665));
MX2X1    g1303(.A(g569), .B(g237), .S0(g18), .Y(n1670));
AND2X1   g1304(.A(g516), .B(g109), .Y(n3144));
MX2X1    g1305(.A(g511), .B(n3144), .S0(n2413), .Y(n1675));
MX2X1    g1306(.A(g575), .B(g248), .S0(g18), .Y(n1680));
NOR2X1   g1307(.A(n2617), .B(n2639_1), .Y(n3147));
XOR2X1   g1308(.A(n3147), .B(n2640), .Y(n3148));
NOR3X1   g1309(.A(n3148), .B(g590), .C(n2249), .Y(n1685));
MX2X1    g1310(.A(g1627), .B(n3126), .S0(n2485_1), .Y(n1695));
AND2X1   g1311(.A(g1292), .B(g109), .Y(n3151));
MX2X1    g1312(.A(g1296), .B(n3151), .S0(n2601), .Y(n1700));
MX2X1    g1313(.A(g131), .B(g290), .S0(n2670), .Y(n1705));
AND2X1   g1314(.A(n2852_1), .B(g1849), .Y(n1710));
NAND3X1  g1315(.A(g762), .B(g766), .C(g758), .Y(n3155));
XOR2X1   g1316(.A(n3155), .B(g770), .Y(n3156));
NOR3X1   g1317(.A(n3156), .B(g590), .C(n2249), .Y(n1715));
MX2X1    g1318(.A(g1424), .B(g1583), .S0(n2574), .Y(n1720));
XOR2X1   g1319(.A(n2518), .B(g466), .Y(n3159));
MX2X1    g1320(.A(g466), .B(n3159), .S0(n2520_1), .Y(n3160));
AND2X1   g1321(.A(n3160), .B(n2523), .Y(n1725));
MX2X1    g1322(.A(g1458), .B(g1561), .S0(n2509), .Y(n1730));
ZERO     g1323(.Y(n1735));
MX2X1    g1324(.A(g1478), .B(g1546), .S0(n2509), .Y(n1740));
MX2X1    g1325(.A(g127), .B(g287), .S0(n2670), .Y(n1745));
MX2X1    g1326(.A(g560), .B(n3069), .S0(n2485_1), .Y(n1750));
AOI22X1  g1327(.A0(n2444), .A1(n2434), .B0(g736), .B1(n2567), .Y(n3167));
XOR2X1   g1328(.A(n3167), .B(g617), .Y(n3168));
NOR2X1   g1329(.A(n3168), .B(n2630), .Y(n1755));
INVX1    g1330(.A(n2841), .Y(n1760));
OAI21X1  g1331(.A0(g754), .A1(n2680), .B0(g336), .Y(n3171));
INVX1    g1332(.A(n2875), .Y(n3172));
INVX1    g1333(.A(g312), .Y(n3173));
NOR4X1   g1334(.A(g466), .B(n3114), .C(n2755), .D(g456), .Y(n3174));
XOR2X1   g1335(.A(n3174), .B(g476), .Y(n3175));
INVX1    g1336(.A(n3175), .Y(n3176));
MX2X1    g1337(.A(n3176), .B(n3173), .S0(n2413), .Y(n3177));
INVX1    g1338(.A(g333), .Y(n3178));
NOR4X1   g1339(.A(g466), .B(n3114), .C(g461), .D(g456), .Y(n3179));
XOR2X1   g1340(.A(n3179), .B(g511), .Y(n3180));
INVX1    g1341(.A(n3180), .Y(n3181));
MX2X1    g1342(.A(n3181), .B(n3178), .S0(n2413), .Y(n3182));
XOR2X1   g1343(.A(n3182), .B(n3117), .Y(n3183));
INVX1    g1344(.A(g327), .Y(n3184));
NOR4X1   g1345(.A(n2728_1), .B(g471), .C(n2755), .D(g456), .Y(n3185));
XOR2X1   g1346(.A(n3185), .B(g501), .Y(n3186));
INVX1    g1347(.A(n3186), .Y(n3187));
MX2X1    g1348(.A(n3187), .B(n3184), .S0(n2413), .Y(n3188));
XOR2X1   g1349(.A(n3188), .B(n3136), .Y(n3189));
XOR2X1   g1350(.A(n3189), .B(n3183), .Y(n3190));
XOR2X1   g1351(.A(n3096_1), .B(n2732), .Y(n3191));
INVX1    g1352(.A(g315), .Y(n3192));
NOR4X1   g1353(.A(g466), .B(g471), .C(n2755), .D(g456), .Y(n3193));
XOR2X1   g1354(.A(n3193), .B(g481), .Y(n3194));
INVX1    g1355(.A(n3194), .Y(n3195));
MX2X1    g1356(.A(n3195), .B(n3192), .S0(n2413), .Y(n3196));
XOR2X1   g1357(.A(n3196), .B(n2759), .Y(n3197));
XOR2X1   g1358(.A(n3197), .B(n3191), .Y(n3198));
XOR2X1   g1359(.A(n3198), .B(n3190), .Y(n3199));
XOR2X1   g1360(.A(n3199), .B(n3177), .Y(n3200));
NOR2X1   g1361(.A(n3200), .B(n3172), .Y(n3201));
NOR4X1   g1362(.A(g466), .B(g471), .C(g461), .D(n2756), .Y(n3202));
NOR4X1   g1363(.A(g506), .B(g516), .C(g501), .D(g511), .Y(n3203));
NOR4X1   g1364(.A(g491), .B(g486), .C(g496), .D(g481), .Y(n3204));
NOR3X1   g1365(.A(g534), .B(g521), .C(g530), .Y(n3205));
NOR4X1   g1366(.A(g476), .B(g542), .C(g538), .D(g525), .Y(n3206));
NAND4X1  g1367(.A(n3205), .B(n3204), .C(n3203), .D(n3206), .Y(n3207));
INVX1    g1368(.A(g521), .Y(n3208));
XOR2X1   g1369(.A(g525), .B(n3208), .Y(n3209));
AND2X1   g1370(.A(n3209), .B(n3207), .Y(n3210));
XOR2X1   g1371(.A(n3210), .B(n3202), .Y(n3211));
MX2X1    g1372(.A(n3211), .B(n2533), .S0(n2413), .Y(n3212));
OAI21X1  g1373(.A0(n3212), .A1(n2875), .B0(n2681), .Y(n3213));
OAI21X1  g1374(.A0(n3213), .A1(n3201), .B0(n3171), .Y(n1765));
XOR2X1   g1375(.A(n2520_1), .B(g456), .Y(n3215));
AND2X1   g1376(.A(n3215), .B(n2523), .Y(n1770));
XOR2X1   g1377(.A(n3212), .B(n3200), .Y(n3217));
MX2X1    g1378(.A(g345), .B(n3217), .S0(n2681), .Y(n1780));
XOR2X1   g1379(.A(g1771), .B(g1766), .Y(n3219));
MX2X1    g1380(.A(g1771), .B(n3219), .S0(n2708_1), .Y(n3220));
AND2X1   g1381(.A(n3220), .B(n2600_1), .Y(n1790));
AND2X1   g1382(.A(n2642), .B(g786), .Y(n3222));
AND2X1   g1383(.A(n3222), .B(g790), .Y(n3223));
XOR2X1   g1384(.A(n3223), .B(g590), .Y(n1795));
MX2X1    g1385(.A(g549), .B(g192), .S0(g18), .Y(n1800));
INVX1    g1386(.A(g1945), .Y(n3226));
OR2X1    g1387(.A(n2336_1), .B(g1936), .Y(n3227));
NAND2X1  g1388(.A(n2339), .B(g1936), .Y(n3228));
MX2X1    g1389(.A(n3227), .B(n3228), .S0(n2326_1), .Y(n3229));
MX2X1    g1390(.A(n2953), .B(n3229), .S0(n2319), .Y(n3230));
XOR2X1   g1391(.A(n3230), .B(g1945), .Y(n3231));
MX2X1    g1392(.A(n3226), .B(n3231), .S0(n2320), .Y(n3232));
OAI21X1  g1393(.A0(n3232), .A1(n2342), .B0(n2348), .Y(n1805));
MX2X1    g1394(.A(g1738), .B(g1766), .S0(n2292), .Y(n1810));
MX2X1    g1395(.A(g1627), .B(g231), .S0(g18), .Y(n3235));
XOR2X1   g1396(.A(n3235), .B(n2611), .Y(n3236));
NOR2X1   g1397(.A(n3236), .B(n2249), .Y(n1815));
MX2X1    g1398(.A(g86), .B(g1035), .S0(g85), .Y(n1820));
XOR2X1   g1399(.A(g1690), .B(g1707), .Y(n3239));
AND2X1   g1400(.A(n3239), .B(g1700), .Y(n1830));
XOR2X1   g1401(.A(n2741), .B(n2612), .Y(n3241));
NOR2X1   g1402(.A(n3241), .B(n2249), .Y(n1835));
NOR3X1   g1403(.A(n2632), .B(g1216), .C(n2249), .Y(n1840));
MX2X1    g1404(.A(g139), .B(g296), .S0(n2670), .Y(n1845));
MX2X1    g1405(.A(g1663), .B(n2960), .S0(n2572), .Y(n1850));
NOR2X1   g1406(.A(n2462), .B(n2511), .Y(n3246));
MX2X1    g1407(.A(n3246), .B(g691), .S0(n2567), .Y(n1855));
MX2X1    g1408(.A(g1762), .B(g1806), .S0(n2292), .Y(n1860));
OAI21X1  g1409(.A0(g754), .A1(n2680), .B0(g360), .Y(n3249));
OAI21X1  g1410(.A0(n3188), .A1(n2682), .B0(n3249), .Y(n1865));
AND2X1   g1411(.A(g1389), .B(g109), .Y(n1870));
MX2X1    g1412(.A(g1657), .B(n2980), .S0(n2572), .Y(n1875));
INVX1    g1413(.A(g727), .Y(n3253));
MX2X1    g1414(.A(n2470_1), .B(n2463), .S0(n2454), .Y(n3254));
MX2X1    g1415(.A(n3253), .B(n3254), .S0(n2445_1), .Y(n3255));
XOR2X1   g1416(.A(n3255), .B(g722), .Y(n3256));
MX2X1    g1417(.A(n2466), .B(n3256), .S0(n2446), .Y(n3257));
OAI21X1  g1418(.A0(n3257), .A1(n2473), .B0(n2478), .Y(n1880));
OR2X1    g1419(.A(n2681), .B(g61), .Y(n1885));
OAI21X1  g1420(.A0(g1703), .A1(g1696), .B0(g566), .Y(n3260));
AOI21X1  g1421(.A0(n2246_1), .A1(g109), .B0(n2591), .Y(n3261));
AND2X1   g1422(.A(n3235), .B(n2592), .Y(n3262));
OAI21X1  g1423(.A0(n3262), .A1(n3261), .B0(n2485_1), .Y(n3263));
NAND2X1  g1424(.A(n3263), .B(n3260), .Y(n1890));
NOR2X1   g1425(.A(g1393), .B(g1394), .Y(n3265));
NOR3X1   g1426(.A(n3265), .B(g115), .C(n2249), .Y(n1895));
MX2X1    g1427(.A(g1089), .B(g357), .S0(n2572), .Y(n1900));
NOR4X1   g1428(.A(n2036), .B(n2091_1), .C(n2177), .D(n2135), .Y(n1905));
MX2X1    g1429(.A(g1071), .B(g339), .S0(n2572), .Y(n1909));
XOR2X1   g1430(.A(n2695), .B(g986), .Y(n3270));
MX2X1    g1431(.A(n2370), .B(n3270), .S0(n639), .Y(n3271));
NOR2X1   g1432(.A(n3271), .B(n2564), .Y(n1914));
XOR2X1   g1433(.A(n639), .B(n2043), .Y(n3273));
NOR2X1   g1434(.A(n3273), .B(n2564), .Y(n1919));
INVX1    g1435(.A(g153), .Y(n3275));
XOR2X1   g1436(.A(g182), .B(g148), .Y(n3276));
XOR2X1   g1437(.A(n3276), .B(n3275), .Y(n3277));
XOR2X1   g1438(.A(n3277), .B(g143), .Y(n3278));
NOR2X1   g1439(.A(n3278), .B(n2249), .Y(n1928));
INVX1    g1440(.A(n2341_1), .Y(n3280));
NOR4X1   g1441(.A(n2343), .B(g1822), .C(n2851), .D(n3280), .Y(n3281));
AND2X1   g1442(.A(n2313), .B(n2308), .Y(n3282));
INVX1    g1443(.A(n3282), .Y(n3283));
AOI21X1  g1444(.A0(n2324), .A1(n3283), .B0(n3280), .Y(n3284));
NOR2X1   g1445(.A(n3284), .B(n3281), .Y(n3285));
XOR2X1   g1446(.A(n3285), .B(g1814), .Y(n3286));
NOR2X1   g1447(.A(n3286), .B(n2630), .Y(n1933));
MX2X1    g1448(.A(g94), .B(g1038), .S0(g85), .Y(n1938));
INVX1    g1449(.A(g1923), .Y(n3289));
NAND2X1  g1450(.A(n2335), .B(n2334), .Y(n3290));
OR2X1    g1451(.A(n2338), .B(n2334), .Y(n3291));
MX2X1    g1452(.A(n3290), .B(n3291), .S0(n2326_1), .Y(n3292));
MX2X1    g1453(.A(n3289), .B(n3292), .S0(n2319), .Y(n3293));
XOR2X1   g1454(.A(n3293), .B(g1918), .Y(n3294));
MX2X1    g1455(.A(n2333), .B(n3294), .S0(n2320), .Y(n3295));
OAI21X1  g1456(.A0(n3295), .A1(n2342), .B0(n2348), .Y(n1947));
NOR3X1   g1457(.A(n2617), .B(n2640), .C(n2639_1), .Y(n3297));
XOR2X1   g1458(.A(n3297), .B(n2641), .Y(n3298));
NOR3X1   g1459(.A(n3298), .B(g590), .C(n2249), .Y(n1952));
AND2X1   g1460(.A(n2341_1), .B(n2344), .Y(n3300));
NOR3X1   g1461(.A(n3280), .B(g1828), .C(n2322), .Y(n3301));
NOR3X1   g1462(.A(n3301), .B(n3300), .C(n3281), .Y(n3302));
XOR2X1   g1463(.A(n3302), .B(g1822), .Y(n3303));
NOR2X1   g1464(.A(n3303), .B(n2630), .Y(n1957));
AND2X1   g1465(.A(g1362), .B(g109), .Y(n1962));
MX2X1    g1466(.A(g92), .B(g1062), .S0(g85), .Y(n1972));
XOR2X1   g1467(.A(n2959), .B(g1458), .Y(n3307));
AND2X1   g1468(.A(n3307), .B(g109), .Y(n1977));
AND2X1   g1469(.A(g148), .B(g109), .Y(n1982));
OAI21X1  g1470(.A0(g754), .A1(n2680), .B0(g366), .Y(n3310));
OAI21X1  g1471(.A0(n3182), .A1(n2682), .B0(n3310), .Y(n1987));
NAND2X1  g1472(.A(g605), .B(g591), .Y(n3312));
NOR3X1   g1473(.A(n3312), .B(n2475_1), .C(g599), .Y(n3313));
AND2X1   g1474(.A(n2472), .B(n2474), .Y(n3314));
NOR3X1   g1475(.A(n2475_1), .B(g605), .C(n2436_1), .Y(n3315));
NOR3X1   g1476(.A(n3315), .B(n3314), .C(n3313), .Y(n3316));
XOR2X1   g1477(.A(n3316), .B(g599), .Y(n3317));
NOR2X1   g1478(.A(n3317), .B(n2630), .Y(n1997));
AOI22X1  g1479(.A0(g1828), .A1(g1814), .B0(g1840), .B1(g1834), .Y(n3319));
OAI21X1  g1480(.A0(n2312), .A1(g1840), .B0(n3319), .Y(n3320));
MX2X1    g1481(.A(n2323), .B(n3320), .S0(n2309), .Y(n3321));
XOR2X1   g1482(.A(n3321), .B(n2740), .Y(n3322));
NAND4X1  g1483(.A(n2347), .B(n2324), .C(n2317), .D(n3319), .Y(n3323));
NAND4X1  g1484(.A(n2852_1), .B(n2345), .C(g1850), .D(n3323), .Y(n3324));
NOR2X1   g1485(.A(n3324), .B(n3322), .Y(n3325));
MX2X1    g1486(.A(n2345), .B(n3325), .S0(g1854), .Y(n3326));
INVX1    g1487(.A(g1806), .Y(n3327));
OAI21X1  g1488(.A0(n3327), .A1(g1690), .B0(n2331_1), .Y(n3328));
OAI22X1  g1489(.A0(n3326), .A1(n2331_1), .B0(n3016), .B1(n3328), .Y(n2002));
MX2X1    g1490(.A(g944), .B(g829), .S0(n2816), .Y(n2007));
NOR2X1   g1491(.A(n2331_1), .B(n3082), .Y(n3331));
MX2X1    g1492(.A(n3331), .B(g1932), .S0(n2766), .Y(n2012));
MX2X1    g1493(.A(g566), .B(g231), .S0(g18), .Y(n2658));
XOR2X1   g1494(.A(n2658), .B(g127), .Y(n3334));
AND2X1   g1495(.A(n3334), .B(g109), .Y(n2017));
AND2X1   g1496(.A(g1515), .B(g109), .Y(n2022));
INVX1    g1497(.A(g691), .Y(n3337));
OR2X1    g1498(.A(g658), .B(g668), .Y(n3338));
OR2X1    g1499(.A(n3338), .B(g677), .Y(n3339));
MX2X1    g1500(.A(n2456), .B(n3339), .S0(n2454), .Y(n3340));
MX2X1    g1501(.A(n3337), .B(n3340), .S0(n2445_1), .Y(n3341));
XOR2X1   g1502(.A(n3341), .B(g686), .Y(n3342));
MX2X1    g1503(.A(n2455_1), .B(n3342), .S0(n2446), .Y(n3343));
OAI21X1  g1504(.A0(n3343), .A1(n2473), .B0(n2478), .Y(n2027));
MX2X1    g1505(.A(g953), .B(g841), .S0(n2816), .Y(n2032));
NAND3X1  g1506(.A(g1776), .B(g1771), .C(g1766), .Y(n3346));
INVX1    g1507(.A(g1781), .Y(n3347));
NAND4X1  g1508(.A(g1690), .B(g1707), .C(g1786), .D(n3347), .Y(n3348));
NAND4X1  g1509(.A(g1796), .B(g1801), .C(g1791), .D(g1806), .Y(n3349));
NOR3X1   g1510(.A(n3349), .B(n3348), .C(n3346), .Y(n2037));
OR2X1    g1511(.A(n2004), .B(n1892), .Y(n3351));
OR2X1    g1512(.A(n2004), .B(n2006), .Y(n3352));
NAND2X1  g1513(.A(n3352), .B(n3351), .Y(n2042));
NOR2X1   g1514(.A(g1610), .B(g1737), .Y(n2047));
INVX1    g1515(.A(n2740), .Y(n3355));
MX2X1    g1516(.A(g1733), .B(n3355), .S0(n2785), .Y(n2052));
AND2X1   g1517(.A(g1270), .B(g109), .Y(n3357));
MX2X1    g1518(.A(g1265), .B(n3357), .S0(n2601), .Y(n2057));
INVX1    g1519(.A(g1610), .Y(n3359));
AOI21X1  g1520(.A0(n2571), .A1(g1696), .B0(n3359), .Y(n2062));
NOR3X1   g1521(.A(n2709), .B(n2496), .C(n2494), .Y(n3361));
XOR2X1   g1522(.A(n3361), .B(n2484), .Y(n3362));
MX2X1    g1523(.A(n2484), .B(n3362), .S0(n2708_1), .Y(n3363));
NOR2X1   g1524(.A(n3363), .B(g1713), .Y(n2067));
MX2X1    g1525(.A(g1791), .B(g1324), .S0(n2907_1), .Y(n2072));
MX2X1    g1526(.A(g1486), .B(g1540), .S0(n2509), .Y(n2077));
AND2X1   g1527(.A(g219), .B(g109), .Y(n2082));
NAND3X1  g1528(.A(g1341), .B(g1336), .C(g1346), .Y(n3368));
NOR2X1   g1529(.A(n3368), .B(n2167), .Y(n2087));
AND2X1   g1530(.A(g491), .B(g109), .Y(n3370));
MX2X1    g1531(.A(g486), .B(n3370), .S0(n2413), .Y(n2091));
AND2X1   g1532(.A(n2852_1), .B(g1848), .Y(n2096));
AND2X1   g1533(.A(g1377), .B(g109), .Y(n2101));
XOR2X1   g1534(.A(n3346), .B(g1781), .Y(n3374));
MX2X1    g1535(.A(n3347), .B(n3374), .S0(n2708_1), .Y(n3375));
NOR2X1   g1536(.A(n3375), .B(g1713), .Y(n2106));
INVX1    g1537(.A(g1905), .Y(n3377));
OR2X1    g1538(.A(g1872), .B(g1882), .Y(n3378));
OR2X1    g1539(.A(n3378), .B(g1891), .Y(n3379));
MX2X1    g1540(.A(n3379), .B(n2657), .S0(n2326_1), .Y(n3380));
MX2X1    g1541(.A(n3377), .B(n3380), .S0(n2319), .Y(n3381));
XOR2X1   g1542(.A(n3381), .B(g1900), .Y(n3382));
MX2X1    g1543(.A(n2656), .B(n3382), .S0(n2320), .Y(n3383));
OAI21X1  g1544(.A0(n3383), .A1(n2342), .B0(n2348), .Y(n2111));
AND2X1   g1545(.A(g1245), .B(g109), .Y(n3385));
MX2X1    g1546(.A(g1240), .B(n3385), .S0(n2601), .Y(n2116));
INVX1    g1547(.A(g627), .Y(n3387));
NAND2X1  g1548(.A(n2841), .B(n3387), .Y(n2126));
MX2X1    g1549(.A(g546), .B(g186), .S0(g18), .Y(n2431));
XOR2X1   g1550(.A(n2431), .B(n3275), .Y(n3390));
NOR2X1   g1551(.A(n3390), .B(n2249), .Y(n2131));
NOR2X1   g1552(.A(n2331_1), .B(n3289), .Y(n3392));
MX2X1    g1553(.A(n3392), .B(g1914), .S0(n2766), .Y(n2141));
NOR2X1   g1554(.A(n2528), .B(n2135), .Y(n2146));
MX2X1    g1555(.A(g1215), .B(g1209), .S0(n2485_1), .Y(n2151));
MX2X1    g1556(.A(g1776), .B(g1314), .S0(n2907_1), .Y(n2156));
XOR2X1   g1557(.A(n2121), .B(n2029), .Y(n3397));
NOR2X1   g1558(.A(n3397), .B(n3052_1), .Y(n2166));
MX2X1    g1559(.A(g153), .B(g272), .S0(n2670), .Y(n2171));
AND2X1   g1560(.A(n2811), .B(g1801), .Y(n3400));
XOR2X1   g1561(.A(n3400), .B(n3327), .Y(n3401));
MX2X1    g1562(.A(n3327), .B(n3401), .S0(n2708_1), .Y(n3402));
NOR2X1   g1563(.A(n3402), .B(g1713), .Y(n2176));
NAND2X1  g1564(.A(n2797_1), .B(g822), .Y(n3404));
XOR2X1   g1565(.A(n3404), .B(g826), .Y(n3405));
NOR4X1   g1566(.A(n2302), .B(n2791), .C(n2249), .D(n3405), .Y(n2181));
MX2X1    g1567(.A(g93), .B(g1065), .S0(g85), .Y(n2186));
NOR2X1   g1568(.A(n2331_1), .B(n2321_1), .Y(n3408));
MX2X1    g1569(.A(n3408), .B(g1878), .S0(n2766), .Y(n2191));
NAND2X1  g1570(.A(n2223), .B(n2006), .Y(n3410));
OAI21X1  g1571(.A0(n2224), .A1(n2006), .B0(n3410), .Y(n2196));
MX2X1    g1572(.A(g968), .B(g861), .S0(n2816), .Y(n2201));
AND2X1   g1573(.A(n2852_1), .B(g1853), .Y(n2206));
AND2X1   g1574(.A(g1137), .B(g109), .Y(n2211));
INVX1    g1575(.A(g1891), .Y(n3415));
NAND2X1  g1576(.A(g1872), .B(g1882), .Y(n3416));
MX2X1    g1577(.A(n3378), .B(n3416), .S0(n2326_1), .Y(n3417));
MX2X1    g1578(.A(n2767_1), .B(n3417), .S0(n2319), .Y(n3418));
XOR2X1   g1579(.A(n3418), .B(g1891), .Y(n3419));
MX2X1    g1580(.A(n3415), .B(n3419), .S0(n2320), .Y(n3420));
OAI21X1  g1581(.A0(n3420), .A1(n2342), .B0(n2348), .Y(n2216));
AND2X1   g1582(.A(g1255), .B(g109), .Y(n3422));
MX2X1    g1583(.A(g1250), .B(n3422), .S0(n2601), .Y(n2221));
NAND3X1  g1584(.A(n2870), .B(n1913), .C(n1887), .Y(n3424));
OR2X1    g1585(.A(n3424), .B(n1919_1), .Y(n2231));
AND2X1   g1586(.A(n2651), .B(n2434), .Y(n3426));
NOR2X1   g1587(.A(g591), .B(n2436_1), .Y(n3427));
AND2X1   g1588(.A(n2472), .B(n3427), .Y(n3428));
NOR3X1   g1589(.A(n3428), .B(n3426), .C(n3313), .Y(n3429));
XOR2X1   g1590(.A(n3429), .B(g591), .Y(n3430));
NOR2X1   g1591(.A(n3430), .B(n2630), .Y(n2236));
NAND2X1  g1592(.A(n2469), .B(g722), .Y(n3432));
MX2X1    g1593(.A(n3432), .B(n2464), .S0(n2454), .Y(n3433));
MX2X1    g1594(.A(n2770), .B(n3433), .S0(n2445_1), .Y(n3434));
XOR2X1   g1595(.A(n3434), .B(g731), .Y(n3435));
MX2X1    g1596(.A(n2467), .B(n3435), .S0(n2446), .Y(n3436));
OAI21X1  g1597(.A0(n3436), .A1(n2473), .B0(n2478), .Y(n2241));
NOR4X1   g1598(.A(g591), .B(g599), .C(g622), .D(n2437), .Y(n3438));
AND2X1   g1599(.A(g255), .B(g622), .Y(n3439));
AOI22X1  g1600(.A0(g591), .A1(g605), .B0(g617), .B1(g611), .Y(n3440));
INVX1    g1601(.A(n3440), .Y(n3441));
OR2X1    g1602(.A(n3441), .B(n2441), .Y(n3442));
MX2X1    g1603(.A(n3427), .B(n3442), .S0(n2435), .Y(n3443));
XOR2X1   g1604(.A(n3443), .B(n3439), .Y(n3444));
OR4X1    g1605(.A(n2477), .B(n3427), .C(n2444), .D(n3441), .Y(n3445));
INVX1    g1606(.A(n3438), .Y(n3446));
NAND4X1  g1607(.A(n3445), .B(n3444), .C(n1236), .D(n3446), .Y(n3447));
MX2X1    g1608(.A(n3438), .B(n3447), .S0(g636), .Y(n3448));
AND2X1   g1609(.A(g798), .B(g794), .Y(n3449));
AND2X1   g1610(.A(g802), .B(g806), .Y(n3450));
OR2X1    g1611(.A(n3450), .B(n3449), .Y(n3451));
OAI22X1  g1612(.A0(n2794), .A1(n2792_1), .B0(n2793), .B1(n2795), .Y(n3452));
NAND3X1  g1613(.A(n3452), .B(n3451), .C(g826), .Y(n3453));
MX2X1    g1614(.A(n3448), .B(n3453), .S0(n2462), .Y(n2246));
XOR2X1   g1615(.A(n2846), .B(g1218), .Y(n3455));
NOR3X1   g1616(.A(n3455), .B(g1212), .C(n2249), .Y(n2251));
INVX1    g1617(.A(n3314), .Y(n3457));
NAND4X1  g1618(.A(n2441), .B(n2434), .C(n2650), .D(n2472), .Y(n3458));
NAND2X1  g1619(.A(n2462), .B(g18), .Y(n3459));
NOR2X1   g1620(.A(n3312), .B(n2436_1), .Y(n3460));
OAI21X1  g1621(.A0(n3460), .A1(n2452), .B0(n2472), .Y(n3461));
NAND4X1  g1622(.A(n3459), .B(n3458), .C(n3457), .D(n3461), .Y(n3462));
XOR2X1   g1623(.A(n3462), .B(n2437), .Y(n3463));
NOR2X1   g1624(.A(n3463), .B(n2630), .Y(n2256));
AND2X1   g1625(.A(n2682), .B(g79), .Y(n2261));
AND2X1   g1626(.A(g178), .B(g109), .Y(n2266));
MX2X1    g1627(.A(g950), .B(g837), .S0(n2816), .Y(n2271));
AND2X1   g1628(.A(g1129), .B(g109), .Y(n2276));
AND2X1   g1629(.A(g448), .B(g109), .Y(n3469));
MX2X1    g1630(.A(g452), .B(n3469), .S0(n2413), .Y(n2286));
AND2X1   g1631(.A(g1828), .B(g1814), .Y(n3471));
AOI22X1  g1632(.A0(n2323), .A1(n2343), .B0(g1822), .B1(n3471), .Y(n3472));
AOI22X1  g1633(.A0(n2331_1), .A1(g18), .B0(n2344), .B1(n2341_1), .Y(n3473));
OAI21X1  g1634(.A0(n3472), .A1(n3280), .B0(n3473), .Y(n3474));
XOR2X1   g1635(.A(n3474), .B(n2343), .Y(n3475));
NOR2X1   g1636(.A(n3475), .B(n2630), .Y(n2291));
MX2X1    g1637(.A(g1727), .B(n2483), .S0(n2785), .Y(n2296));
MX2X1    g1638(.A(g1403), .B(g1592), .S0(n2574), .Y(n2301));
OR2X1    g1639(.A(g1959), .B(n1825), .Y(n2797));
XOR2X1   g1640(.A(g1703), .B(n2707), .Y(n3480));
NOR2X1   g1641(.A(n3480), .B(n2797), .Y(n2306));
NOR2X1   g1642(.A(n2331_1), .B(n2654), .Y(n3482));
MX2X1    g1643(.A(n3482), .B(g1923), .S0(n2766), .Y(n2311));
NOR4X1   g1644(.A(g1110), .B(n2631), .C(g1104), .D(n2672), .Y(n3484));
XOR2X1   g1645(.A(n3484), .B(g1129), .Y(n3485));
MX2X1    g1646(.A(g213), .B(n3485), .S0(n2630), .Y(n3486));
MX2X1    g1647(.A(g1624), .B(n3486), .S0(n2485_1), .Y(n2316));
XOR2X1   g1648(.A(g26), .B(g23), .Y(n2321));
MX2X1    g1649(.A(g1068), .B(g336), .S0(n2572), .Y(n2326));
AND2X1   g1650(.A(g440), .B(g109), .Y(n3490));
MX2X1    g1651(.A(g444), .B(n3490), .S0(n2413), .Y(n2336));
AND2X1   g1652(.A(g476), .B(g109), .Y(n3492));
MX2X1    g1653(.A(g516), .B(n3492), .S0(n2413), .Y(n2341));
AOI21X1  g1654(.A0(g115), .A1(g18), .B0(g119), .Y(n3494));
NOR2X1   g1655(.A(n3494), .B(n2249), .Y(n2346));
INVX1    g1656(.A(g668), .Y(n3496));
INVX1    g1657(.A(g673), .Y(n3497));
INVX1    g1658(.A(g658), .Y(n3498));
XOR2X1   g1659(.A(n2454), .B(n3498), .Y(n3499));
MX2X1    g1660(.A(n3497), .B(n3499), .S0(n2445_1), .Y(n3500));
XOR2X1   g1661(.A(n3500), .B(g668), .Y(n3501));
MX2X1    g1662(.A(n3496), .B(n3501), .S0(n2446), .Y(n3502));
OAI21X1  g1663(.A0(n3502), .A1(n2473), .B0(n2478), .Y(n2351));
XOR2X1   g1664(.A(n1800), .B(n2425), .Y(n3504));
NOR2X1   g1665(.A(n3504), .B(n2249), .Y(n2356));
AND2X1   g1666(.A(g1149), .B(g109), .Y(n2361));
OAI21X1  g1667(.A0(n2111_1), .A1(n2077_1), .B0(n2006), .Y(n3507));
OAI21X1  g1668(.A0(n2112), .A1(n2006), .B0(n3507), .Y(n2366));
NAND2X1  g1669(.A(n2852_1), .B(n2307), .Y(n2371));
MX2X1    g1670(.A(g182), .B(g263), .S0(n2670), .Y(n2376));
NOR3X1   g1671(.A(n2796), .B(n2795), .C(n2793), .Y(n3511));
XOR2X1   g1672(.A(n3511), .B(n2794), .Y(n3512));
NOR4X1   g1673(.A(n2302), .B(n2791), .C(n2249), .D(n3512), .Y(n2381));
MX2X1    g1674(.A(g1747), .B(g1781), .S0(n2292), .Y(n2386));
NOR3X1   g1675(.A(n2302), .B(n2791), .C(n2249), .Y(n3515));
XOR2X1   g1676(.A(n3449), .B(g802), .Y(n3516));
AND2X1   g1677(.A(n3516), .B(n3515), .Y(n2391));
MX2X1    g1678(.A(g158), .B(g275), .S0(n2670), .Y(n2396));
MX2X1    g1679(.A(g1508), .B(g1524), .S0(n2509), .Y(n2401));
MX2X1    g1680(.A(g1419), .B(g1577), .S0(n2574), .Y(n2406));
XOR2X1   g1681(.A(n2796), .B(n2795), .Y(n3521));
AND2X1   g1682(.A(n3521), .B(n3515), .Y(n2411));
AND2X1   g1683(.A(g391), .B(g109), .Y(n3523));
MX2X1    g1684(.A(g386), .B(n3523), .S0(n2413), .Y(n2416));
NOR2X1   g1685(.A(n2445_1), .B(g664), .Y(n3525));
XOR2X1   g1686(.A(n3525), .B(g658), .Y(n3526));
MX2X1    g1687(.A(n3498), .B(n3526), .S0(n2446), .Y(n3527));
OAI21X1  g1688(.A0(n3527), .A1(n2473), .B0(n2478), .Y(n2421));
AND2X1   g1689(.A(g186), .B(g109), .Y(n2426));
OR2X1    g1690(.A(n2871), .B(n1919_1), .Y(n2436));
AND2X1   g1691(.A(g1125), .B(g109), .Y(n2440));
NOR4X1   g1692(.A(g1383), .B(g219), .C(g186), .D(g1386), .Y(n3532));
NOR4X1   g1693(.A(g213), .B(g1377), .C(g207), .D(g1380), .Y(n3533));
AND2X1   g1694(.A(n3533), .B(n3532), .Y(n3534));
INVX1    g1695(.A(n3534), .Y(n3535));
NOR4X1   g1696(.A(g225), .B(g1371), .C(g243), .D(g1368), .Y(n3536));
NOR4X1   g1697(.A(g231), .B(g1365), .C(g1362), .D(g237), .Y(n3537));
AND2X1   g1698(.A(n3537), .B(n3536), .Y(n3538));
INVX1    g1699(.A(n3538), .Y(n3539));
OR4X1    g1700(.A(g192), .B(g1400), .C(g248), .D(g1374), .Y(n3540));
OR4X1    g1701(.A(g201), .B(g1397), .C(g1389), .D(g197), .Y(n3541));
NOR4X1   g1702(.A(n3540), .B(n3539), .C(n3535), .D(n3541), .Y(n3542));
XOR2X1   g1703(.A(g1386), .B(g1389), .Y(n3543));
XOR2X1   g1704(.A(n3543), .B(g197), .Y(n3544));
XOR2X1   g1705(.A(n3544), .B(n2923), .Y(n3545));
XOR2X1   g1706(.A(n3545), .B(n3542), .Y(n3546));
NOR2X1   g1707(.A(n3546), .B(n2249), .Y(n2445));
AND2X1   g1708(.A(g1280), .B(g109), .Y(n3548));
MX2X1    g1709(.A(g1284), .B(n3548), .S0(n2601), .Y(n2450));
MX2X1    g1710(.A(g1083), .B(g351), .S0(n2572), .Y(n2455));
AND2X1   g1711(.A(n2734), .B(n2433), .Y(n3551));
NOR2X1   g1712(.A(g643), .B(g646), .Y(n3552));
XOR2X1   g1713(.A(n3552), .B(g650), .Y(n3553));
MX2X1    g1714(.A(g650), .B(n3553), .S0(g627), .Y(n3554));
AND2X1   g1715(.A(n3554), .B(n3551), .Y(n2460));
MX2X1    g1716(.A(g1636), .B(n2635), .S0(n2485_1), .Y(n2465));
AND2X1   g1717(.A(g421), .B(g109), .Y(n3557));
MX2X1    g1718(.A(g416), .B(n3557), .S0(n2413), .Y(n2475));
NOR2X1   g1719(.A(g590), .B(n2249), .Y(n3559));
XOR2X1   g1720(.A(g762), .B(g758), .Y(n3560));
AND2X1   g1721(.A(n3560), .B(n3559), .Y(n2480));
MX2X1    g1722(.A(g956), .B(g845), .S0(n2816), .Y(n2485));
XOR2X1   g1723(.A(n2530_1), .B(g378), .Y(n3563));
MX2X1    g1724(.A(g378), .B(n3563), .S0(n2580_1), .Y(n3564));
AND2X1   g1725(.A(n3564), .B(n2582), .Y(n2490));
MX2X1    g1726(.A(g1756), .B(g1796), .S0(n2292), .Y(n2495));
MX2X1    g1727(.A(g1035), .B(g1068), .S0(n2485_1), .Y(n3567));
MX2X1    g1728(.A(g1027), .B(n3567), .S0(n2485_1), .Y(n2510));
MX2X1    g1729(.A(g1053), .B(g1086), .S0(n2485_1), .Y(n3569));
MX2X1    g1730(.A(g1003), .B(n3569), .S0(n2485_1), .Y(n2515));
INVX1    g1731(.A(g1432), .Y(n3571));
XOR2X1   g1732(.A(n3486), .B(n3571), .Y(n3572));
NOR2X1   g1733(.A(n3572), .B(n2249), .Y(n2520));
AND2X1   g1734(.A(g1145), .B(g109), .Y(n2525));
NOR3X1   g1735(.A(n2672), .B(g1216), .C(n2249), .Y(n2530));
XOR2X1   g1736(.A(g1223), .B(g1218), .Y(n3576));
MX2X1    g1737(.A(n3576), .B(g1223), .S0(n2846), .Y(n3577));
AND2X1   g1738(.A(n3577), .B(n2844), .Y(n2535));
AND2X1   g1739(.A(g406), .B(g109), .Y(n3579));
MX2X1    g1740(.A(g401), .B(n3579), .S0(n2413), .Y(n2540));
NOR4X1   g1741(.A(n2260), .B(n2393), .C(n2483), .D(n2406_1), .Y(n3581));
NAND4X1  g1742(.A(n2872_1), .B(n3005), .C(g109), .D(n3581), .Y(n3582));
MX2X1    g1743(.A(g1811), .B(n3582), .S0(n2708_1), .Y(n2545));
INVX1    g1744(.A(g1642), .Y(n3584));
AOI21X1  g1745(.A0(n2571), .A1(g1696), .B0(n3584), .Y(n2550));
MX2X1    g1746(.A(g87), .B(g1047), .S0(g85), .Y(n2555));
AOI21X1  g1747(.A0(n1983), .A1(g109), .B0(n2591), .Y(n3587));
AND2X1   g1748(.A(n2990), .B(n2592), .Y(n3588));
OR2X1    g1749(.A(n3588), .B(n3587), .Y(n3589));
MX2X1    g1750(.A(g1654), .B(n3589), .S0(n2572), .Y(n2560));
AND2X1   g1751(.A(g1374), .B(g109), .Y(n2565));
MX2X1    g1752(.A(g1432), .B(g1595), .S0(n2574), .Y(n2570));
MX2X1    g1753(.A(g1490), .B(g1537), .S0(n2509), .Y(n2575));
NOR2X1   g1754(.A(n2462), .B(n3253), .Y(n3594));
MX2X1    g1755(.A(n3594), .B(g718), .S0(n2567), .Y(n2580));
MX2X1    g1756(.A(g1056), .B(g1089), .S0(n2485_1), .Y(n3596));
MX2X1    g1757(.A(g999), .B(n3596), .S0(n2485_1), .Y(n2585));
XOR2X1   g1758(.A(g798), .B(g794), .Y(n3598));
OR4X1    g1759(.A(n2302), .B(n2791), .C(n2249), .D(n3598), .Y(n2590));
INVX1    g1760(.A(n3210), .Y(n3600));
AND2X1   g1761(.A(g481), .B(g109), .Y(n3601));
MX2X1    g1762(.A(n3600), .B(n3601), .S0(n2413), .Y(n2595));
OAI21X1  g1763(.A0(g754), .A1(g750), .B0(g746), .Y(n3603));
AOI21X1  g1764(.A0(g754), .A1(g750), .B0(n3603), .Y(n2600));
MX2X1    g1765(.A(g1801), .B(g1330), .S0(n2907_1), .Y(n2605));
XOR2X1   g1766(.A(n3222), .B(g790), .Y(n3606));
AND2X1   g1767(.A(n3606), .B(n3559), .Y(n2615));
NOR4X1   g1768(.A(n2632), .B(g1101), .C(n2620_1), .D(g1107), .Y(n3608));
XOR2X1   g1769(.A(n3608), .B(g1113), .Y(n3609));
MX2X1    g1770(.A(g1512), .B(n3609), .S0(n2485_1), .Y(n2620));
XOR2X1   g1771(.A(n2802_1), .B(g1486), .Y(n3611));
AND2X1   g1772(.A(n3611), .B(g109), .Y(n2629));
AND2X1   g1773(.A(g1166), .B(g109), .Y(n2634));
MX2X1    g1774(.A(g90), .B(g1056), .S0(g85), .Y(n2639));
OAI21X1  g1775(.A0(g754), .A1(n2680), .B0(g348), .Y(n3615));
OAI21X1  g1776(.A0(n3196), .A1(n2682), .B0(n3615), .Y(n2644));
AND2X1   g1777(.A(g1260), .B(g109), .Y(n3617));
MX2X1    g1778(.A(g1255), .B(n3617), .S0(n2601), .Y(n2653));
XOR2X1   g1779(.A(n1561), .B(g135), .Y(n3619));
AND2X1   g1780(.A(n3619), .B(g109), .Y(n2663));
MX2X1    g1781(.A(g560), .B(g219), .S0(g18), .Y(n2673));
AND2X1   g1782(.A(g521), .B(g109), .Y(n3622));
MX2X1    g1783(.A(g525), .B(n3622), .S0(n2413), .Y(n2678));
MX2X1    g1784(.A(g1781), .B(g1318), .S0(n2907_1), .Y(n2683));
INVX1    g1785(.A(g1872), .Y(n3625));
NOR2X1   g1786(.A(n2319), .B(g1878), .Y(n3626));
XOR2X1   g1787(.A(n3626), .B(g1872), .Y(n3627));
MX2X1    g1788(.A(n3625), .B(n3627), .S0(n2320), .Y(n3628));
OAI21X1  g1789(.A0(n3628), .A1(n2342), .B0(n2348), .Y(n2688));
INVX1    g1790(.A(g677), .Y(n3630));
NAND2X1  g1791(.A(g658), .B(g668), .Y(n3631));
MX2X1    g1792(.A(n3631), .B(n3338), .S0(n2454), .Y(n3632));
MX2X1    g1793(.A(n2713_1), .B(n3632), .S0(n2445_1), .Y(n3633));
XOR2X1   g1794(.A(n3633), .B(g677), .Y(n3634));
MX2X1    g1795(.A(n3630), .B(n3634), .S0(n2446), .Y(n3635));
OAI21X1  g1796(.A0(n3635), .A1(n2473), .B0(n2478), .Y(n2693));
NOR4X1   g1797(.A(n2923), .B(g192), .C(g1397), .D(g1374), .Y(n3637));
NOR4X1   g1798(.A(g1400), .B(g248), .C(g1389), .D(g197), .Y(n3638));
NAND4X1  g1799(.A(n3637), .B(n3538), .C(n3534), .D(n3638), .Y(n3639));
NOR2X1   g1800(.A(n3639), .B(n2249), .Y(n2703));
MX2X1    g1801(.A(g1474), .B(g1549), .S0(n2509), .Y(n2708));
MX2X1    g1802(.A(g947), .B(g833), .S0(n2816), .Y(n2713));
OAI22X1  g1803(.A0(n3283), .A1(n2341_1), .B0(n2765), .B1(n2315), .Y(n3643));
XOR2X1   g1804(.A(n3643), .B(n2316_1), .Y(n3644));
NOR2X1   g1805(.A(n3644), .B(n2630), .Y(n2718));
MX2X1    g1806(.A(g1436), .B(g1598), .S0(n2574), .Y(n2723));
AND2X1   g1807(.A(g1121), .B(g109), .Y(n2728));
MX2X1    g1808(.A(g1786), .B(g1321), .S0(n2907_1), .Y(n2733));
AND2X1   g1809(.A(g506), .B(g109), .Y(n3649));
MX2X1    g1810(.A(g501), .B(n3649), .S0(n2413), .Y(n2738));
MX2X1    g1811(.A(g546), .B(n2595_1), .S0(n2485_1), .Y(n2743));
INVX1    g1812(.A(n2335), .Y(n3652));
MX2X1    g1813(.A(n3652), .B(n2338), .S0(n2326_1), .Y(n3653));
MX2X1    g1814(.A(n3075), .B(n3653), .S0(n2319), .Y(n3654));
XOR2X1   g1815(.A(n3654), .B(g1909), .Y(n3655));
MX2X1    g1816(.A(n2334), .B(n3655), .S0(n2320), .Y(n3656));
OAI21X1  g1817(.A0(n3656), .A1(n2342), .B0(n2348), .Y(n2748));
MX2X1    g1818(.A(g1470), .B(g1552), .S0(n2509), .Y(n2757));
OAI21X1  g1819(.A0(g1703), .A1(g1696), .B0(g1687), .Y(n3659));
NAND2X1  g1820(.A(n3659), .B(n3263), .Y(n2767));
MX2X1    g1821(.A(g1407), .B(g1586), .S0(n2574), .Y(n2772));
AND2X1   g1822(.A(g1141), .B(g109), .Y(n2782));
ZERO     g1823(.Y(n2787));
XOR2X1   g1824(.A(g1341), .B(n2029), .Y(n3664));
MX2X1    g1825(.A(n2081), .B(n3664), .S0(n2121), .Y(n3665));
NOR2X1   g1826(.A(n3665), .B(n3052_1), .Y(n2792));
INVX1    g1827(.A(g1645), .Y(n3667));
AOI21X1  g1828(.A0(n2571), .A1(g1696), .B0(n3667), .Y(n2802));
NAND2X1  g1829(.A(g1394), .B(g109), .Y(n3669));
NOR2X1   g1830(.A(n3669), .B(n3639), .Y(n2807));
XOR2X1   g1831(.A(n1680), .B(g139), .Y(n3671));
AND2X1   g1832(.A(n3671), .B(g109), .Y(n2812));
AND2X1   g1833(.A(g525), .B(g109), .Y(n3673));
MX2X1    g1834(.A(g530), .B(n3673), .S0(n2413), .Y(n2817));
MX2X1    g1835(.A(g1448), .B(g1607), .S0(n2574), .Y(n2827));
OR2X1    g1836(.A(n2681), .B(g67), .Y(n2837));
AND2X1   g1837(.A(g1275), .B(g109), .Y(n3677));
MX2X1    g1838(.A(n2889), .B(n3677), .S0(n2601), .Y(n2842));
MX2X1    g1839(.A(g1771), .B(g1311), .S0(n2907_1), .Y(n2847));
MX2X1    g1840(.A(g1615), .B(n2824), .S0(n2485_1), .Y(n2852));
AOI21X1  g1841(.A0(n2531), .A1(n2949), .B0(g382), .Y(n3681));
NOR3X1   g1842(.A(n3681), .B(g869), .C(n2249), .Y(n2857));
AND2X1   g1843(.A(g201), .B(g109), .Y(n2862));
MX2X1    g1844(.A(g178), .B(g266), .S0(n2670), .Y(n2867));
AND2X1   g1845(.A(g1284), .B(g109), .Y(n3685));
MX2X1    g1846(.A(g1292), .B(n3685), .S0(n2601), .Y(n2872));
AND2X1   g1847(.A(g213), .B(g109), .Y(n2877));
NOR2X1   g1848(.A(n2462), .B(n3497), .Y(n3688));
MX2X1    g1849(.A(n3688), .B(g664), .S0(n2567), .Y(n2882));
AND2X1   g1850(.A(n2852_1), .B(g1850), .Y(n2887));
XOR2X1   g1851(.A(n2673), .B(n2422), .Y(n3691));
NOR2X1   g1852(.A(n3691), .B(n2249), .Y(n2892));
AND2X1   g1853(.A(g411), .B(g109), .Y(n3693));
MX2X1    g1854(.A(g406), .B(n3693), .S0(n2413), .Y(n2897));
AND2X1   g1855(.A(g431), .B(g109), .Y(n3695));
MX2X1    g1856(.A(g435), .B(n3695), .S0(n2413), .Y(n2902));
NOR2X1   g1857(.A(n2331_1), .B(n3377), .Y(n3697));
MX2X1    g1858(.A(n3697), .B(g1896), .S0(n2766), .Y(n2907));
AND2X1   g1859(.A(g1419), .B(g109), .Y(n2912));
MX2X1    g1860(.A(g1630), .B(n2675), .S0(n2485_1), .Y(n2917));
OR2X1    g1861(.A(n2681), .B(g49), .Y(n2922));
MX2X1    g1862(.A(g1050), .B(g1083), .S0(n2485_1), .Y(n3702));
MX2X1    g1863(.A(g991), .B(n3702), .S0(n2485_1), .Y(n2927));
AND2X1   g1864(.A(g1300), .B(g109), .Y(n3704));
MX2X1    g1865(.A(g1304), .B(n3704), .S0(n2601), .Y(n2932));
OAI21X1  g1866(.A0(g754), .A1(n2680), .B0(g339), .Y(n3706));
OAI21X1  g1867(.A0(n3177), .A1(n2682), .B0(n3706), .Y(n2937));
MX2X1    g1868(.A(g1750), .B(g1786), .S0(n2292), .Y(n2947));
INVX1    g1869(.A(g1444), .Y(n3709));
XOR2X1   g1870(.A(n3056), .B(n3709), .Y(n3710));
NOR2X1   g1871(.A(n3710), .B(n2249), .Y(n2957));
MX2X1    g1872(.A(g1666), .B(n2647), .S0(n2572), .Y(n2962));
MX2X1    g1873(.A(g1504), .B(g1528), .S0(n2509), .Y(n2967));
XOR2X1   g1874(.A(n3368), .B(g1351), .Y(n3714));
MX2X1    g1875(.A(n2167), .B(n3714), .S0(n2121), .Y(n3715));
NOR2X1   g1876(.A(n3715), .B(n3052_1), .Y(n2972));
INVX1    g1877(.A(g1648), .Y(n3717));
AOI21X1  g1878(.A0(n2571), .A1(g1696), .B0(n3717), .Y(n2977));
XOR2X1   g1879(.A(n1670), .B(n2420), .Y(n3719));
NOR2X1   g1880(.A(n3719), .B(n2249), .Y(n2982));
NOR4X1   g1881(.A(g1110), .B(n2631), .C(g1104), .D(g1107), .Y(n3721));
NOR4X1   g1882(.A(g1145), .B(g1137), .C(g1133), .D(g1141), .Y(n3722));
NOR4X1   g1883(.A(g1125), .B(g1129), .C(g1117), .D(g1121), .Y(n3723));
NOR3X1   g1884(.A(g1160), .B(g1157), .C(g1153), .Y(n3724));
NOR4X1   g1885(.A(g1166), .B(g1149), .C(g1163), .D(g1113), .Y(n3725));
NAND4X1  g1886(.A(n3724), .B(n3723), .C(n3722), .D(n3725), .Y(n3726));
INVX1    g1887(.A(g1153), .Y(n3727));
XOR2X1   g1888(.A(g1149), .B(n3727), .Y(n3728));
AND2X1   g1889(.A(n3728), .B(n3726), .Y(n3729));
XOR2X1   g1890(.A(n3729), .B(n3721), .Y(n3730));
XOR2X1   g1891(.A(n3730), .B(n2931), .Y(n3731));
XOR2X1   g1892(.A(n3731), .B(n3359), .Y(n3732));
MX2X1    g1893(.A(g1618), .B(n3732), .S0(n2485_1), .Y(n2987));
AND2X1   g1894(.A(g1235), .B(g109), .Y(n3734));
MX2X1    g1895(.A(g1275), .B(n3734), .S0(n2601), .Y(n2992));
MX2X1    g1896(.A(g166), .B(g299), .S0(n2670), .Y(n2997));
AND2X1   g1897(.A(g435), .B(g109), .Y(n3737));
MX2X1    g1898(.A(g440), .B(n3737), .S0(n2413), .Y(n3002));
AND2X1   g1899(.A(n2682), .B(g64), .Y(n3007));
MX2X1    g1900(.A(g1466), .B(g1555), .S0(n2509), .Y(n3012));
MX2X1    g1901(.A(g1047), .B(g1080), .S0(n2485_1), .Y(n3741));
MX2X1    g1902(.A(g995), .B(n3741), .S0(n2485_1), .Y(n3017));
MX2X1    g1903(.A(g1621), .B(n2863), .S0(n2485_1), .Y(n3022));
AND2X1   g1904(.A(g1113), .B(g109), .Y(n3027));
XOR2X1   g1905(.A(g643), .B(n3387), .Y(n3745));
NAND3X1  g1906(.A(n3745), .B(n2734), .C(n2433), .Y(n3032));
XOR2X1   g1907(.A(n2685), .B(g1490), .Y(n3747));
AND2X1   g1908(.A(n3747), .B(g109), .Y(n3037));
MX2X1    g1909(.A(g1415), .B(g1567), .S0(n2574), .Y(n3042));
NOR2X1   g1910(.A(n2462), .B(n3337), .Y(n3750));
MX2X1    g1911(.A(n3750), .B(g682), .S0(n2567), .Y(n3047));
AND2X1   g1912(.A(g534), .B(g109), .Y(n3752));
MX2X1    g1913(.A(g538), .B(n3752), .S0(n2413), .Y(n3052));
AND2X1   g1914(.A(g1771), .B(g1766), .Y(n3754));
XOR2X1   g1915(.A(n3754), .B(n2482), .Y(n3755));
MX2X1    g1916(.A(n2482), .B(n3755), .S0(n2708_1), .Y(n3756));
NOR2X1   g1917(.A(n3756), .B(g1713), .Y(n3057));
MX2X1    g1918(.A(g569), .B(n3589), .S0(n2485_1), .Y(n3062));
AND2X1   g1919(.A(g1160), .B(g109), .Y(n3067));
OR2X1    g1920(.A(n3424), .B(n1962_1), .Y(n3072));
MX2X1    g1921(.A(g88), .B(g1050), .S0(g85), .Y(n3076));
INVX1    g1922(.A(g1), .Y(n3762));
NAND4X1  g1923(.A(g1515), .B(g1520), .C(g1436), .D(g1440), .Y(n3763));
NOR3X1   g1924(.A(n3763), .B(g1411), .C(g1415), .Y(n3764));
NOR4X1   g1925(.A(n3571), .B(n2821), .C(g1407), .D(g1403), .Y(n3765));
NAND2X1  g1926(.A(g1419), .B(g1424), .Y(n3766));
NOR3X1   g1927(.A(n3766), .B(n2629_1), .C(n3709), .Y(n3767));
NAND4X1  g1928(.A(n3765), .B(n3764), .C(n2508), .D(n3767), .Y(n3768));
AOI21X1  g1929(.A0(n3768), .A1(n3762), .B0(n2249), .Y(n3081));
AND2X1   g1930(.A(g511), .B(g109), .Y(n3770));
MX2X1    g1931(.A(g506), .B(n3770), .S0(n2413), .Y(n3086));
MX2X1    g1932(.A(g1724), .B(n2406_1), .S0(n2785), .Y(n3091));
AOI21X1  g1933(.A0(g115), .A1(g18), .B0(g12), .Y(n3773));
NOR2X1   g1934(.A(n3773), .B(n2249), .Y(n3096));
MX2X1    g1935(.A(g1878), .B(g1950), .S0(n2766), .Y(n3775));
OR2X1    g1936(.A(n3775), .B(n2331_1), .Y(n3101));
OR2X1    g1937(.A(n2681), .B(g73), .Y(n3106));
BUFX1    g1938(.A(g18), .Y(g2355));
BUFX1    g1939(.A(g578), .Y(g2601));
BUFX1    g1940(.A(g587), .Y(g2602));
BUFX1    g1941(.A(g588), .Y(g2603));
BUFX1    g1942(.A(g589), .Y(g2604));
BUFX1    g1943(.A(g579), .Y(g2605));
BUFX1    g1944(.A(g580), .Y(g2606));
BUFX1    g1945(.A(g581), .Y(g2607));
BUFX1    g1946(.A(g582), .Y(g2608));
BUFX1    g1947(.A(g583), .Y(g2609));
BUFX1    g1948(.A(g584), .Y(g2610));
BUFX1    g1949(.A(g585), .Y(g2611));
BUFX1    g1950(.A(g586), .Y(g2612));
BUFX1    g1951(.A(g865), .Y(g2648));
BUFX1    g1952(.A(g883), .Y(g2986));
BUFX1    g1953(.A(g878), .Y(g3007));
BUFX1    g1954(.A(g1206), .Y(g3069));
BUFX1    g1955(.A(g754), .Y(g4172));
BUFX1    g1956(.A(g758), .Y(g4173));
BUFX1    g1957(.A(g762), .Y(g4174));
BUFX1    g1958(.A(g766), .Y(g4175));
BUFX1    g1959(.A(g770), .Y(g4176));
BUFX1    g1960(.A(g774), .Y(g4177));
BUFX1    g1961(.A(g778), .Y(g4178));
BUFX1    g1962(.A(g782), .Y(g4179));
BUFX1    g1963(.A(g786), .Y(g4180));
BUFX1    g1964(.A(g790), .Y(g4181));
BUFX1    g1965(.A(g1961), .Y(g4887));
BUFX1    g1966(.A(g1960), .Y(g4888));
BUFX1    g1967(.A(g872), .Y(g5101));
BUFX1    g1968(.A(g873), .Y(g5105));
BUFX1    g1969(.A(g27), .Y(g7744));
BUFX1    g1970(.A(g872), .Y(g8061));
BUFX1    g1971(.A(g873), .Y(g8062));
INVX1    g1972(.A(g1810), .Y(g8271));
MX2X1    g1973(.A(g1654), .B(g1672), .S0(g1690), .Y(g8561));
MX2X1    g1974(.A(g1657), .B(g1675), .S0(g1690), .Y(g8562));
MX2X1    g1975(.A(g1660), .B(g1678), .S0(g1690), .Y(g8563));
MX2X1    g1976(.A(g1663), .B(g1681), .S0(g1690), .Y(g8564));
MX2X1    g1977(.A(g1666), .B(g1684), .S0(g1690), .Y(g8565));
MX2X1    g1978(.A(g1669), .B(g1687), .S0(g1690), .Y(g8566));
BUFX1    g1979(.A(g85), .Y(g6267));
BUFX1    g1980(.A(g42), .Y(g6257));
BUFX1    g1981(.A(g102), .Y(g6282));
BUFX1    g1982(.A(g104), .Y(g6284));
BUFX1    g1983(.A(g101), .Y(g6281));
BUFX1    g1984(.A(g29), .Y(g6253));
BUFX1    g1985(.A(g28), .Y(g6285));
BUFX1    g1986(.A(g103), .Y(g6283));
BUFX1    g1987(.A(g83), .Y(g6265));
BUFX1    g1988(.A(g87), .Y(g6269));
BUFX1    g1989(.A(g922), .Y(g4204));
BUFX1    g1990(.A(g892), .Y(g4193));
BUFX1    g1991(.A(g84), .Y(g6266));
BUFX1    g1992(.A(g919), .Y(g4203));
BUFX1    g1993(.A(g1182), .Y(g4212));
BUFX1    g1994(.A(g925), .Y(g4196));
BUFX1    g1995(.A(g48), .Y(g6263));
BUFX1    g1996(.A(g895), .Y(g4194));
BUFX1    g1997(.A(g889), .Y(g4192));
BUFX1    g1998(.A(g1185), .Y(g4213));
BUFX1    g1999(.A(g41), .Y(g6256));
BUFX1    g2000(.A(g43), .Y(g6258));
BUFX1    g2001(.A(g99), .Y(g6279));
BUFX1    g2002(.A(g1173), .Y(g4209));
BUFX1    g2003(.A(g1203), .Y(g4208));
BUFX1    g2004(.A(g1188), .Y(g4214));
BUFX1    g2005(.A(g1197), .Y(g4206));
BUFX1    g2006(.A(g46), .Y(g6261));
BUFX1    g2007(.A(g31), .Y(g6255));
BUFX1    g2008(.A(g45), .Y(g6260));
BUFX1    g2009(.A(g92), .Y(g6274));
BUFX1    g2010(.A(g89), .Y(g6271));
BUFX1    g2011(.A(g898), .Y(g4195));
BUFX1    g2012(.A(g91), .Y(g6273));
BUFX1    g2013(.A(g93), .Y(g6275));
BUFX1    g2014(.A(g913), .Y(g4201));
BUFX1    g2015(.A(g82), .Y(g6264));
BUFX1    g2016(.A(g88), .Y(g6270));
BUFX1    g2017(.A(g1194), .Y(g4216));
BUFX1    g2018(.A(g47), .Y(g6262));
BUFX1    g2019(.A(g96), .Y(g6278));
BUFX1    g2020(.A(g910), .Y(g4200));
BUFX1    g2021(.A(g95), .Y(g6277));
BUFX1    g2022(.A(g904), .Y(g4198));
BUFX1    g2023(.A(g1176), .Y(g4210));
BUFX1    g2024(.A(g901), .Y(g4197));
BUFX1    g2025(.A(g44), .Y(g6259));
BUFX1    g2026(.A(g916), .Y(g4202));
BUFX1    g2027(.A(g100), .Y(g6280));
BUFX1    g2028(.A(g886), .Y(g4191));
BUFX1    g2029(.A(g30), .Y(g6254));
BUFX1    g2030(.A(g86), .Y(g6268));
BUFX1    g2031(.A(g1170), .Y(g4205));
BUFX1    g2032(.A(g1200), .Y(g4207));
BUFX1    g2033(.A(g1191), .Y(g4215));
BUFX1    g2034(.A(g907), .Y(g4199));
BUFX1    g2035(.A(g90), .Y(g6272));
BUFX1    g2036(.A(g94), .Y(g6276));
BUFX1    g2037(.A(g1179), .Y(g4211));
BUFX1    g2038(.A(g255), .Y(n465));
BUFX1    g2039(.A(g1736), .Y(n579));
BUFX1    g2040(.A(g256), .Y(n659));
BUFX1    g2041(.A(g1713), .Y(n724));
BUFX1    g2042(.A(g794), .Y(n729));
BUFX1    g2043(.A(g104), .Y(n764));
BUFX1    g2044(.A(g260), .Y(n779));
BUFX1    g2045(.A(g1955), .Y(n794));
BUFX1    g2046(.A(g1956), .Y(g1957));
BUFX1    g2047(.A(g746), .Y(n897));
BUFX1    g2048(.A(g878), .Y(n916));
BUFX1    g2049(.A(g29), .Y(n951));
BUFX1    g2050(.A(g883), .Y(n1056));
BUFX1    g2051(.A(g1360), .Y(n1081));
BUFX1    g2052(.A(g102), .Y(n1096));
BUFX1    g2053(.A(g28), .Y(n1201));
BUFX1    g2054(.A(g103), .Y(n1221));
BUFX1    g2055(.A(g755), .Y(n1231));
BUFX1    g2056(.A(g262), .Y(n1326));
BUFX1    g2057(.A(g254), .Y(n1366));
BUFX1    g2058(.A(g103), .Y(n1386));
BUFX1    g2059(.A(g875), .Y(n1391));
BUFX1    g2060(.A(g1206), .Y(n1421));
BUFX1    g2061(.A(g1356), .Y(n1526));
BUFX1    g2062(.A(g257), .Y(n1576));
BUFX1    g2063(.A(g1958), .Y(n1615));
BUFX1    g2064(.A(g261), .Y(n1645));
BUFX1    g2065(.A(g826), .Y(n1690));
BUFX1    g2066(.A(g253), .Y(n1775));
BUFX1    g2067(.A(g636), .Y(n1785));
BUFX1    g2068(.A(g83), .Y(n1924));
BUFX1    g2069(.A(g1217), .Y(n1942));
BUFX1    g2070(.A(g756), .Y(n1967));
BUFX1    g2071(.A(g802), .Y(n1992));
BUFX1    g2072(.A(g798), .Y(n2136));
BUFX1    g2073(.A(g814), .Y(n2161));
BUFX1    g2074(.A(g822), .Y(n2281));
BUFX1    g2075(.A(g101), .Y(n2331));
BUFX1    g2076(.A(g818), .Y(n2470));
BUFX1    g2077(.A(g29), .Y(n2500));
BUFX1    g2078(.A(g806), .Y(n2505));
BUFX1    g2079(.A(g810), .Y(n2610));
BUFX1    g2080(.A(g113), .Y(n2624));
BUFX1    g2081(.A(g874), .Y(n2648));
BUFX1    g2082(.A(g1854), .Y(n2668));
BUFX1    g2083(.A(g28), .Y(n2698));
BUFX1    g2084(.A(g83), .Y(n2753));
BUFX1    g2085(.A(g101), .Y(n2762));
BUFX1    g2086(.A(g259), .Y(n2777));
BUFX1    g2087(.A(g104), .Y(n2822));
BUFX1    g2088(.A(g258), .Y(n2832));
BUFX1    g2089(.A(g102), .Y(n2952));
endmodule
