//Converted to Combinational (Partial output: n3334) , Module name: s38584_n3334 , Timestamp: 2018-12-03T15:51:16.986606 
module s38584_n3334 ( g35, g3614, g3684, g4871, g4983, g4991, g4975, g4966, g4849, g4859, g4843, g4944, g4899, g3654, g3618, g3639, g3610, g3558, g3680, g3562, g3602, g3570, g3632, g3703, g3554, g3625, g3542, g3689, g3574, g3668, g3649, g3550, g3582, g3566, g3598, g3676, g3538, g3672, g3590, g3606, g3546, g3578, g3661, g3594, g3586, n3334 );
input g35, g3614, g3684, g4871, g4983, g4991, g4975, g4966, g4849, g4859, g4843, g4944, g4899, g3654, g3618, g3639, g3610, g3558, g3680, g3562, g3602, g3570, g3632, g3703, g3554, g3625, g3542, g3689, g3574, g3668, g3649, g3550, g3582, g3566, g3598, g3676, g3538, g3672, g3590, g3606, g3546, g3578, g3661, g3594, g3586;
output n3334;
wire n8049, n5930, n5974, n5927, n5928, n5929_1, n5973, n5941, n5956, n5963, n4963, n4960, n4892, n4893, n5965, n5968, n5972_1, n5935, n5940, n5949_1, n5952, n5955, n5962_1, n5957, n5959, n5964, n5966, n5938, n5967_1, n5969, n5970, n5971, n5932, n5933, n5934_1, n5936, n5939_1, n5948, n5943, n5944_1, n5946, n5950, n5951, n5953, n5954_1, n5960, n5961, n5805, n5176_1, n5958_1, n5937, n5945, n5931, n5947, n5942;
MX2X1    g3403(.A(g3614), .B(n8049), .S0(g35), .Y(n3334));
MX2X1    g3402(.A(g3684), .B(n5974), .S0(n5930), .Y(n8049));
AOI21X1  g1290(.A0(n5929_1), .A1(n5928), .B0(n5927), .Y(n5930));
NAND4X1  g1334(.A(n5963), .B(n5956), .C(n5941), .D(n5973), .Y(n5974));
INVX1    g1287(.A(g4871), .Y(n5927));
NOR3X1   g1288(.A(n4963), .B(g4991), .C(g4983), .Y(n5928));
NOR4X1   g1289(.A(g4975), .B(n4893), .C(n4892), .D(n4960), .Y(n5929_1));
NOR3X1   g1333(.A(n5972_1), .B(n5968), .C(n5965), .Y(n5973));
NOR2X1   g1301(.A(n5940), .B(n5935), .Y(n5941));
NOR3X1   g1316(.A(n5955), .B(n5952), .C(n5949_1), .Y(n5956));
AOI21X1  g1323(.A0(n5959), .A1(n5957), .B0(n5962_1), .Y(n5963));
INVX1    g0343(.A(g4966), .Y(n4963));
NAND3X1  g0340(.A(g4843), .B(g4859), .C(g4849), .Y(n4960));
INVX1    g0272(.A(g4944), .Y(n4892));
INVX1    g0273(.A(g4899), .Y(n4893));
NOR2X1   g1325(.A(n5964), .B(n5957), .Y(n5965));
OAI21X1  g1328(.A0(n5967_1), .A1(n5938), .B0(n5966), .Y(n5968));
AOI21X1  g1332(.A0(n5971), .A1(n5970), .B0(n5969), .Y(n5972_1));
AOI21X1  g1295(.A0(n5934_1), .A1(n5933), .B0(n5932), .Y(n5935));
OAI21X1  g1300(.A0(n5939_1), .A1(n5938), .B0(n5936), .Y(n5940));
NAND4X1  g1309(.A(n5946), .B(n5944_1), .C(n5943), .D(n5948), .Y(n5949_1));
OAI21X1  g1312(.A0(n5951), .A1(n5932), .B0(n5950), .Y(n5952));
NAND2X1  g1315(.A(n5954_1), .B(n5953), .Y(n5955));
AOI21X1  g1322(.A0(n5961), .A1(n5960), .B0(n5957), .Y(n5962_1));
XOR2X1   g1317(.A(g3654), .B(n5805), .Y(n5957));
AND2X1   g1319(.A(n5958_1), .B(n5176_1), .Y(n5959));
NAND4X1  g1324(.A(g3610), .B(g3639), .C(g3618), .D(n5937), .Y(n5964));
NAND4X1  g1326(.A(g3654), .B(n5805), .C(g3558), .D(n5176_1), .Y(n5966));
NAND2X1  g1298(.A(n5937), .B(g3639), .Y(n5938));
NAND3X1  g1327(.A(g3562), .B(n5805), .C(g3680), .Y(n5967_1));
INVX1    g1329(.A(n5957), .Y(n5969));
NAND3X1  g1330(.A(n5945), .B(g3602), .C(g3618), .Y(n5970));
NAND4X1  g1331(.A(g3639), .B(g3632), .C(g3570), .D(n5937), .Y(n5971));
NAND2X1  g1292(.A(g3703), .B(n5931), .Y(n5932));
NAND3X1  g1293(.A(n5805), .B(g3625), .C(g3554), .Y(n5933));
NAND3X1  g1294(.A(g3654), .B(g3689), .C(g3542), .Y(n5934_1));
NAND4X1  g1296(.A(g3668), .B(n5805), .C(g3574), .D(n5176_1), .Y(n5936));
NAND3X1  g1299(.A(g3550), .B(n5805), .C(g3649), .Y(n5939_1));
NAND4X1  g1308(.A(n5937), .B(g3582), .C(g3639), .D(n5947), .Y(n5948));
NAND4X1  g1303(.A(g3703), .B(n5931), .C(g3566), .D(n5942), .Y(n5943));
NAND4X1  g1304(.A(g3676), .B(g3689), .C(g3598), .D(n5176_1), .Y(n5944_1));
NAND4X1  g1306(.A(g3538), .B(g3689), .C(g3649), .D(n5945), .Y(n5946));
NAND4X1  g1310(.A(g3590), .B(n5805), .C(g3672), .D(n5945), .Y(n5950));
NAND3X1  g1311(.A(g3676), .B(n5805), .C(g3606), .Y(n5951));
NAND4X1  g1313(.A(g3546), .B(g3689), .C(g3680), .D(n5945), .Y(n5953));
NAND4X1  g1314(.A(g3614), .B(g3689), .C(g3625), .D(n5176_1), .Y(n5954_1));
NAND3X1  g1320(.A(n5945), .B(g3578), .C(g3632), .Y(n5960));
NAND4X1  g1321(.A(g3594), .B(g3661), .C(n5931), .D(g3703), .Y(n5961));
INVX1    g1165(.A(g3689), .Y(n5805));
AND2X1   g0543(.A(g3703), .B(g3639), .Y(n5176_1));
AND2X1   g1318(.A(g3661), .B(g3586), .Y(n5958_1));
INVX1    g1297(.A(g3703), .Y(n5937));
NOR2X1   g1305(.A(g3703), .B(g3639), .Y(n5945));
INVX1    g1291(.A(g3639), .Y(n5931));
AND2X1   g1307(.A(g3689), .B(g3672), .Y(n5947));
AND2X1   g1302(.A(g3668), .B(g3689), .Y(n5942));

endmodule
