//Converted to Combinational (Partial output: Z) , Module name: s420_Z
module s420_Z ( Y_1, Y_13, Y_12, Y_11, Y_10, C_1, C_14, Y_14, C_15, Y_15, C_8, Y_8, C_13, C_12, C_11, C_16, Y_16, Y_4, Y_6, Y_5, Y_7, Y_9, C_10, C_9, Y_3, Y_2, X, C_0, C_2, C_7, C_6, C_5, C_4, C_3, Z );
input Y_1, Y_13, Y_12, Y_11, Y_10, C_1, C_14, Y_14, C_15, Y_15, C_8, Y_8, C_13, C_12, C_11, C_16, Y_16, Y_4, Y_6, Y_5, Y_7, Y_9, C_10, C_9, Y_3, Y_2, X, C_0, C_2, C_7, C_6, C_5, C_4, C_3;
output Z;
wire n82, n112, n117, n81, n72, n73_1, n111, n84, n86, n88_1, n113_1, n114, n116, n80, n110, n90, n92, n93_1, n83_1, n85, n87, n115, n79, n74, n75, n76, n109, n95, n97, n99, n89, n91, n78_1, n108_1, n101, n105, n106, n94, n96, n98_1, n77, n107, n100, n104, n102, n103_1;
NAND3X1  g49(.A(n117), .B(n112), .C(n82), .Y(Z));
OR4X1    g13(.A(Y_13), .B(n73_1), .C(n72), .D(n81), .Y(n82));
NOR4X1   g43(.A(n88_1), .B(n86), .C(n84), .D(n111), .Y(n112));
OAI21X1  g48(.A0(n116), .A1(n114), .B0(n113_1), .Y(n117));
OR4X1    g12(.A(Y_10), .B(Y_11), .C(Y_12), .D(n80), .Y(n81));
INVX1    g03(.A(C_14), .Y(n72));
INVX1    g04(.A(Y_14), .Y(n73_1));
NAND4X1  g42(.A(n93_1), .B(n92), .C(n90), .D(n110), .Y(n111));
NOR2X1   g15(.A(n83_1), .B(n81), .Y(n84));
NOR4X1   g17(.A(n80), .B(Y_10), .C(Y_11), .D(n85), .Y(n86));
NOR3X1   g19(.A(n87), .B(n80), .C(Y_10), .Y(n88_1));
NOR3X1   g44(.A(n81), .B(Y_13), .C(Y_14), .Y(n113_1));
AND2X1   g45(.A(Y_15), .B(C_15), .Y(n114));
NOR2X1   g47(.A(n115), .B(Y_15), .Y(n116));
NAND4X1  g11(.A(n76), .B(n75), .C(n74), .D(n79), .Y(n80));
NOR4X1   g41(.A(n99), .B(n97), .C(n95), .D(n109), .Y(n110));
OR2X1    g21(.A(n89), .B(n80), .Y(n90));
NAND4X1  g23(.A(n79), .B(n75), .C(n74), .D(n91), .Y(n92));
NAND4X1  g24(.A(n75), .B(Y_8), .C(C_8), .D(n79), .Y(n93_1));
NAND2X1  g14(.A(Y_13), .B(C_13), .Y(n83_1));
NAND2X1  g16(.A(Y_12), .B(C_12), .Y(n85));
NAND2X1  g18(.A(Y_11), .B(C_11), .Y(n87));
NAND2X1  g46(.A(Y_16), .B(C_16), .Y(n115));
NOR4X1   g10(.A(Y_5), .B(Y_6), .C(Y_4), .D(n78_1), .Y(n79));
INVX1    g05(.A(Y_8), .Y(n74));
INVX1    g06(.A(Y_7), .Y(n75));
INVX1    g07(.A(Y_9), .Y(n76));
NAND4X1  g40(.A(n106), .B(n105), .C(n101), .D(n108_1), .Y(n109));
AND2X1   g26(.A(n94), .B(n79), .Y(n95));
NOR4X1   g28(.A(n78_1), .B(Y_5), .C(Y_4), .D(n96), .Y(n97));
NOR3X1   g30(.A(n98_1), .B(n78_1), .C(Y_4), .Y(n99));
NAND2X1  g20(.A(Y_10), .B(C_10), .Y(n89));
AND2X1   g22(.A(Y_9), .B(C_9), .Y(n91));
OR4X1    g09(.A(Y_2), .B(Y_3), .C(n77), .D(Y_1), .Y(n78_1));
OAI21X1  g39(.A0(n107), .A1(C_0), .B0(X), .Y(n108_1));
OR2X1    g32(.A(n100), .B(n78_1), .Y(n101));
NAND4X1  g36(.A(n103_1), .B(n102), .C(X), .D(n104), .Y(n105));
NAND4X1  g37(.A(Y_2), .B(C_2), .C(X), .D(n103_1), .Y(n106));
AND2X1   g25(.A(Y_7), .B(C_7), .Y(n94));
NAND2X1  g27(.A(Y_6), .B(C_6), .Y(n96));
NAND2X1  g29(.A(Y_5), .B(C_5), .Y(n98_1));
INVX1    g08(.A(X), .Y(n77));
AND2X1   g38(.A(Y_1), .B(C_1), .Y(n107));
NAND2X1  g31(.A(Y_4), .B(C_4), .Y(n100));
AND2X1   g35(.A(Y_3), .B(C_3), .Y(n104));
INVX1    g33(.A(Y_2), .Y(n102));
INVX1    g34(.A(Y_1), .Y(n103_1));

endmodule
