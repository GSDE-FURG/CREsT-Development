//Converted to Combinational , Module name: s641 , Timestamp: 2018-12-03T15:51:01.880008 
module s641 ( G1, G2, G3, G4, G5, G6, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G64, G65, G66, G67, G68, G69, G70, G71, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G91, G94, G107, G83, G84, G85, G100BF, G98BF, G96BF, G92, G87BF, G89BF, G101BF, G106BF, G97BF, G104BF, G88BF, G99BF, G105BF, G138, G86BF, G95BF, G103BF, G90, n119, n124, n129, n134, n139, n144, n148, n153, n158, n163, n168, n173, n178, n183, n188, n193, n198, n203, n208 );
input G1, G2, G3, G4, G5, G6, G8, G9, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G30, G31, G32, G33, G34, G35, G36, G64, G65, G66, G67, G68, G69, G70, G71, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82;
output G91, G94, G107, G83, G84, G85, G100BF, G98BF, G96BF, G92, G87BF, G89BF, G101BF, G106BF, G97BF, G104BF, G88BF, G99BF, G105BF, G138, G86BF, G95BF, G103BF, G90, n119, n124, n129, n134, n139, n144, n148, n153, n158, n163, n168, n173, n178, n183, n188, n193, n198, n203, n208;
wire n116, n118, n120, n122, n124_1, n128, n129_1, n131, n132, n133, n134_1, n135, n137, n138, n139_1, n140, n141, n142, n145, n146, n147, n148_1, n151, n152, n154, n155, n156, n157, n158_1, n159, n160, n163_1, n164, n167, n168_1, n169, n171, n172, n173_1, n174, n175, n177, n179, n182, n183_1, n184, n185, n186, n188_1, n189, n190, n191, n192, n193_1, n194, n195, n196, n197, n198_1, n199, n204, n209, n210, n211, n212, n214, n215, n216, n218, n219, n220, n222, n223, n224;
NAND2X1  g000(.A(G79), .B(G18), .Y(n116));
NOR2X1   g001(.A(n116), .B(G4), .Y(G107));
NAND2X1  g002(.A(G80), .B(G19), .Y(n118));
NOR2X1   g003(.A(n118), .B(G4), .Y(G83));
NAND2X1  g004(.A(G81), .B(G20), .Y(n120));
NOR2X1   g005(.A(n120), .B(G4), .Y(G84));
NAND2X1  g006(.A(G82), .B(G21), .Y(n122));
NOR2X1   g007(.A(n122), .B(G4), .Y(G85));
INVX1    g008(.A(G4), .Y(n124_1));
NAND3X1  g009(.A(G69), .B(G35), .C(n124_1), .Y(G100BF));
NAND3X1  g010(.A(G71), .B(G33), .C(n124_1), .Y(G98BF));
NAND3X1  g011(.A(G73), .B(G31), .C(n124_1), .Y(G96BF));
NAND2X1  g012(.A(G28), .B(G12), .Y(n128));
NAND2X1  g013(.A(G13), .B(G11), .Y(n129_1));
NOR2X1   g014(.A(n129_1), .B(n128), .Y(G92));
INVX1    g015(.A(G23), .Y(n131));
INVX1    g016(.A(G10), .Y(n132));
NOR4X1   g017(.A(n132), .B(G9), .C(G3), .D(G13), .Y(n133));
NOR2X1   g018(.A(G11), .B(G3), .Y(n134_1));
NOR4X1   g019(.A(n133), .B(G65), .C(n131), .D(n134_1), .Y(n135));
INVX1    g020(.A(n135), .Y(G87BF));
INVX1    g021(.A(G3), .Y(n137));
INVX1    g022(.A(G13), .Y(n138));
NAND4X1  g023(.A(G10), .B(G9), .C(n137), .D(n138), .Y(n139_1));
INVX1    g024(.A(G25), .Y(n140));
NOR3X1   g025(.A(n134_1), .B(G67), .C(n140), .Y(n141));
AND2X1   g026(.A(n141), .B(n139_1), .Y(n142));
INVX1    g027(.A(n142), .Y(G89BF));
NAND4X1  g028(.A(n139_1), .B(G68), .C(G36), .D(n141), .Y(G101BF));
INVX1    g029(.A(G78), .Y(n145));
AOI21X1  g030(.A0(n141), .A1(n139_1), .B0(G3), .Y(n146));
OR2X1    g031(.A(n146), .B(n145), .Y(n147));
INVX1    g032(.A(n147), .Y(n148_1));
NAND2X1  g033(.A(n148_1), .B(G17), .Y(G106BF));
NAND3X1  g034(.A(n135), .B(G72), .C(G32), .Y(G97BF));
OAI21X1  g035(.A0(n135), .A1(G3), .B0(G76), .Y(n151));
INVX1    g036(.A(n151), .Y(n152));
NAND2X1  g037(.A(n152), .B(G15), .Y(G104BF));
INVX1    g038(.A(G2), .Y(n154));
AND2X1   g039(.A(G66), .B(n154), .Y(n155));
OAI21X1  g040(.A0(n146), .A1(n145), .B0(n155), .Y(n156));
INVX1    g041(.A(G9), .Y(n157));
NOR4X1   g042(.A(G10), .B(n157), .C(G3), .D(G13), .Y(n158_1));
OAI21X1  g043(.A0(G11), .A1(G3), .B0(G24), .Y(n159));
NOR2X1   g044(.A(n159), .B(n158_1), .Y(n160));
NAND2X1  g045(.A(n160), .B(n156), .Y(G88BF));
NAND4X1  g046(.A(n156), .B(G70), .C(G34), .D(n160), .Y(G99BF));
INVX1    g047(.A(G77), .Y(n163_1));
AOI21X1  g048(.A0(n160), .A1(n156), .B0(G3), .Y(n164));
NOR2X1   g049(.A(n164), .B(n163_1), .Y(n129));
NAND2X1  g050(.A(n129), .B(G16), .Y(G105BF));
NAND2X1  g051(.A(G69), .B(n124_1), .Y(n167));
INVX1    g052(.A(n167), .Y(n168_1));
NAND3X1  g053(.A(n160), .B(n156), .C(G70), .Y(n169));
NAND2X1  g054(.A(n169), .B(n168_1), .Y(G138));
OAI21X1  g055(.A0(n164), .A1(n163_1), .B0(n147), .Y(n171));
NAND3X1  g056(.A(n151), .B(G64), .C(n154), .Y(n172));
NOR4X1   g057(.A(G10), .B(G9), .C(G3), .D(G13), .Y(n173_1));
OAI21X1  g058(.A0(G11), .A1(G3), .B0(G22), .Y(n174));
NOR2X1   g059(.A(n174), .B(n173_1), .Y(n175));
OAI21X1  g060(.A0(n172), .A1(n171), .B0(n175), .Y(G86BF));
OR2X1    g061(.A(n172), .B(n171), .Y(n177));
NAND4X1  g062(.A(n177), .B(G74), .C(G30), .D(n175), .Y(G95BF));
INVX1    g063(.A(G75), .Y(n179));
AOI21X1  g064(.A0(G86BF), .A1(n137), .B0(n179), .Y(n119));
NAND2X1  g065(.A(n119), .B(G14), .Y(G103BF));
INVX1    g066(.A(G74), .Y(n182));
AND2X1   g067(.A(G73), .B(n124_1), .Y(n183_1));
NAND4X1  g068(.A(n138), .B(n132), .C(n157), .D(n183_1), .Y(n184));
NOR3X1   g069(.A(n184), .B(G86BF), .C(n182), .Y(n185));
NAND3X1  g070(.A(n141), .B(n139_1), .C(G68), .Y(n186));
INVX1    g071(.A(n186), .Y(n139));
AND2X1   g072(.A(n135), .B(G72), .Y(n188_1));
NAND2X1  g073(.A(G71), .B(n124_1), .Y(n189));
NAND3X1  g074(.A(G73), .B(G69), .C(n124_1), .Y(n190));
NOR3X1   g075(.A(n190), .B(n189), .C(G11), .Y(n191));
NAND3X1  g076(.A(n191), .B(n188_1), .C(n139), .Y(n192));
NOR4X1   g077(.A(G86BF), .B(n169), .C(n182), .D(n192), .Y(n193_1));
OR4X1    g078(.A(G13), .B(G10), .C(n157), .D(n167), .Y(n194));
NOR4X1   g079(.A(G13), .B(n132), .C(G9), .D(n189), .Y(n195));
OR4X1    g080(.A(G13), .B(n132), .C(n157), .D(n186), .Y(n196));
NAND3X1  g081(.A(n196), .B(G26), .C(G12), .Y(n197));
AOI21X1  g082(.A0(n195), .A1(n188_1), .B0(n197), .Y(n198_1));
OAI21X1  g083(.A0(n194), .A1(n169), .B0(n198_1), .Y(n199));
NOR3X1   g084(.A(n199), .B(n193_1), .C(n185), .Y(G90));
NOR4X1   g085(.A(n151), .B(n148_1), .C(G2), .D(n129), .Y(n124));
NOR3X1   g086(.A(n146), .B(n145), .C(G2), .Y(n134));
MX2X1    g087(.A(G70), .B(n168_1), .S0(G88BF), .Y(n144));
INVX1    g088(.A(n188_1), .Y(n204));
OAI21X1  g089(.A0(n135), .A1(n189), .B0(n204), .Y(n153));
OR2X1    g090(.A(n188_1), .B(n189), .Y(n158));
MX2X1    g091(.A(G74), .B(n183_1), .S0(G86BF), .Y(n163));
OAI21X1  g092(.A0(G86BF), .A1(n182), .B0(n183_1), .Y(n168));
NAND2X1  g093(.A(n119), .B(n154), .Y(n209));
NAND4X1  g094(.A(n147), .B(n183_1), .C(G8), .D(n151), .Y(n210));
NOR4X1   g095(.A(G86BF), .B(n129), .C(n182), .D(n210), .Y(n211));
AOI21X1  g096(.A0(n119), .A1(G8), .B0(n211), .Y(n212));
NAND2X1  g097(.A(n212), .B(n209), .Y(n173));
NAND3X1  g098(.A(G71), .B(G5), .C(n124_1), .Y(n214));
OR4X1    g099(.A(n129), .B(n204), .C(n148_1), .D(n214), .Y(n215));
OAI21X1  g100(.A0(G5), .A1(n154), .B0(n152), .Y(n216));
OAI21X1  g101(.A0(n215), .A1(n119), .B0(n216), .Y(n178));
NAND4X1  g102(.A(n147), .B(n168_1), .C(G6), .D(n151), .Y(n218));
OR2X1    g103(.A(n218), .B(n169), .Y(n219));
OAI21X1  g104(.A0(G6), .A1(n154), .B0(n129), .Y(n220));
OAI21X1  g105(.A0(n219), .A1(n119), .B0(n220), .Y(n183));
NAND3X1  g106(.A(n151), .B(n139), .C(G1), .Y(n222));
OR2X1    g107(.A(n222), .B(n129), .Y(n223));
OAI21X1  g108(.A0(n154), .A1(G1), .B0(n148_1), .Y(n224));
OAI21X1  g109(.A0(n223), .A1(n119), .B0(n224), .Y(n188));
NOR3X1   g110(.A(n209), .B(n171), .C(n152), .Y(n193));
NOR4X1   g111(.A(n148_1), .B(n163_1), .C(G2), .D(n164), .Y(n203));
BUFX1    g112(.A(G27), .Y(G91));
BUFX1    g113(.A(G29), .Y(G94));
NAND2X1  g114(.A(n169), .B(n168_1), .Y(n148));
NOR4X1   g115(.A(n151), .B(n148_1), .C(G2), .D(n129), .Y(n198));
NOR3X1   g116(.A(n146), .B(n145), .C(G2), .Y(n208));
endmodule
