//Converted to Combinational , Module name: s208
module s208 ( X, Clear, C_8, C_7, C_6, C_5, C_4, C_3, C_2, C_1, C_0, Y_4, Y_3, Y_2, Y_1, Y_8, Y_7, Y_6, Y_5, W, Z, n27, n32, n37, n42, n47, n52, n57, n62 );
input X, Clear, C_8, C_7, C_6, C_5, C_4, C_3, C_2, C_1, C_0, Y_4, Y_3, Y_2, Y_1, Y_8, Y_7, Y_6, Y_5;
output W, Z, n27, n32, n37, n42, n47, n52, n57, n62;
wire n37_1, n38, n40, n41, n42_1, n43, n44, n45, n46, n47_1, n48, n49, n50, n51, n52_1, n53, n54, n55, n56, n57_1, n58, n59, n60, n61, n62_1, n64, n65, n66, n67, n68, n70, n71, n72, n74, n75, n78, n79, n80, n81, n83, n84, n85;
INVX1    g00(.A(Y_8), .Y(n37_1));
NAND3X1  g01(.A(Y_5), .B(Y_6), .C(Y_7), .Y(n38));
NOR2X1   g02(.A(n38), .B(n37_1), .Y(W));
INVX1    g03(.A(Y_4), .Y(n40));
INVX1    g04(.A(Y_5), .Y(n41));
INVX1    g05(.A(X), .Y(n42_1));
NOR4X1   g06(.A(Y_2), .B(Y_3), .C(n42_1), .D(Y_1), .Y(n43));
AND2X1   g07(.A(Y_6), .B(C_6), .Y(n44));
NAND4X1  g08(.A(n43), .B(n41), .C(n40), .D(n44), .Y(n45));
NAND4X1  g09(.A(Y_5), .B(n40), .C(C_5), .D(n43), .Y(n46));
NAND3X1  g10(.A(n43), .B(Y_4), .C(C_4), .Y(n47_1));
NAND2X1  g11(.A(Y_3), .B(C_3), .Y(n48));
NOR4X1   g12(.A(Y_1), .B(Y_2), .C(n42_1), .D(n48), .Y(n49));
NAND2X1  g13(.A(Y_2), .B(C_2), .Y(n50));
NOR3X1   g14(.A(n50), .B(Y_1), .C(n42_1), .Y(n51));
NAND2X1  g15(.A(C_0), .B(X), .Y(n52_1));
NAND3X1  g16(.A(Y_1), .B(C_1), .C(X), .Y(n53));
NAND2X1  g17(.A(n53), .B(n52_1), .Y(n54));
NOR3X1   g18(.A(n54), .B(n51), .C(n49), .Y(n55));
AND2X1   g19(.A(n55), .B(n47_1), .Y(n56));
OR4X1    g20(.A(Y_2), .B(Y_3), .C(n42_1), .D(Y_1), .Y(n57_1));
NOR4X1   g21(.A(Y_5), .B(Y_6), .C(Y_4), .D(n57_1), .Y(n58));
NAND2X1  g22(.A(Y_8), .B(C_8), .Y(n59));
NOR2X1   g23(.A(n59), .B(Y_7), .Y(n60));
AND2X1   g24(.A(Y_7), .B(C_7), .Y(n61));
OAI21X1  g25(.A0(n61), .A1(n60), .B0(n58), .Y(n62_1));
NAND4X1  g26(.A(n56), .B(n46), .C(n45), .D(n62_1), .Y(Z));
INVX1    g27(.A(Clear), .Y(n64));
NAND4X1  g28(.A(Y_2), .B(n64), .C(X), .D(Y_1), .Y(n65));
NAND2X1  g29(.A(Y_3), .B(n40), .Y(n66));
NAND3X1  g30(.A(Y_1), .B(Y_2), .C(Y_3), .Y(n67));
NAND4X1  g31(.A(Y_4), .B(n64), .C(X), .D(n67), .Y(n68));
OAI21X1  g32(.A0(n66), .A1(n65), .B0(n68), .Y(n27));
INVX1    g33(.A(Y_3), .Y(n70));
AND2X1   g34(.A(Y_1), .B(Y_2), .Y(n71));
OR4X1    g35(.A(n70), .B(Clear), .C(n42_1), .D(n71), .Y(n72));
OAI21X1  g36(.A0(n65), .A1(Y_3), .B0(n72), .Y(n32));
INVX1    g37(.A(Y_1), .Y(n74));
NOR3X1   g38(.A(n74), .B(Clear), .C(n42_1), .Y(n75));
NOR3X1   g39(.A(Y_1), .B(Clear), .C(n42_1), .Y(n42));
MX2X1    g40(.A(n75), .B(n42), .S0(Y_2), .Y(n37));
NAND4X1  g41(.A(Y_3), .B(Y_4), .C(n64), .D(n71), .Y(n78));
NOR4X1   g42(.A(n41), .B(n40), .C(Clear), .D(n67), .Y(n79));
NAND4X1  g43(.A(Y_6), .B(Y_7), .C(n37_1), .D(n79), .Y(n80));
NAND2X1  g44(.A(n38), .B(Y_8), .Y(n81));
OAI21X1  g45(.A0(n81), .A1(n78), .B0(n80), .Y(n47));
NAND2X1  g46(.A(n79), .B(Y_6), .Y(n83));
NAND2X1  g47(.A(Y_5), .B(Y_6), .Y(n84));
NAND2X1  g48(.A(n84), .B(Y_7), .Y(n85));
OAI22X1  g49(.A0(n83), .A1(Y_7), .B0(n78), .B1(n85), .Y(n52));
NOR4X1   g50(.A(Y_5), .B(n40), .C(Clear), .D(n67), .Y(n62));
MX2X1    g51(.A(n79), .B(n62), .S0(Y_6), .Y(n57));
endmodule
