//Converted to Combinational , Module name: s38584 , Timestamp: 2018-12-03T15:51:15.799249 
module s38584 ( g35, g36, g6744, g6745, g6746, g6747, g6748, g6749, g6750, g6751, g6752, g6753, g84, g120, g5, g113, g126, g99, g53, g116, g92, g56, g91, g44, g57, g100, g54, g124, g125, g114, g134, g72, g115, g135, g90, g127, g64, g73, g5057, g2771, g1882, g6462, g2299, g4040, g2547, g559, g3017, g3243, g452, g464, g3542, g5232, g5813, g2907, g1744, g5909, g1802, g3554, g6219, g807, g6031, g847, g976, g4172, g4372, g3512, g749, g3490, g6005, g4235, g1600, g1714, g3649, g3155, g3355, g2236, g4555, g3698, g6073, g1736, g1968, g4621, g5607, g2657, g5659, g490, g311, g6069, g772, g5587, g6177, g6377, g3167, g5615, g4567, g3057, g3457, g6287, g1500, g2563, g4776, g4593, g6199, g2295, g1384, g1339, g5180, g2844, g1024, g5591, g3598, g4264, g767, g5853, g3321, g2089, g4933, g4521, g5507, g3625, g6291, g294, g5559, g5794, g6144, g3813, g562, g608, g1205, g3909, g6259, g5905, g921, g2955, g203, g6088, g1099, g4878, g5204, g5630, g3606, g1926, g6215, g3586, g291, g4674, g3570, g640, g5969, g1862, g676, g843, g4132, g4332, g4153, g5666, g6336, g622, g3506, g4558, g6065, g6322, g3111, g117, g2837, g939, g278, g4492, g4864, g1036, g128, g1178, g3239, g718, g6195, g1135, g6137, g6395, g3380, g5343, g554, g496, g3853, g5134, g1422, g3794, g2485, g925, g5555, g878, g1798, g4076, g2941, g3905, g763, g6255, g4375, g4871, g4722, g6692, g1632, g5313, g3100, g1495, g6497, g1437, g6154, g1579, g5567, g1752, g1917, g744, g3040, g4737, g4809, g6267, g3440, g3969, g1442, g5965, g4477, g1233, g4643, g5264, g6329, g2610, g5160, g5360, g5933, g1454, g753, g1296, g3151, g2980, g6727, g3530, g4742, g4104, g1532, g4304, g2177, g3010, g4754, g1189, g2287, g4273, g1389, g1706, g5835, g1171, g4269, g2399, g3372, g4983, g5611, g3618, g4572, g3143, g2898, g3343, g3235, g4543, g3566, g4534, g4961, g6398, g4927, g2259, g2819, g4414, g5802, g2852, g681, g5901, g2886, g3494, g5511, g3518, g1604, g4135, g5092, g4831, g4382, g6386, g479, g3965, g4749, g2008, g736, g3933, g222, g3050, g5736, g1052, g5623, g2122, g2465, g6483, g5889, g4495, g365, g4653, g3179, g1728, g2433, g3835, g6187, g4917, g1070, g822, g6027, g914, g5339, g4164, g969, g2807, g5424, g4054, g6191, g5077, g5523, g3680, g6637, g1682, g1087, g1105, g2342, g6307, g3802, g6159, g2255, g2815, g911, g4012, g1748, g5551, g5742, g3558, g5499, g2960, g3901, g4888, g6251, g6315, g1373, g3092, g2783, g4281, g3574, g2112, g1283, g4297, g5983, g1459, g758, g5712, g4138, g4639, g6537, g5543, g1582, g3736, g5961, g6243, g1227, g3889, g3476, g1664, g1246, g6128, g6629, g4049, g4449, g2932, g4575, g4098, g4498, g528, g5436, g3139, g4584, g5335, g5831, g1216, g2848, g5805, g5022, g4019, g1030, g3672, g3231, g6490, g1430, g4452, g2241, g1564, g5798, g6148, g6649, g884, g3742, g4486, g4504, g5873, g5037, g2319, g5495, g4185, g5208, g2152, g5579, g5869, g5719, g1589, g5752, g6279, g5917, g2975, g6167, g3983, g2599, g1448, g881, g3712, g2370, g5164, g1333, g6549, g4087, g4801, g2984, g3961, g5770, g962, g101, g4226, g6625, g1018, g1418, g4045, g1467, g2461, g5706, g2756, g5990, g471, g1256, g5029, g6519, g4169, g1816, g4369, g3436, g5787, g4578, g4459, g3831, g2514, g3288, g2403, g2145, g1700, g2841, g5297, g3805, g2763, g4793, g952, g1263, g1950, g5138, g2307, g5109, g5791, g3798, g4664, g2223, g5808, g6645, g2016, g5759, g3873, g3632, g2315, g2811, g5957, g2047, g3869, g6358, g3719, g5575, g3752, g3917, g4188, g1585, g4388, g6275, g6311, g4216, g1041, g2595, g2537, g136, g4430, g4564, g3454, g4826, g6239, g3770, g232, g5268, g6545, g2417, g1772, g4741, g5052, g5452, g1890, g2629, g572, g2130, g4108, g4308, g990, g3412, g799, g3706, g3990, g5385, g5881, g1992, g3029, g3171, g3787, g812, g832, g5897, g4165, g4571, g3281, g4455, g2902, g333, g2823, g3684, g3639, g5331, g3338, g5406, g3791, g269, g6040, g5105, g3808, g3759, g4467, g3957, g4093, g1760, g6151, g6351, g5445, g5373, g2279, g3498, g869, g2619, g1183, g1608, g4197, g5283, g1779, g2652, g5459, g2193, g2393, g5767, g661, g4950, g5535, g2834, g1361, g3419, g6235, g1146, g2625, g1696, g6555, g859, g3385, g3881, g6621, g3470, g3897, g3025, g2606, g1472, g6113, g5188, g5689, g1116, g5216, g6494, g4669, g5428, g996, g4531, g2860, g4743, g6593, g2710, g4411, g1413, g4474, g5308, g6641, g3045, g1936, g504, g2587, g4480, g2311, g3602, g5571, g3578, g468, g5448, g3767, g5827, g3582, g6271, g4688, g5774, g2380, g5196, g5396, g3227, g2020, g4000, g1079, g6541, g3203, g1668, g4760, g1840, g70, g5467, g460, g6209, g5290, g3502, g2204, g5256, g4608, g794, g4023, g4423, g3689, g5381, g5685, g703, g5421, g862, g3247, g2040, g4999, g4146, g4633, g1157, g5723, g4732, g5101, g5817, g2151, g2351, g2648, g6736, g4944, g4072, g4443, g3466, g4116, g5041, g5441, g4434, g3827, g6500, g5673, g3133, g3333, g979, g4681, g3774, g2667, g3396, g4210, g1894, g2988, g3538, g827, g1075, g6077, g2555, g5011, g6523, g1526, g4601, g854, g1484, g4922, g5080, g5863, g4581, g3021, g2518, g2567, g3263, g6613, g6044, g6444, g2965, g5857, g1616, g890, g5976, g3562, g4294, g1404, g3723, g3817, g4501, g287, g2724, g4704, g2878, g5220, g1277, g6513, g336, g2882, g933, g1906, g3368, g2799, g887, g5327, g4912, g4157, g2541, g2153, g1945, g5240, g1478, g3080, g3863, g1959, g3480, g6653, g6719, g2864, g4894, g5681, g3857, g3976, g5413, g1002, g776, g1236, g4646, g2476, g1657, g2375, g6012, g896, g967, g3423, g3161, g2384, g3361, g6675, g4616, g4561, g2024, g3451, g2795, g4527, g1844, g5937, g4546, g3103, g2523, g3303, g2643, g6109, g1489, g5390, g2551, g5156, g3072, g1242, g3443, g4277, g1955, g6049, g3034, g2273, g6715, g4771, g6098, g3147, g3347, g2269, g2712, g2729, g5357, g4991, g6019, g4709, g6419, g6052, g2927, g4340, g5929, g4907, g3317, g4035, g2946, g918, g4082, g6486, g2036, g1620, g2831, g930, g3937, g5782, g817, g1249, g837, g3668, g5475, g739, g5949, g6682, g6105, g904, g2873, g1854, g5084, g5603, g4222, g2495, g2437, g2102, g2208, g2579, g4064, g4899, g2719, g4785, g5583, g781, g6173, g6373, g2917, g686, g1252, g2265, g6283, g6369, g5276, g6459, g901, g4194, g5527, g4489, g1974, g1270, g4966, g6415, g6227, g3929, g5503, g4242, g5925, g1124, g4955, g5224, g2012, g6203, g5120, g5320, g2389, g4438, g2429, g2787, g1287, g2675, g4836, g1199, g1399, g5547, g3782, g6428, g2138, g3661, g2338, g4229, g6247, g2791, g3949, g1291, g5945, g5244, g2759, g6741, g785, g1259, g3484, g209, g6609, g5517, g2449, g2575, g2715, g936, g2098, g4462, g6589, g1886, g6466, g6365, g6711, g1870, g4249, g6455, g3004, g1825, g6133, g1008, g4392, g5002, g3546, g5236, g1768, g4854, g3925, g6509, g732, g2504, g1322, g4520, g4219, g2185, g4031, g2070, g4812, g6093, g968, g4176, g4005, g4405, g872, g6181, g6381, g4765, g5563, g1395, g1913, g2331, g6263, g3945, g5731, g4473, g1266, g5489, g714, g2748, g5471, g4540, g6723, g6605, g2445, g2173, g4287, g2491, g4849, g2169, g2283, g6585, g2407, g2868, g2767, g1783, g3310, g1312, g5212, g4245, g4291, g1129, g2227, g6058, g4207, g2246, g1830, g3590, g1592, g6505, g6411, g1221, g5921, g106, g6474, g1932, g1624, g5062, g5462, g2689, g6573, g1677, g2028, g2671, g1576, g4408, g1848, g3089, g3731, g5485, g2741, g802, g2638, g4122, g4322, g5941, g2108, g6000, g1644, g2217, g1319, g2066, g1152, g5252, g2165, g2571, g5176, g5005, g2711, g6023, g1211, g2827, g6423, g875, g4859, g1274, g1426, g2803, g6451, g1821, g2509, g5073, g1280, g4815, g6346, g6633, g5124, g1083, g6303, g5069, g2994, g1636, g3921, g2093, g6732, g1306, g5377, g1061, g3462, g2181, g956, g1756, g5849, g4112, g2685, g2197, g6116, g2421, g1046, g4401, g6434, g1514, g329, g6565, g2950, g4129, g1345, g6533, g3298, g3085, g4727, g6697, g1536, g3941, g5694, g1858, g4932, g3219, g1811, g3431, g6601, g3376, g2441, g1874, g4349, g6581, g6597, g5008, g3610, g2890, g1978, g1612, g2856, g6479, g1982, g6668, g5228, g4119, g6390, g1542, g4258, g4818, g5033, g4717, g1554, g3849, g6704, g3199, g5845, g4975, g790, g5913, g1902, g6163, g4125, g4821, g4939, g1056, g3207, g4483, g3259, g5142, g5248, g2126, g3694, g5481, g1964, g5097, g3215, g4027, g4427, g2779, g4200, g4446, g1720, g1367, g5112, g4145, g2161, g2361, g4191, g2051, g1193, g5401, g3408, g2327, g907, g947, g1834, g3594, g2999, g5727, g2303, g6661, g3065, g699, g723, g5703, g2472, g5953, g3096, g6439, g1740, g3550, g3845, g2116, g5677, g3195, g3913, g4537, g1687, g2681, g2533, g2697, g5747, g4417, g6561, g1141, g1570, g2413, g1710, g6527, g6404, g3255, g1691, g2936, g5644, g5152, g5352, g4213, g6120, g2775, g2922, g1111, g5893, g1311, g3267, g6617, g2060, g4512, g5599, g3401, g4366, g3676, g3129, g3329, g5170, g4456, g5821, g6299, g1239, g3727, g2079, g4698, g3703, g1559, g943, g6140, g3953, g3068, g2704, g6035, g6082, g1300, g4057, g5200, g4843, g5046, g2250, g4549, g2453, g5841, g5763, g3747, g5637, g2912, g2357, g4232, g4253, g5016, g3119, g1351, g1648, g4519, g5115, g3352, g6657, g4552, g3893, g3211, g5654, g929, g3274, g5595, g3614, g2894, g3125, g3325, g3821, g4141, g4570, g5272, g2735, g728, g6295, g5417, g2661, g1988, g5128, g1548, g3106, g4659, g4358, g1792, g2084, g3061, g3187, g4311, g2583, g3003, g1094, g3841, g4284, g3763, g3191, g4239, g3391, g4180, g691, g5366, g2004, g2527, g5456, g4420, g5148, g4507, g5348, g3223, g4931, g2970, g5698, g3416, g5260, g1521, g3522, g3115, g3251, g4628, g1996, g3447, g4515, g4204, g4300, g1724, g1379, g3654, g1878, g5619, g7243, g7245, g7257, g7260, g7540, g7916, g7946, g8132, g8178, g8215, g8235, g8277, g8279, g8283, g8291, g8342, g8344, g8353, g8358, g8398, g8403, g8416, g8475, g8719, g8783, g8784, g8785, g8786, g8787, g8788, g8789, g8839, g8870, g8915, g8916, g8917, g8918, g8919, g8920, g9019, g9048, g9251, g9497, g9553, g9555, g9615, g9617, g9680, g9682, g9741, g9743, g9817, g10122, g10306, g10500, g10527, g11349, g11388, g11418, g11447, g11678, g11770, g12184, g12238, g12300, g12350, g12368, g12422, g12470, g12832, g12919, g12923, g13039, g13049, g13068, g13085, g13099, g13259, g13272, g13865, g13881, g13895, g13906, g13926, g13966, g14096, g14125, g14147, g14167, g14189, g14201, g14217, g14421, g14451, g14518, g14597, g14635, g14662, g14673, g14694, g14705, g14738, g14749, g14779, g14828, g16603, g16624, g16627, g16656, g16659, g16686, g16693, g16718, g16722, g16744, g16748, g16775, g16874, g16924, g16955, g17291, g17316, g17320, g17400, g17404, g17423, g17519, g17577, g17580, g17604, g17607, g17639, g17646, g17649, g17674, g17678, g17685, g17688, g17711, g17715, g17722, g17739, g17743, g17760, g17764, g17778, g17787, g17813, g17819, g17845, g17871, g18092, g18094, g18095, g18096, g18097, g18098, g18099, g18100, g18101, g18881, g19334, g19357, g20049, g20557, g20652, g20654, g20763, g20899, g20901, g21176, g21245, g21270, g21292, g21698, g21727, g23002, g23190, g23612, g23652, g23683, g23759, g24151, g25114, g25167, g25219, g25259, g25582, g25583, g25584, g25585, g25586, g25587, g25588, g25589, g25590, g26801, g26875, g26876, g26877, g27831, g28030, g28041, g28042, g28753, g29210, g29211, g29212, g29213, g29214, g29215, g29216, g29217, g29218, g29219, g29220, g29221, g30327, g30329, g30330, g30331, g30332, g31521, g31656, g31665, g31793, g31860, g31861, g31862, g31863, g32185, g32429, g32454, g32975, g33079, g33435, g33533, g33636, g33659, g33874, g33894, g33935, g33945, g33946, g33947, g33948, g33949, g33950, g33959, g34201, g34221, g34232, g34233, g34234, g34235, g34236, g34237, g34238, g34239, g34240, g34383, g34425, g34435, g34436, g34437, g34597, g34788, g34839, g34913, g34915, g34917, g34919, g34921, g34923, g34925, g34927, g34956, g34972, g24168, g24178, g12833, g24174, g24181, g24172, g24161, g24177, g24171, g24163, g24170, g24185, g24164, g24173, g24162, g24179, g24180, g24175, g24183, g24166, g24176, g24184, g24169, g24182, g24165, g24167, n685, n690, n695, n700, n705, n710, n715, n720, n725, n730, n735, n740, n745, n750, n755, n760, n765, n770, n775, n780, n785, n790, n795, n800, n805, n810, n815, n820, n825, n830, n835, n840, n845, n850, n855, n860, n865, n870, n875, n880, n885, n890, n895, n900, n905, n910, n915, n920, n925, n930, n935, n940, n945, n950, n955, n960, n965, n970, n975, n980, n985, n990, n995, n1000, n1005, n1010, n1015, n1020, n1025, n1030, n1035, n1040, n1045, n1050, n1055, n1060, n1065, n1070, n1075, n1080, n1085, n1090, n1094, n1099, n1104, n1109, n1114, n1119, n1124, n1129, n1134, n1139, n1144, n1149, n1154, n1159, n1164, n1169, n1174, n1179, n1184, n1189, n1194, n1199, n1204, n1209, n1214, n1219, n1224, n1229, n1233, n1238, n1243, n1248, n1253, n1258, n1263, n1268, n1273, n1278, n1283, n1288, n1293, n1298, n1303, n1308, n1313, n1318, n1323, n1328, n1333, n1338, n1343, n1348, n1353, n1358, n1363, n1368, n1373, n1378, n1383, n1388, n1393, n1398, n1403, n1408, n1413, n1418, n1423, n1428, n1433, n1438, n1443, n1448, n1453, n1458, n1463, n1468, n1473, n1478, n1483, n1488, n1493, n1498, n1503, n1508, n1513, n1518, n1523, n1528, n1533, n1538, n1543, n1548, n1553, n1558, n1563, n1568, n1573, n1578, n1583, n1588, n1593, n1598, n1603, n1608, n1613, n1618, n1623, n1628, n1633, n1638, n1643, n1648, n1653, n1658, n1663, n1668, n1673, n1678, n1683, n1688, n1693, n1698, n1703, n1708, n1713, n1718, n1723, n1728, n1733, n1738, n1743, n1748, n1753, n1758, n1763, n1768, n1773, n1778, n1783, n1787, n1792, n1797, n1802, n1807, n1812, n1817, n1822, n1827, n1832, n1837, n1842, n1847, n1852, n1856, n1861, n1866, n1871, n1876, n1881, n1886, n1891, n1896, n1901, n1906, n1911, n1916, n1921, n1926, n1931, n1936, n1941, n1946, n1951, n1956, n1961, n1966, n1971, n1976, n1981, n1986, n1991, n1995, n1999, n2004, n2009, n2014, n2019, n2024, n2029, n2034, n2039, n2044, n2049, n2054, n2059, n2064, n2069, n2074, n2078, n2083, n2088, n2093, n2098, n2103, n2108, n2113, n2118, n2123, n2128, n2133, n2138, n2143, n2148, n2153, n2158, n2163, n2168, n2172, n2177, n2182, n2187, n2192, n2197, n2202, n2206, n2211, n2216, n2221, n2226, n2231, n2236, n2241, n2246, n2251, n2255, n2260, n2264, n2269, n2274, n2279, n2284, n2289, n2294, n2299, n2303, n2308, n2313, n2318, n2323, n2328, n2333, n2338, n2342, n2347, n2352, n2357, n2362, n2367, n2372, n2377, n2382, n2387, n2392, n2397, n2402, n2407, n2412, n2417, n2422, n2427, n2432, n2437, n2442, n2447, n2452, n2457, n2462, n2467, n2472, n2476, n2481, n2486, n2491, n2496, n2501, n2506, n2511, n2516, n2521, n2526, n2530, n2535, n2540, n2545, n2550, n2554, n2559, n2564, n2569, n2574, n2579, n2584, n2589, n2594, n2599, n2604, n2609, n2614, n2619, n2624, n2629, n2634, n2639, n2644, n2649, n2654, n2659, n2664, n2669, n2674, n2678, n2683, n2687, n2691, n2696, n2701, n2705, n2710, n2715, n2720, n2725, n2730, n2735, n2740, n2745, n2750, n2755, n2760, n2765, n2770, n2775, n2779, n2784, n2789, n2794, n2799, n2804, n2809, n2814, n2819, n2824, n2829, n2834, n2839, n2844, n2849, n2854, n2859, n2864, n2869, n2874, n2879, n2884, n2889, n2894, n2899, n2904, n2909, n2914, n2919, n2924, n2929, n2934, n2939, n2944, n2949, n2954, n2959, n2964, n2968, n2973, n2978, n2983, n2988, n2993, n2998, n3003, n3008, n3013, n3018, n3023, n3028, n3032, n3036, n3041, n3046, n3051, n3056, n3061, n3066, n3071, n3076, n3081, n3086, n3091, n3096, n3101, n3106, n3111, n3116, n3121, n3126, n3131, n3136, n3141, n3146, n3151, n3156, n3161, n3166, n3171, n3176, n3181, n3186, n3191, n3196, n3201, n3205, n3210, n3215, n3220, n3225, n3230, n3235, n3240, n3245, n3250, n3255, n3260, n3265, n3270, n3275, n3280, n3285, n3290, n3295, n3300, n3304, n3309, n3314, n3319, n3324, n3329, n3334, n3339, n3344, n3348, n3353, n3358, n3363, n3368, n3373, n3378, n3383, n3388, n3393, n3398, n3403, n3408, n3413, n3418, n3422, n3427, n3431, n3436, n3441, n3446, n3451, n3456, n3461, n3466, n3471, n3476, n3481, n3486, n3491, n3496, n3500, n3505, n3510, n3515, n3520, n3525, n3530, n3535, n3540, n3545, n3550, n3555, n3560, n3565, n3570, n3575, n3580, n3584, n3589, n3594, n3599, n3604, n3609, n3614, n3619, n3624, n3629, n3634, n3639, n3644, n3649, n3654, n3659, n3664, n3669, n3674, n3679, n3684, n3689, n3694, n3699, n3704, n3709, n3714, n3718, n3723, n3728, n3732, n3737, n3742, n3747, n3752, n3757, n3762, n3767, n3772, n3777, n3782, n3787, n3792, n3797, n3802, n3807, n3812, n3817, n3822, n3827, n3832, n3837, n3842, n3847, n3852, n3857, n3862, n3866, n3871, n3876, n3881, n3886, n3891, n3896, n3901, n3906, n3911, n3916, n3921, n3925, n3930, n3935, n3940, n3945, n3950, n3955, n3959, n3964, n3969, n3974, n3979, n3984, n3989, n3994, n3999, n4004, n4009, n4014, n4019, n4024, n4029, n4034, n4039, n4043, n4048, n4053, n4058, n4063, n4068, n4073, n4078, n4082, n4087, n4092, n4097, n4102, n4107, n4112, n4117, n4122, n4127, n4132, n4136, n4141, n4146, n4151, n4156, n4161, n4166, n4171, n4176, n4181, n4186, n4191, n4196, n4201, n4205, n4210, n4215, n4220, n4225, n4230, n4235, n4240, n4245, n4250, n4255, n4260, n4265, n4270, n4275, n4280, n4285, n4290, n4295, n4300, n4305, n4310, n4315, n4320, n4325, n4329, n4334, n4339, n4343, n4348, n4353, n4358, n4363, n4368, n4373, n4378, n4383, n4388, n4393, n4398, n4403, n4407, n4412, n4417, n4422, n4427, n4432, n4437, n4442, n4447, n4452, n4457, n4461, n4465, n4469, n4474, n4479, n4484, n4489, n4494, n4499, n4504, n4509, n4514, n4519, n4524, n4529, n4534, n4539, n4544, n4549, n4554, n4558, n4562, n4566, n4571, n4576, n4581, n4586, n4590, n4595, n4600, n4605, n4610, n4615, n4619, n4622, n4627, n4632, n4637, n4642, n4647, n4652, n4657, n4662, n4667, n4672, n4677, n4682, n4687, n4692, n4697, n4702, n4707, n4712, n4717, n4722, n4727, n4731, n4736, n4741, n4746, n4751, n4756, n4761, n4766, n4770, n4775, n4780, n4784, n4788, n4793, n4798, n4803, n4808, n4812, n4817, n4822, n4827, n4832, n4836, n4841, n4846, n4851, n4856, n4861, n4866, n4871, n4876, n4881, n4886, n4891, n4896, n4901, n4906, n4910, n4915, n4920, n4925, n4930, n4934, n4939, n4944, n4949, n4954, n4959, n4964, n4969, n4974, n4979, n4984, n4988, n4992, n4997, n5002, n5007, n5012, n5017, n5022, n5027, n5032, n5037, n5042, n5047, n5051, n5056, n5061, n5066, n5071, n5076, n5081, n5086, n5091, n5096, n5101, n5106, n5111, n5115, n5120, n5125, n5130, n5135, n5140, n5145, n5149, n5153, n5158, n5162, n5166, n5171, n5176, n5181, n5186, n5191, n5196, n5201, n5206, n5211, n5216, n5221, n5226, n5231, n5236, n5241, n5246, n5250, n5254, n5259, n5264, n5269, n5274, n5279, n5284, n5289, n5294, n5299, n5303, n5308, n5313, n5318, n5322, n5326, n5330, n5335, n5340, n5345, n5350, n5355, n5360, n5365, n5370, n5375, n5380, n5385, n5390, n5395, n5400, n5405, n5410, n5415, n5420, n5425, n5430, n5435, n5440, n5445, n5450, n5455, n5460, n5463, n5467, n5472, n5477, n5482, n5487, n5492, n5497, n5502, n5507, n5511, n5516, n5521, n5526, n5531, n5536, n5541, n5546, n5551, n5555, n5560, n5564, n5568, n5573, n5578, n5583, n5587, n5592, n5597, n5602, n5607, n5611, n5615, n5620, n5625, n5630, n5635, n5640, n5645, n5650, n5655, n5660, n5665, n5669, n5674, n5679, n5684, n5689, n5694, n5699, n5704, n5709, n5713, n5718, n5723, n5728, n5733, n5738, n5743, n5748, n5753, n5758, n5763, n5768, n5773, n5778, n5783, n5787, n5792, n5797, n5802, n5807, n5811, n5816, n5821, n5826, n5831, n5836, n5841, n5845, n5850, n5855, n5860, n5865, n5870, n5875, n5880, n5885, n5890, n5895, n5899, n5904, n5909, n5914, n5919, n5924, n5929, n5934, n5939, n5944, n5949, n5954, n5958, n5962, n5967, n5972, n5977, n5982, n5987, n5992, n5996, n6000, n6005, n6010, n6015, n6020, n6024, n6028, n6033, n6038, n6043, n6048, n6053, n6058, n6063, n6068, n6073, n6078, n6083, n6087, n6092, n6096, n6100, n6105, n6110, n6114, n6118, n6123, n6128, n6132, n6136, n6141, n6146, n6151, n6156, n6161, n6166, n6170, n6174, n6178, n6183, n6187, n6191, n6196, n6201, n6206, n6211, n6216, n6221, n6226, n6231, n6236, n6241, n6246, n6251, n6256, n6261, n6266, n6271, n6276, n6281, n6286, n6291, n6296, n6301, n6306, n6311, n6316, n6321, n6326, n6331, n6336, n6341, n6346, n6351, n6355, n6360, n6365, n6369, n6374, n6379, n6384, n6389, n6394, n6399, n6404, n6409, n6414, n6419, n6424, n6429, n6434, n6439, n6444, n6449, n6453, n6458, n6463, n6468, n6473, n6478, n6483, n6488, n6493, n6498, n6502, n6507, n6512, n6517, n6522, n6526, n6531, n6536, n6541, n6546, n6550, n6555, n6560, n6565, n6570, n6575, n6580, n6585, n6590, n6595, n6600, n6605, n6609, n6613, n6618, n6623, n6628, n6633, n6638, n6643, n6648, n6653, n6658, n6662, n6666, n6671, n6676, n6681, n6685, n6690, n6694, n6699, n6703, n6708, n6713, n6718, n6723, n6728, n6733, n6737, n6742, n6747, n6752, n6757, n6762, n6767, n6772, n6777, n6782, n6787, n6792, n6797, n6801, n6805, n6810, n6815, n6820, n6825, n6830, n6835, n6840, n6844, n6849, n6854, n6859, n6864, n6868, n6872, n6877, n6882, n6886, n6891, n6896, n6901, n6906, n6911, n6916, n6921, n6926, n6931, n6935, n6940, n6945, n6950, n6955, n6960, n6965, n6970, n6975, n6980, n6984, n6988, n6993, n6998, n7003, n7008, n7013, n7017, n7022, n7027, n7032, n7037, n7042, n7047, n7051, n7055, n7060, n7065, n7070, n7075, n7080, n7085, n7089, n7093, n7098, n7103, n7108, n7113, n7118, n7123, n7128, n7132, n7137, n7142, n7147, n7152, n7157, n7162, n7167, n7172, n7177, n7182, n7187, n7192, n7197, n7202, n7207, n7212, n7217, n7221, n7225, n7230, n7234, n7238, n7243, n7248, n7253, n7258, n7263, n7268, n7273, n7278, n7283, n7288, n7293, n7298, n7302, n7306, n7310, n7314, n7319, n7324, n7329, n7333, n7337, n7342, n7347, n7352, n7357, n7362, n7367, n7372, n7377, n7382, n7387, n7392, n7397, n7402, n7407, n7412, n7417, n7422, n7427, n7432, n7437, n7442, n7447, n7452, n7457, n7462, n7467, n7472, n7477, n7481, n7486, n7491, n7496, n7501, n7506, n7511, n7515, n7520, n7525, n7530, n7535, n7540, n7545, n7550, n7555, n7560, n7565, n7570, n7575, n7580, n7585, n7590, n7595, n7600, n7605, n7609, n7613, n7617, n7622, n7627, n7632, n7636, n7641, n7646, n7651, n7656 );
input g1, g58, g86, g341, g194, g215, g191, g79, g121, g316, g218, g392, g405, g160, g429, g401, g319, g324, g475, g457, g59, g433, g153, g146, g164, g150, g157, g355, g351, g142, g298, g301, g182, g174, g168, g344, g347, g441, g437, g446, g111, g102, g424, g411, g417, g93, g671, g650, g645, g110, g74, g637, g255, g246, g239, g262, g225, g283, g71, g63, g305, g513, g667, g65, g655, g499, g43, g112, g12, g370, g385, g376, g358, g85, g55, g51, g568, g604, g50, g550, g94, g49, g534, g586, g613, g48, g542, g577, g617, g47, g546, g582, g46, g590, g626, g52, g199, g599, g45, g595, g538, g632, g518, g7, g31, g6, g8, g28, g9, g19, g16, g34, g482, g66, g22, g25, g37, g35, g36, g6744, g6745, g6746, g6747, g6748, g6749, g6750, g6751, g6752, g6753, g84, g120, g5, g113, g126, g99, g53, g116, g92, g56, g91, g44, g57, g100, g54, g124, g125, g114, g134, g72, g115, g135, g90, g127, g64, g73, g5057, g2771, g1882, g6462, g2299, g4040, g2547, g559, g3017, g3243, g452, g464, g3542, g5232, g5813, g2907, g1744, g5909, g1802, g3554, g6219, g807, g6031, g847, g976, g4172, g4372, g3512, g749, g3490, g6005, g4235, g1600, g1714, g3649, g3155, g3355, g2236, g4555, g3698, g6073, g1736, g1968, g4621, g5607, g2657, g5659, g490, g311, g6069, g772, g5587, g6177, g6377, g3167, g5615, g4567, g3057, g3457, g6287, g1500, g2563, g4776, g4593, g6199, g2295, g1384, g1339, g5180, g2844, g1024, g5591, g3598, g4264, g767, g5853, g3321, g2089, g4933, g4521, g5507, g3625, g6291, g294, g5559, g5794, g6144, g3813, g562, g608, g1205, g3909, g6259, g5905, g921, g2955, g203, g6088, g1099, g4878, g5204, g5630, g3606, g1926, g6215, g3586, g291, g4674, g3570, g640, g5969, g1862, g676, g843, g4132, g4332, g4153, g5666, g6336, g622, g3506, g4558, g6065, g6322, g3111, g117, g2837, g939, g278, g4492, g4864, g1036, g128, g1178, g3239, g718, g6195, g1135, g6137, g6395, g3380, g5343, g554, g496, g3853, g5134, g1422, g3794, g2485, g925, g5555, g878, g1798, g4076, g2941, g3905, g763, g6255, g4375, g4871, g4722, g6692, g1632, g5313, g3100, g1495, g6497, g1437, g6154, g1579, g5567, g1752, g1917, g744, g3040, g4737, g4809, g6267, g3440, g3969, g1442, g5965, g4477, g1233, g4643, g5264, g6329, g2610, g5160, g5360, g5933, g1454, g753, g1296, g3151, g2980, g6727, g3530, g4742, g4104, g1532, g4304, g2177, g3010, g4754, g1189, g2287, g4273, g1389, g1706, g5835, g1171, g4269, g2399, g3372, g4983, g5611, g3618, g4572, g3143, g2898, g3343, g3235, g4543, g3566, g4534, g4961, g6398, g4927, g2259, g2819, g4414, g5802, g2852, g681, g5901, g2886, g3494, g5511, g3518, g1604, g4135, g5092, g4831, g4382, g6386, g479, g3965, g4749, g2008, g736, g3933, g222, g3050, g5736, g1052, g5623, g2122, g2465, g6483, g5889, g4495, g365, g4653, g3179, g1728, g2433, g3835, g6187, g4917, g1070, g822, g6027, g914, g5339, g4164, g969, g2807, g5424, g4054, g6191, g5077, g5523, g3680, g6637, g1682, g1087, g1105, g2342, g6307, g3802, g6159, g2255, g2815, g911, g4012, g1748, g5551, g5742, g3558, g5499, g2960, g3901, g4888, g6251, g6315, g1373, g3092, g2783, g4281, g3574, g2112, g1283, g4297, g5983, g1459, g758, g5712, g4138, g4639, g6537, g5543, g1582, g3736, g5961, g6243, g1227, g3889, g3476, g1664, g1246, g6128, g6629, g4049, g4449, g2932, g4575, g4098, g4498, g528, g5436, g3139, g4584, g5335, g5831, g1216, g2848, g5805, g5022, g4019, g1030, g3672, g3231, g6490, g1430, g4452, g2241, g1564, g5798, g6148, g6649, g884, g3742, g4486, g4504, g5873, g5037, g2319, g5495, g4185, g5208, g2152, g5579, g5869, g5719, g1589, g5752, g6279, g5917, g2975, g6167, g3983, g2599, g1448, g881, g3712, g2370, g5164, g1333, g6549, g4087, g4801, g2984, g3961, g5770, g962, g101, g4226, g6625, g1018, g1418, g4045, g1467, g2461, g5706, g2756, g5990, g471, g1256, g5029, g6519, g4169, g1816, g4369, g3436, g5787, g4578, g4459, g3831, g2514, g3288, g2403, g2145, g1700, g2841, g5297, g3805, g2763, g4793, g952, g1263, g1950, g5138, g2307, g5109, g5791, g3798, g4664, g2223, g5808, g6645, g2016, g5759, g3873, g3632, g2315, g2811, g5957, g2047, g3869, g6358, g3719, g5575, g3752, g3917, g4188, g1585, g4388, g6275, g6311, g4216, g1041, g2595, g2537, g136, g4430, g4564, g3454, g4826, g6239, g3770, g232, g5268, g6545, g2417, g1772, g4741, g5052, g5452, g1890, g2629, g572, g2130, g4108, g4308, g990, g3412, g799, g3706, g3990, g5385, g5881, g1992, g3029, g3171, g3787, g812, g832, g5897, g4165, g4571, g3281, g4455, g2902, g333, g2823, g3684, g3639, g5331, g3338, g5406, g3791, g269, g6040, g5105, g3808, g3759, g4467, g3957, g4093, g1760, g6151, g6351, g5445, g5373, g2279, g3498, g869, g2619, g1183, g1608, g4197, g5283, g1779, g2652, g5459, g2193, g2393, g5767, g661, g4950, g5535, g2834, g1361, g3419, g6235, g1146, g2625, g1696, g6555, g859, g3385, g3881, g6621, g3470, g3897, g3025, g2606, g1472, g6113, g5188, g5689, g1116, g5216, g6494, g4669, g5428, g996, g4531, g2860, g4743, g6593, g2710, g4411, g1413, g4474, g5308, g6641, g3045, g1936, g504, g2587, g4480, g2311, g3602, g5571, g3578, g468, g5448, g3767, g5827, g3582, g6271, g4688, g5774, g2380, g5196, g5396, g3227, g2020, g4000, g1079, g6541, g3203, g1668, g4760, g1840, g70, g5467, g460, g6209, g5290, g3502, g2204, g5256, g4608, g794, g4023, g4423, g3689, g5381, g5685, g703, g5421, g862, g3247, g2040, g4999, g4146, g4633, g1157, g5723, g4732, g5101, g5817, g2151, g2351, g2648, g6736, g4944, g4072, g4443, g3466, g4116, g5041, g5441, g4434, g3827, g6500, g5673, g3133, g3333, g979, g4681, g3774, g2667, g3396, g4210, g1894, g2988, g3538, g827, g1075, g6077, g2555, g5011, g6523, g1526, g4601, g854, g1484, g4922, g5080, g5863, g4581, g3021, g2518, g2567, g3263, g6613, g6044, g6444, g2965, g5857, g1616, g890, g5976, g3562, g4294, g1404, g3723, g3817, g4501, g287, g2724, g4704, g2878, g5220, g1277, g6513, g336, g2882, g933, g1906, g3368, g2799, g887, g5327, g4912, g4157, g2541, g2153, g1945, g5240, g1478, g3080, g3863, g1959, g3480, g6653, g6719, g2864, g4894, g5681, g3857, g3976, g5413, g1002, g776, g1236, g4646, g2476, g1657, g2375, g6012, g896, g967, g3423, g3161, g2384, g3361, g6675, g4616, g4561, g2024, g3451, g2795, g4527, g1844, g5937, g4546, g3103, g2523, g3303, g2643, g6109, g1489, g5390, g2551, g5156, g3072, g1242, g3443, g4277, g1955, g6049, g3034, g2273, g6715, g4771, g6098, g3147, g3347, g2269, g2712, g2729, g5357, g4991, g6019, g4709, g6419, g6052, g2927, g4340, g5929, g4907, g3317, g4035, g2946, g918, g4082, g6486, g2036, g1620, g2831, g930, g3937, g5782, g817, g1249, g837, g3668, g5475, g739, g5949, g6682, g6105, g904, g2873, g1854, g5084, g5603, g4222, g2495, g2437, g2102, g2208, g2579, g4064, g4899, g2719, g4785, g5583, g781, g6173, g6373, g2917, g686, g1252, g2265, g6283, g6369, g5276, g6459, g901, g4194, g5527, g4489, g1974, g1270, g4966, g6415, g6227, g3929, g5503, g4242, g5925, g1124, g4955, g5224, g2012, g6203, g5120, g5320, g2389, g4438, g2429, g2787, g1287, g2675, g4836, g1199, g1399, g5547, g3782, g6428, g2138, g3661, g2338, g4229, g6247, g2791, g3949, g1291, g5945, g5244, g2759, g6741, g785, g1259, g3484, g209, g6609, g5517, g2449, g2575, g2715, g936, g2098, g4462, g6589, g1886, g6466, g6365, g6711, g1870, g4249, g6455, g3004, g1825, g6133, g1008, g4392, g5002, g3546, g5236, g1768, g4854, g3925, g6509, g732, g2504, g1322, g4520, g4219, g2185, g4031, g2070, g4812, g6093, g968, g4176, g4005, g4405, g872, g6181, g6381, g4765, g5563, g1395, g1913, g2331, g6263, g3945, g5731, g4473, g1266, g5489, g714, g2748, g5471, g4540, g6723, g6605, g2445, g2173, g4287, g2491, g4849, g2169, g2283, g6585, g2407, g2868, g2767, g1783, g3310, g1312, g5212, g4245, g4291, g1129, g2227, g6058, g4207, g2246, g1830, g3590, g1592, g6505, g6411, g1221, g5921, g106, g6474, g1932, g1624, g5062, g5462, g2689, g6573, g1677, g2028, g2671, g1576, g4408, g1848, g3089, g3731, g5485, g2741, g802, g2638, g4122, g4322, g5941, g2108, g6000, g1644, g2217, g1319, g2066, g1152, g5252, g2165, g2571, g5176, g5005, g2711, g6023, g1211, g2827, g6423, g875, g4859, g1274, g1426, g2803, g6451, g1821, g2509, g5073, g1280, g4815, g6346, g6633, g5124, g1083, g6303, g5069, g2994, g1636, g3921, g2093, g6732, g1306, g5377, g1061, g3462, g2181, g956, g1756, g5849, g4112, g2685, g2197, g6116, g2421, g1046, g4401, g6434, g1514, g329, g6565, g2950, g4129, g1345, g6533, g3298, g3085, g4727, g6697, g1536, g3941, g5694, g1858, g4932, g3219, g1811, g3431, g6601, g3376, g2441, g1874, g4349, g6581, g6597, g5008, g3610, g2890, g1978, g1612, g2856, g6479, g1982, g6668, g5228, g4119, g6390, g1542, g4258, g4818, g5033, g4717, g1554, g3849, g6704, g3199, g5845, g4975, g790, g5913, g1902, g6163, g4125, g4821, g4939, g1056, g3207, g4483, g3259, g5142, g5248, g2126, g3694, g5481, g1964, g5097, g3215, g4027, g4427, g2779, g4200, g4446, g1720, g1367, g5112, g4145, g2161, g2361, g4191, g2051, g1193, g5401, g3408, g2327, g907, g947, g1834, g3594, g2999, g5727, g2303, g6661, g3065, g699, g723, g5703, g2472, g5953, g3096, g6439, g1740, g3550, g3845, g2116, g5677, g3195, g3913, g4537, g1687, g2681, g2533, g2697, g5747, g4417, g6561, g1141, g1570, g2413, g1710, g6527, g6404, g3255, g1691, g2936, g5644, g5152, g5352, g4213, g6120, g2775, g2922, g1111, g5893, g1311, g3267, g6617, g2060, g4512, g5599, g3401, g4366, g3676, g3129, g3329, g5170, g4456, g5821, g6299, g1239, g3727, g2079, g4698, g3703, g1559, g943, g6140, g3953, g3068, g2704, g6035, g6082, g1300, g4057, g5200, g4843, g5046, g2250, g4549, g2453, g5841, g5763, g3747, g5637, g2912, g2357, g4232, g4253, g5016, g3119, g1351, g1648, g4519, g5115, g3352, g6657, g4552, g3893, g3211, g5654, g929, g3274, g5595, g3614, g2894, g3125, g3325, g3821, g4141, g4570, g5272, g2735, g728, g6295, g5417, g2661, g1988, g5128, g1548, g3106, g4659, g4358, g1792, g2084, g3061, g3187, g4311, g2583, g3003, g1094, g3841, g4284, g3763, g3191, g4239, g3391, g4180, g691, g5366, g2004, g2527, g5456, g4420, g5148, g4507, g5348, g3223, g4931, g2970, g5698, g3416, g5260, g1521, g3522, g3115, g3251, g4628, g1996, g3447, g4515, g4204, g4300, g1724, g1379, g3654, g1878, g5619;
output g7243, g7245, g7257, g7260, g7540, g7916, g7946, g8132, g8178, g8215, g8235, g8277, g8279, g8283, g8291, g8342, g8344, g8353, g8358, g8398, g8403, g8416, g8475, g8719, g8783, g8784, g8785, g8786, g8787, g8788, g8789, g8839, g8870, g8915, g8916, g8917, g8918, g8919, g8920, g9019, g9048, g9251, g9497, g9553, g9555, g9615, g9617, g9680, g9682, g9741, g9743, g9817, g10122, g10306, g10500, g10527, g11349, g11388, g11418, g11447, g11678, g11770, g12184, g12238, g12300, g12350, g12368, g12422, g12470, g12832, g12919, g12923, g13039, g13049, g13068, g13085, g13099, g13259, g13272, g13865, g13881, g13895, g13906, g13926, g13966, g14096, g14125, g14147, g14167, g14189, g14201, g14217, g14421, g14451, g14518, g14597, g14635, g14662, g14673, g14694, g14705, g14738, g14749, g14779, g14828, g16603, g16624, g16627, g16656, g16659, g16686, g16693, g16718, g16722, g16744, g16748, g16775, g16874, g16924, g16955, g17291, g17316, g17320, g17400, g17404, g17423, g17519, g17577, g17580, g17604, g17607, g17639, g17646, g17649, g17674, g17678, g17685, g17688, g17711, g17715, g17722, g17739, g17743, g17760, g17764, g17778, g17787, g17813, g17819, g17845, g17871, g18092, g18094, g18095, g18096, g18097, g18098, g18099, g18100, g18101, g18881, g19334, g19357, g20049, g20557, g20652, g20654, g20763, g20899, g20901, g21176, g21245, g21270, g21292, g21698, g21727, g23002, g23190, g23612, g23652, g23683, g23759, g24151, g25114, g25167, g25219, g25259, g25582, g25583, g25584, g25585, g25586, g25587, g25588, g25589, g25590, g26801, g26875, g26876, g26877, g27831, g28030, g28041, g28042, g28753, g29210, g29211, g29212, g29213, g29214, g29215, g29216, g29217, g29218, g29219, g29220, g29221, g30327, g30329, g30330, g30331, g30332, g31521, g31656, g31665, g31793, g31860, g31861, g31862, g31863, g32185, g32429, g32454, g32975, g33079, g33435, g33533, g33636, g33659, g33874, g33894, g33935, g33945, g33946, g33947, g33948, g33949, g33950, g33959, g34201, g34221, g34232, g34233, g34234, g34235, g34236, g34237, g34238, g34239, g34240, g34383, g34425, g34435, g34436, g34437, g34597, g34788, g34839, g34913, g34915, g34917, g34919, g34921, g34923, g34925, g34927, g34956, g34972, g24168, g24178, g12833, g24174, g24181, g24172, g24161, g24177, g24171, g24163, g24170, g24185, g24164, g24173, g24162, g24179, g24180, g24175, g24183, g24166, g24176, g24184, g24169, g24182, g24165, g24167, n685, n690, n695, n700, n705, n710, n715, n720, n725, n730, n735, n740, n745, n750, n755, n760, n765, n770, n775, n780, n785, n790, n795, n800, n805, n810, n815, n820, n825, n830, n835, n840, n845, n850, n855, n860, n865, n870, n875, n880, n885, n890, n895, n900, n905, n910, n915, n920, n925, n930, n935, n940, n945, n950, n955, n960, n965, n970, n975, n980, n985, n990, n995, n1000, n1005, n1010, n1015, n1020, n1025, n1030, n1035, n1040, n1045, n1050, n1055, n1060, n1065, n1070, n1075, n1080, n1085, n1090, n1094, n1099, n1104, n1109, n1114, n1119, n1124, n1129, n1134, n1139, n1144, n1149, n1154, n1159, n1164, n1169, n1174, n1179, n1184, n1189, n1194, n1199, n1204, n1209, n1214, n1219, n1224, n1229, n1233, n1238, n1243, n1248, n1253, n1258, n1263, n1268, n1273, n1278, n1283, n1288, n1293, n1298, n1303, n1308, n1313, n1318, n1323, n1328, n1333, n1338, n1343, n1348, n1353, n1358, n1363, n1368, n1373, n1378, n1383, n1388, n1393, n1398, n1403, n1408, n1413, n1418, n1423, n1428, n1433, n1438, n1443, n1448, n1453, n1458, n1463, n1468, n1473, n1478, n1483, n1488, n1493, n1498, n1503, n1508, n1513, n1518, n1523, n1528, n1533, n1538, n1543, n1548, n1553, n1558, n1563, n1568, n1573, n1578, n1583, n1588, n1593, n1598, n1603, n1608, n1613, n1618, n1623, n1628, n1633, n1638, n1643, n1648, n1653, n1658, n1663, n1668, n1673, n1678, n1683, n1688, n1693, n1698, n1703, n1708, n1713, n1718, n1723, n1728, n1733, n1738, n1743, n1748, n1753, n1758, n1763, n1768, n1773, n1778, n1783, n1787, n1792, n1797, n1802, n1807, n1812, n1817, n1822, n1827, n1832, n1837, n1842, n1847, n1852, n1856, n1861, n1866, n1871, n1876, n1881, n1886, n1891, n1896, n1901, n1906, n1911, n1916, n1921, n1926, n1931, n1936, n1941, n1946, n1951, n1956, n1961, n1966, n1971, n1976, n1981, n1986, n1991, n1995, n1999, n2004, n2009, n2014, n2019, n2024, n2029, n2034, n2039, n2044, n2049, n2054, n2059, n2064, n2069, n2074, n2078, n2083, n2088, n2093, n2098, n2103, n2108, n2113, n2118, n2123, n2128, n2133, n2138, n2143, n2148, n2153, n2158, n2163, n2168, n2172, n2177, n2182, n2187, n2192, n2197, n2202, n2206, n2211, n2216, n2221, n2226, n2231, n2236, n2241, n2246, n2251, n2255, n2260, n2264, n2269, n2274, n2279, n2284, n2289, n2294, n2299, n2303, n2308, n2313, n2318, n2323, n2328, n2333, n2338, n2342, n2347, n2352, n2357, n2362, n2367, n2372, n2377, n2382, n2387, n2392, n2397, n2402, n2407, n2412, n2417, n2422, n2427, n2432, n2437, n2442, n2447, n2452, n2457, n2462, n2467, n2472, n2476, n2481, n2486, n2491, n2496, n2501, n2506, n2511, n2516, n2521, n2526, n2530, n2535, n2540, n2545, n2550, n2554, n2559, n2564, n2569, n2574, n2579, n2584, n2589, n2594, n2599, n2604, n2609, n2614, n2619, n2624, n2629, n2634, n2639, n2644, n2649, n2654, n2659, n2664, n2669, n2674, n2678, n2683, n2687, n2691, n2696, n2701, n2705, n2710, n2715, n2720, n2725, n2730, n2735, n2740, n2745, n2750, n2755, n2760, n2765, n2770, n2775, n2779, n2784, n2789, n2794, n2799, n2804, n2809, n2814, n2819, n2824, n2829, n2834, n2839, n2844, n2849, n2854, n2859, n2864, n2869, n2874, n2879, n2884, n2889, n2894, n2899, n2904, n2909, n2914, n2919, n2924, n2929, n2934, n2939, n2944, n2949, n2954, n2959, n2964, n2968, n2973, n2978, n2983, n2988, n2993, n2998, n3003, n3008, n3013, n3018, n3023, n3028, n3032, n3036, n3041, n3046, n3051, n3056, n3061, n3066, n3071, n3076, n3081, n3086, n3091, n3096, n3101, n3106, n3111, n3116, n3121, n3126, n3131, n3136, n3141, n3146, n3151, n3156, n3161, n3166, n3171, n3176, n3181, n3186, n3191, n3196, n3201, n3205, n3210, n3215, n3220, n3225, n3230, n3235, n3240, n3245, n3250, n3255, n3260, n3265, n3270, n3275, n3280, n3285, n3290, n3295, n3300, n3304, n3309, n3314, n3319, n3324, n3329, n3334, n3339, n3344, n3348, n3353, n3358, n3363, n3368, n3373, n3378, n3383, n3388, n3393, n3398, n3403, n3408, n3413, n3418, n3422, n3427, n3431, n3436, n3441, n3446, n3451, n3456, n3461, n3466, n3471, n3476, n3481, n3486, n3491, n3496, n3500, n3505, n3510, n3515, n3520, n3525, n3530, n3535, n3540, n3545, n3550, n3555, n3560, n3565, n3570, n3575, n3580, n3584, n3589, n3594, n3599, n3604, n3609, n3614, n3619, n3624, n3629, n3634, n3639, n3644, n3649, n3654, n3659, n3664, n3669, n3674, n3679, n3684, n3689, n3694, n3699, n3704, n3709, n3714, n3718, n3723, n3728, n3732, n3737, n3742, n3747, n3752, n3757, n3762, n3767, n3772, n3777, n3782, n3787, n3792, n3797, n3802, n3807, n3812, n3817, n3822, n3827, n3832, n3837, n3842, n3847, n3852, n3857, n3862, n3866, n3871, n3876, n3881, n3886, n3891, n3896, n3901, n3906, n3911, n3916, n3921, n3925, n3930, n3935, n3940, n3945, n3950, n3955, n3959, n3964, n3969, n3974, n3979, n3984, n3989, n3994, n3999, n4004, n4009, n4014, n4019, n4024, n4029, n4034, n4039, n4043, n4048, n4053, n4058, n4063, n4068, n4073, n4078, n4082, n4087, n4092, n4097, n4102, n4107, n4112, n4117, n4122, n4127, n4132, n4136, n4141, n4146, n4151, n4156, n4161, n4166, n4171, n4176, n4181, n4186, n4191, n4196, n4201, n4205, n4210, n4215, n4220, n4225, n4230, n4235, n4240, n4245, n4250, n4255, n4260, n4265, n4270, n4275, n4280, n4285, n4290, n4295, n4300, n4305, n4310, n4315, n4320, n4325, n4329, n4334, n4339, n4343, n4348, n4353, n4358, n4363, n4368, n4373, n4378, n4383, n4388, n4393, n4398, n4403, n4407, n4412, n4417, n4422, n4427, n4432, n4437, n4442, n4447, n4452, n4457, n4461, n4465, n4469, n4474, n4479, n4484, n4489, n4494, n4499, n4504, n4509, n4514, n4519, n4524, n4529, n4534, n4539, n4544, n4549, n4554, n4558, n4562, n4566, n4571, n4576, n4581, n4586, n4590, n4595, n4600, n4605, n4610, n4615, n4619, n4622, n4627, n4632, n4637, n4642, n4647, n4652, n4657, n4662, n4667, n4672, n4677, n4682, n4687, n4692, n4697, n4702, n4707, n4712, n4717, n4722, n4727, n4731, n4736, n4741, n4746, n4751, n4756, n4761, n4766, n4770, n4775, n4780, n4784, n4788, n4793, n4798, n4803, n4808, n4812, n4817, n4822, n4827, n4832, n4836, n4841, n4846, n4851, n4856, n4861, n4866, n4871, n4876, n4881, n4886, n4891, n4896, n4901, n4906, n4910, n4915, n4920, n4925, n4930, n4934, n4939, n4944, n4949, n4954, n4959, n4964, n4969, n4974, n4979, n4984, n4988, n4992, n4997, n5002, n5007, n5012, n5017, n5022, n5027, n5032, n5037, n5042, n5047, n5051, n5056, n5061, n5066, n5071, n5076, n5081, n5086, n5091, n5096, n5101, n5106, n5111, n5115, n5120, n5125, n5130, n5135, n5140, n5145, n5149, n5153, n5158, n5162, n5166, n5171, n5176, n5181, n5186, n5191, n5196, n5201, n5206, n5211, n5216, n5221, n5226, n5231, n5236, n5241, n5246, n5250, n5254, n5259, n5264, n5269, n5274, n5279, n5284, n5289, n5294, n5299, n5303, n5308, n5313, n5318, n5322, n5326, n5330, n5335, n5340, n5345, n5350, n5355, n5360, n5365, n5370, n5375, n5380, n5385, n5390, n5395, n5400, n5405, n5410, n5415, n5420, n5425, n5430, n5435, n5440, n5445, n5450, n5455, n5460, n5463, n5467, n5472, n5477, n5482, n5487, n5492, n5497, n5502, n5507, n5511, n5516, n5521, n5526, n5531, n5536, n5541, n5546, n5551, n5555, n5560, n5564, n5568, n5573, n5578, n5583, n5587, n5592, n5597, n5602, n5607, n5611, n5615, n5620, n5625, n5630, n5635, n5640, n5645, n5650, n5655, n5660, n5665, n5669, n5674, n5679, n5684, n5689, n5694, n5699, n5704, n5709, n5713, n5718, n5723, n5728, n5733, n5738, n5743, n5748, n5753, n5758, n5763, n5768, n5773, n5778, n5783, n5787, n5792, n5797, n5802, n5807, n5811, n5816, n5821, n5826, n5831, n5836, n5841, n5845, n5850, n5855, n5860, n5865, n5870, n5875, n5880, n5885, n5890, n5895, n5899, n5904, n5909, n5914, n5919, n5924, n5929, n5934, n5939, n5944, n5949, n5954, n5958, n5962, n5967, n5972, n5977, n5982, n5987, n5992, n5996, n6000, n6005, n6010, n6015, n6020, n6024, n6028, n6033, n6038, n6043, n6048, n6053, n6058, n6063, n6068, n6073, n6078, n6083, n6087, n6092, n6096, n6100, n6105, n6110, n6114, n6118, n6123, n6128, n6132, n6136, n6141, n6146, n6151, n6156, n6161, n6166, n6170, n6174, n6178, n6183, n6187, n6191, n6196, n6201, n6206, n6211, n6216, n6221, n6226, n6231, n6236, n6241, n6246, n6251, n6256, n6261, n6266, n6271, n6276, n6281, n6286, n6291, n6296, n6301, n6306, n6311, n6316, n6321, n6326, n6331, n6336, n6341, n6346, n6351, n6355, n6360, n6365, n6369, n6374, n6379, n6384, n6389, n6394, n6399, n6404, n6409, n6414, n6419, n6424, n6429, n6434, n6439, n6444, n6449, n6453, n6458, n6463, n6468, n6473, n6478, n6483, n6488, n6493, n6498, n6502, n6507, n6512, n6517, n6522, n6526, n6531, n6536, n6541, n6546, n6550, n6555, n6560, n6565, n6570, n6575, n6580, n6585, n6590, n6595, n6600, n6605, n6609, n6613, n6618, n6623, n6628, n6633, n6638, n6643, n6648, n6653, n6658, n6662, n6666, n6671, n6676, n6681, n6685, n6690, n6694, n6699, n6703, n6708, n6713, n6718, n6723, n6728, n6733, n6737, n6742, n6747, n6752, n6757, n6762, n6767, n6772, n6777, n6782, n6787, n6792, n6797, n6801, n6805, n6810, n6815, n6820, n6825, n6830, n6835, n6840, n6844, n6849, n6854, n6859, n6864, n6868, n6872, n6877, n6882, n6886, n6891, n6896, n6901, n6906, n6911, n6916, n6921, n6926, n6931, n6935, n6940, n6945, n6950, n6955, n6960, n6965, n6970, n6975, n6980, n6984, n6988, n6993, n6998, n7003, n7008, n7013, n7017, n7022, n7027, n7032, n7037, n7042, n7047, n7051, n7055, n7060, n7065, n7070, n7075, n7080, n7085, n7089, n7093, n7098, n7103, n7108, n7113, n7118, n7123, n7128, n7132, n7137, n7142, n7147, n7152, n7157, n7162, n7167, n7172, n7177, n7182, n7187, n7192, n7197, n7202, n7207, n7212, n7217, n7221, n7225, n7230, n7234, n7238, n7243, n7248, n7253, n7258, n7263, n7268, n7273, n7278, n7283, n7288, n7293, n7298, n7302, n7306, n7310, n7314, n7319, n7324, n7329, n7333, n7337, n7342, n7347, n7352, n7357, n7362, n7367, n7372, n7377, n7382, n7387, n7392, n7397, n7402, n7407, n7412, n7417, n7422, n7427, n7432, n7437, n7442, n7447, n7452, n7457, n7462, n7467, n7472, n7477, n7481, n7486, n7491, n7496, n7501, n7506, n7511, n7515, n7520, n7525, n7530, n7535, n7540, n7545, n7550, n7555, n7560, n7565, n7570, n7575, n7580, n7585, n7590, n7595, n7600, n7605, n7609, n7613, n7617, n7622, n7627, n7632, n7636, n7641, n7646, n7651, n7656;
wire n4620, n4629, n4631, n4642_1, n4643, n4644, n4646, n4647_1, n4649, n4650, n4651, n4652_1, n4653, n4654, n4656, n4657_1, n4658, n4659, n4660, n4661, n4663, n4664, n4665, n4666, n4667_1, n4668, n4670, n4671, n4672_1, n4673, n4674, n4675, n4676, n4677_1, n4678, n4679, n4680, n4681, n4682_1, n4683, n4684, n4685, n4686, n4687_1, n4688, n4689, n4690, n4691, n4692_1, n4693, n4694, n4695, n4696, n4697_1, n4698, n4699, n4700, n4701, n4702_1, n4703, n4704, n4705, n4707_1, n4708, n4709, n4710, n4711, n4712_1, n4713, n4714, n4716, n4717_1, n4719, n4720, n4721, n4722_1, n4723, n4724, n4726, n4727_1, n4728, n4729, n4730, n4731_1, n4732, n4736_1, n4737, n4738, n4739, n4740, n4741_1, n4742, n4743, n4744, n4745, n4746_1, n4747, n4748, n4749, n4750, n4751_1, n4752, n4753, n4754, n4755, n4756_1, n4757, n4758, n4759, n4760, n4761_1, n4762, n4763, n4764, n4765, n4766_1, n4767, n4768, n4769, n4770_1, n4771, n4772, n4773, n4774, n4775_1, n4776, n4777, n4779, n4780_1, n4781, n4782, n4783, n4784_1, n4785, n4786, n4787, n4788_1, n4789, n4790, n4794, n4795, n4796, n4797, n4798_1, n4799, n4800, n4802, n4803_1, n4804, n4805, n4806, n4807, n4809, n4810, n4811, n4812_1, n4813, n4814, n4815, n4816, n4817_1, n4818, n4819, n4820, n4821, n4822_1, n4824, n4825, n4826, n4827_1, n4828, n4829, n4830, n4831, n4832_1, n4833, n4834, n4835, n4836_1, n4837, n4838, n4839, n4840, n4841_1, n4842, n4843, n4844, n4845, n4846_1, n4847, n4848, n4849, n4850, n4851_1, n4852, n4853, n4854, n4855, n4856_1, n4857, n4858, n4859, n4860, n4861_1, n4862, n4863, n4864, n4865, n4866_1, n4867, n4868, n4869, n4870, n4871_1, n4872, n4873, n4874, n4875, n4876_1, n4877, n4879, n4880, n4882, n4883, n4884, n4885, n4886_1, n4888, n4889, n4890, n4891_1, n4892, n4893, n4894, n4895, n4896_1, n4897, n4898, n4899, n4900, n4908, n4909, n4910_1, n4911, n4912, n4913, n4914, n4915_1, n4916, n4917, n4918, n4919, n4920_1, n4921, n4922, n4923, n4924, n4925_1, n4926, n4927, n4928, n4929, n4930_1, n4931, n4932, n4933, n4934_1, n4935, n4936, n4937, n4938, n4939_1, n4940, n4941, n4942, n4943, n4944_1, n4945, n4946, n4947, n4949_1, n4950, n4951, n4952, n4953, n4954_1, n4955, n4956, n4957, n4958, n4959_1, n4960, n4961, n4962, n4963, n4964_1, n4965, n4966, n4967, n4968, n4969_1, n4970, n4971, n4972, n4973, n4976, n4977, n4979_1, n4980, n4981, n4982, n4983, n4984_1, n4985, n4986, n4987, n4988_1, n4989, n4990, n4991, n4992_1, n4993, n4994, n4995, n4996, n4997_1, n4998, n4999, n5000, n5001, n5002_1, n5003, n5004, n5005, n5006, n5007_1, n5008, n5009, n5010, n5011, n5012_1, n5013, n5014, n5015, n5016, n5017_1, n5018, n5019, n5020, n5021, n5022_1, n5023, n5024, n5025, n5026, n5027_1, n5028, n5029, n5030, n5031, n5032_1, n5033, n5034, n5035, n5036, n5037_1, n5038, n5039, n5040, n5041, n5042_1, n5043, n5044, n5045, n5046, n5047_1, n5048, n5049, n5050, n5051_1, n5052, n5053, n5054, n5055, n5056_1, n5057, n5058, n5059, n5060, n5061_1, n5062, n5066_1, n5067, n5068, n5072, n5073, n5074, n5076_1, n5077, n5078, n5079, n5081_1, n5082, n5083, n5085, n5086_1, n5087, n5088, n5089, n5090, n5091_1, n5092, n5093, n5094, n5095, n5096_1, n5097, n5098, n5099, n5100, n5102, n5103, n5104, n5105, n5106_1, n5107, n5110, n5113, n5114, n5115_1, n5116, n5117, n5118, n5120_1, n5121, n5122, n5123, n5124, n5125_1, n5126, n5127, n5129, n5130_1, n5131, n5132, n5133, n5134, n5135_1, n5136, n5137, n5138, n5139, n5140_1, n5141, n5142, n5143, n5144, n5145_1, n5146, n5147, n5148, n5149_1, n5150, n5151, n5152, n5153_1, n5154, n5155, n5156, n5157, n5158_1, n5159, n5160, n5161, n5162_1, n5163, n5164, n5165, n5166_1, n5167, n5168, n5169, n5170, n5173, n5174, n5175, n5176_1, n5177, n5178, n5179, n5180, n5181_1, n5182, n5183, n5184, n5185, n5186_1, n5187, n5188, n5189, n5190, n5191_1, n5192, n5193, n5194, n5195, n5196_1, n5197, n5198, n5199, n5202, n5203, n5204, n5205, n5207, n5215, n5216_1, n5217, n5218, n5219, n5220, n5221_1, n5222, n5223, n5224, n5225, n5226_1, n5227, n5228, n5229, n5230, n5231_1, n5232, n5233, n5234, n5235, n5236_1, n5237, n5238, n5239, n5240, n5241_1, n5242, n5243, n5244, n5245, n5246_1, n5247, n5248, n5250_1, n5251, n5252, n5253, n5254_1, n5255, n5256, n5257, n5258, n5259_1, n5260, n5261, n5262, n5263, n5264_1, n5265, n5266, n5267, n5268, n5269_1, n5270, n5271, n5272, n5273, n5274_1, n5275, n5276, n5277, n5278, n5279_1, n5280, n5282, n5283, n5284_1, n5285, n5286, n5287, n5288, n5289_1, n5290, n5291, n5292, n5293, n5294_1, n5295, n5296, n5297, n5298, n5299_1, n5300, n5301, n5302, n5303_1, n5304, n5305, n5306, n5307, n5308_1, n5310, n5311, n5312, n5313_1, n5314, n5315, n5316, n5317, n5318_1, n5319, n5320, n5321, n5322_1, n5323, n5324, n5325, n5326_1, n5327, n5328, n5329, n5330_1, n5331, n5332, n5333, n5334, n5335_1, n5336, n5337, n5339, n5340_1, n5341, n5342, n5343, n5344, n5345_1, n5346, n5347, n5348, n5349, n5350_1, n5351, n5352, n5353, n5354, n5355_1, n5356, n5357, n5358, n5359, n5360_1, n5361, n5362, n5363, n5364, n5365_1, n5366, n5367, n5368, n5370_1, n5371, n5372, n5373, n5374, n5375_1, n5376, n5377, n5378, n5379, n5380_1, n5381, n5382, n5383, n5384, n5385_1, n5386, n5387, n5388, n5389, n5390_1, n5391, n5392, n5393, n5394, n5395_1, n5396, n5397, n5398, n5399, n5401, n5402, n5403, n5404, n5405_1, n5406, n5407, n5408, n5409, n5410_1, n5411, n5412, n5413, n5414, n5415_1, n5416, n5417, n5418, n5419, n5420_1, n5421, n5422, n5423, n5424, n5425_1, n5428, n5429, n5430_1, n5431, n5432, n5433, n5434, n5435_1, n5436, n5437, n5438, n5439, n5440_1, n5441, n5442, n5443, n5444, n5445_1, n5446, n5447, n5448, n5449, n5450_1, n5451, n5452, n5453, n5454, n5455_1, n5456, n5457, n5461, n5462, n5463_1, n5464, n5465, n5466, n5468, n5469, n5470, n5471, n5472_1, n5476, n5477_1, n5478, n5479, n5480, n5481, n5482_1, n5483, n5484, n5485, n5486, n5487_1, n5488, n5489, n5490, n5491, n5492_1, n5493, n5494, n5495, n5496, n5497_1, n5498, n5499, n5500, n5501, n5502_1, n5503, n5505, n5506, n5507_1, n5508, n5509, n5510, n5511_1, n5512, n5513, n5514, n5516_1, n5517, n5518, n5519, n5520, n5521_1, n5522, n5523, n5524, n5525, n5526_1, n5527, n5528, n5529, n5530, n5531_1, n5532, n5533, n5535, n5536_1, n5537, n5538, n5540, n5541_1, n5542, n5543, n5544, n5545, n5546_1, n5547, n5548, n5549, n5550, n5551_1, n5552, n5553, n5554, n5556, n5557, n5558, n5559, n5560_1, n5562, n5563, n5564_1, n5565, n5566, n5567, n5568_1, n5569, n5570, n5571, n5573_1, n5574, n5575, n5576, n5577, n5578_1, n5579, n5580, n5581, n5582, n5583_1, n5584, n5585, n5586, n5587_1, n5588, n5589, n5591, n5592_1, n5593, n5594, n5595, n5596, n5598, n5599, n5600, n5601, n5602_1, n5604, n5606, n5607_1, n5608, n5610, n5611_1, n5612, n5614, n5616, n5617, n5618, n5620_1, n5621, n5622, n5623, n5624, n5625_1, n5626, n5627, n5628, n5629, n5630_1, n5632, n5633, n5634, n5636, n5637, n5638, n5639, n5640_1, n5642, n5643, n5645_1, n5646, n5647, n5648, n5649, n5651, n5652, n5653, n5654, n5655_1, n5656, n5657, n5658, n5659, n5660_1, n5661, n5662, n5663, n5664, n5665_1, n5666, n5667, n5668, n5669_1, n5670, n5671, n5672, n5673, n5674_1, n5675, n5676, n5677, n5678, n5679_1, n5680, n5681, n5682, n5683, n5684_1, n5685, n5687, n5688, n5689_1, n5691, n5692, n5693, n5694_1, n5697, n5698, n5700, n5701, n5702, n5703, n5704_1, n5705, n5706, n5707, n5708, n5709_1, n5710, n5711, n5712, n5713_1, n5714, n5715, n5716, n5717, n5718_1, n5719, n5720, n5721, n5722, n5723_1, n5724, n5725, n5726, n5727, n5728_1, n5729, n5730, n5732, n5733_1, n5734, n5735, n5736, n5737, n5739, n5741, n5743_1, n5744, n5745, n5746, n5747, n5748_1, n5749, n5750, n5752, n5753_1, n5754, n5755, n5756, n5757, n5758_1, n5759, n5760, n5762, n5763_1, n5765, n5767, n5768_1, n5769, n5770, n5771, n5772, n5773_1, n5774, n5775, n5776, n5777, n5778_1, n5779, n5780, n5781, n5782, n5783_1, n5785, n5786, n5787_1, n5788, n5789, n5790, n5791, n5792_1, n5793, n5794, n5795, n5796, n5797_1, n5798, n5799, n5800, n5802_1, n5803, n5804, n5805, n5806, n5807_1, n5809, n5810, n5811_1, n5812, n5813, n5814, n5815, n5816_1, n5817, n5818, n5819, n5820, n5821_1, n5822, n5823, n5824, n5825, n5826_1, n5827, n5828, n5829, n5830, n5831_1, n5832, n5834, n5835, n5836_1, n5838, n5839, n5840, n5841_1, n5842, n5844, n5845_1, n5846, n5847, n5848, n5849, n5850_1, n5851, n5852, n5854, n5855_1, n5856, n5857, n5859, n5860_1, n5861, n5862, n5863, n5864, n5865_1, n5867, n5868, n5869, n5870_1, n5871, n5872, n5873, n5874, n5876, n5877, n5878, n5879, n5880_1, n5881, n5882, n5883, n5884, n5885_1, n5886, n5889, n5890_1, n5891, n5892, n5893, n5894, n5896, n5897, n5899_1, n5900, n5901, n5903, n5904_1, n5905, n5906, n5907, n5908, n5909_1, n5910, n5911, n5913, n5914_1, n5916, n5917, n5918, n5920, n5921, n5922, n5924_1, n5925, n5927, n5928, n5929_1, n5930, n5931, n5932, n5933, n5934_1, n5935, n5936, n5937, n5938, n5939_1, n5940, n5941, n5942, n5943, n5944_1, n5945, n5946, n5947, n5948, n5949_1, n5950, n5951, n5952, n5953, n5954_1, n5955, n5956, n5957, n5958_1, n5959, n5960, n5961, n5962_1, n5963, n5964, n5965, n5966, n5967_1, n5968, n5969, n5970, n5971, n5972_1, n5973, n5974, n5975, n5976, n5977_1, n5978, n5980, n5981, n5982_1, n5984, n5985, n5986, n5987_1, n5988, n5989, n5990, n5991, n5993, n5994, n5995, n5996_1, n5997, n5998, n5999, n6000_1, n6001, n6002, n6003, n6004, n6005_1, n6007, n6008, n6009, n6010_1, n6011, n6012, n6013, n6014, n6015_1, n6016, n6018, n6019, n6020_1, n6021, n6022, n6023, n6024_1, n6025, n6026, n6027, n6029, n6030, n6032, n6033_1, n6034, n6036, n6037, n6038_1, n6039, n6042, n6043_1, n6044, n6045, n6047, n6049, n6050, n6051, n6052, n6053_1, n6054, n6055, n6056, n6057, n6058_1, n6059, n6060, n6061, n6062, n6064, n6065, n6067, n6068_1, n6069, n6071, n6073_1, n6074, n6077, n6079, n6080, n6081, n6082, n6083_1, n6084, n6085, n6086, n6087_1, n6089, n6090, n6091, n6092_1, n6094, n6097, n6099, n6100_1, n6101, n6103, n6104, n6105_1, n6106, n6107, n6108, n6109, n6110_1, n6111, n6112, n6113, n6114_1, n6115, n6116, n6117, n6118_1, n6119, n6120, n6121, n6122, n6124, n6125, n6129, n6131, n6132_1, n6133, n6134, n6135, n6136_1, n6137, n6138, n6140, n6141_1, n6142, n6143, n6144, n6145, n6146_1, n6147, n6148, n6150, n6152, n6153, n6154, n6156_1, n6157, n6159, n6160, n6162, n6163, n6164, n6165, n6167, n6168, n6169, n6170_1, n6171, n6172, n6173, n6174_1, n6175, n6177, n6178_1, n6180, n6181, n6182, n6183_1, n6184, n6185, n6186, n6188, n6189, n6190, n6192, n6193, n6195, n6196_1, n6197, n6199, n6200, n6202, n6203, n6204, n6205, n6206_1, n6208, n6209, n6211_1, n6212, n6214, n6216_1, n6218, n6219, n6221_1, n6222, n6223, n6224, n6225, n6227, n6228, n6229, n6230, n6231_1, n6232, n6233, n6234, n6235, n6236_1, n6237, n6238, n6239, n6240, n6241_1, n6242, n6243, n6245, n6246_1, n6247, n6248, n6249, n6250, n6252, n6253, n6254, n6256_1, n6257, n6258, n6259, n6260, n6261_1, n6263, n6264, n6265, n6266_1, n6267, n6268, n6269, n6270, n6271_1, n6272, n6273, n6275, n6276_1, n6277, n6278, n6279, n6280, n6281_1, n6282, n6284, n6285, n6286_1, n6287, n6288, n6292, n6293, n6294, n6295, n6297, n6299, n6300, n6301_1, n6302, n6303, n6304, n6305, n6306_1, n6307, n6308, n6309, n6310, n6311_1, n6312, n6313, n6316_1, n6317, n6318, n6319, n6320, n6322, n6323, n6326_1, n6328, n6329, n6330, n6331_1, n6333, n6334, n6335, n6336_1, n6337, n6338, n6339, n6340, n6341_1, n6342, n6343, n6344, n6345, n6346_1, n6347, n6348, n6349, n6350, n6351_1, n6352, n6353, n6354, n6355_1, n6356, n6357, n6358, n6359, n6360_1, n6361, n6362, n6363, n6364, n6365_1, n6366, n6367, n6368, n6369_1, n6370, n6371, n6372, n6373, n6374_1, n6375, n6376, n6377, n6378, n6380, n6382, n6383, n6385, n6386, n6387, n6388, n6389_1, n6390, n6392, n6393, n6394_1, n6396, n6397, n6398, n6399_1, n6400, n6402, n6403, n6404_1, n6406, n6407, n6409_1, n6410, n6411, n6412, n6413, n6414_1, n6415, n6416, n6417, n6418, n6419_1, n6421, n6422, n6424_1, n6425, n6426, n6428, n6429_1, n6430, n6431, n6432, n6433, n6435, n6436, n6438, n6439_1, n6440, n6441, n6444_1, n6445, n6446, n6447, n6449_1, n6450, n6451, n6452, n6453_1, n6454, n6455, n6456, n6457, n6459, n6460, n6462, n6463_1, n6464, n6466, n6467, n6468_1, n6469, n6470, n6471, n6472, n6474, n6475, n6476, n6478_1, n6479, n6480, n6482, n6483_1, n6485, n6487, n6488_1, n6491, n6494, n6495, n6497, n6498_1, n6500, n6501, n6502_1, n6503, n6505, n6506, n6507_1, n6508, n6509, n6510, n6511, n6513, n6514, n6515, n6517_1, n6518, n6519, n6520, n6521, n6522_1, n6523, n6524, n6526_1, n6527, n6528, n6529, n6530, n6531_1, n6532, n6533, n6534, n6535, n6536_1, n6537, n6538, n6539, n6540, n6541_1, n6542, n6543, n6544, n6545, n6546_1, n6547, n6548, n6549, n6550_1, n6551, n6552, n6553, n6554, n6555_1, n6556, n6557, n6558, n6559, n6560_1, n6561, n6562, n6563, n6564, n6565_1, n6566, n6567, n6568, n6569, n6570_1, n6571, n6572, n6574, n6575_1, n6577, n6578, n6579, n6581, n6582, n6584, n6585_1, n6587, n6588, n6589, n6590_1, n6591, n6592, n6593, n6594, n6595_1, n6596, n6597, n6598, n6599, n6601, n6604, n6605_1, n6607, n6608, n6609_1, n6611, n6614, n6616, n6617, n6619, n6621, n6622, n6624, n6625, n6626, n6628_1, n6629, n6630, n6631, n6633_1, n6635, n6636, n6637, n6638_1, n6639, n6640, n6641, n6642, n6643_1, n6644, n6645, n6646, n6647, n6648_1, n6649, n6650, n6651, n6653_1, n6654, n6655, n6656, n6658_1, n6659, n6660, n6661, n6662_1, n6664, n6665, n6667, n6668, n6669, n6670, n6672, n6674, n6675, n6676_1, n6678, n6679, n6680, n6681_1, n6682, n6684, n6685_1, n6686, n6689, n6690_1, n6691, n6692, n6693, n6695, n6697, n6698, n6700, n6701, n6702, n6703_1, n6704, n6705, n6706, n6707, n6708_1, n6709, n6710, n6711, n6713_1, n6714, n6715, n6717, n6718_1, n6720, n6721, n6722, n6723_1, n6724, n6726, n6728_1, n6729, n6730, n6731, n6732, n6734, n6735, n6736, n6738, n6739, n6740, n6742_1, n6744, n6745, n6746, n6747_1, n6748, n6749, n6750, n6752_1, n6753, n6754, n6755, n6756, n6757_1, n6758, n6759, n6760, n6761, n6762_1, n6763, n6765, n6768, n6770, n6771, n6772_1, n6773, n6774, n6775, n6777_1, n6778, n6779, n6780, n6781, n6782_1, n6783, n6785, n6786, n6788, n6789, n6790, n6791, n6792_1, n6793, n6794, n6795, n6796, n6797_1, n6798, n6799, n6800, n6801_1, n6802, n6803, n6804, n6805_1, n6806, n6807, n6808, n6809, n6810_1, n6811, n6812, n6813, n6814, n6816, n6817, n6818, n6820_1, n6821, n6822, n6824, n6825_1, n6826, n6827, n6828, n6829, n6830_1, n6832, n6833, n6835_1, n6836, n6837, n6839, n6840_1, n6842, n6843, n6844_1, n6845, n6846, n6847, n6848, n6849_1, n6850, n6851, n6853, n6854_1, n6855, n6856, n6857, n6858, n6859_1, n6860, n6861, n6862, n6863, n6864_1, n6865, n6866, n6867, n6868_1, n6869, n6870, n6871, n6873, n6874, n6875, n6876, n6877_1, n6878, n6879, n6880, n6881, n6882_1, n6883, n6884, n6885, n6886_1, n6887, n6888, n6889, n6891_1, n6892, n6894, n6895, n6897, n6898, n6899, n6900, n6901_1, n6902, n6903, n6905, n6906_1, n6907, n6908, n6910, n6912, n6914, n6916_1, n6918, n6919, n6921_1, n6922, n6924, n6925, n6926_1, n6928, n6929, n6930, n6932, n6934, n6937, n6939, n6940_1, n6942, n6944, n6945_1, n6946, n6947, n6948, n6949, n6950_1, n6951, n6952, n6953, n6954, n6955_1, n6956, n6957, n6958, n6959, n6960_1, n6961, n6962, n6963, n6964, n6965_1, n6966, n6967, n6968, n6969, n6970_1, n6971, n6972, n6973, n6974, n6975_1, n6976, n6977, n6978, n6979, n6980_1, n6981, n6982, n6983, n6984_1, n6985, n6986, n6987, n6988_1, n6989, n6991, n6992, n6993_1, n6995, n6996, n6997, n6998_1, n6999, n7000, n7001, n7003_1, n7004, n7005, n7006, n7007, n7008_1, n7011, n7013_1, n7014, n7015, n7016, n7017_1, n7018, n7019, n7020, n7021, n7022_1, n7023, n7024, n7025, n7026, n7027_1, n7028, n7029, n7030, n7031, n7032_1, n7033, n7035, n7036, n7037_1, n7039, n7041, n7042_1, n7043, n7044, n7046, n7047_1, n7048, n7049, n7050, n7052, n7053, n7054, n7056, n7057, n7058, n7059, n7060_1, n7061, n7062, n7063, n7064, n7065_1, n7066, n7067, n7068, n7069, n7070_1, n7071, n7072, n7073, n7074, n7075_1, n7076, n7077, n7078, n7079, n7081, n7082, n7083, n7084, n7085_1, n7088, n7089_1, n7090, n7091, n7092, n7094, n7095, n7096, n7097, n7098_1, n7099, n7100, n7101, n7102, n7103_1, n7104, n7106, n7107, n7108_1, n7110, n7111, n7113_1, n7114, n7115, n7118_1, n7119, n7120, n7121, n7123_1, n7124, n7125, n7127, n7128_1, n7129, n7131, n7132_1, n7133, n7134, n7136, n7137_1, n7138, n7140, n7142_1, n7144, n7145, n7146, n7147_1, n7148, n7149, n7150, n7151, n7153, n7154, n7155, n7156, n7157_1, n7158, n7159, n7160, n7161, n7162_1, n7164, n7165, n7166, n7167_1, n7168, n7171, n7172_1, n7173, n7174, n7175, n7176, n7178, n7179, n7180, n7181, n7182_1, n7184, n7185, n7186, n7187_1, n7189, n7190, n7191, n7192_1, n7193, n7195, n7196, n7197_1, n7199, n7200, n7202_1, n7204, n7205, n7206, n7207_1, n7209, n7211, n7212_1, n7213, n7214, n7215, n7216, n7218, n7219, n7220, n7222, n7223, n7224, n7226, n7227, n7228, n7229, n7230_1, n7232, n7233, n7235, n7237, n7238_1, n7239, n7241, n7242, n7243_1, n7244, n7245, n7247, n7248_1, n7249, n7251, n7253_1, n7254, n7256, n7257, n7259, n7260, n7261, n7263_1, n7264, n7266, n7267, n7268_1, n7270, n7272, n7273_1, n7275, n7276, n7277, n7279, n7280, n7282, n7283_1, n7284, n7285, n7286, n7287, n7288_1, n7289, n7290, n7291, n7292, n7295, n7296, n7297, n7298_1, n7299, n7300, n7301, n7302_1, n7303, n7304, n7305, n7306_1, n7307, n7308, n7309, n7310_1, n7311, n7313, n7314_1, n7315, n7317, n7318, n7320, n7321, n7322, n7324_1, n7325, n7326, n7328, n7330, n7331, n7333_1, n7334, n7335, n7337_1, n7338, n7339, n7341, n7343, n7344, n7345, n7347_1, n7348, n7350, n7351, n7352_1, n7353, n7354, n7355, n7356, n7357_1, n7358, n7359, n7360, n7361, n7362_1, n7363, n7364, n7365, n7366, n7367_1, n7368, n7369, n7370, n7371, n7372_1, n7373, n7375, n7376, n7377_1, n7379, n7380, n7381, n7383, n7384, n7385, n7386, n7389, n7390, n7392_1, n7393, n7394, n7396, n7397_1, n7398, n7399, n7400, n7403, n7405, n7406, n7408, n7409, n7411, n7412_1, n7414, n7415, n7416, n7417_1, n7420, n7421, n7422_1, n7423, n7424, n7425, n7426, n7427_1, n7428, n7429, n7430, n7431, n7432_1, n7433, n7434, n7435, n7436, n7437_1, n7438, n7439, n7440, n7441, n7442_1, n7443, n7445, n7446, n7448, n7449, n7451, n7452_1, n7454, n7455, n7456, n7457_1, n7458, n7460, n7462_1, n7464, n7465, n7466, n7467_1, n7468, n7469, n7471, n7472_1, n7473, n7474, n7476, n7477_1, n7478, n7480, n7481_1, n7482, n7484, n7486_1, n7487, n7488, n7489, n7490, n7491_1, n7493, n7494, n7495, n7496_1, n7498, n7499, n7500, n7502, n7503, n7504, n7506_1, n7507, n7508, n7511_1, n7512, n7513, n7514, n7515_1, n7516, n7517, n7518, n7520_1, n7521, n7524, n7525_1, n7526, n7528, n7530_1, n7531, n7532, n7534, n7537, n7538, n7540_1, n7541, n7542, n7543, n7545_1, n7546, n7547, n7548, n7549, n7551, n7552, n7553, n7554, n7556, n7558, n7559, n7561, n7562, n7563, n7566, n7567, n7569, n7571, n7572, n7573, n7574, n7577, n7578, n7579, n7581, n7582, n7584, n7585_1, n7587, n7588, n7589, n7590_1, n7591, n7593, n7595_1, n7596, n7597, n7598, n7599, n7601, n7602, n7603, n7604, n7605_1, n7606, n7608, n7609_1, n7610, n7612, n7613_1, n7614, n7615, n7616, n7617_1, n7618, n7619, n7620, n7621, n7624, n7626, n7628, n7629, n7630, n7632_1, n7633, n7634, n7635, n7637, n7638, n7639, n7640, n7642, n7643, n7644, n7646_1, n7647, n7648, n7649, n7651_1, n7652, n7654, n7655, n7657, n7658, n7659, n7661, n7662, n7664, n7666, n7667, n7668, n7669, n7670, n7671, n7673, n7675, n7676, n7677, n7678, n7679, n7681, n7682, n7683, n7684, n7686, n7687, n7688, n7690, n7692, n7693, n7694, n7695, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7705, n7707, n7708, n7709, n7710, n7711, n7712, n7714, n7715, n7716, n7717, n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7727, n7728, n7730, n7731, n7732, n7733, n7736, n7738, n7739, n7741, n7743, n7744, n7745, n7746, n7748, n7749, n7750, n7753, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7766, n7767, n7768, n7770, n7772, n7773, n7774, n7776, n7777, n7779, n7780, n7782, n7783, n7784, n7785, n7787, n7788, n7789, n7791, n7792, n7793, n7794, n7796, n7797, n7799, n7800, n7801, n7802, n7803, n7805, n7806, n7807, n7808, n7809, n7811, n7812, n7813, n7815, n7816, n7818, n7819, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7831, n7832, n7833, n7835, n7836, n7837, n7839, n7840, n7842, n7843, n7844, n7846, n7847, n7849, n7850, n7851, n7852, n7854, n7855, n7857, n7858, n7859, n7860, n7861, n7863, n7864, n7866, n7867, n7868, n7870, n7872, n7873, n7874, n7875, n7877, n7878, n7880, n7881, n7883, n7884, n7885, n7887, n7888, n7890, n7891, n7892, n7894, n7895, n7898, n7900, n7901, n7902, n7904, n7905, n7906, n7908, n7909, n7910, n7912, n7913, n7915, n7916, n7917, n7920, n7922, n7923, n7924, n7926, n7927, n7928, n7929, n7931, n7933, n7934, n7935, n7937, n7939, n7940, n7941, n7942, n7944, n7945, n7948, n7949, n7950, n7953, n7954, n7956, n7957, n7959, n7961, n7963, n7964, n7965, n7967, n7970, n7971, n7974, n7975, n7976, n7978, n7979, n7980, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7994, n7995, n7996, n7998, n7999, n8000, n8002, n8003, n8004, n8005, n8006, n8007, n8009, n8010, n8011, n8013, n8014, n8016, n8017, n8018, n8019, n8020, n8022, n8023, n8024, n8026, n8027, n8029, n8030, n8032, n8033, n8034, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8044, n8046, n8047, n8049, n8051, n8052, n8053, n8054, n8055, n8057, n8058, n8060, n8061, n8062, n8064, n8065, n8067, n8069, n8071, n8072, n8073, n8075, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8121, n8122, n8124, n8125, n8126, n8128, n8129, n8131, n8132, n8134, n8135, n8136, n8137, n8138, n8140, n8141, n8142, n8144, n8145, n8146, n8147, n8149, n8150, n8151, n8153, n8154, n8155, n8156, n8158, n8160, n8161, n8162, n8164, n8165, n8167, n8168, n8170, n8171, n8172, n8173, n8175, n8176, n8177, n8179, n8180, n8181, n8183, n8184, n8185, n8186, n8188, n8189, n8191, n8193, n8194, n8196, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8208, n8209, n8210, n8213, n8214, n8216, n8217, n8218, n8219, n8221, n8222, n8224, n8225, n8226, n8228, n8229, n8230, n8231, n8233, n8234, n8235, n8237, n8238, n8239, n8241, n8242, n8243, n8246, n8247, n8248, n8249, n8250, n8252, n8253, n8254, n8256, n8257, n8259, n8261, n8262, n8264, n8265, n8267, n8268, n8269, n8271, n8273, n8274, n8275, n8277, n8278, n8279, n8281, n8282, n8284, n8286, n8287, n8288, n8290, n8292, n8294, n8295, n8297, n8298, n8299, n8300, n8301, n8303, n8304, n8305, n8306, n8309, n8310, n8311, n8313, n8315, n8316, n8317, n8319, n8320, n8321, n8324, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8343, n8344, n8346, n8347, n8348, n8350, n8351, n8353, n8354, n8356, n8357, n8359, n8360, n8361, n8363, n8364, n8366, n8367, n8368, n8370, n8371, n8373, n8374, n8376, n8377, n8379, n8382, n8383, n8385, n8387, n8388, n8390, n8391, n8394, n8395, n8396, n8398, n8400, n8401, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8411, n8412, n8414, n8415, n8416, n8418, n8419, n8420, n8422, n8423, n8425, n8426, n8427, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8440, n8442, n8443, n8445, n8447, n8449, n8450, n8451, n8453, n8454, n8455, n8457, n8459, n8461, n8462, n8463, n8465, n8466, n8468, n8469, n8470, n8471, n8472, n8474, n8476, n8477, n8479, n8480, n8481, n8483, n8484, n8485, n8486, n8487, n8489, n8491, n8493, n8494, n8496, n8497, n8498, n8499, n8500, n8502, n8504, n8505, n8506, n8507, n8508, n8510, n8511, n8512, n8513, n8514, n8516, n8517, n8518, n8519, n8520, n8521, n8523, n8526, n8527, n8530, n8531, n8533, n8534, n8536, n8537, n8538, n8540, n8541, n8542, n8544, n8545, n8546, n8547, n8548, n8551, n8552, n8554, n8556, n8557, n8558, n8559, n8561, n8563, n8564, n8565, n8567, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8617, n8618, n8619, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8666, n8667, n8669, n8670, n8671, n8673, n8675, n8676, n8677, n8678, n8679, n8680, n8682, n8683, n8684, n8686, n8687, n8689, n8690, n8694, n8695, n8696, n8697, n8698, n8700, n8701, n8703, n8704, n8705, n8706, n8708, n8709, n8710, n8712, n8714, n8715, n8717, n8718, n8719, n8721, n8722, n8723, n8724, n8726, n8727, n8728, n8729, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8758, n8760, n8761, n8762, n8763, n8765, n8766, n8767, n8769, n8770, n8772, n8773, n8774, n8775, n8776, n8777, n8779, n8780, n8781, n8782, n8785, n8787, n8788, n8789, n8792, n8794, n8795, n8798, n8799, n8800, n8802, n8803, n8804, n8805, n8808, n8809, n8811, n8812, n8813, n8814, n8815, n8816, n8818, n8819, n8821, n8822, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8834, n8835, n8836, n8837, n8838, n8839, n8841, n8842, n8844, n8845, n8847, n8848, n8850, n8851, n8853, n8854, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8866, n8867, n8869, n8870, n8872, n8876, n8877, n8878, n8880, n8882, n8884, n8885, n8886, n8888, n8889, n8890, n8892, n8893, n8894, n8897, n8898, n8899, n8900, n8902, n8903, n8904, n8906, n8908, n8910, n8912, n8913, n8914, n8915, n8917, n8918, n8919, n8921, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8934, n8935, n8937, n8938, n8939, n8941, n8943, n8944, n8945, n8947, n8948, n8949, n8950, n8952, n8953, n8954, n8956, n8957, n8959, n8960, n8961, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8975, n8976, n8977, n8979, n8980, n8982, n8984, n8985, n8987, n8989, n8990, n8992, n8993, n8994, n8996, n8997, n8998, n8999, n9000, n9002, n9004, n9007, n9008, n9009, n9010, n9012, n9013, n9015, n9016, n9017, n9019, n9020, n9021, n9022, n9024, n9025, n9026, n9028, n9029, n9030, n9031, n9032, n9035, n9036, n9038, n9039, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9049, n9050, n9051, n9052, n9054, n9055, n9056, n9058, n9059, n9061, n9062, n9064, n9065, n9066, n9068, n9069, n9070, n9071, n9073, n9074, n9075, n9076, n9077, n9080, n9081, n9083, n9084, n9085, n9087, n9088, n9089, n9091, n9092, n9093, n9095, n9096, n9097, n9099, n9100, n9101, n9102, n9103, n9104, n9106, n9107, n9110, n9112, n9113, n9115, n9116, n9118, n9119, n9120, n9122, n9123, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9136, n9137, n9138, n9140, n9141, n9142, n9144, n9146, n9147, n9148, n9150, n9152, n9153, n9155, n9156, n9157, n9159, n9160, n9161, n9163, n9164, n9165, n9166, n9167, n9169, n9170, n9171, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9184, n9185, n9186, n9188, n9189, n9190, n9191, n9193, n9194, n9195, n9197, n9198, n9200, n9202, n9204, n9206, n9207, n9208, n9210, n9211, n9212, n9215, n9216, n9217, n9219, n9220, n9222, n9223, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9240, n9242, n9243, n9245, n9246, n9248, n9250, n9251, n9252, n9255, n9256, n9257, n9258, n9259, n9260, n9262, n9263, n9265, n9267, n9268, n9269, n9271, n9272, n9274, n9275, n9276, n9277, n9278, n9279, n9281, n9282, n9285, n9287, n9288, n9289, n9291, n9292, n9293, n9295, n9296, n9298, n9299, n9301, n9302, n9304, n9306, n9307, n9309, n9310, n9312, n9314, n9315, n9316, n9318, n9320, n9321, n9322, n9324, n9325, n9327, n9328, n9329, n9331, n9333, n9334, n9335, n9336, n9338, n9339, n9341, n9342, n9344, n9345, n9346, n9347, n9349, n9351, n9352, n9354, n9355, n9358, n9359, n9360, n9363, n9365, n9366, n9367, n9368, n9370, n9371, n9372, n9373, n9374, n9376, n9377, n9378, n9379, n9380, n9381, n9383, n9384, n9385, n9387, n9388, n9390, n9391, n9392, n9394, n9395, n9396, n9397, n9398, n9399, n9401, n9402, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9412, n9413, n9414, n9416, n9417, n9419, n9420, n9423, n9425, n9426, n9427, n9430, n9431, n9433, n9434, n9435, n9437, n9438, n9439, n9441, n9443, n9444, n9445, n9446, n9448, n9450, n9451, n9452, n9454, n9455, n9457, n9458, n9460, n9462, n9463, n9464, n9465, n9466, n9468, n9470, n9471, n9472, n9474, n9475, n9477, n9478, n9479, n9481, n9482, n9484, n9485, n9487, n9488, n9490, n9491, n9493, n9494, n9495, n9497, n9498, n9500, n9501, n9503, n9504, n9505, n9506, n9507, n9509, n9511, n9512, n9514, n9515, n9517, n9518, n9519, n9521, n9522, n9524, n9525, n9527, n9528, n9530, n9532, n9533, n9535, n9536, n9537, n9539, n9540, n9541, n9543, n9544, n9546, n9547, n9549, n9550, n9551, n9553, n9554, n9555, n9557, n9559, n9560, n9562, n9563, n9566, n9567, n9568, n9570, n9571, n9572, n9573, n9575, n9577, n9578, n9579, n9580, n9581, n9582, n9584, n9586, n9587, n9589, n9590, n9592, n9593, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9605, n9606, n9608, n9609, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9632, n9633, n9634, n9636, n9637, n9639, n9640, n9642, n9643, n9644, n9647, n9648, n9650, n9651, n9652, n9653, n9655, n9657, n9659, n9660, n9661, n9663, n9664, n9666, n9667, n9669, n9670, n9671, n9673, n9674, n9675, n9677, n9678, n9680, n9681, n9683, n9684, n9686, n9687, n9688, n9689, n9690, n9691, n9693, n9694, n9696, n9697, n9698, n9699, n9701, n9702, n9703, n9705, n9706, n9707, n9708, n9710, n9711, n9713, n9714, n9716, n9717, n9719, n9720, n9722, n9723, n9725, n9726, n9728, n9729, n9731, n9732, n9733, n9735, n9736, n9737, n9738, n9740, n9741, n9742, n9744, n9745, n9746, n9748, n9749, n9752, n9754, n9756, n9757, n9758, n9760, n9761, n9763, n9764, n9765, n9766, n9767, n9768, n9770, n9771, n9773, n9775, n9777, n9778, n9780, n9782, n9783, n9784, n9786, n9787, n9789, n9790, n9791, n9793, n9795, n9796, n9797, n9799, n9800, n9802, n9803, n9805, n9806, n9807, n9809, n9811, n9812, n9813, n9814, n9816, n9817, n9819, n9820, n9822, n9823, n9824, n9826, n9827, n9828, n9830, n9832, n9833, n9834, n9836, n9837, n9838, n9840, n9841, n9842, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9888, n9890, n9891, n9892, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9903, n9904, n9905, n9906, n9908, n9909, n9910, n9912, n9914, n9915, n9916, n9918, n9920, n9921, n9922, n9924, n9925, n9926, n9927, n9928, n9929, n9931, n9932, n9933, n9935, n9936, n9937, n9939, n9940, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9952, n9954, n9955, n9956, n9957, n9959, n9960, n9962, n9965, n9966, n9967, n9969, n9970, n9972, n9973, n9975, n9976, n9977, n9979, n9980, n9981, n9982, n9984, n9986, n9987, n9990, n9992, n9993, n9995, n9997, n9998, n10001, n10002, n10003, n10004, n10006, n10007, n10009, n10010, n10011, n10012, n10014, n10015, n10016, n10017, n10018, n10020, n10022, n10023, n10025, n10026, n10028, n10029, n10031, n10033, n10034, n10035, n10036, n10037, n10040, n10041, n10043, n10044, n10046, n10047, n10049, n10050, n10052, n10054, n10056, n10058, n10059, n10061, n10062, n10064, n10065, n10066, n10067, n10069, n10071, n10072, n10074, n10075, n10076, n10077, n10078, n10079, n10081, n10082, n10083, n10085, n10087, n10088, n10090, n10091, n10092, n10094, n10095, n10097, n10098, n10099, n10101, n10102, n10104, n10105, n10106, n10107, n10109, n10110, n10112, n10113, n10114, n10115, n10117, n10118, n10119, n10121, n10122, n10123, n10125, n10126, n10127, n10129, n10130, n10132, n10133, n10134, n10136, n10137, n10139, n10140, n10142, n10143, n10144, n10146, n10148, n10150, n10152, n10154, n10156, n10158, n10159, n10160, n10161, n10163, n10164, n10165, n10167, n10168, n10170, n10172, n10173, n10175, n10176, n10177, n10179, n10182, n10183, n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10195, n10197, n10198, n10200, n10201, n10202, n10204, n10205, n10208, n10210, n10211, n10212, n10213, n10214, n10216, n10217, n10219, n10220, n10222, n10223, n10225, n10226, n10227, n10229, n10230, n10231, n10233, n10234, n10236, n10238, n10239, n10241, n10243, n10245, n10246, n10248, n10251, n10252, n10253, n10256, n10257, n10258, n10259, n10260, n10261, n10263, n10265, n10266, n10267, n10268, n10269, n10271, n10272, n10273, n10275, n10276, n10277, n10279, n10280, n10281, n10283, n10284, n10285, n10287, n10288, n10289, n10290, n10292, n10293, n10295, n10296, n10298, n10299, n10302, n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10313, n10314, n10316, n10317, n10319, n10320, n10322, n10324, n10325, n10327, n10328, n10329, n10331, n10333, n10335, n10336, n10337, n10339, n10341, n10342, n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10352, n10353, n10355, n10356, n10357, n10359, n10361, n10362, n10365, n10366, n10368, n10370, n10371, n10373, n10374, n10375, n10376, n10377, n10378, n10380, n10382, n10383, n10385, n10386, n10387, n10389, n10390, n10391, n10393, n10395, n10396, n10398, n10399, n10401, n10402, n10404, n10406, n10407, n10409, n10411, n10412, n10413, n10415, n10416, n10418, n10420, n10422, n10423, n10424, n10425, n10426, n10428, n10429, n10430, n10431, n10433, n10434, n10436, n10437, n10438, n10440, n10441, n10444, n10445, n10446, n10447, n10448, n10451, n10453, n10454, n10456, n10457, n10458, n10460, n10462, n10463, n10465, n10466, n10468, n10469, n10470, n10471, n10472, n10473, n10475, n10477, n10479, n10481, n10482, n10483, n10485, n10487, n10488, n10489, n10490, n10491, n10494, n10496, n10497, n10498, n10499, n10500, n10503, n10505, n10506, n10507, n10509, n10511, n10512, n10513, n10515, n10516, n10518, n10519, n10520, n10521, n10523, n10525, n10526, n10527, n10528, n10530, n10531, n10532, n10534, n10536, n10537, n10538, n10540, n10541, n10543, n10545, n10546, n10547, n10548, n10549, n10551, n10552, n10555, n10556, n10558, n10559, n10561, n10562, n10564, n10565, n10567, n10568, n10569, n10571, n10573, n10575, n10576, n10577, n10579, n10580, n10581, n10584, n10586, n10587, n10589, n10590, n10591, n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10603, n10604, n10605, n10607, n10608, n10610, n10611, n10612, n10614, n10615, n10618, n10621, n10622, n10624, n10625, n10627, n10629, n10631, n10632, n10633, n10635, n10636, n10638, n10639, n10640, n10642, n10644, n10645, n10647, n10648, n10649, n10650, n10652, n10653, n10654, n10656, n10657, n10658, n10659, n10661, n10663, n10664, n10666, n10667, n10668, n10670, n10673, n10674, n10675, n10676, n10677, n10679, n10681, n10682, n10683, n10685, n10686, n10688, n10690, n10691, n10692, n10694, n10696, n10697, n10698, n10699, n10700, n10701, n10703, n10704, n10706, n10708, n10709, n10710, n10712, n10713, n10716, n10718, n10719, n10721, n10722, n10724, n10725, n10728, n10729, n10732, n10734, n10736, n10738, n10740, n10741, n10743, n10745, n10746, n10748, n10749, n10751, n10753, n10754, n10757, n10759, n10761, n10763, n10765, n10766, n10767, n10769, n10770, n10771, n10772, n10774, n10775, n10776, n10778, n10779, n10781, n10782, n10783, n10784, n10785, n10788, n10789, n10791, n10792, n10794, n10795, n10798, n10799, n10800, n10801, n10802, n10803, n10805, n10807, n10810, n10811, n10814, n10815, n10816, n10818, n10819, n10820, n10822, n10823, n10825, n10826, n10827, n10829, n10831, n10832, n10834, n10836, n10838, n10840, n10841, n10842, n10843, n10845, n10847, n10848, n10851, n10854, n10856, n10857, n10859, n10861, n10862, n10863, n10865, n10866, n10868, n10869, n10872, n10873, n10874, n10875, n10877, n10878, n10879, n10882, n10884, n10885, n10886, n10888, n10889, n10890, n10892, n10893, n10894, n10896, n10897, n10898, n10899, n10901, n10902, n10904, n10905, n10908, n10910, n10911;
INVX1    g0000(.A(g35), .Y(n4620));
AND2X1   g0001(.A(g3003), .B(n4620), .Y(g21727));
INVX1    g0002(.A(g37), .Y(g23002));
NOR2X1   g0003(.A(g25), .B(g22), .Y(g23190));
INVX1    g0004(.A(g136), .Y(g23612));
INVX1    g0005(.A(g2834), .Y(g23652));
INVX1    g0006(.A(g2831), .Y(g23759));
ONE      g0007(.Y(g24151));
AND2X1   g0008(.A(g5357), .B(g5297), .Y(g25114));
INVX1    g0009(.A(g1648), .Y(n4629));
NOR2X1   g0010(.A(n4629), .B(g1657), .Y(g25167));
INVX1    g0011(.A(g1668), .Y(n4631));
NOR2X1   g0012(.A(g1636), .B(n4631), .Y(g25259));
ONE      g0013(.Y(g25582));
ONE      g0014(.Y(g25583));
ONE      g0015(.Y(g25584));
ONE      g0016(.Y(g25585));
ONE      g0017(.Y(g25586));
ONE      g0018(.Y(g25587));
ONE      g0019(.Y(g25588));
ONE      g0020(.Y(g25589));
ONE      g0021(.Y(g25590));
INVX1    g0022(.A(g5180), .Y(n4642_1));
INVX1    g0023(.A(g5188), .Y(n4643));
INVX1    g0024(.A(g5176), .Y(n4644));
NOR3X1   g0025(.A(n4644), .B(n4643), .C(n4642_1), .Y(g26801));
OR4X1    g0026(.A(g1830), .B(g2098), .C(g1696), .D(g1964), .Y(n4646));
OR4X1    g0027(.A(g2523), .B(g2255), .C(g2657), .D(g2389), .Y(n4647_1));
NAND3X1  g0028(.A(n4647_1), .B(n4646), .C(g35), .Y(g26875));
NOR4X1   g0029(.A(g1858), .B(g1844), .C(g2112), .D(g1724), .Y(n4649));
NOR4X1   g0030(.A(g2126), .B(g1978), .C(g1992), .D(g1710), .Y(n4650));
AOI21X1  g0031(.A0(n4650), .A1(n4649), .B0(n4620), .Y(n4651));
NOR4X1   g0032(.A(g2283), .B(g2417), .C(g2403), .D(g2671), .Y(n4652_1));
NOR4X1   g0033(.A(g2269), .B(g2551), .C(g2537), .D(g2685), .Y(n4653));
AOI21X1  g0034(.A0(n4653), .A1(n4652_1), .B0(n4620), .Y(n4654));
NAND2X1  g0035(.A(n4654), .B(n4651), .Y(g26876));
NOR4X1   g0036(.A(g1779), .B(g2047), .C(g1798), .D(g1644), .Y(n4656));
NOR4X1   g0037(.A(g1932), .B(g1913), .C(g1664), .D(g2066), .Y(n4657_1));
AOI21X1  g0038(.A0(n4657_1), .A1(n4656), .B0(n4620), .Y(n4658));
NOR4X1   g0039(.A(g2338), .B(g2204), .C(g2625), .D(g2357), .Y(n4659));
NOR4X1   g0040(.A(g2491), .B(g2606), .C(g2223), .D(g2472), .Y(n4660));
AOI21X1  g0041(.A0(n4660), .A1(n4659), .B0(n4620), .Y(n4661));
NAND2X1  g0042(.A(n4661), .B(n4658), .Y(g26877));
INVX1    g0043(.A(g1075), .Y(n4663));
NOR4X1   g0044(.A(g1221), .B(g1216), .C(g1205), .D(g1211), .Y(n4664));
INVX1    g0045(.A(g1171), .Y(n4665));
INVX1    g0046(.A(g979), .Y(n4666));
INVX1    g0047(.A(g1061), .Y(n4667_1));
NOR4X1   g0048(.A(n4666), .B(g1183), .C(n4665), .D(n4667_1), .Y(n4668));
AOI21X1  g0049(.A0(n4668), .A1(n4664), .B0(n4663), .Y(g27831));
OAI21X1  g0050(.A0(g6523), .A1(g6537), .B0(g35), .Y(n4670));
OAI21X1  g0051(.A0(g5845), .A1(g5831), .B0(g35), .Y(n4671));
NAND2X1  g0052(.A(n4671), .B(n4670), .Y(n4672_1));
OAI21X1  g0053(.A0(g6191), .A1(g6177), .B0(g35), .Y(n4673));
INVX1    g0054(.A(n4673), .Y(n4674));
OAI21X1  g0055(.A0(g5485), .A1(g5499), .B0(g35), .Y(n4675));
INVX1    g0056(.A(n4675), .Y(n4676));
OAI21X1  g0057(.A0(g5152), .A1(g5138), .B0(g35), .Y(n4677_1));
OAI21X1  g0058(.A0(g3845), .A1(g3831), .B0(g35), .Y(n4678));
OAI21X1  g0059(.A0(g3129), .A1(g3143), .B0(g35), .Y(n4679));
INVX1    g0060(.A(n4679), .Y(n4680));
OAI21X1  g0061(.A0(g3480), .A1(g3494), .B0(g35), .Y(n4681));
NAND4X1  g0062(.A(n4680), .B(n4678), .C(n4677_1), .D(n4681), .Y(n4682_1));
OR4X1    g0063(.A(n4676), .B(n4674), .C(n4672_1), .D(n4682_1), .Y(n4683));
NOR3X1   g0064(.A(n4676), .B(n4674), .C(n4672_1), .Y(n4684));
INVX1    g0065(.A(n4677_1), .Y(n4685));
NAND2X1  g0066(.A(n4681), .B(n4679), .Y(n4686));
NOR3X1   g0067(.A(n4686), .B(n4678), .C(n4685), .Y(n4687_1));
NAND2X1  g0068(.A(n4678), .B(n4677_1), .Y(n4688));
NOR3X1   g0069(.A(n4681), .B(n4680), .C(n4688), .Y(n4689));
OAI21X1  g0070(.A0(n4689), .A1(n4687_1), .B0(n4684), .Y(n4690));
NAND4X1  g0071(.A(n4679), .B(n4678), .C(n4677_1), .D(n4681), .Y(n4691));
NOR4X1   g0072(.A(n4675), .B(n4674), .C(n4672_1), .D(n4691), .Y(n4692_1));
INVX1    g0073(.A(n4671), .Y(n4693));
NAND4X1  g0074(.A(n4673), .B(n4693), .C(n4670), .D(n4679), .Y(n4694));
NAND2X1  g0075(.A(n4681), .B(n4678), .Y(n4695));
NOR4X1   g0076(.A(n4694), .B(n4685), .C(n4676), .D(n4695), .Y(n4696));
NOR4X1   g0077(.A(n4676), .B(n4674), .C(n4672_1), .D(n4691), .Y(n4697_1));
NAND4X1  g0078(.A(n4679), .B(n4678), .C(n4685), .D(n4681), .Y(n4698));
NOR4X1   g0079(.A(n4676), .B(n4674), .C(n4672_1), .D(n4698), .Y(n4699));
NOR4X1   g0080(.A(n4697_1), .B(n4696), .C(n4692_1), .D(n4699), .Y(n4700));
NOR3X1   g0081(.A(n4685), .B(n4676), .C(n4693), .Y(n4701));
NOR4X1   g0082(.A(n4680), .B(n4674), .C(n4670), .D(n4695), .Y(n4702_1));
INVX1    g0083(.A(n4670), .Y(n4703));
NOR4X1   g0084(.A(n4680), .B(n4673), .C(n4703), .D(n4695), .Y(n4704));
OAI21X1  g0085(.A0(n4704), .A1(n4702_1), .B0(n4701), .Y(n4705));
NAND4X1  g0086(.A(n4700), .B(n4690), .C(n4683), .D(n4705), .Y(g28030));
INVX1    g0087(.A(g1193), .Y(n4707_1));
NOR2X1   g0088(.A(g1008), .B(g969), .Y(n4708));
NOR2X1   g0089(.A(n4708), .B(n4707_1), .Y(n4709));
INVX1    g0090(.A(n4709), .Y(n4710));
INVX1    g0091(.A(g1536), .Y(n4711));
NOR2X1   g0092(.A(g1351), .B(g1312), .Y(n4712_1));
NOR2X1   g0093(.A(n4712_1), .B(n4711), .Y(n4713));
INVX1    g0094(.A(n4713), .Y(n4714));
NAND3X1  g0095(.A(n4714), .B(n4710), .C(g35), .Y(g28041));
INVX1    g0096(.A(g962), .Y(n4716));
INVX1    g0097(.A(g1306), .Y(n4717_1));
NAND3X1  g0098(.A(n4717_1), .B(n4716), .C(g35), .Y(g28042));
INVX1    g0099(.A(g4646), .Y(n4719));
INVX1    g0100(.A(g4776), .Y(n4720));
NOR3X1   g0101(.A(g4793), .B(g4801), .C(n4720), .Y(n4721));
INVX1    g0102(.A(g4698), .Y(n4722_1));
NAND3X1  g0103(.A(g4659), .B(g4669), .C(g4653), .Y(n4723));
NOR4X1   g0104(.A(n4722_1), .B(g4785), .C(g4709), .D(n4723), .Y(n4724));
AOI21X1  g0105(.A0(n4724), .A1(n4721), .B0(n4719), .Y(g28753));
NOR3X1   g0106(.A(g4093), .B(g4087), .C(g4098), .Y(n4726));
NAND3X1  g0107(.A(n4726), .B(g4112), .C(g4076), .Y(n4727_1));
NOR2X1   g0108(.A(g4141), .B(g4082), .Y(n4728));
INVX1    g0109(.A(g4064), .Y(n4729));
INVX1    g0110(.A(g4125), .Y(n4730));
INVX1    g0111(.A(g4057), .Y(n4731_1));
NAND3X1  g0112(.A(n4731_1), .B(n4730), .C(n4729), .Y(n4732));
AOI21X1  g0113(.A0(n4728), .A1(n4727_1), .B0(n4732), .Y(g31521));
NAND2X1  g0114(.A(g2873), .B(g113), .Y(g31656));
NAND2X1  g0115(.A(g2868), .B(g113), .Y(g31665));
AND2X1   g0116(.A(g6163), .B(g35), .Y(n4736_1));
AND2X1   g0117(.A(g5471), .B(g35), .Y(n4737));
AND2X1   g0118(.A(g5817), .B(g35), .Y(n4738));
AND2X1   g0119(.A(g5124), .B(g35), .Y(n4739));
NOR4X1   g0120(.A(n4738), .B(n4737), .C(n4736_1), .D(n4739), .Y(n4740));
OAI21X1  g0121(.A0(g4420), .A1(g4427), .B0(g35), .Y(n4741_1));
OAI21X1  g0122(.A0(g6509), .A1(g3466), .B0(g35), .Y(n4742));
OAI21X1  g0123(.A0(g3115), .A1(g3817), .B0(g35), .Y(n4743));
NAND4X1  g0124(.A(n4742), .B(n4741_1), .C(n4740), .D(n4743), .Y(n4744));
INVX1    g0125(.A(n4744), .Y(n4745));
INVX1    g0126(.A(n4741_1), .Y(n4746_1));
NAND2X1  g0127(.A(n4742), .B(n4737), .Y(n4747));
AND2X1   g0128(.A(g3817), .B(g35), .Y(n4748));
AND2X1   g0129(.A(g3115), .B(g35), .Y(n4749));
OR4X1    g0130(.A(n4748), .B(n4738), .C(n4736_1), .D(n4749), .Y(n4750));
NOR4X1   g0131(.A(n4747), .B(n4746_1), .C(n4739), .D(n4750), .Y(n4751_1));
INVX1    g0132(.A(n4742), .Y(n4752));
INVX1    g0133(.A(n4743), .Y(n4753));
OR2X1    g0134(.A(n4746_1), .B(n4739), .Y(n4754));
OR2X1    g0135(.A(n4754), .B(n4737), .Y(n4755));
INVX1    g0136(.A(g6163), .Y(n4756_1));
NAND3X1  g0137(.A(n4756_1), .B(g5817), .C(g35), .Y(n4757));
NOR4X1   g0138(.A(n4755), .B(n4753), .C(n4752), .D(n4757), .Y(n4758));
OR4X1    g0139(.A(n4738), .B(n4737), .C(n4736_1), .D(n4748), .Y(n4759));
INVX1    g0140(.A(n4749), .Y(n4760));
NAND4X1  g0141(.A(n4742), .B(n4741_1), .C(n4739), .D(n4760), .Y(n4761_1));
NOR2X1   g0142(.A(n4761_1), .B(n4759), .Y(n4762));
NOR4X1   g0143(.A(n4758), .B(n4751_1), .C(n4745), .D(n4762), .Y(n4763));
NOR4X1   g0144(.A(n4748), .B(n4752), .C(n4746_1), .D(n4760), .Y(n4764));
AND2X1   g0145(.A(g6509), .B(g35), .Y(n4765));
NAND2X1  g0146(.A(g3466), .B(g35), .Y(n4766_1));
NOR4X1   g0147(.A(n4766_1), .B(n4765), .C(n4746_1), .D(n4753), .Y(n4767));
OAI21X1  g0148(.A0(n4767), .A1(n4764), .B0(n4740), .Y(n4768));
NOR3X1   g0149(.A(n4753), .B(n4752), .C(n4741_1), .Y(n4769));
INVX1    g0150(.A(n4748), .Y(n4770_1));
NOR4X1   g0151(.A(n4770_1), .B(n4752), .C(n4746_1), .D(n4749), .Y(n4771));
OAI21X1  g0152(.A0(n4771), .A1(n4769), .B0(n4740), .Y(n4772));
NOR4X1   g0153(.A(n4739), .B(n4738), .C(n4737), .D(n4746_1), .Y(n4773));
NOR4X1   g0154(.A(n4752), .B(n4756_1), .C(n4620), .D(n4753), .Y(n4774));
NAND2X1  g0155(.A(n4766_1), .B(n4765), .Y(n4775_1));
NOR4X1   g0156(.A(n4749), .B(n4748), .C(n4736_1), .D(n4775_1), .Y(n4776));
OAI21X1  g0157(.A0(n4776), .A1(n4774), .B0(n4773), .Y(n4777));
NAND4X1  g0158(.A(n4772), .B(n4768), .C(n4763), .D(n4777), .Y(g31793));
NAND2X1  g0159(.A(g2965), .B(g2960), .Y(n4779));
AOI22X1  g0160(.A0(g2950), .A1(g2955), .B0(g2941), .B1(g2936), .Y(n4780_1));
NAND2X1  g0161(.A(n4780_1), .B(n4779), .Y(n4781));
INVX1    g0162(.A(g2975), .Y(n4782));
INVX1    g0163(.A(g2970), .Y(n4783));
NAND2X1  g0164(.A(g2902), .B(g2907), .Y(n4784_1));
OAI21X1  g0165(.A0(n4783), .A1(n4782), .B0(n4784_1), .Y(n4785));
INVX1    g0166(.A(g2927), .Y(n4786));
INVX1    g0167(.A(g2917), .Y(n4787));
INVX1    g0168(.A(g2922), .Y(n4788_1));
INVX1    g0169(.A(g2912), .Y(n4789));
OAI22X1  g0170(.A0(n4788_1), .A1(n4786), .B0(n4787), .B1(n4789), .Y(n4790));
NOR3X1   g0171(.A(n4790), .B(n4785), .C(n4781), .Y(g32185));
ONE      g0172(.Y(g32429));
ONE      g0173(.Y(g32454));
OR2X1    g0174(.A(g2803), .B(g2724), .Y(n4794));
INVX1    g0175(.A(g2807), .Y(n4795));
AOI21X1  g0176(.A0(g2724), .A1(n4795), .B0(g2729), .Y(n4796));
OR2X1    g0177(.A(g2724), .B(g2815), .Y(n4797));
INVX1    g0178(.A(g2819), .Y(n4798_1));
INVX1    g0179(.A(g2729), .Y(n4799));
AOI21X1  g0180(.A0(g2724), .A1(n4798_1), .B0(n4799), .Y(n4800));
AOI22X1  g0181(.A0(n4797), .A1(n4800), .B0(n4796), .B1(n4794), .Y(g33079));
OR2X1    g0182(.A(g2724), .B(g2771), .Y(n4802));
INVX1    g0183(.A(g2775), .Y(n4803_1));
AOI21X1  g0184(.A0(n4803_1), .A1(g2724), .B0(g2729), .Y(n4804));
OR2X1    g0185(.A(g2724), .B(g2783), .Y(n4805));
INVX1    g0186(.A(g2787), .Y(n4806));
AOI21X1  g0187(.A0(n4806), .A1(g2724), .B0(n4799), .Y(n4807));
AOI22X1  g0188(.A0(n4805), .A1(n4807), .B0(n4804), .B1(n4802), .Y(g33435));
AOI21X1  g0189(.A0(g37), .A1(g99), .B0(g134), .Y(n4809));
NAND2X1  g0190(.A(g4815), .B(g4812), .Y(n4810));
NOR2X1   g0191(.A(n4810), .B(n4809), .Y(n4811));
NOR2X1   g0192(.A(g4785), .B(g4709), .Y(n4812_1));
AND2X1   g0193(.A(n4812_1), .B(g4698), .Y(n4813));
INVX1    g0194(.A(g4754), .Y(n4814));
INVX1    g0195(.A(g4709), .Y(n4815));
NOR3X1   g0196(.A(g4785), .B(n4815), .C(n4814), .Y(n4816));
INVX1    g0197(.A(g4743), .Y(n4817_1));
INVX1    g0198(.A(g4785), .Y(n4818));
NOR3X1   g0199(.A(n4818), .B(g4709), .C(n4817_1), .Y(n4819));
AND2X1   g0200(.A(g4785), .B(g4709), .Y(n4820));
AND2X1   g0201(.A(n4820), .B(g4765), .Y(n4821));
NOR4X1   g0202(.A(n4819), .B(n4816), .C(n4813), .D(n4821), .Y(n4822_1));
NAND2X1  g0203(.A(n4822_1), .B(n4811), .Y(g33636));
INVX1    g0204(.A(g113), .Y(n4824));
XOR2X1   g0205(.A(g4104), .B(g73), .Y(n4825));
XOR2X1   g0206(.A(g4108), .B(g72), .Y(n4826));
NOR4X1   g0207(.A(n4825), .B(n4809), .C(n4824), .D(n4826), .Y(n4827_1));
INVX1    g0208(.A(n4827_1), .Y(n4828));
INVX1    g0209(.A(g4098), .Y(n4829));
INVX1    g0210(.A(g4093), .Y(n4830));
OR4X1    g0211(.A(n4825), .B(n4830), .C(n4829), .D(n4826), .Y(n4831));
NOR2X1   g0212(.A(n4831), .B(g4087), .Y(n4832_1));
INVX1    g0213(.A(g3530), .Y(n4833));
INVX1    g0214(.A(g3518), .Y(n4834));
INVX1    g0215(.A(g3522), .Y(n4835));
NOR3X1   g0216(.A(n4835), .B(n4834), .C(n4833), .Y(n4836_1));
OR4X1    g0217(.A(n4825), .B(g4093), .C(g4098), .D(n4826), .Y(n4837));
NOR2X1   g0218(.A(n4837), .B(g4087), .Y(n4838));
AOI22X1  g0219(.A0(n4836_1), .A1(n4832_1), .B0(g26801), .B1(n4838), .Y(n4839));
INVX1    g0220(.A(g4087), .Y(n4840));
OR4X1    g0221(.A(n4825), .B(g4093), .C(n4829), .D(n4826), .Y(n4841_1));
NOR2X1   g0222(.A(n4841_1), .B(n4840), .Y(n4842));
INVX1    g0223(.A(g3167), .Y(n4843));
INVX1    g0224(.A(g3179), .Y(n4844));
INVX1    g0225(.A(g3171), .Y(n4845));
NOR3X1   g0226(.A(n4845), .B(n4844), .C(n4843), .Y(n4846_1));
NOR2X1   g0227(.A(n4831), .B(n4840), .Y(n4847));
INVX1    g0228(.A(g3873), .Y(n4848));
INVX1    g0229(.A(g3869), .Y(n4849));
INVX1    g0230(.A(g3881), .Y(n4850));
NOR3X1   g0231(.A(n4850), .B(n4849), .C(n4848), .Y(n4851_1));
AOI22X1  g0232(.A0(n4847), .A1(n4851_1), .B0(n4846_1), .B1(n4842), .Y(n4852));
NOR2X1   g0233(.A(n4841_1), .B(g4087), .Y(n4853));
INVX1    g0234(.A(g6573), .Y(n4854));
INVX1    g0235(.A(g6565), .Y(n4855));
INVX1    g0236(.A(g6561), .Y(n4856_1));
NOR3X1   g0237(.A(n4856_1), .B(n4855), .C(n4854), .Y(n4857));
OR4X1    g0238(.A(n4825), .B(n4830), .C(g4098), .D(n4826), .Y(n4858));
NOR2X1   g0239(.A(n4858), .B(g4087), .Y(n4859));
INVX1    g0240(.A(g5873), .Y(n4860));
INVX1    g0241(.A(g5869), .Y(n4861_1));
INVX1    g0242(.A(g5881), .Y(n4862));
NOR3X1   g0243(.A(n4862), .B(n4861_1), .C(n4860), .Y(n4863));
AOI22X1  g0244(.A0(n4859), .A1(n4863), .B0(n4857), .B1(n4853), .Y(n4864));
NOR2X1   g0245(.A(n4837), .B(n4840), .Y(n4865));
INVX1    g0246(.A(g5523), .Y(n4866_1));
INVX1    g0247(.A(g5535), .Y(n4867));
INVX1    g0248(.A(g5527), .Y(n4868));
NOR3X1   g0249(.A(n4868), .B(n4867), .C(n4866_1), .Y(n4869));
NOR2X1   g0250(.A(n4858), .B(n4840), .Y(n4870));
INVX1    g0251(.A(g6219), .Y(n4871_1));
INVX1    g0252(.A(g6215), .Y(n4872));
INVX1    g0253(.A(g6227), .Y(n4873));
NOR3X1   g0254(.A(n4873), .B(n4872), .C(n4871_1), .Y(n4874));
AOI22X1  g0255(.A0(n4870), .A1(n4874), .B0(n4869), .B1(n4865), .Y(n4875));
NAND4X1  g0256(.A(n4864), .B(n4852), .C(n4839), .D(n4875), .Y(n4876_1));
NOR2X1   g0257(.A(n4876_1), .B(n4828), .Y(n4877));
INVX1    g0258(.A(n4877), .Y(g33659));
INVX1    g0259(.A(g4507), .Y(n4879));
NOR3X1   g0260(.A(n4809), .B(n4879), .C(g66), .Y(n4880));
INVX1    g0261(.A(n4880), .Y(g33874));
INVX1    g0262(.A(g890), .Y(n4882));
INVX1    g0263(.A(g479), .Y(n4883));
XOR2X1   g0264(.A(g482), .B(g72), .Y(n4884));
XOR2X1   g0265(.A(g490), .B(g73), .Y(n4885));
NOR4X1   g0266(.A(n4884), .B(g528), .C(n4883), .D(n4885), .Y(n4886_1));
NOR2X1   g0267(.A(n4886_1), .B(n4882), .Y(g33894));
NAND2X1  g0268(.A(g5005), .B(g5002), .Y(n4888));
NOR2X1   g0269(.A(n4888), .B(n4809), .Y(n4889));
NOR2X1   g0270(.A(g4975), .B(g4899), .Y(n4890));
AND2X1   g0271(.A(n4890), .B(g4888), .Y(n4891_1));
INVX1    g0272(.A(g4944), .Y(n4892));
INVX1    g0273(.A(g4899), .Y(n4893));
NOR3X1   g0274(.A(g4975), .B(n4893), .C(n4892), .Y(n4894));
INVX1    g0275(.A(g4933), .Y(n4895));
INVX1    g0276(.A(g4975), .Y(n4896_1));
NOR3X1   g0277(.A(n4896_1), .B(g4899), .C(n4895), .Y(n4897));
AND2X1   g0278(.A(g4975), .B(g4899), .Y(n4898));
AND2X1   g0279(.A(n4898), .B(g4955), .Y(n4899));
NOR4X1   g0280(.A(n4897), .B(n4894), .C(n4891_1), .D(n4899), .Y(n4900));
NAND2X1  g0281(.A(n4900), .B(n4889), .Y(g33935));
ONE      g0282(.Y(g33945));
ONE      g0283(.Y(g33946));
ONE      g0284(.Y(g33947));
ONE      g0285(.Y(g33948));
ONE      g0286(.Y(g33949));
ONE      g0287(.Y(g33950));
NOR2X1   g0288(.A(n4809), .B(n4824), .Y(n4908));
INVX1    g0289(.A(g2741), .Y(n4909));
INVX1    g0290(.A(g2756), .Y(n4910_1));
XOR2X1   g0291(.A(g2763), .B(g73), .Y(n4911));
XOR2X1   g0292(.A(g2759), .B(g72), .Y(n4912));
NOR4X1   g0293(.A(n4911), .B(g2748), .C(n4910_1), .D(n4912), .Y(n4913));
NAND2X1  g0294(.A(n4913), .B(n4909), .Y(n4914));
INVX1    g0295(.A(g2748), .Y(n4915_1));
NOR4X1   g0296(.A(n4911), .B(n4915_1), .C(n4910_1), .D(n4912), .Y(n4916));
NAND2X1  g0297(.A(n4916), .B(n4909), .Y(n4917));
NAND2X1  g0298(.A(n4913), .B(g2741), .Y(n4918));
NAND2X1  g0299(.A(n4916), .B(g2741), .Y(n4919));
NAND4X1  g0300(.A(n4918), .B(n4917), .C(n4914), .D(n4919), .Y(n4920_1));
NOR4X1   g0301(.A(n4911), .B(g2748), .C(g2756), .D(n4912), .Y(n4921));
NAND2X1  g0302(.A(n4921), .B(n4909), .Y(n4922));
NOR4X1   g0303(.A(n4911), .B(n4915_1), .C(g2756), .D(n4912), .Y(n4923));
NAND2X1  g0304(.A(n4923), .B(n4909), .Y(n4924));
NAND2X1  g0305(.A(n4921), .B(g2741), .Y(n4925_1));
NAND2X1  g0306(.A(n4923), .B(g2741), .Y(n4926));
NAND4X1  g0307(.A(n4925_1), .B(n4924), .C(n4922), .D(n4926), .Y(n4927));
OAI21X1  g0308(.A0(n4927), .A1(n4920_1), .B0(n4908), .Y(n4928));
INVX1    g0309(.A(g2485), .Y(n4929));
NAND4X1  g0310(.A(n4909), .B(g2476), .C(n4929), .D(n4916), .Y(n4930_1));
NAND3X1  g0311(.A(n4921), .B(g25167), .C(n4909), .Y(n4931));
INVX1    g0312(.A(g2351), .Y(n4932));
NAND4X1  g0313(.A(g2741), .B(n4932), .C(g2342), .D(n4913), .Y(n4933));
INVX1    g0314(.A(g2619), .Y(n4934_1));
NAND4X1  g0315(.A(g2741), .B(n4934_1), .C(g2610), .D(n4916), .Y(n4935));
NAND4X1  g0316(.A(n4933), .B(n4931), .C(n4930_1), .D(n4935), .Y(n4936));
INVX1    g0317(.A(g2217), .Y(n4937));
NAND4X1  g0318(.A(n4937), .B(n4909), .C(g2208), .D(n4913), .Y(n4938));
INVX1    g0319(.A(g1926), .Y(n4939_1));
NAND4X1  g0320(.A(n4909), .B(g1917), .C(n4939_1), .D(n4923), .Y(n4940));
INVX1    g0321(.A(g1792), .Y(n4941));
NAND4X1  g0322(.A(n4941), .B(g2741), .C(g1783), .D(n4921), .Y(n4942));
INVX1    g0323(.A(g2060), .Y(n4943));
NAND4X1  g0324(.A(n4943), .B(g2051), .C(g2741), .D(n4923), .Y(n4944_1));
NAND4X1  g0325(.A(n4942), .B(n4940), .C(n4938), .D(n4944_1), .Y(n4945));
OR2X1    g0326(.A(n4945), .B(n4936), .Y(n4946));
NOR2X1   g0327(.A(n4946), .B(n4928), .Y(n4947));
INVX1    g0328(.A(n4947), .Y(g34201));
INVX1    g0329(.A(g4311), .Y(n4949_1));
INVX1    g0330(.A(g72), .Y(n4950));
XOR2X1   g0331(.A(g4322), .B(n4950), .Y(n4951));
INVX1    g0332(.A(n4951), .Y(n4952));
INVX1    g0333(.A(g73), .Y(n4953));
XOR2X1   g0334(.A(g4332), .B(n4953), .Y(n4954_1));
INVX1    g0335(.A(n4954_1), .Y(n4955));
NOR3X1   g0336(.A(n4955), .B(n4952), .C(n4949_1), .Y(n4956));
NOR3X1   g0337(.A(n4955), .B(n4952), .C(g4311), .Y(n4957));
OAI21X1  g0338(.A0(n4957), .A1(n4956), .B0(n4908), .Y(n4958));
INVX1    g0339(.A(g4878), .Y(n4959_1));
NAND3X1  g0340(.A(g4843), .B(g4859), .C(g4849), .Y(n4960));
NOR2X1   g0341(.A(n4960), .B(n4959_1), .Y(n4961));
INVX1    g0342(.A(g4983), .Y(n4962));
INVX1    g0343(.A(g4966), .Y(n4963));
NOR3X1   g0344(.A(n4963), .B(g4991), .C(n4962), .Y(n4964_1));
NAND3X1  g0345(.A(n4964_1), .B(n4961), .C(n4898), .Y(n4965));
NOR4X1   g0346(.A(n4955), .B(n4952), .C(n4949_1), .D(n4965), .Y(n4966));
INVX1    g0347(.A(g4688), .Y(n4967));
NOR2X1   g0348(.A(n4723), .B(n4967), .Y(n4968));
INVX1    g0349(.A(g4793), .Y(n4969_1));
NOR3X1   g0350(.A(n4969_1), .B(g4801), .C(n4720), .Y(n4970));
NAND3X1  g0351(.A(n4970), .B(n4968), .C(n4820), .Y(n4971));
NOR4X1   g0352(.A(n4955), .B(n4952), .C(g4311), .D(n4971), .Y(n4972));
NOR3X1   g0353(.A(n4972), .B(n4966), .C(n4958), .Y(n4973));
INVX1    g0354(.A(n4973), .Y(g34221));
ONE      g0355(.Y(g34232));
INVX1    g0356(.A(g54), .Y(n4976));
OR2X1    g0357(.A(g34), .B(g53), .Y(n4977));
NOR4X1   g0358(.A(n4976), .B(g57), .C(g56), .D(n4977), .Y(n4383));
INVX1    g0359(.A(g16), .Y(n4979_1));
INVX1    g0360(.A(g19), .Y(n4980));
NOR3X1   g0361(.A(n4980), .B(g9), .C(n4979_1), .Y(n4981));
INVX1    g0362(.A(g28), .Y(n4982));
NOR4X1   g0363(.A(g8), .B(g6), .C(g31), .D(g7), .Y(n4983));
AND2X1   g0364(.A(n4983), .B(n4982), .Y(n4984_1));
NAND3X1  g0365(.A(n4984_1), .B(n4981), .C(n4383), .Y(n4985));
INVX1    g0366(.A(n4985), .Y(n4986));
OR4X1    g0367(.A(n4976), .B(g57), .C(g56), .D(n4977), .Y(n4987));
NAND3X1  g0368(.A(g19), .B(g9), .C(n4979_1), .Y(n4988_1));
NOR3X1   g0369(.A(g7), .B(g8), .C(g6), .Y(n4989));
NAND2X1  g0370(.A(n4989), .B(g31), .Y(n4990));
OR4X1    g0371(.A(n4988_1), .B(n4987), .C(g28), .D(n4990), .Y(n4991));
INVX1    g0372(.A(g6), .Y(n4992_1));
INVX1    g0373(.A(g8), .Y(n4993));
INVX1    g0374(.A(g7), .Y(n4994));
OR4X1    g0375(.A(n4993), .B(n4992_1), .C(g31), .D(n4994), .Y(n4995));
NOR2X1   g0376(.A(g19), .B(g16), .Y(n4996));
NAND2X1  g0377(.A(n4996), .B(g9), .Y(n4997_1));
NOR3X1   g0378(.A(n4997_1), .B(n4995), .C(g28), .Y(n4998));
NOR3X1   g0379(.A(n4995), .B(n4988_1), .C(n4982), .Y(n4999));
NOR3X1   g0380(.A(n4997_1), .B(n4995), .C(n4982), .Y(n5000));
NAND3X1  g0381(.A(n4980), .B(g9), .C(g16), .Y(n5001));
NOR3X1   g0382(.A(n5001), .B(n4995), .C(g28), .Y(n5002_1));
OR4X1    g0383(.A(n5000), .B(n4999), .C(n4998), .D(n5002_1), .Y(n5003));
NAND2X1  g0384(.A(n4983), .B(g28), .Y(n5004));
INVX1    g0385(.A(g9), .Y(n5005));
NAND3X1  g0386(.A(n4980), .B(n5005), .C(g16), .Y(n5006));
NOR2X1   g0387(.A(n5006), .B(n5004), .Y(n5007_1));
OR4X1    g0388(.A(g8), .B(g6), .C(g31), .D(g7), .Y(n5008));
OR2X1    g0389(.A(g19), .B(g16), .Y(n5009));
NOR4X1   g0390(.A(n5008), .B(g28), .C(n5005), .D(n5009), .Y(n5010));
NAND3X1  g0391(.A(n4989), .B(g28), .C(g31), .Y(n5011));
NOR2X1   g0392(.A(n5011), .B(n5006), .Y(n5012_1));
NOR4X1   g0393(.A(n5008), .B(n4982), .C(n5005), .D(n5009), .Y(n5013));
OR4X1    g0394(.A(n5012_1), .B(n5010), .C(n5007_1), .D(n5013), .Y(n5014));
OAI21X1  g0395(.A0(n5014), .A1(n5003), .B0(n4383), .Y(n5015));
NOR3X1   g0396(.A(g19), .B(g9), .C(n4979_1), .Y(n5016));
NAND3X1  g0397(.A(n5016), .B(n4984_1), .C(n4383), .Y(n5017_1));
NAND3X1  g0398(.A(n5017_1), .B(n5015), .C(n4991), .Y(n5018));
NAND2X1  g0399(.A(n4983), .B(n4982), .Y(n5019));
NOR3X1   g0400(.A(n4988_1), .B(n5019), .C(n4987), .Y(n5020));
NAND3X1  g0401(.A(n4989), .B(n4982), .C(g31), .Y(n5021));
NOR3X1   g0402(.A(g19), .B(g9), .C(g16), .Y(n5022_1));
NAND4X1  g0403(.A(n4989), .B(g28), .C(g31), .D(n5022_1), .Y(n5023));
NAND3X1  g0404(.A(g19), .B(n5005), .C(n4979_1), .Y(n5024));
OAI21X1  g0405(.A0(n5024), .A1(n5021), .B0(n5023), .Y(n5025));
NOR4X1   g0406(.A(n5008), .B(g28), .C(g9), .D(n5009), .Y(n5026));
NAND3X1  g0407(.A(n5022_1), .B(n4983), .C(g28), .Y(n5027_1));
OAI21X1  g0408(.A0(n5024), .A1(n5019), .B0(n5027_1), .Y(n5028));
NOR3X1   g0409(.A(n5028), .B(n5026), .C(n5025), .Y(n5029));
OR2X1    g0410(.A(n5029), .B(n4987), .Y(n5030));
NAND3X1  g0411(.A(g19), .B(n5005), .C(g16), .Y(n5031));
NOR3X1   g0412(.A(n5004), .B(n5031), .C(n4987), .Y(n5032_1));
NOR3X1   g0413(.A(n5024), .B(n5004), .C(n4987), .Y(n5033));
NOR2X1   g0414(.A(n4383), .B(g53), .Y(n5034));
NOR2X1   g0415(.A(n5034), .B(n5033), .Y(n5035));
NAND3X1  g0416(.A(n5035), .B(n5032_1), .C(n5030), .Y(n5036));
OR4X1    g0417(.A(n5020), .B(n5018), .C(n4986), .D(n5036), .Y(n5037_1));
NAND3X1  g0418(.A(n5017_1), .B(n5015), .C(n4985), .Y(n5038));
NOR2X1   g0419(.A(n5038), .B(n5032_1), .Y(n5039));
NOR2X1   g0420(.A(n5029), .B(n4987), .Y(n5040));
INVX1    g0421(.A(n5035), .Y(n5041));
NOR4X1   g0422(.A(n5040), .B(n5020), .C(n4991), .D(n5041), .Y(n5042_1));
NAND3X1  g0423(.A(n5035), .B(n5030), .C(n5020), .Y(n5043));
NOR4X1   g0424(.A(n5032_1), .B(n5018), .C(n4986), .D(n5043), .Y(n5044));
AOI21X1  g0425(.A0(n5042_1), .A1(n5039), .B0(n5044), .Y(n5045));
NOR3X1   g0426(.A(n5021), .B(n4988_1), .C(n4987), .Y(n5046));
NOR3X1   g0427(.A(n5006), .B(n5019), .C(n4987), .Y(n5047_1));
NOR3X1   g0428(.A(n4980), .B(n5005), .C(g16), .Y(n5048));
NAND3X1  g0429(.A(n5048), .B(n4984_1), .C(n4383), .Y(n5049));
AND2X1   g0430(.A(n4983), .B(g28), .Y(n5050));
NAND3X1  g0431(.A(n5050), .B(n4981), .C(n4383), .Y(n5051_1));
NAND2X1  g0432(.A(n5051_1), .B(n5049), .Y(n5052));
OR4X1    g0433(.A(n5047_1), .B(n5046), .C(n4986), .D(n5052), .Y(n5053));
NOR4X1   g0434(.A(n5041), .B(n5040), .C(n5015), .D(n5053), .Y(n5054));
NOR4X1   g0435(.A(n5033), .B(n5040), .C(n5047_1), .D(n5034), .Y(n5055));
NAND4X1  g0436(.A(n5015), .B(n4991), .C(n4985), .D(n5051_1), .Y(n5056_1));
NOR2X1   g0437(.A(n5056_1), .B(n5020), .Y(n5057));
AND2X1   g0438(.A(n5057), .B(n5055), .Y(n5058));
NAND3X1  g0439(.A(n5035), .B(n5030), .C(n4986), .Y(n5059));
NOR3X1   g0440(.A(n5059), .B(n5052), .C(n5018), .Y(n5060));
NOR3X1   g0441(.A(n5060), .B(n5058), .C(n5054), .Y(n5061_1));
OR2X1    g0442(.A(n4383), .B(g53), .Y(n5062));
NOR3X1   g0443(.A(n5041), .B(n5040), .C(n5017_1), .Y(n5066_1));
OR4X1    g0444(.A(n5008), .B(n4987), .C(n4982), .D(n5024), .Y(n5067));
NOR4X1   g0445(.A(n5067), .B(n5040), .C(n5047_1), .D(n5034), .Y(n5068));
NAND4X1  g0446(.A(n5061_1), .B(n5045), .C(n5037_1), .D(n5055), .Y(g34233));
OR2X1    g0447(.A(n5014), .B(n5003), .Y(n5072));
AND2X1   g0448(.A(n5072), .B(n4383), .Y(n5073));
NOR4X1   g0449(.A(n5073), .B(n5046), .C(n4986), .D(n5052), .Y(n5074));
NAND2X1  g0450(.A(n5017_1), .B(n5015), .Y(n5076_1));
NOR4X1   g0451(.A(n5052), .B(n5076_1), .C(n5046), .D(n5059), .Y(n5077));
NOR4X1   g0452(.A(n5036), .B(n5020), .C(n5046), .D(n5038), .Y(n5078));
NOR4X1   g0453(.A(n5077), .B(n5058), .C(n5054), .D(n5078), .Y(n5079));
OAI21X1  g0454(.A0(n5068), .A1(n5066_1), .B0(n5074), .Y(n5081_1));
NOR4X1   g0455(.A(n5040), .B(n5049), .C(n5046), .D(n5041), .Y(n5082));
OAI21X1  g0456(.A0(n5082), .A1(n5042_1), .B0(n5039), .Y(n5083));
NAND4X1  g0457(.A(n5081_1), .B(n5122), .C(n5079), .D(n5083), .Y(g34236));
NOR4X1   g0458(.A(n5000), .B(n4999), .C(n4998), .D(n5002_1), .Y(n5085));
NOR3X1   g0459(.A(n5013), .B(n5012_1), .C(n5007_1), .Y(n5086_1));
AOI21X1  g0460(.A0(n5086_1), .A1(n5085), .B0(n4987), .Y(n5087));
NAND2X1  g0461(.A(n5010), .B(n4383), .Y(n5088));
NAND3X1  g0462(.A(n5088), .B(n5049), .C(n4991), .Y(n5089));
NAND3X1  g0463(.A(n5050), .B(n5048), .C(n4383), .Y(n5090));
INVX1    g0464(.A(n5090), .Y(n5091_1));
NOR3X1   g0465(.A(n5091_1), .B(n5089), .C(n5087), .Y(n5092));
AND2X1   g0466(.A(n5092), .B(n5055), .Y(n5093));
NAND4X1  g0467(.A(n5029), .B(n5010), .C(n4383), .D(n5035), .Y(n5094));
NAND3X1  g0468(.A(n5049), .B(n5017_1), .C(n4991), .Y(n5095));
NOR4X1   g0469(.A(n5094), .B(n5091_1), .C(n5087), .D(n5095), .Y(n5096_1));
NAND3X1  g0470(.A(n5087), .B(n5035), .C(n5030), .Y(n5097));
NAND2X1  g0471(.A(n5090), .B(n5088), .Y(n5098));
NOR3X1   g0472(.A(n5098), .B(n5097), .C(n5095), .Y(n5099));
NOR3X1   g0473(.A(n5099), .B(n5096_1), .C(n5093), .Y(n5100));
OR4X1    g0474(.A(n5087), .B(n5047_1), .C(n5046), .D(n5098), .Y(n5102));
NOR2X1   g0475(.A(n5102), .B(n5043), .Y(n5103));
OR4X1    g0476(.A(n5087), .B(n5020), .C(n5047_1), .D(n5098), .Y(n5104));
NOR4X1   g0477(.A(n5041), .B(n5040), .C(n4991), .D(n5104), .Y(n5105));
NOR3X1   g0478(.A(n5105), .B(n5103), .C(n5040), .Y(n5106_1));
INVX1    g0479(.A(n5088), .Y(n5107));
AOI21X1  g0480(.A0(n5092), .A1(n5066_1), .B0(n5091_1), .Y(n5110));
NAND4X1  g0481(.A(n5110), .B(n5106_1), .C(n5100), .D(n5035), .Y(g34237));
NAND3X1  g0482(.A(n5090), .B(n5088), .C(n4985), .Y(n5113));
NOR3X1   g0483(.A(n5113), .B(n5087), .C(n5032_1), .Y(n5114));
AND2X1   g0484(.A(n5114), .B(n5055), .Y(n5115_1));
OR2X1    g0485(.A(n5087), .B(n5047_1), .Y(n5116));
NAND2X1  g0486(.A(n5051_1), .B(n4985), .Y(n5117));
NOR4X1   g0487(.A(n5116), .B(n5094), .C(n5091_1), .D(n5117), .Y(n5118));
NOR4X1   g0488(.A(n5098), .B(n5097), .C(n5047_1), .D(n5117), .Y(n5120_1));
NOR4X1   g0489(.A(n5091_1), .B(n5118), .C(n5115_1), .D(n5120_1), .Y(n5121));
OAI21X1  g0490(.A0(n5040), .A1(n5034), .B0(n5114), .Y(n5122));
OAI21X1  g0491(.A0(n5068), .A1(n5066_1), .B0(n5114), .Y(n5123));
NOR4X1   g0492(.A(n5107), .B(n5087), .C(n5047_1), .D(n5091_1), .Y(n5124));
NOR4X1   g0493(.A(n5032_1), .B(n5040), .C(n4985), .D(n5041), .Y(n5125_1));
NOR4X1   g0494(.A(n5051_1), .B(n5040), .C(n4986), .D(n5041), .Y(n5126));
OAI21X1  g0495(.A0(n5126), .A1(n5125_1), .B0(n5124), .Y(n5127));
NAND4X1  g0496(.A(n5123), .B(n5122), .C(n5121), .D(n5127), .Y(g34239));
INVX1    g0497(.A(g518), .Y(n5129));
INVX1    g0498(.A(g482), .Y(n5130_1));
AOI22X1  g0499(.A0(g490), .A1(n4953), .B0(g72), .B1(n5130_1), .Y(n5131));
INVX1    g0500(.A(g490), .Y(n5132));
AOI22X1  g0501(.A0(n5132), .A1(g73), .B0(n4950), .B1(g482), .Y(n5133));
NAND4X1  g0502(.A(n5131), .B(n5129), .C(g528), .D(n5133), .Y(n5134));
NOR2X1   g0503(.A(n5134), .B(g504), .Y(n5135_1));
INVX1    g0504(.A(g504), .Y(n5136));
NAND4X1  g0505(.A(n5131), .B(g518), .C(g528), .D(n5133), .Y(n5137));
NOR2X1   g0506(.A(n5137), .B(n5136), .Y(n5138));
NOR2X1   g0507(.A(n5134), .B(n5136), .Y(n5139));
NOR2X1   g0508(.A(n5137), .B(g504), .Y(n5140_1));
OR4X1    g0509(.A(n5139), .B(n5138), .C(n5135_1), .D(n5140_1), .Y(n5141));
INVX1    g0510(.A(g528), .Y(n5142));
NAND4X1  g0511(.A(n5131), .B(n5129), .C(n5142), .D(n5133), .Y(n5143));
NOR2X1   g0512(.A(n5143), .B(g504), .Y(n5144));
NAND4X1  g0513(.A(n5131), .B(g518), .C(n5142), .D(n5133), .Y(n5145_1));
NOR2X1   g0514(.A(n5145_1), .B(n5136), .Y(n5146));
NOR2X1   g0515(.A(n5143), .B(n5136), .Y(n5147));
NOR2X1   g0516(.A(n5145_1), .B(g504), .Y(n5148));
OR4X1    g0517(.A(n5147), .B(n5146), .C(n5144), .D(n5148), .Y(n5149_1));
OAI21X1  g0518(.A0(n5149_1), .A1(n5141), .B0(n4908), .Y(n5150));
INVX1    g0519(.A(g2495), .Y(n5151));
NOR2X1   g0520(.A(n5151), .B(g2465), .Y(n5152));
AOI22X1  g0521(.A0(n5144), .A1(g25259), .B0(n5138), .B1(n5152), .Y(n5153_1));
INVX1    g0522(.A(g2361), .Y(n5154));
NOR2X1   g0523(.A(n5154), .B(g2331), .Y(n5155));
INVX1    g0524(.A(g2629), .Y(n5156));
NOR2X1   g0525(.A(n5156), .B(g2599), .Y(n5157));
AOI22X1  g0526(.A0(n5155), .A1(n5139), .B0(n5140_1), .B1(n5157), .Y(n5158_1));
INVX1    g0527(.A(g2227), .Y(n5159));
NOR2X1   g0528(.A(g2197), .B(n5159), .Y(n5160));
INVX1    g0529(.A(g1936), .Y(n5161));
NOR2X1   g0530(.A(g1906), .B(n5161), .Y(n5162_1));
AOI22X1  g0531(.A0(n5160), .A1(n5135_1), .B0(n5146), .B1(n5162_1), .Y(n5163));
INVX1    g0532(.A(g1802), .Y(n5164));
NOR2X1   g0533(.A(g1772), .B(n5164), .Y(n5165));
INVX1    g0534(.A(g2070), .Y(n5166_1));
NOR2X1   g0535(.A(n5166_1), .B(g2040), .Y(n5167));
AOI22X1  g0536(.A0(n5165), .A1(n5147), .B0(n5148), .B1(n5167), .Y(n5168));
NAND4X1  g0537(.A(n5163), .B(n5158_1), .C(n5153_1), .D(n5168), .Y(n5169));
NOR2X1   g0538(.A(n5169), .B(n5150), .Y(n5170));
INVX1    g0539(.A(n5170), .Y(g34383));
INVX1    g0540(.A(g25114), .Y(n5173));
INVX1    g0541(.A(g4349), .Y(n5174));
NAND3X1  g0542(.A(n4956), .B(g4358), .C(n5174), .Y(n5175));
AND2X1   g0543(.A(g3703), .B(g3639), .Y(n5176_1));
INVX1    g0544(.A(n5176_1), .Y(n5177));
NOR2X1   g0545(.A(g4358), .B(g4349), .Y(n5178));
NAND4X1  g0546(.A(n4954_1), .B(n4951), .C(n4949_1), .D(n5178), .Y(n5179));
OAI22X1  g0547(.A0(n5177), .A1(n5175), .B0(n5173), .B1(n5179), .Y(n5180));
INVX1    g0548(.A(g4358), .Y(n5181_1));
NAND3X1  g0549(.A(n4956), .B(n5181_1), .C(g4349), .Y(n5182));
AND2X1   g0550(.A(g3352), .B(g3288), .Y(n5183));
INVX1    g0551(.A(n5183), .Y(n5184));
NAND2X1  g0552(.A(g4358), .B(g4349), .Y(n5185));
OR4X1    g0553(.A(n4955), .B(n4952), .C(n4949_1), .D(n5185), .Y(n5186_1));
AND2X1   g0554(.A(g3990), .B(g4054), .Y(n5187));
INVX1    g0555(.A(n5187), .Y(n5188));
OAI22X1  g0556(.A0(n5186_1), .A1(n5188), .B0(n5184), .B1(n5182), .Y(n5189));
AND2X1   g0557(.A(g6741), .B(g6682), .Y(n5190));
NAND3X1  g0558(.A(n5190), .B(n5178), .C(n4956), .Y(n5191_1));
AND2X1   g0559(.A(g6049), .B(g5990), .Y(n5192));
NAND4X1  g0560(.A(n4957), .B(g4358), .C(n5174), .D(n5192), .Y(n5193));
AND2X1   g0561(.A(g5644), .B(g5703), .Y(n5194));
NAND4X1  g0562(.A(n4957), .B(n5181_1), .C(g4349), .D(n5194), .Y(n5195));
AND2X1   g0563(.A(g6395), .B(g6336), .Y(n5196_1));
NAND4X1  g0564(.A(n4957), .B(g4358), .C(g4349), .D(n5196_1), .Y(n5197));
NAND4X1  g0565(.A(n5195), .B(n5193), .C(n5191_1), .D(n5197), .Y(n5198));
NOR4X1   g0566(.A(n5189), .B(n5180), .C(n4958), .D(n5198), .Y(n5199));
INVX1    g0567(.A(n5199), .Y(g34425));
ZERO     g0568(.Y(g34597));
INVX1    g0569(.A(g4369), .Y(n5202));
INVX1    g0570(.A(g4366), .Y(n5203));
INVX1    g0571(.A(g4332), .Y(n5204));
NOR2X1   g0572(.A(g4311), .B(g4322), .Y(n5205));
INVX1    g0573(.A(g4322), .Y(n5207));
AOI21X1  g0574(.A0(n4957), .A1(n5203), .B0(n5202), .Y(g34839));
NAND2X1  g0575(.A(n5010), .B(g2844), .Y(n5215));
INVX1    g0576(.A(g2848), .Y(n5216_1));
NAND4X1  g0577(.A(n4983), .B(g28), .C(g9), .D(n4996), .Y(n5217));
OR2X1    g0578(.A(n5217), .B(n5216_1), .Y(n5218));
AOI22X1  g0579(.A0(n4998), .A1(g2902), .B0(g2907), .B1(n5000), .Y(n5219));
NAND3X1  g0580(.A(n5219), .B(n5218), .C(n5215), .Y(n5220));
NAND3X1  g0581(.A(n5220), .B(n5072), .C(n4383), .Y(n5221_1));
INVX1    g0582(.A(g632), .Y(n5222));
OR2X1    g0583(.A(n5024), .B(n5019), .Y(n5223));
AOI21X1  g0584(.A0(n5222), .A1(g35), .B0(n5223), .Y(n5224));
INVX1    g0585(.A(g538), .Y(n5225));
NAND3X1  g0586(.A(n5022_1), .B(n4983), .C(n4982), .Y(n5226_1));
NOR2X1   g0587(.A(n5226_1), .B(n5225), .Y(n5227));
INVX1    g0588(.A(g595), .Y(n5228));
OR2X1    g0589(.A(n5024), .B(n5021), .Y(n5229));
AOI21X1  g0590(.A0(n5228), .A1(g35), .B0(n5229), .Y(n5230));
INVX1    g0591(.A(g776), .Y(n5231_1));
AOI21X1  g0592(.A0(n5231_1), .A1(g35), .B0(n5023), .Y(n5232));
OR4X1    g0593(.A(n5230), .B(n5227), .C(n5224), .D(n5232), .Y(n5233));
NAND2X1  g0594(.A(n5233), .B(n5040), .Y(n5234));
INVX1    g0595(.A(g4727), .Y(n5235));
NOR4X1   g0596(.A(n5031), .B(n4987), .C(n5235), .D(n5019), .Y(n5236_1));
INVX1    g0597(.A(g3853), .Y(n5237));
NAND4X1  g0598(.A(n4984_1), .B(n4383), .C(g6199), .D(n5048), .Y(n5238));
OAI21X1  g0599(.A0(n4991), .A1(n5237), .B0(n5238), .Y(n5239));
INVX1    g0600(.A(g45), .Y(n5240));
NAND4X1  g0601(.A(n4981), .B(n4383), .C(g4917), .D(n5050), .Y(n5241_1));
OAI21X1  g0602(.A0(n5062), .A1(n5240), .B0(n5241_1), .Y(n5242));
INVX1    g0603(.A(g1291), .Y(n5243));
NAND2X1  g0604(.A(g1300), .B(n5243), .Y(n5244));
INVX1    g0605(.A(g947), .Y(n5245));
NAND2X1  g0606(.A(n5245), .B(g956), .Y(n5246_1));
OAI22X1  g0607(.A0(n5244), .A1(n5017_1), .B0(n5067), .B1(n5246_1), .Y(n5247));
NOR4X1   g0608(.A(n5242), .B(n5239), .C(n5236_1), .D(n5247), .Y(n5248));
NAND4X1  g0609(.A(n5234), .B(n5221_1), .C(g22), .D(n5248), .Y(g34913));
NOR4X1   g0610(.A(n4993), .B(n4992_1), .C(g31), .D(n4994), .Y(n5250_1));
NAND3X1  g0611(.A(n5250_1), .B(n5048), .C(g28), .Y(n5251));
NAND3X1  g0612(.A(n5016), .B(n5050), .C(g2890), .Y(n5252));
NAND2X1  g0613(.A(n5012_1), .B(g100), .Y(n5253));
INVX1    g0614(.A(g2984), .Y(n5254_1));
OR4X1    g0615(.A(n4995), .B(g28), .C(n5254_1), .D(n5001), .Y(n5255));
NAND4X1  g0616(.A(n5253), .B(n5252), .C(n5251), .D(n5255), .Y(n5256));
NAND2X1  g0617(.A(n5256), .B(n5087), .Y(n5257));
INVX1    g0618(.A(g599), .Y(n5258));
AOI21X1  g0619(.A0(n5258), .A1(g35), .B0(n5223), .Y(n5259_1));
INVX1    g0620(.A(g739), .Y(n5260));
AOI21X1  g0621(.A0(n5260), .A1(g35), .B0(n5023), .Y(n5261));
INVX1    g0622(.A(g562), .Y(n5262));
AOI21X1  g0623(.A0(n5262), .A1(g35), .B0(n5229), .Y(n5263));
NOR2X1   g0624(.A(g781), .B(n4620), .Y(n5264_1));
NAND4X1  g0625(.A(n4983), .B(n4982), .C(g199), .D(n5022_1), .Y(n5265));
OAI21X1  g0626(.A0(n5264_1), .A1(n5027_1), .B0(n5265), .Y(n5266));
OR4X1    g0627(.A(n5263), .B(n5261), .C(n5259_1), .D(n5266), .Y(n5267));
NAND2X1  g0628(.A(n5267), .B(n5040), .Y(n5268));
INVX1    g0629(.A(g2145), .Y(n5269_1));
NOR4X1   g0630(.A(n5019), .B(n4987), .C(n5269_1), .D(n4988_1), .Y(n5270));
INVX1    g0631(.A(g4245), .Y(n5271));
INVX1    g0632(.A(g2704), .Y(n5272));
OAI22X1  g0633(.A0(n4991), .A1(n5272), .B0(n5271), .B1(n5090), .Y(n5273));
INVX1    g0634(.A(g52), .Y(n5274_1));
INVX1    g0635(.A(g4157), .Y(n5275));
OAI22X1  g0636(.A0(n5062), .A1(n5274_1), .B0(n5275), .B1(n5088), .Y(n5276));
INVX1    g0637(.A(g1287), .Y(n5277));
INVX1    g0638(.A(g943), .Y(n5278));
OAI22X1  g0639(.A0(n5017_1), .A1(n5277), .B0(n5278), .B1(n5067), .Y(n5279_1));
NOR4X1   g0640(.A(n5276), .B(n5273), .C(n5270), .D(n5279_1), .Y(n5280));
NAND4X1  g0641(.A(n5268), .B(n5257), .C(g22), .D(n5280), .Y(g34915));
INVX1    g0642(.A(g22), .Y(n5282));
INVX1    g0643(.A(g2999), .Y(n5283));
NOR3X1   g0644(.A(n5006), .B(n5004), .C(n5283), .Y(n5284_1));
NOR2X1   g0645(.A(n5009), .B(n5005), .Y(n5285));
NAND3X1  g0646(.A(n5285), .B(n5250_1), .C(n4982), .Y(n5286));
NAND3X1  g0647(.A(n5285), .B(n5250_1), .C(g28), .Y(n5287));
OAI22X1  g0648(.A0(n5286), .A1(n4787), .B0(n4789), .B1(n5287), .Y(n5288));
NOR2X1   g0649(.A(n5288), .B(n5284_1), .Y(n5289_1));
AOI22X1  g0650(.A0(n5010), .A1(g2852), .B0(g2856), .B1(n5013), .Y(n5290));
AOI21X1  g0651(.A0(n5290), .A1(n5289_1), .B0(n5015), .Y(n5291));
INVX1    g0652(.A(g626), .Y(n5292));
AOI21X1  g0653(.A0(n5292), .A1(g35), .B0(n5223), .Y(n5293));
INVX1    g0654(.A(g772), .Y(n5294_1));
AOI21X1  g0655(.A0(n5294_1), .A1(g35), .B0(n5023), .Y(n5295));
INVX1    g0656(.A(g590), .Y(n5296));
AOI21X1  g0657(.A0(n5296), .A1(g35), .B0(n5229), .Y(n5297));
NOR3X1   g0658(.A(n5297), .B(n5295), .C(n5293), .Y(n5298));
NOR2X1   g0659(.A(n5298), .B(n5030), .Y(n5299_1));
NAND4X1  g0660(.A(n4981), .B(n4383), .C(g4732), .D(n4984_1), .Y(n5300));
AOI22X1  g0661(.A0(n5046), .A1(g3502), .B0(g5853), .B1(n5020), .Y(n5301));
AOI22X1  g0662(.A0(n5032_1), .A1(g4922), .B0(g46), .B1(n5034), .Y(n5302));
INVX1    g0663(.A(g1472), .Y(n5303_1));
NOR2X1   g0664(.A(g1291), .B(n5303_1), .Y(n5304));
INVX1    g0665(.A(g1129), .Y(n5305));
NOR2X1   g0666(.A(g947), .B(n5305), .Y(n5306));
AOI22X1  g0667(.A0(n5304), .A1(n5047_1), .B0(n5033), .B1(n5306), .Y(n5307));
NAND4X1  g0668(.A(n5302), .B(n5301), .C(n5300), .D(n5307), .Y(n5308_1));
OR4X1    g0669(.A(n5299_1), .B(n5291), .C(n5282), .D(n5308_1), .Y(g34917));
NOR3X1   g0670(.A(n5006), .B(n5004), .C(g2994), .Y(n5310));
OAI22X1  g0671(.A0(n5286), .A1(n4786), .B0(n4788_1), .B1(n5287), .Y(n5311));
INVX1    g0672(.A(g2860), .Y(n5312));
INVX1    g0673(.A(g2864), .Y(n5313_1));
NAND4X1  g0674(.A(n4983), .B(n4982), .C(g9), .D(n4996), .Y(n5314));
OAI22X1  g0675(.A0(n5314), .A1(n5312), .B0(n5313_1), .B1(n5217), .Y(n5315));
NOR3X1   g0676(.A(n5315), .B(n5311), .C(n5310), .Y(n5316));
OR2X1    g0677(.A(n5316), .B(n5015), .Y(n5317));
INVX1    g0678(.A(g622), .Y(n5318_1));
AOI21X1  g0679(.A0(n5318_1), .A1(g35), .B0(n5223), .Y(n5319));
INVX1    g0680(.A(g554), .Y(n5320));
AOI21X1  g0681(.A0(n5320), .A1(g35), .B0(n5027_1), .Y(n5321));
INVX1    g0682(.A(g582), .Y(n5322_1));
AOI21X1  g0683(.A0(n5322_1), .A1(g35), .B0(n5229), .Y(n5323));
INVX1    g0684(.A(g546), .Y(n5324));
NOR2X1   g0685(.A(g767), .B(n4620), .Y(n5325));
OAI22X1  g0686(.A0(n5226_1), .A1(n5324), .B0(n5023), .B1(n5325), .Y(n5326_1));
OR4X1    g0687(.A(n5323), .B(n5321), .C(n5319), .D(n5326_1), .Y(n5327));
NAND4X1  g0688(.A(n4981), .B(n4383), .C(g4717), .D(n4984_1), .Y(n5328));
AOI22X1  g0689(.A0(n5046), .A1(g3151), .B0(g5507), .B1(n5020), .Y(n5329));
AOI22X1  g0690(.A0(n5032_1), .A1(g4907), .B0(g47), .B1(n5034), .Y(n5330_1));
INVX1    g0691(.A(g1448), .Y(n5331));
NOR2X1   g0692(.A(g1291), .B(n5331), .Y(n5332));
INVX1    g0693(.A(g1105), .Y(n5333));
NOR2X1   g0694(.A(g947), .B(n5333), .Y(n5334));
AOI22X1  g0695(.A0(n5332), .A1(n5047_1), .B0(n5033), .B1(n5334), .Y(n5335_1));
NAND4X1  g0696(.A(n5330_1), .B(n5329), .C(n5328), .D(n5335_1), .Y(n5336));
AOI21X1  g0697(.A0(n5327), .A1(n5040), .B0(n5336), .Y(n5337));
NAND3X1  g0698(.A(n5337), .B(n5317), .C(g22), .Y(g34919));
NAND4X1  g0699(.A(n5250_1), .B(n4982), .C(g2941), .D(n5285), .Y(n5339));
AOI21X1  g0700(.A0(n5000), .A1(g2936), .B0(n4999), .Y(n5340_1));
INVX1    g0701(.A(g2898), .Y(n5341));
OR2X1    g0702(.A(n5217), .B(n5341), .Y(n5342));
AOI22X1  g0703(.A0(n5007_1), .A1(g2988), .B0(g2894), .B1(n5010), .Y(n5343));
NAND4X1  g0704(.A(n5342), .B(n5340_1), .C(n5339), .D(n5343), .Y(n5344));
INVX1    g0705(.A(g617), .Y(n5345_1));
AOI21X1  g0706(.A0(n5345_1), .A1(g35), .B0(n5223), .Y(n5346));
INVX1    g0707(.A(g807), .Y(n5347));
AOI21X1  g0708(.A0(n5347), .A1(g35), .B0(n5027_1), .Y(n5348));
INVX1    g0709(.A(g577), .Y(n5349));
AOI21X1  g0710(.A0(n5349), .A1(g35), .B0(n5229), .Y(n5350_1));
INVX1    g0711(.A(g542), .Y(n5351));
NOR2X1   g0712(.A(g763), .B(n4620), .Y(n5352));
OAI22X1  g0713(.A0(n5226_1), .A1(n5351), .B0(n5023), .B1(n5352), .Y(n5353));
NOR4X1   g0714(.A(n5350_1), .B(n5348), .C(n5346), .D(n5353), .Y(n5354));
INVX1    g0715(.A(g4912), .Y(n5355_1));
NOR4X1   g0716(.A(n5031), .B(n4987), .C(n5355_1), .D(n5004), .Y(n5356));
INVX1    g0717(.A(g6545), .Y(n5357));
NAND4X1  g0718(.A(n4981), .B(n4383), .C(g4722), .D(n4984_1), .Y(n5358));
OAI21X1  g0719(.A0(n4991), .A1(n5357), .B0(n5358), .Y(n5359));
INVX1    g0720(.A(g48), .Y(n5360_1));
NAND4X1  g0721(.A(n4984_1), .B(n4383), .C(g5160), .D(n5048), .Y(n5361));
OAI21X1  g0722(.A0(n5062), .A1(n5360_1), .B0(n5361), .Y(n5362));
NAND2X1  g0723(.A(n5243), .B(g1478), .Y(n5363));
NAND2X1  g0724(.A(n5245), .B(g1135), .Y(n5364));
OAI22X1  g0725(.A0(n5363), .A1(n5017_1), .B0(n5067), .B1(n5364), .Y(n5365_1));
NOR4X1   g0726(.A(n5362), .B(n5359), .C(n5356), .D(n5365_1), .Y(n5366));
OAI21X1  g0727(.A0(n5354), .A1(n5030), .B0(n5366), .Y(n5367));
AOI21X1  g0728(.A0(n5344), .A1(n5073), .B0(n5367), .Y(n5368));
NAND2X1  g0729(.A(n5368), .B(g22), .Y(g34921));
INVX1    g0730(.A(g2955), .Y(n5370_1));
NOR4X1   g0731(.A(n4995), .B(g28), .C(n5370_1), .D(n4997_1), .Y(n5371));
NAND4X1  g0732(.A(n5250_1), .B(g2950), .C(g28), .D(n5285), .Y(n5372));
NAND2X1  g0733(.A(n5372), .B(n5251), .Y(n5373));
INVX1    g0734(.A(g2882), .Y(n5374));
NOR2X1   g0735(.A(n5217), .B(n5374), .Y(n5375_1));
NAND3X1  g0736(.A(n5016), .B(n5050), .C(g2868), .Y(n5376));
OR4X1    g0737(.A(n4990), .B(g23002), .C(n4982), .D(n5006), .Y(n5377));
NAND2X1  g0738(.A(n5377), .B(n5376), .Y(n5378));
OR4X1    g0739(.A(n5375_1), .B(n5373), .C(n5371), .D(n5378), .Y(n5379));
NAND2X1  g0740(.A(n5379), .B(n5087), .Y(n5380_1));
INVX1    g0741(.A(g613), .Y(n5381));
AOI21X1  g0742(.A0(n5381), .A1(g35), .B0(n5223), .Y(n5382));
INVX1    g0743(.A(g794), .Y(n5383));
AOI21X1  g0744(.A0(n5383), .A1(g35), .B0(n5027_1), .Y(n5384));
INVX1    g0745(.A(g586), .Y(n5385_1));
AOI21X1  g0746(.A0(n5385_1), .A1(g35), .B0(n5229), .Y(n5386));
INVX1    g0747(.A(g534), .Y(n5387));
NOR2X1   g0748(.A(g758), .B(n4620), .Y(n5388));
OAI22X1  g0749(.A0(n5226_1), .A1(n5387), .B0(n5023), .B1(n5388), .Y(n5389));
OR4X1    g0750(.A(n5386), .B(n5384), .C(n5382), .D(n5389), .Y(n5390_1));
NAND4X1  g0751(.A(n5048), .B(n4383), .C(g4300), .D(n5050), .Y(n5391));
INVX1    g0752(.A(n5391), .Y(n5392));
INVX1    g0753(.A(g4172), .Y(n5393));
OAI22X1  g0754(.A0(n5051_1), .A1(g4927), .B0(n5393), .B1(n5088), .Y(n5394));
INVX1    g0755(.A(g49), .Y(n5395_1));
OAI22X1  g0756(.A0(n4985), .A1(g4737), .B0(n5395_1), .B1(n5062), .Y(n5396));
OAI22X1  g0757(.A0(n5017_1), .A1(n5243), .B0(n5245), .B1(n5067), .Y(n5397));
OR4X1    g0758(.A(n5396), .B(n5394), .C(n5392), .D(n5397), .Y(n5398));
AOI21X1  g0759(.A0(n5390_1), .A1(n5040), .B0(n5398), .Y(n5399));
NAND3X1  g0760(.A(n5399), .B(n5380_1), .C(g22), .Y(g34923));
NAND3X1  g0761(.A(n5016), .B(n5050), .C(g2873), .Y(n5401));
AOI22X1  g0762(.A0(n4998), .A1(g2965), .B0(g2960), .B1(n5000), .Y(n5402));
AOI22X1  g0763(.A0(n5012_1), .A1(g94), .B0(g2878), .B1(n5013), .Y(n5403));
NAND3X1  g0764(.A(n5403), .B(n5402), .C(n5401), .Y(n5404));
AND2X1   g0765(.A(n5404), .B(n5087), .Y(n5405_1));
INVX1    g0766(.A(g608), .Y(n5406));
AOI21X1  g0767(.A0(n5406), .A1(g35), .B0(n5223), .Y(n5407));
INVX1    g0768(.A(g790), .Y(n5408));
AOI21X1  g0769(.A0(n5408), .A1(g35), .B0(n5027_1), .Y(n5409));
INVX1    g0770(.A(g572), .Y(n5410_1));
AOI21X1  g0771(.A0(n5410_1), .A1(g35), .B0(n5229), .Y(n5411));
NOR2X1   g0772(.A(g749), .B(n4620), .Y(n5412));
OAI22X1  g0773(.A0(n5226_1), .A1(g550), .B0(n5023), .B1(n5412), .Y(n5413));
NOR4X1   g0774(.A(n5411), .B(n5409), .C(n5407), .D(n5413), .Y(n5414));
INVX1    g0775(.A(g2130), .Y(n5415_1));
NOR4X1   g0776(.A(n5019), .B(n4987), .C(n5415_1), .D(n4988_1), .Y(n5416));
INVX1    g0777(.A(g2689), .Y(n5417));
NAND4X1  g0778(.A(n5048), .B(n4383), .C(g4253), .D(n5050), .Y(n5418));
OAI21X1  g0779(.A0(n4991), .A1(n5417), .B0(n5418), .Y(n5419));
INVX1    g0780(.A(g50), .Y(n5420_1));
NAND3X1  g0781(.A(n5010), .B(n4383), .C(g4176), .Y(n5421));
OAI21X1  g0782(.A0(n5062), .A1(n5420_1), .B0(n5421), .Y(n5422));
OAI22X1  g0783(.A0(n5017_1), .A1(g1296), .B0(g952), .B1(n5067), .Y(n5423));
NOR4X1   g0784(.A(n5422), .B(n5419), .C(n5416), .D(n5423), .Y(n5424));
OAI21X1  g0785(.A0(n5414), .A1(n5030), .B0(n5424), .Y(n5425_1));
OR2X1    g0786(.A(n5425_1), .B(n5405_1), .Y(n6708));
OR2X1    g0787(.A(n6708), .B(n5282), .Y(g34925));
INVX1    g0788(.A(g2980), .Y(n5428));
OR4X1    g0789(.A(n4995), .B(g28), .C(n5428), .D(n5001), .Y(n5429));
AOI22X1  g0790(.A0(n4998), .A1(g2975), .B0(g2970), .B1(n5000), .Y(n5430_1));
INVX1    g0791(.A(g2886), .Y(n5431));
OR2X1    g0792(.A(n5217), .B(n5431), .Y(n5432));
AOI22X1  g0793(.A0(n5007_1), .A1(g127), .B0(g92), .B1(n5012_1), .Y(n5433));
NAND4X1  g0794(.A(n5432), .B(n5430_1), .C(n5429), .D(n5433), .Y(n5434));
AND2X1   g0795(.A(n5434), .B(n5087), .Y(n5435_1));
INVX1    g0796(.A(g604), .Y(n5436));
AOI21X1  g0797(.A0(n5436), .A1(g35), .B0(n5223), .Y(n5437));
INVX1    g0798(.A(g785), .Y(n5438));
AOI21X1  g0799(.A0(n5438), .A1(g35), .B0(n5027_1), .Y(n5439));
INVX1    g0800(.A(g568), .Y(n5440_1));
AOI21X1  g0801(.A0(n5440_1), .A1(g35), .B0(n5229), .Y(n5441));
NOR2X1   g0802(.A(g744), .B(n4620), .Y(n5442));
OAI22X1  g0803(.A0(n5226_1), .A1(g23612), .B0(n5023), .B1(n5442), .Y(n5443));
NOR4X1   g0804(.A(n5441), .B(n5439), .C(n5437), .D(n5443), .Y(n5444));
INVX1    g0805(.A(g2138), .Y(n5445_1));
NOR4X1   g0806(.A(n5019), .B(n4987), .C(n5445_1), .D(n4988_1), .Y(n5446));
INVX1    g0807(.A(g2697), .Y(n5447));
NAND4X1  g0808(.A(n5048), .B(n4383), .C(g4249), .D(n5050), .Y(n5448));
OAI21X1  g0809(.A0(n4991), .A1(n5447), .B0(n5448), .Y(n5449));
INVX1    g0810(.A(g51), .Y(n5450_1));
NAND3X1  g0811(.A(n5010), .B(n4383), .C(g4146), .Y(n5451));
OAI21X1  g0812(.A0(n5062), .A1(n5450_1), .B0(n5451), .Y(n5452));
INVX1    g0813(.A(g939), .Y(n5453));
INVX1    g0814(.A(g1283), .Y(n5454));
OAI22X1  g0815(.A0(n5017_1), .A1(n5454), .B0(n5453), .B1(n5067), .Y(n5455_1));
NOR4X1   g0816(.A(n5452), .B(n5449), .C(n5446), .D(n5455_1), .Y(n5456));
OAI21X1  g0817(.A0(n5444), .A1(n5030), .B0(n5456), .Y(n5457));
OR2X1    g0818(.A(n5457), .B(n5435_1), .Y(n4586));
OR2X1    g0819(.A(n4586), .B(n5282), .Y(g34927));
NAND3X1  g0820(.A(n5280), .B(n5268), .C(n5257), .Y(n3220));
XOR2X1   g0821(.A(n4586), .B(n3220), .Y(n5461));
AND2X1   g0822(.A(n5399), .B(n5380_1), .Y(n5462));
XOR2X1   g0823(.A(n6708), .B(n5462), .Y(n5463_1));
XOR2X1   g0824(.A(n5463_1), .B(n5461), .Y(n5464));
AND2X1   g0825(.A(n5337), .B(n5317), .Y(n5465));
XOR2X1   g0826(.A(n5368), .B(n5465), .Y(n5466));
NAND3X1  g0827(.A(n5248), .B(n5234), .C(n5221_1), .Y(n3747));
NOR3X1   g0828(.A(n5308_1), .B(n5299_1), .C(n5291), .Y(n5468));
XOR2X1   g0829(.A(n5468), .B(n3747), .Y(n5469));
XOR2X1   g0830(.A(n5469), .B(n5466), .Y(n5470));
XOR2X1   g0831(.A(n5470), .B(n5464), .Y(n5471));
OAI21X1  g0832(.A0(n4976), .A1(g56), .B0(g55), .Y(n5472_1));
XOR2X1   g0833(.A(n5472_1), .B(n5471), .Y(n5962));
OR2X1    g0834(.A(n5962), .B(n5282), .Y(g34972));
INVX1    g0835(.A(g5), .Y(g12833));
INVX1    g0836(.A(g5057), .Y(n5476));
INVX1    g0837(.A(g5052), .Y(n5477_1));
INVX1    g0838(.A(g5046), .Y(n5478));
INVX1    g0839(.A(g5029), .Y(n5479));
INVX1    g0840(.A(g5062), .Y(n5480));
INVX1    g0841(.A(g5033), .Y(n5481));
INVX1    g0842(.A(g5016), .Y(n5482_1));
NOR4X1   g0843(.A(n5481), .B(n5480), .C(n5479), .D(n5482_1), .Y(n5483));
NAND3X1  g0844(.A(n5483), .B(g5041), .C(g5037), .Y(n5484));
NOR2X1   g0845(.A(n5484), .B(n5478), .Y(n5485));
INVX1    g0846(.A(g5037), .Y(n5486));
INVX1    g0847(.A(g5041), .Y(n5487_1));
INVX1    g0848(.A(g5022), .Y(n5488));
NOR4X1   g0849(.A(g5033), .B(g5029), .C(n5488), .D(g5016), .Y(n5489));
NAND3X1  g0850(.A(n5489), .B(n5487_1), .C(n5486), .Y(n5490));
NOR2X1   g0851(.A(n5490), .B(g5046), .Y(n5491));
MX2X1    g0852(.A(n5485), .B(n5491), .S0(n5477_1), .Y(n5492_1));
NOR2X1   g0853(.A(n5480), .B(g5057), .Y(n5493));
NOR3X1   g0854(.A(n5478), .B(n5477_1), .C(g84), .Y(n5494));
INVX1    g0855(.A(g84), .Y(n5495));
NOR3X1   g0856(.A(n5478), .B(n5487_1), .C(n5495), .Y(n5496));
OAI21X1  g0857(.A0(n5496), .A1(n5494), .B0(n5493), .Y(n5497_1));
AND2X1   g0858(.A(g5022), .B(g5057), .Y(n5498));
NAND4X1  g0859(.A(n5478), .B(n5487_1), .C(g84), .D(n5498), .Y(n5499));
NAND4X1  g0860(.A(n5478), .B(n5477_1), .C(n5495), .D(n5498), .Y(n5500));
NAND3X1  g0861(.A(n5500), .B(n5499), .C(n5497_1), .Y(n5501));
NOR2X1   g0862(.A(n5501), .B(n5476), .Y(n5502_1));
MX2X1    g0863(.A(n5502_1), .B(n5476), .S0(n5492_1), .Y(n5503));
MX2X1    g0864(.A(g5052), .B(n5503), .S0(g35), .Y(n685));
INVX1    g0865(.A(g2771), .Y(n5505));
NOR2X1   g0866(.A(n4809), .B(g113), .Y(n5506));
AND2X1   g0867(.A(n5506), .B(g85), .Y(n5507_1));
INVX1    g0868(.A(g2735), .Y(n5508));
NOR4X1   g0869(.A(n4909), .B(n4915_1), .C(n4910_1), .D(n5508), .Y(n5509));
NOR2X1   g0870(.A(g2729), .B(g2724), .Y(n5510));
AND2X1   g0871(.A(n5510), .B(n5509), .Y(n5511_1));
INVX1    g0872(.A(g2767), .Y(n5512));
OAI21X1  g0873(.A0(n5506), .A1(n5512), .B0(n5511_1), .Y(n5513));
OAI22X1  g0874(.A0(n5511_1), .A1(n5505), .B0(n5507_1), .B1(n5513), .Y(n5514));
MX2X1    g0875(.A(g2775), .B(n5514), .S0(g35), .Y(n690));
INVX1    g0876(.A(g691), .Y(n5516_1));
NOR2X1   g0877(.A(n5516_1), .B(g209), .Y(n5517));
AOI21X1  g0878(.A0(n5517), .A1(n4709), .B0(g134), .Y(n5518));
NAND2X1  g0879(.A(g2138), .B(g2130), .Y(n5519));
NOR2X1   g0880(.A(n5519), .B(g2145), .Y(n5520));
NOR3X1   g0881(.A(n5520), .B(n5518), .C(n5306), .Y(n5521_1));
INVX1    g0882(.A(g1242), .Y(n5522));
OR4X1    g0883(.A(n5518), .B(n5306), .C(n5522), .D(n5520), .Y(n5523));
INVX1    g0884(.A(g4180), .Y(n5524));
NOR3X1   g0885(.A(n5518), .B(n5306), .C(n5524), .Y(n5525));
OAI21X1  g0886(.A0(n5525), .A1(n5521_1), .B0(n5523), .Y(n5526_1));
INVX1    g0887(.A(g1862), .Y(n5527));
INVX1    g0888(.A(n4664), .Y(n5528));
NAND4X1  g0889(.A(g979), .B(g1183), .C(g1171), .D(g1061), .Y(n5529));
OAI21X1  g0890(.A0(n5529), .A1(n5528), .B0(g1083), .Y(n5530));
AND2X1   g0891(.A(n5530), .B(n5521_1), .Y(n5531_1));
NOR3X1   g0892(.A(n5531_1), .B(n5161), .C(n5527), .Y(n5532));
MX2X1    g0893(.A(g1882), .B(n5526_1), .S0(n5532), .Y(n5533));
MX2X1    g0894(.A(g1886), .B(n5533), .S0(g35), .Y(n695));
INVX1    g0895(.A(g6459), .Y(n5535));
NOR2X1   g0896(.A(g6455), .B(n5535), .Y(n5536_1));
NOR2X1   g0897(.A(g6451), .B(n5535), .Y(n5537));
MX2X1    g0898(.A(n5536_1), .B(n5537), .S0(g6466), .Y(n5538));
MX2X1    g0899(.A(g6459), .B(n5538), .S0(g35), .Y(n700));
INVX1    g0900(.A(g1585), .Y(n5540));
NOR4X1   g0901(.A(n5516_1), .B(n4711), .C(g209), .D(n4712_1), .Y(n5541_1));
OAI22X1  g0902(.A0(g1291), .A1(n5331), .B0(g134), .B1(n5541_1), .Y(n5542));
NAND2X1  g0903(.A(g2704), .B(g2689), .Y(n5543));
NOR2X1   g0904(.A(n5543), .B(g2697), .Y(n5544));
NOR2X1   g0905(.A(n5544), .B(n5542), .Y(n5545));
OR2X1    g0906(.A(n5542), .B(n5524), .Y(n5546_1));
MX2X1    g0907(.A(n5546_1), .B(n5540), .S0(n5545), .Y(n5547));
OR4X1    g0908(.A(g1559), .B(g1554), .C(g1564), .D(g1548), .Y(n5548));
INVX1    g0909(.A(g1514), .Y(n5549));
NAND4X1  g0910(.A(g1322), .B(g1404), .C(g1526), .D(n5549), .Y(n5550));
OAI21X1  g0911(.A0(n5550), .A1(n5548), .B0(g1422), .Y(n5551_1));
AND2X1   g0912(.A(n5551_1), .B(n5545), .Y(n5552));
NOR3X1   g0913(.A(n5552), .B(g2361), .C(g2287), .Y(n5553));
MX2X1    g0914(.A(g2299), .B(n5547), .S0(n5553), .Y(n5554));
MX2X1    g0915(.A(g2380), .B(n5554), .S0(g35), .Y(n705));
INVX1    g0916(.A(g3969), .Y(n5556));
INVX1    g0917(.A(g3983), .Y(n5557));
NAND2X1  g0918(.A(g4005), .B(g4012), .Y(n5558));
NOR3X1   g0919(.A(n5558), .B(n5557), .C(n5556), .Y(n5559));
XOR2X1   g0920(.A(n5559), .B(g4040), .Y(n5560_1));
MX2X1    g0921(.A(g4031), .B(n5560_1), .S0(g35), .Y(n710));
INVX1    g0922(.A(g2453), .Y(n5562));
INVX1    g0923(.A(g2815), .Y(n5563));
INVX1    g0924(.A(n5510), .Y(n5564_1));
OR2X1    g0925(.A(g2748), .B(g2756), .Y(n5565));
NOR3X1   g0926(.A(n5565), .B(n5508), .C(g2741), .Y(n5566));
AOI21X1  g0927(.A0(n5566), .A1(n5563), .B0(n5564_1), .Y(n5567));
INVX1    g0928(.A(g2715), .Y(n5568_1));
NAND2X1  g0929(.A(n5568_1), .B(g2719), .Y(n5569));
NOR4X1   g0930(.A(n5567), .B(n5562), .C(n4929), .D(n5569), .Y(n5570));
MX2X1    g0931(.A(g2547), .B(g2541), .S0(n5570), .Y(n5571));
MX2X1    g0932(.A(g2541), .B(n5571), .S0(g35), .Y(n715));
INVX1    g0933(.A(g3050), .Y(n5573_1));
NOR2X1   g0934(.A(g3045), .B(n5573_1), .Y(n5574));
INVX1    g0935(.A(g3040), .Y(n5575));
INVX1    g0936(.A(g3034), .Y(n5576));
NOR3X1   g0937(.A(n5576), .B(n5575), .C(g84), .Y(n5577));
INVX1    g0938(.A(g3029), .Y(n5578_1));
NOR3X1   g0939(.A(n5576), .B(n5578_1), .C(n5495), .Y(n5579));
OAI21X1  g0940(.A0(n5579), .A1(n5577), .B0(n5574), .Y(n5580));
AND2X1   g0941(.A(g3045), .B(g3010), .Y(n5581));
NAND4X1  g0942(.A(n5576), .B(n5578_1), .C(g84), .D(n5581), .Y(n5582));
NAND4X1  g0943(.A(n5576), .B(n5575), .C(n5495), .D(n5581), .Y(n5583_1));
NAND3X1  g0944(.A(n5583_1), .B(n5582), .C(n5580), .Y(n5584));
INVX1    g0945(.A(g3017), .Y(n5585));
MX2X1    g0946(.A(g3010), .B(g3050), .S0(g3004), .Y(n5586));
OR2X1    g0947(.A(n5586), .B(n5585), .Y(n5587_1));
NAND2X1  g0948(.A(n5586), .B(n5585), .Y(n5588));
OAI21X1  g0949(.A0(n5587_1), .A1(n5584), .B0(n5588), .Y(n5589));
MX2X1    g0950(.A(g3004), .B(n5589), .S0(g35), .Y(n725));
NOR2X1   g0951(.A(n5524), .B(g4284), .Y(n5591));
INVX1    g0952(.A(n5591), .Y(n5592_1));
INVX1    g0953(.A(g3161), .Y(n5593));
NAND2X1  g0954(.A(g3171), .B(g3179), .Y(n5594));
NOR3X1   g0955(.A(n5594), .B(n5593), .C(g3155), .Y(n5595));
MX2X1    g0956(.A(g3243), .B(n5592_1), .S0(n5595), .Y(n5596));
MX2X1    g0957(.A(g3227), .B(n5596), .S0(g35), .Y(n730));
INVX1    g0958(.A(g358), .Y(n5598));
INVX1    g0959(.A(g376), .Y(n5599));
INVX1    g0960(.A(g385), .Y(n5600));
NOR4X1   g0961(.A(n5599), .B(g370), .C(n5598), .D(n5600), .Y(n5601));
MX2X1    g0962(.A(g452), .B(g460), .S0(n5601), .Y(n5602_1));
MX2X1    g0963(.A(g460), .B(n5602_1), .S0(g35), .Y(n735));
MX2X1    g0964(.A(g464), .B(g471), .S0(n5601), .Y(n5604));
MX2X1    g0965(.A(g471), .B(n5604), .S0(g35), .Y(n740));
NOR3X1   g0966(.A(g3518), .B(g3506), .C(g3512), .Y(n5606));
NAND3X1  g0967(.A(n5606), .B(g3522), .C(n4833), .Y(n5607_1));
MX2X1    g0968(.A(n5592_1), .B(g3542), .S0(n5607_1), .Y(n5608));
MX2X1    g0969(.A(g3546), .B(n5608), .S0(g35), .Y(n745));
INVX1    g0970(.A(g5164), .Y(n5610));
NOR4X1   g0971(.A(n4643), .B(n5610), .C(g5180), .D(g5170), .Y(n5611_1));
MX2X1    g0972(.A(g5232), .B(n5592_1), .S0(n5611_1), .Y(n5612));
MX2X1    g0973(.A(g5208), .B(n5612), .S0(g35), .Y(n750));
MX2X1    g0974(.A(g5813), .B(g5849), .S0(n4863), .Y(n5614));
MX2X1    g0975(.A(g5849), .B(n5614), .S0(g35), .Y(n755));
INVX1    g0976(.A(g12), .Y(n5616));
NOR4X1   g0977(.A(n4995), .B(n5616), .C(n4982), .D(n4997_1), .Y(n5617));
MX2X1    g0978(.A(g2907), .B(n3747), .S0(n5617), .Y(n5618));
MX2X1    g0979(.A(g2984), .B(n5618), .S0(g35), .Y(n760));
NOR3X1   g0980(.A(g2138), .B(n5415_1), .C(n5269_1), .Y(n5620_1));
NOR3X1   g0981(.A(n5620_1), .B(n5518), .C(n5334), .Y(n5621));
OR4X1    g0982(.A(n5518), .B(n5334), .C(g1242), .D(n5620_1), .Y(n5622));
NOR3X1   g0983(.A(n5518), .B(n5334), .C(n5524), .Y(n5623));
OAI21X1  g0984(.A0(n5623), .A1(n5621), .B0(n5622), .Y(n5624));
INVX1    g0985(.A(g1772), .Y(n5625_1));
NAND4X1  g0986(.A(g979), .B(g1183), .C(n4665), .D(g1061), .Y(n5626));
OAI21X1  g0987(.A0(n5626), .A1(n5528), .B0(g1079), .Y(n5627));
AND2X1   g0988(.A(n5627), .B(n5621), .Y(n5628));
NOR3X1   g0989(.A(n5628), .B(n5625_1), .C(g1802), .Y(n5629));
MX2X1    g0990(.A(g1744), .B(n5624), .S0(n5629), .Y(n5630_1));
MX2X1    g0991(.A(g1736), .B(n5630_1), .S0(g35), .Y(n765));
NOR3X1   g0992(.A(g5857), .B(g5863), .C(g5869), .Y(n5632));
NAND3X1  g0993(.A(n5632), .B(g5881), .C(g5873), .Y(n5633));
MX2X1    g0994(.A(n5592_1), .B(g5909), .S0(n5633), .Y(n5634));
MX2X1    g0995(.A(g5913), .B(n5634), .S0(g35), .Y(n770));
INVX1    g0996(.A(n5628), .Y(n5636));
INVX1    g0997(.A(n4809), .Y(n5637));
NAND4X1  g0998(.A(n5637), .B(g112), .C(n4824), .D(n5147), .Y(n5638));
NAND3X1  g0999(.A(n5638), .B(n5636), .C(g1772), .Y(n5639));
OAI21X1  g1000(.A0(n5636), .A1(n5164), .B0(n5639), .Y(n5640_1));
MX2X1    g1001(.A(g1772), .B(n5640_1), .S0(g35), .Y(n775));
NOR3X1   g1002(.A(n4835), .B(n4834), .C(g3530), .Y(n5642));
MX2X1    g1003(.A(g3554), .B(n5592_1), .S0(n5642), .Y(n5643));
MX2X1    g1004(.A(g3602), .B(n5643), .S0(g35), .Y(n780));
NAND3X1  g1005(.A(n5637), .B(g43), .C(n4824), .Y(n5645_1));
NOR3X1   g1006(.A(n5645_1), .B(n4858), .C(n4840), .Y(n5646));
NAND2X1  g1007(.A(g6215), .B(n4871_1), .Y(n5647));
NAND2X1  g1008(.A(n4872), .B(g6219), .Y(n5648));
AOI21X1  g1009(.A0(n5648), .A1(n5647), .B0(n5646), .Y(n5649));
MX2X1    g1010(.A(g6215), .B(n5649), .S0(g35), .Y(n785));
INVX1    g1011(.A(g802), .Y(n5651));
NOR2X1   g1012(.A(n5651), .B(g736), .Y(n5652));
INVX1    g1013(.A(g781), .Y(n5653));
NAND2X1  g1014(.A(n5651), .B(g799), .Y(n5654));
INVX1    g1015(.A(n5601), .Y(n5655_1));
NOR2X1   g1016(.A(g499), .B(g518), .Y(n5656));
NAND4X1  g1017(.A(n5130_1), .B(n5142), .C(n5132), .D(n5656), .Y(n5657));
NOR3X1   g1018(.A(g655), .B(g753), .C(g718), .Y(n5658));
NAND3X1  g1019(.A(g655), .B(g753), .C(g718), .Y(n5659));
OAI21X1  g1020(.A0(n5320), .A1(n5347), .B0(n5659), .Y(n5660_1));
NOR4X1   g1021(.A(n5658), .B(n5657), .C(n5655_1), .D(n5660_1), .Y(n5661));
INVX1    g1022(.A(g736), .Y(n5662));
AOI21X1  g1023(.A0(g802), .A1(n5662), .B0(n5260), .Y(n5663));
INVX1    g1024(.A(g744), .Y(n5664));
AOI21X1  g1025(.A0(g802), .A1(n5662), .B0(n5664), .Y(n5665_1));
NAND4X1  g1026(.A(n5663), .B(n5661), .C(n5654), .D(n5665_1), .Y(n5666));
INVX1    g1027(.A(g749), .Y(n5667));
AOI21X1  g1028(.A0(g802), .A1(n5662), .B0(n5667), .Y(n5668));
INVX1    g1029(.A(n5668), .Y(n5669_1));
INVX1    g1030(.A(g758), .Y(n5670));
AOI21X1  g1031(.A0(g802), .A1(n5662), .B0(n5670), .Y(n5671));
INVX1    g1032(.A(n5671), .Y(n5672));
NOR3X1   g1033(.A(n5672), .B(n5669_1), .C(n5666), .Y(n5673));
INVX1    g1034(.A(g763), .Y(n5674_1));
AOI21X1  g1035(.A0(g802), .A1(n5662), .B0(n5674_1), .Y(n5675));
INVX1    g1036(.A(g767), .Y(n5676));
AOI21X1  g1037(.A0(g802), .A1(n5662), .B0(n5676), .Y(n5677));
AOI21X1  g1038(.A0(g802), .A1(n5662), .B0(n5294_1), .Y(n5678));
NAND4X1  g1039(.A(n5677), .B(n5675), .C(n5673), .D(n5678), .Y(n5679_1));
OR4X1    g1040(.A(n5652), .B(n5653), .C(n5231_1), .D(n5679_1), .Y(n5680));
NOR4X1   g1041(.A(n5652), .B(n5408), .C(n5438), .D(n5680), .Y(n5681));
AOI21X1  g1042(.A0(g802), .A1(n5662), .B0(n5383), .Y(n5682));
NAND2X1  g1043(.A(n5682), .B(n5681), .Y(n5683));
AOI21X1  g1044(.A0(g802), .A1(n5662), .B0(n5347), .Y(n5684_1));
MX2X1    g1045(.A(n5347), .B(n5684_1), .S0(n5683), .Y(n5685));
MX2X1    g1046(.A(g794), .B(n5685), .S0(g35), .Y(n790));
INVX1    g1047(.A(g370), .Y(n5687));
NOR4X1   g1048(.A(n5599), .B(n5687), .C(n5598), .D(n5600), .Y(n5688));
MX2X1    g1049(.A(g847), .B(g854), .S0(n5688), .Y(n5689_1));
MX2X1    g1050(.A(g854), .B(n5689_1), .S0(g35), .Y(n800));
INVX1    g1051(.A(g1227), .Y(n5691));
NOR3X1   g1052(.A(g1061), .B(n5691), .C(g1052), .Y(n5692));
NOR2X1   g1053(.A(n4667_1), .B(g1227), .Y(n5693));
OAI21X1  g1054(.A0(n5693), .A1(n5692), .B0(g1056), .Y(n5694_1));
MX2X1    g1055(.A(g1061), .B(n5694_1), .S0(g35), .Y(n805));
INVX1    g1056(.A(n5462), .Y(n2447));
NOR2X1   g1057(.A(n5314), .B(n5616), .Y(n5697));
OAI21X1  g1058(.A0(g4153), .A1(g4172), .B0(g35), .Y(n5698));
AOI21X1  g1059(.A0(n5697), .A1(n2447), .B0(n5698), .Y(n810));
INVX1    g1060(.A(g2994), .Y(n5700));
NOR2X1   g1061(.A(g73), .B(g72), .Y(n5701));
INVX1    g1062(.A(n5701), .Y(n5702));
AOI21X1  g1063(.A0(n5700), .A1(g90), .B0(n5702), .Y(n5703));
NOR2X1   g1064(.A(n5703), .B(g4311), .Y(n5704_1));
OAI21X1  g1065(.A0(n5703), .A1(n4949_1), .B0(n5207), .Y(n5705));
NOR2X1   g1066(.A(n5705), .B(n5704_1), .Y(n5706));
AOI21X1  g1067(.A0(n5701), .A1(g4515), .B0(g4311), .Y(n5707));
AOI21X1  g1068(.A0(n5701), .A1(g4515), .B0(n4949_1), .Y(n5708));
NOR3X1   g1069(.A(n5708), .B(n5707), .C(n5207), .Y(n5709_1));
NOR3X1   g1070(.A(n5709_1), .B(n5706), .C(g4332), .Y(n5710));
NOR3X1   g1071(.A(n4949_1), .B(g4322), .C(n5204), .Y(n5711));
NOR4X1   g1072(.A(n5710), .B(g4349), .C(g4340), .D(n5711), .Y(n5712));
INVX1    g1073(.A(g4340), .Y(n5713_1));
INVX1    g1074(.A(g4584), .Y(n5714));
AOI21X1  g1075(.A0(g4608), .A1(n5714), .B0(g4616), .Y(n5715));
INVX1    g1076(.A(g4608), .Y(n5716));
XOR2X1   g1077(.A(g4601), .B(g4593), .Y(n5717));
AOI21X1  g1078(.A0(n5716), .A1(g4584), .B0(n5717), .Y(n5718_1));
NAND2X1  g1079(.A(n5718_1), .B(n5715), .Y(n5719));
INVX1    g1080(.A(g4593), .Y(n5720));
NOR4X1   g1081(.A(g4608), .B(n5714), .C(n5720), .D(g4601), .Y(n5721));
NOR3X1   g1082(.A(n5716), .B(g4584), .C(g4593), .Y(n5722));
NOR2X1   g1083(.A(n5722), .B(n5721), .Y(n5723_1));
AOI21X1  g1084(.A0(n5723_1), .A1(n5719), .B0(g135), .Y(n5724));
AOI21X1  g1085(.A0(n5724), .A1(n5713_1), .B0(n5174), .Y(n5725));
OR2X1    g1086(.A(n5725), .B(g4358), .Y(n5726));
AOI21X1  g1087(.A0(n5724), .A1(n5713_1), .B0(g4349), .Y(n5727));
NOR3X1   g1088(.A(n5724), .B(n5174), .C(g4340), .Y(n5728_1));
OR2X1    g1089(.A(n5728_1), .B(n5181_1), .Y(n5729));
OAI22X1  g1090(.A0(n5727), .A1(n5729), .B0(n5726), .B1(n5712), .Y(n5730));
MX2X1    g1091(.A(g4366), .B(n5730), .S0(g35), .Y(n815));
NOR3X1   g1092(.A(n5645_1), .B(n4831), .C(g4087), .Y(n5732));
INVX1    g1093(.A(g3512), .Y(n5733_1));
NAND2X1  g1094(.A(g3506), .B(n5733_1), .Y(n5734));
INVX1    g1095(.A(g3506), .Y(n5735));
NAND2X1  g1096(.A(n5735), .B(g3512), .Y(n5736));
AOI21X1  g1097(.A0(n5736), .A1(n5734), .B0(n5732), .Y(n5737));
MX2X1    g1098(.A(g3506), .B(n5737), .S0(g35), .Y(n820));
MX2X1    g1099(.A(n5667), .B(n5668), .S0(n5666), .Y(n5739));
MX2X1    g1100(.A(g744), .B(n5739), .S0(g35), .Y(n825));
MX2X1    g1101(.A(g3490), .B(g3484), .S0(n4836_1), .Y(n5741));
MX2X1    g1102(.A(g3484), .B(n5741), .S0(g35), .Y(n830));
INVX1    g1103(.A(g5969), .Y(n5743_1));
INVX1    g1104(.A(g5983), .Y(n5744));
OAI22X1  g1105(.A0(n5744), .A1(g6005), .B0(n5743_1), .B1(g6012), .Y(n5745));
MX2X1    g1106(.A(g6000), .B(n5743_1), .S0(g5976), .Y(n5746));
INVX1    g1107(.A(g6005), .Y(n5747));
INVX1    g1108(.A(g6012), .Y(n5748_1));
NOR4X1   g1109(.A(n5744), .B(n5743_1), .C(n5747), .D(n5748_1), .Y(n5749));
OAI21X1  g1110(.A0(n5748_1), .A1(g5983), .B0(g35), .Y(n5750));
NOR4X1   g1111(.A(n5749), .B(n5746), .C(n5745), .D(n5750), .Y(n835));
INVX1    g1112(.A(n5518), .Y(n5752));
NAND3X1  g1113(.A(n5445_1), .B(g2130), .C(n5269_1), .Y(n5753_1));
NAND3X1  g1114(.A(n5753_1), .B(n5752), .C(n5364), .Y(n5754));
NAND3X1  g1115(.A(n5752), .B(n5364), .C(g4180), .Y(n5755));
MX2X1    g1116(.A(g1242), .B(n5755), .S0(n5754), .Y(n5756));
INVX1    g1117(.A(g1592), .Y(n5757));
NOR2X1   g1118(.A(n5754), .B(g27831), .Y(n5758_1));
NOR3X1   g1119(.A(n5758_1), .B(g1636), .C(n5757), .Y(n5759));
MX2X1    g1120(.A(g1600), .B(n5756), .S0(n5759), .Y(n5760));
MX2X1    g1121(.A(g1604), .B(n5760), .S0(g35), .Y(n845));
NOR3X1   g1122(.A(n5758_1), .B(g1592), .C(g1668), .Y(n5762));
XOR2X1   g1123(.A(n5762), .B(g1714), .Y(n5763_1));
MX2X1    g1124(.A(g1710), .B(n5763_1), .S0(g35), .Y(n850));
NOR3X1   g1125(.A(n5645_1), .B(n4841_1), .C(n4840), .Y(n5765));
NOR4X1   g1126(.A(g3167), .B(g3155), .C(n4620), .D(n5765), .Y(n860));
INVX1    g1127(.A(g3401), .Y(n5767));
NOR2X1   g1128(.A(n5767), .B(g3396), .Y(n5768_1));
INVX1    g1129(.A(g3385), .Y(n5769));
INVX1    g1130(.A(g3391), .Y(n5770));
NOR3X1   g1131(.A(n5770), .B(n5769), .C(g84), .Y(n5771));
INVX1    g1132(.A(g3380), .Y(n5772));
NOR3X1   g1133(.A(n5769), .B(n5772), .C(n5495), .Y(n5773_1));
OAI21X1  g1134(.A0(n5773_1), .A1(n5771), .B0(n5768_1), .Y(n5774));
AND2X1   g1135(.A(g3361), .B(g3396), .Y(n5775));
NAND4X1  g1136(.A(n5769), .B(n5772), .C(g84), .D(n5775), .Y(n5776));
NAND4X1  g1137(.A(n5770), .B(n5769), .C(n5495), .D(n5775), .Y(n5777));
NAND3X1  g1138(.A(n5777), .B(n5776), .C(n5774), .Y(n5778_1));
INVX1    g1139(.A(g3355), .Y(n5779));
OAI21X1  g1140(.A0(g3401), .A1(g3361), .B0(n5779), .Y(n5780));
INVX1    g1141(.A(g3361), .Y(n5781));
NAND3X1  g1142(.A(n5767), .B(n5781), .C(g3355), .Y(n5782));
OAI21X1  g1143(.A0(n5780), .A1(n5778_1), .B0(n5782), .Y(n5783_1));
MX2X1    g1144(.A(g3361), .B(n5783_1), .S0(g35), .Y(n865));
INVX1    g1145(.A(g2803), .Y(n5785));
AOI21X1  g1146(.A0(n5566), .A1(n5785), .B0(n5564_1), .Y(n5786));
OR2X1    g1147(.A(g2715), .B(g2719), .Y(n5787_1));
NOR2X1   g1148(.A(n5787_1), .B(n5786), .Y(n5788));
INVX1    g1149(.A(g2185), .Y(n5789));
NAND3X1  g1150(.A(n4937), .B(g2173), .C(n5789), .Y(n5790));
NAND3X1  g1151(.A(g2161), .B(n5789), .C(g2208), .Y(n5791));
AND2X1   g1152(.A(n5791), .B(n5790), .Y(n5792_1));
AND2X1   g1153(.A(g2217), .B(g2185), .Y(n5793));
NOR2X1   g1154(.A(n4937), .B(g2208), .Y(n5794));
AOI22X1  g1155(.A0(n5793), .A1(g2165), .B0(g2169), .B1(n5794), .Y(n5795));
NAND3X1  g1156(.A(g2181), .B(n4937), .C(g2208), .Y(n5796));
INVX1    g1157(.A(g2208), .Y(n5797_1));
NAND3X1  g1158(.A(g2185), .B(n5797_1), .C(g2177), .Y(n5798));
NAND4X1  g1159(.A(n5796), .B(n5795), .C(n5792_1), .D(n5798), .Y(n5799));
MX2X1    g1160(.A(g2236), .B(n5799), .S0(n5788), .Y(n5800));
MX2X1    g1161(.A(g2217), .B(n5800), .S0(g35), .Y(n870));
INVX1    g1162(.A(g3694), .Y(n5802_1));
INVX1    g1163(.A(g3618), .Y(n5803));
INVX1    g1164(.A(g3632), .Y(n5804));
INVX1    g1165(.A(g3689), .Y(n5805));
NAND2X1  g1166(.A(g3654), .B(g3661), .Y(n5806));
NOR4X1   g1167(.A(n5805), .B(n5804), .C(n5803), .D(n5806), .Y(n5807_1));
AOI21X1  g1168(.A0(n5807_1), .A1(g35), .B0(n5802_1), .Y(n880));
INVX1    g1169(.A(g6098), .Y(n5809));
NOR2X1   g1170(.A(g6093), .B(n5809), .Y(n5810));
INVX1    g1171(.A(g6088), .Y(n5811_1));
INVX1    g1172(.A(g6082), .Y(n5812));
NOR3X1   g1173(.A(n5812), .B(n5811_1), .C(g84), .Y(n5813));
INVX1    g1174(.A(g6077), .Y(n5814));
NOR3X1   g1175(.A(n5812), .B(n5814), .C(n5495), .Y(n5815));
OAI21X1  g1176(.A0(n5815), .A1(n5813), .B0(n5810), .Y(n5816_1));
AND2X1   g1177(.A(g6058), .B(g6093), .Y(n5817));
NAND4X1  g1178(.A(n5812), .B(n5814), .C(g84), .D(n5817), .Y(n5818));
NAND4X1  g1179(.A(n5812), .B(n5811_1), .C(n5495), .D(n5817), .Y(n5819));
NAND3X1  g1180(.A(n5819), .B(n5818), .C(n5816_1), .Y(n5820));
INVX1    g1181(.A(g6069), .Y(n5821_1));
INVX1    g1182(.A(g6065), .Y(n5822));
INVX1    g1183(.A(g6052), .Y(n5823));
NOR4X1   g1184(.A(n5809), .B(n5822), .C(n5821_1), .D(n5823), .Y(n5824));
INVX1    g1185(.A(n5824), .Y(n5825));
INVX1    g1186(.A(g6058), .Y(n5826_1));
NOR4X1   g1187(.A(g6052), .B(g6065), .C(g6069), .D(n5826_1), .Y(n5827));
INVX1    g1188(.A(n5827), .Y(n5828));
NAND3X1  g1189(.A(n5828), .B(n5825), .C(g6073), .Y(n5829));
INVX1    g1190(.A(g6073), .Y(n5830));
OAI21X1  g1191(.A0(n5827), .A1(n5824), .B0(n5830), .Y(n5831_1));
OAI21X1  g1192(.A0(n5829), .A1(n5820), .B0(n5831_1), .Y(n5832));
MX2X1    g1193(.A(g6069), .B(n5832), .S0(g35), .Y(n885));
INVX1    g1194(.A(g1728), .Y(n5834));
NOR3X1   g1195(.A(n5628), .B(g1772), .C(n5834), .Y(n5835));
MX2X1    g1196(.A(g1736), .B(n5624), .S0(n5835), .Y(n5836_1));
MX2X1    g1197(.A(g1740), .B(n5836_1), .S0(g35), .Y(n890));
INVX1    g1198(.A(g1894), .Y(n5838));
INVX1    g1199(.A(g2783), .Y(n5839));
AOI21X1  g1200(.A0(n5566), .A1(n5839), .B0(n5564_1), .Y(n5840));
NOR4X1   g1201(.A(n5569), .B(n5838), .C(n4939_1), .D(n5840), .Y(n5841_1));
XOR2X1   g1202(.A(n5841_1), .B(g1968), .Y(n5842));
MX2X1    g1203(.A(g1964), .B(n5842), .S0(g35), .Y(n895));
INVX1    g1204(.A(g4643), .Y(n5844));
OAI21X1  g1205(.A0(n5702), .A1(n5506), .B0(g65), .Y(n5845_1));
AND2X1   g1206(.A(n5845_1), .B(n5844), .Y(n5846));
INVX1    g1207(.A(n5846), .Y(n5847));
INVX1    g1208(.A(g4621), .Y(n5848));
NAND4X1  g1209(.A(g4639), .B(n5844), .C(n5848), .D(n5845_1), .Y(n5849));
INVX1    g1210(.A(g4639), .Y(n5850_1));
NAND2X1  g1211(.A(n5850_1), .B(g4621), .Y(n5851));
OAI21X1  g1212(.A0(n5851), .A1(n5847), .B0(n5849), .Y(n5852));
MX2X1    g1213(.A(g4639), .B(n5852), .S0(g35), .Y(n900));
INVX1    g1214(.A(g5511), .Y(n5854));
INVX1    g1215(.A(g5517), .Y(n5855_1));
NOR4X1   g1216(.A(n4868), .B(g5535), .C(n5854), .D(n5855_1), .Y(n5856));
MX2X1    g1217(.A(g5607), .B(n5592_1), .S0(n5856), .Y(n5857));
MX2X1    g1218(.A(g5591), .B(n5857), .S0(g35), .Y(n905));
XOR2X1   g1219(.A(g2648), .B(g2652), .Y(n5859));
INVX1    g1220(.A(g2610), .Y(n5860_1));
NOR4X1   g1221(.A(n5508), .B(g2741), .C(g2819), .D(n5565), .Y(n5861));
AND2X1   g1222(.A(g2715), .B(g2719), .Y(n5862));
OAI21X1  g1223(.A0(n5861), .A1(n5564_1), .B0(n5862), .Y(n5863));
NOR3X1   g1224(.A(n5863), .B(g2587), .C(n5860_1), .Y(n5864));
MX2X1    g1225(.A(g2657), .B(n5859), .S0(n5864), .Y(n5865_1));
MX2X1    g1226(.A(g2652), .B(n5865_1), .S0(g35), .Y(n910));
INVX1    g1227(.A(g5623), .Y(n5867));
INVX1    g1228(.A(g5637), .Y(n5868));
OAI22X1  g1229(.A0(n5867), .A1(g5666), .B0(g5659), .B1(n5868), .Y(n5869));
MX2X1    g1230(.A(g5654), .B(n5867), .S0(g5630), .Y(n5870_1));
INVX1    g1231(.A(g5659), .Y(n5871));
INVX1    g1232(.A(g5666), .Y(n5872));
NOR4X1   g1233(.A(n5867), .B(n5872), .C(n5871), .D(n5868), .Y(n5873));
OAI21X1  g1234(.A0(g5637), .A1(n5872), .B0(g35), .Y(n5874));
NOR4X1   g1235(.A(n5873), .B(n5870_1), .C(n5869), .D(n5874), .Y(n915));
INVX1    g1236(.A(g667), .Y(n5876));
OAI21X1  g1237(.A0(g686), .A1(n5876), .B0(g490), .Y(n5877));
NOR3X1   g1238(.A(n5130_1), .B(g528), .C(n5132), .Y(n5878));
INVX1    g1239(.A(n5878), .Y(n5879));
NOR3X1   g1240(.A(n5600), .B(g376), .C(n5598), .Y(n5880_1));
NOR2X1   g1241(.A(n5129), .B(g513), .Y(n5881));
NAND2X1  g1242(.A(n5881), .B(n5880_1), .Y(n5882));
AOI21X1  g1243(.A0(n5879), .A1(n5142), .B0(n5882), .Y(n5883));
NAND2X1  g1244(.A(n5883), .B(g482), .Y(n5884));
OAI21X1  g1245(.A0(g686), .A1(n5876), .B0(n5132), .Y(n5885_1));
MX2X1    g1246(.A(n5877), .B(n5885_1), .S0(n5884), .Y(n5886));
MX2X1    g1247(.A(g482), .B(n5886), .S0(g35), .Y(n920));
MX2X1    g1248(.A(g305), .B(g6744), .S0(g35), .Y(n925));
NOR3X1   g1249(.A(n5823), .B(n5809), .C(n5822), .Y(n5889));
NOR3X1   g1250(.A(n5826_1), .B(g6052), .C(g6065), .Y(n5890_1));
OAI21X1  g1251(.A0(n5890_1), .A1(n5889), .B0(n5821_1), .Y(n5891));
NOR2X1   g1252(.A(n5890_1), .B(n5889), .Y(n5892));
NAND2X1  g1253(.A(n5892), .B(g6069), .Y(n5893));
OAI21X1  g1254(.A0(n5893), .A1(n5820), .B0(n5891), .Y(n5894));
MX2X1    g1255(.A(g6065), .B(n5894), .S0(g35), .Y(n930));
NAND3X1  g1256(.A(n5677), .B(n5675), .C(n5673), .Y(n5896));
MX2X1    g1257(.A(n5294_1), .B(n5678), .S0(n5896), .Y(n5897));
MX2X1    g1258(.A(g767), .B(n5897), .S0(g35), .Y(n935));
OR2X1    g1259(.A(g5527), .B(g5535), .Y(n5899_1));
NOR3X1   g1260(.A(n5899_1), .B(n5855_1), .C(g5511), .Y(n5900));
MX2X1    g1261(.A(g5587), .B(n5592_1), .S0(n5900), .Y(n5901));
MX2X1    g1262(.A(g5571), .B(n5901), .S0(g35), .Y(n940));
INVX1    g1263(.A(g6167), .Y(n5903));
XOR2X1   g1264(.A(g6173), .B(n5903), .Y(n5904_1));
INVX1    g1265(.A(g4765), .Y(n5905));
NOR4X1   g1266(.A(n5905), .B(n4818), .C(n4815), .D(n4723), .Y(n5906));
AOI21X1  g1267(.A0(n5906), .A1(n4721), .B0(n4967), .Y(n5907));
INVX1    g1268(.A(n5907), .Y(n5908));
NAND4X1  g1269(.A(g6395), .B(g6322), .C(g6336), .D(g6381), .Y(n5909_1));
NOR2X1   g1270(.A(n5909_1), .B(n5908), .Y(n5910));
MX2X1    g1271(.A(g6177), .B(n5904_1), .S0(n5910), .Y(n5911));
MX2X1    g1272(.A(g6173), .B(n5911), .S0(g35), .Y(n945));
INVX1    g1273(.A(g3155), .Y(n5913));
NOR4X1   g1274(.A(n5593), .B(g3167), .C(n5913), .D(n5765), .Y(n5914_1));
MX2X1    g1275(.A(g3161), .B(n5914_1), .S0(g35), .Y(n955));
NAND2X1  g1276(.A(g5527), .B(g5535), .Y(n5916));
NOR3X1   g1277(.A(n5916), .B(n5855_1), .C(n5854), .Y(n5917));
MX2X1    g1278(.A(g5615), .B(n5592_1), .S0(n5917), .Y(n5918));
MX2X1    g1279(.A(g5599), .B(n5918), .S0(g35), .Y(n960));
INVX1    g1280(.A(g4575), .Y(n5920));
NAND3X1  g1281(.A(n5920), .B(g73), .C(n4950), .Y(n5921));
MX2X1    g1282(.A(g4543), .B(n5921), .S0(g4581), .Y(n5922));
MX2X1    g1283(.A(g4543), .B(n5922), .S0(g35), .Y(n965));
INVX1    g1284(.A(g3045), .Y(n5924_1));
NAND3X1  g1285(.A(n5583_1), .B(n5582), .C(g35), .Y(n5925));
OAI21X1  g1286(.A0(n5924_1), .A1(g35), .B0(n5925), .Y(n970));
INVX1    g1287(.A(g4871), .Y(n5927));
NOR3X1   g1288(.A(n4963), .B(g4991), .C(g4983), .Y(n5928));
NOR4X1   g1289(.A(g4975), .B(n4893), .C(n4892), .D(n4960), .Y(n5929_1));
AOI21X1  g1290(.A0(n5929_1), .A1(n5928), .B0(n5927), .Y(n5930));
INVX1    g1291(.A(g3639), .Y(n5931));
NAND2X1  g1292(.A(g3703), .B(n5931), .Y(n5932));
NAND3X1  g1293(.A(n5805), .B(g3625), .C(g3554), .Y(n5933));
NAND3X1  g1294(.A(g3654), .B(g3689), .C(g3542), .Y(n5934_1));
AOI21X1  g1295(.A0(n5934_1), .A1(n5933), .B0(n5932), .Y(n5935));
NAND4X1  g1296(.A(g3668), .B(n5805), .C(g3574), .D(n5176_1), .Y(n5936));
INVX1    g1297(.A(g3703), .Y(n5937));
NAND2X1  g1298(.A(n5937), .B(g3639), .Y(n5938));
NAND3X1  g1299(.A(g3550), .B(n5805), .C(g3649), .Y(n5939_1));
OAI21X1  g1300(.A0(n5939_1), .A1(n5938), .B0(n5936), .Y(n5940));
NOR2X1   g1301(.A(n5940), .B(n5935), .Y(n5941));
AND2X1   g1302(.A(g3668), .B(g3689), .Y(n5942));
NAND4X1  g1303(.A(g3703), .B(n5931), .C(g3566), .D(n5942), .Y(n5943));
NAND4X1  g1304(.A(g3676), .B(g3689), .C(g3598), .D(n5176_1), .Y(n5944_1));
NOR2X1   g1305(.A(g3703), .B(g3639), .Y(n5945));
NAND4X1  g1306(.A(g3538), .B(g3689), .C(g3649), .D(n5945), .Y(n5946));
AND2X1   g1307(.A(g3689), .B(g3672), .Y(n5947));
NAND4X1  g1308(.A(n5937), .B(g3582), .C(g3639), .D(n5947), .Y(n5948));
NAND4X1  g1309(.A(n5946), .B(n5944_1), .C(n5943), .D(n5948), .Y(n5949_1));
NAND4X1  g1310(.A(g3590), .B(n5805), .C(g3672), .D(n5945), .Y(n5950));
NAND3X1  g1311(.A(g3676), .B(n5805), .C(g3606), .Y(n5951));
OAI21X1  g1312(.A0(n5951), .A1(n5932), .B0(n5950), .Y(n5952));
NAND4X1  g1313(.A(g3546), .B(g3689), .C(g3680), .D(n5945), .Y(n5953));
NAND4X1  g1314(.A(g3614), .B(g3689), .C(g3625), .D(n5176_1), .Y(n5954_1));
NAND2X1  g1315(.A(n5954_1), .B(n5953), .Y(n5955));
NOR3X1   g1316(.A(n5955), .B(n5952), .C(n5949_1), .Y(n5956));
XOR2X1   g1317(.A(g3654), .B(n5805), .Y(n5957));
AND2X1   g1318(.A(g3661), .B(g3586), .Y(n5958_1));
AND2X1   g1319(.A(n5958_1), .B(n5176_1), .Y(n5959));
NAND3X1  g1320(.A(n5945), .B(g3578), .C(g3632), .Y(n5960));
NAND4X1  g1321(.A(g3594), .B(g3661), .C(n5931), .D(g3703), .Y(n5961));
AOI21X1  g1322(.A0(n5961), .A1(n5960), .B0(n5957), .Y(n5962_1));
AOI21X1  g1323(.A0(n5959), .A1(n5957), .B0(n5962_1), .Y(n5963));
NAND4X1  g1324(.A(g3610), .B(g3639), .C(g3618), .D(n5937), .Y(n5964));
NOR2X1   g1325(.A(n5964), .B(n5957), .Y(n5965));
NAND4X1  g1326(.A(g3654), .B(n5805), .C(g3558), .D(n5176_1), .Y(n5966));
NAND3X1  g1327(.A(g3562), .B(n5805), .C(g3680), .Y(n5967_1));
OAI21X1  g1328(.A0(n5967_1), .A1(n5938), .B0(n5966), .Y(n5968));
INVX1    g1329(.A(n5957), .Y(n5969));
NAND3X1  g1330(.A(n5945), .B(g3602), .C(g3618), .Y(n5970));
NAND4X1  g1331(.A(g3639), .B(g3632), .C(g3570), .D(n5937), .Y(n5971));
AOI21X1  g1332(.A0(n5971), .A1(n5970), .B0(n5969), .Y(n5972_1));
NOR3X1   g1333(.A(n5972_1), .B(n5968), .C(n5965), .Y(n5973));
NAND4X1  g1334(.A(n5963), .B(n5956), .C(n5941), .D(n5973), .Y(n5974));
NAND4X1  g1335(.A(g3689), .B(g3639), .C(g3625), .D(g3703), .Y(n5975));
AND2X1   g1336(.A(n5975), .B(g3457), .Y(n5976));
XOR2X1   g1337(.A(n5976), .B(n5974), .Y(n5977_1));
MX2X1    g1338(.A(g3457), .B(n5977_1), .S0(n5930), .Y(n5978));
MX2X1    g1339(.A(g3462), .B(n5978), .S0(g35), .Y(n975));
INVX1    g1340(.A(g6209), .Y(n5980));
NOR4X1   g1341(.A(n4873), .B(n5980), .C(g6219), .D(g6203), .Y(n5981));
MX2X1    g1342(.A(g6287), .B(n5592_1), .S0(n5981), .Y(n5982_1));
MX2X1    g1343(.A(g6271), .B(n5982_1), .S0(g35), .Y(n980));
XOR2X1   g1344(.A(g1322), .B(g1339), .Y(n5984));
NOR2X1   g1345(.A(g1322), .B(g1333), .Y(n5985));
INVX1    g1346(.A(n5985), .Y(n5986));
XOR2X1   g1347(.A(g1322), .B(g1579), .Y(n5987_1));
NAND4X1  g1348(.A(n5986), .B(n5984), .C(n4712_1), .D(n5987_1), .Y(n5988));
OR2X1    g1349(.A(g1582), .B(g1459), .Y(n5989));
OR4X1    g1350(.A(g1399), .B(g1333), .C(g1500), .D(n5989), .Y(n5990));
XOR2X1   g1351(.A(n5990), .B(n5988), .Y(n5991));
MX2X1    g1352(.A(g1339), .B(n5991), .S0(g35), .Y(n985));
OAI21X1  g1353(.A0(n5541_1), .A1(g134), .B0(n5244), .Y(n5993));
NOR2X1   g1354(.A(n5543), .B(n5447), .Y(n5994));
NOR2X1   g1355(.A(n5994), .B(n5993), .Y(n5995));
INVX1    g1356(.A(n5995), .Y(n5996_1));
AOI21X1  g1357(.A0(n5994), .A1(n5524), .B0(n5993), .Y(n5997));
OAI21X1  g1358(.A0(n5996_1), .A1(g1585), .B0(n5997), .Y(n5998));
INVX1    g1359(.A(g2555), .Y(n5999));
INVX1    g1360(.A(g1526), .Y(n6000_1));
NAND4X1  g1361(.A(g1322), .B(g1404), .C(n6000_1), .D(n5549), .Y(n6001));
OAI21X1  g1362(.A0(n6001), .A1(n5548), .B0(g1430), .Y(n6002));
AND2X1   g1363(.A(n6002), .B(n5995), .Y(n6003));
NOR3X1   g1364(.A(n6003), .B(n5999), .C(g2599), .Y(n6004));
MX2X1    g1365(.A(g2563), .B(n5998), .S0(n6004), .Y(n6005_1));
MX2X1    g1366(.A(g2567), .B(n6005_1), .S0(g35), .Y(n990));
NAND3X1  g1367(.A(n5506), .B(n4957), .C(g63), .Y(n6007));
NOR4X1   g1368(.A(n4967), .B(n4969_1), .C(n4720), .D(n4723), .Y(n6008));
INVX1    g1369(.A(n6008), .Y(n6009));
AND2X1   g1370(.A(n6009), .B(n6007), .Y(n6010_1));
INVX1    g1371(.A(g4801), .Y(n6011));
NOR4X1   g1372(.A(n4967), .B(n4969_1), .C(n6011), .D(n4723), .Y(n6012));
AND2X1   g1373(.A(n6012), .B(n4720), .Y(n6013));
NOR2X1   g1374(.A(n6012), .B(n4720), .Y(n6014));
OAI21X1  g1375(.A0(n6014), .A1(n6013), .B0(n6010_1), .Y(n6015_1));
NAND2X1  g1376(.A(g4801), .B(n4620), .Y(n6016));
OAI21X1  g1377(.A0(n6015_1), .A1(n4620), .B0(n6016), .Y(n995));
INVX1    g1378(.A(g4628), .Y(n6018));
NAND3X1  g1379(.A(g4358), .B(g4349), .C(g4340), .Y(n6019));
NOR4X1   g1380(.A(n6018), .B(g4639), .C(n5848), .D(n6019), .Y(n6020_1));
NAND3X1  g1381(.A(n6020_1), .B(g4322), .C(g4332), .Y(n6021));
NAND3X1  g1382(.A(n6020_1), .B(g4616), .C(g4584), .Y(n6022));
OAI21X1  g1383(.A0(n6022), .A1(n6021), .B0(n5845_1), .Y(n6023));
NAND4X1  g1384(.A(g4322), .B(g4584), .C(g4332), .D(n6020_1), .Y(n6024_1));
NAND2X1  g1385(.A(n6024_1), .B(g4593), .Y(n6025));
OR2X1    g1386(.A(n6024_1), .B(g4593), .Y(n6026));
AOI21X1  g1387(.A0(n6026), .A1(n6025), .B0(n6023), .Y(n6027));
MX2X1    g1388(.A(g4584), .B(n6027), .S0(g35), .Y(n1000));
NOR3X1   g1389(.A(n4988_1), .B(n5019), .C(n5616), .Y(n6029));
MX2X1    g1390(.A(g6199), .B(n3747), .S0(n6029), .Y(n6030));
AND2X1   g1391(.A(n6030), .B(g35), .Y(n1005));
INVX1    g1392(.A(g2287), .Y(n6032));
NOR3X1   g1393(.A(n5552), .B(g2331), .C(n6032), .Y(n6033_1));
MX2X1    g1394(.A(g2295), .B(n5547), .S0(n6033_1), .Y(n6034));
MX2X1    g1395(.A(g2299), .B(n6034), .S0(g35), .Y(n1010));
INVX1    g1396(.A(g1351), .Y(n6036));
NOR2X1   g1397(.A(n6036), .B(g1384), .Y(n6037));
OAI21X1  g1398(.A0(g1322), .A1(g1333), .B0(n5984), .Y(n6038_1));
MX2X1    g1399(.A(n6037), .B(g1384), .S0(n6038_1), .Y(n6039));
MX2X1    g1400(.A(g1379), .B(n6039), .S0(g35), .Y(n1015));
MX2X1    g1401(.A(g1579), .B(g1570), .S0(g35), .Y(n1020));
NOR3X1   g1402(.A(n5645_1), .B(n4837), .C(g4087), .Y(n6042));
NAND2X1  g1403(.A(g5176), .B(n4642_1), .Y(n6043_1));
NAND2X1  g1404(.A(n4644), .B(g5180), .Y(n6044));
AOI21X1  g1405(.A0(n6044), .A1(n6043_1), .B0(n6042), .Y(n6045));
MX2X1    g1406(.A(g5176), .B(n6045), .S0(g35), .Y(n1025));
MX2X1    g1407(.A(g2844), .B(n3747), .S0(n5697), .Y(n6047));
MX2X1    g1408(.A(g2890), .B(n6047), .S0(g35), .Y(n1030));
INVX1    g1409(.A(g1008), .Y(n6049));
XOR2X1   g1410(.A(g979), .B(g996), .Y(n6050));
AOI21X1  g1411(.A0(n6050), .A1(n6049), .B0(g969), .Y(n6051));
INVX1    g1412(.A(g1046), .Y(n6052));
NAND3X1  g1413(.A(g1008), .B(g1018), .C(g1030), .Y(n6053_1));
MX2X1    g1414(.A(n6053_1), .B(n6052), .S0(n6050), .Y(n6054));
NAND2X1  g1415(.A(n6054), .B(n6051), .Y(n6055));
NOR2X1   g1416(.A(n6055), .B(g1024), .Y(n6056));
NOR2X1   g1417(.A(n6055), .B(g1018), .Y(n6057));
NOR2X1   g1418(.A(g979), .B(g990), .Y(n6058_1));
INVX1    g1419(.A(n6058_1), .Y(n6059));
OAI21X1  g1420(.A0(n6055), .A1(g1002), .B0(n6059), .Y(n6060));
NOR2X1   g1421(.A(n6060), .B(n6057), .Y(n6061));
MX2X1    g1422(.A(g1024), .B(n6056), .S0(n6061), .Y(n6062));
MX2X1    g1423(.A(g1018), .B(n6062), .S0(g35), .Y(n1035));
NOR4X1   g1424(.A(n4868), .B(g5535), .C(g5511), .D(n5855_1), .Y(n6064));
MX2X1    g1425(.A(g5591), .B(n5592_1), .S0(n6064), .Y(n6065));
MX2X1    g1426(.A(g5575), .B(n6065), .S0(g35), .Y(n1040));
OR2X1    g1427(.A(g3522), .B(g3530), .Y(n6067));
NOR3X1   g1428(.A(n6067), .B(n5735), .C(n5733_1), .Y(n6068_1));
MX2X1    g1429(.A(g3598), .B(n5592_1), .S0(n6068_1), .Y(n6069));
MX2X1    g1430(.A(g3582), .B(n6069), .S0(g35), .Y(n1045));
XOR2X1   g1431(.A(g4258), .B(g4264), .Y(n6071));
MX2X1    g1432(.A(g4258), .B(n6071), .S0(g35), .Y(n1050));
AND2X1   g1433(.A(n5675), .B(n5673), .Y(n6073_1));
MX2X1    g1434(.A(n5677), .B(n5676), .S0(n6073_1), .Y(n6074));
MX2X1    g1435(.A(g763), .B(n6074), .S0(g35), .Y(n1055));
INVX1    g1436(.A(n5468), .Y(n6676));
MX2X1    g1437(.A(g5853), .B(n6676), .S0(n6029), .Y(n6077));
AND2X1   g1438(.A(n6077), .B(g35), .Y(n1060));
INVX1    g1439(.A(g1183), .Y(n6079));
NAND4X1  g1440(.A(g979), .B(n6079), .C(n4665), .D(g1061), .Y(n6080));
OAI21X1  g1441(.A0(n6080), .A1(n5528), .B0(g1087), .Y(n6081));
NAND2X1  g1442(.A(n5752), .B(n5246_1), .Y(n6082));
NOR2X1   g1443(.A(n5519), .B(n5269_1), .Y(n6083_1));
NOR2X1   g1444(.A(n6083_1), .B(n6082), .Y(n6084));
AND2X1   g1445(.A(n6084), .B(n6081), .Y(n6085));
NOR3X1   g1446(.A(n6085), .B(g1996), .C(g2070), .Y(n6086));
MX2X1    g1447(.A(g2089), .B(g2084), .S0(n6086), .Y(n6087_1));
MX2X1    g1448(.A(g2084), .B(n6087_1), .S0(g35), .Y(n1070));
NOR3X1   g1449(.A(n4809), .B(g5008), .C(g4999), .Y(n6089));
AOI21X1  g1450(.A0(n4964_1), .A1(n4890), .B0(n6089), .Y(n6090));
MX2X1    g1451(.A(g4939), .B(g71), .S0(n6089), .Y(n6091));
MX2X1    g1452(.A(n6091), .B(g4933), .S0(n6090), .Y(n6092_1));
MX2X1    g1453(.A(g4939), .B(n6092_1), .S0(g35), .Y(n1075));
NAND2X1  g1454(.A(g4581), .B(g4531), .Y(n6094));
MX2X1    g1455(.A(g4512), .B(n6094), .S0(g35), .Y(n1080));
INVX1    g1456(.A(n5465), .Y(n4447));
MX2X1    g1457(.A(g5507), .B(n4447), .S0(n6029), .Y(n6097));
AND2X1   g1458(.A(n6097), .B(g35), .Y(n1085));
NAND2X1  g1459(.A(g6227), .B(g6219), .Y(n6099));
NOR3X1   g1460(.A(n6099), .B(g6203), .C(n5980), .Y(n6100_1));
MX2X1    g1461(.A(g6291), .B(n5592_1), .S0(n6100_1), .Y(n6101));
MX2X1    g1462(.A(g6275), .B(n6101), .S0(g35), .Y(n1094));
INVX1    g1463(.A(g294), .Y(n6103));
INVX1    g1464(.A(g283), .Y(n6104));
INVX1    g1465(.A(g225), .Y(n6105_1));
INVX1    g1466(.A(g232), .Y(n6106));
INVX1    g1467(.A(g269), .Y(n6107));
INVX1    g1468(.A(g262), .Y(n6108));
NOR4X1   g1469(.A(n6107), .B(g239), .C(g246), .D(n6108), .Y(n6109));
NAND4X1  g1470(.A(g255), .B(n6106), .C(n6105_1), .D(n6109), .Y(n6110_1));
NAND4X1  g1471(.A(n6107), .B(g239), .C(g246), .D(n6108), .Y(n6111));
OR4X1    g1472(.A(g255), .B(n6106), .C(n6105_1), .D(n6111), .Y(n6112));
MX2X1    g1473(.A(n6110_1), .B(n6112), .S0(g278), .Y(n6113));
OR4X1    g1474(.A(n5661), .B(n5516_1), .C(n6104), .D(n6113), .Y(n6114_1));
INVX1    g1475(.A(g287), .Y(n6115));
OR4X1    g1476(.A(n5661), .B(n5516_1), .C(n6115), .D(n6113), .Y(n6116));
NOR2X1   g1477(.A(n6116), .B(n6114_1), .Y(n6117));
INVX1    g1478(.A(g291), .Y(n6118_1));
NOR4X1   g1479(.A(n5661), .B(n5516_1), .C(n6118_1), .D(n6113), .Y(n6119));
AND2X1   g1480(.A(n6119), .B(n6117), .Y(n6120));
NOR4X1   g1481(.A(n5661), .B(n5516_1), .C(n6103), .D(n6113), .Y(n6121));
MX2X1    g1482(.A(n6121), .B(n6103), .S0(n6120), .Y(n6122));
MX2X1    g1483(.A(g291), .B(n6122), .S0(g35), .Y(n1099));
NOR3X1   g1484(.A(n4868), .B(g5535), .C(n4866_1), .Y(n6124));
MX2X1    g1485(.A(g5559), .B(n5592_1), .S0(n6124), .Y(n6125));
MX2X1    g1486(.A(g5607), .B(n6125), .S0(g35), .Y(n1104));
AND2X1   g1487(.A(g5881), .B(g35), .Y(n1109));
MX2X1    g1488(.A(g6098), .B(g6381), .S0(g35), .Y(n1114));
MX2X1    g1489(.A(g3813), .B(g3849), .S0(n4851_1), .Y(n6129));
MX2X1    g1490(.A(g3849), .B(n6129), .S0(g35), .Y(n1119));
INVX1    g1491(.A(g637), .Y(n6131));
OAI21X1  g1492(.A0(n6131), .A1(g640), .B0(g74), .Y(n6132_1));
INVX1    g1493(.A(g559), .Y(n6133));
AND2X1   g1494(.A(g640), .B(n6133), .Y(n6134));
AND2X1   g1495(.A(g626), .B(g632), .Y(n6135));
NOR3X1   g1496(.A(n6135), .B(n6134), .C(n5262), .Y(n6136_1));
NOR3X1   g1497(.A(n6135), .B(n6134), .C(g562), .Y(n6137));
MX2X1    g1498(.A(n6137), .B(n6136_1), .S0(n6132_1), .Y(n6138));
MX2X1    g1499(.A(g559), .B(n6138), .S0(g35), .Y(n1124));
NOR4X1   g1500(.A(n6132_1), .B(n5440_1), .C(n5262), .D(n6134), .Y(n6140));
AOI21X1  g1501(.A0(g640), .A1(n6133), .B0(n5410_1), .Y(n6141_1));
AOI21X1  g1502(.A0(g640), .A1(n6133), .B0(n5385_1), .Y(n6142));
NAND3X1  g1503(.A(n6142), .B(n6141_1), .C(n6140), .Y(n6143));
OR4X1    g1504(.A(n6134), .B(n5322_1), .C(n5349), .D(n6143), .Y(n6144));
OR4X1    g1505(.A(n6134), .B(n5228), .C(n5296), .D(n6144), .Y(n6145));
OR4X1    g1506(.A(n6134), .B(n5436), .C(n5258), .D(n6145), .Y(n6146_1));
AOI21X1  g1507(.A0(g640), .A1(n6133), .B0(n5406), .Y(n6147));
MX2X1    g1508(.A(n5406), .B(n6147), .S0(n6146_1), .Y(n6148));
MX2X1    g1509(.A(g604), .B(n6148), .S0(g35), .Y(n1129));
XOR2X1   g1510(.A(g1087), .B(g1205), .Y(n6150));
MX2X1    g1511(.A(g1087), .B(n6150), .S0(g35), .Y(n1134));
NOR3X1   g1512(.A(g3857), .B(g3863), .C(g3869), .Y(n6152));
NAND3X1  g1513(.A(n6152), .B(g3881), .C(g3873), .Y(n6153));
MX2X1    g1514(.A(n5592_1), .B(g3909), .S0(n6153), .Y(n6154));
MX2X1    g1515(.A(g3913), .B(n6154), .S0(g35), .Y(n1139));
NOR3X1   g1516(.A(n4873), .B(n4872), .C(g6219), .Y(n6156_1));
MX2X1    g1517(.A(g6259), .B(n5592_1), .S0(n6156_1), .Y(n6157));
MX2X1    g1518(.A(g6303), .B(n6157), .S0(g35), .Y(n1144));
NOR3X1   g1519(.A(g5881), .B(n4861_1), .C(n4860), .Y(n6159));
MX2X1    g1520(.A(g5905), .B(n5592_1), .S0(n6159), .Y(n6160));
MX2X1    g1521(.A(g5953), .B(n6160), .S0(g35), .Y(n1149));
INVX1    g1522(.A(g921), .Y(n6162));
AND2X1   g1523(.A(g904), .B(g1227), .Y(n6163));
AND2X1   g1524(.A(g1227), .B(g921), .Y(n6164));
MX2X1    g1525(.A(n6164), .B(n6162), .S0(n6163), .Y(n6165));
MX2X1    g1526(.A(g904), .B(n6165), .S0(g35), .Y(n1154));
NOR3X1   g1527(.A(n5462), .B(n5286), .C(n5616), .Y(n6167));
OAI21X1  g1528(.A0(n4647_1), .A1(n4646), .B0(g35), .Y(n6168));
INVX1    g1529(.A(n6168), .Y(n6169));
NOR2X1   g1530(.A(n4654), .B(n4651), .Y(n6170_1));
INVX1    g1531(.A(n6170_1), .Y(n6171));
OR4X1    g1532(.A(n6169), .B(g2946), .C(g2955), .D(n6171), .Y(n6172));
NAND2X1  g1533(.A(n4745), .B(n4697_1), .Y(n6173));
OAI21X1  g1534(.A0(n6173), .A1(n6172), .B0(g35), .Y(n6174_1));
NAND2X1  g1535(.A(g2941), .B(n4620), .Y(n6175));
OAI21X1  g1536(.A0(n6174_1), .A1(n6167), .B0(n6175), .Y(n1159));
INVX1    g1537(.A(g365), .Y(n6177));
NOR3X1   g1538(.A(n5600), .B(n5599), .C(n6177), .Y(n6178_1));
MX2X1    g1539(.A(g385), .B(n6178_1), .S0(g35), .Y(n1164));
NAND3X1  g1540(.A(n5824), .B(g6077), .C(g6073), .Y(n6180));
NOR2X1   g1541(.A(n6180), .B(n5812), .Y(n6181));
NAND3X1  g1542(.A(n5827), .B(n5814), .C(n5830), .Y(n6182));
NOR2X1   g1543(.A(n6182), .B(g6082), .Y(n6183_1));
OAI21X1  g1544(.A0(n6183_1), .A1(n6181), .B0(n5811_1), .Y(n6184));
OR4X1    g1545(.A(n6181), .B(n5820), .C(n5811_1), .D(n6183_1), .Y(n6185));
NAND2X1  g1546(.A(n6185), .B(n6184), .Y(n6186));
MX2X1    g1547(.A(g6082), .B(n6186), .S0(g35), .Y(n1169));
INVX1    g1548(.A(g1116), .Y(n6188));
NOR3X1   g1549(.A(n6188), .B(g1183), .C(g1171), .Y(n6189));
MX2X1    g1550(.A(g1099), .B(g1152), .S0(n6189), .Y(n6190));
MX2X1    g1551(.A(g1152), .B(n6190), .S0(g35), .Y(n1174));
NAND3X1  g1552(.A(n5506), .B(n4956), .C(g63), .Y(n6192));
INVX1    g1553(.A(n6192), .Y(n6193));
AOI21X1  g1554(.A0(n6193), .A1(g35), .B0(n5927), .Y(n1179));
OR2X1    g1555(.A(g5188), .B(g5180), .Y(n6195));
NOR2X1   g1556(.A(n6195), .B(n4644), .Y(n6196_1));
MX2X1    g1557(.A(g5204), .B(n5592_1), .S0(n6196_1), .Y(n6197));
MX2X1    g1558(.A(g5256), .B(n6197), .S0(g35), .Y(n1184));
NOR4X1   g1559(.A(n4833), .B(n5735), .C(n5733_1), .D(g3522), .Y(n6199));
MX2X1    g1560(.A(g3606), .B(n5592_1), .S0(n6199), .Y(n6200));
MX2X1    g1561(.A(g3590), .B(n6200), .S0(g35), .Y(n1194));
NOR2X1   g1562(.A(n5840), .B(n5569), .Y(n6202));
INVX1    g1563(.A(g1917), .Y(n6203));
NAND3X1  g1564(.A(n5637), .B(g110), .C(n4824), .Y(n6204));
OAI21X1  g1565(.A0(n6204), .A1(n4924), .B0(n6203), .Y(n6205));
MX2X1    g1566(.A(g1926), .B(n6205), .S0(n6202), .Y(n6206_1));
MX2X1    g1567(.A(g1932), .B(n6206_1), .S0(g35), .Y(n1199));
INVX1    g1568(.A(g6203), .Y(n6208));
NOR4X1   g1569(.A(n6208), .B(n5980), .C(g6215), .D(n5646), .Y(n6209));
MX2X1    g1570(.A(g6209), .B(n6209), .S0(g35), .Y(n1204));
NOR4X1   g1571(.A(g3530), .B(g3506), .C(n5733_1), .D(n4835), .Y(n6211_1));
MX2X1    g1572(.A(g3586), .B(n5592_1), .S0(n6211_1), .Y(n6212));
MX2X1    g1573(.A(g3570), .B(n6212), .S0(g35), .Y(n1209));
MX2X1    g1574(.A(n6119), .B(n6118_1), .S0(n6117), .Y(n6214));
MX2X1    g1575(.A(g287), .B(n6214), .S0(g35), .Y(n1214));
INVX1    g1576(.A(n6007), .Y(n6216_1));
AOI21X1  g1577(.A0(n6216_1), .A1(g35), .B0(n4719), .Y(n1219));
NOR4X1   g1578(.A(g3530), .B(n5735), .C(g3512), .D(n4835), .Y(n6218));
MX2X1    g1579(.A(g3570), .B(n5592_1), .S0(n6218), .Y(n6219));
MX2X1    g1580(.A(g3542), .B(n6219), .S0(g35), .Y(n1224));
NAND3X1  g1581(.A(n5530), .B(n5521_1), .C(g1862), .Y(n6221_1));
INVX1    g1582(.A(n5531_1), .Y(n6222));
NAND4X1  g1583(.A(n5637), .B(g112), .C(n4824), .D(n5146), .Y(n6223));
AOI21X1  g1584(.A0(g1906), .A1(n5527), .B0(g1936), .Y(n6224));
NAND3X1  g1585(.A(n6224), .B(n6223), .C(n6222), .Y(n6225));
AOI21X1  g1586(.A0(n6225), .A1(n6221_1), .B0(n4620), .Y(n1238));
XOR2X1   g1587(.A(g728), .B(g661), .Y(n6227));
XOR2X1   g1588(.A(g655), .B(g718), .Y(n6228));
INVX1    g1589(.A(g699), .Y(n6229));
OR2X1    g1590(.A(n6229), .B(g645), .Y(n6230));
INVX1    g1591(.A(g681), .Y(n6231_1));
OR2X1    g1592(.A(g650), .B(n6231_1), .Y(n6232));
NOR4X1   g1593(.A(n6230), .B(n6228), .C(n6227), .D(n6232), .Y(n6233));
INVX1    g1594(.A(g499), .Y(n6234));
INVX1    g1595(.A(n5688), .Y(n6235));
NOR4X1   g1596(.A(n6235), .B(n6234), .C(g504), .D(n5879), .Y(n6236_1));
NAND2X1  g1597(.A(n6236_1), .B(n6233), .Y(n6237));
NAND2X1  g1598(.A(n6237), .B(g703), .Y(n6238));
NAND2X1  g1599(.A(n6236_1), .B(g671), .Y(n6239));
NAND2X1  g1600(.A(n6239), .B(g676), .Y(n6240));
INVX1    g1601(.A(g676), .Y(n6241_1));
NAND3X1  g1602(.A(n6236_1), .B(g671), .C(n6241_1), .Y(n6242));
AOI21X1  g1603(.A0(n6242), .A1(n6240), .B0(n6238), .Y(n6243));
MX2X1    g1604(.A(g671), .B(n6243), .S0(g35), .Y(n1243));
AND2X1   g1605(.A(g376), .B(g358), .Y(n6245));
NAND4X1  g1606(.A(g385), .B(g370), .C(g847), .D(n6245), .Y(n6246_1));
INVX1    g1607(.A(g837), .Y(n6247));
NOR2X1   g1608(.A(n6247), .B(g843), .Y(n6248));
AND2X1   g1609(.A(g837), .B(g843), .Y(n6249));
MX2X1    g1610(.A(n6248), .B(n6249), .S0(n6246_1), .Y(n6250));
MX2X1    g1611(.A(g837), .B(n6250), .S0(g35), .Y(n1248));
NOR3X1   g1612(.A(g4141), .B(g4082), .C(g4076), .Y(n6252));
NAND4X1  g1613(.A(n4726), .B(n4731_1), .C(g4064), .D(n6252), .Y(n6253));
MX2X1    g1614(.A(g4164), .B(g4132), .S0(n6253), .Y(n6254));
MX2X1    g1615(.A(g4129), .B(n6254), .S0(g35), .Y(n1253));
AND2X1   g1616(.A(n6021), .B(n5845_1), .Y(n6256_1));
NAND3X1  g1617(.A(n6020_1), .B(g4311), .C(g4322), .Y(n6257));
AND2X1   g1618(.A(n6257), .B(g4332), .Y(n6258));
NOR2X1   g1619(.A(n6257), .B(g4332), .Y(n6259));
OAI21X1  g1620(.A0(n6259), .A1(n6258), .B0(n6256_1), .Y(n6260));
NAND2X1  g1621(.A(g4322), .B(n4620), .Y(n6261_1));
OAI21X1  g1622(.A0(n6260), .A1(n4620), .B0(n6261_1), .Y(n1258));
INVX1    g1623(.A(g116), .Y(n6263));
MX2X1    g1624(.A(n6263), .B(g115), .S0(n5275), .Y(n6264));
MX2X1    g1625(.A(g114), .B(g116), .S0(g4157), .Y(n6265));
OR2X1    g1626(.A(n6265), .B(n6264), .Y(n6266_1));
MX2X1    g1627(.A(g120), .B(g124), .S0(g4146), .Y(n6267));
INVX1    g1628(.A(n6267), .Y(n6268));
INVX1    g1629(.A(g126), .Y(n6269));
MX2X1    g1630(.A(n6269), .B(g124), .S0(g4146), .Y(n6270));
OR2X1    g1631(.A(n6270), .B(n6268), .Y(n6271_1));
AOI22X1  g1632(.A0(n6268), .A1(n6270), .B0(n6265), .B1(n6264), .Y(n6272));
NAND3X1  g1633(.A(n6272), .B(n6271_1), .C(n6266_1), .Y(n6273));
MX2X1    g1634(.A(g4122), .B(n6273), .S0(g35), .Y(n1263));
NOR4X1   g1635(.A(n4955), .B(n4952), .C(g4311), .D(n5185), .Y(n6275));
NAND4X1  g1636(.A(n5506), .B(n6275), .C(g93), .D(n5907), .Y(n6276_1));
INVX1    g1637(.A(g6395), .Y(n6277));
NOR3X1   g1638(.A(n5908), .B(n6277), .C(g6336), .Y(n6278));
INVX1    g1639(.A(g6336), .Y(n6279));
AOI21X1  g1640(.A0(n5907), .A1(g6395), .B0(n6279), .Y(n6280));
OAI21X1  g1641(.A0(n6280), .A1(n6278), .B0(n6276_1), .Y(n6281_1));
NAND2X1  g1642(.A(g6395), .B(n4620), .Y(n6282));
OAI21X1  g1643(.A0(n6281_1), .A1(n4620), .B0(n6282), .Y(n1273));
NOR4X1   g1644(.A(n6134), .B(n5381), .C(n5406), .D(n6146_1), .Y(n6284));
AOI21X1  g1645(.A0(g640), .A1(n6133), .B0(n5345_1), .Y(n6285));
AND2X1   g1646(.A(n6285), .B(n6284), .Y(n6286_1));
AOI21X1  g1647(.A0(g640), .A1(n6133), .B0(n5318_1), .Y(n6287));
MX2X1    g1648(.A(n6287), .B(n5318_1), .S0(n6286_1), .Y(n6288));
MX2X1    g1649(.A(g617), .B(n6288), .S0(g35), .Y(n1278));
NOR4X1   g1650(.A(g3518), .B(g3506), .C(n4620), .D(n5732), .Y(n1283));
MX2X1    g1651(.A(g4555), .B(g6748), .S0(g35), .Y(n1288));
MX2X1    g1652(.A(g6058), .B(g6098), .S0(g6052), .Y(n6292));
OR2X1    g1653(.A(n6292), .B(n5822), .Y(n6293));
NAND2X1  g1654(.A(n6292), .B(n5822), .Y(n6294));
OAI21X1  g1655(.A0(n6293), .A1(n5820), .B0(n6294), .Y(n6295));
MX2X1    g1656(.A(g6052), .B(n6295), .S0(g35), .Y(n1293));
MX2X1    g1657(.A(g3111), .B(g3147), .S0(n4846_1), .Y(n6297));
MX2X1    g1658(.A(g3147), .B(n6297), .S0(g35), .Y(n1303));
NAND2X1  g1659(.A(g2638), .B(g2715), .Y(n6299));
NAND2X1  g1660(.A(n6299), .B(g2719), .Y(n6300));
AOI21X1  g1661(.A0(g2504), .A1(n5568_1), .B0(n6300), .Y(n6301_1));
NAND2X1  g1662(.A(n5568_1), .B(g2236), .Y(n6302));
AOI21X1  g1663(.A0(g2715), .A1(g2370), .B0(g2719), .Y(n6303));
AND2X1   g1664(.A(n6303), .B(n6302), .Y(n6304));
NOR4X1   g1665(.A(n5564_1), .B(g2735), .C(g2741), .D(n5565), .Y(n6305));
OR2X1    g1666(.A(n6305), .B(n6304), .Y(n6306_1));
INVX1    g1667(.A(g2719), .Y(n6307));
OAI21X1  g1668(.A0(n5568_1), .A1(g2807), .B0(n6307), .Y(n6308));
AOI21X1  g1669(.A0(n5785), .A1(n5568_1), .B0(n6308), .Y(n6309));
NOR2X1   g1670(.A(g2715), .B(g2815), .Y(n6310));
OAI21X1  g1671(.A0(n5568_1), .A1(g2819), .B0(g2719), .Y(n6311_1));
OAI21X1  g1672(.A0(n6311_1), .A1(n6310), .B0(n6305), .Y(n6312));
OAI22X1  g1673(.A0(n6309), .A1(n6312), .B0(n6306_1), .B1(n6301_1), .Y(n6313));
MX2X1    g1674(.A(g2834), .B(n6313), .S0(g35), .Y(n1308));
AND2X1   g1675(.A(g125), .B(g35), .Y(n1313));
OR2X1    g1676(.A(n5024), .B(n5004), .Y(n6316_1));
OAI21X1  g1677(.A0(n5457), .A1(n5435_1), .B0(g12), .Y(n6317));
NOR2X1   g1678(.A(n6317), .B(n6316_1), .Y(n6318));
OAI21X1  g1679(.A0(g933), .A1(g939), .B0(g35), .Y(n6319));
NAND2X1  g1680(.A(g952), .B(n4620), .Y(n6320));
OAI21X1  g1681(.A0(n6319), .A1(n6318), .B0(n6320), .Y(n1318));
INVX1    g1682(.A(g278), .Y(n6322));
NAND2X1  g1683(.A(n6112), .B(g35), .Y(n6323));
AOI21X1  g1684(.A0(n6110_1), .A1(n6322), .B0(n6323), .Y(n1323));
MX2X1    g1685(.A(g4489), .B(g6750), .S0(g35), .Y(n1328));
INVX1    g1686(.A(g4836), .Y(n6326_1));
AOI21X1  g1687(.A0(n6193), .A1(g35), .B0(n6326_1), .Y(n1333));
NOR2X1   g1688(.A(n6055), .B(g1030), .Y(n6328));
NOR4X1   g1689(.A(n6060), .B(n6057), .C(n6056), .D(n6328), .Y(n6329));
NOR2X1   g1690(.A(n6055), .B(g1036), .Y(n6330));
MX2X1    g1691(.A(g1036), .B(n6330), .S0(n6329), .Y(n6331_1));
MX2X1    g1692(.A(g1030), .B(n6331_1), .S0(g35), .Y(n1338));
INVX1    g1693(.A(g5297), .Y(n6333));
NAND2X1  g1694(.A(g5357), .B(n6333), .Y(n6334));
INVX1    g1695(.A(g5343), .Y(n6335));
NAND3X1  g1696(.A(g5212), .B(g5283), .C(n6335), .Y(n6336_1));
NAND3X1  g1697(.A(g5200), .B(g5313), .C(g5343), .Y(n6337));
AOI21X1  g1698(.A0(n6337), .A1(n6336_1), .B0(n6334), .Y(n6338));
NAND4X1  g1699(.A(g5327), .B(n6335), .C(g5232), .D(g25114), .Y(n6339));
INVX1    g1700(.A(g5357), .Y(n6340));
NAND2X1  g1701(.A(n6340), .B(g5297), .Y(n6341_1));
NAND3X1  g1702(.A(g5308), .B(g5208), .C(n6335), .Y(n6342));
OAI21X1  g1703(.A0(n6342), .A1(n6341_1), .B0(n6339), .Y(n6343));
NOR2X1   g1704(.A(n6343), .B(n6338), .Y(n6344));
AND2X1   g1705(.A(g5327), .B(g5343), .Y(n6345));
NAND4X1  g1706(.A(g5224), .B(g5357), .C(n6333), .D(n6345), .Y(n6346_1));
NAND4X1  g1707(.A(g5256), .B(g5335), .C(g5343), .D(g25114), .Y(n6347));
NOR2X1   g1708(.A(g5357), .B(g5297), .Y(n6348));
NAND4X1  g1709(.A(g5196), .B(g5308), .C(g5343), .D(n6348), .Y(n6349));
AND2X1   g1710(.A(g5331), .B(g5343), .Y(n6350));
NAND4X1  g1711(.A(n6340), .B(g5240), .C(g5297), .D(n6350), .Y(n6351_1));
NAND4X1  g1712(.A(n6349), .B(n6347), .C(n6346_1), .D(n6351_1), .Y(n6352));
NAND4X1  g1713(.A(g5248), .B(g5331), .C(n6335), .D(n6348), .Y(n6353));
NAND3X1  g1714(.A(g5335), .B(g5264), .C(n6335), .Y(n6354));
OAI21X1  g1715(.A0(n6354), .A1(n6334), .B0(n6353), .Y(n6355_1));
NAND4X1  g1716(.A(g5339), .B(g5343), .C(g5204), .D(n6348), .Y(n6356));
NAND4X1  g1717(.A(g5272), .B(g5283), .C(g5343), .D(g25114), .Y(n6357));
NAND2X1  g1718(.A(n6357), .B(n6356), .Y(n6358));
NOR3X1   g1719(.A(n6358), .B(n6355_1), .C(n6352), .Y(n6359));
XOR2X1   g1720(.A(g5313), .B(n6335), .Y(n6360_1));
AND2X1   g1721(.A(g5244), .B(g5320), .Y(n6361));
AND2X1   g1722(.A(n6361), .B(g25114), .Y(n6362));
NAND3X1  g1723(.A(n6348), .B(g5236), .C(g5290), .Y(n6363));
NAND4X1  g1724(.A(g5320), .B(g5357), .C(n6333), .D(g5252), .Y(n6364));
AOI21X1  g1725(.A0(n6364), .A1(n6363), .B0(n6360_1), .Y(n6365_1));
AOI21X1  g1726(.A0(n6362), .A1(n6360_1), .B0(n6365_1), .Y(n6366));
NAND4X1  g1727(.A(n6340), .B(g5268), .C(g5297), .D(g5276), .Y(n6367));
NOR2X1   g1728(.A(n6367), .B(n6360_1), .Y(n6368));
NAND4X1  g1729(.A(g5216), .B(g5313), .C(n6335), .D(g25114), .Y(n6369_1));
NAND3X1  g1730(.A(g5220), .B(g5339), .C(n6335), .Y(n6370));
OAI21X1  g1731(.A0(n6370), .A1(n6341_1), .B0(n6369_1), .Y(n6371));
INVX1    g1732(.A(n6360_1), .Y(n6372));
NAND3X1  g1733(.A(n6348), .B(g5260), .C(g5276), .Y(n6373));
NAND4X1  g1734(.A(n6340), .B(g5290), .C(g5297), .D(g5228), .Y(n6374_1));
AOI21X1  g1735(.A0(n6374_1), .A1(n6373), .B0(n6372), .Y(n6375));
NOR3X1   g1736(.A(n6375), .B(n6371), .C(n6368), .Y(n6376));
NAND4X1  g1737(.A(n6366), .B(n6359), .C(n6344), .D(n6376), .Y(n6377));
MX2X1    g1738(.A(g128), .B(n6377), .S0(g28753), .Y(n6378));
MX2X1    g1739(.A(g5272), .B(n6378), .S0(g35), .Y(n1343));
MX2X1    g1740(.A(g1178), .B(g996), .S0(g1157), .Y(n6380));
MX2X1    g1741(.A(g1183), .B(n6380), .S0(g35), .Y(n1348));
NOR4X1   g1742(.A(g3171), .B(n4844), .C(g3155), .D(n5593), .Y(n6382));
MX2X1    g1743(.A(g3239), .B(n5592_1), .S0(n6382), .Y(n6383));
MX2X1    g1744(.A(g3223), .B(n6383), .S0(g35), .Y(n1353));
INVX1    g1745(.A(g417), .Y(n6385));
NOR3X1   g1746(.A(g411), .B(g424), .C(n6385), .Y(n6386));
OR2X1    g1747(.A(n6386), .B(g691), .Y(n6387));
OAI21X1  g1748(.A0(g499), .A1(g518), .B0(g691), .Y(n6388));
NAND3X1  g1749(.A(n6388), .B(n6387), .C(n5601), .Y(n6389_1));
MX2X1    g1750(.A(g655), .B(g718), .S0(n6389_1), .Y(n6390));
MX2X1    g1751(.A(g655), .B(n6390), .S0(g35), .Y(n1358));
INVX1    g1752(.A(g6195), .Y(n6392));
OAI22X1  g1753(.A0(n5524), .A1(g4284), .B0(n6392), .B1(n4874), .Y(n6393));
OR4X1    g1754(.A(n5524), .B(g4284), .C(n6392), .D(n4874), .Y(n6394_1));
AOI21X1  g1755(.A0(n6394_1), .A1(n6393), .B0(n4620), .Y(n1363));
INVX1    g1756(.A(g1152), .Y(n6396));
NAND2X1  g1757(.A(n6396), .B(g1099), .Y(n6397));
NOR4X1   g1758(.A(n6188), .B(g1183), .C(n4665), .D(n6397), .Y(n6398));
XOR2X1   g1759(.A(g1094), .B(g1135), .Y(n6399_1));
MX2X1    g1760(.A(g1135), .B(n6399_1), .S0(n6398), .Y(n6400));
MX2X1    g1761(.A(g1094), .B(n6400), .S0(g35), .Y(n1368));
AND2X1   g1762(.A(g6120), .B(g6128), .Y(n6402));
AND2X1   g1763(.A(n6402), .B(g6133), .Y(n6403));
XOR2X1   g1764(.A(n6403), .B(g6137), .Y(n6404_1));
MX2X1    g1765(.A(g6133), .B(n6404_1), .S0(g35), .Y(n1373));
NAND3X1  g1766(.A(n6276_1), .B(n5907), .C(n6277), .Y(n6406));
OAI21X1  g1767(.A0(n5907), .A1(n6277), .B0(n6406), .Y(n6407));
MX2X1    g1768(.A(g6390), .B(n6407), .S0(g35), .Y(n1378));
INVX1    g1769(.A(g3376), .Y(n6409_1));
INVX1    g1770(.A(g3372), .Y(n6410));
INVX1    g1771(.A(g3368), .Y(n6411));
NOR4X1   g1772(.A(n6411), .B(n6410), .C(n5779), .D(n5767), .Y(n6412));
INVX1    g1773(.A(n6412), .Y(n6413));
NOR4X1   g1774(.A(g3368), .B(g3372), .C(g3355), .D(n5781), .Y(n6414_1));
INVX1    g1775(.A(n6414_1), .Y(n6415));
MX2X1    g1776(.A(n6413), .B(n6415), .S0(n6409_1), .Y(n6416));
OR2X1    g1777(.A(n6416), .B(g3380), .Y(n6417));
NAND2X1  g1778(.A(n6416), .B(g3380), .Y(n6418));
OAI21X1  g1779(.A0(n6418), .A1(n5778_1), .B0(n6417), .Y(n6419_1));
MX2X1    g1780(.A(g3376), .B(n6419_1), .S0(g35), .Y(n1383));
NAND4X1  g1781(.A(g5276), .B(g5290), .C(g5313), .D(g5320), .Y(n6421));
XOR2X1   g1782(.A(n6421), .B(n6335), .Y(n6422));
MX2X1    g1783(.A(g5339), .B(n6422), .S0(g35), .Y(n1388));
NAND3X1  g1784(.A(n5684_1), .B(n5682), .C(n5681), .Y(n6424_1));
AOI21X1  g1785(.A0(g802), .A1(n5662), .B0(n5320), .Y(n6425));
MX2X1    g1786(.A(n5320), .B(n6425), .S0(n6424_1), .Y(n6426));
MX2X1    g1787(.A(g807), .B(n6426), .S0(g35), .Y(n1393));
AOI21X1  g1788(.A0(g262), .A1(g72), .B0(g73), .Y(n6428));
OAI21X1  g1789(.A0(n6107), .A1(g72), .B0(n6428), .Y(n6429_1));
INVX1    g1790(.A(g255), .Y(n6430));
OAI21X1  g1791(.A0(n6430), .A1(g72), .B0(g73), .Y(n6431));
NAND3X1  g1792(.A(n6431), .B(n6429_1), .C(g35), .Y(n6432));
NAND2X1  g1793(.A(g102), .B(n4620), .Y(n6433));
NAND2X1  g1794(.A(n6433), .B(n6432), .Y(n1398));
NOR3X1   g1795(.A(n5021), .B(n4988_1), .C(n5616), .Y(n6435));
MX2X1    g1796(.A(g3853), .B(n3747), .S0(n6435), .Y(n6436));
AND2X1   g1797(.A(n6436), .B(g35), .Y(n1403));
INVX1    g1798(.A(g28753), .Y(n6438));
NAND4X1  g1799(.A(g5283), .B(g5297), .C(g5343), .D(g5357), .Y(n6439_1));
NOR2X1   g1800(.A(n6439_1), .B(n6438), .Y(n6440));
MX2X1    g1801(.A(g5134), .B(g5128), .S0(n6440), .Y(n6441));
MX2X1    g1802(.A(g5128), .B(n6441), .S0(g35), .Y(n1408));
AND2X1   g1803(.A(g3881), .B(g35), .Y(n1418));
NOR2X1   g1804(.A(n5569), .B(n5567), .Y(n6444_1));
INVX1    g1805(.A(g2476), .Y(n6445));
OAI21X1  g1806(.A0(n6204), .A1(n4917), .B0(n6445), .Y(n6446));
MX2X1    g1807(.A(g2485), .B(n6446), .S0(n6444_1), .Y(n6447));
MX2X1    g1808(.A(g2491), .B(n6447), .S0(g35), .Y(n1423));
INVX1    g1809(.A(g925), .Y(n6449_1));
INVX1    g1810(.A(g914), .Y(n6450));
INVX1    g1811(.A(g911), .Y(n6451));
INVX1    g1812(.A(g907), .Y(n6452));
NAND4X1  g1813(.A(g904), .B(g1227), .C(g921), .D(g936), .Y(n6453_1));
NOR4X1   g1814(.A(n6452), .B(n6451), .C(n6450), .D(n6453_1), .Y(n6454));
NAND2X1  g1815(.A(n6454), .B(g918), .Y(n6455));
AND2X1   g1816(.A(g1227), .B(g925), .Y(n6456));
MX2X1    g1817(.A(n6449_1), .B(n6456), .S0(n6455), .Y(n6457));
MX2X1    g1818(.A(g918), .B(n6457), .S0(g35), .Y(n1428));
OR2X1    g1819(.A(n5368), .B(g22), .Y(n6459));
OR2X1    g1820(.A(n5368), .B(n5282), .Y(n6460));
NAND2X1  g1821(.A(n6460), .B(n6459), .Y(n1433));
NOR3X1   g1822(.A(g5517), .B(g5523), .C(g5511), .Y(n6462));
NAND3X1  g1823(.A(n6462), .B(n4868), .C(g5535), .Y(n6463_1));
MX2X1    g1824(.A(n5592_1), .B(g5555), .S0(n6463_1), .Y(n6464));
MX2X1    g1825(.A(g5559), .B(n6464), .S0(g35), .Y(n1438));
INVX1    g1826(.A(n5506), .Y(n6466));
AOI21X1  g1827(.A0(n5566), .A1(n4803_1), .B0(n5564_1), .Y(n6467));
NAND2X1  g1828(.A(g2715), .B(n6307), .Y(n6468_1));
NOR4X1   g1829(.A(n6467), .B(n6466), .C(n4925_1), .D(n6468_1), .Y(n6469));
NOR2X1   g1830(.A(n4941), .B(g1783), .Y(n6470));
XOR2X1   g1831(.A(n6470), .B(g110), .Y(n6471));
MX2X1    g1832(.A(g1798), .B(n6471), .S0(n6469), .Y(n6472));
MX2X1    g1833(.A(g1783), .B(n6472), .S0(g35), .Y(n1448));
NAND4X1  g1834(.A(g4057), .B(g4064), .C(g4082), .D(g4141), .Y(n6474));
XOR2X1   g1835(.A(n6474), .B(g4076), .Y(n6475));
NAND2X1  g1836(.A(n6475), .B(g4169), .Y(n6476));
MX2X1    g1837(.A(g4082), .B(n6476), .S0(g35), .Y(n1453));
NOR3X1   g1838(.A(n5368), .B(n5286), .C(n5616), .Y(n6478_1));
NOR3X1   g1839(.A(g4072), .B(g2941), .C(g4153), .Y(n6479));
OR2X1    g1840(.A(n6479), .B(n4620), .Y(n6480));
OAI22X1  g1841(.A0(n6478_1), .A1(n6480), .B0(n4786), .B1(g35), .Y(n1458));
NOR3X1   g1842(.A(g3881), .B(n4849), .C(n4848), .Y(n6482));
MX2X1    g1843(.A(g3905), .B(n5592_1), .S0(n6482), .Y(n6483_1));
MX2X1    g1844(.A(g3953), .B(n6483_1), .S0(g35), .Y(n1463));
MX2X1    g1845(.A(n5675), .B(n5674_1), .S0(n5673), .Y(n6485));
MX2X1    g1846(.A(g758), .B(n6485), .S0(g35), .Y(n1468));
NOR4X1   g1847(.A(g6203), .B(g6209), .C(g6215), .D(n6099), .Y(n6487));
MX2X1    g1848(.A(g6255), .B(n5592_1), .S0(n6487), .Y(n6488_1));
MX2X1    g1849(.A(g6259), .B(n6488_1), .S0(g35), .Y(n1473));
MX2X1    g1850(.A(g4427), .B(g4423), .S0(g35), .Y(n1478));
INVX1    g1851(.A(g4864), .Y(n6491));
AOI21X1  g1852(.A0(n6193), .A1(g35), .B0(n6491), .Y(n1483));
INVX1    g1853(.A(n5368), .Y(n3393));
NOR3X1   g1854(.A(n5019), .B(n5031), .C(n5616), .Y(n6494));
MX2X1    g1855(.A(g4722), .B(n3393), .S0(n6494), .Y(n6495));
MX2X1    g1856(.A(g4717), .B(n6495), .S0(g35), .Y(n1488));
AOI21X1  g1857(.A0(g640), .A1(n6133), .B0(n5296), .Y(n6497));
MX2X1    g1858(.A(n5296), .B(n6497), .S0(n6144), .Y(n6498_1));
MX2X1    g1859(.A(g582), .B(n6498_1), .S0(g35), .Y(n1493));
NAND2X1  g1860(.A(g1636), .B(n5757), .Y(n6500));
AOI21X1  g1861(.A0(n5566), .A1(n5505), .B0(n5564_1), .Y(n6501));
NOR4X1   g1862(.A(n5787_1), .B(n4629), .C(g1657), .D(n6501), .Y(n6502_1));
MX2X1    g1863(.A(g1632), .B(n6500), .S0(n6502_1), .Y(n6503));
MX2X1    g1864(.A(g1612), .B(n6503), .S0(g35), .Y(n1503));
INVX1    g1865(.A(n6421), .Y(n6505));
INVX1    g1866(.A(g5290), .Y(n6506));
INVX1    g1867(.A(g5276), .Y(n6507_1));
OAI22X1  g1868(.A0(n6507_1), .A1(g5320), .B0(n6506), .B1(g5313), .Y(n6508));
MX2X1    g1869(.A(g5308), .B(n6507_1), .S0(g5283), .Y(n6509));
INVX1    g1870(.A(g5320), .Y(n6510));
OAI21X1  g1871(.A0(n6510), .A1(g5290), .B0(g35), .Y(n6511));
NOR4X1   g1872(.A(n6509), .B(n6508), .C(n6505), .D(n6511), .Y(n1508));
INVX1    g1873(.A(g1459), .Y(n6513));
NOR3X1   g1874(.A(g1514), .B(g1526), .C(n6513), .Y(n6514));
MX2X1    g1875(.A(g1495), .B(g1489), .S0(n6514), .Y(n6515));
MX2X1    g1876(.A(g1489), .B(n6515), .S0(g35), .Y(n1518));
INVX1    g1877(.A(g1437), .Y(n6517_1));
INVX1    g1878(.A(g1478), .Y(n6518));
NOR3X1   g1879(.A(n4712_1), .B(n4711), .C(g1319), .Y(n6519));
XOR2X1   g1880(.A(n6519), .B(n6518), .Y(n6520));
OR2X1    g1881(.A(g1489), .B(g1442), .Y(n6521));
AOI21X1  g1882(.A0(n6521), .A1(n6517_1), .B0(n6520), .Y(n6522_1));
NOR3X1   g1883(.A(n5549), .B(g1526), .C(n6513), .Y(n6523));
MX2X1    g1884(.A(g1437), .B(n6522_1), .S0(n6523), .Y(n6524));
MX2X1    g1885(.A(g1442), .B(n6524), .S0(g35), .Y(n1528));
NAND2X1  g1886(.A(g6395), .B(n6279), .Y(n6526_1));
INVX1    g1887(.A(g6381), .Y(n6527));
NAND3X1  g1888(.A(n6527), .B(g6251), .C(g6322), .Y(n6528));
NAND3X1  g1889(.A(g6381), .B(g6351), .C(g6239), .Y(n6529));
AOI21X1  g1890(.A0(n6529), .A1(n6528), .B0(n6526_1), .Y(n6530));
NAND4X1  g1891(.A(n6527), .B(g6365), .C(g6271), .D(n5196_1), .Y(n6531_1));
NAND2X1  g1892(.A(n6277), .B(g6336), .Y(n6532));
NAND3X1  g1893(.A(g6346), .B(n6527), .C(g6247), .Y(n6533));
OAI21X1  g1894(.A0(n6533), .A1(n6532), .B0(n6531_1), .Y(n6534));
NOR2X1   g1895(.A(n6534), .B(n6530), .Y(n6535));
AND2X1   g1896(.A(g6381), .B(g6365), .Y(n6536_1));
NAND4X1  g1897(.A(g6263), .B(g6395), .C(n6279), .D(n6536_1), .Y(n6537));
NAND4X1  g1898(.A(g6295), .B(g6381), .C(g6373), .D(n5196_1), .Y(n6538));
NOR2X1   g1899(.A(g6395), .B(g6336), .Y(n6539));
NAND4X1  g1900(.A(g6346), .B(g6381), .C(g6235), .D(n6539), .Y(n6540));
AND2X1   g1901(.A(g6381), .B(g6369), .Y(n6541_1));
NAND4X1  g1902(.A(g6279), .B(n6277), .C(g6336), .D(n6541_1), .Y(n6542));
NAND4X1  g1903(.A(n6540), .B(n6538), .C(n6537), .D(n6542), .Y(n6543));
NAND4X1  g1904(.A(n6527), .B(g6369), .C(g6287), .D(n6539), .Y(n6544));
NAND3X1  g1905(.A(g6303), .B(n6527), .C(g6373), .Y(n6545));
OAI21X1  g1906(.A0(n6545), .A1(n6526_1), .B0(n6544), .Y(n6546_1));
NAND4X1  g1907(.A(g6381), .B(g6243), .C(g6377), .D(n6539), .Y(n6547));
NAND4X1  g1908(.A(g6381), .B(g6311), .C(g6322), .D(n5196_1), .Y(n6548));
NAND2X1  g1909(.A(n6548), .B(n6547), .Y(n6549));
NOR3X1   g1910(.A(n6549), .B(n6546_1), .C(n6543), .Y(n6550_1));
INVX1    g1911(.A(g6351), .Y(n6551));
XOR2X1   g1912(.A(g6381), .B(n6551), .Y(n6552));
AND2X1   g1913(.A(g6283), .B(g6358), .Y(n6553));
AND2X1   g1914(.A(n6553), .B(n5196_1), .Y(n6554));
NAND3X1  g1915(.A(n6539), .B(g6275), .C(g6329), .Y(n6555_1));
NAND4X1  g1916(.A(g6395), .B(n6279), .C(g6291), .D(g6358), .Y(n6556));
AOI21X1  g1917(.A0(n6556), .A1(n6555_1), .B0(n6552), .Y(n6557));
AOI21X1  g1918(.A0(n6554), .A1(n6552), .B0(n6557), .Y(n6558));
NAND4X1  g1919(.A(g6307), .B(n6277), .C(g6336), .D(g6315), .Y(n6559));
NOR2X1   g1920(.A(n6559), .B(n6552), .Y(n6560_1));
NAND4X1  g1921(.A(n6527), .B(g6351), .C(g6255), .D(n5196_1), .Y(n6561));
NAND3X1  g1922(.A(n6527), .B(g6259), .C(g6377), .Y(n6562));
OAI21X1  g1923(.A0(n6562), .A1(n6532), .B0(n6561), .Y(n6563));
INVX1    g1924(.A(n6552), .Y(n6564));
NAND3X1  g1925(.A(n6539), .B(g6299), .C(g6315), .Y(n6565_1));
NAND4X1  g1926(.A(g6267), .B(n6277), .C(g6336), .D(g6329), .Y(n6566));
AOI21X1  g1927(.A0(n6566), .A1(n6565_1), .B0(n6564), .Y(n6567));
NOR3X1   g1928(.A(n6567), .B(n6563), .C(n6560_1), .Y(n6568));
NAND4X1  g1929(.A(n6558), .B(n6550_1), .C(n6535), .D(n6568), .Y(n6569));
AND2X1   g1930(.A(n5909_1), .B(g6154), .Y(n6570_1));
XOR2X1   g1931(.A(n6570_1), .B(n6569), .Y(n6571));
MX2X1    g1932(.A(g6154), .B(n6571), .S0(n5907), .Y(n6572));
MX2X1    g1933(.A(g6159), .B(n6572), .S0(g35), .Y(n1533));
NOR3X1   g1934(.A(g5527), .B(n4867), .C(n4866_1), .Y(n6574));
MX2X1    g1935(.A(g5567), .B(n5592_1), .S0(n6574), .Y(n6575_1));
MX2X1    g1936(.A(g5611), .B(n6575_1), .S0(g35), .Y(n1543));
NAND2X1  g1937(.A(g1772), .B(n5834), .Y(n6577));
AOI21X1  g1938(.A0(n5627), .A1(n5621), .B0(n6577), .Y(n6578));
MX2X1    g1939(.A(g1752), .B(n5624), .S0(n6578), .Y(n6579));
MX2X1    g1940(.A(g1756), .B(n6579), .S0(g35), .Y(n1548));
OAI21X1  g1941(.A0(n6204), .A1(n4924), .B0(n5838), .Y(n6581));
MX2X1    g1942(.A(g1917), .B(n6581), .S0(n6202), .Y(n6582));
MX2X1    g1943(.A(g1894), .B(n6582), .S0(g35), .Y(n1553));
NAND3X1  g1944(.A(n5663), .B(n5661), .C(n5654), .Y(n6584));
MX2X1    g1945(.A(n5664), .B(n5665_1), .S0(n6584), .Y(n6585_1));
MX2X1    g1946(.A(g739), .B(n6585_1), .S0(g35), .Y(n1558));
INVX1    g1947(.A(g3021), .Y(n6587));
INVX1    g1948(.A(g3004), .Y(n6588));
NOR4X1   g1949(.A(n6587), .B(n5573_1), .C(n5585), .D(n6588), .Y(n6589));
NAND3X1  g1950(.A(n6589), .B(g3025), .C(g3029), .Y(n6590_1));
NOR2X1   g1951(.A(n6590_1), .B(n5576), .Y(n6591));
INVX1    g1952(.A(g3025), .Y(n6592));
INVX1    g1953(.A(g3010), .Y(n6593));
NOR4X1   g1954(.A(g3021), .B(n6593), .C(g3017), .D(g3004), .Y(n6594));
NAND3X1  g1955(.A(n6594), .B(n6592), .C(n5578_1), .Y(n6595_1));
NOR2X1   g1956(.A(n6595_1), .B(g3034), .Y(n6596));
OAI21X1  g1957(.A0(n6596), .A1(n6591), .B0(n5575), .Y(n6597));
OR4X1    g1958(.A(n6591), .B(n5584), .C(n5575), .D(n6596), .Y(n6598));
NAND2X1  g1959(.A(n6598), .B(n6597), .Y(n6599));
MX2X1    g1960(.A(g3034), .B(n6599), .S0(g35), .Y(n1563));
MX2X1    g1961(.A(g4737), .B(n5462), .S0(n6494), .Y(n6601));
MX2X1    g1962(.A(g4722), .B(n6601), .S0(g35), .Y(n1568));
AND2X1   g1963(.A(g113), .B(g35), .Y(n1573));
NOR4X1   g1964(.A(g6227), .B(g6209), .C(n4871_1), .D(n6208), .Y(n6604));
MX2X1    g1965(.A(g6267), .B(n5592_1), .S0(n6604), .Y(n6605_1));
MX2X1    g1966(.A(g6239), .B(n6605_1), .S0(g35), .Y(n1578));
AND2X1   g1967(.A(g3431), .B(g3423), .Y(n6607));
AND2X1   g1968(.A(n6607), .B(g3436), .Y(n6608));
XOR2X1   g1969(.A(n6608), .B(g3440), .Y(n6609_1));
MX2X1    g1970(.A(g3436), .B(n6609_1), .S0(g35), .Y(n1583));
MX2X1    g1971(.A(g1442), .B(g1495), .S0(n6514), .Y(n6611));
MX2X1    g1972(.A(g1495), .B(n6611), .S0(g35), .Y(n1593));
MX2X1    g1973(.A(g5965), .B(n5592_1), .S0(n4863), .Y(n6614));
MX2X1    g1974(.A(g5961), .B(n6614), .S0(g35), .Y(n1598));
NAND2X1  g1975(.A(g4474), .B(g35), .Y(n6616));
NAND2X1  g1976(.A(g4474), .B(n4620), .Y(n6617));
NAND2X1  g1977(.A(n6617), .B(n6616), .Y(n1603));
MX2X1    g1978(.A(g1233), .B(g1227), .S0(g1083), .Y(n6619));
MX2X1    g1979(.A(g1246), .B(n6619), .S0(g35), .Y(n1608));
INVX1    g1980(.A(g4633), .Y(n6621));
NAND4X1  g1981(.A(n5850_1), .B(g4621), .C(g35), .D(g4633), .Y(n6622));
OAI22X1  g1982(.A0(n5847), .A1(n6622), .B0(n6621), .B1(g35), .Y(n1613));
INVX1    g1983(.A(g5170), .Y(n6624));
NOR4X1   g1984(.A(n4643), .B(n5610), .C(g5180), .D(n6624), .Y(n6625));
MX2X1    g1985(.A(g5264), .B(n5592_1), .S0(n6625), .Y(n6626));
MX2X1    g1986(.A(g5248), .B(n6626), .S0(g35), .Y(n1618));
INVX1    g1987(.A(n5863), .Y(n6628_1));
INVX1    g1988(.A(g2587), .Y(n6629));
OAI21X1  g1989(.A0(n6204), .A1(n4919), .B0(n6629), .Y(n6630));
MX2X1    g1990(.A(g2610), .B(n6630), .S0(n6628_1), .Y(n6631));
MX2X1    g1991(.A(g2587), .B(n6631), .S0(g35), .Y(n1628));
MX2X1    g1992(.A(g5160), .B(n3393), .S0(n6029), .Y(n6633_1));
AND2X1   g1993(.A(n6633_1), .B(g35), .Y(n1633));
INVX1    g1994(.A(g5406), .Y(n6635));
NOR2X1   g1995(.A(g5401), .B(n6635), .Y(n6636));
INVX1    g1996(.A(g5396), .Y(n6637));
INVX1    g1997(.A(g5390), .Y(n6638_1));
NOR3X1   g1998(.A(n6638_1), .B(n6637), .C(g84), .Y(n6639));
INVX1    g1999(.A(g5385), .Y(n6640));
NOR3X1   g2000(.A(n6638_1), .B(n6640), .C(n5495), .Y(n6641));
OAI21X1  g2001(.A0(n6641), .A1(n6639), .B0(n6636), .Y(n6642));
AND2X1   g2002(.A(g5366), .B(g5401), .Y(n6643_1));
NAND4X1  g2003(.A(n6638_1), .B(n6640), .C(g84), .D(n6643_1), .Y(n6644));
NAND4X1  g2004(.A(n6638_1), .B(n6637), .C(n5495), .D(n6643_1), .Y(n6645));
NAND3X1  g2005(.A(n6645), .B(n6644), .C(n6642), .Y(n6646));
INVX1    g2006(.A(g5360), .Y(n6647));
OAI21X1  g2007(.A0(g5366), .A1(g5406), .B0(n6647), .Y(n6648_1));
INVX1    g2008(.A(g5366), .Y(n6649));
NAND3X1  g2009(.A(n6649), .B(n6635), .C(g5360), .Y(n6650));
OAI21X1  g2010(.A0(n6648_1), .A1(n6646), .B0(n6650), .Y(n6651));
MX2X1    g2011(.A(g5366), .B(n6651), .S0(g35), .Y(n1638));
INVX1    g2012(.A(g5863), .Y(n6653_1));
OR2X1    g2013(.A(g5881), .B(g5873), .Y(n6654));
NOR3X1   g2014(.A(n6654), .B(g5857), .C(n6653_1), .Y(n6655));
MX2X1    g2015(.A(g5933), .B(n5592_1), .S0(n6655), .Y(n6656));
MX2X1    g2016(.A(g5917), .B(n6656), .S0(g35), .Y(n1643));
INVX1    g2017(.A(g1454), .Y(n6658_1));
XOR2X1   g2018(.A(n6519), .B(n5331), .Y(n6659));
AOI21X1  g2019(.A0(n6521), .A1(n6658_1), .B0(n6659), .Y(n6660));
NOR3X1   g2020(.A(g1514), .B(n6000_1), .C(n6513), .Y(n6661));
MX2X1    g2021(.A(g1454), .B(n6660), .S0(n6661), .Y(n6662_1));
MX2X1    g2022(.A(g1478), .B(n6662_1), .S0(g35), .Y(n1648));
NOR2X1   g2023(.A(n5657), .B(n5655_1), .Y(n6664));
MX2X1    g2024(.A(g753), .B(g732), .S0(n6664), .Y(n6665));
MX2X1    g2025(.A(g732), .B(n6665), .S0(g35), .Y(n1653));
NAND2X1  g2026(.A(n5016), .B(n4984_1), .Y(n6667));
OAI21X1  g2027(.A0(n5425_1), .A1(n5405_1), .B0(g12), .Y(n6668));
NOR2X1   g2028(.A(n6668), .B(n6667), .Y(n6669));
OAI21X1  g2029(.A0(n4717_1), .A1(g1296), .B0(g35), .Y(n6670));
OAI22X1  g2030(.A0(n6669), .A1(n6670), .B0(n5243), .B1(g35), .Y(n1658));
MX2X1    g2031(.A(g3151), .B(n4447), .S0(n6435), .Y(n6672));
AND2X1   g2032(.A(n6672), .B(g35), .Y(n1663));
NOR4X1   g2033(.A(n4995), .B(n5616), .C(g28), .D(n5001), .Y(n6674));
AND2X1   g2034(.A(n6674), .B(n4586), .Y(n6675));
OAI21X1  g2035(.A0(g34), .A1(g2980), .B0(g35), .Y(n6676_1));
OAI22X1  g2036(.A0(n6675), .A1(n6676_1), .B0(n5431), .B1(g35), .Y(n1668));
INVX1    g2037(.A(g6675), .Y(n6678));
INVX1    g2038(.A(g6704), .Y(n6679));
NAND2X1  g2039(.A(g6661), .B(g6697), .Y(n6680));
NOR3X1   g2040(.A(n6680), .B(n6679), .C(n6678), .Y(n6681_1));
XOR2X1   g2041(.A(n6681_1), .B(g6727), .Y(n6682));
MX2X1    g2042(.A(g6723), .B(n6682), .S0(g35), .Y(n1673));
OAI21X1  g2043(.A0(n4835), .A1(n4834), .B0(g3530), .Y(n6684));
NAND3X1  g2044(.A(g3522), .B(g3518), .C(n4833), .Y(n6685_1));
AOI21X1  g2045(.A0(n6685_1), .A1(n6684), .B0(n5732), .Y(n6686));
MX2X1    g2046(.A(g3522), .B(n6686), .S0(g35), .Y(n1678));
AND2X1   g2047(.A(g4741), .B(n4620), .Y(n1683));
INVX1    g2048(.A(g4076), .Y(n6689));
NOR4X1   g2049(.A(n4830), .B(n4840), .C(n6689), .D(n6474), .Y(n6690_1));
NAND3X1  g2050(.A(n6690_1), .B(g4108), .C(g4098), .Y(n6691));
XOR2X1   g2051(.A(n6691), .B(g4104), .Y(n6692));
NAND2X1  g2052(.A(n6692), .B(g4169), .Y(n6693));
MX2X1    g2053(.A(g4108), .B(n6693), .S0(g35), .Y(n1688));
MX2X1    g2054(.A(g1532), .B(g1521), .S0(g1500), .Y(n6695));
MX2X1    g2055(.A(g1306), .B(n6695), .S0(g35), .Y(n1693));
XOR2X1   g2056(.A(g4308), .B(g4304), .Y(n6697));
XOR2X1   g2057(.A(n6697), .B(g4304), .Y(n6698));
NOR2X1   g2058(.A(n6698), .B(n4620), .Y(n1698));
OAI21X1  g2059(.A0(n5541_1), .A1(g134), .B0(n5363), .Y(n6700));
NOR3X1   g2060(.A(g2704), .B(g2697), .C(n5417), .Y(n6701));
NOR2X1   g2061(.A(n6701), .B(n6700), .Y(n6702));
INVX1    g2062(.A(n6702), .Y(n6703_1));
AOI21X1  g2063(.A0(n6701), .A1(n5524), .B0(n6700), .Y(n6704));
OAI21X1  g2064(.A0(n6703_1), .A1(n5540), .B0(n6704), .Y(n6705));
NAND4X1  g2065(.A(g1322), .B(g1404), .C(n6000_1), .D(g1514), .Y(n6706));
OAI21X1  g2066(.A0(n6706), .A1(n5548), .B0(g1418), .Y(n6707));
INVX1    g2067(.A(g2153), .Y(n6708_1));
NAND2X1  g2068(.A(g2197), .B(n6708_1), .Y(n6709));
AOI21X1  g2069(.A0(n6707), .A1(n6702), .B0(n6709), .Y(n6710));
MX2X1    g2070(.A(g2177), .B(n6705), .S0(n6710), .Y(n6711));
MX2X1    g2071(.A(g2181), .B(n6711), .S0(g35), .Y(n1703));
INVX1    g2072(.A(g3103), .Y(n6713_1));
AOI21X1  g2073(.A0(g3096), .A1(n6713_1), .B0(g3010), .Y(n6714));
OR2X1    g2074(.A(g3092), .B(n4620), .Y(n6715));
OAI22X1  g2075(.A0(n6714), .A1(n6715), .B0(n6713_1), .B1(g35), .Y(n1708));
NAND2X1  g2076(.A(n3220), .B(n5282), .Y(n6717));
NAND2X1  g2077(.A(n3220), .B(g22), .Y(n6718_1));
NAND2X1  g2078(.A(n6718_1), .B(n6717), .Y(n1713));
NOR2X1   g2079(.A(n4818), .B(g4709), .Y(n6720));
NOR3X1   g2080(.A(n4809), .B(g4818), .C(g4809), .Y(n6721));
AOI21X1  g2081(.A0(n4970), .A1(n6720), .B0(n6721), .Y(n6722));
MX2X1    g2082(.A(g4760), .B(g101), .S0(n6721), .Y(n6723_1));
MX2X1    g2083(.A(n6723_1), .B(g4754), .S0(n6722), .Y(n6724));
MX2X1    g2084(.A(g4760), .B(n6724), .S0(g35), .Y(n1718));
MX2X1    g2085(.A(g1189), .B(g1178), .S0(g1157), .Y(n6726));
MX2X1    g2086(.A(g962), .B(n6726), .S0(g35), .Y(n1723));
NAND3X1  g2087(.A(n5551_1), .B(n5545), .C(g2287), .Y(n6728_1));
INVX1    g2088(.A(n5552), .Y(n6729));
NAND4X1  g2089(.A(n5637), .B(g112), .C(n4824), .D(n5139), .Y(n6730));
AOI21X1  g2090(.A0(g2331), .A1(n6032), .B0(g2361), .Y(n6731));
NAND3X1  g2091(.A(n6731), .B(n6730), .C(n6729), .Y(n6732));
AOI21X1  g2092(.A0(n6732), .A1(n6728_1), .B0(n4620), .Y(n1728));
AND2X1   g2093(.A(g4258), .B(g4264), .Y(n6734));
AND2X1   g2094(.A(n6734), .B(g4269), .Y(n6735));
XOR2X1   g2095(.A(n6735), .B(g4273), .Y(n6736));
MX2X1    g2096(.A(g4269), .B(n6736), .S0(g35), .Y(n1733));
OR4X1    g2097(.A(n6037), .B(n6036), .C(g1389), .D(n6038_1), .Y(n6738));
OAI21X1  g2098(.A0(n6038_1), .A1(n6037), .B0(g1389), .Y(n6739));
NAND2X1  g2099(.A(n6739), .B(n6738), .Y(n6740));
MX2X1    g2100(.A(g1384), .B(n6740), .S0(g35), .Y(n1738));
MX2X1    g2101(.A(g1706), .B(g1700), .S0(n5762), .Y(n6742_1));
MX2X1    g2102(.A(g1700), .B(n6742_1), .S0(g35), .Y(n1743));
INVX1    g2103(.A(g4681), .Y(n6744));
NOR4X1   g2104(.A(g4785), .B(n4815), .C(n4814), .D(n4723), .Y(n6745));
AOI21X1  g2105(.A0(n6745), .A1(n4721), .B0(n6744), .Y(n6746));
INVX1    g2106(.A(n6746), .Y(n6747_1));
NAND4X1  g2107(.A(g6049), .B(g5976), .C(g5990), .D(g6035), .Y(n6748));
NOR2X1   g2108(.A(n6748), .B(n6747_1), .Y(n6749));
XOR2X1   g2109(.A(n6749), .B(g5835), .Y(n6750));
MX2X1    g2110(.A(g5831), .B(n6750), .S0(g35), .Y(n1748));
INVX1    g2111(.A(g1157), .Y(n6752_1));
NAND2X1  g2112(.A(g1183), .B(n4665), .Y(n6753));
INVX1    g2113(.A(n4708), .Y(n6754));
NAND3X1  g2114(.A(g1002), .B(g1036), .C(g1024), .Y(n6755));
NOR3X1   g2115(.A(n6755), .B(n6058_1), .C(n6050), .Y(n6756));
INVX1    g2116(.A(g1178), .Y(n6757_1));
INVX1    g2117(.A(g996), .Y(n6758));
NOR4X1   g2118(.A(n6758), .B(g1189), .C(n6757_1), .D(n6752_1), .Y(n6759));
OAI21X1  g2119(.A0(n6756), .A1(n6754), .B0(n6759), .Y(n6760));
AOI21X1  g2120(.A0(n6753), .A1(g1193), .B0(n6760), .Y(n6761));
OAI21X1  g2121(.A0(n6761), .A1(g1171), .B0(n6752_1), .Y(n6762_1));
OAI21X1  g2122(.A0(n6761), .A1(n4665), .B0(g1157), .Y(n6763));
AOI21X1  g2123(.A0(n6763), .A1(n6762_1), .B0(n4620), .Y(n1753));
XOR2X1   g2124(.A(n6734), .B(g4269), .Y(n6765));
MX2X1    g2125(.A(g4264), .B(n6765), .S0(g35), .Y(n1758));
MX2X1    g2126(.A(g2399), .B(g2393), .S0(n5553), .Y(n6768));
MX2X1    g2127(.A(g2393), .B(n6768), .S0(g35), .Y(n1763));
NOR3X1   g2128(.A(n5767), .B(n6411), .C(n5779), .Y(n6770));
NOR3X1   g2129(.A(n5781), .B(g3368), .C(g3355), .Y(n6771));
OAI21X1  g2130(.A0(n6771), .A1(n6770), .B0(n6410), .Y(n6772_1));
NOR2X1   g2131(.A(n6771), .B(n6770), .Y(n6773));
NAND2X1  g2132(.A(n6773), .B(g3372), .Y(n6774));
OAI21X1  g2133(.A0(n6774), .A1(n5778_1), .B0(n6772_1), .Y(n6775));
MX2X1    g2134(.A(g3368), .B(n6775), .S0(g35), .Y(n1768));
NOR4X1   g2135(.A(n4963), .B(n4962), .C(n4959_1), .D(n4960), .Y(n6777_1));
INVX1    g2136(.A(n6777_1), .Y(n6778));
AND2X1   g2137(.A(n6778), .B(n6192), .Y(n6779));
NOR2X1   g2138(.A(n4961), .B(n4962), .Y(n6780));
NOR3X1   g2139(.A(n4960), .B(g4983), .C(n4959_1), .Y(n6781));
OAI21X1  g2140(.A0(n6781), .A1(n6780), .B0(n6779), .Y(n6782_1));
NAND2X1  g2141(.A(g5008), .B(n4620), .Y(n6783));
OAI21X1  g2142(.A0(n6782_1), .A1(n4620), .B0(n6783), .Y(n1773));
NOR4X1   g2143(.A(g5527), .B(n4867), .C(n5854), .D(n5855_1), .Y(n6785));
MX2X1    g2144(.A(g5611), .B(n5592_1), .S0(n6785), .Y(n6786));
MX2X1    g2145(.A(g5595), .B(n6786), .S0(g35), .Y(n1778));
AOI22X1  g2146(.A0(g5011), .A1(g4836), .B0(g3684), .B1(g4871), .Y(n6788));
INVX1    g2147(.A(n6788), .Y(n6789));
OAI22X1  g2148(.A0(g3333), .A1(n6491), .B0(n4959_1), .B1(g4035), .Y(n6790));
NOR4X1   g2149(.A(g4871), .B(g4864), .C(g4878), .D(g4836), .Y(n6791));
INVX1    g2150(.A(n6791), .Y(n6792_1));
OAI21X1  g2151(.A0(n6790), .A1(n6789), .B0(n6792_1), .Y(n6793));
INVX1    g2152(.A(n5928), .Y(n6794));
INVX1    g2153(.A(n4900), .Y(n6795));
NOR2X1   g2154(.A(g4975), .B(n4893), .Y(n6796));
AOI22X1  g2155(.A0(n4890), .A1(g4912), .B0(g4922), .B1(n6796), .Y(n6797_1));
NOR2X1   g2156(.A(n4896_1), .B(g4899), .Y(n6798));
AOI22X1  g2157(.A0(n6798), .A1(g4907), .B0(g4917), .B1(n4898), .Y(n6799));
AND2X1   g2158(.A(n6799), .B(n6797_1), .Y(n6800));
XOR2X1   g2159(.A(n6800), .B(n6795), .Y(n6801_1));
INVX1    g2160(.A(g4991), .Y(n6802));
NAND2X1  g2161(.A(n4963), .B(g4983), .Y(n6803));
OR2X1    g2162(.A(g4966), .B(g4991), .Y(n6804));
OAI22X1  g2163(.A0(n6803), .A1(n6802), .B0(n4962), .B1(n6804), .Y(n6805_1));
INVX1    g2164(.A(n4964_1), .Y(n6806));
INVX1    g2165(.A(g4927), .Y(n6807));
XOR2X1   g2166(.A(g4975), .B(g4899), .Y(n6808));
AOI21X1  g2167(.A0(n4898), .A1(n6807), .B0(n6808), .Y(n6809));
OR4X1    g2168(.A(g4966), .B(g4991), .C(g4983), .D(n6809), .Y(n6810_1));
NAND2X1  g2169(.A(n6810_1), .B(n6806), .Y(n6811));
AOI21X1  g2170(.A0(n6805_1), .A1(n6795), .B0(n6811), .Y(n6812));
OAI21X1  g2171(.A0(n6801_1), .A1(n6794), .B0(n6812), .Y(n6813));
NAND2X1  g2172(.A(n6813), .B(n6791), .Y(n6814));
AOI21X1  g2173(.A0(n6814), .A1(n6793), .B0(n4620), .Y(n1787));
INVX1    g2174(.A(g3139), .Y(n6816));
XOR2X1   g2175(.A(g3133), .B(n6816), .Y(n6817));
MX2X1    g2176(.A(g3143), .B(n6817), .S0(n4846_1), .Y(n6818));
MX2X1    g2177(.A(g3139), .B(n6818), .S0(g35), .Y(n1792));
NOR3X1   g2178(.A(n5368), .B(n5217), .C(n5616), .Y(n6820_1));
NAND2X1  g2179(.A(n4697_1), .B(n5341), .Y(n6821));
NAND2X1  g2180(.A(n6821), .B(g35), .Y(n6822));
OAI22X1  g2181(.A0(n6820_1), .A1(n6822), .B0(n5313_1), .B1(g35), .Y(n1797));
INVX1    g2182(.A(g3338), .Y(n6824));
INVX1    g2183(.A(g3281), .Y(n6825_1));
INVX1    g2184(.A(g3310), .Y(n6826));
NAND2X1  g2185(.A(g3267), .B(g3303), .Y(n6827));
NOR4X1   g2186(.A(n6826), .B(n6824), .C(n6825_1), .D(n6827), .Y(n6828));
INVX1    g2187(.A(g3347), .Y(n6829));
NAND2X1  g2188(.A(n6829), .B(g35), .Y(n6830_1));
OAI22X1  g2189(.A0(n6828), .A1(n6830_1), .B0(n6824), .B1(g35), .Y(n1802));
NOR4X1   g2190(.A(n4845), .B(g3179), .C(g3155), .D(n5593), .Y(n6832));
MX2X1    g2191(.A(g3235), .B(n5592_1), .S0(n6832), .Y(n6833));
MX2X1    g2192(.A(g3219), .B(n6833), .S0(g35), .Y(n1807));
INVX1    g2193(.A(g4578), .Y(n6835_1));
NAND3X1  g2194(.A(n6835_1), .B(g73), .C(n4950), .Y(n6836));
MX2X1    g2195(.A(g4540), .B(n6836), .S0(g4581), .Y(n6837));
MX2X1    g2196(.A(g4540), .B(n6837), .S0(g35), .Y(n1812));
NOR3X1   g2197(.A(n6067), .B(n5735), .C(g3512), .Y(n6839));
MX2X1    g2198(.A(g3566), .B(n5592_1), .S0(n6839), .Y(n6840_1));
MX2X1    g2199(.A(g3538), .B(n6840_1), .S0(g35), .Y(n1817));
INVX1    g2200(.A(g4552), .Y(n6842));
NOR3X1   g2201(.A(g4575), .B(g73), .C(g72), .Y(n6843));
MX2X1    g2202(.A(n6842), .B(n6843), .S0(g4581), .Y(n6844_1));
AND2X1   g2203(.A(n6844_1), .B(n5702), .Y(n6845));
NAND2X1  g2204(.A(g4561), .B(g4555), .Y(n6846));
NAND2X1  g2205(.A(g4564), .B(g4558), .Y(n6847));
NOR2X1   g2206(.A(n6847), .B(n6846), .Y(n6848));
OR2X1    g2207(.A(n5702), .B(g2988), .Y(n6849_1));
OAI21X1  g2208(.A0(n6849_1), .A1(n6848), .B0(g35), .Y(n6850));
NAND2X1  g2209(.A(g4564), .B(n4620), .Y(n6851));
OAI21X1  g2210(.A0(n6850), .A1(n6845), .B0(n6851), .Y(n1822));
INVX1    g2211(.A(g4961), .Y(n6853));
INVX1    g2212(.A(g4955), .Y(n6854_1));
NOR4X1   g2213(.A(n4896_1), .B(n6854_1), .C(n4893), .D(n4960), .Y(n6855));
AOI21X1  g2214(.A0(n6855), .A1(n5928), .B0(n4959_1), .Y(n6856));
OR2X1    g2215(.A(n6856), .B(n6853), .Y(n6857));
INVX1    g2216(.A(g4045), .Y(n6858));
INVX1    g2217(.A(g4054), .Y(n6859_1));
NAND2X1  g2218(.A(g3990), .B(n6859_1), .Y(n6860));
OAI21X1  g2219(.A0(n6860), .A1(n6858), .B0(n6853), .Y(n6861));
NOR2X1   g2220(.A(g3990), .B(g4054), .Y(n6862));
INVX1    g2221(.A(n6862), .Y(n6863));
INVX1    g2222(.A(g4049), .Y(n6864_1));
INVX1    g2223(.A(g3990), .Y(n6865));
NAND2X1  g2224(.A(n6865), .B(g4054), .Y(n6866));
MX2X1    g2225(.A(n5188), .B(n6866), .S0(n6864_1), .Y(n6867));
OAI21X1  g2226(.A0(n6863), .A1(g4045), .B0(n6867), .Y(n6868_1));
INVX1    g2227(.A(n6856), .Y(n6869));
NOR4X1   g2228(.A(n6806), .B(g4975), .C(n4893), .D(n6869), .Y(n6870));
OAI21X1  g2229(.A0(n6868_1), .A1(n6861), .B0(n6870), .Y(n6871));
AOI21X1  g2230(.A0(n6871), .A1(n6857), .B0(n4620), .Y(n1827));
INVX1    g2231(.A(g6444), .Y(n6873));
NOR2X1   g2232(.A(g6439), .B(n6873), .Y(n6874));
INVX1    g2233(.A(g6428), .Y(n6875));
INVX1    g2234(.A(g6434), .Y(n6876));
NOR3X1   g2235(.A(n6876), .B(n6875), .C(g84), .Y(n6877_1));
INVX1    g2236(.A(g6423), .Y(n6878));
NOR3X1   g2237(.A(n6878), .B(n6875), .C(n5495), .Y(n6879));
OAI21X1  g2238(.A0(n6879), .A1(n6877_1), .B0(n6874), .Y(n6880));
AND2X1   g2239(.A(g6404), .B(g6439), .Y(n6881));
NAND4X1  g2240(.A(n6878), .B(n6875), .C(g84), .D(n6881), .Y(n6882_1));
NAND4X1  g2241(.A(n6876), .B(n6875), .C(n5495), .D(n6881), .Y(n6883));
NAND3X1  g2242(.A(n6883), .B(n6882_1), .C(n6880), .Y(n6884));
INVX1    g2243(.A(g6398), .Y(n6885));
OAI21X1  g2244(.A0(g6404), .A1(g6444), .B0(n6885), .Y(n6886_1));
INVX1    g2245(.A(g6404), .Y(n6887));
NAND3X1  g2246(.A(n6887), .B(n6873), .C(g6398), .Y(n6888));
OAI21X1  g2247(.A0(n6886_1), .A1(n6884), .B0(n6888), .Y(n6889));
MX2X1    g2248(.A(g6404), .B(n6889), .S0(g35), .Y(n1832));
NOR3X1   g2249(.A(n5004), .B(n5031), .C(n5616), .Y(n6891_1));
MX2X1    g2250(.A(g4927), .B(n5462), .S0(n6891_1), .Y(n6892));
MX2X1    g2251(.A(g4912), .B(n6892), .S0(g35), .Y(n1837));
NOR4X1   g2252(.A(n5786), .B(n4937), .C(n5789), .D(n5787_1), .Y(n6894));
XOR2X1   g2253(.A(n6894), .B(g2259), .Y(n6895));
MX2X1    g2254(.A(g2255), .B(n6895), .S0(g35), .Y(n1842));
AND2X1   g2255(.A(n5506), .B(g111), .Y(n6897));
INVX1    g2256(.A(g2724), .Y(n6898));
INVX1    g2257(.A(n5509), .Y(n6899));
NOR3X1   g2258(.A(n6899), .B(n4799), .C(n6898), .Y(n6900));
OAI21X1  g2259(.A0(n4809), .A1(g113), .B0(g2827), .Y(n6901_1));
NAND4X1  g2260(.A(n5509), .B(g2729), .C(g2724), .D(n6901_1), .Y(n6902));
OAI22X1  g2261(.A0(n6900), .A1(n4798_1), .B0(n6897), .B1(n6902), .Y(n6903));
MX2X1    g2262(.A(g2827), .B(n6903), .S0(g35), .Y(n1847));
OR2X1    g2263(.A(g4405), .B(g4375), .Y(n6905));
NOR4X1   g2264(.A(g4408), .B(g4411), .C(g4414), .D(n6905), .Y(n6906_1));
AND2X1   g2265(.A(g4382), .B(g4375), .Y(n6907));
MX2X1    g2266(.A(n6907), .B(g4392), .S0(n6906_1), .Y(n6908));
MX2X1    g2267(.A(g4375), .B(n6908), .S0(g35), .Y(n1852));
MX2X1    g2268(.A(g2852), .B(n6676), .S0(n5697), .Y(n6910));
MX2X1    g2269(.A(g2844), .B(n6910), .S0(g35), .Y(n1861));
MX2X1    g2270(.A(g417), .B(g446), .S0(n5688), .Y(n6912));
AND2X1   g2271(.A(n6912), .B(g35), .Y(n1866));
MX2X1    g2272(.A(g645), .B(g681), .S0(n6389_1), .Y(n6914));
MX2X1    g2273(.A(g645), .B(n6914), .S0(g35), .Y(n1871));
MX2X1    g2274(.A(g437), .B(g441), .S0(n5688), .Y(n6916_1));
MX2X1    g2275(.A(g441), .B(n6916_1), .S0(g35), .Y(n1876));
INVX1    g2276(.A(g347), .Y(n6918));
NAND3X1  g2277(.A(n6918), .B(g344), .C(g35), .Y(n6919));
OAI21X1  g2278(.A0(n6918), .A1(g35), .B0(n6919), .Y(n1881));
NAND3X1  g2279(.A(n5632), .B(g5881), .C(n4860), .Y(n6921_1));
MX2X1    g2280(.A(n5592_1), .B(g5901), .S0(n6921_1), .Y(n6922));
MX2X1    g2281(.A(g5905), .B(n6922), .S0(g35), .Y(n1886));
NOR2X1   g2282(.A(n6317), .B(n5217), .Y(n6924));
OAI21X1  g2283(.A0(g2946), .A1(g2886), .B0(g35), .Y(n6925));
NAND2X1  g2284(.A(g2878), .B(n4620), .Y(n6926_1));
OAI21X1  g2285(.A0(n6925), .A1(n6924), .B0(n6926_1), .Y(n1891));
INVX1    g2286(.A(g3490), .Y(n6928));
XOR2X1   g2287(.A(g3484), .B(n6928), .Y(n6929));
MX2X1    g2288(.A(g3494), .B(n6929), .S0(n4836_1), .Y(n6930));
MX2X1    g2289(.A(g3490), .B(n6930), .S0(g35), .Y(n1896));
NOR3X1   g2290(.A(n5645_1), .B(n4837), .C(n4840), .Y(n6932));
NOR4X1   g2291(.A(g5523), .B(g5511), .C(n4620), .D(n6932), .Y(n1901));
NOR4X1   g2292(.A(g3518), .B(n5735), .C(n5733_1), .D(n5732), .Y(n6934));
MX2X1    g2293(.A(g3512), .B(n6934), .S0(g35), .Y(n1906));
MX2X1    g2294(.A(g1604), .B(n5756), .S0(n5762), .Y(n6937));
MX2X1    g2295(.A(g1687), .B(n6937), .S0(g35), .Y(n1911));
NAND4X1  g2296(.A(n4726), .B(g4057), .C(n4729), .D(n6252), .Y(n6939));
MX2X1    g2297(.A(g4164), .B(g4135), .S0(n6939), .Y(n6940_1));
MX2X1    g2298(.A(g4132), .B(n6940_1), .S0(g35), .Y(n1916));
XOR2X1   g2299(.A(g5084), .B(g5092), .Y(n6942));
MX2X1    g2300(.A(g5084), .B(n6942), .S0(g35), .Y(n1921));
INVX1    g2301(.A(g5990), .Y(n6944));
NAND2X1  g2302(.A(g6049), .B(n6944), .Y(n6945_1));
INVX1    g2303(.A(g6035), .Y(n6946));
NAND3X1  g2304(.A(n6946), .B(g5976), .C(g5905), .Y(n6947));
NAND3X1  g2305(.A(g6035), .B(g5893), .C(g6005), .Y(n6948));
AOI21X1  g2306(.A0(n6948), .A1(n6947), .B0(n6945_1), .Y(n6949));
NAND4X1  g2307(.A(n6946), .B(g5925), .C(g6019), .D(n5192), .Y(n6950_1));
INVX1    g2308(.A(g6049), .Y(n6951));
NAND2X1  g2309(.A(n6951), .B(g5990), .Y(n6952));
NAND3X1  g2310(.A(n6946), .B(g6000), .C(g5901), .Y(n6953));
OAI21X1  g2311(.A0(n6953), .A1(n6952), .B0(n6950_1), .Y(n6954));
NOR2X1   g2312(.A(n6954), .B(n6949), .Y(n6955_1));
AND2X1   g2313(.A(g6035), .B(g6019), .Y(n6956));
NAND4X1  g2314(.A(g6049), .B(n6944), .C(g5917), .D(n6956), .Y(n6957));
NAND4X1  g2315(.A(g6035), .B(g5949), .C(g6027), .D(n5192), .Y(n6958));
NOR2X1   g2316(.A(g6049), .B(g5990), .Y(n6959));
NAND4X1  g2317(.A(g6035), .B(g6000), .C(g5889), .D(n6959), .Y(n6960_1));
AND2X1   g2318(.A(g6035), .B(g6023), .Y(n6961));
NAND4X1  g2319(.A(n6951), .B(g5990), .C(g5933), .D(n6961), .Y(n6962));
NAND4X1  g2320(.A(n6960_1), .B(n6958), .C(n6957), .D(n6962), .Y(n6963));
NAND4X1  g2321(.A(n6946), .B(g6023), .C(g5941), .D(n6959), .Y(n6964));
NAND3X1  g2322(.A(n6946), .B(g5957), .C(g6027), .Y(n6965_1));
OAI21X1  g2323(.A0(n6965_1), .A1(n6945_1), .B0(n6964), .Y(n6966));
NAND4X1  g2324(.A(g6035), .B(g5897), .C(g6031), .D(n6959), .Y(n6967));
NAND4X1  g2325(.A(g6035), .B(g5976), .C(g5965), .D(n5192), .Y(n6968));
NAND2X1  g2326(.A(n6968), .B(n6967), .Y(n6969));
NOR3X1   g2327(.A(n6969), .B(n6966), .C(n6963), .Y(n6970_1));
XOR2X1   g2328(.A(g6035), .B(n5747), .Y(n6971));
AND2X1   g2329(.A(g5937), .B(g6012), .Y(n6972));
AND2X1   g2330(.A(n6972), .B(n5192), .Y(n6973));
NAND3X1  g2331(.A(n6959), .B(g5929), .C(g5983), .Y(n6974));
NAND4X1  g2332(.A(g6049), .B(g6012), .C(n6944), .D(g5945), .Y(n6975_1));
AOI21X1  g2333(.A0(n6975_1), .A1(n6974), .B0(n6971), .Y(n6976));
AOI21X1  g2334(.A0(n6973), .A1(n6971), .B0(n6976), .Y(n6977));
NAND4X1  g2335(.A(g5990), .B(g5961), .C(g5969), .D(n6951), .Y(n6978));
NOR2X1   g2336(.A(n6978), .B(n6971), .Y(n6979));
NAND4X1  g2337(.A(n6946), .B(g6005), .C(g5909), .D(n5192), .Y(n6980_1));
NAND3X1  g2338(.A(n6946), .B(g5913), .C(g6031), .Y(n6981));
OAI21X1  g2339(.A0(n6981), .A1(n6952), .B0(n6980_1), .Y(n6982));
INVX1    g2340(.A(n6971), .Y(n6983));
NAND3X1  g2341(.A(n6959), .B(g5953), .C(g5969), .Y(n6984_1));
NAND4X1  g2342(.A(n6951), .B(g5990), .C(g5983), .D(g5921), .Y(n6985));
AOI21X1  g2343(.A0(n6985), .A1(n6984_1), .B0(n6983), .Y(n6986));
NOR3X1   g2344(.A(n6986), .B(n6982), .C(n6979), .Y(n6987));
NAND4X1  g2345(.A(n6977), .B(n6970_1), .C(n6955_1), .D(n6987), .Y(n6988_1));
MX2X1    g2346(.A(g4831), .B(n6988_1), .S0(n6746), .Y(n6989));
MX2X1    g2347(.A(g5965), .B(n6989), .S0(g35), .Y(n1926));
XOR2X1   g2348(.A(g4382), .B(g4375), .Y(n6991));
NOR2X1   g2349(.A(g4417), .B(g4392), .Y(n6992));
MX2X1    g2350(.A(n6991), .B(n6992), .S0(n6906_1), .Y(n6993_1));
MX2X1    g2351(.A(g4388), .B(n6993_1), .S0(g35), .Y(n1931));
INVX1    g2352(.A(g6329), .Y(n6995));
INVX1    g2353(.A(g6315), .Y(n6996));
INVX1    g2354(.A(g6358), .Y(n6997));
NOR4X1   g2355(.A(n6997), .B(n6996), .C(n6995), .D(n6551), .Y(n6998_1));
AND2X1   g2356(.A(n6998_1), .B(g6381), .Y(n6999));
INVX1    g2357(.A(g6390), .Y(n7000));
NAND2X1  g2358(.A(n7000), .B(g35), .Y(n7001));
OAI22X1  g2359(.A0(n6999), .A1(n7001), .B0(n6527), .B1(g35), .Y(n1936));
NAND4X1  g2360(.A(g168), .B(g174), .C(g203), .D(n5881), .Y(n7003_1));
INVX1    g2361(.A(g513), .Y(n7004));
AND2X1   g2362(.A(g182), .B(g203), .Y(n7005));
NAND4X1  g2363(.A(g518), .B(g168), .C(n7004), .D(n7005), .Y(n7006));
NAND4X1  g2364(.A(g518), .B(n7004), .C(g174), .D(n7005), .Y(n7007));
AND2X1   g2365(.A(n7007), .B(n7006), .Y(n7008_1));
AOI21X1  g2366(.A0(n7008_1), .A1(n7003_1), .B0(n4620), .Y(n1941));
MX2X1    g2367(.A(g3965), .B(n5592_1), .S0(n4851_1), .Y(n7011));
MX2X1    g2368(.A(g3961), .B(n7011), .S0(g35), .Y(n1946));
INVX1    g2369(.A(g4749), .Y(n7013_1));
INVX1    g2370(.A(g4674), .Y(n7014));
NOR4X1   g2371(.A(n4818), .B(g4709), .C(n4817_1), .D(n4723), .Y(n7015));
AOI21X1  g2372(.A0(n7015), .A1(n4721), .B0(n7014), .Y(n7016));
OR2X1    g2373(.A(n7016), .B(n7013_1), .Y(n7017_1));
INVX1    g2374(.A(g5694), .Y(n7018));
INVX1    g2375(.A(g5703), .Y(n7019));
NAND2X1  g2376(.A(g5644), .B(n7019), .Y(n7020));
OAI21X1  g2377(.A0(n7020), .A1(n7018), .B0(n7013_1), .Y(n7021));
NOR2X1   g2378(.A(g5644), .B(g5703), .Y(n7022_1));
INVX1    g2379(.A(n7022_1), .Y(n7023));
INVX1    g2380(.A(g5698), .Y(n7024));
INVX1    g2381(.A(n5194), .Y(n7025));
INVX1    g2382(.A(g5644), .Y(n7026));
NAND2X1  g2383(.A(n7026), .B(g5703), .Y(n7027_1));
MX2X1    g2384(.A(n7025), .B(n7027_1), .S0(n7024), .Y(n7028));
OAI21X1  g2385(.A0(n7023), .A1(g5694), .B0(n7028), .Y(n7029));
INVX1    g2386(.A(n4970), .Y(n7030));
INVX1    g2387(.A(n7016), .Y(n7031));
NOR4X1   g2388(.A(n7030), .B(g4785), .C(g4709), .D(n7031), .Y(n7032_1));
OAI21X1  g2389(.A0(n7029), .A1(n7021), .B0(n7032_1), .Y(n7033));
AOI21X1  g2390(.A0(n7033), .A1(n7017_1), .B0(n4620), .Y(n1951));
INVX1    g2391(.A(n6084), .Y(n7035));
AOI21X1  g2392(.A0(n6083_1), .A1(n5524), .B0(n6082), .Y(n7036));
OAI21X1  g2393(.A0(n7035), .A1(g1242), .B0(n7036), .Y(n7037_1));
MX2X1    g2394(.A(g2008), .B(n7037_1), .S0(n6086), .Y(n7039));
MX2X1    g2395(.A(g2089), .B(n7039), .S0(g35), .Y(n1956));
INVX1    g2396(.A(g3863), .Y(n7041));
OR2X1    g2397(.A(g3881), .B(g3873), .Y(n7042_1));
NOR3X1   g2398(.A(n7042_1), .B(g3857), .C(n7041), .Y(n7043));
MX2X1    g2399(.A(g3933), .B(n5592_1), .S0(n7043), .Y(n7044));
MX2X1    g2400(.A(g3917), .B(n7044), .S0(g35), .Y(n1966));
INVX1    g2401(.A(g301), .Y(n7046));
INVX1    g2402(.A(g298), .Y(n7047_1));
NOR4X1   g2403(.A(n5661), .B(n5516_1), .C(n7047_1), .D(n6113), .Y(n7048));
NAND4X1  g2404(.A(n6121), .B(n6119), .C(n6117), .D(n7048), .Y(n7049));
NAND2X1  g2405(.A(g142), .B(g35), .Y(n7050));
OAI22X1  g2406(.A0(n7049), .A1(n7050), .B0(n7046), .B1(g35), .Y(n1971));
INVX1    g2407(.A(g3100), .Y(n7052));
AOI21X1  g2408(.A0(g3092), .A1(n7052), .B0(g3050), .Y(n7053));
OR2X1    g2409(.A(g3096), .B(n4620), .Y(n7054));
OAI22X1  g2410(.A0(n7053), .A1(n7054), .B0(n7052), .B1(g35), .Y(n1976));
INVX1    g2411(.A(g5736), .Y(n7056));
INVX1    g2412(.A(g5719), .Y(n7057));
INVX1    g2413(.A(g5752), .Y(n7058));
INVX1    g2414(.A(g5706), .Y(n7059));
INVX1    g2415(.A(g5723), .Y(n7060_1));
NOR4X1   g2416(.A(n7059), .B(n7058), .C(n7057), .D(n7060_1), .Y(n7061));
NAND3X1  g2417(.A(n7061), .B(g5727), .C(g5731), .Y(n7062));
INVX1    g2418(.A(g5731), .Y(n7063));
INVX1    g2419(.A(g5727), .Y(n7064));
INVX1    g2420(.A(g5712), .Y(n7065_1));
NOR4X1   g2421(.A(g5706), .B(g5719), .C(n7065_1), .D(g5723), .Y(n7066));
NAND3X1  g2422(.A(n7066), .B(n7064), .C(n7063), .Y(n7067));
AND2X1   g2423(.A(n7067), .B(n7062), .Y(n7068));
NOR2X1   g2424(.A(g5747), .B(n7058), .Y(n7069));
INVX1    g2425(.A(g5742), .Y(n7070_1));
NOR3X1   g2426(.A(n7070_1), .B(n7056), .C(g84), .Y(n7071));
NOR3X1   g2427(.A(n7063), .B(n7056), .C(n5495), .Y(n7072));
OAI21X1  g2428(.A0(n7072), .A1(n7071), .B0(n7069), .Y(n7073));
AND2X1   g2429(.A(g5747), .B(g5712), .Y(n7074));
NAND4X1  g2430(.A(n7063), .B(n7056), .C(g84), .D(n7074), .Y(n7075_1));
NAND4X1  g2431(.A(n7070_1), .B(n7056), .C(n5495), .D(n7074), .Y(n7076));
NAND3X1  g2432(.A(n7076), .B(n7075_1), .C(n7073), .Y(n7077));
NOR2X1   g2433(.A(n7077), .B(n7056), .Y(n7078));
MX2X1    g2434(.A(n7056), .B(n7078), .S0(n7068), .Y(n7079));
MX2X1    g2435(.A(g5731), .B(n7079), .S0(g35), .Y(n1981));
INVX1    g2436(.A(g1052), .Y(n7081));
NOR3X1   g2437(.A(g1056), .B(g1157), .C(g990), .Y(n7082));
OAI21X1  g2438(.A0(n7082), .A1(n5691), .B0(n7081), .Y(n7083));
NOR3X1   g2439(.A(n7082), .B(n5691), .C(n7081), .Y(n7084));
NOR3X1   g2440(.A(n7084), .B(g979), .C(n4620), .Y(n7085_1));
AND2X1   g2441(.A(n7085_1), .B(n7083), .Y(n1986));
ZERO     g2442(.Y(n1991));
INVX1    g2443(.A(g2028), .Y(n7088));
NOR4X1   g2444(.A(n5508), .B(g2741), .C(g2787), .D(n5565), .Y(n7089_1));
OAI21X1  g2445(.A0(n7089_1), .A1(n5564_1), .B0(n5862), .Y(n7090));
NOR3X1   g2446(.A(n7090), .B(n4943), .C(n7088), .Y(n7091));
MX2X1    g2447(.A(g2122), .B(g2116), .S0(n7091), .Y(n7092));
MX2X1    g2448(.A(g2116), .B(n7092), .S0(g35), .Y(n1999));
INVX1    g2449(.A(g2465), .Y(n7094));
NAND4X1  g2450(.A(g1322), .B(g1404), .C(g1526), .D(g1514), .Y(n7095));
OAI21X1  g2451(.A0(n7095), .A1(n5548), .B0(g1426), .Y(n7096));
OAI22X1  g2452(.A0(g1291), .A1(n5303_1), .B0(g134), .B1(n5541_1), .Y(n7097));
NOR3X1   g2453(.A(g2704), .B(n5447), .C(n5417), .Y(n7098_1));
NOR2X1   g2454(.A(n7098_1), .B(n7097), .Y(n7099));
AND2X1   g2455(.A(n7099), .B(n7096), .Y(n7100));
INVX1    g2456(.A(n7100), .Y(n7101));
NAND4X1  g2457(.A(n5637), .B(g112), .C(n4824), .D(n5138), .Y(n7102));
NAND3X1  g2458(.A(n7102), .B(n7101), .C(g2421), .Y(n7103_1));
OAI21X1  g2459(.A0(n7101), .A1(n7094), .B0(n7103_1), .Y(n7104));
MX2X1    g2460(.A(g2472), .B(n7104), .S0(g35), .Y(n2004));
AND2X1   g2461(.A(g6474), .B(g6466), .Y(n7106));
AND2X1   g2462(.A(n7106), .B(g6479), .Y(n7107));
XOR2X1   g2463(.A(n7107), .B(g6483), .Y(n7108_1));
MX2X1    g2464(.A(g6479), .B(n7108_1), .S0(g35), .Y(n2009));
NOR4X1   g2465(.A(g5857), .B(g5863), .C(g5869), .D(n6654), .Y(n7110));
MX2X1    g2466(.A(g5889), .B(n5592_1), .S0(n7110), .Y(n7111));
MX2X1    g2467(.A(g5881), .B(n7111), .S0(g35), .Y(n2014));
INVX1    g2468(.A(g4572), .Y(n7113_1));
NAND3X1  g2469(.A(n7113_1), .B(g73), .C(n4950), .Y(n7114));
MX2X1    g2470(.A(g4480), .B(n7114), .S0(g4581), .Y(n7115));
MX2X1    g2471(.A(g4480), .B(n7115), .S0(g35), .Y(n2019));
NOR3X1   g2472(.A(g358), .B(g365), .C(n4620), .Y(n2024));
INVX1    g2473(.A(g4653), .Y(n7118_1));
NOR4X1   g2474(.A(n4968), .B(g4688), .C(n7118_1), .D(n6216_1), .Y(n7119));
NOR4X1   g2475(.A(n4968), .B(n4967), .C(g4653), .D(n6216_1), .Y(n7120));
OR2X1    g2476(.A(n7120), .B(n7119), .Y(n7121));
MX2X1    g2477(.A(g4688), .B(n7121), .S0(g35), .Y(n2029));
OAI21X1  g2478(.A0(n4845), .A1(n4843), .B0(g3179), .Y(n7123_1));
NAND3X1  g2479(.A(g3171), .B(n4844), .C(g3167), .Y(n7124));
AOI21X1  g2480(.A0(n7124), .A1(n7123_1), .B0(n5765), .Y(n7125));
MX2X1    g2481(.A(g3171), .B(n7125), .S0(g35), .Y(n2034));
NAND3X1  g2482(.A(n5627), .B(n5621), .C(g1728), .Y(n7127));
AOI21X1  g2483(.A0(g1772), .A1(n5834), .B0(g1802), .Y(n7128_1));
NAND3X1  g2484(.A(n7128_1), .B(n5638), .C(n5636), .Y(n7129));
AOI21X1  g2485(.A0(n7129), .A1(n7127), .B0(n4620), .Y(n2039));
OR2X1    g2486(.A(n7097), .B(n5524), .Y(n7131));
MX2X1    g2487(.A(n7131), .B(g1585), .S0(n7099), .Y(n7132_1));
NOR3X1   g2488(.A(n7100), .B(g2421), .C(g2495), .Y(n7133));
MX2X1    g2489(.A(g2433), .B(n7132_1), .S0(n7133), .Y(n7134));
MX2X1    g2490(.A(g2514), .B(n7134), .S0(g35), .Y(n2044));
NAND4X1  g2491(.A(g3990), .B(g4054), .C(g4040), .D(g3976), .Y(n7136));
NOR2X1   g2492(.A(n7136), .B(n6869), .Y(n7137_1));
XOR2X1   g2493(.A(n7137_1), .B(g3835), .Y(n7138));
MX2X1    g2494(.A(g3831), .B(n7138), .S0(g35), .Y(n2049));
MX2X1    g2495(.A(g6187), .B(g6181), .S0(n4874), .Y(n7140));
MX2X1    g2496(.A(g6181), .B(n7140), .S0(g35), .Y(n2054));
MX2X1    g2497(.A(g4917), .B(n3747), .S0(n6891_1), .Y(n7142_1));
AND2X1   g2498(.A(n7142_1), .B(g35), .Y(n2059));
INVX1    g2499(.A(g1070), .Y(n7144));
NOR3X1   g2500(.A(n6758), .B(g1189), .C(n6757_1), .Y(n7145));
NOR3X1   g2501(.A(n7145), .B(n6753), .C(n6752_1), .Y(n7146));
NAND3X1  g2502(.A(n7146), .B(g1199), .C(n7144), .Y(n7147_1));
INVX1    g2503(.A(g1199), .Y(n7148));
INVX1    g2504(.A(n7146), .Y(n7149));
OAI21X1  g2505(.A0(n7149), .A1(n7148), .B0(g1070), .Y(n7150));
AOI21X1  g2506(.A0(n7150), .A1(n7147_1), .B0(n6761), .Y(n7151));
MX2X1    g2507(.A(g1199), .B(n7151), .S0(g35), .Y(n2064));
INVX1    g2508(.A(g832), .Y(n7153));
NAND4X1  g2509(.A(g385), .B(g370), .C(g817), .D(n6245), .Y(n7154));
NOR2X1   g2510(.A(n7154), .B(n7153), .Y(n7155));
INVX1    g2511(.A(g847), .Y(n7156));
INVX1    g2512(.A(g812), .Y(n7157_1));
AOI21X1  g2513(.A0(g837), .A1(n7157_1), .B0(n7156), .Y(n7158));
NOR2X1   g2514(.A(n7158), .B(g822), .Y(n7159));
INVX1    g2515(.A(g822), .Y(n7160));
NOR2X1   g2516(.A(n7158), .B(n7160), .Y(n7161));
MX2X1    g2517(.A(n7161), .B(n7159), .S0(n7155), .Y(n7162_1));
MX2X1    g2518(.A(g832), .B(n7162_1), .S0(g35), .Y(n2069));
INVX1    g2519(.A(g936), .Y(n7164));
NAND3X1  g2520(.A(g904), .B(g1227), .C(g921), .Y(n7165));
OR4X1    g2521(.A(n6452), .B(n7164), .C(n6451), .D(n7165), .Y(n7166));
AND2X1   g2522(.A(g1227), .B(g914), .Y(n7167_1));
MX2X1    g2523(.A(n6450), .B(n7167_1), .S0(n7166), .Y(n7168));
MX2X1    g2524(.A(g911), .B(n7168), .S0(g35), .Y(n2078));
MX2X1    g2525(.A(g4153), .B(n6265), .S0(g35), .Y(n2088));
OR2X1    g2526(.A(n6755), .B(g1008), .Y(n7171));
OAI22X1  g2527(.A0(n6053_1), .A1(g1046), .B0(n6050), .B1(n7171), .Y(n7172_1));
INVX1    g2528(.A(g969), .Y(n7173));
AOI21X1  g2529(.A0(n6053_1), .A1(n7173), .B0(n6050), .Y(n7174));
OAI21X1  g2530(.A0(n7174), .A1(n7172_1), .B0(n6059), .Y(n7175));
NAND2X1  g2531(.A(n6058_1), .B(g969), .Y(n7176));
AOI21X1  g2532(.A0(n7176), .A1(n7175), .B0(n4620), .Y(n2093));
INVX1    g2533(.A(g2811), .Y(n7178));
NOR2X1   g2534(.A(n5506), .B(n7178), .Y(n7179));
NOR3X1   g2535(.A(n6899), .B(g2729), .C(n6898), .Y(n7180));
OR4X1    g2536(.A(n6899), .B(g2729), .C(n6898), .D(n6897), .Y(n7181));
OAI22X1  g2537(.A0(n7180), .A1(n4795), .B0(n7179), .B1(n7181), .Y(n7182_1));
MX2X1    g2538(.A(g2815), .B(n7182_1), .S0(g35), .Y(n2098));
INVX1    g2539(.A(g5421), .Y(n7184));
NOR2X1   g2540(.A(g5417), .B(n7184), .Y(n7185));
NOR2X1   g2541(.A(g5413), .B(n7184), .Y(n7186));
MX2X1    g2542(.A(n7185), .B(n7186), .S0(g5428), .Y(n7187_1));
MX2X1    g2543(.A(g5421), .B(n7187_1), .S0(g35), .Y(n2103));
OR2X1    g2544(.A(n6856), .B(n6859_1), .Y(n7189));
NAND2X1  g2545(.A(n5506), .B(g93), .Y(n7190));
NOR3X1   g2546(.A(n6869), .B(n7190), .C(n5186_1), .Y(n7191));
NAND2X1  g2547(.A(n6856), .B(n6859_1), .Y(n7192_1));
OAI21X1  g2548(.A0(n7192_1), .A1(n7191), .B0(n7189), .Y(n7193));
MX2X1    g2549(.A(g4049), .B(n7193), .S0(g35), .Y(n2108));
INVX1    g2550(.A(g6187), .Y(n7195));
XOR2X1   g2551(.A(g6181), .B(n7195), .Y(n7196));
MX2X1    g2552(.A(g6191), .B(n7196), .S0(n4874), .Y(n7197_1));
MX2X1    g2553(.A(g6187), .B(n7197_1), .S0(g35), .Y(n2113));
INVX1    g2554(.A(g5073), .Y(n7199));
INVX1    g2555(.A(g5069), .Y(n7200));
AOI21X1  g2556(.A0(n7200), .A1(g35), .B0(n7199), .Y(n2118));
NOR4X1   g2557(.A(n5855_1), .B(g5523), .C(n5854), .D(n6932), .Y(n7202_1));
MX2X1    g2558(.A(g5517), .B(n7202_1), .S0(g35), .Y(n2123));
INVX1    g2559(.A(g6555), .Y(n7204));
NAND2X1  g2560(.A(g6565), .B(g6573), .Y(n7205));
NOR3X1   g2561(.A(n7205), .B(n7204), .C(g6549), .Y(n7206));
MX2X1    g2562(.A(g6637), .B(n5592_1), .S0(n7206), .Y(n7207_1));
MX2X1    g2563(.A(g6621), .B(n7207_1), .S0(g35), .Y(n2133));
MX2X1    g2564(.A(g174), .B(g182), .S0(n5601), .Y(n7209));
MX2X1    g2565(.A(g182), .B(n7209), .S0(g35), .Y(n2138));
INVX1    g2566(.A(n5758_1), .Y(n7211));
MX2X1    g2567(.A(g1246), .B(n5755), .S0(n5754), .Y(n7212_1));
OR2X1    g2568(.A(g1592), .B(g1668), .Y(n7213));
AND2X1   g2569(.A(n7213), .B(g1682), .Y(n7214));
XOR2X1   g2570(.A(n7214), .B(n7212_1), .Y(n7215));
MX2X1    g2571(.A(g1682), .B(n7215), .S0(n7211), .Y(n7216));
MX2X1    g2572(.A(g1668), .B(n7216), .S0(g35), .Y(n2143));
INVX1    g2573(.A(g351), .Y(n7218));
OR2X1    g2574(.A(g333), .B(g355), .Y(n7219));
NAND3X1  g2575(.A(n7219), .B(n7218), .C(g35), .Y(n7220));
OAI21X1  g2576(.A0(n7218), .A1(g35), .B0(n7220), .Y(n2148));
NOR3X1   g2577(.A(n6397), .B(n6753), .C(n6188), .Y(n7222));
XOR2X1   g2578(.A(g1111), .B(g1105), .Y(n7223));
MX2X1    g2579(.A(g1105), .B(n7223), .S0(n7222), .Y(n7224));
MX2X1    g2580(.A(g1111), .B(n7224), .S0(g35), .Y(n2158));
OR4X1    g2581(.A(n5508), .B(g2741), .C(g2807), .D(n5565), .Y(n7226));
AOI21X1  g2582(.A0(n7226), .A1(n5510), .B0(n6468_1), .Y(n7227));
INVX1    g2583(.A(g2319), .Y(n7228));
OAI21X1  g2584(.A0(n6204), .A1(n4918), .B0(n7228), .Y(n7229));
MX2X1    g2585(.A(g2342), .B(n7229), .S0(n7227), .Y(n7230_1));
MX2X1    g2586(.A(g2319), .B(n7230_1), .S0(g35), .Y(n2163));
NOR3X1   g2587(.A(n6099), .B(n6208), .C(n5980), .Y(n7232));
MX2X1    g2588(.A(g6307), .B(n5592_1), .S0(n7232), .Y(n7233));
MX2X1    g2589(.A(g6291), .B(n7233), .S0(g35), .Y(n2168));
MX2X1    g2590(.A(g6159), .B(g6195), .S0(n4874), .Y(n7235));
MX2X1    g2591(.A(g6195), .B(n7235), .S0(g35), .Y(n2177));
XOR2X1   g2592(.A(g2250), .B(g2246), .Y(n7237));
NOR4X1   g2593(.A(n5786), .B(g2185), .C(n5797_1), .D(n5787_1), .Y(n7238_1));
MX2X1    g2594(.A(g2255), .B(n7237), .S0(n7238_1), .Y(n7239));
MX2X1    g2595(.A(g2250), .B(n7239), .S0(g35), .Y(n2182));
INVX1    g2596(.A(g2823), .Y(n7241));
NOR2X1   g2597(.A(n5506), .B(n7241), .Y(n7242));
NOR3X1   g2598(.A(n6899), .B(n4799), .C(g2724), .Y(n7243_1));
OR4X1    g2599(.A(n6899), .B(n4799), .C(g2724), .D(n6897), .Y(n7244));
OAI22X1  g2600(.A0(n7243_1), .A1(n5563), .B0(n7242), .B1(n7244), .Y(n7245));
MX2X1    g2601(.A(g2819), .B(n7245), .S0(g35), .Y(n2187));
NOR2X1   g2602(.A(n6453_1), .B(n6452), .Y(n7247));
AND2X1   g2603(.A(g1227), .B(g911), .Y(n7248_1));
MX2X1    g2604(.A(n7248_1), .B(n6451), .S0(n7247), .Y(n7249));
MX2X1    g2605(.A(g907), .B(n7249), .S0(g35), .Y(n2192));
NAND2X1  g2606(.A(n4876_1), .B(n4828), .Y(n7251));
OAI21X1  g2607(.A0(n4877), .A1(n4828), .B0(n7251), .Y(n2197));
NOR3X1   g2608(.A(n5628), .B(n5834), .C(n5164), .Y(n7253_1));
MX2X1    g2609(.A(g1748), .B(n5624), .S0(n7253_1), .Y(n7254));
MX2X1    g2610(.A(g1752), .B(n7254), .S0(g35), .Y(n2206));
NOR2X1   g2611(.A(n5899_1), .B(n4866_1), .Y(n7256));
MX2X1    g2612(.A(g5551), .B(n5592_1), .S0(n7256), .Y(n7257));
MX2X1    g2613(.A(g5603), .B(n7257), .S0(g35), .Y(n2211));
MX2X1    g2614(.A(n7062), .B(n7067), .S0(n7056), .Y(n7259));
NOR2X1   g2615(.A(n7077), .B(n7070_1), .Y(n7260));
MX2X1    g2616(.A(n7070_1), .B(n7260), .S0(n7259), .Y(n7261));
MX2X1    g2617(.A(g5736), .B(n7261), .S0(g35), .Y(n2216));
NAND3X1  g2618(.A(n5606), .B(g3522), .C(g3530), .Y(n7263_1));
MX2X1    g2619(.A(n5592_1), .B(g3558), .S0(n7263_1), .Y(n7264));
MX2X1    g2620(.A(g3562), .B(n7264), .S0(g35), .Y(n2221));
INVX1    g2621(.A(g5495), .Y(n7266));
XOR2X1   g2622(.A(g5489), .B(n7266), .Y(n7267));
MX2X1    g2623(.A(g5499), .B(n7267), .S0(n4869), .Y(n7268_1));
MX2X1    g2624(.A(g5495), .B(n7268_1), .S0(g35), .Y(n2226));
MX2X1    g2625(.A(g2960), .B(n6708), .S0(n5617), .Y(n7270));
MX2X1    g2626(.A(g2950), .B(n7270), .S0(g35), .Y(n2231));
NAND3X1  g2627(.A(n6152), .B(g3881), .C(n4848), .Y(n7272));
MX2X1    g2628(.A(n5592_1), .B(g3901), .S0(n7272), .Y(n7273_1));
MX2X1    g2629(.A(g3905), .B(n7273_1), .S0(g35), .Y(n2236));
AOI21X1  g2630(.A0(n4964_1), .A1(n4898), .B0(n6089), .Y(n7275));
MX2X1    g2631(.A(g4894), .B(g71), .S0(n6089), .Y(n7276));
MX2X1    g2632(.A(n7276), .B(g4888), .S0(n7275), .Y(n7277));
MX2X1    g2633(.A(g4894), .B(n7277), .S0(g35), .Y(n2241));
NOR3X1   g2634(.A(g6227), .B(n4872), .C(n4871_1), .Y(n7279));
MX2X1    g2635(.A(g6251), .B(n5592_1), .S0(n7279), .Y(n7280));
MX2X1    g2636(.A(g6299), .B(n7280), .S0(g35), .Y(n2246));
AOI21X1  g2637(.A0(n5984), .A1(n6036), .B0(g1312), .Y(n7282));
INVX1    g2638(.A(g1389), .Y(n7283_1));
NAND3X1  g2639(.A(g1351), .B(g1361), .C(g1373), .Y(n7284));
MX2X1    g2640(.A(n7284), .B(n7283_1), .S0(n5984), .Y(n7285));
NAND2X1  g2641(.A(n7285), .B(n7282), .Y(n7286));
NOR2X1   g2642(.A(n7286), .B(g1373), .Y(n7287));
NOR2X1   g2643(.A(n7286), .B(g1367), .Y(n7288_1));
NOR2X1   g2644(.A(n7286), .B(g1361), .Y(n7289));
NOR2X1   g2645(.A(n7286), .B(g1345), .Y(n7290));
OR4X1    g2646(.A(n7289), .B(n7288_1), .C(n5985), .D(n7290), .Y(n7291));
MX2X1    g2647(.A(n7287), .B(g1373), .S0(n7291), .Y(n7292));
MX2X1    g2648(.A(g1367), .B(n7292), .S0(g35), .Y(n2255));
AND2X1   g2649(.A(g3179), .B(g35), .Y(n2260));
INVX1    g2650(.A(g157), .Y(n7295));
INVX1    g2651(.A(g150), .Y(n7296));
INVX1    g2652(.A(g164), .Y(n7297));
INVX1    g2653(.A(g203), .Y(n7298_1));
NOR3X1   g2654(.A(n5129), .B(g513), .C(n7298_1), .Y(n7299));
INVX1    g2655(.A(n7299), .Y(n7300));
NOR3X1   g2656(.A(g182), .B(g168), .C(g174), .Y(n7301));
OAI21X1  g2657(.A0(n7301), .A1(n7300), .B0(g691), .Y(n7302_1));
NOR2X1   g2658(.A(n7302_1), .B(n5661), .Y(n7303));
INVX1    g2659(.A(n7303), .Y(n7304));
NAND3X1  g2660(.A(n7303), .B(n7299), .C(g146), .Y(n7305));
NOR4X1   g2661(.A(n7304), .B(n7297), .C(n7296), .D(n7305), .Y(n7306_1));
INVX1    g2662(.A(g153), .Y(n7307));
NOR3X1   g2663(.A(n7302_1), .B(n5661), .C(n7307), .Y(n7308));
NAND2X1  g2664(.A(n7308), .B(n7306_1), .Y(n7309));
NOR3X1   g2665(.A(n7302_1), .B(n5661), .C(n7295), .Y(n7310_1));
MX2X1    g2666(.A(n7295), .B(n7310_1), .S0(n7309), .Y(n7311));
MX2X1    g2667(.A(g153), .B(n7311), .S0(g35), .Y(n2264));
INVX1    g2668(.A(g2791), .Y(n7313));
OAI21X1  g2669(.A0(n5506), .A1(n7313), .B0(n7243_1), .Y(n7314_1));
OAI22X1  g2670(.A0(n7243_1), .A1(n5839), .B0(n5507_1), .B1(n7314_1), .Y(n7315));
MX2X1    g2671(.A(g2787), .B(n7315), .S0(g35), .Y(n2269));
NOR4X1   g2672(.A(n4833), .B(n5735), .C(g3512), .D(g3522), .Y(n7317));
MX2X1    g2673(.A(g3574), .B(n5592_1), .S0(n7317), .Y(n7318));
MX2X1    g2674(.A(g3550), .B(n7318), .S0(g35), .Y(n2279));
INVX1    g2675(.A(g2102), .Y(n7320));
XOR2X1   g2676(.A(g2108), .B(n7320), .Y(n7321));
MX2X1    g2677(.A(g2112), .B(n7321), .S0(n6086), .Y(n7322));
MX2X1    g2678(.A(g2108), .B(n7322), .S0(g35), .Y(n2284));
NOR2X1   g2679(.A(n6317), .B(n6667), .Y(n7324_1));
OAI21X1  g2680(.A0(g1277), .A1(g1283), .B0(g35), .Y(n7325));
NAND2X1  g2681(.A(g1296), .B(n4620), .Y(n7326));
OAI21X1  g2682(.A0(n7325), .A1(n7324_1), .B0(n7326), .Y(n2289));
MX2X1    g2683(.A(g433), .B(g269), .S0(n5688), .Y(n7328));
MX2X1    g2684(.A(g437), .B(n7328), .S0(g35), .Y(n2294));
OR2X1    g2685(.A(n5669_1), .B(n5666), .Y(n7330));
MX2X1    g2686(.A(n5670), .B(n5671), .S0(n7330), .Y(n7331));
MX2X1    g2687(.A(g749), .B(n7331), .S0(g35), .Y(n2313));
INVX1    g2688(.A(g5805), .Y(n7333_1));
AOI21X1  g2689(.A0(g5798), .A1(n7333_1), .B0(g5712), .Y(n7334));
OR2X1    g2690(.A(g5794), .B(n4620), .Y(n7335));
OAI22X1  g2691(.A0(n7334), .A1(n7335), .B0(n7333_1), .B1(g35), .Y(n2318));
AND2X1   g2692(.A(g4057), .B(g4064), .Y(n7337_1));
NAND3X1  g2693(.A(n7337_1), .B(n6252), .C(n4726), .Y(n7338));
MX2X1    g2694(.A(g4164), .B(g4138), .S0(n7338), .Y(n7339));
MX2X1    g2695(.A(g4135), .B(n7339), .S0(g35), .Y(n2323));
INVX1    g2696(.A(n5845_1), .Y(n7341));
NOR4X1   g2697(.A(g4639), .B(g4643), .C(n4620), .D(n7341), .Y(n2328));
INVX1    g2698(.A(g6533), .Y(n7343));
XOR2X1   g2699(.A(g6527), .B(n7343), .Y(n7344));
MX2X1    g2700(.A(g6537), .B(n7344), .S0(n4857), .Y(n7345));
MX2X1    g2701(.A(g6533), .B(n7345), .S0(g35), .Y(n2333));
NOR4X1   g2702(.A(g5517), .B(g5523), .C(g5511), .D(n5899_1), .Y(n7347_1));
MX2X1    g2703(.A(g5543), .B(n5592_1), .S0(n7347_1), .Y(n7348));
MX2X1    g2704(.A(g5535), .B(n7348), .S0(g35), .Y(n2338));
INVX1    g2705(.A(g3736), .Y(n7350));
INVX1    g2706(.A(g3719), .Y(n7351));
INVX1    g2707(.A(g3752), .Y(n7352_1));
INVX1    g2708(.A(g3706), .Y(n7353));
INVX1    g2709(.A(g3723), .Y(n7354));
NOR4X1   g2710(.A(n7353), .B(n7352_1), .C(n7351), .D(n7354), .Y(n7355));
NAND3X1  g2711(.A(n7355), .B(g3727), .C(g3731), .Y(n7356));
INVX1    g2712(.A(g3731), .Y(n7357_1));
INVX1    g2713(.A(g3727), .Y(n7358));
INVX1    g2714(.A(g3712), .Y(n7359));
NOR4X1   g2715(.A(g3706), .B(g3719), .C(n7359), .D(g3723), .Y(n7360));
NAND3X1  g2716(.A(n7360), .B(n7358), .C(n7357_1), .Y(n7361));
AND2X1   g2717(.A(n7361), .B(n7356), .Y(n7362_1));
NOR2X1   g2718(.A(g3747), .B(n7352_1), .Y(n7363));
INVX1    g2719(.A(g3742), .Y(n7364));
NOR3X1   g2720(.A(n7364), .B(n7350), .C(g84), .Y(n7365));
NOR3X1   g2721(.A(n7357_1), .B(n7350), .C(n5495), .Y(n7366));
OAI21X1  g2722(.A0(n7366), .A1(n7365), .B0(n7363), .Y(n7367_1));
AND2X1   g2723(.A(g3747), .B(g3712), .Y(n7368));
NAND4X1  g2724(.A(n7357_1), .B(n7350), .C(g84), .D(n7368), .Y(n7369));
NAND4X1  g2725(.A(n7364), .B(n7350), .C(n5495), .D(n7368), .Y(n7370));
NAND3X1  g2726(.A(n7370), .B(n7369), .C(n7367_1), .Y(n7371));
NOR2X1   g2727(.A(n7371), .B(n7350), .Y(n7372_1));
MX2X1    g2728(.A(n7350), .B(n7372_1), .S0(n7362_1), .Y(n7373));
MX2X1    g2729(.A(g3731), .B(n7373), .S0(g35), .Y(n2347));
INVX1    g2730(.A(g5857), .Y(n7375));
NOR4X1   g2731(.A(n6653_1), .B(n4862), .C(n4860), .D(n7375), .Y(n7376));
MX2X1    g2732(.A(g5961), .B(n5592_1), .S0(n7376), .Y(n7377_1));
MX2X1    g2733(.A(g5945), .B(n7377_1), .S0(g35), .Y(n2352));
OR2X1    g2734(.A(g6227), .B(g6219), .Y(n7379));
NOR2X1   g2735(.A(n7379), .B(n4872), .Y(n7380));
MX2X1    g2736(.A(g6243), .B(n5592_1), .S0(n7380), .Y(n7381));
MX2X1    g2737(.A(g6295), .B(n7381), .S0(g35), .Y(n2357));
AOI21X1  g2738(.A0(g640), .A1(n6133), .B0(n5292), .Y(n7383));
NAND4X1  g2739(.A(n6287), .B(n6285), .C(n6284), .D(n7383), .Y(n7384));
AOI21X1  g2740(.A0(g640), .A1(n6133), .B0(n5222), .Y(n7385));
MX2X1    g2741(.A(n5222), .B(n7385), .S0(n7384), .Y(n7386));
MX2X1    g2742(.A(g626), .B(n7386), .S0(g35), .Y(n2362));
MX2X1    g2743(.A(g1211), .B(g102), .S0(g35), .Y(n2367));
NOR4X1   g2744(.A(g3857), .B(g3863), .C(g3869), .D(n7042_1), .Y(n7389));
MX2X1    g2745(.A(g3889), .B(n5592_1), .S0(n7389), .Y(n7390));
MX2X1    g2746(.A(g3881), .B(n7390), .S0(g35), .Y(n2372));
INVX1    g2747(.A(n5930), .Y(n7392_1));
NOR2X1   g2748(.A(n5975), .B(n7392_1), .Y(n7393));
MX2X1    g2749(.A(g3476), .B(g3470), .S0(n7393), .Y(n7394));
MX2X1    g2750(.A(g3470), .B(n7394), .S0(g35), .Y(n2377));
NOR4X1   g2751(.A(n5787_1), .B(n6466), .C(n4922), .D(n6501), .Y(n7396));
INVX1    g2752(.A(g1657), .Y(n7397_1));
NOR2X1   g2753(.A(g1648), .B(n7397_1), .Y(n7398));
XOR2X1   g2754(.A(n7398), .B(g110), .Y(n7399));
MX2X1    g2755(.A(g1664), .B(n7399), .S0(n7396), .Y(n7400));
MX2X1    g2756(.A(g1648), .B(n7400), .S0(g35), .Y(n2382));
MX2X1    g2757(.A(g1242), .B(g1227), .S0(g35), .Y(n2387));
XOR2X1   g2758(.A(g6120), .B(g6128), .Y(n7403));
MX2X1    g2759(.A(g6120), .B(n7403), .S0(g35), .Y(n2392));
NOR4X1   g2760(.A(g6573), .B(n7204), .C(g6549), .D(n4855), .Y(n7405));
MX2X1    g2761(.A(g6629), .B(n5592_1), .S0(n7405), .Y(n7406));
MX2X1    g2762(.A(g6613), .B(n7406), .S0(g35), .Y(n2397));
NOR3X1   g2763(.A(g896), .B(n4882), .C(g862), .Y(n7408));
MX2X1    g2764(.A(g246), .B(g887), .S0(n7408), .Y(n7409));
MX2X1    g2765(.A(g269), .B(n7409), .S0(g35), .Y(n2402));
INVX1    g2766(.A(g4040), .Y(n7411));
NOR4X1   g2767(.A(n5557), .B(n5556), .C(n7411), .D(n5558), .Y(n7412_1));
AOI21X1  g2768(.A0(n7412_1), .A1(g35), .B0(n6858), .Y(n2407));
OR2X1    g2769(.A(g4438), .B(g4443), .Y(n7414));
NOR4X1   g2770(.A(g4446), .B(g4452), .C(g4449), .D(n7414), .Y(n7415));
AND2X1   g2771(.A(g4438), .B(g4382), .Y(n7416));
MX2X1    g2772(.A(n7416), .B(g4392), .S0(n7415), .Y(n7417_1));
MX2X1    g2773(.A(g4438), .B(n7417_1), .S0(g35), .Y(n2412));
MX2X1    g2774(.A(g4308), .B(n6697), .S0(g35), .Y(n2417));
AOI22X1  g2775(.A0(g4681), .A1(g4831), .B0(g128), .B1(g4646), .Y(n7420));
INVX1    g2776(.A(n7420), .Y(n7421));
OAI22X1  g2777(.A0(n4967), .A1(g4826), .B0(n7014), .B1(g4821), .Y(n7422_1));
NOR4X1   g2778(.A(g4681), .B(g4688), .C(g4674), .D(g4646), .Y(n7423));
INVX1    g2779(.A(n7423), .Y(n7424));
OAI21X1  g2780(.A0(n7422_1), .A1(n7421), .B0(n7424), .Y(n7425));
INVX1    g2781(.A(n4721), .Y(n7426));
INVX1    g2782(.A(n4822_1), .Y(n7427_1));
NOR2X1   g2783(.A(g4785), .B(n4815), .Y(n7428));
AOI22X1  g2784(.A0(n4812_1), .A1(g4722), .B0(g4732), .B1(n7428), .Y(n7429));
AOI22X1  g2785(.A0(n6720), .A1(g4717), .B0(g4727), .B1(n4820), .Y(n7430));
AND2X1   g2786(.A(n7430), .B(n7429), .Y(n7431));
XOR2X1   g2787(.A(n7431), .B(n7427_1), .Y(n7432_1));
NAND2X1  g2788(.A(g4793), .B(g4801), .Y(n7433));
OR2X1    g2789(.A(g4801), .B(g4776), .Y(n7434));
OAI22X1  g2790(.A0(n7433), .A1(g4776), .B0(n4969_1), .B1(n7434), .Y(n7435));
INVX1    g2791(.A(g4737), .Y(n7436));
XOR2X1   g2792(.A(g4785), .B(g4709), .Y(n7437_1));
AOI21X1  g2793(.A0(n4820), .A1(n7436), .B0(n7437_1), .Y(n7438));
OR4X1    g2794(.A(g4793), .B(g4801), .C(g4776), .D(n7438), .Y(n7439));
NAND2X1  g2795(.A(n7439), .B(n7030), .Y(n7440));
AOI21X1  g2796(.A0(n7435), .A1(n7427_1), .B0(n7440), .Y(n7441));
OAI21X1  g2797(.A0(n7432_1), .A1(n7426), .B0(n7441), .Y(n7442_1));
NAND2X1  g2798(.A(n7442_1), .B(n7423), .Y(n7443));
AOI21X1  g2799(.A0(n7443), .A1(n7425), .B0(n4620), .Y(n7656));
INVX1    g2800(.A(g59), .Y(n7445));
NOR2X1   g2801(.A(n7445), .B(g35), .Y(n7446));
OR2X1    g2802(.A(n7446), .B(n7656), .Y(n2422));
XOR2X1   g2803(.A(n6690_1), .B(n4829), .Y(n7448));
NAND2X1  g2804(.A(n7448), .B(g4169), .Y(n7449));
MX2X1    g2805(.A(g4093), .B(n7449), .S0(g35), .Y(n2427));
NAND3X1  g2806(.A(n7445), .B(g73), .C(n4950), .Y(n7451));
MX2X1    g2807(.A(g4495), .B(n7451), .S0(g4581), .Y(n7452_1));
MX2X1    g2808(.A(g4495), .B(n7452_1), .S0(g35), .Y(n2432));
OAI21X1  g2809(.A0(g686), .A1(n5876), .B0(n5142), .Y(n7454));
NOR2X1   g2810(.A(n7454), .B(n5878), .Y(n7455));
INVX1    g2811(.A(g686), .Y(n7456));
AOI21X1  g2812(.A0(n7456), .A1(g667), .B0(n5142), .Y(n7457_1));
MX2X1    g2813(.A(n7455), .B(n7457_1), .S0(n5882), .Y(n7458));
MX2X1    g2814(.A(g518), .B(n7458), .S0(g35), .Y(n2437));
XOR2X1   g2815(.A(g5428), .B(g5436), .Y(n7460));
MX2X1    g2816(.A(g5428), .B(n7460), .S0(g35), .Y(n2442));
MX2X1    g2817(.A(g3139), .B(g3133), .S0(n4846_1), .Y(n7462_1));
MX2X1    g2818(.A(g3133), .B(n7462_1), .S0(g35), .Y(n2452));
NAND2X1  g2819(.A(g246), .B(n4950), .Y(n7464));
AOI21X1  g2820(.A0(g239), .A1(g72), .B0(g73), .Y(n7465));
AND2X1   g2821(.A(n7465), .B(n7464), .Y(n7466));
NOR2X1   g2822(.A(n6106), .B(g72), .Y(n7467_1));
OAI21X1  g2823(.A0(n6105_1), .A1(n4950), .B0(g73), .Y(n7468));
OAI21X1  g2824(.A0(n7468), .A1(n7467_1), .B0(g35), .Y(n7469));
OAI22X1  g2825(.A0(n7466), .A1(n7469), .B0(n4883), .B1(g35), .Y(n2457));
INVX1    g2826(.A(n6020_1), .Y(n7471));
OAI21X1  g2827(.A0(n6021), .A1(n7471), .B0(g4584), .Y(n7472_1));
NAND4X1  g2828(.A(g4322), .B(n5714), .C(g4332), .D(n6020_1), .Y(n7473));
AOI21X1  g2829(.A0(n7473), .A1(n7472_1), .B0(n6023), .Y(n7474));
MX2X1    g2830(.A(g4332), .B(n7474), .S0(g35), .Y(n2462));
INVX1    g2831(.A(g142), .Y(n7476));
NOR4X1   g2832(.A(n5661), .B(n5516_1), .C(n7476), .D(n6113), .Y(n7477_1));
MX2X1    g2833(.A(n7476), .B(n7477_1), .S0(n7049), .Y(n7478));
MX2X1    g2834(.A(g298), .B(n7478), .S0(g35), .Y(n2467));
INVX1    g2835(.A(g5821), .Y(n7480));
XOR2X1   g2836(.A(n7480), .B(g5827), .Y(n7481_1));
MX2X1    g2837(.A(g5831), .B(n7481_1), .S0(n6749), .Y(n7482));
MX2X1    g2838(.A(g5827), .B(n7482), .S0(g35), .Y(n2476));
MX2X1    g2839(.A(g239), .B(g881), .S0(n7408), .Y(n7484));
MX2X1    g2840(.A(g262), .B(n7484), .S0(g35), .Y(n2481));
NAND4X1  g2841(.A(g1221), .B(g1087), .C(g1205), .D(g1211), .Y(n7486_1));
INVX1    g2842(.A(n7486_1), .Y(n7487));
NAND3X1  g2843(.A(g1221), .B(g1087), .C(g1205), .Y(n7488));
OR2X1    g2844(.A(n7488), .B(g1216), .Y(n7489));
NAND2X1  g2845(.A(n7488), .B(g1216), .Y(n7490));
AOI21X1  g2846(.A0(n7490), .A1(n7489), .B0(n7487), .Y(n7491_1));
MX2X1    g2847(.A(g1221), .B(n7491_1), .S0(g35), .Y(n2486));
NOR2X1   g2848(.A(n5217), .B(n5616), .Y(n7493));
OAI21X1  g2849(.A0(n6169), .A1(g2848), .B0(g35), .Y(n7494));
AOI21X1  g2850(.A0(n7493), .A1(n3747), .B0(n7494), .Y(n7495));
AND2X1   g2851(.A(g94), .B(n4620), .Y(n7496_1));
OR2X1    g2852(.A(n7496_1), .B(n7495), .Y(n2491));
INVX1    g2853(.A(g5112), .Y(n7498));
AOI21X1  g2854(.A0(n7498), .A1(g5105), .B0(g5022), .Y(n7499));
OR2X1    g2855(.A(g5101), .B(n4620), .Y(n7500));
OAI22X1  g2856(.A0(n7499), .A1(n7500), .B0(n7498), .B1(g35), .Y(n2501));
NOR2X1   g2857(.A(n6055), .B(g1002), .Y(n7502));
OR4X1    g2858(.A(n7502), .B(n6057), .C(n6056), .D(n6058_1), .Y(n7503));
MX2X1    g2859(.A(n6328), .B(g1030), .S0(n7503), .Y(n7504));
MX2X1    g2860(.A(g1024), .B(n7504), .S0(g35), .Y(n2511));
OR2X1    g2861(.A(g3171), .B(g3179), .Y(n7506_1));
NOR3X1   g2862(.A(n7506_1), .B(n5593), .C(g3155), .Y(n7507));
MX2X1    g2863(.A(g3231), .B(n5592_1), .S0(n7507), .Y(n7508));
MX2X1    g2864(.A(g3215), .B(n7508), .S0(g35), .Y(n2521));
MX2X1    g2865(.A(g6444), .B(g6727), .S0(g35), .Y(n2526));
AND2X1   g2866(.A(n6707), .B(n6702), .Y(n7511_1));
INVX1    g2867(.A(n7511_1), .Y(n7512));
INVX1    g2868(.A(g1589), .Y(n7513));
NOR2X1   g2869(.A(n6700), .B(n5524), .Y(n7514));
MX2X1    g2870(.A(n7514), .B(n7513), .S0(n6702), .Y(n7515_1));
OAI21X1  g2871(.A0(g2227), .A1(g2153), .B0(g2241), .Y(n7516));
XOR2X1   g2872(.A(n7516), .B(n7515_1), .Y(n7517));
MX2X1    g2873(.A(g2241), .B(n7517), .S0(n7512), .Y(n7518));
MX2X1    g2874(.A(g2227), .B(n7518), .S0(g35), .Y(n2540));
AND2X1   g2875(.A(g1548), .B(g1430), .Y(n7520_1));
XOR2X1   g2876(.A(n7520_1), .B(g1564), .Y(n7521));
MX2X1    g2877(.A(g1548), .B(n7521), .S0(g35), .Y(n2545));
MX2X1    g2878(.A(g5752), .B(g6035), .S0(g35), .Y(n2550));
INVX1    g2879(.A(g6549), .Y(n7524));
NOR4X1   g2880(.A(n4854), .B(n7204), .C(n7524), .D(g6565), .Y(n7525_1));
MX2X1    g2881(.A(g6649), .B(n5592_1), .S0(n7525_1), .Y(n7526));
MX2X1    g2882(.A(g6633), .B(n7526), .S0(g35), .Y(n2559));
NAND2X1  g2883(.A(n4946), .B(n4928), .Y(n7528));
OAI21X1  g2884(.A0(n4947), .A1(n4928), .B0(n7528), .Y(n2564));
MX2X1    g2885(.A(n7356), .B(n7361), .S0(n7350), .Y(n7530_1));
NOR2X1   g2886(.A(n7371), .B(n7364), .Y(n7531));
MX2X1    g2887(.A(n7364), .B(n7531), .S0(n7530_1), .Y(n7532));
MX2X1    g2888(.A(g3736), .B(n7532), .S0(g35), .Y(n2574));
MX2X1    g2889(.A(g225), .B(g859), .S0(n7408), .Y(n7534));
MX2X1    g2890(.A(g872), .B(n7534), .S0(g35), .Y(n2579));
MX2X1    g2891(.A(g4483), .B(g6748), .S0(g35), .Y(n2584));
NAND3X1  g2892(.A(n7445), .B(n4953), .C(g72), .Y(n7537));
MX2X1    g2893(.A(g4501), .B(n7537), .S0(g4581), .Y(n7538));
MX2X1    g2894(.A(g4501), .B(n7538), .S0(g35), .Y(n2589));
NOR3X1   g2895(.A(n5645_1), .B(n4858), .C(g4087), .Y(n7540_1));
NAND2X1  g2896(.A(g5869), .B(n4860), .Y(n7541));
NAND2X1  g2897(.A(n4861_1), .B(g5873), .Y(n7542));
AOI21X1  g2898(.A0(n7542), .A1(n7541), .B0(n7540_1), .Y(n7543));
MX2X1    g2899(.A(g5869), .B(n7543), .S0(g35), .Y(n2594));
INVX1    g2900(.A(n5483), .Y(n7545_1));
INVX1    g2901(.A(n5489), .Y(n7546));
NAND3X1  g2902(.A(n7546), .B(n7545_1), .C(g5037), .Y(n7547));
OAI21X1  g2903(.A0(n5489), .A1(n5483), .B0(n5486), .Y(n7548));
OAI21X1  g2904(.A0(n7547), .A1(n5501), .B0(n7548), .Y(n7549));
MX2X1    g2905(.A(g5033), .B(n7549), .S0(g35), .Y(n2599));
INVX1    g2906(.A(g2342), .Y(n7551));
OAI21X1  g2907(.A0(g2319), .A1(n7551), .B0(n4932), .Y(n7552));
OAI21X1  g2908(.A0(n6204), .A1(n4918), .B0(n7552), .Y(n7553));
MX2X1    g2909(.A(g2319), .B(n7553), .S0(n7227), .Y(n7554));
MX2X1    g2910(.A(g2327), .B(n7554), .S0(g35), .Y(n2604));
MX2X1    g2911(.A(g5495), .B(g5489), .S0(n4869), .Y(n7556));
MX2X1    g2912(.A(g5489), .B(n7556), .S0(g35), .Y(n2609));
MX2X1    g2913(.A(g4145), .B(g4164), .S0(g4253), .Y(n7558));
INVX1    g2914(.A(n7558), .Y(n7559));
MX2X1    g2915(.A(g4180), .B(n7559), .S0(g35), .Y(n2614));
NOR3X1   g2916(.A(g5170), .B(g5176), .C(g5164), .Y(n7561));
NAND3X1  g2917(.A(n7561), .B(g5188), .C(n4642_1), .Y(n7562));
MX2X1    g2918(.A(n5592_1), .B(g5208), .S0(n7562), .Y(n7563));
MX2X1    g2919(.A(g5212), .B(n7563), .S0(g35), .Y(n2619));
AND2X1   g2920(.A(g2151), .B(n4620), .Y(n2624));
NOR4X1   g2921(.A(g5527), .B(n4867), .C(n5854), .D(g5517), .Y(n7566));
MX2X1    g2922(.A(g5579), .B(n5592_1), .S0(n7566), .Y(n7567));
MX2X1    g2923(.A(g5555), .B(n7567), .S0(g35), .Y(n2629));
NOR4X1   g2924(.A(n7375), .B(n6653_1), .C(g5869), .D(n7540_1), .Y(n7569));
MX2X1    g2925(.A(g5863), .B(n7569), .S0(g35), .Y(n2634));
MX2X1    g2926(.A(g5712), .B(g5752), .S0(g5706), .Y(n7571));
OR2X1    g2927(.A(n7571), .B(n7057), .Y(n7572));
NAND2X1  g2928(.A(n7571), .B(n7057), .Y(n7573));
OAI21X1  g2929(.A0(n7572), .A1(n7077), .B0(n7573), .Y(n7574));
MX2X1    g2930(.A(g5706), .B(n7574), .S0(g35), .Y(n2639));
MX2X1    g2931(.A(g1585), .B(g1570), .S0(g35), .Y(n2644));
INVX1    g2932(.A(g5802), .Y(n7577));
AOI21X1  g2933(.A0(n7577), .A1(g5794), .B0(g5752), .Y(n7578));
OR2X1    g2934(.A(g5798), .B(n4620), .Y(n7579));
OAI22X1  g2935(.A0(n7578), .A1(n7579), .B0(n7577), .B1(g35), .Y(n2649));
NOR3X1   g2936(.A(n7379), .B(g6203), .C(n5980), .Y(n7581));
MX2X1    g2937(.A(g6279), .B(n5592_1), .S0(n7581), .Y(n7582));
MX2X1    g2938(.A(g6263), .B(n7582), .S0(g35), .Y(n2654));
NOR3X1   g2939(.A(n6654), .B(n7375), .C(g5863), .Y(n7584));
MX2X1    g2940(.A(g5917), .B(n5592_1), .S0(n7584), .Y(n7585_1));
MX2X1    g2941(.A(g5889), .B(n7585_1), .S0(g35), .Y(n2659));
NOR4X1   g2942(.A(n4995), .B(n5616), .C(g28), .D(n4997_1), .Y(n7587));
AND2X1   g2943(.A(n7587), .B(n4586), .Y(n7588));
AOI21X1  g2944(.A0(g1306), .A1(g962), .B0(n4620), .Y(n7589));
OAI21X1  g2945(.A0(n7589), .A1(g2975), .B0(g35), .Y(n7590_1));
NAND2X1  g2946(.A(g2965), .B(n4620), .Y(n7591));
OAI21X1  g2947(.A0(n7590_1), .A1(n7588), .B0(n7591), .Y(n2664));
XOR2X1   g2948(.A(n4874), .B(g6167), .Y(n7593));
MX2X1    g2949(.A(g6163), .B(n7593), .S0(g35), .Y(n2669));
INVX1    g2950(.A(g2599), .Y(n7595_1));
INVX1    g2951(.A(n6003), .Y(n7596));
NAND4X1  g2952(.A(n5637), .B(g112), .C(n4824), .D(n5140_1), .Y(n7597));
NAND3X1  g2953(.A(n7597), .B(n7596), .C(g2555), .Y(n7598));
OAI21X1  g2954(.A0(n7596), .A1(n7595_1), .B0(n7598), .Y(n7599));
MX2X1    g2955(.A(g2606), .B(n7599), .S0(g35), .Y(n2678));
NAND2X1  g2956(.A(n5549), .B(g1526), .Y(n7601));
INVX1    g2957(.A(g1495), .Y(n7602));
NAND2X1  g2958(.A(g1442), .B(n7602), .Y(n7603));
NOR3X1   g2959(.A(n7603), .B(n7601), .C(n6513), .Y(n7604));
XOR2X1   g2960(.A(g1448), .B(g1454), .Y(n7605_1));
MX2X1    g2961(.A(g1448), .B(n7605_1), .S0(n7604), .Y(n7606));
MX2X1    g2962(.A(g1454), .B(n7606), .S0(g35), .Y(n2683));
INVX1    g2963(.A(g3805), .Y(n7608));
AOI21X1  g2964(.A0(g3798), .A1(n7608), .B0(g3712), .Y(n7609_1));
OR2X1    g2965(.A(g3794), .B(n4620), .Y(n7610));
OAI22X1  g2966(.A0(n7609_1), .A1(n7610), .B0(n7608), .B1(g35), .Y(n2691));
NAND3X1  g2967(.A(n4932), .B(g2307), .C(n7228), .Y(n7612));
NAND3X1  g2968(.A(n7228), .B(g2342), .C(g2295), .Y(n7613_1));
AND2X1   g2969(.A(n7613_1), .B(n7612), .Y(n7614));
AND2X1   g2970(.A(g2351), .B(g2319), .Y(n7615));
NOR2X1   g2971(.A(n4932), .B(g2342), .Y(n7616));
AOI22X1  g2972(.A0(n7615), .A1(g2299), .B0(g2303), .B1(n7616), .Y(n7617_1));
NAND3X1  g2973(.A(n4932), .B(g2315), .C(g2342), .Y(n7618));
NAND3X1  g2974(.A(g2311), .B(g2319), .C(n7551), .Y(n7619));
NAND4X1  g2975(.A(n7618), .B(n7617_1), .C(n7614), .D(n7619), .Y(n7620));
MX2X1    g2976(.A(g2370), .B(n7620), .S0(n7227), .Y(n7621));
MX2X1    g2977(.A(g2351), .B(n7621), .S0(g35), .Y(n2696));
NOR4X1   g2978(.A(g5176), .B(g5164), .C(n4620), .D(n6042), .Y(n2701));
MX2X1    g2979(.A(n7308), .B(n7307), .S0(n7306_1), .Y(n7624));
MX2X1    g2980(.A(g150), .B(n7624), .S0(g35), .Y(n2710));
NOR3X1   g2981(.A(n5645_1), .B(n4841_1), .C(g4087), .Y(n7626));
NOR4X1   g2982(.A(g6561), .B(g6549), .C(n4620), .D(n7626), .Y(n2715));
NOR2X1   g2983(.A(n6474), .B(n6689), .Y(n7628));
XOR2X1   g2984(.A(n7628), .B(n4840), .Y(n7629));
NAND2X1  g2985(.A(g4169), .B(g35), .Y(n7630));
OAI22X1  g2986(.A0(n7629), .A1(n7630), .B0(n6689), .B1(g35), .Y(n2720));
NOR4X1   g2987(.A(n4967), .B(n4969_1), .C(g4801), .D(n4723), .Y(n7632_1));
AOI21X1  g2988(.A0(n4968), .A1(g4793), .B0(n6011), .Y(n7633));
OAI21X1  g2989(.A0(n7633), .A1(n7632_1), .B0(n6010_1), .Y(n7634));
NAND2X1  g2990(.A(g4793), .B(n4620), .Y(n7635));
OAI21X1  g2991(.A0(n7634), .A1(n4620), .B0(n7635), .Y(n2725));
NOR3X1   g2992(.A(g54), .B(g56), .C(g53), .Y(n7637));
AOI21X1  g2993(.A0(n7637), .A1(n5962), .B0(g2984), .Y(n7638));
NAND2X1  g2994(.A(n6674), .B(n3220), .Y(n7639));
NAND2X1  g2995(.A(n7639), .B(g35), .Y(n7640));
OAI22X1  g2996(.A0(n7638), .A1(n7640), .B0(n5428), .B1(g35), .Y(n2730));
INVX1    g2997(.A(g3857), .Y(n7642));
NOR4X1   g2998(.A(n7041), .B(n4850), .C(n4848), .D(n7642), .Y(n7643));
MX2X1    g2999(.A(g3961), .B(n5592_1), .S0(n7643), .Y(n7644));
MX2X1    g3000(.A(g3945), .B(n7644), .S0(g35), .Y(n2735));
INVX1    g3001(.A(g5767), .Y(n7646_1));
NOR2X1   g3002(.A(g5763), .B(n7646_1), .Y(n7647));
NOR2X1   g3003(.A(n7646_1), .B(g5759), .Y(n7648));
MX2X1    g3004(.A(n7647), .B(n7648), .S0(g5774), .Y(n7649));
MX2X1    g3005(.A(g5767), .B(n7649), .S0(g35), .Y(n2740));
NAND3X1  g3006(.A(g1157), .B(g1183), .C(g1171), .Y(n7651_1));
MX2X1    g3007(.A(g996), .B(g962), .S0(n7651_1), .Y(n7652));
MX2X1    g3008(.A(g1178), .B(n7652), .S0(g35), .Y(n2745));
NOR2X1   g3009(.A(n4822_1), .B(n4811), .Y(n7654));
NOR3X1   g3010(.A(n4822_1), .B(n4810), .C(n4809), .Y(n7655));
OR2X1    g3011(.A(n7655), .B(n7654), .Y(n2750));
OR2X1    g3012(.A(g6565), .B(g6573), .Y(n7657));
NOR3X1   g3013(.A(n7657), .B(n7204), .C(g6549), .Y(n7658));
MX2X1    g3014(.A(g6625), .B(n5592_1), .S0(n7658), .Y(n7659));
MX2X1    g3015(.A(g6609), .B(n7659), .S0(g35), .Y(n2760));
OAI21X1  g3016(.A0(n5457), .A1(n5435_1), .B0(n5282), .Y(n7661));
OAI21X1  g3017(.A0(n5457), .A1(n5435_1), .B0(g22), .Y(n7662));
NAND2X1  g3018(.A(n7662), .B(n7661), .Y(n2765));
MX2X1    g3019(.A(n6057), .B(g1018), .S0(n6060), .Y(n7664));
MX2X1    g3020(.A(g1002), .B(n7664), .S0(g35), .Y(n2770));
NAND3X1  g3021(.A(n5986), .B(n5984), .C(n4712_1), .Y(n7666));
INVX1    g3022(.A(g1564), .Y(n7667));
INVX1    g3023(.A(g1554), .Y(n7668));
INVX1    g3024(.A(n7520_1), .Y(n7669));
NOR3X1   g3025(.A(n7669), .B(n7668), .C(n7667), .Y(n7670));
OR4X1    g3026(.A(g1418), .B(g1422), .C(n4620), .D(g1426), .Y(n7671));
AOI21X1  g3027(.A0(n7670), .A1(n7666), .B0(n7671), .Y(n2775));
NAND2X1  g3028(.A(n6864_1), .B(g35), .Y(n7673));
OAI22X1  g3029(.A0(n7412_1), .A1(n7673), .B0(n7411), .B1(g35), .Y(n2779));
INVX1    g3030(.A(g1467), .Y(n7675));
XOR2X1   g3031(.A(n6519), .B(n5303_1), .Y(n7676));
AOI21X1  g3032(.A0(n6521), .A1(n7675), .B0(n7676), .Y(n7677));
NOR3X1   g3033(.A(n5549), .B(n6000_1), .C(n6513), .Y(n7678));
MX2X1    g3034(.A(g1467), .B(n7677), .S0(n7678), .Y(n7679));
MX2X1    g3035(.A(g1448), .B(n7679), .S0(g35), .Y(n2784));
INVX1    g3036(.A(g2421), .Y(n7681));
NAND2X1  g3037(.A(n7681), .B(g2465), .Y(n7682));
NOR4X1   g3038(.A(n5567), .B(n6445), .C(g2485), .D(n5569), .Y(n7683));
MX2X1    g3039(.A(g2461), .B(n7682), .S0(n7683), .Y(n7684));
MX2X1    g3040(.A(g2441), .B(n7684), .S0(g35), .Y(n2789));
OAI21X1  g3041(.A0(g5752), .A1(g5712), .B0(n7059), .Y(n7686));
NAND3X1  g3042(.A(g5706), .B(n7058), .C(n7065_1), .Y(n7687));
OAI21X1  g3043(.A0(n7686), .A1(n7077), .B0(n7687), .Y(n7688));
MX2X1    g3044(.A(g5712), .B(n7688), .S0(g35), .Y(n2794));
MX2X1    g3045(.A(g457), .B(g452), .S0(n5601), .Y(n7690));
MX2X1    g3046(.A(g452), .B(n7690), .S0(g35), .Y(n2799));
NAND4X1  g3047(.A(g2719), .B(g2729), .C(g2724), .D(g2715), .Y(n7692));
NOR4X1   g3048(.A(n5508), .B(n4909), .C(n4915_1), .D(n7692), .Y(n7693));
XOR2X1   g3049(.A(n7693), .B(n4910_1), .Y(n7694));
NAND2X1  g3050(.A(n7694), .B(g2841), .Y(n7695));
MX2X1    g3051(.A(g2748), .B(n7695), .S0(g35), .Y(n2804));
INVX1    g3052(.A(g93), .Y(n7697));
NAND3X1  g3053(.A(n4957), .B(g4358), .C(n5174), .Y(n7698));
OR4X1    g3054(.A(n6466), .B(n7698), .C(n7697), .D(n6747_1), .Y(n7699));
NOR3X1   g3055(.A(n6747_1), .B(n6951), .C(g5990), .Y(n7700));
AOI21X1  g3056(.A0(n6746), .A1(g6049), .B0(n6944), .Y(n7701));
OAI21X1  g3057(.A0(n7701), .A1(n7700), .B0(n7699), .Y(n7702));
NAND2X1  g3058(.A(g6049), .B(n4620), .Y(n7703));
OAI21X1  g3059(.A0(n7702), .A1(n4620), .B0(n7703), .Y(n2809));
MX2X1    g3060(.A(g471), .B(g269), .S0(n5601), .Y(n7705));
MX2X1    g3061(.A(g457), .B(n7705), .S0(g35), .Y(n2814));
INVX1    g3062(.A(g1256), .Y(n7707));
INVX1    g3063(.A(g1252), .Y(n7708));
NAND4X1  g3064(.A(g1280), .B(g1266), .C(g1249), .D(g1570), .Y(n7709));
NOR2X1   g3065(.A(n7709), .B(n7708), .Y(n7710));
AND2X1   g3066(.A(g1570), .B(g1256), .Y(n7711));
MX2X1    g3067(.A(n7711), .B(n7707), .S0(n7710), .Y(n7712));
MX2X1    g3068(.A(g1252), .B(n7712), .S0(g35), .Y(n2819));
MX2X1    g3069(.A(g5022), .B(g5062), .S0(g5016), .Y(n7714));
OR2X1    g3070(.A(n7714), .B(n5479), .Y(n7715));
NAND2X1  g3071(.A(n7714), .B(n5479), .Y(n7716));
OAI21X1  g3072(.A0(n7715), .A1(n5501), .B0(n7716), .Y(n7717));
MX2X1    g3073(.A(g5016), .B(n7717), .S0(g35), .Y(n2824));
INVX1    g3074(.A(g4888), .Y(n7719));
NOR4X1   g3075(.A(g4975), .B(g4899), .C(n7719), .D(n4960), .Y(n7720));
AOI21X1  g3076(.A0(n7720), .A1(n5928), .B0(n6326_1), .Y(n7721));
INVX1    g3077(.A(n7721), .Y(n7722));
NAND4X1  g3078(.A(g6741), .B(g6682), .C(g6727), .D(g6668), .Y(n7723));
NOR2X1   g3079(.A(n7723), .B(n7722), .Y(n7724));
MX2X1    g3080(.A(g6519), .B(g6513), .S0(n7724), .Y(n7725));
MX2X1    g3081(.A(g6513), .B(n7725), .S0(g35), .Y(n2829));
NAND2X1  g3082(.A(g4165), .B(g35), .Y(n7727));
NAND2X1  g3083(.A(g4165), .B(n4620), .Y(n7728));
NAND2X1  g3084(.A(n7728), .B(n7727), .Y(n2834));
MX2X1    g3085(.A(n5623), .B(g1246), .S0(n5621), .Y(n7730));
OAI21X1  g3086(.A0(g1728), .A1(g1802), .B0(g1816), .Y(n7731));
XOR2X1   g3087(.A(n7731), .B(n7730), .Y(n7732));
MX2X1    g3088(.A(g1816), .B(n7732), .S0(n5636), .Y(n7733));
MX2X1    g3089(.A(g1802), .B(n7733), .S0(g35), .Y(n2839));
MX2X1    g3090(.A(g4459), .B(g4473), .S0(g35), .Y(n2844));
XOR2X1   g3091(.A(n6607), .B(g3436), .Y(n7736));
MX2X1    g3092(.A(g3431), .B(n7736), .S0(g35), .Y(n2849));
AND2X1   g3093(.A(g5782), .B(g5774), .Y(n7738));
XOR2X1   g3094(.A(n7738), .B(g5787), .Y(n7739));
MX2X1    g3095(.A(g5782), .B(n7739), .S0(g35), .Y(n2854));
NOR2X1   g3096(.A(n7113_1), .B(g35), .Y(n7741));
OR2X1    g3097(.A(n7741), .B(n1787), .Y(n2859));
INVX1    g3098(.A(g4477), .Y(n7743));
OAI21X1  g3099(.A0(n4809), .A1(g4507), .B0(n5701), .Y(n7744));
NAND3X1  g3100(.A(n7744), .B(g4474), .C(n7743), .Y(n7745));
AND2X1   g3101(.A(g4462), .B(g4467), .Y(n7746));
AOI21X1  g3102(.A0(n7746), .A1(n7745), .B0(n4620), .Y(n2864));
INVX1    g3103(.A(g3821), .Y(n7748));
XOR2X1   g3104(.A(n7748), .B(g3827), .Y(n7749));
MX2X1    g3105(.A(g3831), .B(n7749), .S0(n7137_1), .Y(n7750));
MX2X1    g3106(.A(g3827), .B(n7750), .S0(g35), .Y(n2869));
MX2X1    g3107(.A(g2514), .B(g2509), .S0(n7133), .Y(n7753));
MX2X1    g3108(.A(g2509), .B(n7753), .S0(g35), .Y(n2874));
NOR4X1   g3109(.A(n4896_1), .B(g4899), .C(n4895), .D(n4960), .Y(n7755));
AOI21X1  g3110(.A0(n7755), .A1(n5928), .B0(n6491), .Y(n7756));
INVX1    g3111(.A(n7756), .Y(n7757));
OR4X1    g3112(.A(n6466), .B(n5182), .C(n7697), .D(n7757), .Y(n7758));
INVX1    g3113(.A(g3352), .Y(n7759));
NOR3X1   g3114(.A(n7757), .B(n7759), .C(g3288), .Y(n7760));
INVX1    g3115(.A(g3288), .Y(n7761));
AOI21X1  g3116(.A0(n7756), .A1(g3352), .B0(n7761), .Y(n7762));
OAI21X1  g3117(.A0(n7762), .A1(n7760), .B0(n7758), .Y(n7763));
NAND2X1  g3118(.A(g3352), .B(n4620), .Y(n7764));
OAI21X1  g3119(.A0(n7763), .A1(n4620), .B0(n7764), .Y(n2879));
INVX1    g3120(.A(g2399), .Y(n7766));
XOR2X1   g3121(.A(g2393), .B(n7766), .Y(n7767));
MX2X1    g3122(.A(g2403), .B(n7767), .S0(n5553), .Y(n7768));
MX2X1    g3123(.A(g2399), .B(n7768), .S0(g35), .Y(n2884));
MX2X1    g3124(.A(g2145), .B(n3220), .S0(n6029), .Y(n7770));
MX2X1    g3125(.A(g2138), .B(n7770), .S0(g35), .Y(n2889));
INVX1    g3126(.A(g1624), .Y(n7772));
NOR4X1   g3127(.A(n5787_1), .B(n7772), .C(n7397_1), .D(n6501), .Y(n7773));
XOR2X1   g3128(.A(n7773), .B(g1700), .Y(n7774));
MX2X1    g3129(.A(g1696), .B(n7774), .S0(g35), .Y(n2894));
AOI21X1  g3130(.A0(n7456), .A1(g667), .B0(n5136), .Y(n7776));
MX2X1    g3131(.A(g513), .B(n7776), .S0(n5880_1), .Y(n7777));
MX2X1    g3132(.A(g504), .B(n7777), .S0(g35), .Y(n2899));
NAND2X1  g3133(.A(g2837), .B(g35), .Y(n7779));
NAND2X1  g3134(.A(g2837), .B(n4620), .Y(n7780));
NAND2X1  g3135(.A(n7780), .B(n7779), .Y(n2904));
NOR3X1   g3136(.A(n7190), .B(n5179), .C(n6438), .Y(n7782));
NAND3X1  g3137(.A(g28753), .B(g5357), .C(n6333), .Y(n7783));
OAI21X1  g3138(.A0(n6438), .A1(n6340), .B0(g5297), .Y(n7784));
AOI21X1  g3139(.A0(n7784), .A1(n7783), .B0(n7782), .Y(n7785));
MX2X1    g3140(.A(g5357), .B(n7785), .S0(g35), .Y(n2909));
NAND3X1  g3141(.A(n7693), .B(g2759), .C(g2756), .Y(n7787));
XOR2X1   g3142(.A(n7787), .B(g2763), .Y(n7788));
NAND2X1  g3143(.A(n7788), .B(g2841), .Y(n7789));
MX2X1    g3144(.A(g2759), .B(n7789), .S0(g35), .Y(n2919));
NOR2X1   g3145(.A(n4968), .B(n4969_1), .Y(n7791));
NOR3X1   g3146(.A(n4723), .B(n4967), .C(g4793), .Y(n7792));
OAI21X1  g3147(.A0(n7792), .A1(n7791), .B0(n6010_1), .Y(n7793));
NAND2X1  g3148(.A(g4818), .B(n4620), .Y(n7794));
OAI21X1  g3149(.A0(n7793), .A1(n4620), .B0(n7794), .Y(n2924));
NOR2X1   g3150(.A(n6668), .B(n6316_1), .Y(n7796));
OAI21X1  g3151(.A0(g952), .A1(n4716), .B0(g35), .Y(n7797));
OAI22X1  g3152(.A0(n7796), .A1(n7797), .B0(n5245), .B1(g35), .Y(n2929));
INVX1    g3153(.A(g1263), .Y(n7799));
INVX1    g3154(.A(g1259), .Y(n7800));
NOR4X1   g3155(.A(n7800), .B(n7708), .C(n7707), .D(n7709), .Y(n7801));
AND2X1   g3156(.A(g1570), .B(g1263), .Y(n7802));
MX2X1    g3157(.A(n7802), .B(n7799), .S0(n7801), .Y(n7803));
MX2X1    g3158(.A(g1259), .B(n7803), .S0(g35), .Y(n2934));
INVX1    g3159(.A(g1246), .Y(n7805));
MX2X1    g3160(.A(n5525), .B(n7805), .S0(n5521_1), .Y(n7806));
OAI21X1  g3161(.A0(g1936), .A1(g1862), .B0(g1950), .Y(n7807));
XOR2X1   g3162(.A(n7807), .B(n7806), .Y(n7808));
MX2X1    g3163(.A(g1950), .B(n7808), .S0(n6222), .Y(n7809));
MX2X1    g3164(.A(g1936), .B(n7809), .S0(g35), .Y(n2939));
INVX1    g3165(.A(g5128), .Y(n7811));
XOR2X1   g3166(.A(n7811), .B(g5134), .Y(n7812));
MX2X1    g3167(.A(g5138), .B(n7812), .S0(n6440), .Y(n7813));
MX2X1    g3168(.A(g5134), .B(n7813), .S0(g35), .Y(n2944));
NOR3X1   g3169(.A(n5552), .B(n5154), .C(n6032), .Y(n7815));
MX2X1    g3170(.A(g2307), .B(n5547), .S0(n7815), .Y(n7816));
MX2X1    g3171(.A(g2311), .B(n7816), .S0(g35), .Y(n2949));
AND2X1   g3172(.A(n7738), .B(g5787), .Y(n7818));
XOR2X1   g3173(.A(n7818), .B(g5791), .Y(n7819));
MX2X1    g3174(.A(g5787), .B(n7819), .S0(g35), .Y(n2959));
MX2X1    g3175(.A(g3752), .B(g4040), .S0(g35), .Y(n2964));
NOR2X1   g3176(.A(n6216_1), .B(n4968), .Y(n7822));
INVX1    g3177(.A(g4664), .Y(n7823));
AND2X1   g3178(.A(g4688), .B(g4653), .Y(n7824));
AOI21X1  g3179(.A0(n7824), .A1(g4659), .B0(n7823), .Y(n7825));
INVX1    g3180(.A(g4659), .Y(n7826));
NOR4X1   g3181(.A(n4967), .B(g4664), .C(n7118_1), .D(n7826), .Y(n7827));
OAI21X1  g3182(.A0(n7827), .A1(n7825), .B0(n7822), .Y(n7828));
NAND2X1  g3183(.A(g4659), .B(n4620), .Y(n7829));
OAI21X1  g3184(.A0(n7828), .A1(n4620), .B0(n7829), .Y(n2968));
NOR4X1   g3185(.A(n5786), .B(n6466), .C(n4914), .D(n5787_1), .Y(n7831));
XOR2X1   g3186(.A(n5794), .B(g110), .Y(n7832));
MX2X1    g3187(.A(g2223), .B(n7832), .S0(n7831), .Y(n7833));
MX2X1    g3188(.A(g2208), .B(n7833), .S0(g35), .Y(n2973));
AND2X1   g3189(.A(n6748), .B(g5808), .Y(n7835));
XOR2X1   g3190(.A(n7835), .B(n6988_1), .Y(n7836));
MX2X1    g3191(.A(g5808), .B(n7836), .S0(n6746), .Y(n7837));
MX2X1    g3192(.A(g5813), .B(n7837), .S0(g35), .Y(n2978));
NOR4X1   g3193(.A(g6573), .B(n7204), .C(n7524), .D(n4855), .Y(n7839));
MX2X1    g3194(.A(g6645), .B(n5592_1), .S0(n7839), .Y(n7840));
MX2X1    g3195(.A(g6629), .B(n7840), .S0(g35), .Y(n2983));
INVX1    g3196(.A(g1996), .Y(n7842));
NOR3X1   g3197(.A(n6085), .B(n7842), .C(n5166_1), .Y(n7843));
MX2X1    g3198(.A(g2016), .B(n7037_1), .S0(n7843), .Y(n7844));
MX2X1    g3199(.A(g2020), .B(n7844), .S0(g35), .Y(n2988));
INVX1    g3200(.A(g5747), .Y(n7846));
NAND3X1  g3201(.A(n7076), .B(n7075_1), .C(g35), .Y(n7847));
OAI21X1  g3202(.A0(n7846), .A1(g35), .B0(n7847), .Y(n2993));
NOR3X1   g3203(.A(n5645_1), .B(n4831), .C(n4840), .Y(n7849));
NAND2X1  g3204(.A(g3869), .B(n4848), .Y(n7850));
NAND2X1  g3205(.A(n4849), .B(g3873), .Y(n7851));
AOI21X1  g3206(.A0(n7851), .A1(n7850), .B0(n7849), .Y(n7852));
MX2X1    g3207(.A(g3869), .B(n7852), .S0(g35), .Y(n2998));
NOR3X1   g3208(.A(n5552), .B(n5154), .C(g2331), .Y(n7854));
MX2X1    g3209(.A(g2315), .B(n5547), .S0(n7854), .Y(n7855));
MX2X1    g3210(.A(g2303), .B(n7855), .S0(g35), .Y(n3008));
INVX1    g3211(.A(g2799), .Y(n7857));
INVX1    g3212(.A(g2327), .Y(n7858));
AOI21X1  g3213(.A0(n4915_1), .A1(n4910_1), .B0(n5509), .Y(n7859));
AOI21X1  g3214(.A0(n7859), .A1(n7858), .B0(g2811), .Y(n7860));
OAI21X1  g3215(.A0(n5565), .A1(n4909), .B0(g35), .Y(n7861));
OAI22X1  g3216(.A0(n7860), .A1(n7861), .B0(n7857), .B1(g35), .Y(n3013));
NOR4X1   g3217(.A(n6653_1), .B(n4862), .C(g5873), .D(n7375), .Y(n7863));
MX2X1    g3218(.A(g5957), .B(n5592_1), .S0(n7863), .Y(n7864));
MX2X1    g3219(.A(g5941), .B(n7864), .S0(g35), .Y(n3018));
NOR4X1   g3220(.A(n6466), .B(n5145_1), .C(g504), .D(n6081), .Y(n7866));
XOR2X1   g3221(.A(n5167), .B(g112), .Y(n7867));
MX2X1    g3222(.A(g2047), .B(n7867), .S0(n7866), .Y(n7868));
MX2X1    g3223(.A(g1996), .B(n7868), .S0(g35), .Y(n3023));
NOR4X1   g3224(.A(n7642), .B(n7041), .C(g3869), .D(n7849), .Y(n7870));
MX2X1    g3225(.A(g3863), .B(n7870), .S0(g35), .Y(n3028));
MX2X1    g3226(.A(g3712), .B(g3752), .S0(g3706), .Y(n7872));
OR2X1    g3227(.A(n7872), .B(n7351), .Y(n7873));
NAND2X1  g3228(.A(n7872), .B(n7351), .Y(n7874));
OAI21X1  g3229(.A0(n7873), .A1(n7371), .B0(n7874), .Y(n7875));
MX2X1    g3230(.A(g3706), .B(n7875), .S0(g35), .Y(n3036));
NOR4X1   g3231(.A(n4868), .B(g5535), .C(n5854), .D(g5517), .Y(n7877));
MX2X1    g3232(.A(g5575), .B(n5592_1), .S0(n7877), .Y(n7878));
MX2X1    g3233(.A(g5547), .B(n7878), .S0(g35), .Y(n3041));
OR2X1    g3234(.A(n5468), .B(g22), .Y(n7880));
OR2X1    g3235(.A(n5468), .B(n5282), .Y(n7881));
NAND2X1  g3236(.A(n7881), .B(n7880), .Y(n3046));
INVX1    g3237(.A(g3802), .Y(n7883));
AOI21X1  g3238(.A0(n7883), .A1(g3794), .B0(g3752), .Y(n7884));
OR2X1    g3239(.A(g3798), .B(n4620), .Y(n7885));
OAI22X1  g3240(.A0(n7884), .A1(n7885), .B0(n7883), .B1(g35), .Y(n3051));
NOR3X1   g3241(.A(n7042_1), .B(n7642), .C(g3863), .Y(n7887));
MX2X1    g3242(.A(g3917), .B(n5592_1), .S0(n7887), .Y(n7888));
MX2X1    g3243(.A(g3889), .B(n7888), .S0(g35), .Y(n3056));
INVX1    g3244(.A(g4411), .Y(n7890));
NAND3X1  g3245(.A(n6906_1), .B(g4401), .C(g4392), .Y(n7891));
NAND2X1  g3246(.A(n7891), .B(n7890), .Y(n7892));
MX2X1    g3247(.A(g4401), .B(n7892), .S0(g35), .Y(n3071));
NOR3X1   g3248(.A(n6099), .B(n6208), .C(g6209), .Y(n7894));
MX2X1    g3249(.A(g6275), .B(n5592_1), .S0(n7894), .Y(n7895));
MX2X1    g3250(.A(g6255), .B(n7895), .S0(g35), .Y(n3076));
MX2X1    g3251(.A(g6311), .B(n5592_1), .S0(n4874), .Y(n7898));
MX2X1    g3252(.A(g6307), .B(n7898), .S0(g35), .Y(n3081));
NOR2X1   g3253(.A(n6049), .B(g1041), .Y(n7900));
OAI21X1  g3254(.A0(g979), .A1(g990), .B0(n6050), .Y(n7901));
MX2X1    g3255(.A(n7900), .B(g1041), .S0(n7901), .Y(n7902));
MX2X1    g3256(.A(g1036), .B(n7902), .S0(g35), .Y(n3091));
NAND2X1  g3257(.A(n5999), .B(g2599), .Y(n7904));
NOR3X1   g3258(.A(n5863), .B(g2619), .C(n5860_1), .Y(n7905));
MX2X1    g3259(.A(g2595), .B(n7904), .S0(n7905), .Y(n7906));
MX2X1    g3260(.A(g2575), .B(n7906), .S0(g35), .Y(n3096));
INVX1    g3261(.A(g2533), .Y(n7908));
XOR2X1   g3262(.A(g2527), .B(n7908), .Y(n7909));
MX2X1    g3263(.A(g2537), .B(n7909), .S0(n7133), .Y(n7910));
MX2X1    g3264(.A(g2533), .B(n7910), .S0(g35), .Y(n3101));
NOR2X1   g3265(.A(n5226_1), .B(n5616), .Y(n7912));
MX2X1    g3266(.A(g136), .B(n4586), .S0(n7912), .Y(n7913));
MX2X1    g3267(.A(g550), .B(n7913), .S0(g35), .Y(n3106));
INVX1    g3268(.A(g4443), .Y(n7915));
NAND3X1  g3269(.A(n7415), .B(g4392), .C(g4434), .Y(n7916));
NAND2X1  g3270(.A(n7916), .B(n7915), .Y(n7917));
MX2X1    g3271(.A(g4434), .B(n7917), .S0(g35), .Y(n3111));
MX2X1    g3272(.A(g4561), .B(g6750), .S0(g35), .Y(n3116));
MX2X1    g3273(.A(g4826), .B(n6569), .S0(n5907), .Y(n7920));
MX2X1    g3274(.A(g6311), .B(n7920), .S0(g35), .Y(n3126));
NOR3X1   g3275(.A(g6203), .B(g6209), .C(g6215), .Y(n7922));
NAND3X1  g3276(.A(n7922), .B(n4873), .C(g6219), .Y(n7923));
MX2X1    g3277(.A(n5592_1), .B(g6239), .S0(n7923), .Y(n7924));
MX2X1    g3278(.A(g6243), .B(n7924), .S0(g35), .Y(n3131));
INVX1    g3279(.A(g3767), .Y(n7926));
NOR2X1   g3280(.A(g3763), .B(n7926), .Y(n7927));
NOR2X1   g3281(.A(n7926), .B(g3759), .Y(n7928));
MX2X1    g3282(.A(n7927), .B(n7928), .S0(g3774), .Y(n7929));
MX2X1    g3283(.A(g3767), .B(n7929), .S0(g35), .Y(n3136));
MX2X1    g3284(.A(g232), .B(g875), .S0(n7408), .Y(n7931));
MX2X1    g3285(.A(g255), .B(n7931), .S0(g35), .Y(n3141));
NAND2X1  g3286(.A(g5188), .B(g5180), .Y(n7933));
NOR3X1   g3287(.A(n7933), .B(n6624), .C(n5610), .Y(n7934));
MX2X1    g3288(.A(g5268), .B(n5592_1), .S0(n7934), .Y(n7935));
MX2X1    g3289(.A(g5252), .B(n7935), .S0(g35), .Y(n3146));
MX2X1    g3290(.A(n5357), .B(n5368), .S0(n6435), .Y(n7937));
NOR2X1   g3291(.A(n7937), .B(n4620), .Y(n3151));
INVX1    g3292(.A(g2407), .Y(n7939));
XOR2X1   g3293(.A(g2413), .B(n7939), .Y(n7940));
AND2X1   g3294(.A(n7615), .B(n7227), .Y(n7941));
MX2X1    g3295(.A(g2417), .B(n7940), .S0(n7941), .Y(n7942));
MX2X1    g3296(.A(g2413), .B(n7942), .S0(g35), .Y(n3156));
NAND3X1  g3297(.A(n5638), .B(n5636), .C(g1728), .Y(n7944));
OAI21X1  g3298(.A0(n5636), .A1(n5625_1), .B0(n7944), .Y(n7945));
MX2X1    g3299(.A(g1779), .B(n7945), .S0(g35), .Y(n3161));
NOR2X1   g3300(.A(n7436), .B(g35), .Y(n3166));
OAI21X1  g3301(.A0(n5491), .A1(n5485), .B0(n5477_1), .Y(n7948));
OR4X1    g3302(.A(n5491), .B(n5485), .C(n5477_1), .D(n5501), .Y(n7949));
NAND2X1  g3303(.A(n7949), .B(n7948), .Y(n7950));
MX2X1    g3304(.A(g5046), .B(n7950), .S0(g35), .Y(n3171));
MX2X1    g3305(.A(g5406), .B(g5689), .S0(g35), .Y(n3176));
NOR3X1   g3306(.A(n5531_1), .B(g1906), .C(n5161), .Y(n7953));
MX2X1    g3307(.A(g1890), .B(n5526_1), .S0(n7953), .Y(n7954));
MX2X1    g3308(.A(g1878), .B(n7954), .S0(g35), .Y(n3181));
NAND3X1  g3309(.A(n7597), .B(n7596), .C(g2599), .Y(n7956));
OAI21X1  g3310(.A0(n7596), .A1(n5156), .B0(n7956), .Y(n7957));
MX2X1    g3311(.A(g2599), .B(n7957), .S0(g35), .Y(n3186));
MX2X1    g3312(.A(n6141_1), .B(n5410_1), .S0(n6140), .Y(n7959));
MX2X1    g3313(.A(g568), .B(n7959), .S0(g35), .Y(n3191));
MX2X1    g3314(.A(g2130), .B(n6708), .S0(n6029), .Y(n7961));
AND2X1   g3315(.A(n7961), .B(g35), .Y(n3196));
NAND2X1  g3316(.A(n6690_1), .B(g4098), .Y(n7963));
XOR2X1   g3317(.A(n7963), .B(g4108), .Y(n7964));
NAND2X1  g3318(.A(n7964), .B(g4169), .Y(n7965));
MX2X1    g3319(.A(g4098), .B(n7965), .S0(g35), .Y(n3201));
MX2X1    g3320(.A(g475), .B(g246), .S0(n5688), .Y(n7967));
MX2X1    g3321(.A(g424), .B(n7967), .S0(g35), .Y(n3210));
MX2X1    g3322(.A(g3408), .B(n5774), .S0(g35), .Y(n3225));
NAND2X1  g3323(.A(n3747), .B(n5282), .Y(n7970));
NAND2X1  g3324(.A(n3747), .B(g22), .Y(n7971));
NAND2X1  g3325(.A(n7971), .B(n7970), .Y(n3230));
MX2X1    g3326(.A(g753), .B(g64), .S0(g35), .Y(n3235));
OAI21X1  g3327(.A0(g3752), .A1(g3712), .B0(n7353), .Y(n7974));
NAND3X1  g3328(.A(g3706), .B(n7352_1), .C(n7359), .Y(n7975));
OAI21X1  g3329(.A0(n7974), .A1(n7371), .B0(n7975), .Y(n7976));
MX2X1    g3330(.A(g3712), .B(n7976), .S0(g35), .Y(n3240));
NAND3X1  g3331(.A(n6856), .B(n6865), .C(g4054), .Y(n7978));
OAI21X1  g3332(.A0(n6869), .A1(n6859_1), .B0(g3990), .Y(n7979));
AOI21X1  g3333(.A0(n7979), .A1(n7978), .B0(n7191), .Y(n7980));
MX2X1    g3334(.A(g4054), .B(n7980), .S0(g35), .Y(n3245));
INVX1    g3335(.A(g5381), .Y(n7982));
INVX1    g3336(.A(g5373), .Y(n7983));
INVX1    g3337(.A(g5377), .Y(n7984));
NOR4X1   g3338(.A(n7983), .B(n6635), .C(n6647), .D(n7984), .Y(n7985));
INVX1    g3339(.A(n7985), .Y(n7986));
NOR4X1   g3340(.A(g5377), .B(g5373), .C(g5360), .D(n6649), .Y(n7987));
INVX1    g3341(.A(n7987), .Y(n7988));
MX2X1    g3342(.A(n7986), .B(n7988), .S0(n7982), .Y(n7989));
OR2X1    g3343(.A(n7989), .B(g5385), .Y(n7990));
NAND2X1  g3344(.A(n7989), .B(g5385), .Y(n7991));
OAI21X1  g3345(.A0(n7991), .A1(n6646), .B0(n7990), .Y(n7992));
MX2X1    g3346(.A(g5381), .B(n7992), .S0(g35), .Y(n3250));
OAI21X1  g3347(.A0(n4861_1), .A1(n4860), .B0(g5881), .Y(n7994));
NAND3X1  g3348(.A(n4862), .B(g5869), .C(g5873), .Y(n7995));
AOI21X1  g3349(.A0(n7995), .A1(n7994), .B0(n7540_1), .Y(n7996));
MX2X1    g3350(.A(g5873), .B(n7996), .S0(g35), .Y(n3255));
INVX1    g3351(.A(g1982), .Y(n7998));
XOR2X1   g3352(.A(g1988), .B(n7998), .Y(n7999));
MX2X1    g3353(.A(g1992), .B(n7999), .S0(n5841_1), .Y(n8000));
MX2X1    g3354(.A(g1988), .B(n8000), .S0(g35), .Y(n3260));
INVX1    g3355(.A(n6589), .Y(n8002));
INVX1    g3356(.A(n6594), .Y(n8003));
MX2X1    g3357(.A(n8002), .B(n8003), .S0(n6592), .Y(n8004));
OR2X1    g3358(.A(n8004), .B(g3029), .Y(n8005));
NAND2X1  g3359(.A(n8004), .B(g3029), .Y(n8006));
OAI21X1  g3360(.A0(n8006), .A1(n5584), .B0(n8005), .Y(n8007));
MX2X1    g3361(.A(g3025), .B(n8007), .S0(g35), .Y(n3265));
NAND2X1  g3362(.A(n4845), .B(g3167), .Y(n8009));
NAND2X1  g3363(.A(g3171), .B(n4843), .Y(n8010));
AOI21X1  g3364(.A0(n8010), .A1(n8009), .B0(n5765), .Y(n8011));
MX2X1    g3365(.A(g3167), .B(n8011), .S0(g35), .Y(n3270));
AND2X1   g3366(.A(g3782), .B(g3774), .Y(n8013));
XOR2X1   g3367(.A(n8013), .B(g3787), .Y(n8014));
MX2X1    g3368(.A(g3782), .B(n8014), .S0(g35), .Y(n3275));
INVX1    g3369(.A(g843), .Y(n8016));
OR4X1    g3370(.A(n6247), .B(g812), .C(n8016), .D(n6246_1), .Y(n8017));
AND2X1   g3371(.A(g837), .B(g812), .Y(n8018));
OAI21X1  g3372(.A0(n6246_1), .A1(n8016), .B0(n8018), .Y(n8019));
NAND2X1  g3373(.A(n8019), .B(n8017), .Y(n8020));
MX2X1    g3374(.A(g843), .B(n8020), .S0(g35), .Y(n3280));
NOR2X1   g3375(.A(n7158), .B(g832), .Y(n8022));
NOR2X1   g3376(.A(n7158), .B(n7153), .Y(n8023));
MX2X1    g3377(.A(n8022), .B(n8023), .S0(n7154), .Y(n8024));
MX2X1    g3378(.A(g817), .B(n8024), .S0(g35), .Y(n3285));
NOR2X1   g3379(.A(n6654), .B(n4861_1), .Y(n8026));
MX2X1    g3380(.A(g5897), .B(n5592_1), .S0(n8026), .Y(n8027));
MX2X1    g3381(.A(g5949), .B(n8027), .S0(g35), .Y(n3290));
NAND2X1  g3382(.A(g4456), .B(g35), .Y(n8029));
NAND2X1  g3383(.A(g4456), .B(n4620), .Y(n8030));
NAND2X1  g3384(.A(n8030), .B(n8029), .Y(n3309));
AND2X1   g3385(.A(n7587), .B(n3747), .Y(n8032));
OR4X1    g3386(.A(g209), .B(g301), .C(g2902), .D(n5516_1), .Y(n8033));
NAND2X1  g3387(.A(n8033), .B(g35), .Y(n8034));
OAI22X1  g3388(.A0(n8032), .A1(n8034), .B0(n4783), .B1(g35), .Y(n3314));
MX2X1    g3389(.A(g311), .B(g305), .S0(g324), .Y(n8036));
NOR4X1   g3390(.A(g329), .B(g305), .C(g311), .D(g319), .Y(n8037));
AOI21X1  g3391(.A0(n8036), .A1(g319), .B0(n8037), .Y(n8038));
INVX1    g3392(.A(g336), .Y(n8039));
NAND3X1  g3393(.A(n8036), .B(n8039), .C(g311), .Y(n8040));
NAND3X1  g3394(.A(n8036), .B(g305), .C(g336), .Y(n8041));
NAND3X1  g3395(.A(n8041), .B(n8040), .C(n8038), .Y(n8042));
MX2X1    g3396(.A(g329), .B(n8042), .S0(g35), .Y(n3319));
MX2X1    g3397(.A(g168), .B(g174), .S0(n5601), .Y(n8044));
MX2X1    g3398(.A(g174), .B(n8044), .S0(g35), .Y(n3324));
INVX1    g3399(.A(g2461), .Y(n8046));
AOI21X1  g3400(.A0(n7859), .A1(n8046), .B0(g2823), .Y(n8047));
OAI22X1  g3401(.A0(n7861), .A1(n8047), .B0(n7178), .B1(g35), .Y(n3329));
MX2X1    g3402(.A(g3684), .B(n5974), .S0(n5930), .Y(n8049));
MX2X1    g3403(.A(g3614), .B(n8049), .S0(g35), .Y(n3334));
OR4X1    g3404(.A(n6466), .B(n5175), .C(n7697), .D(n7392_1), .Y(n8051));
NOR3X1   g3405(.A(n7392_1), .B(n5937), .C(g3639), .Y(n8052));
AOI21X1  g3406(.A0(n5930), .A1(g3703), .B0(n5931), .Y(n8053));
OAI21X1  g3407(.A0(n8053), .A1(n8052), .B0(n8051), .Y(n8054));
NAND2X1  g3408(.A(g3703), .B(n4620), .Y(n8055));
OAI21X1  g3409(.A0(n8054), .A1(n4620), .B0(n8055), .Y(n3339));
NOR3X1   g3410(.A(n6827), .B(n6826), .C(n6825_1), .Y(n8057));
XOR2X1   g3411(.A(n8057), .B(g3338), .Y(n8058));
MX2X1    g3412(.A(g3329), .B(n8058), .S0(g35), .Y(n3348));
INVX1    g3413(.A(g5456), .Y(n8060));
AOI21X1  g3414(.A0(n8060), .A1(g5448), .B0(g5406), .Y(n8061));
OR2X1    g3415(.A(g5452), .B(n4620), .Y(n8062));
OAI22X1  g3416(.A0(n8061), .A1(n8062), .B0(n8060), .B1(g35), .Y(n3353));
AND2X1   g3417(.A(n8013), .B(g3787), .Y(n8064));
XOR2X1   g3418(.A(n8064), .B(g3791), .Y(n8065));
MX2X1    g3419(.A(g3787), .B(n8065), .S0(g35), .Y(n3358));
MX2X1    g3420(.A(g269), .B(g884), .S0(n7408), .Y(n8067));
MX2X1    g3421(.A(g239), .B(n8067), .S0(g35), .Y(n3363));
MX2X1    g3422(.A(g401), .B(g429), .S0(n5688), .Y(n8069));
MX2X1    g3423(.A(g429), .B(n8069), .S0(g35), .Y(n3368));
AND2X1   g3424(.A(n5749), .B(g6035), .Y(n8071));
INVX1    g3425(.A(g6044), .Y(n8072));
NAND2X1  g3426(.A(n8072), .B(g35), .Y(n8073));
OAI22X1  g3427(.A0(n8071), .A1(n8073), .B0(n6946), .B1(g35), .Y(n3373));
MX2X1    g3428(.A(g441), .B(g475), .S0(n5688), .Y(n8075));
MX2X1    g3429(.A(g475), .B(n8075), .S0(g35), .Y(n3378));
MX2X1    g3430(.A(g5062), .B(g5343), .S0(g35), .Y(n3383));
NAND3X1  g3431(.A(g3976), .B(g3905), .C(n7411), .Y(n8078));
NAND3X1  g3432(.A(g3893), .B(g4005), .C(g4040), .Y(n8079));
AOI21X1  g3433(.A0(n8079), .A1(n8078), .B0(n6866), .Y(n8080));
NAND4X1  g3434(.A(g3925), .B(g4019), .C(n7411), .D(n5187), .Y(n8081));
NAND3X1  g3435(.A(g4000), .B(g3901), .C(n7411), .Y(n8082));
OAI21X1  g3436(.A0(n8082), .A1(n6860), .B0(n8081), .Y(n8083));
NOR2X1   g3437(.A(n8083), .B(n8080), .Y(n8084));
AND2X1   g3438(.A(g4019), .B(g4040), .Y(n8085));
NAND4X1  g3439(.A(n6865), .B(g3917), .C(g4054), .D(n8085), .Y(n8086));
NAND4X1  g3440(.A(g4027), .B(g3949), .C(g4040), .D(n5187), .Y(n8087));
NAND4X1  g3441(.A(g4000), .B(g3889), .C(g4040), .D(n6862), .Y(n8088));
AND2X1   g3442(.A(g4023), .B(g4040), .Y(n8089));
NAND4X1  g3443(.A(g3990), .B(n6859_1), .C(g3933), .D(n8089), .Y(n8090));
NAND4X1  g3444(.A(n8088), .B(n8087), .C(n8086), .D(n8090), .Y(n8091));
NAND4X1  g3445(.A(g3941), .B(g4023), .C(n7411), .D(n6862), .Y(n8092));
NAND3X1  g3446(.A(g4027), .B(g3957), .C(n7411), .Y(n8093));
OAI21X1  g3447(.A0(n8093), .A1(n6866), .B0(n8092), .Y(n8094));
NAND4X1  g3448(.A(g4031), .B(g3897), .C(g4040), .D(n6862), .Y(n8095));
NAND4X1  g3449(.A(g3976), .B(g3965), .C(g4040), .D(n5187), .Y(n8096));
NAND2X1  g3450(.A(n8096), .B(n8095), .Y(n8097));
NOR3X1   g3451(.A(n8097), .B(n8094), .C(n8091), .Y(n8098));
XOR2X1   g3452(.A(g4005), .B(n7411), .Y(n8099));
AND2X1   g3453(.A(g3937), .B(g4012), .Y(n8100));
AND2X1   g3454(.A(n8100), .B(n5187), .Y(n8101));
NAND3X1  g3455(.A(n6862), .B(g3929), .C(g3983), .Y(n8102));
NAND4X1  g3456(.A(n6865), .B(g4012), .C(g4054), .D(g3945), .Y(n8103));
AOI21X1  g3457(.A0(n8103), .A1(n8102), .B0(n8099), .Y(n8104));
AOI21X1  g3458(.A0(n8101), .A1(n8099), .B0(n8104), .Y(n8105));
NAND4X1  g3459(.A(g3961), .B(n6859_1), .C(g3969), .D(g3990), .Y(n8106));
NOR2X1   g3460(.A(n8106), .B(n8099), .Y(n8107));
NAND4X1  g3461(.A(g4005), .B(g3909), .C(n7411), .D(n5187), .Y(n8108));
NAND3X1  g3462(.A(g3913), .B(g4031), .C(n7411), .Y(n8109));
OAI21X1  g3463(.A0(n8109), .A1(n6860), .B0(n8108), .Y(n8110));
INVX1    g3464(.A(n8099), .Y(n8111));
NAND3X1  g3465(.A(n6862), .B(g3953), .C(g3969), .Y(n8112));
NAND4X1  g3466(.A(g3990), .B(g3983), .C(n6859_1), .D(g3921), .Y(n8113));
AOI21X1  g3467(.A0(n8113), .A1(n8112), .B0(n8111), .Y(n8114));
NOR3X1   g3468(.A(n8114), .B(n8110), .C(n8107), .Y(n8115));
NAND4X1  g3469(.A(n8105), .B(n8098), .C(n8084), .D(n8115), .Y(n8116));
AND2X1   g3470(.A(n7136), .B(g3808), .Y(n8117));
XOR2X1   g3471(.A(n8117), .B(n8116), .Y(n8118));
MX2X1    g3472(.A(g3808), .B(n8118), .S0(n6856), .Y(n8119));
MX2X1    g3473(.A(g3813), .B(n8119), .S0(g35), .Y(n3388));
INVX1    g3474(.A(g3747), .Y(n8121));
NAND3X1  g3475(.A(n7370), .B(n7369), .C(g35), .Y(n8122));
OAI21X1  g3476(.A0(n8121), .A1(g35), .B0(n8122), .Y(n3398));
AOI21X1  g3477(.A0(g4473), .A1(g4467), .B0(g4462), .Y(n8124));
NAND2X1  g3478(.A(n8124), .B(n7745), .Y(n8125));
OR2X1    g3479(.A(g4581), .B(n4620), .Y(n8126));
MX2X1    g3480(.A(n8125), .B(n8126), .S0(n4620), .Y(n3403));
NOR4X1   g3481(.A(n7041), .B(n4850), .C(g3873), .D(n7642), .Y(n8128));
MX2X1    g3482(.A(g3957), .B(n5592_1), .S0(n8128), .Y(n8129));
MX2X1    g3483(.A(g3941), .B(n8129), .S0(g35), .Y(n3408));
NOR3X1   g3484(.A(n6474), .B(n4840), .C(n6689), .Y(n8131));
XOR2X1   g3485(.A(n8131), .B(n4830), .Y(n8132));
OAI22X1  g3486(.A0(n7630), .A1(n8132), .B0(n4840), .B1(g35), .Y(n3413));
NOR2X1   g3487(.A(n6468_1), .B(n6467), .Y(n8134));
INVX1    g3488(.A(g1783), .Y(n8135));
OAI21X1  g3489(.A0(n8135), .A1(g1760), .B0(n4941), .Y(n8136));
OAI21X1  g3490(.A0(n6204), .A1(n4925_1), .B0(n8136), .Y(n8137));
MX2X1    g3491(.A(g1760), .B(n8137), .S0(n8134), .Y(n8138));
MX2X1    g3492(.A(g1768), .B(n8138), .S0(g35), .Y(n3418));
OAI22X1  g3493(.A0(g6358), .A1(n6996), .B0(n6995), .B1(g6351), .Y(n8140));
MX2X1    g3494(.A(g6346), .B(n6996), .S0(g6322), .Y(n8141));
OAI21X1  g3495(.A0(n6997), .A1(g6329), .B0(g35), .Y(n8142));
NOR4X1   g3496(.A(n8141), .B(n8140), .C(n6998_1), .D(n8142), .Y(n3427));
INVX1    g3497(.A(g160), .Y(n8144));
NAND3X1  g3498(.A(n7310_1), .B(n7308), .C(n7306_1), .Y(n8145));
NOR3X1   g3499(.A(n7302_1), .B(n5661), .C(n8144), .Y(n8146));
MX2X1    g3500(.A(n8144), .B(n8146), .S0(n8145), .Y(n8147));
MX2X1    g3501(.A(g157), .B(n8147), .S0(g35), .Y(n3431));
AND2X1   g3502(.A(g5428), .B(g5436), .Y(n8149));
AND2X1   g3503(.A(n8149), .B(g5441), .Y(n8150));
XOR2X1   g3504(.A(n8150), .B(g5445), .Y(n8151));
MX2X1    g3505(.A(g5441), .B(n8151), .S0(g35), .Y(n3436));
MX2X1    g3506(.A(g5366), .B(g5406), .S0(g5360), .Y(n8153));
OR2X1    g3507(.A(n8153), .B(n7983), .Y(n8154));
NAND2X1  g3508(.A(n8153), .B(n7983), .Y(n8155));
OAI21X1  g3509(.A0(n8154), .A1(n6646), .B0(n8155), .Y(n8156));
MX2X1    g3510(.A(g5360), .B(n8156), .S0(g35), .Y(n3441));
MX2X1    g3511(.A(g2279), .B(g2273), .S0(n6894), .Y(n8158));
MX2X1    g3512(.A(g2273), .B(n8158), .S0(g35), .Y(n3446));
INVX1    g3513(.A(g3498), .Y(n8160));
OAI22X1  g3514(.A0(n5524), .A1(g4284), .B0(n8160), .B1(n4836_1), .Y(n8161));
OR4X1    g3515(.A(n5524), .B(g4284), .C(n8160), .D(n4836_1), .Y(n8162));
AOI21X1  g3516(.A0(n8162), .A1(n8161), .B0(n4620), .Y(n3451));
NAND2X1  g3517(.A(n6141_1), .B(n6140), .Y(n8164));
MX2X1    g3518(.A(n5385_1), .B(n6142), .S0(n8164), .Y(n8165));
MX2X1    g3519(.A(g572), .B(n8165), .S0(g35), .Y(n3456));
OAI21X1  g3520(.A0(n6204), .A1(n4919), .B0(n5860_1), .Y(n8167));
MX2X1    g3521(.A(g2619), .B(n8167), .S0(n6628_1), .Y(n8168));
MX2X1    g3522(.A(g2625), .B(n8168), .S0(g35), .Y(n3466));
AND2X1   g3523(.A(g1157), .B(g1171), .Y(n8170));
OAI21X1  g3524(.A0(n6761), .A1(n6079), .B0(n8170), .Y(n8171));
OAI22X1  g3525(.A0(n6752_1), .A1(n4665), .B0(g1183), .B1(n6761), .Y(n8172));
NAND2X1  g3526(.A(n8172), .B(n8171), .Y(n8173));
MX2X1    g3527(.A(g1171), .B(n8173), .S0(g35), .Y(n3471));
INVX1    g3528(.A(g1636), .Y(n8175));
NOR3X1   g3529(.A(n5758_1), .B(n8175), .C(g1668), .Y(n8176));
MX2X1    g3530(.A(g1608), .B(n5756), .S0(n8176), .Y(n8177));
MX2X1    g3531(.A(g1600), .B(n8177), .S0(g35), .Y(n3476));
NOR4X1   g3532(.A(n6466), .B(n5143), .C(n5136), .D(n5627), .Y(n8179));
XOR2X1   g3533(.A(n5165), .B(g112), .Y(n8180));
MX2X1    g3534(.A(g1779), .B(n8180), .S0(n8179), .Y(n8181));
MX2X1    g3535(.A(g1728), .B(n8181), .S0(g35), .Y(n3491));
INVX1    g3536(.A(g2652), .Y(n8183));
AOI21X1  g3537(.A0(n6629), .A1(g2610), .B0(n8183), .Y(n8184));
XOR2X1   g3538(.A(n8184), .B(g2638), .Y(n8185));
MX2X1    g3539(.A(n8185), .B(g2652), .S0(n5863), .Y(n8186));
MX2X1    g3540(.A(g2638), .B(n8186), .S0(g35), .Y(n3496));
NOR4X1   g3541(.A(n5786), .B(g2217), .C(n5797_1), .D(n5787_1), .Y(n8188));
MX2X1    g3542(.A(g2193), .B(n6709), .S0(n8188), .Y(n8189));
MX2X1    g3543(.A(g2173), .B(n8189), .S0(g35), .Y(n3505));
XOR2X1   g3544(.A(n7941), .B(g2393), .Y(n8191));
MX2X1    g3545(.A(g2389), .B(n8191), .S0(g35), .Y(n3510));
INVX1    g3546(.A(g5759), .Y(n8193));
INVX1    g3547(.A(g5763), .Y(n8194));
AOI21X1  g3548(.A0(n8193), .A1(g35), .B0(n8194), .Y(n3515));
MX2X1    g3549(.A(g718), .B(g661), .S0(n6389_1), .Y(n8196));
MX2X1    g3550(.A(g718), .B(n8196), .S0(g35), .Y(n3520));
INVX1    g3551(.A(g4950), .Y(n8198));
OR2X1    g3552(.A(n5930), .B(n8198), .Y(n8199));
OAI21X1  g3553(.A0(n5938), .A1(n5802_1), .B0(n8198), .Y(n8200));
NAND2X1  g3554(.A(n5945), .B(n5802_1), .Y(n8201));
INVX1    g3555(.A(g3698), .Y(n8202));
MX2X1    g3556(.A(n5177), .B(n5932), .S0(n8202), .Y(n8203));
NAND2X1  g3557(.A(n8203), .B(n8201), .Y(n8204));
NOR4X1   g3558(.A(n6806), .B(n4896_1), .C(g4899), .D(n7392_1), .Y(n8205));
OAI21X1  g3559(.A0(n8204), .A1(n8200), .B0(n8205), .Y(n8206));
AOI21X1  g3560(.A0(n8206), .A1(n8199), .B0(n4620), .Y(n3525));
OAI21X1  g3561(.A0(n4868), .A1(n4866_1), .B0(g5535), .Y(n8208));
NAND3X1  g3562(.A(g5527), .B(n4867), .C(g5523), .Y(n8209));
AOI21X1  g3563(.A0(n8209), .A1(n8208), .B0(n6932), .Y(n8210));
MX2X1    g3564(.A(g5527), .B(n8210), .S0(g35), .Y(n3530));
MX2X1    g3565(.A(g2803), .B(n6313), .S0(g35), .Y(n3535));
OAI21X1  g3566(.A0(n7286), .A1(g1345), .B0(n5986), .Y(n8213));
MX2X1    g3567(.A(n7289), .B(g1361), .S0(n8213), .Y(n8214));
MX2X1    g3568(.A(g1345), .B(n8214), .S0(g35), .Y(n3540));
INVX1    g3569(.A(g3416), .Y(n8216));
NOR2X1   g3570(.A(n8216), .B(g3412), .Y(n8217));
NOR2X1   g3571(.A(n8216), .B(g3408), .Y(n8218));
MX2X1    g3572(.A(n8217), .B(n8218), .S0(g3423), .Y(n8219));
MX2X1    g3573(.A(g3416), .B(n8219), .S0(g35), .Y(n3545));
NOR4X1   g3574(.A(g6203), .B(g6209), .C(g6215), .D(n7379), .Y(n8221));
MX2X1    g3575(.A(g6235), .B(n5592_1), .S0(n8221), .Y(n8222));
MX2X1    g3576(.A(g6227), .B(n8222), .S0(g35), .Y(n3550));
INVX1    g3577(.A(g1146), .Y(n8224));
OAI21X1  g3578(.A0(g1152), .A1(n8224), .B0(g1099), .Y(n8225));
MX2X1    g3579(.A(g1146), .B(n8225), .S0(n6189), .Y(n8226));
AND2X1   g3580(.A(n8226), .B(g35), .Y(n3555));
NOR3X1   g3581(.A(n5863), .B(n6466), .C(n4919), .Y(n8228));
NOR2X1   g3582(.A(n4934_1), .B(g2610), .Y(n8229));
XOR2X1   g3583(.A(n8229), .B(g110), .Y(n8230));
MX2X1    g3584(.A(g2625), .B(n8230), .S0(n8228), .Y(n8231));
MX2X1    g3585(.A(g2610), .B(n8231), .S0(g35), .Y(n3560));
NOR3X1   g3586(.A(n7305), .B(n7304), .C(n7297), .Y(n8233));
NOR3X1   g3587(.A(n7302_1), .B(n5661), .C(n7296), .Y(n8234));
MX2X1    g3588(.A(n8234), .B(n7296), .S0(n8233), .Y(n8235));
MX2X1    g3589(.A(g164), .B(n8235), .S0(g35), .Y(n3565));
XOR2X1   g3590(.A(g1691), .B(g1687), .Y(n8237));
NOR4X1   g3591(.A(n5787_1), .B(n4629), .C(g1624), .D(n6501), .Y(n8238));
MX2X1    g3592(.A(g1696), .B(n8237), .S0(n8238), .Y(n8239));
MX2X1    g3593(.A(g1691), .B(n8239), .S0(g35), .Y(n3570));
NAND2X1  g3594(.A(g6555), .B(n7524), .Y(n8241));
NAND2X1  g3595(.A(n7204), .B(g6549), .Y(n8242));
AOI21X1  g3596(.A0(n8242), .A1(n8241), .B0(n7626), .Y(n8243));
MX2X1    g3597(.A(g6549), .B(n8243), .S0(g35), .Y(n3575));
AND2X1   g3598(.A(g106), .B(g35), .Y(n3580));
NAND3X1  g3599(.A(n6412), .B(g3376), .C(g3380), .Y(n8246));
NAND3X1  g3600(.A(n6414_1), .B(n6409_1), .C(n5772), .Y(n8247));
AND2X1   g3601(.A(n8247), .B(n8246), .Y(n8248));
NOR2X1   g3602(.A(n5778_1), .B(n5769), .Y(n8249));
MX2X1    g3603(.A(n5769), .B(n8249), .S0(n8248), .Y(n8250));
MX2X1    g3604(.A(g3380), .B(n8250), .S0(g35), .Y(n3584));
OAI21X1  g3605(.A0(n4849), .A1(n4848), .B0(g3881), .Y(n8252));
NAND3X1  g3606(.A(n4850), .B(g3869), .C(g3873), .Y(n8253));
AOI21X1  g3607(.A0(n8253), .A1(n8252), .B0(n7849), .Y(n8254));
MX2X1    g3608(.A(g3873), .B(n8254), .S0(g35), .Y(n3589));
NOR3X1   g3609(.A(n7205), .B(g6555), .C(n7524), .Y(n8256));
MX2X1    g3610(.A(g6621), .B(n5592_1), .S0(n8256), .Y(n8257));
MX2X1    g3611(.A(g6601), .B(n8257), .S0(g35), .Y(n3594));
XOR2X1   g3612(.A(n4836_1), .B(g3470), .Y(n8259));
MX2X1    g3613(.A(g3466), .B(n8259), .S0(g35), .Y(n3599));
NOR2X1   g3614(.A(n7042_1), .B(n4849), .Y(n8261));
MX2X1    g3615(.A(g3897), .B(n5592_1), .S0(n8261), .Y(n8262));
MX2X1    g3616(.A(g3949), .B(n8262), .S0(g35), .Y(n3604));
AOI21X1  g3617(.A0(n7456), .A1(g667), .B0(n7004), .Y(n8264));
MX2X1    g3618(.A(g518), .B(n8264), .S0(n5880_1), .Y(n8265));
MX2X1    g3619(.A(g513), .B(n8265), .S0(g35), .Y(n3609));
NAND3X1  g3620(.A(n8003), .B(n8002), .C(g3025), .Y(n8267));
OAI21X1  g3621(.A0(n6594), .A1(n6589), .B0(n6592), .Y(n8268));
OAI21X1  g3622(.A0(n8267), .A1(n5584), .B0(n8268), .Y(n8269));
MX2X1    g3623(.A(g3021), .B(n8269), .S0(g35), .Y(n3614));
OAI21X1  g3624(.A0(g209), .A1(g538), .B0(g35), .Y(n8271));
AOI21X1  g3625(.A0(n7912), .A1(n3747), .B0(n8271), .Y(n3619));
NOR4X1   g3626(.A(n6466), .B(n5137), .C(g504), .D(n6002), .Y(n8273));
XOR2X1   g3627(.A(n5157), .B(g112), .Y(n8274));
MX2X1    g3628(.A(g2606), .B(n8274), .S0(n8273), .Y(n8275));
MX2X1    g3629(.A(g2555), .B(n8275), .S0(g35), .Y(n3624));
NOR4X1   g3630(.A(n5549), .B(n6000_1), .C(n6513), .D(n7603), .Y(n8277));
XOR2X1   g3631(.A(g1472), .B(g1467), .Y(n8278));
MX2X1    g3632(.A(g1472), .B(n8278), .S0(n8277), .Y(n8279));
MX2X1    g3633(.A(g1467), .B(n8279), .S0(g35), .Y(n3629));
INVX1    g3634(.A(g6109), .Y(n8281));
INVX1    g3635(.A(g6105), .Y(n8282));
AOI21X1  g3636(.A0(n8282), .A1(g35), .B0(n8281), .Y(n3634));
OAI21X1  g3637(.A0(n5516_1), .A1(g542), .B0(g35), .Y(n8284));
OAI22X1  g3638(.A0(n5652), .A1(n8284), .B0(n5324), .B1(g35), .Y(n3639));
OAI21X1  g3639(.A0(n4644), .A1(n4642_1), .B0(g5188), .Y(n8286));
NAND3X1  g3640(.A(g5176), .B(n4643), .C(g5180), .Y(n8287));
AOI21X1  g3641(.A0(n8287), .A1(n8286), .B0(n6042), .Y(n8288));
MX2X1    g3642(.A(g5180), .B(n8288), .S0(g35), .Y(n3644));
XOR2X1   g3643(.A(n5873), .B(g5689), .Y(n8290));
MX2X1    g3644(.A(g5685), .B(n8290), .S0(g35), .Y(n3649));
MX2X1    g3645(.A(g405), .B(g392), .S0(n5688), .Y(n8292));
MX2X1    g3646(.A(g392), .B(n8292), .S0(g35), .Y(n3659));
NOR4X1   g3647(.A(g5170), .B(g5176), .C(g5164), .D(n7933), .Y(n8294));
MX2X1    g3648(.A(g5216), .B(n5592_1), .S0(n8294), .Y(n8295));
MX2X1    g3649(.A(g5220), .B(n8295), .S0(g35), .Y(n3664));
NAND4X1  g3650(.A(g4688), .B(g4664), .C(g4653), .D(g4659), .Y(n8297));
NOR2X1   g3651(.A(n8297), .B(g4669), .Y(n8298));
AND2X1   g3652(.A(n8297), .B(g4669), .Y(n8299));
OAI21X1  g3653(.A0(n8299), .A1(n8298), .B0(n7822), .Y(n8300));
NAND2X1  g3654(.A(g4664), .B(n4620), .Y(n8301));
OAI21X1  g3655(.A0(n8300), .A1(n4620), .B0(n8301), .Y(n3674));
OR2X1    g3656(.A(g5428), .B(g5424), .Y(n8303));
INVX1    g3657(.A(g5417), .Y(n8304));
AOI22X1  g3658(.A0(g5421), .A1(n8304), .B0(g5428), .B1(g5424), .Y(n8305));
OAI21X1  g3659(.A0(n8303), .A1(n7186), .B0(n8305), .Y(n8306));
MX2X1    g3660(.A(g5424), .B(n8306), .S0(g35), .Y(n3679));
MX2X1    g3661(.A(g1236), .B(g1227), .S0(g35), .Y(n3684));
NAND2X1  g3662(.A(n5205), .B(n5204), .Y(n8309));
NAND4X1  g3663(.A(n5713_1), .B(g4643), .C(g35), .D(n5178), .Y(n8310));
NAND2X1  g3664(.A(g66), .B(n4620), .Y(n8311));
OAI21X1  g3665(.A0(n8310), .A1(n8309), .B0(n8311), .Y(n3689));
MX2X1    g3666(.A(g2860), .B(n4447), .S0(n5697), .Y(n8313));
MX2X1    g3667(.A(g2852), .B(n8313), .S0(g35), .Y(n3694));
AOI21X1  g3668(.A0(n4970), .A1(n4812_1), .B0(n6721), .Y(n8315));
MX2X1    g3669(.A(g4749), .B(g101), .S0(n6721), .Y(n8316));
MX2X1    g3670(.A(n8316), .B(g4743), .S0(n8315), .Y(n8317));
MX2X1    g3671(.A(g4749), .B(n8317), .S0(g35), .Y(n3699));
NOR3X1   g3672(.A(g6561), .B(g6555), .C(g6549), .Y(n8319));
NAND3X1  g3673(.A(n8319), .B(n4855), .C(g6573), .Y(n8320));
MX2X1    g3674(.A(n5592_1), .B(g6593), .S0(n8320), .Y(n8321));
MX2X1    g3675(.A(g6597), .B(n8321), .S0(g35), .Y(n3704));
NOR2X1   g3676(.A(n5272), .B(g35), .Y(n3709));
INVX1    g3677(.A(g218), .Y(n8324));
MX2X1    g3678(.A(g209), .B(n8324), .S0(g35), .Y(n3714));
INVX1    g3679(.A(n4712_1), .Y(n8326));
NAND3X1  g3680(.A(g1379), .B(g1367), .C(g1345), .Y(n8327));
NOR3X1   g3681(.A(n8327), .B(n5985), .C(n5984), .Y(n8328));
INVX1    g3682(.A(g1500), .Y(n8329));
NAND2X1  g3683(.A(g1521), .B(g1339), .Y(n8330));
NOR3X1   g3684(.A(n8330), .B(g1532), .C(n8329), .Y(n8331));
OAI21X1  g3685(.A0(n8328), .A1(n8326), .B0(n8331), .Y(n8332));
AOI21X1  g3686(.A0(n7601), .A1(g1536), .B0(n8332), .Y(n8333));
INVX1    g3687(.A(g1413), .Y(n8334));
NOR2X1   g3688(.A(n8330), .B(g1532), .Y(n8335));
NOR3X1   g3689(.A(n8335), .B(n7601), .C(n8329), .Y(n8336));
NAND3X1  g3690(.A(n8336), .B(g1542), .C(n8334), .Y(n8337));
INVX1    g3691(.A(g1542), .Y(n8338));
INVX1    g3692(.A(n8336), .Y(n8339));
OAI21X1  g3693(.A0(n8339), .A1(n8338), .B0(g1413), .Y(n8340));
AOI21X1  g3694(.A0(n8340), .A1(n8337), .B0(n8333), .Y(n8341));
MX2X1    g3695(.A(g1542), .B(n8341), .S0(g35), .Y(n3723));
NOR3X1   g3696(.A(n7657), .B(n7204), .C(n7524), .Y(n8343));
MX2X1    g3697(.A(g6641), .B(n5592_1), .S0(n8343), .Y(n8344));
MX2X1    g3698(.A(g6625), .B(n8344), .S0(g35), .Y(n3737));
MX2X1    g3699(.A(n6591), .B(n6596), .S0(n5575), .Y(n8346));
NOR2X1   g3700(.A(n5584), .B(n5924_1), .Y(n8347));
MX2X1    g3701(.A(n8347), .B(n5924_1), .S0(n8346), .Y(n8348));
MX2X1    g3702(.A(g3040), .B(n8348), .S0(g35), .Y(n3742));
NAND3X1  g3703(.A(n6223), .B(n6222), .C(g1906), .Y(n8350));
OAI21X1  g3704(.A0(n6222), .A1(n5161), .B0(n8350), .Y(n8351));
MX2X1    g3705(.A(g1906), .B(n8351), .S0(g35), .Y(n3752));
NAND2X1  g3706(.A(n5962), .B(n5282), .Y(n8353));
NAND2X1  g3707(.A(n5962), .B(g22), .Y(n8354));
NAND2X1  g3708(.A(n8354), .B(n8353), .Y(n3757));
OAI21X1  g3709(.A0(g686), .A1(n5876), .B0(n6234), .Y(n8356));
MX2X1    g3710(.A(g504), .B(n8356), .S0(n5880_1), .Y(n8357));
MX2X1    g3711(.A(g499), .B(n8357), .S0(g35), .Y(n3762));
OAI21X1  g3712(.A0(g2587), .A1(n5860_1), .B0(n4934_1), .Y(n8359));
OAI21X1  g3713(.A0(n6204), .A1(n4919), .B0(n8359), .Y(n8360));
MX2X1    g3714(.A(g2587), .B(n8360), .S0(n6628_1), .Y(n8361));
MX2X1    g3715(.A(g2595), .B(n8361), .S0(g35), .Y(n3767));
NAND3X1  g3716(.A(n7445), .B(g73), .C(g72), .Y(n8363));
MX2X1    g3717(.A(g4372), .B(n8363), .S0(g4581), .Y(n8364));
MX2X1    g3718(.A(g4477), .B(n8364), .S0(g35), .Y(n3772));
NAND2X1  g3719(.A(g2331), .B(n6032), .Y(n8366));
AOI21X1  g3720(.A0(n5551_1), .A1(n5545), .B0(n8366), .Y(n8367));
MX2X1    g3721(.A(g2311), .B(n5547), .S0(n8367), .Y(n8368));
MX2X1    g3722(.A(g2315), .B(n8368), .S0(g35), .Y(n3777));
NOR4X1   g3723(.A(g3530), .B(n5735), .C(n5733_1), .D(n4835), .Y(n8370));
MX2X1    g3724(.A(g3602), .B(n5592_1), .S0(n8370), .Y(n8371));
MX2X1    g3725(.A(g3586), .B(n8371), .S0(g35), .Y(n3782));
NOR3X1   g3726(.A(n5899_1), .B(g5517), .C(n5854), .Y(n8373));
MX2X1    g3727(.A(g5571), .B(n5592_1), .S0(n8373), .Y(n8374));
MX2X1    g3728(.A(g5543), .B(n8374), .S0(g35), .Y(n3787));
NOR4X1   g3729(.A(n4833), .B(n5735), .C(g3512), .D(n4835), .Y(n8376));
MX2X1    g3730(.A(g3578), .B(n5592_1), .S0(n8376), .Y(n8377));
MX2X1    g3731(.A(g3558), .B(n8377), .S0(g35), .Y(n3792));
MX2X1    g3732(.A(g468), .B(g464), .S0(n5601), .Y(n8379));
MX2X1    g3733(.A(g464), .B(n8379), .S0(g35), .Y(n3797));
AND2X1   g3734(.A(g5535), .B(g35), .Y(n3802));
INVX1    g3735(.A(g3759), .Y(n8382));
INVX1    g3736(.A(g3763), .Y(n8383));
AOI21X1  g3737(.A0(n8382), .A1(g35), .B0(n8383), .Y(n3807));
MX2X1    g3738(.A(g5827), .B(g5821), .S0(n6749), .Y(n8385));
MX2X1    g3739(.A(g5821), .B(n8385), .S0(g35), .Y(n3812));
NOR3X1   g3740(.A(n6067), .B(g3506), .C(n5733_1), .Y(n8387));
MX2X1    g3741(.A(g3582), .B(n5592_1), .S0(n8387), .Y(n8388));
MX2X1    g3742(.A(g3566), .B(n8388), .S0(g35), .Y(n3817));
NOR4X1   g3743(.A(n4873), .B(g6209), .C(g6219), .D(n6208), .Y(n8390));
MX2X1    g3744(.A(g6271), .B(n5592_1), .S0(n8390), .Y(n8391));
MX2X1    g3745(.A(g6247), .B(n8391), .S0(g35), .Y(n3822));
AOI21X1  g3746(.A0(n6216_1), .A1(g35), .B0(n6744), .Y(n3827));
OR2X1    g3747(.A(g5774), .B(g5770), .Y(n8394));
AOI22X1  g3748(.A0(g5774), .A1(g5770), .B0(g5767), .B1(n8194), .Y(n8395));
OAI21X1  g3749(.A0(n8394), .A1(n7648), .B0(n8395), .Y(n8396));
MX2X1    g3750(.A(g5770), .B(n8396), .S0(g35), .Y(n3832));
MX2X1    g3751(.A(g2380), .B(g2375), .S0(n5553), .Y(n8398));
MX2X1    g3752(.A(g2375), .B(n8398), .S0(g35), .Y(n3837));
NOR4X1   g3753(.A(g5170), .B(g5176), .C(g5164), .D(n6195), .Y(n8400));
MX2X1    g3754(.A(g5196), .B(n5592_1), .S0(n8400), .Y(n8401));
MX2X1    g3755(.A(g5188), .B(n8401), .S0(g35), .Y(n3842));
NAND3X1  g3756(.A(n7985), .B(g5381), .C(g5385), .Y(n8403));
NOR2X1   g3757(.A(n8403), .B(n6638_1), .Y(n8404));
NAND3X1  g3758(.A(n7987), .B(n7982), .C(n6640), .Y(n8405));
NOR2X1   g3759(.A(n8405), .B(g5390), .Y(n8406));
OAI21X1  g3760(.A0(n8406), .A1(n8404), .B0(n6637), .Y(n8407));
OR4X1    g3761(.A(n8404), .B(n6646), .C(n6637), .D(n8406), .Y(n8408));
NAND2X1  g3762(.A(n8408), .B(n8407), .Y(n8409));
MX2X1    g3763(.A(g5390), .B(n8409), .S0(g35), .Y(n3847));
NOR3X1   g3764(.A(n5594), .B(g3161), .C(n5913), .Y(n8411));
MX2X1    g3765(.A(g3227), .B(n5592_1), .S0(n8411), .Y(n8412));
MX2X1    g3766(.A(g3207), .B(n8412), .S0(g35), .Y(n3852));
NAND2X1  g3767(.A(n7842), .B(g2040), .Y(n8414));
AOI21X1  g3768(.A0(n6084), .A1(n6081), .B0(n8414), .Y(n8415));
MX2X1    g3769(.A(g2020), .B(n7037_1), .S0(n8415), .Y(n8416));
MX2X1    g3770(.A(g2024), .B(n8416), .S0(g35), .Y(n3857));
INVX1    g3771(.A(g6541), .Y(n8418));
OAI22X1  g3772(.A0(n5524), .A1(g4284), .B0(n8418), .B1(n4857), .Y(n8419));
OR4X1    g3773(.A(n5524), .B(g4284), .C(n8418), .D(n4857), .Y(n8420));
AOI21X1  g3774(.A0(n8420), .A1(n8419), .B0(n4620), .Y(n3871));
NOR3X1   g3775(.A(n4845), .B(g3179), .C(n4843), .Y(n8422));
MX2X1    g3776(.A(g3203), .B(n5592_1), .S0(n8422), .Y(n8423));
MX2X1    g3777(.A(g3251), .B(n8423), .S0(g35), .Y(n3876));
NAND4X1  g3778(.A(n5637), .B(g112), .C(n4824), .D(n5144), .Y(n8425));
NAND3X1  g3779(.A(n8425), .B(n7211), .C(g1636), .Y(n8426));
OAI21X1  g3780(.A0(n7211), .A1(n4631), .B0(n8426), .Y(n8427));
MX2X1    g3781(.A(g1636), .B(n8427), .S0(g35), .Y(n3881));
INVX1    g3782(.A(g4760), .Y(n8429));
OR2X1    g3783(.A(n6746), .B(n8429), .Y(n8430));
INVX1    g3784(.A(g6040), .Y(n8431));
OAI21X1  g3785(.A0(n6952), .A1(n8431), .B0(n8429), .Y(n8432));
NAND2X1  g3786(.A(n6959), .B(n8431), .Y(n8433));
NAND3X1  g3787(.A(g6049), .B(n8072), .C(n6944), .Y(n8434));
NAND3X1  g3788(.A(g6049), .B(g6044), .C(g5990), .Y(n8435));
NAND3X1  g3789(.A(n8435), .B(n8434), .C(n8433), .Y(n8436));
OR2X1    g3790(.A(n8436), .B(n8432), .Y(n8437));
NAND4X1  g3791(.A(n6746), .B(n4970), .C(n6720), .D(n8437), .Y(n8438));
AOI21X1  g3792(.A0(n8438), .A1(n8430), .B0(n4620), .Y(n3886));
MX2X1    g3793(.A(g262), .B(g878), .S0(n7408), .Y(n8440));
MX2X1    g3794(.A(g232), .B(n8440), .S0(g35), .Y(n3891));
NOR3X1   g3795(.A(n5628), .B(g1728), .C(g1802), .Y(n8442));
MX2X1    g3796(.A(g1840), .B(g1834), .S0(n8442), .Y(n8443));
MX2X1    g3797(.A(g1834), .B(n8443), .S0(g35), .Y(n3896));
MX2X1    g3798(.A(g5467), .B(g5503), .S0(n4869), .Y(n8445));
MX2X1    g3799(.A(g5503), .B(n8445), .S0(g35), .Y(n3906));
MX2X1    g3800(.A(g460), .B(g246), .S0(n5601), .Y(n8447));
MX2X1    g3801(.A(g168), .B(n8447), .S0(g35), .Y(n3911));
NAND2X1  g3802(.A(n6208), .B(g6209), .Y(n8449));
NAND2X1  g3803(.A(g6203), .B(n5980), .Y(n8450));
AOI21X1  g3804(.A0(n8450), .A1(n8449), .B0(n5646), .Y(n8451));
MX2X1    g3805(.A(g6203), .B(n8451), .S0(g35), .Y(n3916));
NOR2X1   g3806(.A(n7219), .B(n7218), .Y(n8453));
OAI21X1  g3807(.A0(g74), .A1(g351), .B0(g35), .Y(n8454));
NAND2X1  g3808(.A(g355), .B(n4620), .Y(n8455));
OAI21X1  g3809(.A0(n8454), .A1(n8453), .B0(n8455), .Y(n3921));
MX2X1    g3810(.A(g650), .B(g655), .S0(n6389_1), .Y(n8457));
MX2X1    g3811(.A(g650), .B(n8457), .S0(g35), .Y(n3930));
MX2X1    g3812(.A(g3502), .B(n6676), .S0(n6435), .Y(n8459));
AND2X1   g3813(.A(n8459), .B(g35), .Y(n3935));
NOR4X1   g3814(.A(n6466), .B(n5134), .C(g504), .D(n6707), .Y(n8461));
XOR2X1   g3815(.A(n5160), .B(g112), .Y(n8462));
MX2X1    g3816(.A(g2204), .B(n8462), .S0(n8461), .Y(n8463));
MX2X1    g3817(.A(g2153), .B(n8463), .S0(g35), .Y(n3940));
NOR3X1   g3818(.A(n6195), .B(n6624), .C(n5610), .Y(n8465));
MX2X1    g3819(.A(g5256), .B(n5592_1), .S0(n8465), .Y(n8466));
MX2X1    g3820(.A(g5240), .B(n8466), .S0(g35), .Y(n3945));
INVX1    g3821(.A(g4601), .Y(n8468));
NOR3X1   g3822(.A(n6024_1), .B(n8468), .C(n5720), .Y(n8469));
NOR2X1   g3823(.A(n6023), .B(n5716), .Y(n8470));
NOR2X1   g3824(.A(n6023), .B(g4608), .Y(n8471));
MX2X1    g3825(.A(n8470), .B(n8471), .S0(n8469), .Y(n8472));
MX2X1    g3826(.A(g4601), .B(n8472), .S0(g35), .Y(n3950));
MX2X1    g3827(.A(n5682), .B(n5383), .S0(n5681), .Y(n8474));
MX2X1    g3828(.A(g790), .B(n8474), .S0(g35), .Y(n3955));
NOR3X1   g3829(.A(n5806), .B(n5804), .C(n5803), .Y(n8476));
XOR2X1   g3830(.A(n8476), .B(g3689), .Y(n8477));
MX2X1    g3831(.A(g3680), .B(n8477), .S0(g35), .Y(n3969));
NAND3X1  g3832(.A(n7988), .B(n7986), .C(g5381), .Y(n8479));
OAI21X1  g3833(.A0(n7987), .A1(n7985), .B0(n7982), .Y(n8480));
OAI21X1  g3834(.A0(n8479), .A1(n6646), .B0(n8480), .Y(n8481));
MX2X1    g3835(.A(g5377), .B(n8481), .S0(g35), .Y(n3974));
NAND4X1  g3836(.A(g817), .B(g822), .C(n7156), .D(g723), .Y(n8483));
NAND2X1  g3837(.A(g703), .B(n7156), .Y(n8484));
OAI21X1  g3838(.A0(n6247), .A1(n7157_1), .B0(g703), .Y(n8485));
NAND3X1  g3839(.A(n8485), .B(n8484), .C(n8483), .Y(n8486));
MX2X1    g3840(.A(g703), .B(n8486), .S0(n5688), .Y(n8487));
MX2X1    g3841(.A(g847), .B(n8487), .S0(g35), .Y(n3984));
INVX1    g3842(.A(g5413), .Y(n8489));
AOI21X1  g3843(.A0(n8489), .A1(g35), .B0(n8304), .Y(n3989));
MX2X1    g3844(.A(g862), .B(n4882), .S0(g896), .Y(n8491));
MX2X1    g3845(.A(g890), .B(n8491), .S0(g35), .Y(n3994));
NOR3X1   g3846(.A(n7506_1), .B(n5593), .C(n5913), .Y(n8493));
MX2X1    g3847(.A(g3247), .B(n5592_1), .S0(n8493), .Y(n8494));
MX2X1    g3848(.A(g3231), .B(n8494), .S0(g35), .Y(n3999));
INVX1    g3849(.A(g2040), .Y(n8496));
INVX1    g3850(.A(n6085), .Y(n8497));
NAND4X1  g3851(.A(n5637), .B(g112), .C(n4824), .D(n5148), .Y(n8498));
NAND3X1  g3852(.A(n8498), .B(n8497), .C(g1996), .Y(n8499));
OAI21X1  g3853(.A0(n8497), .A1(n8496), .B0(n8499), .Y(n8500));
MX2X1    g3854(.A(g2047), .B(n8500), .S0(g35), .Y(n4004));
MX2X1    g3855(.A(g4146), .B(n4586), .S0(n5697), .Y(n8502));
MX2X1    g3856(.A(g4176), .B(n8502), .S0(g35), .Y(n4014));
NAND3X1  g3857(.A(g4628), .B(g4639), .C(g4621), .Y(n8504));
NOR2X1   g3858(.A(n8504), .B(g4633), .Y(n8505));
AND2X1   g3859(.A(n8504), .B(g4633), .Y(n8506));
OAI21X1  g3860(.A0(n8506), .A1(n8505), .B0(n5846), .Y(n8507));
NAND2X1  g3861(.A(g4628), .B(n4620), .Y(n8508));
OAI21X1  g3862(.A0(n8507), .A1(n4620), .B0(n8508), .Y(n4019));
XOR2X1   g3863(.A(g1236), .B(g979), .Y(n8510));
NAND4X1  g3864(.A(n6059), .B(n6050), .C(n4708), .D(n8510), .Y(n8511));
OR2X1    g3865(.A(g1239), .B(g1116), .Y(n8512));
OR4X1    g3866(.A(g1056), .B(g1157), .C(g990), .D(n8512), .Y(n8513));
XOR2X1   g3867(.A(n8513), .B(n8511), .Y(n8514));
MX2X1    g3868(.A(g996), .B(n8514), .S0(g35), .Y(n4024));
NOR3X1   g3869(.A(n7059), .B(n7058), .C(n7057), .Y(n8516));
NOR3X1   g3870(.A(g5706), .B(g5719), .C(n7065_1), .Y(n8517));
OAI21X1  g3871(.A0(n8517), .A1(n8516), .B0(n7060_1), .Y(n8518));
NOR2X1   g3872(.A(n8517), .B(n8516), .Y(n8519));
NAND2X1  g3873(.A(n8519), .B(g5723), .Y(n8520));
OAI21X1  g3874(.A0(n8520), .A1(n7077), .B0(n8518), .Y(n8521));
MX2X1    g3875(.A(g5719), .B(n8521), .S0(g35), .Y(n4029));
MX2X1    g3876(.A(g4732), .B(n6676), .S0(n6494), .Y(n8523));
MX2X1    g3877(.A(g4727), .B(n8523), .S0(g35), .Y(n4034));
AND2X1   g3878(.A(g5188), .B(g35), .Y(n4039));
XOR2X1   g3879(.A(g5808), .B(g5813), .Y(n8526));
MX2X1    g3880(.A(g5817), .B(n8526), .S0(n6749), .Y(n8527));
MX2X1    g3881(.A(g5808), .B(n8527), .S0(g35), .Y(n4043));
NOR2X1   g3882(.A(n5269_1), .B(g35), .Y(n4048));
OAI21X1  g3883(.A0(n6204), .A1(n4918), .B0(n7551), .Y(n8530));
MX2X1    g3884(.A(g2351), .B(n8530), .S0(n7227), .Y(n8531));
MX2X1    g3885(.A(g2357), .B(n8531), .S0(g35), .Y(n4053));
NOR3X1   g3886(.A(n6003), .B(g2555), .C(g2629), .Y(n8533));
MX2X1    g3887(.A(g2648), .B(g2643), .S0(n8533), .Y(n8534));
MX2X1    g3888(.A(g2643), .B(n8534), .S0(g35), .Y(n4058));
INVX1    g3889(.A(g6732), .Y(n8536));
INVX1    g3890(.A(g6727), .Y(n8537));
NOR4X1   g3891(.A(n6679), .B(n6678), .C(n8537), .D(n6680), .Y(n8538));
AOI21X1  g3892(.A0(n8538), .A1(g35), .B0(n8536), .Y(n4063));
AOI21X1  g3893(.A0(n4964_1), .A1(n6798), .B0(n6089), .Y(n8540));
MX2X1    g3894(.A(g4950), .B(g71), .S0(n6089), .Y(n8541));
MX2X1    g3895(.A(n8541), .B(g4944), .S0(n8540), .Y(n8542));
MX2X1    g3896(.A(g4950), .B(n8542), .S0(g35), .Y(n4068));
NAND4X1  g3897(.A(n4729), .B(g4098), .C(g4076), .D(n4731_1), .Y(n8544));
NAND3X1  g3898(.A(n4728), .B(n4830), .C(g4087), .Y(n8545));
NOR2X1   g3899(.A(n8545), .B(n8544), .Y(n8546));
INVX1    g3900(.A(g4169), .Y(n8547));
NAND2X1  g3901(.A(n8547), .B(g35), .Y(n8548));
OAI22X1  g3902(.A0(n8546), .A1(n8548), .B0(n4730), .B1(g35), .Y(n4073));
MX2X1    g3903(.A(g333), .B(n6918), .S0(g35), .Y(n4078));
XOR2X1   g3904(.A(g3462), .B(g3457), .Y(n8551));
MX2X1    g3905(.A(g3466), .B(n8551), .S0(n7393), .Y(n8552));
MX2X1    g3906(.A(g3457), .B(n8552), .S0(g35), .Y(n4087));
MX2X1    g3907(.A(g4145), .B(g4116), .S0(n6253), .Y(n8554));
MX2X1    g3908(.A(g4112), .B(n8554), .S0(g35), .Y(n4092));
MX2X1    g3909(.A(n7545_1), .B(n7546), .S0(n5486), .Y(n8556));
OR2X1    g3910(.A(n8556), .B(g5041), .Y(n8557));
NAND2X1  g3911(.A(n8556), .B(g5041), .Y(n8558));
OAI21X1  g3912(.A0(n8558), .A1(n5501), .B0(n8557), .Y(n8559));
MX2X1    g3913(.A(g5037), .B(n8559), .S0(g35), .Y(n4097));
XOR2X1   g3914(.A(n8149), .B(g5441), .Y(n8561));
MX2X1    g3915(.A(g5436), .B(n8561), .S0(g35), .Y(n4102));
INVX1    g3916(.A(g4452), .Y(n8563));
INVX1    g3917(.A(g4392), .Y(n8564));
NAND3X1  g3918(.A(n7415), .B(n8564), .C(g4430), .Y(n8565));
OAI21X1  g3919(.A0(n8565), .A1(n4620), .B0(n8563), .Y(n4107));
MX2X1    g3920(.A(g3827), .B(g3821), .S0(n7137_1), .Y(n8567));
MX2X1    g3921(.A(g3821), .B(n8567), .S0(g35), .Y(n4112));
INVX1    g3922(.A(g6682), .Y(n8569));
NAND2X1  g3923(.A(g6741), .B(n8569), .Y(n8570));
NAND3X1  g3924(.A(g6668), .B(g6597), .C(n8537), .Y(n8571));
NAND3X1  g3925(.A(g6697), .B(g6585), .C(g6727), .Y(n8572));
AOI21X1  g3926(.A0(n8572), .A1(n8571), .B0(n8570), .Y(n8573));
NAND4X1  g3927(.A(g6617), .B(g6711), .C(n8537), .D(n5190), .Y(n8574));
INVX1    g3928(.A(g6741), .Y(n8575));
NAND2X1  g3929(.A(n8575), .B(g6682), .Y(n8576));
NAND3X1  g3930(.A(g6593), .B(n8537), .C(g6692), .Y(n8577));
OAI21X1  g3931(.A0(n8577), .A1(n8576), .B0(n8574), .Y(n8578));
NOR2X1   g3932(.A(n8578), .B(n8573), .Y(n8579));
AND2X1   g3933(.A(g6711), .B(g6727), .Y(n8580));
NAND4X1  g3934(.A(g6609), .B(g6741), .C(n8569), .D(n8580), .Y(n8581));
NAND4X1  g3935(.A(g6719), .B(g6641), .C(g6727), .D(n5190), .Y(n8582));
NOR2X1   g3936(.A(g6741), .B(g6682), .Y(n8583));
NAND4X1  g3937(.A(g6581), .B(g6727), .C(g6692), .D(n8583), .Y(n8584));
AND2X1   g3938(.A(g6715), .B(g6727), .Y(n8585));
NAND4X1  g3939(.A(n8575), .B(g6682), .C(g6625), .D(n8585), .Y(n8586));
NAND4X1  g3940(.A(n8584), .B(n8582), .C(n8581), .D(n8586), .Y(n8587));
NAND4X1  g3941(.A(g6633), .B(g6715), .C(n8537), .D(n8583), .Y(n8588));
NAND3X1  g3942(.A(g6719), .B(g6649), .C(n8537), .Y(n8589));
OAI21X1  g3943(.A0(n8589), .A1(n8570), .B0(n8588), .Y(n8590));
NAND4X1  g3944(.A(g6723), .B(g6589), .C(g6727), .D(n8583), .Y(n8591));
NAND4X1  g3945(.A(g6657), .B(g6668), .C(g6727), .D(n5190), .Y(n8592));
NAND2X1  g3946(.A(n8592), .B(n8591), .Y(n8593));
NOR3X1   g3947(.A(n8593), .B(n8590), .C(n8587), .Y(n8594));
XOR2X1   g3948(.A(g6697), .B(n8537), .Y(n8595));
AND2X1   g3949(.A(g6704), .B(g6629), .Y(n8596));
AND2X1   g3950(.A(n8596), .B(n5190), .Y(n8597));
NAND3X1  g3951(.A(n8583), .B(g6675), .C(g6621), .Y(n8598));
NAND4X1  g3952(.A(g6741), .B(n8569), .C(g6637), .D(g6704), .Y(n8599));
AOI21X1  g3953(.A0(n8599), .A1(n8598), .B0(n8595), .Y(n8600));
AOI21X1  g3954(.A0(n8597), .A1(n8595), .B0(n8600), .Y(n8601));
NAND4X1  g3955(.A(n8575), .B(g6682), .C(g6653), .D(g6661), .Y(n8602));
NOR2X1   g3956(.A(n8602), .B(n8595), .Y(n8603));
NAND4X1  g3957(.A(g6601), .B(g6697), .C(n8537), .D(n5190), .Y(n8604));
NAND3X1  g3958(.A(g6605), .B(g6723), .C(n8537), .Y(n8605));
OAI21X1  g3959(.A0(n8605), .A1(n8576), .B0(n8604), .Y(n8606));
INVX1    g3960(.A(n8595), .Y(n8607));
NAND3X1  g3961(.A(n8583), .B(g6661), .C(g6645), .Y(n8608));
NAND4X1  g3962(.A(g6682), .B(g6675), .C(g6613), .D(n8575), .Y(n8609));
AOI21X1  g3963(.A0(n8609), .A1(n8608), .B0(n8607), .Y(n8610));
NOR3X1   g3964(.A(n8610), .B(n8606), .C(n8603), .Y(n8611));
NAND4X1  g3965(.A(n8601), .B(n8594), .C(n8579), .D(n8611), .Y(n8612));
AND2X1   g3966(.A(n7723), .B(g6500), .Y(n8613));
XOR2X1   g3967(.A(n8613), .B(n8612), .Y(n8614));
MX2X1    g3968(.A(g6500), .B(n8614), .S0(n7721), .Y(n8615));
MX2X1    g3969(.A(g6505), .B(n8615), .S0(g35), .Y(n4117));
NAND4X1  g3970(.A(g3352), .B(g3338), .C(g3288), .D(g3274), .Y(n8617));
NOR2X1   g3971(.A(n8617), .B(n7757), .Y(n8618));
XOR2X1   g3972(.A(n8618), .B(g3133), .Y(n8619));
MX2X1    g3973(.A(g3129), .B(n8619), .S0(g35), .Y(n4127));
NAND2X1  g3974(.A(g3352), .B(n7761), .Y(n8621));
NAND3X1  g3975(.A(g3274), .B(g3203), .C(n6824), .Y(n8622));
NAND3X1  g3976(.A(g3191), .B(g3303), .C(g3338), .Y(n8623));
AOI21X1  g3977(.A0(n8623), .A1(n8622), .B0(n8621), .Y(n8624));
NAND4X1  g3978(.A(g3223), .B(g3317), .C(n6824), .D(n5183), .Y(n8625));
NAND2X1  g3979(.A(n7759), .B(g3288), .Y(n8626));
NAND3X1  g3980(.A(g3199), .B(g3298), .C(n6824), .Y(n8627));
OAI21X1  g3981(.A0(n8627), .A1(n8626), .B0(n8625), .Y(n8628));
NOR2X1   g3982(.A(n8628), .B(n8624), .Y(n8629));
AND2X1   g3983(.A(g3317), .B(g3338), .Y(n8630));
NAND4X1  g3984(.A(g3352), .B(g3215), .C(n7761), .D(n8630), .Y(n8631));
NAND4X1  g3985(.A(g3325), .B(g3247), .C(g3338), .D(n5183), .Y(n8632));
NOR2X1   g3986(.A(g3352), .B(g3288), .Y(n8633));
NAND4X1  g3987(.A(g3187), .B(g3298), .C(g3338), .D(n8633), .Y(n8634));
AND2X1   g3988(.A(g3338), .B(g3321), .Y(n8635));
NAND4X1  g3989(.A(n7759), .B(g3288), .C(g3231), .D(n8635), .Y(n8636));
NAND4X1  g3990(.A(n8634), .B(n8632), .C(n8631), .D(n8636), .Y(n8637));
NAND4X1  g3991(.A(n6824), .B(g3239), .C(g3321), .D(n8633), .Y(n8638));
NAND3X1  g3992(.A(g3325), .B(g3255), .C(n6824), .Y(n8639));
OAI21X1  g3993(.A0(n8639), .A1(n8621), .B0(n8638), .Y(n8640));
NAND4X1  g3994(.A(g3329), .B(g3195), .C(g3338), .D(n8633), .Y(n8641));
NAND4X1  g3995(.A(g3274), .B(g3263), .C(g3338), .D(n5183), .Y(n8642));
NAND2X1  g3996(.A(n8642), .B(n8641), .Y(n8643));
NOR3X1   g3997(.A(n8643), .B(n8640), .C(n8637), .Y(n8644));
XOR2X1   g3998(.A(g3303), .B(n6824), .Y(n8645));
AND2X1   g3999(.A(g3310), .B(g3235), .Y(n8646));
AND2X1   g4000(.A(n8646), .B(n5183), .Y(n8647));
NAND3X1  g4001(.A(n8633), .B(g3227), .C(g3281), .Y(n8648));
NAND4X1  g4002(.A(g3310), .B(n7761), .C(g3243), .D(g3352), .Y(n8649));
AOI21X1  g4003(.A0(n8649), .A1(n8648), .B0(n8645), .Y(n8650));
AOI21X1  g4004(.A0(n8647), .A1(n8645), .B0(n8650), .Y(n8651));
NAND4X1  g4005(.A(g3267), .B(g3259), .C(g3288), .D(n7759), .Y(n8652));
NOR2X1   g4006(.A(n8652), .B(n8645), .Y(n8653));
NAND4X1  g4007(.A(g3207), .B(g3303), .C(n6824), .D(n5183), .Y(n8654));
NAND3X1  g4008(.A(g3211), .B(g3329), .C(n6824), .Y(n8655));
OAI21X1  g4009(.A0(n8655), .A1(n8626), .B0(n8654), .Y(n8656));
INVX1    g4010(.A(n8645), .Y(n8657));
NAND3X1  g4011(.A(n8633), .B(g3251), .C(g3267), .Y(n8658));
NAND4X1  g4012(.A(g3219), .B(g3281), .C(g3288), .D(n7759), .Y(n8659));
AOI21X1  g4013(.A0(n8659), .A1(n8658), .B0(n8657), .Y(n8660));
NOR3X1   g4014(.A(n8660), .B(n8656), .C(n8653), .Y(n8661));
NAND4X1  g4015(.A(n8651), .B(n8644), .C(n8629), .D(n8661), .Y(n8662));
MX2X1    g4016(.A(g3333), .B(n8662), .S0(n7756), .Y(n8663));
MX2X1    g4017(.A(g3263), .B(n8663), .S0(g35), .Y(n4132));
AOI21X1  g4018(.A0(n6216_1), .A1(g35), .B0(n7014), .Y(n4141));
NAND3X1  g4019(.A(n6121), .B(n6119), .C(n6117), .Y(n8666));
MX2X1    g4020(.A(n7047_1), .B(n7048), .S0(n8666), .Y(n8667));
MX2X1    g4021(.A(g294), .B(n8667), .S0(g35), .Y(n4146));
OR2X1    g4022(.A(g3774), .B(g3770), .Y(n8669));
AOI22X1  g4023(.A0(g3774), .A1(g3770), .B0(g3767), .B1(n8383), .Y(n8670));
OAI21X1  g4024(.A0(n8669), .A1(n7928), .B0(n8670), .Y(n8671));
MX2X1    g4025(.A(g3770), .B(n8671), .S0(g35), .Y(n4151));
MX2X1    g4026(.A(g2667), .B(g2661), .S0(n8533), .Y(n8673));
MX2X1    g4027(.A(g2661), .B(n8673), .S0(g35), .Y(n4156));
INVX1    g4028(.A(g3396), .Y(n8675));
NOR3X1   g4029(.A(n8246), .B(n5770), .C(n5769), .Y(n8676));
NOR3X1   g4030(.A(n8247), .B(g3391), .C(g3385), .Y(n8677));
OR4X1    g4031(.A(n8676), .B(n5778_1), .C(n8675), .D(n8677), .Y(n8678));
OAI21X1  g4032(.A0(n8677), .A1(n8676), .B0(n8675), .Y(n8679));
NAND2X1  g4033(.A(n8679), .B(n8678), .Y(n8680));
MX2X1    g4034(.A(g3391), .B(n8680), .S0(g35), .Y(n4161));
OAI21X1  g4035(.A0(g1894), .A1(n6203), .B0(n4939_1), .Y(n8682));
OAI21X1  g4036(.A0(n6204), .A1(n4924), .B0(n8682), .Y(n8683));
MX2X1    g4037(.A(g1894), .B(n8683), .S0(n6202), .Y(n8684));
MX2X1    g4038(.A(g1902), .B(n8684), .S0(g35), .Y(n4171));
NOR3X1   g4039(.A(n5006), .B(n5004), .C(n5616), .Y(n8686));
MX2X1    g4040(.A(g2988), .B(n3393), .S0(n8686), .Y(n8687));
MX2X1    g4041(.A(g2994), .B(n8687), .S0(g35), .Y(n4176));
NOR4X1   g4042(.A(g3518), .B(g3506), .C(g3512), .D(n6067), .Y(n8689));
MX2X1    g4043(.A(g3538), .B(n5592_1), .S0(n8689), .Y(n8690));
MX2X1    g4044(.A(g3530), .B(n8690), .S0(g35), .Y(n4181));
AOI21X1  g4045(.A0(n8145), .A1(g35), .B0(n8144), .Y(n4186));
MX2X1    g4046(.A(g106), .B(g316), .S0(g35), .Y(n4191));
NOR3X1   g4047(.A(n7154), .B(n7153), .C(n7160), .Y(n8694));
NOR2X1   g4048(.A(n7158), .B(g827), .Y(n8695));
INVX1    g4049(.A(g827), .Y(n8696));
NOR2X1   g4050(.A(n7158), .B(n8696), .Y(n8697));
MX2X1    g4051(.A(n8697), .B(n8695), .S0(n8694), .Y(n8698));
MX2X1    g4052(.A(g822), .B(n8698), .S0(g35), .Y(n4196));
NAND3X1  g4053(.A(n6059), .B(n6050), .C(n4708), .Y(n8700));
OR4X1    g4054(.A(g1075), .B(g1079), .C(n4620), .D(g1083), .Y(n8701));
AOI21X1  g4055(.A0(n8700), .A1(n7487), .B0(n8701), .Y(n4201));
MX2X1    g4056(.A(n5825), .B(n5828), .S0(n5830), .Y(n8703));
OR2X1    g4057(.A(n8703), .B(g6077), .Y(n8704));
NAND2X1  g4058(.A(n8703), .B(g6077), .Y(n8705));
OAI21X1  g4059(.A0(n8705), .A1(n5820), .B0(n8704), .Y(n8706));
MX2X1    g4060(.A(g6073), .B(n8706), .S0(g35), .Y(n4205));
NAND3X1  g4061(.A(n6002), .B(n5995), .C(g2555), .Y(n8708));
AOI21X1  g4062(.A0(n5999), .A1(g2599), .B0(g2629), .Y(n8709));
NAND3X1  g4063(.A(n8709), .B(n7597), .C(n7596), .Y(n8710));
AOI21X1  g4064(.A0(n8710), .A1(n8708), .B0(n4620), .Y(n4210));
MX2X1    g4065(.A(g5011), .B(n8612), .S0(n7721), .Y(n8712));
MX2X1    g4066(.A(g6657), .B(n8712), .S0(g35), .Y(n4215));
AND2X1   g4067(.A(n7912), .B(n3220), .Y(n8714));
OAI21X1  g4068(.A0(g199), .A1(g222), .B0(g35), .Y(n8715));
OAI22X1  g4069(.A0(n8714), .A1(n8715), .B0(g23612), .B1(g35), .Y(n4220));
INVX1    g4070(.A(g6513), .Y(n8717));
XOR2X1   g4071(.A(n8717), .B(g6519), .Y(n8718));
MX2X1    g4072(.A(g6523), .B(n8718), .S0(n7724), .Y(n8719));
MX2X1    g4073(.A(g6519), .B(n8719), .S0(g35), .Y(n4225));
AND2X1   g4074(.A(g1514), .B(g1500), .Y(n8721));
OAI21X1  g4075(.A0(n8333), .A1(n6000_1), .B0(n8721), .Y(n8722));
OAI22X1  g4076(.A0(n5549), .A1(n8329), .B0(g1526), .B1(n8333), .Y(n8723));
NAND2X1  g4077(.A(n8723), .B(n8722), .Y(n8724));
MX2X1    g4078(.A(g1514), .B(n8724), .S0(g35), .Y(n4230));
NOR2X1   g4079(.A(n6024_1), .B(n5720), .Y(n8726));
NOR3X1   g4080(.A(n8726), .B(n6023), .C(n8468), .Y(n8727));
NOR4X1   g4081(.A(n6023), .B(g4601), .C(n5720), .D(n6024_1), .Y(n8728));
OR2X1    g4082(.A(n8728), .B(n8727), .Y(n8729));
MX2X1    g4083(.A(g4593), .B(n8729), .S0(g35), .Y(n4235));
INVX1    g4084(.A(g854), .Y(n8731));
XOR2X1   g4085(.A(g392), .B(g405), .Y(n8732));
NAND3X1  g4086(.A(g392), .B(g405), .C(g401), .Y(n8733));
INVX1    g4087(.A(g392), .Y(n8734));
NAND2X1  g4088(.A(g424), .B(n8734), .Y(n8735));
OAI21X1  g4089(.A0(n8735), .A1(g405), .B0(n8733), .Y(n8736));
AOI21X1  g4090(.A0(n8732), .A1(g437), .B0(n8736), .Y(n8737));
XOR2X1   g4091(.A(n8737), .B(g417), .Y(n8738));
MX2X1    g4092(.A(g174), .B(g452), .S0(g392), .Y(n8739));
NOR2X1   g4093(.A(n8739), .B(g182), .Y(n8740));
AND2X1   g4094(.A(n8739), .B(g182), .Y(n8741));
AND2X1   g4095(.A(g411), .B(n8734), .Y(n8742));
NAND2X1  g4096(.A(g392), .B(g441), .Y(n8743));
NAND3X1  g4097(.A(n8743), .B(n5516_1), .C(n6385), .Y(n8744));
NOR4X1   g4098(.A(n8742), .B(n8741), .C(n8740), .D(n8744), .Y(n8745));
NOR2X1   g4099(.A(n8745), .B(n8738), .Y(n8746));
NOR4X1   g4100(.A(n5599), .B(n5687), .C(n6177), .D(g385), .Y(n8747));
MX2X1    g4101(.A(n8731), .B(n8746), .S0(n8747), .Y(n8748));
NOR2X1   g4102(.A(n8748), .B(n4620), .Y(n4240));
INVX1    g4103(.A(g1442), .Y(n8750));
INVX1    g4104(.A(g1489), .Y(n8751));
XOR2X1   g4105(.A(n6519), .B(g1300), .Y(n8752));
NAND3X1  g4106(.A(n8752), .B(n8751), .C(n8750), .Y(n8753));
NAND3X1  g4107(.A(n8752), .B(n6521), .C(g1484), .Y(n8754));
NAND2X1  g4108(.A(n8754), .B(n8753), .Y(n8755));
MX2X1    g4109(.A(g1484), .B(n8755), .S0(n6514), .Y(n8756));
MX2X1    g4110(.A(g1472), .B(n8756), .S0(g35), .Y(n4245));
MX2X1    g4111(.A(g4922), .B(n6676), .S0(n6891_1), .Y(n8758));
MX2X1    g4112(.A(g4917), .B(n8758), .S0(g35), .Y(n4250));
INVX1    g4113(.A(g5077), .Y(n8760));
NOR2X1   g4114(.A(g5073), .B(n8760), .Y(n8761));
NOR2X1   g4115(.A(g5069), .B(n8760), .Y(n8762));
MX2X1    g4116(.A(n8761), .B(n8762), .S0(g5084), .Y(n8763));
MX2X1    g4117(.A(g5077), .B(n8763), .S0(g35), .Y(n4255));
NAND2X1  g4118(.A(n7375), .B(g5863), .Y(n8765));
NAND2X1  g4119(.A(g5857), .B(n6653_1), .Y(n8766));
AOI21X1  g4120(.A0(n8766), .A1(n8765), .B0(n7540_1), .Y(n8767));
MX2X1    g4121(.A(g5857), .B(n8767), .S0(g35), .Y(n4260));
INVX1    g4122(.A(g4462), .Y(n8769));
OR2X1    g4123(.A(g4473), .B(n4620), .Y(n8770));
OAI22X1  g4124(.A0(n8769), .A1(g35), .B0(g4467), .B1(n8770), .Y(n4265));
NOR3X1   g4125(.A(n6588), .B(n5573_1), .C(n5585), .Y(n8772));
NOR3X1   g4126(.A(g3004), .B(n6593), .C(g3017), .Y(n8773));
OAI21X1  g4127(.A0(n8773), .A1(n8772), .B0(n6587), .Y(n8774));
NOR2X1   g4128(.A(n8773), .B(n8772), .Y(n8775));
NAND2X1  g4129(.A(n8775), .B(g3021), .Y(n8776));
OAI21X1  g4130(.A0(n8776), .A1(n5584), .B0(n8774), .Y(n8777));
MX2X1    g4131(.A(g3017), .B(n8777), .S0(g35), .Y(n4270));
INVX1    g4132(.A(g2518), .Y(n8779));
AOI21X1  g4133(.A0(n5562), .A1(g2476), .B0(n8779), .Y(n8780));
XOR2X1   g4134(.A(n8780), .B(g2504), .Y(n8781));
MX2X1    g4135(.A(g2518), .B(n8781), .S0(n6444_1), .Y(n8782));
MX2X1    g4136(.A(g2504), .B(n8782), .S0(g35), .Y(n4275));
MX2X1    g4137(.A(g2567), .B(n5998), .S0(n8533), .Y(n8785));
MX2X1    g4138(.A(g2648), .B(n8785), .S0(g35), .Y(n4280));
NOR3X1   g4139(.A(n6134), .B(n6132_1), .C(n5262), .Y(n8787));
AOI21X1  g4140(.A0(g640), .A1(n6133), .B0(n5440_1), .Y(n8788));
MX2X1    g4141(.A(n8788), .B(n5440_1), .S0(n8787), .Y(n8789));
MX2X1    g4142(.A(g562), .B(n8789), .S0(g35), .Y(n4285));
MX2X1    g4143(.A(g3263), .B(n5592_1), .S0(n4846_1), .Y(n8792));
MX2X1    g4144(.A(g3259), .B(n8792), .S0(g35), .Y(n4290));
NOR4X1   g4145(.A(g6573), .B(g6555), .C(n7524), .D(n4855), .Y(n8794));
MX2X1    g4146(.A(g6613), .B(n5592_1), .S0(n8794), .Y(n8795));
MX2X1    g4147(.A(g6585), .B(n8795), .S0(g35), .Y(n4295));
AOI21X1  g4148(.A0(n8071), .A1(g35), .B0(n8431), .Y(n4300));
INVX1    g4149(.A(g6494), .Y(n8798));
AOI21X1  g4150(.A0(g6486), .A1(n8798), .B0(g6444), .Y(n8799));
OR2X1    g4151(.A(g6490), .B(n4620), .Y(n8800));
OAI22X1  g4152(.A0(n8799), .A1(n8800), .B0(n8798), .B1(g35), .Y(n4305));
AND2X1   g4153(.A(n7587), .B(n6708), .Y(n8802));
INVX1    g4154(.A(g91), .Y(n8803));
OR4X1    g4155(.A(n4658), .B(g2965), .C(n8803), .D(n4661), .Y(n8804));
NAND2X1  g4156(.A(n8804), .B(g35), .Y(n8805));
OAI22X1  g4157(.A0(n8802), .A1(n8805), .B0(n5370_1), .B1(g35), .Y(n4310));
NOR4X1   g4158(.A(g5857), .B(g5869), .C(n4620), .D(n7540_1), .Y(n4315));
NOR2X1   g4159(.A(n6500), .B(n5758_1), .Y(n8808));
MX2X1    g4160(.A(g1616), .B(n5756), .S0(n8808), .Y(n8809));
MX2X1    g4161(.A(g1620), .B(n8809), .S0(g35), .Y(n4320));
INVX1    g4162(.A(n8747), .Y(n8811));
NOR3X1   g4163(.A(n8811), .B(n8746), .C(g703), .Y(n8812));
INVX1    g4164(.A(g862), .Y(n8813));
OR2X1    g4165(.A(n6178_1), .B(n8813), .Y(n8814));
MX2X1    g4166(.A(n8813), .B(n4882), .S0(g896), .Y(n8815));
OAI21X1  g4167(.A0(n8814), .A1(n8812), .B0(n8815), .Y(n8816));
MX2X1    g4168(.A(g446), .B(n8816), .S0(g35), .Y(n4325));
NOR3X1   g4169(.A(g3522), .B(n4834), .C(n4833), .Y(n8818));
MX2X1    g4170(.A(g3562), .B(n5592_1), .S0(n8818), .Y(n8819));
MX2X1    g4171(.A(g3606), .B(n8819), .S0(g35), .Y(n4334));
INVX1    g4172(.A(g4239), .Y(n8821));
OR2X1    g4173(.A(g4294), .B(n4620), .Y(n8822));
OAI22X1  g4174(.A0(n8821), .A1(g35), .B0(g4297), .B1(n8822), .Y(n4339));
INVX1    g4175(.A(g1395), .Y(n8824));
INVX1    g4176(.A(g1570), .Y(n8825));
NOR3X1   g4177(.A(g1399), .B(g1333), .C(g1500), .Y(n8826));
NOR3X1   g4178(.A(n8826), .B(n8825), .C(n8824), .Y(n8827));
NOR2X1   g4179(.A(n8827), .B(g1404), .Y(n8828));
INVX1    g4180(.A(g1404), .Y(n8829));
OR4X1    g4181(.A(n8825), .B(n8824), .C(n8829), .D(n8826), .Y(n8830));
NOR2X1   g4182(.A(g1322), .B(n4620), .Y(n8831));
NAND2X1  g4183(.A(n8831), .B(n8830), .Y(n8832));
OAI22X1  g4184(.A0(n8828), .A1(n8832), .B0(n8824), .B1(g35), .Y(n4343));
NOR3X1   g4185(.A(n7353), .B(n7352_1), .C(n7351), .Y(n8834));
NOR3X1   g4186(.A(g3706), .B(g3719), .C(n7359), .Y(n8835));
OAI21X1  g4187(.A0(n8835), .A1(n8834), .B0(n7354), .Y(n8836));
NOR2X1   g4188(.A(n8835), .B(n8834), .Y(n8837));
NAND2X1  g4189(.A(n8837), .B(g3723), .Y(n8838));
OAI21X1  g4190(.A0(n8838), .A1(n7371), .B0(n8836), .Y(n8839));
MX2X1    g4191(.A(g3719), .B(n8839), .S0(g35), .Y(n4348));
XOR2X1   g4192(.A(g3808), .B(g3813), .Y(n8841));
MX2X1    g4193(.A(g3817), .B(n8841), .S0(n7137_1), .Y(n8842));
MX2X1    g4194(.A(g3808), .B(n8842), .S0(g35), .Y(n4353));
OR2X1    g4195(.A(n5189), .B(n5180), .Y(n8844));
OAI21X1  g4196(.A0(n5198), .A1(n8844), .B0(n4958), .Y(n8845));
OAI21X1  g4197(.A0(n5199), .A1(n4958), .B0(n8845), .Y(n4358));
NAND3X1  g4198(.A(n7113_1), .B(n4953), .C(g72), .Y(n8847));
MX2X1    g4199(.A(g4498), .B(n8847), .S0(g4581), .Y(n8848));
MX2X1    g4200(.A(g4498), .B(n8848), .S0(g35), .Y(n4363));
NOR4X1   g4201(.A(n5661), .B(n5516_1), .C(n6115), .D(n6113), .Y(n8850));
MX2X1    g4202(.A(n6115), .B(n8850), .S0(n6114_1), .Y(n8851));
MX2X1    g4203(.A(g283), .B(n8851), .S0(g35), .Y(n4368));
XOR2X1   g4204(.A(n5862), .B(n6898), .Y(n8853));
NAND2X1  g4205(.A(g2841), .B(g35), .Y(n8854));
OAI22X1  g4206(.A0(n8853), .A1(n8854), .B0(n6307), .B1(g35), .Y(n4373));
INVX1    g4207(.A(g4704), .Y(n8856));
OR2X1    g4208(.A(g28753), .B(n8856), .Y(n8857));
NAND3X1  g4209(.A(g5348), .B(n6340), .C(g5297), .Y(n8858));
INVX1    g4210(.A(g5348), .Y(n8859));
NAND2X1  g4211(.A(n6348), .B(n8859), .Y(n8860));
INVX1    g4212(.A(g5352), .Y(n8861));
MX2X1    g4213(.A(n5173), .B(n6334), .S0(n8861), .Y(n8862));
NAND4X1  g4214(.A(n8860), .B(n8858), .C(n8856), .D(n8862), .Y(n8863));
NAND4X1  g4215(.A(n4970), .B(n4820), .C(g28753), .D(n8863), .Y(n8864));
AOI21X1  g4216(.A0(n8864), .A1(n8857), .B0(n4620), .Y(n4378));
NOR2X1   g4217(.A(n6668), .B(n5217), .Y(n8866));
OAI21X1  g4218(.A0(g2878), .A1(n8803), .B0(g35), .Y(n8867));
OAI22X1  g4219(.A0(n8866), .A1(n8867), .B0(n5374), .B1(g35), .Y(n4388));
NOR3X1   g4220(.A(n4644), .B(n4643), .C(g5180), .Y(n8869));
MX2X1    g4221(.A(g5220), .B(n5592_1), .S0(n8869), .Y(n8870));
MX2X1    g4222(.A(g5264), .B(n8870), .S0(g35), .Y(n4393));
MX2X1    g4223(.A(n6285), .B(n5345_1), .S0(n6284), .Y(n8872));
MX2X1    g4224(.A(g613), .B(n8872), .S0(g35), .Y(n4398));
AND2X1   g4225(.A(g64), .B(g35), .Y(n4403));
MX2X1    g4226(.A(g324), .B(n8036), .S0(g35), .Y(n4407));
INVX1    g4227(.A(g1274), .Y(n8876));
NAND3X1  g4228(.A(n7801), .B(g1270), .C(g1263), .Y(n8877));
OR4X1    g4229(.A(n4713), .B(n8876), .C(n4620), .D(n8877), .Y(n8878));
OAI21X1  g4230(.A0(n8876), .A1(g35), .B0(n8878), .Y(n4412));
XOR2X1   g4231(.A(n4857), .B(g6513), .Y(n8880));
MX2X1    g4232(.A(g6509), .B(n8880), .S0(g35), .Y(n4417));
MX2X1    g4233(.A(g336), .B(g305), .S0(n8036), .Y(n8882));
MX2X1    g4234(.A(g311), .B(n8882), .S0(g35), .Y(n4422));
NOR3X1   g4235(.A(n5462), .B(n5217), .C(n5616), .Y(n8884));
NOR3X1   g4236(.A(n4661), .B(n4658), .C(g2882), .Y(n8885));
OR2X1    g4237(.A(n8885), .B(n4620), .Y(n8886));
OAI22X1  g4238(.A0(n8884), .A1(n8886), .B0(n5341), .B1(g35), .Y(n4427));
INVX1    g4239(.A(g930), .Y(n8888));
NAND3X1  g4240(.A(n6454), .B(g918), .C(g925), .Y(n8889));
OR4X1    g4241(.A(n4709), .B(n8888), .C(n4620), .D(n8889), .Y(n8890));
OAI21X1  g4242(.A0(n8888), .A1(g35), .B0(n8890), .Y(n4432));
INVX1    g4243(.A(g1906), .Y(n8892));
NAND3X1  g4244(.A(n6223), .B(n6222), .C(g1862), .Y(n8893));
OAI21X1  g4245(.A0(n6222), .A1(n8892), .B0(n8893), .Y(n8894));
MX2X1    g4246(.A(g1913), .B(n8894), .S0(g35), .Y(n4437));
AND2X1   g4247(.A(g6745), .B(g35), .Y(n4442));
MX2X1    g4248(.A(g3361), .B(g3401), .S0(g3355), .Y(n8897));
OR2X1    g4249(.A(n8897), .B(n6411), .Y(n8898));
NAND2X1  g4250(.A(n8897), .B(n6411), .Y(n8899));
OAI21X1  g4251(.A0(n8898), .A1(n5778_1), .B0(n8899), .Y(n8900));
MX2X1    g4252(.A(g3355), .B(n8900), .S0(g35), .Y(n4452));
INVX1    g4253(.A(g2193), .Y(n8902));
AOI21X1  g4254(.A0(n7859), .A1(n8902), .B0(g2799), .Y(n8903));
NAND2X1  g4255(.A(g121), .B(n4620), .Y(n8904));
OAI21X1  g4256(.A0(n8903), .A1(n7861), .B0(n8904), .Y(n4457));
MX2X1    g4257(.A(g4912), .B(n3393), .S0(n6891_1), .Y(n8906));
MX2X1    g4258(.A(g4907), .B(n8906), .S0(g35), .Y(n4469));
MX2X1    g4259(.A(g4157), .B(n3220), .S0(n5697), .Y(n8908));
MX2X1    g4260(.A(g4146), .B(n8908), .S0(g35), .Y(n4474));
XOR2X1   g4261(.A(n7133), .B(g2541), .Y(n8910));
MX2X1    g4262(.A(g2537), .B(n8910), .S0(g35), .Y(n4479));
NAND3X1  g4263(.A(n6707), .B(n6702), .C(g2153), .Y(n8912));
NAND4X1  g4264(.A(n5637), .B(g112), .C(n4824), .D(n5135_1), .Y(n8913));
AOI21X1  g4265(.A0(g2197), .A1(n6708_1), .B0(g2227), .Y(n8914));
NAND3X1  g4266(.A(n8914), .B(n8913), .C(n7512), .Y(n8915));
AOI21X1  g4267(.A0(n8915), .A1(n8912), .B0(n4620), .Y(n4484));
AND2X1   g4268(.A(n7912), .B(n6708), .Y(n8917));
INVX1    g4269(.A(g79), .Y(n8918));
OAI21X1  g4270(.A0(n8918), .A1(g550), .B0(g35), .Y(n8919));
OAI22X1  g4271(.A0(n8917), .A1(n8919), .B0(n5387), .B1(g35), .Y(n4489));
MX2X1    g4272(.A(g255), .B(g869), .S0(n7408), .Y(n8921));
MX2X1    g4273(.A(g225), .B(n8921), .S0(g35), .Y(n4494));
NAND3X1  g4274(.A(n5838), .B(n4939_1), .C(g1882), .Y(n8923));
NAND3X1  g4275(.A(g1870), .B(n5838), .C(g1917), .Y(n8924));
AND2X1   g4276(.A(n8924), .B(n8923), .Y(n8925));
AND2X1   g4277(.A(g1894), .B(g1926), .Y(n8926));
NOR2X1   g4278(.A(g1917), .B(n4939_1), .Y(n8927));
AOI22X1  g4279(.A0(n8926), .A1(g1874), .B0(g1878), .B1(n8927), .Y(n8928));
NAND3X1  g4280(.A(g1890), .B(g1917), .C(n4939_1), .Y(n8929));
NAND3X1  g4281(.A(g1886), .B(g1894), .C(n6203), .Y(n8930));
NAND4X1  g4282(.A(n8929), .B(n8928), .C(n8925), .D(n8930), .Y(n8931));
MX2X1    g4283(.A(g1945), .B(n8931), .S0(n6202), .Y(n8932));
MX2X1    g4284(.A(g1926), .B(n8932), .S0(g35), .Y(n4499));
NOR3X1   g4285(.A(n6195), .B(n6624), .C(g5164), .Y(n8934));
MX2X1    g4286(.A(g5240), .B(n5592_1), .S0(n8934), .Y(n8935));
MX2X1    g4287(.A(g5224), .B(n8935), .S0(g35), .Y(n4504));
NOR4X1   g4288(.A(n5549), .B(g1526), .C(n6513), .D(n7603), .Y(n8937));
XOR2X1   g4289(.A(g1478), .B(g1437), .Y(n8938));
MX2X1    g4290(.A(g1478), .B(n8938), .S0(n8937), .Y(n8939));
MX2X1    g4291(.A(g1437), .B(n8939), .S0(g35), .Y(n4509));
XOR2X1   g4292(.A(g3072), .B(g3080), .Y(n8941));
MX2X1    g4293(.A(g3072), .B(n8941), .S0(g35), .Y(n4514));
NAND2X1  g4294(.A(n7642), .B(g3863), .Y(n8943));
NAND2X1  g4295(.A(g3857), .B(n7041), .Y(n8944));
AOI21X1  g4296(.A0(n8944), .A1(n8943), .B0(n7849), .Y(n8945));
MX2X1    g4297(.A(g3857), .B(n8945), .S0(g35), .Y(n4519));
INVX1    g4298(.A(g1945), .Y(n8947));
OAI21X1  g4299(.A0(g1894), .A1(n6203), .B0(g1959), .Y(n8948));
XOR2X1   g4300(.A(n8948), .B(n8947), .Y(n8949));
MX2X1    g4301(.A(g1959), .B(n8949), .S0(n6202), .Y(n8950));
MX2X1    g4302(.A(g1945), .B(n8950), .S0(g35), .Y(n4524));
INVX1    g4303(.A(g3476), .Y(n8952));
XOR2X1   g4304(.A(g3470), .B(n8952), .Y(n8953));
MX2X1    g4305(.A(g3480), .B(n8953), .S0(n7393), .Y(n8954));
MX2X1    g4306(.A(g3476), .B(n8954), .S0(g35), .Y(n4529));
NOR3X1   g4307(.A(n7205), .B(n7204), .C(n7524), .Y(n8956));
MX2X1    g4308(.A(g6653), .B(n5592_1), .S0(n8956), .Y(n8957));
MX2X1    g4309(.A(g6637), .B(n8957), .S0(g35), .Y(n4534));
NOR3X1   g4310(.A(n5465), .B(n5217), .C(n5616), .Y(n8959));
OAI21X1  g4311(.A0(n4744), .A1(g2864), .B0(g35), .Y(n8960));
NAND2X1  g4312(.A(g2856), .B(n4620), .Y(n8961));
OAI21X1  g4313(.A0(n8960), .A1(n8959), .B0(n8961), .Y(n4544));
INVX1    g4314(.A(g4894), .Y(n8963));
OR2X1    g4315(.A(n7721), .B(n8963), .Y(n8964));
OAI21X1  g4316(.A0(n8576), .A1(n8536), .B0(n8963), .Y(n8965));
NAND2X1  g4317(.A(n8583), .B(n8536), .Y(n8966));
INVX1    g4318(.A(g6736), .Y(n8967));
NAND3X1  g4319(.A(g6741), .B(n8569), .C(n8967), .Y(n8968));
NAND3X1  g4320(.A(g6741), .B(g6682), .C(g6736), .Y(n8969));
NAND3X1  g4321(.A(n8969), .B(n8968), .C(n8966), .Y(n8970));
OR2X1    g4322(.A(n8970), .B(n8965), .Y(n8971));
NAND4X1  g4323(.A(n7721), .B(n4964_1), .C(n4898), .D(n8971), .Y(n8972));
AOI21X1  g4324(.A0(n8972), .A1(n8964), .B0(n4620), .Y(n4549));
NOR4X1   g4325(.A(g3857), .B(g3869), .C(n4620), .D(n7849), .Y(n4558));
OAI21X1  g4326(.A0(g686), .A1(n5876), .B0(g518), .Y(n8975));
AOI21X1  g4327(.A0(g499), .A1(n7004), .B0(n8975), .Y(n8976));
MX2X1    g4328(.A(n6234), .B(n8976), .S0(n5880_1), .Y(n8977));
NOR2X1   g4329(.A(n8977), .B(n4620), .Y(n4566));
INVX1    g4330(.A(g5401), .Y(n8979));
NAND3X1  g4331(.A(n6645), .B(n6644), .C(g35), .Y(n8980));
OAI21X1  g4332(.A0(n8979), .A1(g35), .B0(n8980), .Y(n4571));
MX2X1    g4333(.A(g1002), .B(n7502), .S0(n6059), .Y(n8982));
MX2X1    g4334(.A(g1008), .B(n8982), .S0(g35), .Y(n4576));
AOI21X1  g4335(.A0(g802), .A1(n5662), .B0(n5231_1), .Y(n8984));
MX2X1    g4336(.A(n5231_1), .B(n8984), .S0(n5679_1), .Y(n8985));
MX2X1    g4337(.A(g772), .B(n8985), .S0(g35), .Y(n4581));
NAND4X1  g4338(.A(n6744), .B(n7014), .C(g35), .D(n4719), .Y(n8987));
NOR3X1   g4339(.A(n8987), .B(n6216_1), .C(n4968), .Y(n4595));
OAI21X1  g4340(.A0(n6204), .A1(n4917), .B0(n5562), .Y(n8989));
MX2X1    g4341(.A(g2476), .B(n8989), .S0(n6444_1), .Y(n8990));
MX2X1    g4342(.A(g2453), .B(n8990), .S0(g35), .Y(n4600));
NOR2X1   g4343(.A(n6501), .B(n5787_1), .Y(n8992));
OAI21X1  g4344(.A0(n6204), .A1(n4922), .B0(n4629), .Y(n8993));
MX2X1    g4345(.A(g1657), .B(n8993), .S0(n8992), .Y(n8994));
MX2X1    g4346(.A(g1664), .B(n8994), .S0(g35), .Y(n4605));
NOR2X1   g4347(.A(n5542), .B(n5524), .Y(n8996));
MX2X1    g4348(.A(n8996), .B(g1589), .S0(n5545), .Y(n8997));
OAI21X1  g4349(.A0(g2361), .A1(g2287), .B0(g2375), .Y(n8998));
XOR2X1   g4350(.A(n8998), .B(n8997), .Y(n8999));
MX2X1    g4351(.A(n8999), .B(g2375), .S0(n5552), .Y(n9000));
MX2X1    g4352(.A(g2361), .B(n9000), .S0(g35), .Y(n4610));
OAI21X1  g4353(.A0(n4972), .A1(n4966), .B0(n4958), .Y(n9002));
OAI21X1  g4354(.A0(n4973), .A1(n4958), .B0(n9002), .Y(n4615));
XOR2X1   g4355(.A(g890), .B(n8813), .Y(n9004));
MX2X1    g4356(.A(g862), .B(n9004), .S0(g35), .Y(n4627));
NOR2X1   g4357(.A(n5278), .B(g35), .Y(n4632));
OR2X1    g4358(.A(g3423), .B(g3419), .Y(n9007));
INVX1    g4359(.A(g3412), .Y(n9008));
AOI22X1  g4360(.A0(g3423), .A1(g3419), .B0(n9008), .B1(g3416), .Y(n9009));
OAI21X1  g4361(.A0(n9007), .A1(n8218), .B0(n9009), .Y(n9010));
MX2X1    g4362(.A(g3419), .B(n9010), .S0(g35), .Y(n4637));
NAND2X1  g4363(.A(n6104), .B(g35), .Y(n9012));
OR4X1    g4364(.A(n6113), .B(n5661), .C(n5516_1), .D(n9012), .Y(n9013));
OAI21X1  g4365(.A0(n6322), .A1(g35), .B0(n9013), .Y(n4642));
NAND2X1  g4366(.A(g3161), .B(n5913), .Y(n9015));
NAND2X1  g4367(.A(n5593), .B(g3155), .Y(n9016));
AOI21X1  g4368(.A0(n9016), .A1(n9015), .B0(n5765), .Y(n9017));
MX2X1    g4369(.A(g3155), .B(n9017), .S0(g35), .Y(n4647));
INVX1    g4370(.A(g2384), .Y(n9019));
AOI21X1  g4371(.A0(n7228), .A1(g2342), .B0(n9019), .Y(n9020));
XOR2X1   g4372(.A(n9020), .B(g2370), .Y(n9021));
MX2X1    g4373(.A(g2384), .B(n9021), .S0(n7227), .Y(n9022));
MX2X1    g4374(.A(g2370), .B(n9022), .S0(g35), .Y(n4652));
INVX1    g4375(.A(g3454), .Y(n9024));
AOI21X1  g4376(.A0(g3447), .A1(n9024), .B0(g3361), .Y(n9025));
OR2X1    g4377(.A(g3443), .B(n4620), .Y(n9026));
OAI22X1  g4378(.A0(n9025), .A1(n9026), .B0(n9024), .B1(g35), .Y(n4657));
NOR4X1   g4379(.A(n8468), .B(n5716), .C(n5720), .D(n6024_1), .Y(n9028));
INVX1    g4380(.A(g4616), .Y(n9029));
NOR2X1   g4381(.A(n6023), .B(n9029), .Y(n9030));
NOR2X1   g4382(.A(n6023), .B(g4616), .Y(n9031));
MX2X1    g4383(.A(n9030), .B(n9031), .S0(n9028), .Y(n9032));
MX2X1    g4384(.A(g4608), .B(n9032), .S0(g35), .Y(n4667));
MX2X1    g4385(.A(g4558), .B(g6749), .S0(g35), .Y(n4672));
NOR3X1   g4386(.A(n6085), .B(n5166_1), .C(g2040), .Y(n9035));
MX2X1    g4387(.A(g2024), .B(n7037_1), .S0(n9035), .Y(n9036));
MX2X1    g4388(.A(g2012), .B(n9036), .S0(g35), .Y(n4677));
INVX1    g4389(.A(g2036), .Y(n9038));
AOI21X1  g4390(.A0(n7859), .A1(n9038), .B0(g2795), .Y(n9039));
OAI22X1  g4391(.A0(n7861), .A1(n9039), .B0(n7313), .B1(g35), .Y(n4687));
NOR3X1   g4392(.A(n6143), .B(n6134), .C(n5349), .Y(n9041));
AOI21X1  g4393(.A0(g640), .A1(n6133), .B0(n5322_1), .Y(n9042));
NAND3X1  g4394(.A(n6497), .B(n9042), .C(n9041), .Y(n9043));
OR4X1    g4395(.A(n6134), .B(n5228), .C(n5258), .D(n9043), .Y(n9044));
OR4X1    g4396(.A(n6134), .B(n5436), .C(n5406), .D(n9044), .Y(n9045));
AOI21X1  g4397(.A0(g640), .A1(n6133), .B0(n5381), .Y(n9046));
MX2X1    g4398(.A(n5381), .B(n9046), .S0(n9045), .Y(n9047));
MX2X1    g4399(.A(g608), .B(n9047), .S0(g35), .Y(n4692));
NAND4X1  g4400(.A(g4489), .B(g4486), .C(g4492), .D(g4483), .Y(n9049));
INVX1    g4401(.A(n9049), .Y(n9050));
XOR2X1   g4402(.A(n9050), .B(g4527), .Y(n9051));
MX2X1    g4403(.A(n5724), .B(n9051), .S0(g4521), .Y(n9052));
MX2X1    g4404(.A(g4521), .B(n9052), .S0(g35), .Y(n4697));
INVX1    g4405(.A(g1840), .Y(n9054));
XOR2X1   g4406(.A(g1834), .B(n9054), .Y(n9055));
MX2X1    g4407(.A(g1844), .B(n9055), .S0(n8442), .Y(n9056));
MX2X1    g4408(.A(g1840), .B(n9056), .S0(g35), .Y(n4702));
NOR4X1   g4409(.A(n6653_1), .B(g5881), .C(n4860), .D(g5857), .Y(n9058));
MX2X1    g4410(.A(g5937), .B(n5592_1), .S0(n9058), .Y(n9059));
MX2X1    g4411(.A(g5921), .B(n9059), .S0(g35), .Y(n4707));
NAND3X1  g4412(.A(n6835_1), .B(n4953), .C(g72), .Y(n9061));
MX2X1    g4413(.A(g4567), .B(n9061), .S0(g4581), .Y(n9062));
MX2X1    g4414(.A(g4567), .B(n9062), .S0(g35), .Y(n4712));
XOR2X1   g4415(.A(g2518), .B(g2514), .Y(n9064));
NOR4X1   g4416(.A(n5567), .B(g2453), .C(n6445), .D(n5569), .Y(n9065));
MX2X1    g4417(.A(g2523), .B(n9064), .S0(n9065), .Y(n9066));
MX2X1    g4418(.A(g2518), .B(n9066), .S0(g35), .Y(n4722));
INVX1    g4419(.A(g3267), .Y(n9068));
OAI22X1  g4420(.A0(g3310), .A1(n9068), .B0(g3303), .B1(n6825_1), .Y(n9069));
MX2X1    g4421(.A(g3298), .B(n9068), .S0(g3274), .Y(n9070));
OAI21X1  g4422(.A0(n6826), .A1(g3281), .B0(g35), .Y(n9071));
NOR4X1   g4423(.A(n9070), .B(n9069), .C(n8057), .D(n9071), .Y(n4727));
NOR2X1   g4424(.A(n5993), .B(n5524), .Y(n9073));
MX2X1    g4425(.A(n9073), .B(g1589), .S0(n5995), .Y(n9074));
OAI21X1  g4426(.A0(g2555), .A1(g2629), .B0(g2643), .Y(n9075));
XOR2X1   g4427(.A(n9075), .B(n9074), .Y(n9076));
MX2X1    g4428(.A(n9076), .B(g2643), .S0(n6003), .Y(n9077));
MX2X1    g4429(.A(g2629), .B(n9077), .S0(g35), .Y(n4731));
MX2X1    g4430(.A(g6105), .B(n5816_1), .S0(g35), .Y(n4736));
AOI21X1  g4431(.A0(g1489), .A1(n7602), .B0(n8750), .Y(n9080));
MX2X1    g4432(.A(n8751), .B(n9080), .S0(n6514), .Y(n9081));
NOR2X1   g4433(.A(n9081), .B(n4620), .Y(n4741));
AND2X1   g4434(.A(n8405), .B(n8403), .Y(n9083));
NOR2X1   g4435(.A(n6646), .B(n6638_1), .Y(n9084));
MX2X1    g4436(.A(n6638_1), .B(n9084), .S0(n9083), .Y(n9085));
MX2X1    g4437(.A(g5385), .B(n9085), .S0(g35), .Y(n4746));
INVX1    g4438(.A(g191), .Y(n9087));
AND2X1   g4439(.A(g218), .B(g215), .Y(n9088));
MX2X1    g4440(.A(g194), .B(n9087), .S0(n9088), .Y(n9089));
MX2X1    g4441(.A(g222), .B(n9089), .S0(g35), .Y(n4751));
INVX1    g4442(.A(g2547), .Y(n9091));
XOR2X1   g4443(.A(g2541), .B(n9091), .Y(n9092));
MX2X1    g4444(.A(g2551), .B(n9092), .S0(n5570), .Y(n9093));
MX2X1    g4445(.A(g2547), .B(n9093), .S0(g35), .Y(n4756));
INVX1    g4446(.A(g5156), .Y(n9095));
OAI22X1  g4447(.A0(n5524), .A1(g4284), .B0(n9095), .B1(g26801), .Y(n9096));
OR4X1    g4448(.A(n5524), .B(g4284), .C(n9095), .D(g26801), .Y(n9097));
AOI21X1  g4449(.A0(n9097), .A1(n9096), .B0(n4620), .Y(n4761));
INVX1    g4450(.A(g3065), .Y(n9099));
NOR2X1   g4451(.A(n9099), .B(g3057), .Y(n9100));
OR2X1    g4452(.A(g3068), .B(g3072), .Y(n9101));
INVX1    g4453(.A(g3061), .Y(n9102));
AOI22X1  g4454(.A0(g3068), .A1(g3072), .B0(g3065), .B1(n9102), .Y(n9103));
OAI21X1  g4455(.A0(n9101), .A1(n9100), .B0(n9103), .Y(n9104));
MX2X1    g4456(.A(g3068), .B(n9104), .S0(g35), .Y(n4766));
AOI21X1  g4457(.A0(n5337), .A1(n5317), .B0(g22), .Y(n9106));
AOI21X1  g4458(.A0(n5337), .A1(n5317), .B0(n5282), .Y(n9107));
OR2X1    g4459(.A(n9107), .B(n9106), .Y(n4775));
AND2X1   g4460(.A(g3530), .B(g35), .Y(n4780));
OR2X1    g4461(.A(g4281), .B(n4620), .Y(n9110));
OAI21X1  g4462(.A0(n5271), .A1(g35), .B0(n9110), .Y(n4784));
NOR3X1   g4463(.A(n5531_1), .B(g1936), .C(g1862), .Y(n9112));
MX2X1    g4464(.A(g1955), .B(g1950), .S0(n9112), .Y(n9113));
MX2X1    g4465(.A(g1950), .B(n9113), .S0(g35), .Y(n4788));
NAND3X1  g4466(.A(n7699), .B(n6746), .C(n6951), .Y(n9115));
OAI21X1  g4467(.A0(n6746), .A1(n6951), .B0(n9115), .Y(n9116));
MX2X1    g4468(.A(g6044), .B(n9116), .S0(g35), .Y(n4793));
AND2X1   g4469(.A(n6595_1), .B(n6590_1), .Y(n9118));
NOR2X1   g4470(.A(n5584), .B(n5576), .Y(n9119));
MX2X1    g4471(.A(n5576), .B(n9119), .S0(n9118), .Y(n9120));
MX2X1    g4472(.A(g3029), .B(n9120), .S0(g35), .Y(n4798));
NOR3X1   g4473(.A(n7511_1), .B(g2227), .C(g2153), .Y(n9122));
XOR2X1   g4474(.A(n9122), .B(g2273), .Y(n9123));
MX2X1    g4475(.A(g2269), .B(n9123), .S0(g35), .Y(n4803));
INVX1    g4476(.A(g4771), .Y(n9125));
OR2X1    g4477(.A(n5907), .B(n9125), .Y(n9126));
INVX1    g4478(.A(g6386), .Y(n9127));
OAI21X1  g4479(.A0(n6532), .A1(n9127), .B0(n9125), .Y(n9128));
NAND2X1  g4480(.A(n6539), .B(n9127), .Y(n9129));
NAND3X1  g4481(.A(n7000), .B(g6395), .C(n6279), .Y(n9130));
NAND3X1  g4482(.A(g6390), .B(g6395), .C(g6336), .Y(n9131));
NAND3X1  g4483(.A(n9131), .B(n9130), .C(n9129), .Y(n9132));
OR2X1    g4484(.A(n9132), .B(n9128), .Y(n9133));
NAND4X1  g4485(.A(n5907), .B(n4970), .C(n7428), .D(n9133), .Y(n9134));
AOI21X1  g4486(.A0(n9134), .A1(n9126), .B0(n4620), .Y(n4812));
INVX1    g4487(.A(g6148), .Y(n9136));
AOI21X1  g4488(.A0(g6140), .A1(n9136), .B0(g6098), .Y(n9137));
OR2X1    g4489(.A(g6144), .B(n4620), .Y(n9138));
OAI22X1  g4490(.A0(n9137), .A1(n9138), .B0(n9136), .B1(g35), .Y(n4817));
INVX1    g4491(.A(g3147), .Y(n9140));
OAI22X1  g4492(.A0(n5524), .A1(g4284), .B0(n9140), .B1(n4846_1), .Y(n9141));
OR4X1    g4493(.A(n5524), .B(g4284), .C(n9140), .D(n4846_1), .Y(n9142));
AOI21X1  g4494(.A0(n9142), .A1(n9141), .B0(n4620), .Y(n4822));
INVX1    g4495(.A(g3343), .Y(n9144));
AOI21X1  g4496(.A0(n6828), .A1(g35), .B0(n9144), .Y(n4827));
INVX1    g4497(.A(g2259), .Y(n9146));
XOR2X1   g4498(.A(g2265), .B(n9146), .Y(n9147));
MX2X1    g4499(.A(g2269), .B(n9147), .S0(n9122), .Y(n9148));
MX2X1    g4500(.A(g2265), .B(n9148), .S0(g35), .Y(n4832));
INVX1    g4501(.A(g2841), .Y(n9150));
OAI22X1  g4502(.A0(g2712), .A1(n7779), .B0(n9150), .B1(g35), .Y(n4841));
NAND3X1  g4503(.A(n6287), .B(n6285), .C(n6284), .Y(n9152));
MX2X1    g4504(.A(n5292), .B(n7383), .S0(n9152), .Y(n9153));
MX2X1    g4505(.A(g622), .B(n9153), .S0(g35), .Y(n4846));
NAND3X1  g4506(.A(g2715), .B(g2719), .C(g2724), .Y(n9155));
XOR2X1   g4507(.A(n9155), .B(g2729), .Y(n9156));
NAND2X1  g4508(.A(n9156), .B(g2841), .Y(n9157));
MX2X1    g4509(.A(g2724), .B(n9157), .S0(g35), .Y(n4851));
OR2X1    g4510(.A(g28753), .B(n6340), .Y(n9159));
NAND2X1  g4511(.A(g28753), .B(n6340), .Y(n9160));
OAI21X1  g4512(.A0(n9160), .A1(n7782), .B0(n9159), .Y(n9161));
MX2X1    g4513(.A(g5352), .B(n9161), .S0(g35), .Y(n4856));
NOR4X1   g4514(.A(g4991), .B(n4962), .C(n4959_1), .D(n4960), .Y(n9163));
NOR3X1   g4515(.A(n4960), .B(n4962), .C(n4959_1), .Y(n9164));
NOR2X1   g4516(.A(n9164), .B(n6802), .Y(n9165));
OAI21X1  g4517(.A0(n9165), .A1(n9163), .B0(n6779), .Y(n9166));
NAND2X1  g4518(.A(g4983), .B(n4620), .Y(n9167));
OAI21X1  g4519(.A0(n9166), .A1(n4620), .B0(n9167), .Y(n4861));
NAND3X1  g4520(.A(n6008), .B(g4785), .C(n4815), .Y(n9169));
OAI21X1  g4521(.A0(n6009), .A1(n4818), .B0(g4709), .Y(n9170));
AOI21X1  g4522(.A0(n9170), .A1(n9169), .B0(n6216_1), .Y(n9171));
MX2X1    g4523(.A(g4785), .B(n9171), .S0(g35), .Y(n4871));
INVX1    g4524(.A(g6415), .Y(n9173));
INVX1    g4525(.A(g6411), .Y(n9174));
NOR4X1   g4526(.A(n9173), .B(n6873), .C(n6885), .D(n9174), .Y(n9175));
INVX1    g4527(.A(n9175), .Y(n9176));
NOR4X1   g4528(.A(g6411), .B(g6415), .C(g6398), .D(n6887), .Y(n9177));
INVX1    g4529(.A(n9177), .Y(n9178));
NAND3X1  g4530(.A(n9178), .B(n9176), .C(g6419), .Y(n9179));
INVX1    g4531(.A(g6419), .Y(n9180));
OAI21X1  g4532(.A0(n9177), .A1(n9175), .B0(n9180), .Y(n9181));
OAI21X1  g4533(.A0(n9179), .A1(n6884), .B0(n9181), .Y(n9182));
MX2X1    g4534(.A(g6415), .B(n9182), .S0(g35), .Y(n4876));
OAI21X1  g4535(.A0(g6058), .A1(g6098), .B0(n5823), .Y(n9184));
NAND3X1  g4536(.A(n5826_1), .B(g6052), .C(n5809), .Y(n9185));
OAI21X1  g4537(.A0(n9184), .A1(n5820), .B0(n9185), .Y(n9186));
MX2X1    g4538(.A(g6058), .B(n9186), .S0(g35), .Y(n4881));
NOR3X1   g4539(.A(n5465), .B(n5286), .C(n5616), .Y(n9188));
INVX1    g4540(.A(g44), .Y(n9189));
OR2X1    g4541(.A(g2927), .B(g2932), .Y(n9190));
OAI21X1  g4542(.A0(n9190), .A1(n9189), .B0(g35), .Y(n9191));
OAI22X1  g4543(.A0(n9188), .A1(n9191), .B0(n4787), .B1(g35), .Y(n4886));
OAI21X1  g4544(.A0(n5851), .A1(n6018), .B0(n5845_1), .Y(n9193));
NAND2X1  g4545(.A(n5845_1), .B(g4340), .Y(n9194));
MX2X1    g4546(.A(g4340), .B(n9194), .S0(n9193), .Y(n9195));
MX2X1    g4547(.A(g4643), .B(n9195), .S0(g35), .Y(n4891));
NOR4X1   g4548(.A(g5863), .B(n4862), .C(n4860), .D(n7375), .Y(n9197));
MX2X1    g4549(.A(g5929), .B(n5592_1), .S0(n9197), .Y(n9198));
MX2X1    g4550(.A(g5909), .B(n9198), .S0(g35), .Y(n4896));
MX2X1    g4551(.A(g4907), .B(n4447), .S0(n6891_1), .Y(n9200));
MX2X1    g4552(.A(g4922), .B(n9200), .S0(g35), .Y(n4901));
MX2X1    g4553(.A(g4035), .B(n8116), .S0(n6856), .Y(n9202));
MX2X1    g4554(.A(g3965), .B(n9202), .S0(g35), .Y(n4910));
XOR2X1   g4555(.A(g4291), .B(g4287), .Y(n9204));
MX2X1    g4556(.A(g4291), .B(n9204), .S0(g35), .Y(n4915));
INVX1    g4557(.A(g918), .Y(n9206));
AND2X1   g4558(.A(g918), .B(g1227), .Y(n9207));
MX2X1    g4559(.A(n9207), .B(n9206), .S0(n6454), .Y(n9208));
MX2X1    g4560(.A(g914), .B(n9208), .S0(g35), .Y(n4920));
NAND3X1  g4561(.A(g4141), .B(g4057), .C(g4064), .Y(n9210));
XOR2X1   g4562(.A(n9210), .B(g4082), .Y(n9211));
NAND2X1  g4563(.A(n9211), .B(g4169), .Y(n9212));
MX2X1    g4564(.A(g4141), .B(n9212), .S0(g35), .Y(n4925));
AND2X1   g4565(.A(g6573), .B(g35), .Y(n4930));
INVX1    g4566(.A(g2051), .Y(n9215));
NOR3X1   g4567(.A(n7090), .B(g2060), .C(n9215), .Y(n9216));
MX2X1    g4568(.A(g2036), .B(n8414), .S0(n9216), .Y(n9217));
MX2X1    g4569(.A(g2016), .B(n9217), .S0(g35), .Y(n4934));
AOI21X1  g4570(.A0(g640), .A1(n6133), .B0(n5349), .Y(n9219));
MX2X1    g4571(.A(n5349), .B(n9219), .S0(n6143), .Y(n9220));
MX2X1    g4572(.A(g586), .B(n9220), .S0(g35), .Y(n4939));
NOR3X1   g4573(.A(n5758_1), .B(g1636), .C(n4631), .Y(n9222));
MX2X1    g4574(.A(g1620), .B(n5756), .S0(n9222), .Y(n9223));
MX2X1    g4575(.A(g1608), .B(n9223), .S0(g35), .Y(n4944));
NAND2X1  g4576(.A(g1677), .B(n5568_1), .Y(n9225));
AOI21X1  g4577(.A0(g1811), .A1(g2715), .B0(g2719), .Y(n9226));
AND2X1   g4578(.A(n9226), .B(n9225), .Y(n9227));
NOR2X1   g4579(.A(g2715), .B(n8947), .Y(n9228));
NAND2X1  g4580(.A(g2079), .B(g2715), .Y(n9229));
NAND2X1  g4581(.A(n9229), .B(g2719), .Y(n9230));
NOR2X1   g4582(.A(n9230), .B(n9228), .Y(n9231));
OR2X1    g4583(.A(n9231), .B(n6305), .Y(n9232));
OAI21X1  g4584(.A0(g2775), .A1(n5568_1), .B0(n6307), .Y(n9233));
AOI21X1  g4585(.A0(n5568_1), .A1(n5505), .B0(n9233), .Y(n9234));
NOR2X1   g4586(.A(g2715), .B(g2783), .Y(n9235));
OAI21X1  g4587(.A0(n5568_1), .A1(g2787), .B0(g2719), .Y(n9236));
OAI21X1  g4588(.A0(n9236), .A1(n9235), .B0(n6305), .Y(n9237));
OAI22X1  g4589(.A0(n9234), .A1(n9237), .B0(n9232), .B1(n9227), .Y(n9238));
MX2X1    g4590(.A(g2771), .B(n9238), .S0(g35), .Y(n4949));
MX2X1    g4591(.A(g667), .B(g686), .S0(n5880_1), .Y(n9240));
MX2X1    g4592(.A(g686), .B(n9240), .S0(g35), .Y(n4954));
AND2X1   g4593(.A(g930), .B(g1227), .Y(n9242));
MX2X1    g4594(.A(n8888), .B(n9242), .S0(n8889), .Y(n9243));
MX2X1    g4595(.A(g925), .B(n9243), .S0(g35), .Y(n4959));
NOR4X1   g4596(.A(n7041), .B(g3881), .C(n4848), .D(g3857), .Y(n9245));
MX2X1    g4597(.A(g3937), .B(n5592_1), .S0(n9245), .Y(n9246));
MX2X1    g4598(.A(g3921), .B(n9246), .S0(g35), .Y(n4964));
XOR2X1   g4599(.A(g5782), .B(g5774), .Y(n9248));
MX2X1    g4600(.A(g5774), .B(n9248), .S0(g35), .Y(n4969));
OR2X1    g4601(.A(n6235), .B(g817), .Y(n9250));
NAND2X1  g4602(.A(n6235), .B(g817), .Y(n9251));
AOI21X1  g4603(.A0(n9251), .A1(n9250), .B0(n7158), .Y(n9252));
MX2X1    g4604(.A(g812), .B(n9252), .S0(g35), .Y(n4974));
NOR3X1   g4605(.A(n8825), .B(g1249), .C(n4620), .Y(n4979));
AOI21X1  g4606(.A0(g827), .A1(g832), .B0(n6247), .Y(n9255));
NAND2X1  g4607(.A(n9255), .B(n7156), .Y(n9256));
NOR2X1   g4608(.A(g837), .B(n7156), .Y(n9257));
AOI22X1  g4609(.A0(n9257), .A1(g703), .B0(n7157_1), .B1(n9255), .Y(n9258));
NAND2X1  g4610(.A(n9258), .B(n9256), .Y(n9259));
MX2X1    g4611(.A(n9259), .B(g837), .S0(n6235), .Y(n9260));
MX2X1    g4612(.A(g703), .B(n9260), .S0(g35), .Y(n4984));
AOI21X1  g4613(.A0(g640), .A1(n6133), .B0(n5258), .Y(n9262));
MX2X1    g4614(.A(n5258), .B(n9262), .S0(n6145), .Y(n9263));
MX2X1    g4615(.A(g595), .B(n9263), .S0(g35), .Y(n4992));
XOR2X1   g4616(.A(n4869), .B(g5475), .Y(n9265));
MX2X1    g4617(.A(g5471), .B(n9265), .S0(g35), .Y(n4997));
NAND2X1  g4618(.A(n5661), .B(n5654), .Y(n9267));
AOI21X1  g4619(.A0(g802), .A1(n5662), .B0(g739), .Y(n9268));
MX2X1    g4620(.A(n9268), .B(n5663), .S0(n9267), .Y(n9269));
MX2X1    g4621(.A(g736), .B(n9269), .S0(g35), .Y(n5002));
NOR3X1   g4622(.A(n6654), .B(n7375), .C(n6653_1), .Y(n9271));
MX2X1    g4623(.A(g5949), .B(n5592_1), .S0(n9271), .Y(n9272));
MX2X1    g4624(.A(g5933), .B(n9272), .S0(g35), .Y(n5007));
NOR3X1   g4625(.A(n4809), .B(n7697), .C(g113), .Y(n9274));
NAND4X1  g4626(.A(n9274), .B(n5178), .C(n4956), .D(n7721), .Y(n9275));
NOR3X1   g4627(.A(n7722), .B(n8575), .C(g6682), .Y(n9276));
AOI21X1  g4628(.A0(n7721), .A1(g6741), .B0(n8569), .Y(n9277));
OAI21X1  g4629(.A0(n9277), .A1(n9276), .B0(n9275), .Y(n9278));
NAND2X1  g4630(.A(g6741), .B(n4620), .Y(n9279));
OAI21X1  g4631(.A0(n9278), .A1(n4620), .B0(n9279), .Y(n5012));
INVX1    g4632(.A(g6093), .Y(n9281));
NAND3X1  g4633(.A(n5819), .B(n5818), .C(g35), .Y(n9282));
OAI21X1  g4634(.A0(n9281), .A1(g35), .B0(n9282), .Y(n5017));
NOR3X1   g4635(.A(g904), .B(n5691), .C(n4620), .Y(n5022));
MX2X1    g4636(.A(g2873), .B(n6708), .S0(n8686), .Y(n9285));
MX2X1    g4637(.A(g2868), .B(n9285), .S0(g35), .Y(n5027));
INVX1    g4638(.A(g1760), .Y(n9287));
NOR4X1   g4639(.A(n6467), .B(n4941), .C(n9287), .D(n6468_1), .Y(n9288));
MX2X1    g4640(.A(g1854), .B(g1848), .S0(n9288), .Y(n9289));
MX2X1    g4641(.A(g1848), .B(n9289), .S0(g35), .Y(n5032));
OR2X1    g4642(.A(g5084), .B(g5080), .Y(n9291));
AOI22X1  g4643(.A0(g5084), .A1(g5080), .B0(g5077), .B1(n7199), .Y(n9292));
OAI21X1  g4644(.A0(n9291), .A1(n8762), .B0(n9292), .Y(n9293));
MX2X1    g4645(.A(g5080), .B(n9293), .S0(g35), .Y(n5037));
NOR3X1   g4646(.A(n5899_1), .B(n5855_1), .C(n5854), .Y(n9295));
MX2X1    g4647(.A(g5603), .B(n5592_1), .S0(n9295), .Y(n9296));
MX2X1    g4648(.A(g5587), .B(n9296), .S0(g35), .Y(n5042));
NAND3X1  g4649(.A(n7102), .B(n7101), .C(g2465), .Y(n9298));
OAI21X1  g4650(.A0(n7101), .A1(n5151), .B0(n9298), .Y(n9299));
MX2X1    g4651(.A(g2465), .B(n9299), .S0(g35), .Y(n5051));
NOR3X1   g4652(.A(n7100), .B(g2495), .C(n7094), .Y(n9301));
MX2X1    g4653(.A(g2437), .B(n7132_1), .S0(n9301), .Y(n9302));
MX2X1    g4654(.A(g2429), .B(n9302), .S0(g35), .Y(n5056));
XOR2X1   g4655(.A(n7091), .B(g2102), .Y(n9304));
MX2X1    g4656(.A(g2098), .B(n9304), .S0(g35), .Y(n5061));
OAI21X1  g4657(.A0(n6204), .A1(n4914), .B0(n5789), .Y(n9306));
MX2X1    g4658(.A(g2208), .B(n9306), .S0(n5788), .Y(n9307));
MX2X1    g4659(.A(g2185), .B(n9307), .S0(g35), .Y(n5066));
AOI21X1  g4660(.A0(n6002), .A1(n5995), .B0(n7904), .Y(n9309));
MX2X1    g4661(.A(g2579), .B(n5998), .S0(n9309), .Y(n9310));
MX2X1    g4662(.A(g2583), .B(n9310), .S0(g35), .Y(n5071));
NAND2X1  g4663(.A(g4064), .B(g4169), .Y(n9312));
MX2X1    g4664(.A(g4072), .B(n9312), .S0(g35), .Y(n5076));
NAND3X1  g4665(.A(n6777_1), .B(g4975), .C(n4893), .Y(n9314));
OAI21X1  g4666(.A0(n6778), .A1(n4896_1), .B0(g4899), .Y(n9315));
AOI21X1  g4667(.A0(n9315), .A1(n9314), .B0(n6193), .Y(n9316));
MX2X1    g4668(.A(g4975), .B(n9316), .S0(g35), .Y(n5081));
NAND3X1  g4669(.A(n6468_1), .B(n5569), .C(g2841), .Y(n9318));
MX2X1    g4670(.A(g2715), .B(n9318), .S0(g35), .Y(n5086));
NAND3X1  g4671(.A(n6008), .B(n6007), .C(n4818), .Y(n9320));
NAND3X1  g4672(.A(n6009), .B(n6007), .C(g4785), .Y(n9321));
NAND2X1  g4673(.A(n9321), .B(n9320), .Y(n9322));
MX2X1    g4674(.A(g4776), .B(n9322), .S0(g35), .Y(n5091));
NOR3X1   g4675(.A(n5916), .B(g5517), .C(n5854), .Y(n9324));
MX2X1    g4676(.A(g5583), .B(n5592_1), .S0(n9324), .Y(n9325));
MX2X1    g4677(.A(g5563), .B(n9325), .S0(g35), .Y(n5096));
NAND4X1  g4678(.A(n5678), .B(n5677), .C(n6073_1), .D(n8984), .Y(n9327));
AOI21X1  g4679(.A0(g802), .A1(n5662), .B0(n5653), .Y(n9328));
MX2X1    g4680(.A(n5653), .B(n9328), .S0(n9327), .Y(n9329));
MX2X1    g4681(.A(g776), .B(n9329), .S0(g35), .Y(n5101));
MX2X1    g4682(.A(g6173), .B(g6167), .S0(n5910), .Y(n9331));
MX2X1    g4683(.A(g6167), .B(n9331), .S0(g35), .Y(n5106));
NOR3X1   g4684(.A(n5468), .B(n5286), .C(n5616), .Y(n9333));
AOI21X1  g4685(.A0(n4713), .A1(n4709), .B0(n4620), .Y(n9334));
OAI21X1  g4686(.A0(n9334), .A1(g2917), .B0(g35), .Y(n9335));
NAND2X1  g4687(.A(g2902), .B(n4620), .Y(n9336));
OAI21X1  g4688(.A0(n9335), .A1(n9333), .B0(n9336), .Y(n5115));
NAND3X1  g4689(.A(n6233), .B(n5516_1), .C(g703), .Y(n9338));
MX2X1    g4690(.A(g686), .B(n9338), .S0(n5880_1), .Y(n9339));
MX2X1    g4691(.A(g691), .B(n9339), .S0(g35), .Y(n5120));
AND2X1   g4692(.A(g1570), .B(g1252), .Y(n9341));
MX2X1    g4693(.A(n7708), .B(n9341), .S0(n7709), .Y(n9342));
MX2X1    g4694(.A(g1280), .B(n9342), .S0(g35), .Y(n5125));
INVX1    g4695(.A(g671), .Y(n9344));
OR2X1    g4696(.A(n6236_1), .B(n9344), .Y(n9345));
NAND2X1  g4697(.A(n6236_1), .B(n9344), .Y(n9346));
AOI21X1  g4698(.A0(n9346), .A1(n9345), .B0(n6238), .Y(n9347));
MX2X1    g4699(.A(g667), .B(n9347), .S0(g35), .Y(n5130));
MX2X1    g4700(.A(g2265), .B(g2259), .S0(n9122), .Y(n9349));
MX2X1    g4701(.A(g2259), .B(n9349), .S0(g35), .Y(n5135));
NOR4X1   g4702(.A(g6227), .B(n5980), .C(n4871_1), .D(g6203), .Y(n9351));
MX2X1    g4703(.A(g6283), .B(n5592_1), .S0(n9351), .Y(n9352));
MX2X1    g4704(.A(g6267), .B(n9352), .S0(g35), .Y(n5140));
INVX1    g4705(.A(g6455), .Y(n9354));
INVX1    g4706(.A(g6451), .Y(n9355));
AOI21X1  g4707(.A0(n9355), .A1(g35), .B0(n9354), .Y(n5153));
AND2X1   g4708(.A(g896), .B(n4620), .Y(n5158));
NAND2X1  g4709(.A(n4868), .B(g5523), .Y(n9358));
NAND2X1  g4710(.A(g5527), .B(n4866_1), .Y(n9359));
AOI21X1  g4711(.A0(n9359), .A1(n9358), .B0(n6932), .Y(n9360));
MX2X1    g4712(.A(g5523), .B(n9360), .S0(g35), .Y(n5166));
MX2X1    g4713(.A(g4486), .B(g6749), .S0(g35), .Y(n5171));
MX2X1    g4714(.A(g1974), .B(g1968), .S0(n9112), .Y(n9363));
MX2X1    g4715(.A(g1968), .B(n9363), .S0(g35), .Y(n5176));
INVX1    g4716(.A(g1270), .Y(n9365));
NAND2X1  g4717(.A(n7801), .B(g1263), .Y(n9366));
AND2X1   g4718(.A(g1570), .B(g1270), .Y(n9367));
MX2X1    g4719(.A(n9365), .B(n9367), .S0(n9366), .Y(n9368));
MX2X1    g4720(.A(g1263), .B(n9368), .S0(g35), .Y(n5181));
INVX1    g4721(.A(n4961), .Y(n9370));
NOR4X1   g4722(.A(g4966), .B(n6802), .C(n4962), .D(n9370), .Y(n9371));
AOI21X1  g4723(.A0(n9164), .A1(g4991), .B0(n4963), .Y(n9372));
OAI21X1  g4724(.A0(n9372), .A1(n9371), .B0(n6779), .Y(n9373));
NAND2X1  g4725(.A(g4991), .B(n4620), .Y(n9374));
OAI21X1  g4726(.A0(n9373), .A1(n4620), .B0(n9374), .Y(n5186));
NOR3X1   g4727(.A(n9174), .B(n6873), .C(n6885), .Y(n9376));
NOR3X1   g4728(.A(n6887), .B(g6411), .C(g6398), .Y(n9377));
OAI21X1  g4729(.A0(n9377), .A1(n9376), .B0(n9173), .Y(n9378));
NOR2X1   g4730(.A(n9377), .B(n9376), .Y(n9379));
NAND2X1  g4731(.A(n9379), .B(g6415), .Y(n9380));
OAI21X1  g4732(.A0(n9380), .A1(n6884), .B0(n9378), .Y(n9381));
MX2X1    g4733(.A(g6411), .B(n9381), .S0(g35), .Y(n5191));
OAI21X1  g4734(.A0(n4872), .A1(n4871_1), .B0(g6227), .Y(n9383));
NAND3X1  g4735(.A(n4873), .B(g6215), .C(g6219), .Y(n9384));
AOI21X1  g4736(.A0(n9384), .A1(n9383), .B0(n5646), .Y(n9385));
MX2X1    g4737(.A(g6219), .B(n9385), .S0(g35), .Y(n5196));
NOR4X1   g4738(.A(g3863), .B(n4850), .C(n4848), .D(n7642), .Y(n9387));
MX2X1    g4739(.A(g3929), .B(n5592_1), .S0(n9387), .Y(n9388));
MX2X1    g4740(.A(g3909), .B(n9388), .S0(g35), .Y(n5201));
INVX1    g4741(.A(g5503), .Y(n9390));
OAI22X1  g4742(.A0(n5524), .A1(g4284), .B0(n9390), .B1(n4869), .Y(n9391));
OR4X1    g4743(.A(n5524), .B(g4284), .C(n9390), .D(n4869), .Y(n9392));
AOI21X1  g4744(.A0(n9392), .A1(n9391), .B0(n4620), .Y(n5206));
NOR3X1   g4745(.A(g4229), .B(g4226), .C(g4185), .Y(n9394));
OR4X1    g4746(.A(g4213), .B(g4216), .C(g4235), .D(g4232), .Y(n9395));
NOR3X1   g4747(.A(n9395), .B(g4219), .C(g4222), .Y(n9396));
XOR2X1   g4748(.A(g4222), .B(g4235), .Y(n9397));
AOI21X1  g4749(.A0(n9396), .A1(n9394), .B0(n9397), .Y(n9398));
XOR2X1   g4750(.A(n9398), .B(n7558), .Y(n9399));
MX2X1    g4751(.A(g4235), .B(n9399), .S0(g35), .Y(n5211));
NOR4X1   g4752(.A(g5863), .B(n4862), .C(g5873), .D(n7375), .Y(n9401));
MX2X1    g4753(.A(g5925), .B(n5592_1), .S0(n9401), .Y(n9402));
MX2X1    g4754(.A(g5901), .B(n9402), .S0(g35), .Y(n5216));
INVX1    g4755(.A(g1124), .Y(n9404));
NOR3X1   g4756(.A(n4708), .B(n4707_1), .C(g976), .Y(n9405));
XOR2X1   g4757(.A(n9405), .B(n5305), .Y(n9406));
OR2X1    g4758(.A(g1146), .B(g1099), .Y(n9407));
AOI21X1  g4759(.A0(n9407), .A1(n9404), .B0(n9406), .Y(n9408));
NOR3X1   g4760(.A(n6188), .B(n6079), .C(n4665), .Y(n9409));
MX2X1    g4761(.A(g1124), .B(n9408), .S0(n9409), .Y(n9410));
MX2X1    g4762(.A(g1105), .B(n9410), .S0(g35), .Y(n5221));
AOI21X1  g4763(.A0(n4964_1), .A1(n6796), .B0(n6089), .Y(n9412));
MX2X1    g4764(.A(g4961), .B(g71), .S0(n6089), .Y(n9413));
MX2X1    g4765(.A(n9413), .B(g4955), .S0(n9412), .Y(n9414));
MX2X1    g4766(.A(g4961), .B(n9414), .S0(g35), .Y(n5226));
NOR3X1   g4767(.A(n6195), .B(g5170), .C(n5610), .Y(n9416));
MX2X1    g4768(.A(g5224), .B(n5592_1), .S0(n9416), .Y(n9417));
MX2X1    g4769(.A(g5196), .B(n9417), .S0(g35), .Y(n5231));
NOR3X1   g4770(.A(n6085), .B(g2070), .C(n8496), .Y(n9419));
MX2X1    g4771(.A(g2012), .B(n7037_1), .S0(n9419), .Y(n9420));
MX2X1    g4772(.A(g2004), .B(n9420), .S0(g35), .Y(n5236));
NOR4X1   g4773(.A(g6203), .B(g6215), .C(n4620), .D(n5646), .Y(n5241));
MX2X1    g4774(.A(g5120), .B(g5156), .S0(g26801), .Y(n9423));
MX2X1    g4775(.A(g5156), .B(n9423), .S0(g35), .Y(n5246));
XOR2X1   g4776(.A(g2384), .B(g2380), .Y(n9425));
NAND3X1  g4777(.A(n7227), .B(n7228), .C(g2342), .Y(n9426));
MX2X1    g4778(.A(n9425), .B(g2389), .S0(n9426), .Y(n9427));
MX2X1    g4779(.A(g2384), .B(n9427), .S0(g35), .Y(n5254));
AND2X1   g4780(.A(g4423), .B(g35), .Y(n5259));
NOR3X1   g4781(.A(n7100), .B(n7681), .C(g2465), .Y(n9430));
MX2X1    g4782(.A(g2429), .B(n7132_1), .S0(n9430), .Y(n9431));
MX2X1    g4783(.A(g2433), .B(n9431), .S0(g35), .Y(n5264));
OAI21X1  g4784(.A0(n4809), .A1(g113), .B0(g2795), .Y(n9433));
NAND4X1  g4785(.A(n5509), .B(g2729), .C(g2724), .D(n9433), .Y(n9434));
OAI22X1  g4786(.A0(n6900), .A1(n4806), .B0(n5507_1), .B1(n9434), .Y(n9435));
MX2X1    g4787(.A(g2795), .B(n9435), .S0(g35), .Y(n5269));
NAND2X1  g4788(.A(n3220), .B(g12), .Y(n9437));
NOR2X1   g4789(.A(n9437), .B(n6667), .Y(n9438));
OAI21X1  g4790(.A0(n4714), .A1(g1287), .B0(g35), .Y(n9439));
OAI22X1  g4791(.A0(n9438), .A1(n9439), .B0(n5454), .B1(g35), .Y(n5274));
XOR2X1   g4792(.A(n8533), .B(g2675), .Y(n9441));
MX2X1    g4793(.A(g2671), .B(n9441), .S0(g35), .Y(n5279));
NOR4X1   g4794(.A(g4322), .B(g4616), .C(g4608), .D(g4311), .Y(n9443));
NAND4X1  g4795(.A(n5178), .B(n5714), .C(n5204), .D(n9443), .Y(n9444));
NOR4X1   g4796(.A(g4601), .B(g4593), .C(n4620), .D(n5713_1), .Y(n9445));
NAND4X1  g4797(.A(g4633), .B(n5850_1), .C(g4621), .D(n9445), .Y(n9446));
OAI22X1  g4798(.A0(n9444), .A1(n9446), .B0(n5181_1), .B1(g35), .Y(n5284));
NAND4X1  g4799(.A(n5927), .B(n6491), .C(g35), .D(n6326_1), .Y(n9448));
NOR3X1   g4800(.A(n9448), .B(n6193), .C(n4961), .Y(n5289));
OR2X1    g4801(.A(n7146), .B(n7148), .Y(n9450));
OR4X1    g4802(.A(n6753), .B(g1199), .C(n6752_1), .D(n7145), .Y(n9451));
AOI21X1  g4803(.A0(n9451), .A1(n9450), .B0(n6761), .Y(n9452));
MX2X1    g4804(.A(g1193), .B(n9452), .S0(g35), .Y(n5294));
INVX1    g4805(.A(g1333), .Y(n9454));
XOR2X1   g4806(.A(n5988), .B(n9454), .Y(n9455));
MX2X1    g4807(.A(g1333), .B(n9455), .S0(g35), .Y(n5299));
NAND3X1  g4808(.A(n6462), .B(g5527), .C(n4867), .Y(n9457));
MX2X1    g4809(.A(n5592_1), .B(g5547), .S0(n9457), .Y(n9458));
MX2X1    g4810(.A(g5551), .B(n9458), .S0(g35), .Y(n5303));
XOR2X1   g4811(.A(g3782), .B(g3774), .Y(n9460));
MX2X1    g4812(.A(g3774), .B(n9460), .S0(g35), .Y(n5308));
NAND3X1  g4813(.A(n9175), .B(g6423), .C(g6419), .Y(n9462));
NAND3X1  g4814(.A(n9177), .B(n6878), .C(n9180), .Y(n9463));
AND2X1   g4815(.A(n9463), .B(n9462), .Y(n9464));
NOR2X1   g4816(.A(n6884), .B(n6875), .Y(n9465));
MX2X1    g4817(.A(n6875), .B(n9465), .S0(n9464), .Y(n9466));
MX2X1    g4818(.A(g6423), .B(n9466), .S0(g35), .Y(n5313));
MX2X1    g4819(.A(g2138), .B(n4586), .S0(n6029), .Y(n9468));
MX2X1    g4820(.A(g2130), .B(n9468), .S0(g35), .Y(n5318));
NOR4X1   g4821(.A(n6466), .B(n5134), .C(n5136), .D(n5551_1), .Y(n9470));
XOR2X1   g4822(.A(n5155), .B(g112), .Y(n9471));
MX2X1    g4823(.A(g2338), .B(n9471), .S0(n9470), .Y(n9472));
MX2X1    g4824(.A(g2287), .B(n9472), .S0(g35), .Y(n5326));
NAND3X1  g4825(.A(n7922), .B(g6227), .C(n4871_1), .Y(n9474));
MX2X1    g4826(.A(n5592_1), .B(g6247), .S0(n9474), .Y(n9475));
MX2X1    g4827(.A(g6251), .B(n9475), .S0(g35), .Y(n5335));
INVX1    g4828(.A(g2779), .Y(n9477));
INVX1    g4829(.A(g1902), .Y(n9478));
AOI21X1  g4830(.A0(n7859), .A1(n9478), .B0(g2791), .Y(n9479));
OAI22X1  g4831(.A0(n7861), .A1(n9479), .B0(n9477), .B1(g35), .Y(n5340));
NOR3X1   g4832(.A(n7042_1), .B(n7642), .C(n7041), .Y(n9481));
MX2X1    g4833(.A(g3949), .B(n5592_1), .S0(n9481), .Y(n9482));
MX2X1    g4834(.A(g3933), .B(n9482), .S0(g35), .Y(n5345));
OAI21X1  g4835(.A0(n6667), .A1(n5616), .B0(g1291), .Y(n9484));
OR4X1    g4836(.A(n5006), .B(n5019), .C(n5616), .D(n5462), .Y(n9485));
AOI21X1  g4837(.A0(n9485), .A1(n9484), .B0(n4620), .Y(n5350));
NOR4X1   g4838(.A(n6653_1), .B(n4862), .C(n4860), .D(g5857), .Y(n9487));
MX2X1    g4839(.A(g5945), .B(n5592_1), .S0(n9487), .Y(n9488));
MX2X1    g4840(.A(g5929), .B(n9488), .S0(g35), .Y(n5355));
NOR4X1   g4841(.A(g5188), .B(g5164), .C(n4642_1), .D(n6624), .Y(n9490));
MX2X1    g4842(.A(g5244), .B(n5592_1), .S0(n9490), .Y(n9491));
MX2X1    g4843(.A(g5228), .B(n9491), .S0(g35), .Y(n5360));
NAND2X1  g4844(.A(n7693), .B(g2756), .Y(n9493));
XOR2X1   g4845(.A(n9493), .B(g2759), .Y(n9494));
NAND2X1  g4846(.A(n9494), .B(g2841), .Y(n9495));
MX2X1    g4847(.A(g2756), .B(n9495), .S0(g35), .Y(n5365));
NAND3X1  g4848(.A(n9275), .B(n7721), .C(n8575), .Y(n9497));
OAI21X1  g4849(.A0(n7721), .A1(n8575), .B0(n9497), .Y(n9498));
MX2X1    g4850(.A(g6736), .B(n9498), .S0(g35), .Y(n5370));
AOI21X1  g4851(.A0(g802), .A1(n5662), .B0(n5438), .Y(n9500));
MX2X1    g4852(.A(n5438), .B(n9500), .S0(n5680), .Y(n9501));
MX2X1    g4853(.A(g781), .B(n9501), .S0(g35), .Y(n5375));
INVX1    g4854(.A(g1280), .Y(n9503));
NAND3X1  g4855(.A(g1570), .B(g1266), .C(g1249), .Y(n9504));
OR4X1    g4856(.A(n9503), .B(n7708), .C(n7707), .D(n9504), .Y(n9505));
AND2X1   g4857(.A(g1570), .B(g1259), .Y(n9506));
MX2X1    g4858(.A(n7800), .B(n9506), .S0(n9505), .Y(n9507));
MX2X1    g4859(.A(g1256), .B(n9507), .S0(g35), .Y(n5380));
XOR2X1   g4860(.A(n7393), .B(g3484), .Y(n9509));
MX2X1    g4861(.A(g3480), .B(n9509), .S0(g35), .Y(n5385));
XOR2X1   g4862(.A(g191), .B(g194), .Y(n9511));
MX2X1    g4863(.A(g209), .B(n9511), .S0(n9088), .Y(n9512));
MX2X1    g4864(.A(g191), .B(n9512), .S0(g35), .Y(n5390));
NOR3X1   g4865(.A(n7657), .B(g6555), .C(n7524), .Y(n9514));
MX2X1    g4866(.A(g6609), .B(n5592_1), .S0(n9514), .Y(n9515));
MX2X1    g4867(.A(g6581), .B(n9515), .S0(g35), .Y(n5395));
NAND2X1  g4868(.A(g5517), .B(n5854), .Y(n9517));
NAND2X1  g4869(.A(n5855_1), .B(g5511), .Y(n9518));
AOI21X1  g4870(.A0(n9518), .A1(n9517), .B0(n6932), .Y(n9519));
MX2X1    g4871(.A(g5511), .B(n9519), .S0(g35), .Y(n5400));
NOR3X1   g4872(.A(n7100), .B(n5151), .C(g2465), .Y(n9521));
MX2X1    g4873(.A(g2449), .B(n7132_1), .S0(n9521), .Y(n9522));
MX2X1    g4874(.A(g2437), .B(n9522), .S0(g35), .Y(n5405));
NOR3X1   g4875(.A(n6003), .B(n5999), .C(n5156), .Y(n9524));
MX2X1    g4876(.A(g2575), .B(n5998), .S0(n9524), .Y(n9525));
MX2X1    g4877(.A(g2579), .B(n9525), .S0(g35), .Y(n5410));
OR2X1    g4878(.A(n4809), .B(n4879), .Y(n9527));
OAI21X1  g4879(.A0(n4809), .A1(n4879), .B0(g66), .Y(n9528));
OAI21X1  g4880(.A0(n4880), .A1(n9527), .B0(n9528), .Y(n5415));
NAND2X1  g4881(.A(g2715), .B(g2841), .Y(n9530));
MX2X1    g4882(.A(g2712), .B(n9530), .S0(g35), .Y(n5420));
AND2X1   g4883(.A(g936), .B(g1227), .Y(n9532));
MX2X1    g4884(.A(n7164), .B(n9532), .S0(n7165), .Y(n9533));
MX2X1    g4885(.A(g921), .B(n9533), .S0(g35), .Y(n5425));
XOR2X1   g4886(.A(g2093), .B(g2089), .Y(n9535));
NOR3X1   g4887(.A(n7090), .B(n9215), .C(g2028), .Y(n9536));
MX2X1    g4888(.A(g2098), .B(n9535), .S0(n9536), .Y(n9537));
MX2X1    g4889(.A(g2093), .B(n9537), .S0(g35), .Y(n5430));
NAND3X1  g4890(.A(g4473), .B(g4462), .C(n5844), .Y(n9539));
OAI21X1  g4891(.A0(n8769), .A1(g4467), .B0(g4473), .Y(n9540));
NAND3X1  g4892(.A(n9540), .B(n9539), .C(n7745), .Y(n9541));
MX2X1    g4893(.A(g4473), .B(n9541), .S0(g35), .Y(n5435));
AOI21X1  g4894(.A0(g640), .A1(n6133), .B0(n5436), .Y(n9543));
MX2X1    g4895(.A(n5436), .B(n9543), .S0(n9044), .Y(n9544));
MX2X1    g4896(.A(g599), .B(n9544), .S0(g35), .Y(n5440));
NOR2X1   g4897(.A(n7657), .B(n4856_1), .Y(n9546));
MX2X1    g4898(.A(g6589), .B(n5592_1), .S0(n9546), .Y(n9547));
MX2X1    g4899(.A(g6641), .B(n9547), .S0(g35), .Y(n5445));
NAND2X1  g4900(.A(g1906), .B(n5527), .Y(n9549));
AOI21X1  g4901(.A0(n5530), .A1(n5521_1), .B0(n9549), .Y(n9550));
MX2X1    g4902(.A(g1886), .B(n5526_1), .S0(n9550), .Y(n9551));
MX2X1    g4903(.A(g1890), .B(n9551), .S0(g35), .Y(n5450));
OR2X1    g4904(.A(g6466), .B(g6462), .Y(n9553));
AOI22X1  g4905(.A0(g6466), .A1(g6462), .B0(g6459), .B1(n9354), .Y(n9554));
OAI21X1  g4906(.A0(n9553), .A1(n5537), .B0(n9554), .Y(n9555));
MX2X1    g4907(.A(g6462), .B(n9555), .S0(g35), .Y(n5455));
MX2X1    g4908(.A(g429), .B(g433), .S0(n5688), .Y(n9557));
MX2X1    g4909(.A(g433), .B(n9557), .S0(g35), .Y(n5467));
NOR3X1   g4910(.A(n5531_1), .B(g1906), .C(n5527), .Y(n9559));
MX2X1    g4911(.A(g1870), .B(n5526_1), .S0(n9559), .Y(n9560));
MX2X1    g4912(.A(g1874), .B(n9560), .S0(g35), .Y(n5472));
NOR3X1   g4913(.A(n5004), .B(n4988_1), .C(n5616), .Y(n9562));
MX2X1    g4914(.A(g4249), .B(n4586), .S0(n9562), .Y(n9563));
MX2X1    g4915(.A(g4253), .B(n9563), .S0(g35), .Y(n5477));
MX2X1    g4916(.A(g6451), .B(n6880), .S0(g35), .Y(n5482));
OAI21X1  g4917(.A0(g3050), .A1(g3010), .B0(n6588), .Y(n9566));
NAND3X1  g4918(.A(g3004), .B(n5573_1), .C(n6593), .Y(n9567));
OAI21X1  g4919(.A0(n9566), .A1(n5584), .B0(n9567), .Y(n9568));
MX2X1    g4920(.A(g3010), .B(n9568), .S0(g35), .Y(n5487));
INVX1    g4921(.A(g1825), .Y(n9570));
AOI21X1  g4922(.A0(g1783), .A1(n9287), .B0(n9570), .Y(n9571));
XOR2X1   g4923(.A(n9571), .B(g1811), .Y(n9572));
MX2X1    g4924(.A(g1825), .B(n9572), .S0(n8134), .Y(n9573));
MX2X1    g4925(.A(g1811), .B(n9573), .S0(g35), .Y(n5492));
XOR2X1   g4926(.A(n6402), .B(g6133), .Y(n9575));
MX2X1    g4927(.A(g6128), .B(n9575), .S0(g35), .Y(n5497));
NAND2X1  g4928(.A(g1018), .B(g1030), .Y(n9577));
NAND4X1  g4929(.A(n6050), .B(n6052), .C(g1008), .D(n9577), .Y(n9578));
NAND2X1  g4930(.A(n9577), .B(g1008), .Y(n9579));
MX2X1    g4931(.A(n9579), .B(n7173), .S0(n6050), .Y(n9580));
NAND2X1  g4932(.A(n9580), .B(n9578), .Y(n9581));
MX2X1    g4933(.A(g1008), .B(n9581), .S0(n6059), .Y(n9582));
MX2X1    g4934(.A(g969), .B(n9582), .S0(g35), .Y(n5502));
MX2X1    g4935(.A(g4392), .B(n6992), .S0(n6906_1), .Y(n9584));
MX2X1    g4936(.A(g4417), .B(n9584), .S0(g35), .Y(n5507));
NOR2X1   g4937(.A(n6067), .B(n4834), .Y(n9586));
MX2X1    g4938(.A(g3546), .B(n5592_1), .S0(n9586), .Y(n9587));
MX2X1    g4939(.A(g3598), .B(n9587), .S0(g35), .Y(n5516));
NOR3X1   g4940(.A(n7933), .B(g5170), .C(n5610), .Y(n9589));
MX2X1    g4941(.A(g5236), .B(n5592_1), .S0(n9589), .Y(n9590));
MX2X1    g4942(.A(g5216), .B(n9590), .S0(g35), .Y(n5521));
NOR4X1   g4943(.A(n6467), .B(g1792), .C(n8135), .D(n6468_1), .Y(n9592));
MX2X1    g4944(.A(g1768), .B(n6577), .S0(n9592), .Y(n9593));
MX2X1    g4945(.A(g1748), .B(n9593), .S0(g35), .Y(n5526));
AND2X1   g4946(.A(n6192), .B(n9370), .Y(n9595));
INVX1    g4947(.A(g4854), .Y(n9596));
AND2X1   g4948(.A(g4843), .B(g4878), .Y(n9597));
AOI21X1  g4949(.A0(n9597), .A1(g4849), .B0(n9596), .Y(n9598));
INVX1    g4950(.A(g4849), .Y(n9599));
INVX1    g4951(.A(g4843), .Y(n9600));
NOR4X1   g4952(.A(n9599), .B(g4854), .C(n4959_1), .D(n9600), .Y(n9601));
OAI21X1  g4953(.A0(n9601), .A1(n9598), .B0(n9595), .Y(n9602));
NAND2X1  g4954(.A(g4849), .B(n4620), .Y(n9603));
OAI21X1  g4955(.A0(n9602), .A1(n4620), .B0(n9603), .Y(n5531));
NOR4X1   g4956(.A(g3863), .B(n4850), .C(g3873), .D(n7642), .Y(n9605));
MX2X1    g4957(.A(g3925), .B(n5592_1), .S0(n9605), .Y(n9606));
MX2X1    g4958(.A(g3901), .B(n9606), .S0(g35), .Y(n5536));
XOR2X1   g4959(.A(g6505), .B(g6500), .Y(n9608));
MX2X1    g4960(.A(g6509), .B(n9608), .S0(n7724), .Y(n9609));
MX2X1    g4961(.A(g6500), .B(n9609), .S0(g35), .Y(n5541));
XOR2X1   g4962(.A(g255), .B(g232), .Y(n9611));
XOR2X1   g4963(.A(n9611), .B(n6105_1), .Y(n9612));
XOR2X1   g4964(.A(g262), .B(g239), .Y(n9613));
XOR2X1   g4965(.A(g269), .B(g246), .Y(n9614));
XOR2X1   g4966(.A(n9614), .B(n9613), .Y(n9615));
XOR2X1   g4967(.A(n9615), .B(n9612), .Y(n9616));
OAI21X1  g4968(.A0(n5657), .A1(n5655_1), .B0(g732), .Y(n9617));
XOR2X1   g4969(.A(n9617), .B(n9616), .Y(n9618));
AND2X1   g4970(.A(g496), .B(g35), .Y(n9619));
MX2X1    g4971(.A(n9618), .B(n9619), .S0(n4620), .Y(n5546));
NAND3X1  g4972(.A(n5562), .B(g2441), .C(n4929), .Y(n9621));
NAND3X1  g4973(.A(n5562), .B(g2429), .C(g2476), .Y(n9622));
AND2X1   g4974(.A(n9622), .B(n9621), .Y(n9623));
AND2X1   g4975(.A(g2453), .B(g2485), .Y(n9624));
NOR2X1   g4976(.A(g2476), .B(n4929), .Y(n9625));
AOI22X1  g4977(.A0(n9624), .A1(g2433), .B0(g2437), .B1(n9625), .Y(n9626));
NAND3X1  g4978(.A(g2449), .B(g2476), .C(n4929), .Y(n9627));
NAND3X1  g4979(.A(g2453), .B(g2445), .C(n6445), .Y(n9628));
NAND4X1  g4980(.A(n9627), .B(n9626), .C(n9623), .D(n9628), .Y(n9629));
MX2X1    g4981(.A(g2504), .B(n9629), .S0(n6444_1), .Y(n9630));
MX2X1    g4982(.A(g2485), .B(n9630), .S0(g35), .Y(n5551));
OAI21X1  g4983(.A0(g2185), .A1(n5797_1), .B0(n4937), .Y(n9632));
OAI21X1  g4984(.A0(n6204), .A1(n4914), .B0(n9632), .Y(n9633));
MX2X1    g4985(.A(g2185), .B(n9633), .S0(n5788), .Y(n9634));
MX2X1    g4986(.A(g2193), .B(n9634), .S0(g35), .Y(n5568));
NOR3X1   g4987(.A(n5011), .B(n5006), .C(n5616), .Y(n9636));
MX2X1    g4988(.A(g37), .B(n2447), .S0(n9636), .Y(n9637));
MX2X1    g4989(.A(g2894), .B(n9637), .S0(g35), .Y(n5573));
NAND3X1  g4990(.A(n8498), .B(n8497), .C(g2040), .Y(n9639));
OAI21X1  g4991(.A0(n8497), .A1(n5166_1), .B0(n9639), .Y(n9640));
MX2X1    g4992(.A(g2040), .B(n9640), .S0(g35), .Y(n5583));
MX2X1    g4993(.A(n6181), .B(n6183_1), .S0(n5811_1), .Y(n9642));
NOR2X1   g4994(.A(n5820), .B(n9281), .Y(n9643));
MX2X1    g4995(.A(n9643), .B(n9281), .S0(n9642), .Y(n9644));
MX2X1    g4996(.A(g6088), .B(n9644), .S0(g35), .Y(n5592));
AND2X1   g4997(.A(g967), .B(n4620), .Y(n5597));
AND2X1   g4998(.A(n5697), .B(n6708), .Y(n9647));
OAI21X1  g4999(.A0(g4176), .A1(g4072), .B0(g35), .Y(n9648));
OAI22X1  g5000(.A0(n9647), .A1(n9648), .B0(n5393), .B1(g35), .Y(n5602));
OAI22X1  g5001(.A0(n5557), .A1(g4005), .B0(g4012), .B1(n5556), .Y(n9650));
MX2X1    g5002(.A(g4000), .B(n5556), .S0(g3976), .Y(n9651));
INVX1    g5003(.A(g4012), .Y(n9652));
OAI21X1  g5004(.A0(g3983), .A1(n9652), .B0(g35), .Y(n9653));
NOR4X1   g5005(.A(n9651), .B(n9650), .C(n5559), .D(n9653), .Y(n5607));
XOR2X1   g5006(.A(n5910), .B(g6181), .Y(n9655));
MX2X1    g5007(.A(g6177), .B(n9655), .S0(g35), .Y(n5620));
XOR2X1   g5008(.A(n6998_1), .B(g6381), .Y(n9657));
MX2X1    g5009(.A(g6377), .B(n9657), .S0(g35), .Y(n5625));
AOI21X1  g5010(.A0(n4970), .A1(n7428), .B0(n6721), .Y(n9659));
MX2X1    g5011(.A(g4771), .B(g101), .S0(n6721), .Y(n9660));
MX2X1    g5012(.A(n9660), .B(g4765), .S0(n9659), .Y(n9661));
MX2X1    g5013(.A(g4771), .B(n9661), .S0(g35), .Y(n5630));
NOR4X1   g5014(.A(g5517), .B(g5523), .C(g5511), .D(n5916), .Y(n9663));
MX2X1    g5015(.A(g5563), .B(n5592_1), .S0(n9663), .Y(n9664));
MX2X1    g5016(.A(g5567), .B(n9664), .S0(g35), .Y(n5635));
OAI21X1  g5017(.A0(n8826), .A1(n8825), .B0(n8824), .Y(n9666));
NOR3X1   g5018(.A(n8827), .B(g1322), .C(n4620), .Y(n9667));
AND2X1   g5019(.A(n9667), .B(n9666), .Y(n5640));
NOR4X1   g5020(.A(n6466), .B(n5145_1), .C(n5136), .D(n5530), .Y(n9669));
XOR2X1   g5021(.A(n5162_1), .B(g112), .Y(n9670));
MX2X1    g5022(.A(g1913), .B(n9670), .S0(n9669), .Y(n9671));
MX2X1    g5023(.A(g1862), .B(n9671), .S0(g35), .Y(n5645));
INVX1    g5024(.A(g2331), .Y(n9673));
NAND3X1  g5025(.A(n6730), .B(n6729), .C(g2287), .Y(n9674));
OAI21X1  g5026(.A0(n6729), .A1(n9673), .B0(n9674), .Y(n9675));
MX2X1    g5027(.A(g2338), .B(n9675), .S0(g35), .Y(n5650));
NOR3X1   g5028(.A(n7379), .B(n6208), .C(g6209), .Y(n9677));
MX2X1    g5029(.A(g6263), .B(n5592_1), .S0(n9677), .Y(n9678));
MX2X1    g5030(.A(g6235), .B(n9678), .S0(g35), .Y(n5655));
OAI21X1  g5031(.A0(n5425_1), .A1(n5405_1), .B0(n5282), .Y(n9680));
OAI21X1  g5032(.A0(n5425_1), .A1(n5405_1), .B0(g22), .Y(n9681));
NAND2X1  g5033(.A(n9681), .B(n9680), .Y(n5660));
NOR4X1   g5034(.A(n7041), .B(n4850), .C(n4848), .D(g3857), .Y(n9683));
MX2X1    g5035(.A(g3945), .B(n5592_1), .S0(n9683), .Y(n9684));
MX2X1    g5036(.A(g3929), .B(n9684), .S0(g35), .Y(n5665));
INVX1    g5037(.A(n7061), .Y(n9686));
INVX1    g5038(.A(n7066), .Y(n9687));
MX2X1    g5039(.A(n9686), .B(n9687), .S0(n7064), .Y(n9688));
OR2X1    g5040(.A(n9688), .B(g5731), .Y(n9689));
NAND2X1  g5041(.A(n9688), .B(g5731), .Y(n9690));
OAI21X1  g5042(.A0(n9690), .A1(n7077), .B0(n9689), .Y(n9691));
MX2X1    g5043(.A(g5727), .B(n9691), .S0(g35), .Y(n5674));
AOI21X1  g5044(.A0(g4473), .A1(n8769), .B0(g4459), .Y(n9693));
NAND2X1  g5045(.A(n9693), .B(n7745), .Y(n9694));
MX2X1    g5046(.A(g4369), .B(n9694), .S0(g35), .Y(n5679));
INVX1    g5047(.A(g1266), .Y(n9696));
AND2X1   g5048(.A(g1570), .B(g1249), .Y(n9697));
AND2X1   g5049(.A(g1570), .B(g1266), .Y(n9698));
MX2X1    g5050(.A(n9698), .B(n9696), .S0(n9697), .Y(n9699));
MX2X1    g5051(.A(g1249), .B(n9699), .S0(g35), .Y(n5684));
NAND4X1  g5052(.A(g5703), .B(g5689), .C(g5630), .D(g5644), .Y(n9701));
NOR2X1   g5053(.A(n9701), .B(n7031), .Y(n9702));
XOR2X1   g5054(.A(n9702), .B(g5489), .Y(n9703));
MX2X1    g5055(.A(g5485), .B(n9703), .S0(g35), .Y(n5689));
OAI21X1  g5056(.A0(n6239), .A1(n6241_1), .B0(g714), .Y(n9705));
INVX1    g5057(.A(g714), .Y(n9706));
NAND4X1  g5058(.A(n9706), .B(g671), .C(g676), .D(n6236_1), .Y(n9707));
AOI21X1  g5059(.A0(n9707), .A1(n9705), .B0(n6238), .Y(n9708));
MX2X1    g5060(.A(g676), .B(n9708), .S0(g35), .Y(n5694));
NOR3X1   g5061(.A(n7692), .B(n5508), .C(n4909), .Y(n9710));
XOR2X1   g5062(.A(n9710), .B(n4915_1), .Y(n9711));
OAI22X1  g5063(.A0(n8854), .A1(n9711), .B0(n4909), .B1(g35), .Y(n5699));
XOR2X1   g5064(.A(g5462), .B(g5467), .Y(n9713));
MX2X1    g5065(.A(g5471), .B(n9713), .S0(n9702), .Y(n9714));
MX2X1    g5066(.A(g5462), .B(n9714), .S0(g35), .Y(n5704));
NAND3X1  g5067(.A(n5920), .B(g73), .C(g72), .Y(n9716));
MX2X1    g5068(.A(g4372), .B(n9716), .S0(g4581), .Y(n9717));
MX2X1    g5069(.A(g4423), .B(n9717), .S0(g35), .Y(n5709));
NOR3X1   g5070(.A(n4856_1), .B(g6565), .C(n4854), .Y(n9719));
MX2X1    g5071(.A(g6605), .B(n5592_1), .S0(n9719), .Y(n9720));
MX2X1    g5072(.A(g6649), .B(n9720), .S0(g35), .Y(n5718));
AOI21X1  g5073(.A0(n7099), .A1(n7096), .B0(n7682), .Y(n9722));
MX2X1    g5074(.A(g2445), .B(n7132_1), .S0(n9722), .Y(n9723));
MX2X1    g5075(.A(g2449), .B(n9723), .S0(g35), .Y(n5723));
NOR3X1   g5076(.A(n7511_1), .B(n5159), .C(n6708_1), .Y(n9725));
MX2X1    g5077(.A(g2173), .B(n6705), .S0(n9725), .Y(n9726));
MX2X1    g5078(.A(g2177), .B(n9726), .S0(g35), .Y(n5728));
INVX1    g5079(.A(g4287), .Y(n9728));
XOR2X1   g5080(.A(n9204), .B(n9728), .Y(n9729));
MX2X1    g5081(.A(g4284), .B(n9729), .S0(g35), .Y(n5733));
NOR4X1   g5082(.A(n5567), .B(n6466), .C(n4917), .D(n5569), .Y(n9731));
XOR2X1   g5083(.A(n9625), .B(g110), .Y(n9732));
MX2X1    g5084(.A(g2491), .B(n9732), .S0(n9731), .Y(n9733));
MX2X1    g5085(.A(g2476), .B(n9733), .S0(g35), .Y(n5738));
AND2X1   g5086(.A(n9597), .B(n9599), .Y(n9735));
NOR2X1   g5087(.A(n9597), .B(n9599), .Y(n9736));
OAI21X1  g5088(.A0(n9736), .A1(n9735), .B0(n9595), .Y(n9737));
NAND2X1  g5089(.A(g4843), .B(n4620), .Y(n9738));
OAI21X1  g5090(.A0(n9737), .A1(n4620), .B0(n9738), .Y(n5743));
INVX1    g5091(.A(g2197), .Y(n9740));
NOR3X1   g5092(.A(n7511_1), .B(n9740), .C(g2227), .Y(n9741));
MX2X1    g5093(.A(g2169), .B(n6705), .S0(n9741), .Y(n9742));
MX2X1    g5094(.A(g2161), .B(n9742), .S0(g35), .Y(n5748));
INVX1    g5095(.A(g2279), .Y(n9744));
XOR2X1   g5096(.A(g2273), .B(n9744), .Y(n9745));
MX2X1    g5097(.A(g2283), .B(n9745), .S0(n6894), .Y(n9746));
MX2X1    g5098(.A(g2279), .B(n9746), .S0(g35), .Y(n5753));
NAND3X1  g5099(.A(n8319), .B(g6565), .C(n4854), .Y(n9748));
MX2X1    g5100(.A(n5592_1), .B(g6585), .S0(n9748), .Y(n9749));
MX2X1    g5101(.A(g6589), .B(n9749), .S0(g35), .Y(n5758));
MX2X1    g5102(.A(g2831), .B(n9238), .S0(g35), .Y(n5763));
XOR2X1   g5103(.A(n5553), .B(g2407), .Y(n9752));
MX2X1    g5104(.A(g2403), .B(n9752), .S0(g35), .Y(n5768));
MX2X1    g5105(.A(g2868), .B(n2447), .S0(n8686), .Y(n9754));
MX2X1    g5106(.A(g2988), .B(n9754), .S0(g35), .Y(n5773));
INVX1    g5107(.A(g1632), .Y(n9756));
AOI21X1  g5108(.A0(n7859), .A1(n9756), .B0(g2767), .Y(n9757));
NAND2X1  g5109(.A(g2763), .B(n4620), .Y(n9758));
OAI21X1  g5110(.A0(n9757), .A1(n7861), .B0(n9758), .Y(n5778));
OAI21X1  g5111(.A0(n6204), .A1(n4925_1), .B0(n9287), .Y(n9760));
MX2X1    g5112(.A(g1783), .B(n9760), .S0(n8134), .Y(n9761));
MX2X1    g5113(.A(g1760), .B(n9761), .S0(g35), .Y(n5783));
OR2X1    g5114(.A(n8327), .B(g1351), .Y(n9763));
OAI22X1  g5115(.A0(n7284), .A1(g1389), .B0(n5984), .B1(n9763), .Y(n9764));
INVX1    g5116(.A(g1312), .Y(n9765));
AOI21X1  g5117(.A0(n7284), .A1(n9765), .B0(n5984), .Y(n9766));
OAI21X1  g5118(.A0(n9766), .A1(n9764), .B0(n5986), .Y(n9767));
NAND2X1  g5119(.A(n5985), .B(g1312), .Y(n9768));
AOI21X1  g5120(.A0(n9768), .A1(n9767), .B0(n4620), .Y(n5792));
NOR3X1   g5121(.A(n4644), .B(g5188), .C(n4642_1), .Y(n9770));
MX2X1    g5122(.A(g5212), .B(n5592_1), .S0(n9770), .Y(n9771));
MX2X1    g5123(.A(g5260), .B(n9771), .S0(g35), .Y(n5797));
MX2X1    g5124(.A(g4245), .B(n3220), .S0(n9562), .Y(n9773));
MX2X1    g5125(.A(g4249), .B(n9773), .S0(g35), .Y(n5802));
MX2X1    g5126(.A(g446), .B(g645), .S0(n6389_1), .Y(n9775));
AND2X1   g5127(.A(n9775), .B(g35), .Y(n5807));
OR2X1    g5128(.A(g728), .B(g661), .Y(n9777));
MX2X1    g5129(.A(g79), .B(n9777), .S0(n6236_1), .Y(n9778));
MX2X1    g5130(.A(g728), .B(n9778), .S0(g35), .Y(n5816));
MX2X1    g5131(.A(g182), .B(g446), .S0(n5601), .Y(n9780));
MX2X1    g5132(.A(g405), .B(n9780), .S0(g35), .Y(n5821));
NOR4X1   g5133(.A(n6188), .B(n6079), .C(n4665), .D(n6397), .Y(n9782));
XOR2X1   g5134(.A(g1129), .B(g1124), .Y(n9783));
MX2X1    g5135(.A(g1129), .B(n9783), .S0(n9782), .Y(n9784));
MX2X1    g5136(.A(g1124), .B(n9784), .S0(g35), .Y(n5826));
NAND3X1  g5137(.A(n8913), .B(n7512), .C(g2197), .Y(n9786));
OAI21X1  g5138(.A0(n7512), .A1(n5159), .B0(n9786), .Y(n9787));
MX2X1    g5139(.A(g2197), .B(n9787), .S0(g35), .Y(n5831));
INVX1    g5140(.A(g6151), .Y(n9789));
AOI21X1  g5141(.A0(n9789), .A1(g6144), .B0(g6058), .Y(n9790));
OR2X1    g5142(.A(g6140), .B(n4620), .Y(n9791));
OAI22X1  g5143(.A0(n9790), .A1(n9791), .B0(n9789), .B1(g35), .Y(n5836));
MX2X1    g5144(.A(g2246), .B(g2241), .S0(n9122), .Y(n9793));
MX2X1    g5145(.A(g2241), .B(n9793), .S0(g35), .Y(n5845));
XOR2X1   g5146(.A(g1821), .B(g1825), .Y(n9795));
NOR4X1   g5147(.A(n6467), .B(n8135), .C(g1760), .D(n6468_1), .Y(n9796));
MX2X1    g5148(.A(g1830), .B(n9795), .S0(n9796), .Y(n9797));
MX2X1    g5149(.A(g1825), .B(n9797), .S0(g35), .Y(n5850));
NOR4X1   g5150(.A(n4833), .B(g3506), .C(n5733_1), .D(g3522), .Y(n9799));
MX2X1    g5151(.A(g3590), .B(n5592_1), .S0(n9799), .Y(n9800));
MX2X1    g5152(.A(g3574), .B(n9800), .S0(g35), .Y(n5855));
NOR2X1   g5153(.A(n8731), .B(g703), .Y(n9802));
MX2X1    g5154(.A(g392), .B(n9802), .S0(n5688), .Y(n9803));
MX2X1    g5155(.A(g401), .B(n9803), .S0(g35), .Y(n5860));
NAND2X1  g5156(.A(n5758_1), .B(g1592), .Y(n9805));
AOI21X1  g5157(.A0(g1636), .A1(n5757), .B0(g1668), .Y(n9806));
NAND3X1  g5158(.A(n9806), .B(n8425), .C(n7211), .Y(n9807));
AOI21X1  g5159(.A0(n9807), .A1(n9805), .B0(n4620), .Y(n5865));
MX2X1    g5160(.A(g6505), .B(g6541), .S0(n4857), .Y(n9809));
MX2X1    g5161(.A(g6541), .B(n9809), .S0(g35), .Y(n5870));
MX2X1    g5162(.A(g6404), .B(g6444), .S0(g6398), .Y(n9811));
OR2X1    g5163(.A(n9811), .B(n9174), .Y(n9812));
NAND2X1  g5164(.A(n9811), .B(n9174), .Y(n9813));
OAI21X1  g5165(.A0(n9812), .A1(n6884), .B0(n9813), .Y(n9814));
MX2X1    g5166(.A(g6398), .B(n9814), .S0(g35), .Y(n5875));
AND2X1   g5167(.A(g1087), .B(g1205), .Y(n9816));
XOR2X1   g5168(.A(n9816), .B(g1221), .Y(n9817));
MX2X1    g5169(.A(g1205), .B(n9817), .S0(g35), .Y(n5880));
NOR4X1   g5170(.A(g5863), .B(g5881), .C(n4860), .D(n7375), .Y(n9819));
MX2X1    g5171(.A(g5921), .B(n5592_1), .S0(n9819), .Y(n9820));
MX2X1    g5172(.A(g5893), .B(n9820), .S0(g35), .Y(n5885));
INVX1    g5173(.A(g329), .Y(n9822));
OR4X1    g5174(.A(n9822), .B(g341), .C(n4620), .D(n8036), .Y(n9823));
NAND2X1  g5175(.A(g74), .B(n4620), .Y(n9824));
NAND2X1  g5176(.A(n9824), .B(n9823), .Y(n5890));
OR4X1    g5177(.A(n7300), .B(n5661), .C(g146), .D(n7302_1), .Y(n9826));
NAND3X1  g5178(.A(n7303), .B(n7300), .C(g146), .Y(n9827));
NAND2X1  g5179(.A(n9827), .B(n9826), .Y(n9828));
MX2X1    g5180(.A(g142), .B(n9828), .S0(g35), .Y(n5895));
XOR2X1   g5181(.A(g6474), .B(g6466), .Y(n9830));
MX2X1    g5182(.A(g6466), .B(n9830), .S0(g35), .Y(n5904));
NOR4X1   g5183(.A(n5569), .B(n6466), .C(n4924), .D(n5840), .Y(n9832));
XOR2X1   g5184(.A(n8927), .B(g110), .Y(n9833));
MX2X1    g5185(.A(g1932), .B(n9833), .S0(n9832), .Y(n9834));
MX2X1    g5186(.A(g1917), .B(n9834), .S0(g35), .Y(n5909));
OAI21X1  g5187(.A0(n4629), .A1(g1624), .B0(n7397_1), .Y(n9836));
OAI21X1  g5188(.A0(n6204), .A1(n4922), .B0(n9836), .Y(n9837));
MX2X1    g5189(.A(g1624), .B(n9837), .S0(n8992), .Y(n9838));
MX2X1    g5190(.A(g1632), .B(n9838), .S0(g35), .Y(n5914));
INVX1    g5191(.A(g5109), .Y(n9840));
AOI21X1  g5192(.A0(g5101), .A1(n9840), .B0(g5062), .Y(n9841));
OR2X1    g5193(.A(g5105), .B(n4620), .Y(n9842));
OAI22X1  g5194(.A0(n9841), .A1(n9842), .B0(n9840), .B1(g35), .Y(n5919));
INVX1    g5195(.A(g5689), .Y(n9844));
NAND3X1  g5196(.A(n9844), .B(g5630), .C(g5559), .Y(n9845));
NAND3X1  g5197(.A(g5547), .B(g5689), .C(g5659), .Y(n9846));
AOI21X1  g5198(.A0(n9846), .A1(n9845), .B0(n7027_1), .Y(n9847));
NAND4X1  g5199(.A(g5673), .B(n9844), .C(g5579), .D(n5194), .Y(n9848));
NAND3X1  g5200(.A(g5654), .B(n9844), .C(g5555), .Y(n9849));
OAI21X1  g5201(.A0(n9849), .A1(n7020), .B0(n9848), .Y(n9850));
NOR2X1   g5202(.A(n9850), .B(n9847), .Y(n9851));
AND2X1   g5203(.A(g5673), .B(g5689), .Y(n9852));
NAND4X1  g5204(.A(n7026), .B(g5703), .C(g5571), .D(n9852), .Y(n9853));
NAND4X1  g5205(.A(g5603), .B(g5681), .C(g5689), .D(n5194), .Y(n9854));
NAND4X1  g5206(.A(g5654), .B(g5689), .C(g5543), .D(n7022_1), .Y(n9855));
AND2X1   g5207(.A(g5677), .B(g5689), .Y(n9856));
NAND4X1  g5208(.A(g5644), .B(n7019), .C(g5587), .D(n9856), .Y(n9857));
NAND4X1  g5209(.A(n9855), .B(n9854), .C(n9853), .D(n9857), .Y(n9858));
NAND4X1  g5210(.A(g5595), .B(g5677), .C(n9844), .D(n7022_1), .Y(n9859));
NAND3X1  g5211(.A(g5681), .B(n9844), .C(g5611), .Y(n9860));
OAI21X1  g5212(.A0(n9860), .A1(n7027_1), .B0(n9859), .Y(n9861));
NAND4X1  g5213(.A(g5685), .B(g5689), .C(g5551), .D(n7022_1), .Y(n9862));
NAND4X1  g5214(.A(g5619), .B(g5689), .C(g5630), .D(n5194), .Y(n9863));
NAND2X1  g5215(.A(n9863), .B(n9862), .Y(n9864));
NOR3X1   g5216(.A(n9864), .B(n9861), .C(n9858), .Y(n9865));
XOR2X1   g5217(.A(g5689), .B(n5871), .Y(n9866));
AND2X1   g5218(.A(g5666), .B(g5591), .Y(n9867));
AND2X1   g5219(.A(n9867), .B(n5194), .Y(n9868));
NAND3X1  g5220(.A(n7022_1), .B(g5637), .C(g5583), .Y(n9869));
NAND4X1  g5221(.A(n7026), .B(g5703), .C(g5666), .D(g5599), .Y(n9870));
AOI21X1  g5222(.A0(n9870), .A1(n9869), .B0(n9866), .Y(n9871));
AOI21X1  g5223(.A0(n9868), .A1(n9866), .B0(n9871), .Y(n9872));
NAND4X1  g5224(.A(n7019), .B(g5623), .C(g5615), .D(g5644), .Y(n9873));
NOR2X1   g5225(.A(n9873), .B(n9866), .Y(n9874));
NAND4X1  g5226(.A(g5563), .B(n9844), .C(g5659), .D(n5194), .Y(n9875));
NAND3X1  g5227(.A(g5685), .B(n9844), .C(g5567), .Y(n9876));
OAI21X1  g5228(.A0(n9876), .A1(n7020), .B0(n9875), .Y(n9877));
INVX1    g5229(.A(n9866), .Y(n9878));
NAND3X1  g5230(.A(n7022_1), .B(g5623), .C(g5607), .Y(n9879));
NAND4X1  g5231(.A(g5644), .B(n7019), .C(g5575), .D(g5637), .Y(n9880));
AOI21X1  g5232(.A0(n9880), .A1(n9879), .B0(n9878), .Y(n9881));
NOR3X1   g5233(.A(n9881), .B(n9877), .C(n9874), .Y(n9882));
NAND4X1  g5234(.A(n9872), .B(n9865), .C(n9851), .D(n9882), .Y(n9883));
AND2X1   g5235(.A(n9701), .B(g5462), .Y(n9884));
XOR2X1   g5236(.A(n9884), .B(n9883), .Y(n9885));
MX2X1    g5237(.A(g5462), .B(n9885), .S0(n7016), .Y(n9886));
MX2X1    g5238(.A(g5467), .B(n9886), .S0(g35), .Y(n5924));
MX2X1    g5239(.A(g2689), .B(n6708), .S0(n6435), .Y(n9888));
AND2X1   g5240(.A(n9888), .B(g35), .Y(n5929));
OAI21X1  g5241(.A0(n4856_1), .A1(n4855), .B0(g6573), .Y(n9890));
NAND3X1  g5242(.A(g6561), .B(g6565), .C(n4854), .Y(n9891));
AOI21X1  g5243(.A0(n9891), .A1(n9890), .B0(n7626), .Y(n9892));
MX2X1    g5244(.A(g6565), .B(n9892), .S0(g35), .Y(n5934));
NAND3X1  g5245(.A(g1612), .B(n7772), .C(n7397_1), .Y(n9894));
NAND3X1  g5246(.A(g1648), .B(n7772), .C(g1600), .Y(n9895));
AND2X1   g5247(.A(g1624), .B(g1657), .Y(n9896));
AOI22X1  g5248(.A0(n7398), .A1(g1608), .B0(g1604), .B1(n9896), .Y(n9897));
AND2X1   g5249(.A(n4629), .B(g1616), .Y(n9898));
AOI22X1  g5250(.A0(g25167), .A1(g1620), .B0(g1624), .B1(n9898), .Y(n9899));
NAND4X1  g5251(.A(n9897), .B(n9895), .C(n9894), .D(n9899), .Y(n9900));
MX2X1    g5252(.A(g1677), .B(n9900), .S0(n8992), .Y(n9901));
MX2X1    g5253(.A(g1657), .B(n9901), .S0(g35), .Y(n5939));
INVX1    g5254(.A(n7090), .Y(n9903));
OAI21X1  g5255(.A0(n9215), .A1(g2028), .B0(n4943), .Y(n9904));
OAI21X1  g5256(.A0(n6204), .A1(n4926), .B0(n9904), .Y(n9905));
MX2X1    g5257(.A(g2028), .B(n9905), .S0(n9903), .Y(n9906));
MX2X1    g5258(.A(g2036), .B(n9906), .S0(g35), .Y(n5944));
INVX1    g5259(.A(g2667), .Y(n9908));
XOR2X1   g5260(.A(g2661), .B(n9908), .Y(n9909));
MX2X1    g5261(.A(g2671), .B(n9909), .S0(n8533), .Y(n9910));
MX2X1    g5262(.A(g2667), .B(n9910), .S0(g35), .Y(n5949));
MX2X1    g5263(.A(g1576), .B(g1570), .S0(g1426), .Y(n9912));
MX2X1    g5264(.A(g1589), .B(n9912), .S0(g35), .Y(n5954));
INVX1    g5265(.A(g4375), .Y(n9914));
NOR2X1   g5266(.A(g4382), .B(n9914), .Y(n9915));
MX2X1    g5267(.A(n9915), .B(n8564), .S0(n6906_1), .Y(n9916));
MX2X1    g5268(.A(g4411), .B(n9916), .S0(g35), .Y(n5958));
XOR2X1   g5269(.A(n8442), .B(g1848), .Y(n9918));
MX2X1    g5270(.A(g1844), .B(n9918), .S0(g35), .Y(n5967));
AND2X1   g5271(.A(g3072), .B(g3080), .Y(n9920));
AND2X1   g5272(.A(n9920), .B(g3085), .Y(n9921));
XOR2X1   g5273(.A(n9921), .B(g3089), .Y(n9922));
MX2X1    g5274(.A(g3085), .B(n9922), .S0(g35), .Y(n5972));
INVX1    g5275(.A(n7355), .Y(n9924));
INVX1    g5276(.A(n7360), .Y(n9925));
MX2X1    g5277(.A(n9924), .B(n9925), .S0(n7358), .Y(n9926));
OR2X1    g5278(.A(n9926), .B(g3731), .Y(n9927));
NAND2X1  g5279(.A(n9926), .B(g3731), .Y(n9928));
OAI21X1  g5280(.A0(n9928), .A1(n7371), .B0(n9927), .Y(n9929));
MX2X1    g5281(.A(g3727), .B(n9929), .S0(g35), .Y(n5977));
AND2X1   g5282(.A(g5084), .B(g5092), .Y(n9931));
AND2X1   g5283(.A(n9931), .B(g5097), .Y(n9932));
XOR2X1   g5284(.A(n9932), .B(g86), .Y(n9933));
MX2X1    g5285(.A(g5097), .B(n9933), .S0(g35), .Y(n5982));
INVX1    g5286(.A(g5475), .Y(n9935));
XOR2X1   g5287(.A(g5481), .B(n9935), .Y(n9936));
MX2X1    g5288(.A(g5485), .B(n9936), .S0(n9702), .Y(n9937));
MX2X1    g5289(.A(g5481), .B(n9937), .S0(g35), .Y(n5987));
NOR2X1   g5290(.A(n7692), .B(n5508), .Y(n9939));
XOR2X1   g5291(.A(n9939), .B(n4909), .Y(n9940));
OAI22X1  g5292(.A0(n8854), .A1(n9940), .B0(n5508), .B1(g35), .Y(n5992));
NAND3X1  g5293(.A(g2575), .B(n6629), .C(n4934_1), .Y(n9942));
NAND3X1  g5294(.A(n6629), .B(g2610), .C(g2563), .Y(n9943));
AND2X1   g5295(.A(n9943), .B(n9942), .Y(n9944));
AND2X1   g5296(.A(g2587), .B(g2619), .Y(n9945));
AOI22X1  g5297(.A0(n8229), .A1(g2571), .B0(g2567), .B1(n9945), .Y(n9946));
NAND3X1  g5298(.A(g2583), .B(n4934_1), .C(g2610), .Y(n9947));
NAND3X1  g5299(.A(g2579), .B(g2587), .C(n5860_1), .Y(n9948));
NAND4X1  g5300(.A(n9947), .B(n9946), .C(n9944), .D(n9948), .Y(n9949));
MX2X1    g5301(.A(g2638), .B(n9949), .S0(n6628_1), .Y(n9950));
MX2X1    g5302(.A(g2619), .B(n9950), .S0(g35), .Y(n6000));
MX2X1    g5303(.A(g4145), .B(g4122), .S0(n7338), .Y(n9952));
MX2X1    g5304(.A(g4119), .B(n9952), .S0(g35), .Y(n6005));
AOI21X1  g5305(.A0(n6020_1), .A1(g4311), .B0(n5207), .Y(n9954));
NOR3X1   g5306(.A(n7471), .B(n4949_1), .C(g4322), .Y(n9955));
OAI21X1  g5307(.A0(n9955), .A1(n9954), .B0(n6256_1), .Y(n9956));
NAND2X1  g5308(.A(g4311), .B(n4620), .Y(n9957));
OAI21X1  g5309(.A0(n9956), .A1(n4620), .B0(n9957), .Y(n6010));
NOR4X1   g5310(.A(n6653_1), .B(n4862), .C(g5873), .D(g5857), .Y(n9959));
MX2X1    g5311(.A(g5941), .B(n5592_1), .S0(n9959), .Y(n9960));
MX2X1    g5312(.A(g5925), .B(n9960), .S0(g35), .Y(n6015));
MX2X1    g5313(.A(g2108), .B(g2102), .S0(n6086), .Y(n9962));
MX2X1    g5314(.A(g2102), .B(n9962), .S0(g35), .Y(n6020));
OR2X1    g5315(.A(g12), .B(g25), .Y(n6028));
NAND3X1  g5316(.A(n5506), .B(n5144), .C(g27831), .Y(n9965));
XOR2X1   g5317(.A(g25259), .B(g112), .Y(n9966));
MX2X1    g5318(.A(n9966), .B(g1644), .S0(n9965), .Y(n9967));
MX2X1    g5319(.A(g1592), .B(n9967), .S0(g35), .Y(n6033));
AOI21X1  g5320(.A0(g640), .A1(n6133), .B0(n5228), .Y(n9969));
MX2X1    g5321(.A(n5228), .B(n9969), .S0(n9043), .Y(n9970));
MX2X1    g5322(.A(g590), .B(n9970), .S0(g35), .Y(n6038));
OAI21X1  g5323(.A0(n6204), .A1(n4914), .B0(n5797_1), .Y(n9972));
MX2X1    g5324(.A(g2217), .B(n9972), .S0(n5788), .Y(n9973));
MX2X1    g5325(.A(g2223), .B(n9973), .S0(g35), .Y(n6043));
NOR3X1   g5326(.A(n8825), .B(g1395), .C(g1404), .Y(n9975));
NOR2X1   g5327(.A(g1570), .B(n8829), .Y(n9976));
OAI21X1  g5328(.A0(n9976), .A1(n9975), .B0(g1399), .Y(n9977));
MX2X1    g5329(.A(g1404), .B(n9977), .S0(g35), .Y(n6048));
NOR3X1   g5330(.A(n7090), .B(n6466), .C(n4926), .Y(n9979));
NOR2X1   g5331(.A(n4943), .B(g2051), .Y(n9980));
XOR2X1   g5332(.A(n9980), .B(g110), .Y(n9981));
MX2X1    g5333(.A(g2066), .B(n9981), .S0(n9979), .Y(n9982));
MX2X1    g5334(.A(g2051), .B(n9982), .S0(g35), .Y(n6053));
MX2X1    g5335(.A(g1152), .B(g1146), .S0(n6189), .Y(n9984));
MX2X1    g5336(.A(g1146), .B(n9984), .S0(g35), .Y(n6058));
NOR3X1   g5337(.A(n7933), .B(n6624), .C(g5164), .Y(n9986));
MX2X1    g5338(.A(g5252), .B(n5592_1), .S0(n9986), .Y(n9987));
MX2X1    g5339(.A(g5236), .B(n9987), .S0(g35), .Y(n6063));
MX2X1    g5340(.A(g2165), .B(n6705), .S0(n9122), .Y(n9990));
MX2X1    g5341(.A(g2246), .B(n9990), .S0(g35), .Y(n6068));
NOR3X1   g5342(.A(n6003), .B(g2629), .C(n7595_1), .Y(n9992));
MX2X1    g5343(.A(g2571), .B(n5998), .S0(n9992), .Y(n9993));
MX2X1    g5344(.A(g2563), .B(n9993), .S0(g35), .Y(n6073));
NOR4X1   g5345(.A(n6624), .B(g5176), .C(n5610), .D(n6042), .Y(n9995));
MX2X1    g5346(.A(g5170), .B(n9995), .S0(g35), .Y(n6078));
NAND2X1  g5347(.A(g901), .B(g35), .Y(n9997));
NAND2X1  g5348(.A(g901), .B(n4620), .Y(n9998));
NAND2X1  g5349(.A(n9998), .B(n9997), .Y(n6083));
AND2X1   g5350(.A(g2710), .B(n4620), .Y(n6092));
NAND4X1  g5351(.A(g1216), .B(g1087), .C(g1205), .D(g1221), .Y(n10001));
NOR2X1   g5352(.A(n7487), .B(g1211), .Y(n10002));
AND2X1   g5353(.A(n7486_1), .B(g1211), .Y(n10003));
MX2X1    g5354(.A(n10002), .B(n10003), .S0(n10001), .Y(n10004));
MX2X1    g5355(.A(g1216), .B(n10004), .S0(g35), .Y(n6100));
INVX1    g5356(.A(g2595), .Y(n10006));
AOI21X1  g5357(.A0(n7859), .A1(n10006), .B0(g2827), .Y(n10007));
OAI22X1  g5358(.A0(n7861), .A1(n10007), .B0(n7241), .B1(g35), .Y(n6105));
MX2X1    g5359(.A(n9176), .B(n9178), .S0(n9180), .Y(n10009));
OR2X1    g5360(.A(n10009), .B(g6423), .Y(n10010));
NAND2X1  g5361(.A(n10009), .B(g6423), .Y(n10011));
OAI21X1  g5362(.A0(n10011), .A1(n6884), .B0(n10010), .Y(n10012));
MX2X1    g5363(.A(g6419), .B(n10012), .S0(g35), .Y(n6110));
NAND4X1  g5364(.A(g4849), .B(g4854), .C(g4878), .D(g4843), .Y(n10014));
NOR2X1   g5365(.A(n10014), .B(g4859), .Y(n10015));
AND2X1   g5366(.A(n10014), .B(g4859), .Y(n10016));
OAI21X1  g5367(.A0(n10016), .A1(n10015), .B0(n9595), .Y(n10017));
NAND2X1  g5368(.A(g4854), .B(n4620), .Y(n10018));
OAI21X1  g5369(.A0(n10017), .A1(n4620), .B0(n10018), .Y(n6118));
MX2X1    g5370(.A(g424), .B(g411), .S0(n5688), .Y(n10020));
MX2X1    g5371(.A(g411), .B(n10020), .S0(g35), .Y(n6123));
AND2X1   g5372(.A(g1570), .B(g1274), .Y(n10022));
MX2X1    g5373(.A(n8876), .B(n10022), .S0(n8877), .Y(n10023));
MX2X1    g5374(.A(g1270), .B(n10023), .S0(g35), .Y(n6128));
OAI21X1  g5375(.A0(n5506), .A1(n7857), .B0(n5511_1), .Y(n10025));
OAI22X1  g5376(.A0(n6897), .A1(n10025), .B0(n5511_1), .B1(n5785), .Y(n10026));
MX2X1    g5377(.A(g2807), .B(n10026), .S0(g35), .Y(n6141));
INVX1    g5378(.A(g6439), .Y(n10028));
NAND3X1  g5379(.A(n6883), .B(n6882_1), .C(g35), .Y(n10029));
OAI21X1  g5380(.A0(n10028), .A1(g35), .B0(n10029), .Y(n6146));
MX2X1    g5381(.A(g1821), .B(g1816), .S0(n8442), .Y(n10031));
MX2X1    g5382(.A(g1816), .B(n10031), .S0(g35), .Y(n6151));
NOR2X1   g5383(.A(n7097), .B(n5524), .Y(n10033));
MX2X1    g5384(.A(n10033), .B(n7513), .S0(n7099), .Y(n10034));
OAI21X1  g5385(.A0(g2421), .A1(g2495), .B0(g2509), .Y(n10035));
XOR2X1   g5386(.A(n10035), .B(n10034), .Y(n10036));
MX2X1    g5387(.A(n10036), .B(g2509), .S0(n7100), .Y(n10037));
MX2X1    g5388(.A(g2495), .B(n10037), .S0(g35), .Y(n6156));
MX2X1    g5389(.A(g5069), .B(n5497_1), .S0(g35), .Y(n6161));
AND2X1   g5390(.A(g1570), .B(g1280), .Y(n10040));
MX2X1    g5391(.A(n9503), .B(n10040), .S0(n9504), .Y(n10041));
MX2X1    g5392(.A(g1266), .B(n10041), .S0(g35), .Y(n6166));
NOR4X1   g5393(.A(n4854), .B(n7204), .C(g6549), .D(g6565), .Y(n10043));
MX2X1    g5394(.A(g6633), .B(n5592_1), .S0(n10043), .Y(n10044));
MX2X1    g5395(.A(g6617), .B(n10044), .S0(g35), .Y(n6178));
XOR2X1   g5396(.A(g5115), .B(g5120), .Y(n10046));
MX2X1    g5397(.A(g5124), .B(n10046), .S0(n6440), .Y(n10047));
MX2X1    g5398(.A(g5115), .B(n10047), .S0(g35), .Y(n6183));
NOR4X1   g5399(.A(n4873), .B(n5980), .C(g6219), .D(n6208), .Y(n10049));
MX2X1    g5400(.A(g6303), .B(n5592_1), .S0(n10049), .Y(n10050));
MX2X1    g5401(.A(g6287), .B(n10050), .S0(g35), .Y(n6191));
NAND3X1  g5402(.A(n5500), .B(n5499), .C(g35), .Y(n10052));
OAI21X1  g5403(.A0(n5476), .A1(g35), .B0(n10052), .Y(n6196));
MX2X1    g5404(.A(g2994), .B(n5465), .S0(n8686), .Y(n10054));
MX2X1    g5405(.A(g2999), .B(n10054), .S0(g35), .Y(n6201));
MX2X1    g5406(.A(g681), .B(g650), .S0(n6389_1), .Y(n10056));
MX2X1    g5407(.A(g699), .B(n10056), .S0(g35), .Y(n6206));
NAND3X1  g5408(.A(n8425), .B(n7211), .C(g1592), .Y(n10058));
OAI21X1  g5409(.A0(n7211), .A1(n8175), .B0(n10058), .Y(n10059));
MX2X1    g5410(.A(g1644), .B(n10059), .S0(g35), .Y(n6211));
NOR4X1   g5411(.A(g3863), .B(g3881), .C(n4848), .D(n7642), .Y(n10061));
MX2X1    g5412(.A(g3921), .B(n5592_1), .S0(n10061), .Y(n10062));
MX2X1    g5413(.A(g3893), .B(n10062), .S0(g35), .Y(n6216));
INVX1    g5414(.A(g2093), .Y(n10064));
AOI21X1  g5415(.A0(g2051), .A1(n7088), .B0(n10064), .Y(n10065));
XOR2X1   g5416(.A(n10065), .B(g2079), .Y(n10066));
MX2X1    g5417(.A(n10066), .B(g2093), .S0(n7090), .Y(n10067));
MX2X1    g5418(.A(g2079), .B(n10067), .S0(g35), .Y(n6221));
NAND2X1  g5419(.A(n8967), .B(g35), .Y(n10069));
OAI22X1  g5420(.A0(n8538), .A1(n10069), .B0(n8537), .B1(g35), .Y(n6226));
NAND3X1  g5421(.A(g1514), .B(g1526), .C(g1500), .Y(n10071));
MX2X1    g5422(.A(g1339), .B(g1306), .S0(n10071), .Y(n10072));
MX2X1    g5423(.A(g1521), .B(n10072), .S0(g35), .Y(n6231));
NOR3X1   g5424(.A(n7983), .B(n6635), .C(n6647), .Y(n10074));
NOR3X1   g5425(.A(n6649), .B(g5373), .C(g5360), .Y(n10075));
OAI21X1  g5426(.A0(n10075), .A1(n10074), .B0(n7984), .Y(n10076));
NOR2X1   g5427(.A(n10075), .B(n10074), .Y(n10077));
NAND2X1  g5428(.A(n10077), .B(g5377), .Y(n10078));
OAI21X1  g5429(.A0(n10078), .A1(n6646), .B0(n10076), .Y(n10079));
MX2X1    g5430(.A(g5373), .B(n10079), .S0(g35), .Y(n6236));
NOR2X1   g5431(.A(n7084), .B(g1061), .Y(n10081));
OR4X1    g5432(.A(n4667_1), .B(n5691), .C(n7081), .D(n7082), .Y(n10082));
NAND3X1  g5433(.A(n10082), .B(n4666), .C(g35), .Y(n10083));
OAI22X1  g5434(.A0(n10081), .A1(n10083), .B0(n7081), .B1(g35), .Y(n6241));
MX2X1    g5435(.A(g3462), .B(g3498), .S0(n4836_1), .Y(n10085));
MX2X1    g5436(.A(g3498), .B(n10085), .S0(g35), .Y(n6246));
NOR3X1   g5437(.A(n7511_1), .B(g2197), .C(n5159), .Y(n10087));
MX2X1    g5438(.A(g2181), .B(n6705), .S0(n10087), .Y(n10088));
MX2X1    g5439(.A(g2169), .B(n10088), .S0(g35), .Y(n6251));
NOR4X1   g5440(.A(n6188), .B(g1183), .C(g1171), .D(n6397), .Y(n10090));
XOR2X1   g5441(.A(g1141), .B(g956), .Y(n10091));
MX2X1    g5442(.A(g956), .B(n10091), .S0(n10090), .Y(n10092));
MX2X1    g5443(.A(g1141), .B(n10092), .S0(g35), .Y(n6256));
NOR3X1   g5444(.A(n5628), .B(g1772), .C(n5164), .Y(n10094));
MX2X1    g5445(.A(g1756), .B(n5624), .S0(n10094), .Y(n10095));
MX2X1    g5446(.A(g1744), .B(n10095), .S0(g35), .Y(n6261));
INVX1    g5447(.A(g5849), .Y(n10097));
OAI22X1  g5448(.A0(n5524), .A1(g4284), .B0(n10097), .B1(n4863), .Y(n10098));
OR4X1    g5449(.A(n5524), .B(g4284), .C(n10097), .D(n4863), .Y(n10099));
AOI21X1  g5450(.A0(n10099), .A1(n10098), .B0(n4620), .Y(n6266));
NAND4X1  g5451(.A(n4726), .B(n4731_1), .C(n4729), .D(n6252), .Y(n10101));
MX2X1    g5452(.A(g4145), .B(g4112), .S0(n10101), .Y(n10102));
MX2X1    g5453(.A(g4145), .B(n10102), .S0(g35), .Y(n6271));
INVX1    g5454(.A(g2675), .Y(n10104));
XOR2X1   g5455(.A(g2681), .B(n10104), .Y(n10105));
NOR3X1   g5456(.A(n5863), .B(n6629), .C(n4934_1), .Y(n10106));
MX2X1    g5457(.A(g2685), .B(n10105), .S0(n10106), .Y(n10107));
MX2X1    g5458(.A(g2681), .B(n10107), .S0(g35), .Y(n6276));
NAND3X1  g5459(.A(n8913), .B(n7512), .C(g2153), .Y(n10109));
OAI21X1  g5460(.A0(n7512), .A1(n9740), .B0(n10109), .Y(n10110));
MX2X1    g5461(.A(g2204), .B(n10110), .S0(g35), .Y(n6281));
INVX1    g5462(.A(g6113), .Y(n10112));
NOR2X1   g5463(.A(g6109), .B(n10112), .Y(n10113));
NOR2X1   g5464(.A(g6105), .B(n10112), .Y(n10114));
MX2X1    g5465(.A(n10113), .B(n10114), .S0(g6120), .Y(n10115));
MX2X1    g5466(.A(g6113), .B(n10115), .S0(g35), .Y(n6286));
NAND3X1  g5467(.A(n7099), .B(n7096), .C(g2421), .Y(n10117));
AOI21X1  g5468(.A0(n7681), .A1(g2465), .B0(g2495), .Y(n10118));
NAND3X1  g5469(.A(n10118), .B(n7102), .C(n7101), .Y(n10119));
AOI21X1  g5470(.A0(n10119), .A1(n10117), .B0(n4620), .Y(n6291));
OR4X1    g5471(.A(n7900), .B(g1046), .C(n6049), .D(n7901), .Y(n10121));
OAI21X1  g5472(.A0(n7901), .A1(n7900), .B0(g1046), .Y(n10122));
NAND2X1  g5473(.A(n10122), .B(n10121), .Y(n10123));
MX2X1    g5474(.A(g1041), .B(n10123), .S0(g35), .Y(n6296));
OAI21X1  g5475(.A0(g686), .A1(n5876), .B0(n5130_1), .Y(n10125));
OAI21X1  g5476(.A0(g686), .A1(n5876), .B0(g482), .Y(n10126));
MX2X1    g5477(.A(n10125), .B(n10126), .S0(n5883), .Y(n10127));
MX2X1    g5478(.A(g528), .B(n10127), .S0(g35), .Y(n6301));
INVX1    g5479(.A(g4405), .Y(n10129));
NAND3X1  g5480(.A(n6906_1), .B(n8564), .C(g4388), .Y(n10130));
OAI21X1  g5481(.A0(n10130), .A1(n4620), .B0(n10129), .Y(n6306));
MX2X1    g5482(.A(n9462), .B(n9463), .S0(n6875), .Y(n10132));
NOR2X1   g5483(.A(n6884), .B(n6876), .Y(n10133));
MX2X1    g5484(.A(n6876), .B(n10133), .S0(n10132), .Y(n10134));
MX2X1    g5485(.A(g6428), .B(n10134), .S0(g35), .Y(n6311));
OAI21X1  g5486(.A0(n8333), .A1(g1514), .B0(n8329), .Y(n10136));
OAI21X1  g5487(.A0(n8333), .A1(n5549), .B0(g1500), .Y(n10137));
AOI21X1  g5488(.A0(n10137), .A1(n10136), .B0(n4620), .Y(n6316));
NAND2X1  g5489(.A(g319), .B(g35), .Y(n10139));
NAND2X1  g5490(.A(g319), .B(n4620), .Y(n10140));
NAND2X1  g5491(.A(n10140), .B(n10139), .Y(n6321));
NAND2X1  g5492(.A(g6561), .B(n4855), .Y(n10142));
NAND2X1  g5493(.A(n4856_1), .B(g6565), .Y(n10143));
AOI21X1  g5494(.A0(n10143), .A1(n10142), .B0(n7626), .Y(n10144));
MX2X1    g5495(.A(g6561), .B(n10144), .S0(g35), .Y(n6326));
MX2X1    g5496(.A(g2950), .B(n2447), .S0(n5617), .Y(n10146));
MX2X1    g5497(.A(g2936), .B(n10146), .S0(g35), .Y(n6331));
MX2X1    g5498(.A(g4164), .B(g4129), .S0(n10101), .Y(n10148));
MX2X1    g5499(.A(g4164), .B(n10148), .S0(g35), .Y(n6336));
MX2X1    g5500(.A(g1345), .B(n7290), .S0(n5986), .Y(n10150));
MX2X1    g5501(.A(g1351), .B(n10150), .S0(g35), .Y(n6341));
MX2X1    g5502(.A(g6533), .B(g6527), .S0(n4857), .Y(n10152));
MX2X1    g5503(.A(g6527), .B(n10152), .S0(g35), .Y(n6346));
XOR2X1   g5504(.A(n9920), .B(g3085), .Y(n10154));
MX2X1    g5505(.A(g3080), .B(n10154), .S0(g35), .Y(n6355));
MX2X1    g5506(.A(g4727), .B(n3747), .S0(n6494), .Y(n10156));
AND2X1   g5507(.A(n10156), .B(g35), .Y(n6360));
INVX1    g5508(.A(g6661), .Y(n10158));
OAI22X1  g5509(.A0(g6704), .A1(n10158), .B0(g6697), .B1(n6678), .Y(n10159));
MX2X1    g5510(.A(g6692), .B(n10158), .S0(g6668), .Y(n10160));
OAI21X1  g5511(.A0(n6679), .A1(g6675), .B0(g35), .Y(n10161));
NOR4X1   g5512(.A(n10160), .B(n10159), .C(n6681_1), .D(n10161), .Y(n6365));
OR2X1    g5513(.A(n8332), .B(g1536), .Y(n10163));
NOR3X1   g5514(.A(n8339), .B(n8338), .C(n8334), .Y(n10164));
OAI21X1  g5515(.A0(n10164), .A1(n4711), .B0(n10163), .Y(n10165));
MX2X1    g5516(.A(g1532), .B(n10165), .S0(g35), .Y(n6369));
NOR4X1   g5517(.A(n7041), .B(n4850), .C(g3873), .D(g3857), .Y(n10167));
MX2X1    g5518(.A(g3941), .B(n5592_1), .S0(n10167), .Y(n10168));
MX2X1    g5519(.A(g3925), .B(n10168), .S0(g35), .Y(n6374));
XOR2X1   g5520(.A(n6178_1), .B(g370), .Y(n10170));
MX2X1    g5521(.A(g358), .B(n10170), .S0(g35), .Y(n6379));
AND2X1   g5522(.A(n5873), .B(g5689), .Y(n10172));
NAND2X1  g5523(.A(n7024), .B(g35), .Y(n10173));
OAI22X1  g5524(.A0(n10172), .A1(n10173), .B0(n9844), .B1(g35), .Y(n6384));
INVX1    g5525(.A(g1854), .Y(n10175));
XOR2X1   g5526(.A(g1848), .B(n10175), .Y(n10176));
MX2X1    g5527(.A(g1858), .B(n10176), .S0(n9288), .Y(n10177));
MX2X1    g5528(.A(g1854), .B(n10177), .S0(g35), .Y(n6389));
MX2X1    g5529(.A(g446), .B(g872), .S0(n7408), .Y(n10179));
MX2X1    g5530(.A(g246), .B(n10179), .S0(g35), .Y(n6394));
AND2X1   g5531(.A(g4931), .B(n4620), .Y(n6399));
NOR4X1   g5532(.A(n4845), .B(g3179), .C(n5913), .D(g3161), .Y(n10182));
MX2X1    g5533(.A(g3219), .B(n5592_1), .S0(n10182), .Y(n10183));
MX2X1    g5534(.A(g3191), .B(n10183), .S0(g35), .Y(n6404));
NAND3X1  g5535(.A(n4941), .B(n9287), .C(g1748), .Y(n10185));
NAND3X1  g5536(.A(g1783), .B(n9287), .C(g1736), .Y(n10186));
AND2X1   g5537(.A(n10186), .B(n10185), .Y(n10187));
AND2X1   g5538(.A(g1792), .B(g1760), .Y(n10188));
AOI22X1  g5539(.A0(n6470), .A1(g1744), .B0(g1740), .B1(n10188), .Y(n10189));
NAND3X1  g5540(.A(n4941), .B(g1756), .C(g1783), .Y(n10190));
NAND3X1  g5541(.A(n8135), .B(g1760), .C(g1752), .Y(n10191));
NAND4X1  g5542(.A(n10190), .B(n10189), .C(n10187), .D(n10191), .Y(n10192));
MX2X1    g5543(.A(g1811), .B(n10192), .S0(n8134), .Y(n10193));
MX2X1    g5544(.A(g1792), .B(n10193), .S0(g35), .Y(n6409));
XOR2X1   g5545(.A(g3431), .B(g3423), .Y(n10195));
MX2X1    g5546(.A(g3423), .B(n10195), .S0(g35), .Y(n6414));
NOR4X1   g5547(.A(g6561), .B(g6555), .C(g6549), .D(n7205), .Y(n10197));
MX2X1    g5548(.A(g6601), .B(n5592_1), .S0(n10197), .Y(n10198));
MX2X1    g5549(.A(g6605), .B(n10198), .S0(g35), .Y(n6419));
NAND3X1  g5550(.A(n6415), .B(n6413), .C(g3376), .Y(n10200));
OAI21X1  g5551(.A0(n6414_1), .A1(n6412), .B0(n6409_1), .Y(n10201));
OAI21X1  g5552(.A0(n10200), .A1(n5778_1), .B0(n10201), .Y(n10202));
MX2X1    g5553(.A(g3372), .B(n10202), .S0(g35), .Y(n6424));
NOR3X1   g5554(.A(n7100), .B(n7681), .C(n5151), .Y(n10204));
MX2X1    g5555(.A(g2441), .B(n7132_1), .S0(n10204), .Y(n10205));
MX2X1    g5556(.A(g2445), .B(n10205), .S0(g35), .Y(n6429));
MX2X1    g5557(.A(g1874), .B(n5526_1), .S0(n9112), .Y(n10208));
MX2X1    g5558(.A(g1955), .B(n10208), .S0(g35), .Y(n6434));
NOR4X1   g5559(.A(n5713_1), .B(g4639), .C(n5848), .D(n6018), .Y(n10210));
NAND3X1  g5560(.A(n10210), .B(n5845_1), .C(n5174), .Y(n10211));
INVX1    g5561(.A(n10210), .Y(n10212));
NAND3X1  g5562(.A(n10212), .B(n5845_1), .C(g4349), .Y(n10213));
NAND2X1  g5563(.A(n10213), .B(n10211), .Y(n10214));
MX2X1    g5564(.A(g4340), .B(n10214), .S0(g35), .Y(n6439));
NOR4X1   g5565(.A(g6561), .B(g6555), .C(g6549), .D(n7657), .Y(n10216));
MX2X1    g5566(.A(g6581), .B(n5592_1), .S0(n10216), .Y(n10217));
MX2X1    g5567(.A(g6573), .B(n10217), .S0(g35), .Y(n6444));
NOR3X1   g5568(.A(n4856_1), .B(n4855), .C(g6573), .Y(n10219));
MX2X1    g5569(.A(g6597), .B(n5592_1), .S0(n10219), .Y(n10220));
MX2X1    g5570(.A(g6645), .B(n10220), .S0(g35), .Y(n6449));
NOR4X1   g5571(.A(n4833), .B(n5735), .C(n5733_1), .D(n4835), .Y(n10222));
MX2X1    g5572(.A(g3610), .B(n5592_1), .S0(n10222), .Y(n10223));
MX2X1    g5573(.A(g3594), .B(n10223), .S0(g35), .Y(n6458));
OAI21X1  g5574(.A0(g2890), .A1(n9189), .B0(g35), .Y(n10225));
AOI21X1  g5575(.A0(n8686), .A1(n3220), .B0(n10225), .Y(n10226));
AND2X1   g5576(.A(g2873), .B(n4620), .Y(n10227));
OR2X1    g5577(.A(n10227), .B(n10226), .Y(n6463));
INVX1    g5578(.A(g1968), .Y(n10229));
XOR2X1   g5579(.A(g1974), .B(n10229), .Y(n10230));
MX2X1    g5580(.A(g1978), .B(n10230), .S0(n9112), .Y(n10231));
MX2X1    g5581(.A(g1974), .B(n10231), .S0(g35), .Y(n6468));
NOR3X1   g5582(.A(n5758_1), .B(n5757), .C(n4631), .Y(n10233));
MX2X1    g5583(.A(g1612), .B(n5756), .S0(n10233), .Y(n10234));
MX2X1    g5584(.A(g1616), .B(n10234), .S0(g35), .Y(n6473));
NAND2X1  g5585(.A(n5169), .B(n5150), .Y(n10236));
OAI21X1  g5586(.A0(n5170), .A1(n5150), .B0(n10236), .Y(n6478));
NOR3X1   g5587(.A(n5468), .B(n5217), .C(n5616), .Y(n10238));
OAI21X1  g5588(.A0(n6171), .A1(g2856), .B0(g35), .Y(n10239));
OAI22X1  g5589(.A0(n10238), .A1(n10239), .B0(n5216_1), .B1(g35), .Y(n6483));
XOR2X1   g5590(.A(n7106), .B(g6479), .Y(n10241));
MX2X1    g5591(.A(g6474), .B(n10241), .S0(g35), .Y(n6488));
XOR2X1   g5592(.A(n9112), .B(g1982), .Y(n10243));
MX2X1    g5593(.A(g1978), .B(n10243), .S0(g35), .Y(n6493));
NOR4X1   g5594(.A(g5188), .B(n5610), .C(n4642_1), .D(g5170), .Y(n10245));
MX2X1    g5595(.A(g5228), .B(n5592_1), .S0(n10245), .Y(n10246));
MX2X1    g5596(.A(g5200), .B(n10246), .S0(g35), .Y(n6502));
MX2X1    g5597(.A(g4145), .B(g4119), .S0(n6939), .Y(n10248));
MX2X1    g5598(.A(g4116), .B(n10248), .S0(g35), .Y(n6507));
AOI21X1  g5599(.A0(n6999), .A1(g35), .B0(n9127), .Y(n6512));
OR2X1    g5600(.A(n8336), .B(n8338), .Y(n10251));
OR4X1    g5601(.A(n7601), .B(g1542), .C(n8329), .D(n8335), .Y(n10252));
AOI21X1  g5602(.A0(n10252), .A1(n10251), .B0(n8333), .Y(n10253));
MX2X1    g5603(.A(g1536), .B(n10253), .S0(g35), .Y(n6517));
NOR2X1   g5604(.A(g4258), .B(n4620), .Y(n6522));
NOR3X1   g5605(.A(n5482_1), .B(n5480), .C(n5479), .Y(n10256));
NOR3X1   g5606(.A(g5016), .B(g5029), .C(n5488), .Y(n10257));
OAI21X1  g5607(.A0(n10257), .A1(n10256), .B0(n5481), .Y(n10258));
NOR2X1   g5608(.A(n10257), .B(n10256), .Y(n10259));
NAND2X1  g5609(.A(n10259), .B(g5033), .Y(n10260));
OAI21X1  g5610(.A0(n10260), .A1(n5501), .B0(n10258), .Y(n10261));
MX2X1    g5611(.A(g5029), .B(n10261), .S0(g35), .Y(n6531));
MX2X1    g5612(.A(g4717), .B(n4447), .S0(n6494), .Y(n10263));
MX2X1    g5613(.A(g4732), .B(n10263), .S0(g35), .Y(n6536));
INVX1    g5614(.A(g1559), .Y(n10265));
NOR3X1   g5615(.A(n7669), .B(n10265), .C(n7667), .Y(n10266));
NAND4X1  g5616(.A(g1559), .B(n7668), .C(g1564), .D(n7520_1), .Y(n10267));
OAI21X1  g5617(.A0(n7669), .A1(n7667), .B0(g1554), .Y(n10268));
OAI21X1  g5618(.A0(n10268), .A1(n10266), .B0(n10267), .Y(n10269));
MX2X1    g5619(.A(g1559), .B(n10269), .S0(g35), .Y(n6541));
INVX1    g5620(.A(g3849), .Y(n10271));
OAI22X1  g5621(.A0(n5524), .A1(g4284), .B0(n10271), .B1(n4851_1), .Y(n10272));
OR4X1    g5622(.A(n5524), .B(g4284), .C(n10271), .D(n4851_1), .Y(n10273));
AOI21X1  g5623(.A0(n10273), .A1(n10272), .B0(n4620), .Y(n6546));
NOR3X1   g5624(.A(g3161), .B(g3167), .C(g3155), .Y(n10275));
NAND3X1  g5625(.A(n10275), .B(n4845), .C(g3179), .Y(n10276));
MX2X1    g5626(.A(n5592_1), .B(g3199), .S0(n10276), .Y(n10277));
MX2X1    g5627(.A(g3203), .B(n10277), .S0(g35), .Y(n6555));
INVX1    g5628(.A(g5835), .Y(n10279));
XOR2X1   g5629(.A(g5841), .B(n10279), .Y(n10280));
MX2X1    g5630(.A(g5845), .B(n10280), .S0(n4863), .Y(n10281));
MX2X1    g5631(.A(g5841), .B(n10281), .S0(g35), .Y(n6560));
NAND3X1  g5632(.A(n6777_1), .B(n6192), .C(n4896_1), .Y(n10283));
NAND3X1  g5633(.A(n6778), .B(n6192), .C(g4975), .Y(n10284));
NAND2X1  g5634(.A(n10284), .B(n10283), .Y(n10285));
MX2X1    g5635(.A(g4966), .B(n10285), .S0(g35), .Y(n6565));
INVX1    g5636(.A(n9500), .Y(n10287));
OR2X1    g5637(.A(n10287), .B(n5680), .Y(n10288));
AOI21X1  g5638(.A0(g802), .A1(n5662), .B0(n5408), .Y(n10289));
MX2X1    g5639(.A(n5408), .B(n10289), .S0(n10288), .Y(n10290));
MX2X1    g5640(.A(g785), .B(n10290), .S0(g35), .Y(n6570));
NOR3X1   g5641(.A(n4862), .B(n4861_1), .C(g5873), .Y(n10292));
MX2X1    g5642(.A(g5913), .B(n5592_1), .S0(n10292), .Y(n10293));
MX2X1    g5643(.A(g5957), .B(n10293), .S0(g35), .Y(n6575));
NOR4X1   g5644(.A(n5569), .B(n6203), .C(g1926), .D(n5840), .Y(n10295));
MX2X1    g5645(.A(g1902), .B(n9549), .S0(n10295), .Y(n10296));
MX2X1    g5646(.A(g1882), .B(n10296), .S0(g35), .Y(n6580));
XOR2X1   g5647(.A(g6159), .B(g6154), .Y(n10298));
MX2X1    g5648(.A(g6163), .B(n10298), .S0(n5910), .Y(n10299));
MX2X1    g5649(.A(g6154), .B(n10299), .S0(g35), .Y(n6585));
OAI22X1  g5650(.A0(g4125), .A1(n7727), .B0(n8547), .B1(g35), .Y(n6590));
MX2X1    g5651(.A(g4821), .B(n9883), .S0(n7016), .Y(n10302));
MX2X1    g5652(.A(g5619), .B(n10302), .S0(g35), .Y(n6595));
INVX1    g5653(.A(g4939), .Y(n10304));
OR2X1    g5654(.A(n7756), .B(n10304), .Y(n10305));
OAI21X1  g5655(.A0(n8626), .A1(n9144), .B0(n10304), .Y(n10306));
NAND2X1  g5656(.A(n8633), .B(n9144), .Y(n10307));
MX2X1    g5657(.A(n5184), .B(n8621), .S0(n6829), .Y(n10308));
NAND2X1  g5658(.A(n10308), .B(n10307), .Y(n10309));
NOR4X1   g5659(.A(n6806), .B(g4975), .C(g4899), .D(n7757), .Y(n10310));
OAI21X1  g5660(.A0(n10309), .A1(n10306), .B0(n10310), .Y(n10311));
AOI21X1  g5661(.A0(n10311), .A1(n10305), .B0(n4620), .Y(n6600));
INVX1    g5662(.A(g990), .Y(n10313));
XOR2X1   g5663(.A(n8511), .B(n10313), .Y(n10314));
MX2X1    g5664(.A(g990), .B(n10314), .S0(g35), .Y(n6605));
NOR4X1   g5665(.A(g3161), .B(g3167), .C(g3155), .D(n5594), .Y(n10316));
MX2X1    g5666(.A(g3207), .B(n5592_1), .S0(n10316), .Y(n10317));
MX2X1    g5667(.A(g3211), .B(n10317), .S0(g35), .Y(n6609));
NOR3X1   g5668(.A(n5594), .B(n5593), .C(n5913), .Y(n10319));
MX2X1    g5669(.A(g3259), .B(n5592_1), .S0(n10319), .Y(n10320));
MX2X1    g5670(.A(g3243), .B(n10320), .S0(g35), .Y(n6618));
XOR2X1   g5671(.A(n6440), .B(g5142), .Y(n10322));
MX2X1    g5672(.A(g5138), .B(n10322), .S0(g35), .Y(n6623));
NOR4X1   g5673(.A(n4643), .B(g5164), .C(g5180), .D(n6624), .Y(n10324));
MX2X1    g5674(.A(g5248), .B(n5592_1), .S0(n10324), .Y(n10325));
MX2X1    g5675(.A(g5232), .B(n10325), .S0(g35), .Y(n6628));
INVX1    g5676(.A(g2122), .Y(n10327));
XOR2X1   g5677(.A(g2116), .B(n10327), .Y(n10328));
MX2X1    g5678(.A(g2126), .B(n10328), .S0(n7091), .Y(n10329));
MX2X1    g5679(.A(g2122), .B(n10329), .S0(g35), .Y(n6633));
NAND2X1  g5680(.A(n8202), .B(g35), .Y(n10331));
OAI22X1  g5681(.A0(n5807_1), .A1(n10331), .B0(n5805), .B1(g35), .Y(n6638));
MX2X1    g5682(.A(g5481), .B(g5475), .S0(n9702), .Y(n10333));
MX2X1    g5683(.A(g5475), .B(n10333), .S0(g35), .Y(n6643));
XOR2X1   g5684(.A(g1955), .B(g1959), .Y(n10335));
NOR4X1   g5685(.A(n5569), .B(g1894), .C(n6203), .D(n5840), .Y(n10336));
MX2X1    g5686(.A(g1964), .B(n10335), .S0(n10336), .Y(n10337));
MX2X1    g5687(.A(g1959), .B(n10337), .S0(g35), .Y(n6648));
XOR2X1   g5688(.A(n9931), .B(g5097), .Y(n10339));
MX2X1    g5689(.A(g5092), .B(n10339), .S0(g35), .Y(n6653));
NOR3X1   g5690(.A(n7506_1), .B(g3161), .C(n5913), .Y(n10341));
MX2X1    g5691(.A(g3215), .B(n5592_1), .S0(n10341), .Y(n10342));
MX2X1    g5692(.A(g3187), .B(n10342), .S0(g35), .Y(n6658));
INVX1    g5693(.A(g4430), .Y(n10344));
INVX1    g5694(.A(g4434), .Y(n10345));
AOI22X1  g5695(.A0(n10345), .A1(g4401), .B0(n10344), .B1(g4388), .Y(n10346));
INVX1    g5696(.A(g4388), .Y(n10347));
INVX1    g5697(.A(g4401), .Y(n10348));
AOI22X1  g5698(.A0(g4434), .A1(n10348), .B0(g4430), .B1(n10347), .Y(n10349));
NAND2X1  g5699(.A(n10349), .B(n10346), .Y(n10350));
MX2X1    g5700(.A(g4430), .B(n10350), .S0(g35), .Y(n6671));
INVX1    g5701(.A(g1768), .Y(n10352));
AOI21X1  g5702(.A0(n7859), .A1(n10352), .B0(g2779), .Y(n10353));
OAI22X1  g5703(.A0(n7861), .A1(n10353), .B0(n5512), .B1(g35), .Y(n6681));
INVX1    g5704(.A(g4438), .Y(n10355));
NOR2X1   g5705(.A(n10355), .B(g4382), .Y(n10356));
MX2X1    g5706(.A(n10356), .B(n8564), .S0(n7415), .Y(n10357));
MX2X1    g5707(.A(g4443), .B(n10357), .S0(g35), .Y(n6690));
MX2X1    g5708(.A(g1720), .B(g1714), .S0(n7773), .Y(n10359));
MX2X1    g5709(.A(g1714), .B(n10359), .S0(g35), .Y(n6694));
NOR2X1   g5710(.A(n8213), .B(n7289), .Y(n10361));
MX2X1    g5711(.A(g1367), .B(n7288_1), .S0(n10361), .Y(n10362));
MX2X1    g5712(.A(g1361), .B(n10362), .S0(g35), .Y(n6699));
MX2X1    g5713(.A(g4104), .B(n6267), .S0(g35), .Y(n6713));
NOR3X1   g5714(.A(n7511_1), .B(g2197), .C(n6708_1), .Y(n10365));
MX2X1    g5715(.A(g2161), .B(n6705), .S0(n10365), .Y(n10366));
MX2X1    g5716(.A(g2165), .B(n10366), .S0(g35), .Y(n6718));
XOR2X1   g5717(.A(g376), .B(g358), .Y(n10368));
MX2X1    g5718(.A(g370), .B(n10368), .S0(g35), .Y(n6723));
NAND3X1  g5719(.A(n6730), .B(n6729), .C(g2331), .Y(n10370));
OAI21X1  g5720(.A0(n6729), .A1(n5154), .B0(n10370), .Y(n10371));
MX2X1    g5721(.A(g2331), .B(n10371), .S0(g35), .Y(n6728));
NOR3X1   g5722(.A(g4191), .B(g4200), .C(g4197), .Y(n10373));
NOR2X1   g5723(.A(g4204), .B(g4207), .Y(n10374));
NOR4X1   g5724(.A(g4194), .B(g4210), .C(g4188), .D(g4180), .Y(n10375));
NAND3X1  g5725(.A(n10375), .B(n10374), .C(n10373), .Y(n10376));
XOR2X1   g5726(.A(n5524), .B(g4200), .Y(n10377));
NAND2X1  g5727(.A(n10377), .B(n10376), .Y(n10378));
MX2X1    g5728(.A(g2946), .B(n10378), .S0(g35), .Y(n6733));
MX2X1    g5729(.A(n9042), .B(n5322_1), .S0(n9041), .Y(n10380));
MX2X1    g5730(.A(g577), .B(n10380), .S0(g35), .Y(n6737));
OAI21X1  g5731(.A0(n6204), .A1(n4926), .B0(n7088), .Y(n10382));
MX2X1    g5732(.A(g2051), .B(n10382), .S0(n9903), .Y(n10383));
MX2X1    g5733(.A(g2028), .B(n10383), .S0(g35), .Y(n6742));
OR2X1    g5734(.A(n6760), .B(g1193), .Y(n10385));
NOR3X1   g5735(.A(n7149), .B(n7148), .C(n7144), .Y(n10386));
OAI21X1  g5736(.A0(n10386), .A1(n4707_1), .B0(n10385), .Y(n10387));
MX2X1    g5737(.A(g1189), .B(n10387), .S0(g35), .Y(n6747));
MX2X1    g5738(.A(n8404), .B(n8406), .S0(n6637), .Y(n10389));
NOR2X1   g5739(.A(n6646), .B(n8979), .Y(n10390));
MX2X1    g5740(.A(n10390), .B(n8979), .S0(n10389), .Y(n10391));
MX2X1    g5741(.A(g5396), .B(n10391), .S0(g35), .Y(n6752));
NAND3X1  g5742(.A(n5777), .B(n5776), .C(g35), .Y(n10393));
OAI21X1  g5743(.A0(n8675), .A1(g35), .B0(n10393), .Y(n6757));
NAND3X1  g5744(.A(n7227), .B(n4932), .C(g2342), .Y(n10395));
MX2X1    g5745(.A(n8366), .B(g2327), .S0(n10395), .Y(n10396));
MX2X1    g5746(.A(g2307), .B(n10396), .S0(g35), .Y(n6762));
AND2X1   g5747(.A(g907), .B(g1227), .Y(n10398));
MX2X1    g5748(.A(n6452), .B(n10398), .S0(n6453_1), .Y(n10399));
MX2X1    g5749(.A(g936), .B(n10399), .S0(g35), .Y(n6767));
OAI21X1  g5750(.A0(n6316_1), .A1(n5616), .B0(g947), .Y(n10401));
OR4X1    g5751(.A(n5024), .B(n5004), .C(n5616), .D(n5462), .Y(n10402));
AOI21X1  g5752(.A0(n10402), .A1(n10401), .B0(n4620), .Y(n6772));
XOR2X1   g5753(.A(n9288), .B(g1834), .Y(n10404));
MX2X1    g5754(.A(g1830), .B(n10404), .S0(g35), .Y(n6777));
NOR4X1   g5755(.A(n4833), .B(g3506), .C(n5733_1), .D(n4835), .Y(n10406));
MX2X1    g5756(.A(g3594), .B(n5592_1), .S0(n10406), .Y(n10407));
MX2X1    g5757(.A(g3578), .B(n10407), .S0(g35), .Y(n6782));
OAI21X1  g5758(.A0(g2999), .A1(g2932), .B0(g35), .Y(n10409));
AOI21X1  g5759(.A0(n8686), .A1(n6676), .B0(n10409), .Y(n6787));
NAND3X1  g5760(.A(n9687), .B(n9686), .C(g5727), .Y(n10411));
OAI21X1  g5761(.A0(n7066), .A1(n7061), .B0(n7064), .Y(n10412));
OAI21X1  g5762(.A0(n10411), .A1(n7077), .B0(n10412), .Y(n10413));
MX2X1    g5763(.A(g5723), .B(n10413), .S0(g35), .Y(n6792));
NOR3X1   g5764(.A(n5552), .B(g2361), .C(n9673), .Y(n10415));
MX2X1    g5765(.A(g2303), .B(n5547), .S0(n10415), .Y(n10416));
MX2X1    g5766(.A(g2295), .B(n10416), .S0(g35), .Y(n6797));
INVX1    g5767(.A(g3057), .Y(n10418));
AOI21X1  g5768(.A0(n10418), .A1(g35), .B0(n9102), .Y(n6805));
OAI21X1  g5769(.A0(n5688), .A1(n6229), .B0(n6389_1), .Y(n10420));
MX2X1    g5770(.A(g681), .B(n10420), .S0(g35), .Y(n6810));
OR4X1    g5771(.A(n8696), .B(n7153), .C(n7160), .D(n7154), .Y(n10422));
NOR2X1   g5772(.A(n7158), .B(g723), .Y(n10423));
INVX1    g5773(.A(g723), .Y(n10424));
NOR2X1   g5774(.A(n7158), .B(n10424), .Y(n10425));
MX2X1    g5775(.A(n10423), .B(n10425), .S0(n10422), .Y(n10426));
MX2X1    g5776(.A(g827), .B(n10426), .S0(g35), .Y(n6815));
AND2X1   g5777(.A(n7016), .B(n9274), .Y(n10428));
NAND4X1  g5778(.A(n4957), .B(n5181_1), .C(g4349), .D(n10428), .Y(n10429));
NAND3X1  g5779(.A(n10429), .B(n7016), .C(n7019), .Y(n10430));
OAI21X1  g5780(.A0(n7016), .A1(n7019), .B0(n10430), .Y(n10431));
MX2X1    g5781(.A(g5698), .B(n10431), .S0(g35), .Y(n6820));
NOR3X1   g5782(.A(n5465), .B(n5226_1), .C(n5616), .Y(n10433));
OAI21X1  g5783(.A0(n5516_1), .A1(g546), .B0(g35), .Y(n10434));
OAI22X1  g5784(.A0(n10433), .A1(n10434), .B0(n5225), .B1(g35), .Y(n6825));
NOR4X1   g5785(.A(n6466), .B(n5137), .C(n5136), .D(n7096), .Y(n10436));
XOR2X1   g5786(.A(n5152), .B(g112), .Y(n10437));
MX2X1    g5787(.A(g2472), .B(n10437), .S0(n10436), .Y(n10438));
MX2X1    g5788(.A(g2421), .B(n10438), .S0(g35), .Y(n6830));
NOR4X1   g5789(.A(n6653_1), .B(g5881), .C(n4860), .D(n7375), .Y(n10440));
MX2X1    g5790(.A(g5953), .B(n5592_1), .S0(n10440), .Y(n10441));
MX2X1    g5791(.A(g5937), .B(n10441), .S0(g35), .Y(n6835));
MX2X1    g5792(.A(g3050), .B(g3338), .S0(g35), .Y(n6840));
NOR3X1   g5793(.A(n9462), .B(n6876), .C(n6875), .Y(n10444));
NOR3X1   g5794(.A(n9463), .B(g6434), .C(g6428), .Y(n10445));
OR4X1    g5795(.A(n10444), .B(n6884), .C(n10028), .D(n10445), .Y(n10446));
OAI21X1  g5796(.A0(n10445), .A1(n10444), .B0(n10028), .Y(n10447));
NAND2X1  g5797(.A(n10447), .B(n10446), .Y(n10448));
MX2X1    g5798(.A(g6434), .B(n10448), .S0(g35), .Y(n6844));
MX2X1    g5799(.A(g1740), .B(n5624), .S0(n8442), .Y(n10451));
MX2X1    g5800(.A(g1821), .B(n10451), .S0(g35), .Y(n6849));
NAND3X1  g5801(.A(n5606), .B(n4835), .C(g3530), .Y(n10453));
MX2X1    g5802(.A(n5592_1), .B(g3550), .S0(n10453), .Y(n10454));
MX2X1    g5803(.A(g3554), .B(n10454), .S0(g35), .Y(n6854));
INVX1    g5804(.A(g3835), .Y(n10456));
XOR2X1   g5805(.A(g3841), .B(n10456), .Y(n10457));
MX2X1    g5806(.A(g3845), .B(n10457), .S0(n4851_1), .Y(n10458));
MX2X1    g5807(.A(g3841), .B(n10458), .S0(g35), .Y(n6859));
XOR2X1   g5808(.A(n6086), .B(g2116), .Y(n10460));
MX2X1    g5809(.A(g2112), .B(n10460), .S0(g35), .Y(n6864));
NOR2X1   g5810(.A(n7506_1), .B(n4843), .Y(n10462));
MX2X1    g5811(.A(g3195), .B(n5592_1), .S0(n10462), .Y(n10463));
MX2X1    g5812(.A(g3247), .B(n10463), .S0(g35), .Y(n6872));
NOR3X1   g5813(.A(n4850), .B(n4849), .C(g3873), .Y(n10465));
MX2X1    g5814(.A(g3913), .B(n5592_1), .S0(n10465), .Y(n10466));
MX2X1    g5815(.A(g3957), .B(n10466), .S0(g35), .Y(n6877));
INVX1    g5816(.A(g4512), .Y(n10468));
NOR3X1   g5817(.A(g59), .B(g73), .C(g72), .Y(n10469));
MX2X1    g5818(.A(n10468), .B(n10469), .S0(g4581), .Y(n10470));
AND2X1   g5819(.A(n10470), .B(n5702), .Y(n10471));
OAI21X1  g5820(.A0(n9050), .A1(n6849_1), .B0(g35), .Y(n10472));
NAND2X1  g5821(.A(g4492), .B(n4620), .Y(n10473));
OAI21X1  g5822(.A0(n10472), .A1(n10471), .B0(n10473), .Y(n6882));
MX2X1    g5823(.A(g1687), .B(g1682), .S0(n5762), .Y(n10475));
MX2X1    g5824(.A(g1682), .B(n10475), .S0(g35), .Y(n6886));
MX2X1    g5825(.A(g2681), .B(g2675), .S0(n10106), .Y(n10477));
MX2X1    g5826(.A(g2675), .B(n10477), .S0(g35), .Y(n6891));
MX2X1    g5827(.A(g2533), .B(g2527), .S0(n7133), .Y(n10479));
MX2X1    g5828(.A(g2527), .B(n10479), .S0(g35), .Y(n6896));
INVX1    g5829(.A(g305), .Y(n10481));
INVX1    g5830(.A(g324), .Y(n10482));
OAI21X1  g5831(.A0(n10482), .A1(g311), .B0(n10481), .Y(n10483));
MX2X1    g5832(.A(g336), .B(n10483), .S0(g35), .Y(n6901));
MX2X1    g5833(.A(g2697), .B(n4586), .S0(n6435), .Y(n10485));
MX2X1    g5834(.A(g2689), .B(n10485), .S0(g35), .Y(n6906));
NOR3X1   g5835(.A(n7062), .B(n7070_1), .C(n7056), .Y(n10487));
NOR3X1   g5836(.A(n7067), .B(g5742), .C(g5736), .Y(n10488));
OR4X1    g5837(.A(n10487), .B(n7077), .C(n7846), .D(n10488), .Y(n10489));
OAI21X1  g5838(.A0(n10488), .A1(n10487), .B0(n7846), .Y(n10490));
NAND2X1  g5839(.A(n10490), .B(n10489), .Y(n10491));
MX2X1    g5840(.A(g5742), .B(n10491), .S0(g35), .Y(n6911));
MX2X1    g5841(.A(g4382), .B(n5506), .S0(g35), .Y(n6916));
NOR4X1   g5842(.A(g6561), .B(n7204), .C(n7524), .D(n7626), .Y(n10494));
MX2X1    g5843(.A(g6555), .B(n10494), .S0(g35), .Y(n6921));
INVX1    g5844(.A(g1141), .Y(n10496));
OR4X1    g5845(.A(n4707_1), .B(g956), .C(g976), .D(n4708), .Y(n10497));
OAI21X1  g5846(.A0(n4710), .A1(g976), .B0(g956), .Y(n10498));
AOI22X1  g5847(.A0(n10497), .A1(n10498), .B0(n9407), .B1(n10496), .Y(n10499));
MX2X1    g5848(.A(g1141), .B(n10499), .S0(n6189), .Y(n10500));
MX2X1    g5849(.A(g1129), .B(n10500), .S0(g35), .Y(n6926));
MX2X1    g5850(.A(g1554), .B(g496), .S0(g35), .Y(n6931));
MX2X1    g5851(.A(g2413), .B(g2407), .S0(n7941), .Y(n10503));
MX2X1    g5852(.A(g2407), .B(n10503), .S0(g35), .Y(n6935));
INVX1    g5853(.A(g1706), .Y(n10505));
XOR2X1   g5854(.A(g1700), .B(n10505), .Y(n10506));
MX2X1    g5855(.A(g1710), .B(n10506), .S0(n5762), .Y(n10507));
MX2X1    g5856(.A(g1706), .B(n10507), .S0(g35), .Y(n6940));
XOR2X1   g5857(.A(n7724), .B(g6527), .Y(n10509));
MX2X1    g5858(.A(g6523), .B(n10509), .S0(g35), .Y(n6945));
INVX1    g5859(.A(g6497), .Y(n10511));
AOI21X1  g5860(.A0(g6490), .A1(n10511), .B0(g6404), .Y(n10512));
OR2X1    g5861(.A(g6486), .B(n4620), .Y(n10513));
OAI22X1  g5862(.A0(n10512), .A1(n10513), .B0(n10511), .B1(g35), .Y(n6950));
NOR4X1   g5863(.A(g3171), .B(n4844), .C(n5913), .D(n5593), .Y(n10515));
MX2X1    g5864(.A(g3255), .B(n5592_1), .S0(n10515), .Y(n10516));
MX2X1    g5865(.A(g3239), .B(n10516), .S0(g35), .Y(n6955));
INVX1    g5866(.A(g1691), .Y(n10518));
AOI21X1  g5867(.A0(g1648), .A1(n7772), .B0(n10518), .Y(n10519));
XOR2X1   g5868(.A(n10519), .B(g1677), .Y(n10520));
MX2X1    g5869(.A(g1691), .B(n10520), .S0(n8992), .Y(n10521));
MX2X1    g5870(.A(g1677), .B(n10521), .S0(g35), .Y(n6960));
MX2X1    g5871(.A(g2936), .B(n3393), .S0(n5617), .Y(n10523));
MX2X1    g5872(.A(g2922), .B(n10523), .S0(g35), .Y(n6965));
NOR3X1   g5873(.A(n7031), .B(g5644), .C(n7019), .Y(n10525));
AOI21X1  g5874(.A0(n7016), .A1(g5703), .B0(n7026), .Y(n10526));
OAI21X1  g5875(.A0(n10526), .A1(n10525), .B0(n10429), .Y(n10527));
NAND2X1  g5876(.A(g5703), .B(n4620), .Y(n10528));
OAI21X1  g5877(.A0(n10527), .A1(n4620), .B0(n10528), .Y(n6970));
INVX1    g5878(.A(g5142), .Y(n10530));
XOR2X1   g5879(.A(g5148), .B(n10530), .Y(n10531));
MX2X1    g5880(.A(g5152), .B(n10531), .S0(g26801), .Y(n10532));
MX2X1    g5881(.A(g5148), .B(n10532), .S0(g35), .Y(n6975));
NOR2X1   g5882(.A(n6421), .B(n6335), .Y(n10534));
AOI21X1  g5883(.A0(n10534), .A1(g35), .B0(n8859), .Y(n6980));
OR2X1    g5884(.A(g6120), .B(g6116), .Y(n10536));
AOI22X1  g5885(.A0(g6116), .A1(g6120), .B0(n8281), .B1(g6113), .Y(n10537));
OAI21X1  g5886(.A0(n10536), .A1(n10114), .B0(n10537), .Y(n10538));
MX2X1    g5887(.A(g6116), .B(n10538), .S0(g35), .Y(n6988));
OAI21X1  g5888(.A0(n5506), .A1(n9477), .B0(n7180), .Y(n10540));
OAI22X1  g5889(.A0(n7180), .A1(n4803_1), .B0(n5507_1), .B1(n10540), .Y(n10541));
MX2X1    g5890(.A(g2783), .B(n10541), .S0(g35), .Y(n6993));
MX2X1    g5891(.A(g2922), .B(n4447), .S0(n5617), .Y(n10543));
MX2X1    g5892(.A(g2912), .B(n10543), .S0(g35), .Y(n6998));
NOR3X1   g5893(.A(n6188), .B(n6079), .C(g1171), .Y(n10545));
INVX1    g5894(.A(g1111), .Y(n10546));
XOR2X1   g5895(.A(n9405), .B(n5333), .Y(n10547));
AOI21X1  g5896(.A0(n9407), .A1(n10546), .B0(n10547), .Y(n10548));
MX2X1    g5897(.A(g1111), .B(n10548), .S0(n10545), .Y(n10549));
MX2X1    g5898(.A(g1135), .B(n10549), .S0(g35), .Y(n7003));
NAND3X1  g5899(.A(n5632), .B(n4862), .C(g5873), .Y(n10551));
MX2X1    g5900(.A(n5592_1), .B(g5893), .S0(n10551), .Y(n10552));
MX2X1    g5901(.A(g5897), .B(n10552), .S0(g35), .Y(n7008));
NOR2X1   g5902(.A(n5277), .B(g35), .Y(n7013));
NOR4X1   g5903(.A(n4854), .B(g6555), .C(n7524), .D(g6565), .Y(n10555));
MX2X1    g5904(.A(g6617), .B(n5592_1), .S0(n10555), .Y(n10556));
MX2X1    g5905(.A(g6593), .B(n10556), .S0(g35), .Y(n7022));
OAI21X1  g5906(.A0(n6204), .A1(n4926), .B0(n9215), .Y(n10558));
MX2X1    g5907(.A(g2060), .B(n10558), .S0(n9903), .Y(n10559));
MX2X1    g5908(.A(g2066), .B(n10559), .S0(g35), .Y(n7027));
NAND3X1  g5909(.A(n7113_1), .B(n4953), .C(n4950), .Y(n10561));
MX2X1    g5910(.A(g4504), .B(n10561), .S0(g4581), .Y(n10562));
MX2X1    g5911(.A(g4504), .B(n10562), .S0(g35), .Y(n7032));
NOR3X1   g5912(.A(n5916), .B(n5855_1), .C(g5511), .Y(n10564));
MX2X1    g5913(.A(g5599), .B(n5592_1), .S0(n10564), .Y(n10565));
MX2X1    g5914(.A(g5583), .B(n10565), .S0(g35), .Y(n7037));
INVX1    g5915(.A(g3451), .Y(n10567));
AOI21X1  g5916(.A0(g3443), .A1(n10567), .B0(g3401), .Y(n10568));
OR2X1    g5917(.A(g3447), .B(n4620), .Y(n10569));
OAI22X1  g5918(.A0(n10568), .A1(n10569), .B0(n10567), .B1(g35), .Y(n7042));
NOR4X1   g5919(.A(n6621), .B(g4639), .C(n5848), .D(n6019), .Y(n10571));
AOI21X1  g5920(.A0(n10571), .A1(n5724), .B0(n4620), .Y(n7047));
MX2X1    g5921(.A(g94), .B(n6708), .S0(n9636), .Y(n10573));
MX2X1    g5922(.A(g37), .B(n10573), .S0(g35), .Y(n7055));
INVX1    g5923(.A(g3119), .Y(n10575));
XOR2X1   g5924(.A(g3125), .B(n10575), .Y(n10576));
MX2X1    g5925(.A(g3129), .B(n10576), .S0(n8618), .Y(n10577));
MX2X1    g5926(.A(g3125), .B(n10577), .S0(g35), .Y(n7060));
NAND2X1  g5927(.A(n6624), .B(g5164), .Y(n10579));
NAND2X1  g5928(.A(g5170), .B(n5610), .Y(n10580));
AOI21X1  g5929(.A0(n10580), .A1(n10579), .B0(n6042), .Y(n10581));
MX2X1    g5930(.A(g5164), .B(n10581), .S0(g35), .Y(n7070));
NOR2X1   g5931(.A(n8564), .B(g35), .Y(n7075));
XOR2X1   g5932(.A(n4863), .B(g5821), .Y(n10584));
MX2X1    g5933(.A(g5817), .B(n10584), .S0(g35), .Y(n7080));
NOR4X1   g5934(.A(g6227), .B(n5980), .C(n4871_1), .D(n6208), .Y(n10586));
MX2X1    g5935(.A(g6299), .B(n5592_1), .S0(n10586), .Y(n10587));
MX2X1    g5936(.A(g6283), .B(n10587), .S0(g35), .Y(n7085));
NAND3X1  g5937(.A(n9925), .B(n9924), .C(g3727), .Y(n10589));
OAI21X1  g5938(.A0(n7360), .A1(n7355), .B0(n7358), .Y(n10590));
OAI21X1  g5939(.A0(n10589), .A1(n7371), .B0(n10590), .Y(n10591));
MX2X1    g5940(.A(g3723), .B(n10591), .S0(g35), .Y(n7093));
NAND3X1  g5941(.A(n4943), .B(n7088), .C(g2016), .Y(n10593));
NAND3X1  g5942(.A(g2004), .B(g2051), .C(n7088), .Y(n10594));
AND2X1   g5943(.A(n10594), .B(n10593), .Y(n10595));
AND2X1   g5944(.A(g2060), .B(g2028), .Y(n10596));
AOI22X1  g5945(.A0(n10596), .A1(g2008), .B0(g2012), .B1(n9980), .Y(n10597));
NAND3X1  g5946(.A(n4943), .B(g2051), .C(g2024), .Y(n10598));
NAND3X1  g5947(.A(n9215), .B(g2028), .C(g2020), .Y(n10599));
NAND4X1  g5948(.A(n10598), .B(n10597), .C(n10595), .D(n10599), .Y(n10600));
MX2X1    g5949(.A(g2079), .B(n10600), .S0(n9903), .Y(n10601));
MX2X1    g5950(.A(g2060), .B(n10601), .S0(g35), .Y(n7098));
AOI21X1  g5951(.A0(n4970), .A1(n4820), .B0(n6721), .Y(n10603));
MX2X1    g5952(.A(g4704), .B(g101), .S0(n6721), .Y(n10604));
MX2X1    g5953(.A(n10604), .B(g4698), .S0(n10603), .Y(n10605));
MX2X1    g5954(.A(g4704), .B(n10605), .S0(g35), .Y(n7103));
NAND3X1  g5955(.A(n8051), .B(n5930), .C(n5937), .Y(n10607));
OAI21X1  g5956(.A0(n5930), .A1(n5937), .B0(n10607), .Y(n10608));
MX2X1    g5957(.A(g3698), .B(n10608), .S0(g35), .Y(n7108));
NAND3X1  g5958(.A(n7520_1), .B(n10265), .C(g1564), .Y(n10610));
OAI21X1  g5959(.A0(n7669), .A1(n7667), .B0(g1559), .Y(n10611));
AOI21X1  g5960(.A0(n10611), .A1(n10610), .B0(n7670), .Y(n10612));
MX2X1    g5961(.A(g1564), .B(n10612), .S0(g35), .Y(n7113));
NOR2X1   g5962(.A(n9437), .B(n6316_1), .Y(n10614));
OAI21X1  g5963(.A0(n4710), .A1(g943), .B0(g35), .Y(n10615));
OAI22X1  g5964(.A0(n10614), .A1(n10615), .B0(n5453), .B1(g35), .Y(n7118));
MX2X1    g5965(.A(n8737), .B(g411), .S0(n6235), .Y(n10618));
MX2X1    g5966(.A(g417), .B(n10618), .S0(g35), .Y(n7123));
AND2X1   g5967(.A(g6227), .B(g35), .Y(n7128));
NOR4X1   g5968(.A(n7041), .B(g3881), .C(n4848), .D(n7642), .Y(n10621));
MX2X1    g5969(.A(g3953), .B(n5592_1), .S0(n10621), .Y(n10622));
MX2X1    g5970(.A(g3937), .B(n10622), .S0(g35), .Y(n7132));
NOR2X1   g5971(.A(g3061), .B(n9099), .Y(n10624));
MX2X1    g5972(.A(n10624), .B(n9100), .S0(g3072), .Y(n10625));
MX2X1    g5973(.A(g3065), .B(n10625), .S0(g35), .Y(n7137));
MX2X1    g5974(.A(g2704), .B(n3220), .S0(n6435), .Y(n10627));
MX2X1    g5975(.A(g2697), .B(n10627), .S0(g35), .Y(n7142));
XOR2X1   g5976(.A(n5749), .B(g6035), .Y(n10629));
MX2X1    g5977(.A(g6031), .B(n10629), .S0(g35), .Y(n7147));
AND2X1   g5978(.A(n6182), .B(n6180), .Y(n10631));
NOR2X1   g5979(.A(n5820), .B(n5812), .Y(n10632));
MX2X1    g5980(.A(n5812), .B(n10632), .S0(n10631), .Y(n10633));
MX2X1    g5981(.A(g6077), .B(n10633), .S0(g35), .Y(n7152));
AOI21X1  g5982(.A0(n5399), .A1(n5380_1), .B0(g22), .Y(n10635));
AOI21X1  g5983(.A0(n5399), .A1(n5380_1), .B0(n5282), .Y(n10636));
OR2X1    g5984(.A(n10636), .B(n10635), .Y(n7157));
NOR4X1   g5985(.A(g1514), .B(g1526), .C(n6513), .D(n7603), .Y(n10638));
XOR2X1   g5986(.A(g1300), .B(g1484), .Y(n10639));
MX2X1    g5987(.A(g1300), .B(n10639), .S0(n10638), .Y(n10640));
MX2X1    g5988(.A(g1484), .B(n10640), .S0(g35), .Y(n7162));
XOR2X1   g5989(.A(g4057), .B(n4729), .Y(n10642));
OAI22X1  g5990(.A0(n7630), .A1(n10642), .B0(n4729), .B1(g35), .Y(n7167));
NAND3X1  g5991(.A(n7561), .B(n4643), .C(g5180), .Y(n10644));
MX2X1    g5992(.A(n5592_1), .B(g5200), .S0(n10644), .Y(n10645));
MX2X1    g5993(.A(g5204), .B(n10645), .S0(g35), .Y(n7172));
NOR2X1   g5994(.A(n9600), .B(g4878), .Y(n10647));
NOR2X1   g5995(.A(g4843), .B(n4959_1), .Y(n10648));
OAI21X1  g5996(.A0(n10648), .A1(n10647), .B0(n9595), .Y(n10649));
NAND2X1  g5997(.A(g4878), .B(n4620), .Y(n10650));
OAI21X1  g5998(.A0(n10649), .A1(n4620), .B0(n10650), .Y(n7177));
AND2X1   g5999(.A(n5490), .B(n5484), .Y(n10652));
NOR2X1   g6000(.A(n5501), .B(n5478), .Y(n10653));
MX2X1    g6001(.A(n5478), .B(n10653), .S0(n10652), .Y(n10654));
MX2X1    g6002(.A(g5041), .B(n10654), .S0(g35), .Y(n7182));
INVX1    g6003(.A(g2250), .Y(n10656));
AOI21X1  g6004(.A0(n5789), .A1(g2208), .B0(n10656), .Y(n10657));
XOR2X1   g6005(.A(n10657), .B(g2236), .Y(n10658));
MX2X1    g6006(.A(g2250), .B(n10658), .S0(n5788), .Y(n10659));
MX2X1    g6007(.A(g2236), .B(n10659), .S0(g35), .Y(n7187));
OR2X1    g6008(.A(g305), .B(g311), .Y(n10661));
MX2X1    g6009(.A(g316), .B(n10661), .S0(g35), .Y(n7192));
NAND3X1  g6010(.A(n5920), .B(n4953), .C(g72), .Y(n10663));
MX2X1    g6011(.A(g4546), .B(n10663), .S0(g4581), .Y(n10664));
MX2X1    g6012(.A(g4546), .B(n10664), .S0(g35), .Y(n7197));
OAI21X1  g6013(.A0(g2453), .A1(n6445), .B0(n4929), .Y(n10666));
OAI21X1  g6014(.A0(n6204), .A1(n4917), .B0(n10666), .Y(n10667));
MX2X1    g6015(.A(g2453), .B(n10667), .S0(n6444_1), .Y(n10668));
MX2X1    g6016(.A(g2461), .B(n10668), .S0(g35), .Y(n7202));
MX2X1    g6017(.A(g5841), .B(g5835), .S0(n4863), .Y(n10670));
MX2X1    g6018(.A(g5835), .B(n10670), .S0(g35), .Y(n7207));
MX2X1    g6019(.A(g5759), .B(n7073), .S0(g35), .Y(n7212));
NOR3X1   g6020(.A(n7356), .B(n7364), .C(n7350), .Y(n10673));
NOR3X1   g6021(.A(n7361), .B(g3742), .C(g3736), .Y(n10674));
OR4X1    g6022(.A(n10673), .B(n7371), .C(n8121), .D(n10674), .Y(n10675));
OAI21X1  g6023(.A0(n10674), .A1(n10673), .B0(n8121), .Y(n10676));
NAND2X1  g6024(.A(n10676), .B(n10675), .Y(n10677));
MX2X1    g6025(.A(g3742), .B(n10677), .S0(g35), .Y(n7217));
MX2X1    g6026(.A(g2912), .B(n6676), .S0(n5617), .Y(n10679));
MX2X1    g6027(.A(g2907), .B(n10679), .S0(g35), .Y(n7225));
NAND4X1  g6028(.A(n5506), .B(n4913), .C(g2741), .D(n7227), .Y(n10681));
XOR2X1   g6029(.A(n7616), .B(g110), .Y(n10682));
MX2X1    g6030(.A(n10682), .B(g2357), .S0(n10681), .Y(n10683));
MX2X1    g6031(.A(g2342), .B(n10683), .S0(g35), .Y(n7230));
NOR3X1   g6032(.A(n7302_1), .B(n5661), .C(n7297), .Y(n10685));
MX2X1    g6033(.A(n7297), .B(n10685), .S0(n7305), .Y(n10686));
MX2X1    g6034(.A(g146), .B(n10686), .S0(g35), .Y(n7238));
MX2X1    g6035(.A(g4253), .B(n6708), .S0(n9562), .Y(n10688));
MX2X1    g6036(.A(g4300), .B(n10688), .S0(g35), .Y(n7243));
OAI21X1  g6037(.A0(g5062), .A1(g5022), .B0(n5482_1), .Y(n10690));
NAND3X1  g6038(.A(g5016), .B(n5480), .C(n5488), .Y(n10691));
OAI21X1  g6039(.A0(n10690), .A1(n5501), .B0(n10691), .Y(n10692));
MX2X1    g6040(.A(g5022), .B(n10692), .S0(g35), .Y(n7248));
XOR2X1   g6041(.A(n4846_1), .B(g3119), .Y(n10694));
MX2X1    g6042(.A(g3115), .B(n10694), .S0(g35), .Y(n7253));
NAND2X1  g6043(.A(g1361), .B(g1373), .Y(n10696));
NAND4X1  g6044(.A(n5984), .B(g1351), .C(n7283_1), .D(n10696), .Y(n10697));
NAND2X1  g6045(.A(n10696), .B(g1351), .Y(n10698));
MX2X1    g6046(.A(n10698), .B(n9765), .S0(n5984), .Y(n10699));
NAND2X1  g6047(.A(n10699), .B(n10697), .Y(n10700));
MX2X1    g6048(.A(g1351), .B(n10700), .S0(n5986), .Y(n10701));
MX2X1    g6049(.A(g1312), .B(n10701), .S0(g35), .Y(n7258));
OAI21X1  g6050(.A0(n6204), .A1(n4922), .B0(n7772), .Y(n10703));
MX2X1    g6051(.A(g1648), .B(n10703), .S0(n8992), .Y(n10704));
MX2X1    g6052(.A(g1624), .B(n10704), .S0(g35), .Y(n7263));
NAND2X1  g6053(.A(g4515), .B(n4620), .Y(n10706));
OAI21X1  g6054(.A0(n10470), .A1(n4620), .B0(n10706), .Y(n7268));
AND2X1   g6055(.A(n6439_1), .B(g5115), .Y(n10708));
XOR2X1   g6056(.A(n10708), .B(n6377), .Y(n10709));
MX2X1    g6057(.A(g5115), .B(n10709), .S0(g28753), .Y(n10710));
MX2X1    g6058(.A(g5120), .B(n10710), .S0(g35), .Y(n7273));
NAND3X1  g6059(.A(n7758), .B(n7756), .C(n7759), .Y(n10712));
OAI21X1  g6060(.A0(n7756), .A1(n7759), .B0(n10712), .Y(n10713));
MX2X1    g6061(.A(g3347), .B(n10713), .S0(g35), .Y(n7278));
MX2X1    g6062(.A(g6657), .B(n5592_1), .S0(n4857), .Y(n10716));
MX2X1    g6063(.A(g6653), .B(n10716), .S0(g35), .Y(n7283));
NAND3X1  g6064(.A(n6835_1), .B(n4953), .C(n4950), .Y(n10718));
MX2X1    g6065(.A(g4549), .B(n10718), .S0(g4581), .Y(n10719));
MX2X1    g6066(.A(g4549), .B(n10719), .S0(g35), .Y(n7288));
NAND3X1  g6067(.A(n6152), .B(n4850), .C(g3873), .Y(n10721));
MX2X1    g6068(.A(n5592_1), .B(g3893), .S0(n10721), .Y(n10722));
MX2X1    g6069(.A(g3897), .B(n10722), .S0(g35), .Y(n7293));
NOR3X1   g6070(.A(g3171), .B(n4844), .C(n4843), .Y(n10724));
MX2X1    g6071(.A(g3211), .B(n5592_1), .S0(n10724), .Y(n10725));
MX2X1    g6072(.A(g3255), .B(n10725), .S0(g35), .Y(n7298));
AND2X1   g6073(.A(g1311), .B(n4620), .Y(n7306));
NOR4X1   g6074(.A(g5527), .B(n4867), .C(g5511), .D(n5855_1), .Y(n10728));
MX2X1    g6075(.A(g5595), .B(n5592_1), .S0(n10728), .Y(n10729));
MX2X1    g6076(.A(g5579), .B(n10729), .S0(g35), .Y(n7314));
MX2X1    g6077(.A(g3614), .B(n5592_1), .S0(n4836_1), .Y(n10732));
MX2X1    g6078(.A(g3610), .B(n10732), .S0(g35), .Y(n7319));
MX2X1    g6079(.A(g2894), .B(n3393), .S0(n5697), .Y(n10734));
MX2X1    g6080(.A(g2860), .B(n10734), .S0(g35), .Y(n7324));
MX2X1    g6081(.A(g3125), .B(g3119), .S0(n8618), .Y(n10736));
MX2X1    g6082(.A(g3119), .B(n10736), .S0(g35), .Y(n7329));
XOR2X1   g6083(.A(n4851_1), .B(g3821), .Y(n10738));
MX2X1    g6084(.A(g3817), .B(n10738), .S0(g35), .Y(n7337));
INVX1    g6085(.A(g4141), .Y(n10740));
XOR2X1   g6086(.A(n7337_1), .B(n10740), .Y(n10741));
OAI22X1  g6087(.A0(n7630), .A1(n10741), .B0(n4731_1), .B1(g35), .Y(n7342));
NAND2X1  g6088(.A(g4552), .B(n4620), .Y(n10743));
OAI21X1  g6089(.A0(n6844_1), .A1(n4620), .B0(n10743), .Y(n7347));
NOR2X1   g6090(.A(n7933), .B(n4644), .Y(n10745));
MX2X1    g6091(.A(g5272), .B(n5592_1), .S0(n10745), .Y(n10746));
MX2X1    g6092(.A(g5268), .B(n10746), .S0(g35), .Y(n7352));
XOR2X1   g6093(.A(n7692), .B(g2735), .Y(n10748));
NAND2X1  g6094(.A(n10748), .B(g2841), .Y(n10749));
MX2X1    g6095(.A(g2729), .B(n10749), .S0(g35), .Y(n7357));
MX2X1    g6096(.A(g661), .B(g728), .S0(n6389_1), .Y(n10751));
MX2X1    g6097(.A(g661), .B(n10751), .S0(g35), .Y(n7362));
NOR3X1   g6098(.A(n7379), .B(n6208), .C(n5980), .Y(n10753));
MX2X1    g6099(.A(g6295), .B(n5592_1), .S0(n10753), .Y(n10754));
MX2X1    g6100(.A(g6279), .B(n10754), .S0(g35), .Y(n7367));
MX2X1    g6101(.A(g5413), .B(n6642), .S0(g35), .Y(n7372));
XOR2X1   g6102(.A(n10106), .B(g2661), .Y(n10757));
MX2X1    g6103(.A(g2657), .B(n10757), .S0(g35), .Y(n7377));
MX2X1    g6104(.A(g1988), .B(g1982), .S0(n5841_1), .Y(n10759));
MX2X1    g6105(.A(g1982), .B(n10759), .S0(g35), .Y(n7382));
XOR2X1   g6106(.A(g26801), .B(g5128), .Y(n10761));
MX2X1    g6107(.A(g5124), .B(n10761), .S0(g35), .Y(n7387));
XOR2X1   g6108(.A(g1548), .B(g1430), .Y(n10763));
MX2X1    g6109(.A(g1430), .B(n10763), .S0(g35), .Y(n7392));
AND2X1   g6110(.A(n8617), .B(g3106), .Y(n10765));
XOR2X1   g6111(.A(n10765), .B(n8662), .Y(n10766));
MX2X1    g6112(.A(g3106), .B(n10766), .S0(n7756), .Y(n10767));
MX2X1    g6113(.A(g3111), .B(n10767), .S0(g35), .Y(n7397));
AND2X1   g6114(.A(n7824), .B(n7826), .Y(n10769));
NOR2X1   g6115(.A(n7824), .B(n7826), .Y(n10770));
OAI21X1  g6116(.A0(n10770), .A1(n10769), .B0(n7822), .Y(n10771));
NAND2X1  g6117(.A(g4653), .B(n4620), .Y(n10772));
OAI21X1  g6118(.A0(n10771), .A1(n4620), .B0(n10772), .Y(n7402));
NAND3X1  g6119(.A(n10210), .B(n5181_1), .C(g4349), .Y(n10774));
OAI21X1  g6120(.A0(n10212), .A1(n5174), .B0(g4358), .Y(n10775));
AOI21X1  g6121(.A0(n10775), .A1(n10774), .B0(n7341), .Y(n10776));
MX2X1    g6122(.A(g4349), .B(n10776), .S0(g35), .Y(n7407));
OAI21X1  g6123(.A0(n6204), .A1(n4925_1), .B0(n8135), .Y(n10778));
MX2X1    g6124(.A(g1792), .B(n10778), .S0(n8134), .Y(n10779));
MX2X1    g6125(.A(g1798), .B(n10779), .S0(g35), .Y(n7412));
NOR2X1   g6126(.A(n6082), .B(n5524), .Y(n10781));
MX2X1    g6127(.A(n10781), .B(g1246), .S0(n6084), .Y(n10782));
OAI21X1  g6128(.A0(g1996), .A1(g2070), .B0(g2084), .Y(n10783));
XOR2X1   g6129(.A(n10783), .B(n10782), .Y(n10784));
MX2X1    g6130(.A(g2084), .B(n10784), .S0(n8497), .Y(n10785));
MX2X1    g6131(.A(g2070), .B(n10785), .S0(g35), .Y(n7417));
MX2X1    g6132(.A(g3057), .B(n5580), .S0(g35), .Y(n7422));
NOR4X1   g6133(.A(g3161), .B(g3167), .C(g3155), .D(n7506_1), .Y(n10788));
MX2X1    g6134(.A(g3187), .B(n5592_1), .S0(n10788), .Y(n10789));
MX2X1    g6135(.A(g3179), .B(n10789), .S0(g35), .Y(n7427));
NAND4X1  g6136(.A(n7471), .B(n5845_1), .C(g4311), .D(n6021), .Y(n10791));
NAND4X1  g6137(.A(n6020_1), .B(n5845_1), .C(n4949_1), .D(n6021), .Y(n10792));
AOI21X1  g6138(.A0(n10792), .A1(n10791), .B0(n4620), .Y(n7432));
NOR3X1   g6139(.A(n6003), .B(n5156), .C(g2599), .Y(n10794));
MX2X1    g6140(.A(g2583), .B(n5998), .S0(n10794), .Y(n10795));
MX2X1    g6141(.A(g2571), .B(n10795), .S0(g35), .Y(n7437));
NOR2X1   g6142(.A(n4782), .B(g35), .Y(n7442));
NOR3X1   g6143(.A(n6188), .B(g1183), .C(n4665), .Y(n10798));
INVX1    g6144(.A(g1094), .Y(n10799));
OR4X1    g6145(.A(n4707_1), .B(g1135), .C(g976), .D(n4708), .Y(n10800));
OAI21X1  g6146(.A0(n4710), .A1(g976), .B0(g1135), .Y(n10801));
AOI22X1  g6147(.A0(n10800), .A1(n10801), .B0(n9407), .B1(n10799), .Y(n10802));
MX2X1    g6148(.A(g1094), .B(n10802), .S0(n10798), .Y(n10803));
MX2X1    g6149(.A(g1099), .B(n10803), .S0(g35), .Y(n7447));
MX2X1    g6150(.A(g3841), .B(g3835), .S0(n4851_1), .Y(n10805));
MX2X1    g6151(.A(g3835), .B(n10805), .S0(g35), .Y(n7452));
XOR2X1   g6152(.A(g4277), .B(g4281), .Y(n10807));
MX2X1    g6153(.A(g4281), .B(n10807), .S0(g35), .Y(n7457));
MX2X1    g6154(.A(g3759), .B(n7367_1), .S0(g35), .Y(n7462));
NAND3X1  g6155(.A(n10275), .B(g3171), .C(n4844), .Y(n10810));
MX2X1    g6156(.A(n5592_1), .B(g3191), .S0(n10810), .Y(n10811));
MX2X1    g6157(.A(g3195), .B(n10811), .S0(g35), .Y(n7467));
MX2X1    g6158(.A(g4273), .B(n8821), .S0(g35), .Y(n7472));
MX2X1    g6159(.A(n8246), .B(n8247), .S0(n5769), .Y(n10814));
NOR2X1   g6160(.A(n5778_1), .B(n5770), .Y(n10815));
MX2X1    g6161(.A(n5770), .B(n10815), .S0(n10814), .Y(n10816));
MX2X1    g6162(.A(g3385), .B(n10816), .S0(g35), .Y(n7477));
NAND3X1  g6163(.A(g691), .B(n9706), .C(g703), .Y(n10818));
OAI21X1  g6164(.A0(n9338), .A1(g691), .B0(n10818), .Y(n10819));
MX2X1    g6165(.A(g691), .B(n10819), .S0(n5880_1), .Y(n10820));
MX2X1    g6166(.A(g79), .B(n10820), .S0(g35), .Y(n7486));
NOR3X1   g6167(.A(n5462), .B(n5226_1), .C(n5616), .Y(n10822));
OAI21X1  g6168(.A0(g534), .A1(g301), .B0(g35), .Y(n10823));
OAI22X1  g6169(.A0(n10822), .A1(n10823), .B0(n5351), .B1(g35), .Y(n7491));
INVX1    g6170(.A(g5459), .Y(n10825));
AOI21X1  g6171(.A0(n10825), .A1(g5452), .B0(g5366), .Y(n10826));
OR2X1    g6172(.A(g5448), .B(n4620), .Y(n10827));
OAI22X1  g6173(.A0(n10826), .A1(n10827), .B0(n10825), .B1(g35), .Y(n7496));
XOR2X1   g6174(.A(n6245), .B(g385), .Y(n10829));
MX2X1    g6175(.A(g376), .B(n10829), .S0(g35), .Y(n7501));
NOR3X1   g6176(.A(n6085), .B(n7842), .C(g2040), .Y(n10831));
MX2X1    g6177(.A(g2004), .B(n7037_1), .S0(n10831), .Y(n10832));
MX2X1    g6178(.A(g2008), .B(n10832), .S0(g35), .Y(n7506));
XOR2X1   g6179(.A(n5570), .B(g2527), .Y(n10834));
MX2X1    g6180(.A(g2523), .B(n10834), .S0(g35), .Y(n7511));
XOR2X1   g6181(.A(g4537), .B(g4534), .Y(n10836));
MX2X1    g6182(.A(g4534), .B(n10836), .S0(g35), .Y(n7520));
MX2X1    g6183(.A(g5148), .B(g5142), .S0(g26801), .Y(n10838));
MX2X1    g6184(.A(g5142), .B(n10838), .S0(g35), .Y(n7525));
INVX1    g6185(.A(g4459), .Y(n10840));
NAND2X1  g6186(.A(g4473), .B(n10840), .Y(n10841));
MX2X1    g6187(.A(g113), .B(g4507), .S0(n10841), .Y(n10842));
OR2X1    g6188(.A(g70), .B(n4620), .Y(n10843));
MX2X1    g6189(.A(n10842), .B(n10843), .S0(n4620), .Y(n7530));
NAND2X1  g6190(.A(n8861), .B(g35), .Y(n10845));
OAI22X1  g6191(.A0(n10534), .A1(n10845), .B0(n6335), .B1(g35), .Y(n7535));
NOR4X1   g6192(.A(g3171), .B(n4844), .C(n5913), .D(g3161), .Y(n10847));
MX2X1    g6193(.A(g3223), .B(n5592_1), .S0(n10847), .Y(n10848));
MX2X1    g6194(.A(g3199), .B(n10848), .S0(g35), .Y(n7540));
NOR2X1   g6195(.A(n6807), .B(g35), .Y(n7545));
MX2X1    g6196(.A(g2970), .B(n4586), .S0(n5617), .Y(n10851));
MX2X1    g6197(.A(g2960), .B(n10851), .S0(g35), .Y(n7550));
AOI21X1  g6198(.A0(n10172), .A1(g35), .B0(n7018), .Y(n7555));
INVX1    g6199(.A(g3408), .Y(n10854));
AOI21X1  g6200(.A0(n10854), .A1(g35), .B0(n9008), .Y(n7560));
NOR4X1   g6201(.A(g5188), .B(n5610), .C(n4642_1), .D(n6624), .Y(n10856));
MX2X1    g6202(.A(g5260), .B(n5592_1), .S0(n10856), .Y(n10857));
MX2X1    g6203(.A(g5244), .B(n10857), .S0(g35), .Y(n7565));
MX2X1    g6204(.A(g1521), .B(g1339), .S0(g1500), .Y(n10859));
MX2X1    g6205(.A(g1526), .B(n10859), .S0(g35), .Y(n7570));
NAND2X1  g6206(.A(n4835), .B(g3518), .Y(n10861));
NAND2X1  g6207(.A(g3522), .B(n4834), .Y(n10862));
AOI21X1  g6208(.A0(n10862), .A1(n10861), .B0(n5732), .Y(n10863));
MX2X1    g6209(.A(g3518), .B(n10863), .S0(g35), .Y(n7575));
XOR2X1   g6210(.A(g3106), .B(g3111), .Y(n10865));
MX2X1    g6211(.A(g3115), .B(n10865), .S0(n8618), .Y(n10866));
MX2X1    g6212(.A(g3106), .B(n10866), .S0(g35), .Y(n7580));
NOR4X1   g6213(.A(n4845), .B(g3179), .C(n5913), .D(n5593), .Y(n10868));
MX2X1    g6214(.A(g3251), .B(n5592_1), .S0(n10868), .Y(n10869));
MX2X1    g6215(.A(g3235), .B(n10869), .S0(g35), .Y(n7585));
MX2X1    g6216(.A(g4455), .B(n9584), .S0(g35), .Y(n7590));
NOR3X1   g6217(.A(g4628), .B(n5850_1), .C(n5848), .Y(n10872));
AOI21X1  g6218(.A0(g4639), .A1(g4621), .B0(n6018), .Y(n10873));
OAI21X1  g6219(.A0(n10873), .A1(n10872), .B0(n5846), .Y(n10874));
NAND2X1  g6220(.A(g4621), .B(n4620), .Y(n10875));
OAI21X1  g6221(.A0(n10874), .A1(n4620), .B0(n10875), .Y(n7595));
NAND3X1  g6222(.A(n6084), .B(n6081), .C(g1996), .Y(n10877));
AOI21X1  g6223(.A0(n7842), .A1(g2040), .B0(g2070), .Y(n10878));
NAND3X1  g6224(.A(n10878), .B(n8498), .C(n8497), .Y(n10879));
AOI21X1  g6225(.A0(n10879), .A1(n10877), .B0(n4620), .Y(n7600));
MX2X1    g6226(.A(g3401), .B(g3689), .S0(g35), .Y(n7605));
MX2X1    g6227(.A(n9051), .B(g4515), .S0(g4521), .Y(n10882));
MX2X1    g6228(.A(g4527), .B(n10882), .S0(g35), .Y(n7609));
NOR4X1   g6229(.A(n5004), .B(n4988_1), .C(n5616), .D(n5462), .Y(n10884));
OAI21X1  g6230(.A0(g4300), .A1(g4242), .B0(g35), .Y(n10885));
NAND2X1  g6231(.A(g4297), .B(n4620), .Y(n10886));
OAI21X1  g6232(.A0(n10885), .A1(n10884), .B0(n10886), .Y(n7617));
INVX1    g6233(.A(g1714), .Y(n10888));
XOR2X1   g6234(.A(g1720), .B(n10888), .Y(n10889));
MX2X1    g6235(.A(g1724), .B(n10889), .S0(n7773), .Y(n10890));
MX2X1    g6236(.A(g1720), .B(n10890), .S0(g35), .Y(n7622));
NOR4X1   g6237(.A(n7289), .B(n7288_1), .C(n7287), .D(n8213), .Y(n10892));
NOR2X1   g6238(.A(n7286), .B(g1379), .Y(n10893));
MX2X1    g6239(.A(g1379), .B(n10893), .S0(n10892), .Y(n10894));
MX2X1    g6240(.A(g1373), .B(n10894), .S0(g35), .Y(n7627));
OAI22X1  g6241(.A0(g3661), .A1(n5803), .B0(n5804), .B1(g3654), .Y(n10896));
MX2X1    g6242(.A(g3649), .B(n5803), .S0(g3625), .Y(n10897));
INVX1    g6243(.A(g3661), .Y(n10898));
OAI21X1  g6244(.A0(n10898), .A1(g3632), .B0(g35), .Y(n10899));
NOR4X1   g6245(.A(n10897), .B(n10896), .C(n8476), .D(n10899), .Y(n7632));
INVX1    g6246(.A(g56), .Y(n10901));
NAND4X1  g6247(.A(g58), .B(n4976), .C(n10901), .D(n5616), .Y(n10902));
NOR4X1   g6248(.A(n4977), .B(n4976), .C(g57), .D(n10902), .Y(n7636));
NOR3X1   g6249(.A(n5531_1), .B(n8892), .C(g1936), .Y(n10904));
MX2X1    g6250(.A(g1878), .B(n5526_1), .S0(n10904), .Y(n10905));
MX2X1    g6251(.A(g1870), .B(n10905), .S0(g35), .Y(n7641));
MX2X1    g6252(.A(g5619), .B(n5592_1), .S0(n4869), .Y(n10908));
MX2X1    g6253(.A(g5615), .B(n10908), .S0(g35), .Y(n7646));
NOR2X1   g6254(.A(n4900), .B(n4889), .Y(n10910));
NOR3X1   g6255(.A(n4900), .B(n4888), .C(n4809), .Y(n10911));
OR2X1    g6256(.A(n10911), .B(n10910), .Y(n7651));
BUFX1    g6257(.A(g4408), .Y(g7243));
BUFX1    g6258(.A(g4446), .Y(g7245));
BUFX1    g6259(.A(g4414), .Y(g7257));
BUFX1    g6260(.A(g4449), .Y(g7260));
BUFX1    g6261(.A(g344), .Y(g7540));
BUFX1    g6262(.A(g1157), .Y(g7916));
BUFX1    g6263(.A(g1500), .Y(g7946));
BUFX1    g6264(.A(g4809), .Y(g8132));
BUFX1    g6265(.A(g4999), .Y(g8178));
BUFX1    g6266(.A(g3092), .Y(g8215));
BUFX1    g6267(.A(g4812), .Y(g8235));
BUFX1    g6268(.A(g3096), .Y(g8277));
BUFX1    g6269(.A(g3443), .Y(g8279));
BUFX1    g6270(.A(g5002), .Y(g8283));
BUFX1    g6271(.A(g215), .Y(g8291));
BUFX1    g6272(.A(g3447), .Y(g8342));
BUFX1    g6273(.A(g3794), .Y(g8344));
BUFX1    g6274(.A(g4815), .Y(g8353));
BUFX1    g6275(.A(g194), .Y(g8358));
BUFX1    g6276(.A(g3798), .Y(g8398));
BUFX1    g6277(.A(g5005), .Y(g8403));
BUFX1    g6278(.A(g1239), .Y(g8416));
BUFX1    g6279(.A(g1582), .Y(g8475));
BUFX1    g6280(.A(g365), .Y(g8719));
BUFX1    g6281(.A(g4188), .Y(g8783));
BUFX1    g6282(.A(g4194), .Y(g8784));
BUFX1    g6283(.A(g4197), .Y(g8785));
BUFX1    g6284(.A(g4200), .Y(g8786));
BUFX1    g6285(.A(g4204), .Y(g8787));
BUFX1    g6286(.A(g4207), .Y(g8788));
BUFX1    g6287(.A(g4210), .Y(g8789));
BUFX1    g6288(.A(g4277), .Y(g8839));
BUFX1    g6289(.A(g4222), .Y(g8870));
BUFX1    g6290(.A(g4213), .Y(g8915));
BUFX1    g6291(.A(g4216), .Y(g8916));
BUFX1    g6292(.A(g4219), .Y(g8917));
BUFX1    g6293(.A(g4226), .Y(g8918));
BUFX1    g6294(.A(g4229), .Y(g8919));
BUFX1    g6295(.A(g4232), .Y(g8920));
BUFX1    g6296(.A(g4287), .Y(g9019));
BUFX1    g6297(.A(g640), .Y(g9048));
BUFX1    g6298(.A(g4304), .Y(g9251));
BUFX1    g6299(.A(g5101), .Y(g9497));
BUFX1    g6300(.A(g5105), .Y(g9553));
BUFX1    g6301(.A(g5448), .Y(g9555));
BUFX1    g6302(.A(g5452), .Y(g9615));
BUFX1    g6303(.A(g5794), .Y(g9617));
BUFX1    g6304(.A(g5798), .Y(g9680));
BUFX1    g6305(.A(g6140), .Y(g9682));
BUFX1    g6306(.A(g6144), .Y(g9741));
BUFX1    g6307(.A(g6486), .Y(g9743));
BUFX1    g6308(.A(g6490), .Y(g9817));
BUFX1    g6309(.A(g4294), .Y(g10122));
BUFX1    g6310(.A(g4537), .Y(g10306));
BUFX1    g6311(.A(g1233), .Y(g10500));
BUFX1    g6312(.A(g1576), .Y(g10527));
BUFX1    g6313(.A(g3303), .Y(g11349));
BUFX1    g6314(.A(g3654), .Y(g11388));
BUFX1    g6315(.A(g4005), .Y(g11418));
BUFX1    g6316(.A(g4191), .Y(g11447));
BUFX1    g6317(.A(g802), .Y(g11678));
BUFX1    g6318(.A(g4185), .Y(g11770));
BUFX1    g6319(.A(g799), .Y(g12184));
BUFX1    g6320(.A(g5313), .Y(g12238));
BUFX1    g6321(.A(g5659), .Y(g12300));
BUFX1    g6322(.A(g6005), .Y(g12350));
BUFX1    g6323(.A(g637), .Y(g12368));
BUFX1    g6324(.A(g6351), .Y(g12422));
BUFX1    g6325(.A(g6697), .Y(g12470));
BUFX1    g6326(.A(g1), .Y(g12832));
BUFX1    g6327(.A(g1227), .Y(g12919));
BUFX1    g6328(.A(g1570), .Y(g12923));
BUFX1    g6329(.A(g5308), .Y(g13039));
BUFX1    g6330(.A(g5654), .Y(g13049));
BUFX1    g6331(.A(g6000), .Y(g13068));
BUFX1    g6332(.A(g6346), .Y(g13085));
BUFX1    g6333(.A(g6692), .Y(g13099));
BUFX1    g6334(.A(g1116), .Y(g13259));
BUFX1    g6335(.A(g1459), .Y(g13272));
BUFX1    g6336(.A(g3321), .Y(g13865));
BUFX1    g6337(.A(g3672), .Y(g13881));
BUFX1    g6338(.A(g3281), .Y(g13895));
BUFX1    g6339(.A(g4023), .Y(g13906));
BUFX1    g6340(.A(g3632), .Y(g13926));
BUFX1    g6341(.A(g3983), .Y(g13966));
BUFX1    g6342(.A(g878), .Y(g14096));
BUFX1    g6343(.A(g881), .Y(g14125));
BUFX1    g6344(.A(g884), .Y(g14147));
BUFX1    g6345(.A(g887), .Y(g14167));
BUFX1    g6346(.A(g859), .Y(g14189));
BUFX1    g6347(.A(g869), .Y(g14201));
BUFX1    g6348(.A(g875), .Y(g14217));
BUFX1    g6349(.A(g3298), .Y(g14421));
BUFX1    g6350(.A(g3649), .Y(g14451));
BUFX1    g6351(.A(g4000), .Y(g14518));
BUFX1    g6352(.A(g5331), .Y(g14597));
BUFX1    g6353(.A(g5677), .Y(g14635));
BUFX1    g6354(.A(g5290), .Y(g14662));
BUFX1    g6355(.A(g6023), .Y(g14673));
BUFX1    g6356(.A(g5637), .Y(g14694));
BUFX1    g6357(.A(g6369), .Y(g14705));
BUFX1    g6358(.A(g5983), .Y(g14738));
BUFX1    g6359(.A(g6715), .Y(g14749));
BUFX1    g6360(.A(g6329), .Y(g14779));
BUFX1    g6361(.A(g6675), .Y(g14828));
BUFX1    g6362(.A(g3267), .Y(g16603));
BUFX1    g6363(.A(g3274), .Y(g16624));
BUFX1    g6364(.A(g3618), .Y(g16627));
BUFX1    g6365(.A(g3625), .Y(g16656));
BUFX1    g6366(.A(g3969), .Y(g16659));
BUFX1    g6367(.A(g3325), .Y(g16686));
BUFX1    g6368(.A(g3976), .Y(g16693));
BUFX1    g6369(.A(g3310), .Y(g16718));
BUFX1    g6370(.A(g3676), .Y(g16722));
BUFX1    g6371(.A(g3661), .Y(g16744));
BUFX1    g6372(.A(g4027), .Y(g16748));
BUFX1    g6373(.A(g4012), .Y(g16775));
BUFX1    g6374(.A(g3317), .Y(g16874));
BUFX1    g6375(.A(g3668), .Y(g16924));
BUFX1    g6376(.A(g4019), .Y(g16955));
BUFX1    g6377(.A(g1075), .Y(g17291));
BUFX1    g6378(.A(g1079), .Y(g17316));
BUFX1    g6379(.A(g1418), .Y(g17320));
BUFX1    g6380(.A(g1083), .Y(g17400));
BUFX1    g6381(.A(g1422), .Y(g17404));
BUFX1    g6382(.A(g1426), .Y(g17423));
BUFX1    g6383(.A(g5276), .Y(g17519));
BUFX1    g6384(.A(g5283), .Y(g17577));
BUFX1    g6385(.A(g5623), .Y(g17580));
BUFX1    g6386(.A(g5630), .Y(g17604));
BUFX1    g6387(.A(g5969), .Y(g17607));
BUFX1    g6388(.A(g5335), .Y(g17639));
BUFX1    g6389(.A(g5976), .Y(g17646));
BUFX1    g6390(.A(g6315), .Y(g17649));
BUFX1    g6391(.A(g5320), .Y(g17674));
BUFX1    g6392(.A(g5681), .Y(g17678));
BUFX1    g6393(.A(g6322), .Y(g17685));
BUFX1    g6394(.A(g6661), .Y(g17688));
BUFX1    g6395(.A(g5666), .Y(g17711));
BUFX1    g6396(.A(g6027), .Y(g17715));
BUFX1    g6397(.A(g6668), .Y(g17722));
BUFX1    g6398(.A(g6012), .Y(g17739));
BUFX1    g6399(.A(g6373), .Y(g17743));
BUFX1    g6400(.A(g6358), .Y(g17760));
BUFX1    g6401(.A(g6719), .Y(g17764));
BUFX1    g6402(.A(g6704), .Y(g17778));
BUFX1    g6403(.A(g5327), .Y(g17787));
BUFX1    g6404(.A(g5673), .Y(g17813));
BUFX1    g6405(.A(g6019), .Y(g17819));
BUFX1    g6406(.A(g6365), .Y(g17845));
BUFX1    g6407(.A(g6711), .Y(g17871));
BUFX1    g6408(.A(g6753), .Y(g18092));
BUFX1    g6409(.A(g6748), .Y(g18094));
BUFX1    g6410(.A(g6749), .Y(g18095));
BUFX1    g6411(.A(g6750), .Y(g18096));
BUFX1    g6412(.A(g6747), .Y(g18097));
BUFX1    g6413(.A(g6744), .Y(g18098));
BUFX1    g6414(.A(g6745), .Y(g18099));
BUFX1    g6415(.A(g6751), .Y(g18100));
BUFX1    g6416(.A(g6746), .Y(g18101));
BUFX1    g6417(.A(g66), .Y(g18881));
BUFX1    g6418(.A(g1056), .Y(g19334));
BUFX1    g6419(.A(g1399), .Y(g19357));
BUFX1    g6420(.A(g59), .Y(g20049));
BUFX1    g6421(.A(g86), .Y(g20557));
BUFX1    g6422(.A(g94), .Y(g20652));
BUFX1    g6423(.A(g121), .Y(g20654));
BUFX1    g6424(.A(g74), .Y(g20763));
BUFX1    g6425(.A(g79), .Y(g20899));
BUFX1    g6426(.A(g102), .Y(g20901));
BUFX1    g6427(.A(g106), .Y(g21176));
BUFX1    g6428(.A(g128), .Y(g21245));
BUFX1    g6429(.A(g117), .Y(g21270));
BUFX1    g6430(.A(g136), .Y(g21292));
BUFX1    g6431(.A(g36), .Y(g21698));
BUFX1    g6432(.A(g1242), .Y(g23683));
BUFX1    g6433(.A(g5343), .Y(g25219));
BUFX1    g6434(.A(g59), .Y(g29210));
BUFX1    g6435(.A(g74), .Y(g29211));
BUFX1    g6436(.A(g79), .Y(g29212));
BUFX1    g6437(.A(g86), .Y(g29213));
BUFX1    g6438(.A(g94), .Y(g29214));
BUFX1    g6439(.A(g102), .Y(g29215));
BUFX1    g6440(.A(g106), .Y(g29216));
BUFX1    g6441(.A(g117), .Y(g29217));
BUFX1    g6442(.A(g66), .Y(g29218));
BUFX1    g6443(.A(g121), .Y(g29219));
BUFX1    g6444(.A(g128), .Y(g29220));
BUFX1    g6445(.A(g136), .Y(g29221));
INVX1    g6446(.A(g37), .Y(g30327));
INVX1    g6447(.A(g136), .Y(g30329));
INVX1    g6448(.A(g2834), .Y(g30330));
INVX1    g6449(.A(g2831), .Y(g30331));
BUFX1    g6450(.A(g1242), .Y(g30332));
AND2X1   g6451(.A(g5357), .B(g5297), .Y(g31860));
BUFX1    g6452(.A(g5343), .Y(g31861));
NOR2X1   g6453(.A(g1636), .B(n4631), .Y(g31862));
NOR2X1   g6454(.A(n4629), .B(g1657), .Y(g31863));
NOR3X1   g6455(.A(n4644), .B(n4643), .C(n4642_1), .Y(g32975));
AOI21X1  g6456(.A0(n4668), .A1(n4664), .B0(n4663), .Y(g33533));
AOI21X1  g6457(.A0(n4724), .A1(n4721), .B0(n4719), .Y(g33959));
NAND4X1  g6458(.A(n5061_1), .B(n5045), .C(n5037_1), .D(n5055), .Y(g34234));
NAND4X1  g6459(.A(n5061_1), .B(n5045), .C(n5037_1), .D(n5055), .Y(g34235));
NAND4X1  g6460(.A(n5110), .B(n5106_1), .C(n5100), .D(n5035), .Y(g34238));
NAND4X1  g6461(.A(n5110), .B(n5106_1), .C(n5100), .D(n5035), .Y(g34240));
AOI21X1  g6462(.A0(n4728), .A1(n4727_1), .B0(n4732), .Y(g34435));
NAND2X1  g6463(.A(g2873), .B(g113), .Y(g34436));
NAND2X1  g6464(.A(g2868), .B(g113), .Y(g34437));
NOR2X1   g6465(.A(n4886_1), .B(n4882), .Y(g34788));
AOI21X1  g6466(.A0(n4957), .A1(n5203), .B0(n5202), .Y(g34956));
BUFX1    g6467(.A(g84), .Y(g24168));
BUFX1    g6468(.A(g120), .Y(g24178));
BUFX1    g6469(.A(g113), .Y(g24174));
BUFX1    g6470(.A(g126), .Y(g24181));
BUFX1    g6471(.A(g99), .Y(g24172));
BUFX1    g6472(.A(g53), .Y(g24161));
BUFX1    g6473(.A(g116), .Y(g24177));
BUFX1    g6474(.A(g92), .Y(g24171));
BUFX1    g6475(.A(g56), .Y(g24163));
BUFX1    g6476(.A(g91), .Y(g24170));
BUFX1    g6477(.A(g44), .Y(g24185));
BUFX1    g6478(.A(g57), .Y(g24164));
BUFX1    g6479(.A(g100), .Y(g24173));
BUFX1    g6480(.A(g54), .Y(g24162));
BUFX1    g6481(.A(g124), .Y(g24179));
BUFX1    g6482(.A(g125), .Y(g24180));
BUFX1    g6483(.A(g114), .Y(g24175));
BUFX1    g6484(.A(g134), .Y(g24183));
BUFX1    g6485(.A(g72), .Y(g24166));
BUFX1    g6486(.A(g115), .Y(g24176));
BUFX1    g6487(.A(g135), .Y(g24184));
BUFX1    g6488(.A(g90), .Y(g24169));
BUFX1    g6489(.A(g127), .Y(g24182));
BUFX1    g6490(.A(g64), .Y(g24165));
BUFX1    g6491(.A(g73), .Y(g24167));
BUFX1    g6492(.A(g640), .Y(n720));
BUFX1    g6493(.A(g6027), .Y(n795));
BUFX1    g6494(.A(g4232), .Y(n840));
BUFX1    g6495(.A(g3625), .Y(n855));
BUFX1    g6496(.A(g4571), .Y(n875));
BUFX1    g6497(.A(g6373), .Y(n950));
BUFX1    g6498(.A(g3317), .Y(n1065));
BUFX1    g6499(.A(g3618), .Y(n1090));
BUFX1    g6500(.A(g5623), .Y(n1189));
BUFX1    g6501(.A(g637), .Y(n1229));
BUFX1    g6502(.A(g6012), .Y(n1233));
BUFX1    g6503(.A(g5637), .Y(n1268));
BUFX1    g6504(.A(g6315), .Y(n1298));
BUFX1    g6505(.A(g1418), .Y(n1413));
BUFX1    g6506(.A(g875), .Y(n1443));
BUFX1    g6507(.A(g6668), .Y(n1498));
BUFX1    g6508(.A(g3092), .Y(n1513));
BUFX1    g6509(.A(g6490), .Y(n1523));
BUFX1    g6510(.A(g1576), .Y(n1538));
BUFX1    g6511(.A(g4012), .Y(n1588));
BUFX1    g6512(.A(g6351), .Y(n1623));
BUFX1    g6513(.A(g3661), .Y(n1783));
BUFX1    g6514(.A(g5794), .Y(n1856));
BUFX1    g6515(.A(g802), .Y(n1961));
BUFX1    g6516(.A(g5666), .Y(n1995));
BUFX1    g6517(.A(g6023), .Y(n2074));
BUFX1    g6518(.A(g5335), .Y(n2083));
BUFX1    g6519(.A(g3676), .Y(n2128));
BUFX1    g6520(.A(g1083), .Y(n2153));
BUFX1    g6521(.A(g3794), .Y(n2172));
BUFX1    g6522(.A(g3983), .Y(n2202));
BUFX1    g6523(.A(g6358), .Y(n2251));
BUFX1    g6524(.A(g4277), .Y(n2274));
BUFX1    g6525(.A(g4294), .Y(n2299));
BUFX1    g6526(.A(g6005), .Y(n2303));
BUFX1    g6527(.A(g1399), .Y(n2308));
BUFX1    g6528(.A(g1500), .Y(n2342));
BUFX1    g6529(.A(g5331), .Y(n2472));
BUFX1    g6530(.A(g5798), .Y(n2496));
BUFX1    g6531(.A(g4000), .Y(n2506));
BUFX1    g6532(.A(g3668), .Y(n2516));
BUFX1    g6533(.A(g1426), .Y(n2530));
BUFX1    g6534(.A(g4446), .Y(n2535));
BUFX1    g6535(.A(g6140), .Y(n2554));
BUFX1    g6536(.A(g881), .Y(n2569));
BUFX1    g6537(.A(g4005), .Y(n2674));
BUFX1    g6538(.A(g878), .Y(n2687));
BUFX1    g6539(.A(g1582), .Y(n2705));
BUFX1    g6540(.A(g4222), .Y(n2755));
BUFX1    g6541(.A(g3798), .Y(n2914));
BUFX1    g6542(.A(g5101), .Y(n2954));
BUFX1    g6543(.A(g3654), .Y(n3003));
BUFX1    g6544(.A(g6329), .Y(n3032));
BUFX1    g6545(.A(g4191), .Y(n3061));
BUFX1    g6546(.A(g1570), .Y(n3066));
BUFX1    g6547(.A(g4213), .Y(n3086));
BUFX1    g6548(.A(g3447), .Y(n3121));
BUFX1    g6549(.A(g4304), .Y(n3205));
BUFX1    g6550(.A(g1239), .Y(n3215));
AND2X1   g6551(.A(g125), .B(g35), .Y(n3295));
BUFX1    g6552(.A(g4570), .Y(n3300));
BUFX1    g6553(.A(g3303), .Y(n3304));
BUFX1    g6554(.A(g5327), .Y(n3344));
BUFX1    g6555(.A(g6144), .Y(n3422));
BUFX1    g6556(.A(g859), .Y(n3461));
BUFX1    g6557(.A(g4194), .Y(n3481));
BUFX1    g6558(.A(g5276), .Y(n3486));
BUFX1    g6559(.A(g5452), .Y(n3500));
BUFX1    g6560(.A(g1056), .Y(n3654));
BUFX1    g6561(.A(g6486), .Y(n3669));
BUFX1    g6562(.A(g4414), .Y(n3718));
BUFX1    g6563(.A(g4467), .Y(n3728));
BUFX1    g6564(.A(g5283), .Y(n3732));
BUFX1    g6565(.A(g3976), .Y(n3862));
BUFX1    g6566(.A(g1075), .Y(n3866));
BUFX1    g6567(.A(g6752), .Y(n3901));
BUFX1    g6568(.A(g5313), .Y(n3925));
BUFX1    g6569(.A(g4019), .Y(n3959));
BUFX1    g6570(.A(g4537), .Y(n3964));
BUFX1    g6571(.A(g5681), .Y(n3979));
AND2X1   g6572(.A(g113), .B(g35), .Y(n4009));
BUFX1    g6573(.A(g4449), .Y(n4082));
BUFX1    g6574(.A(g5654), .Y(n4122));
BUFX1    g6575(.A(g1116), .Y(n4136));
BUFX1    g6576(.A(g4207), .Y(n4166));
BUFX1    g6577(.A(g5969), .Y(n4329));
BUFX1    g6578(.A(g884), .Y(n4461));
BUFX1    g6579(.A(g5308), .Y(n4465));
BUFX1    g6580(.A(g6715), .Y(n4539));
BUFX1    g6581(.A(g5677), .Y(n4554));
BUFX1    g6582(.A(g3969), .Y(n4562));
BUFX1    g6583(.A(g1233), .Y(n4590));
BUFX1    g6584(.A(g5983), .Y(n4619));
BUFX1    g6585(.A(g365), .Y(n4622));
BUFX1    g6586(.A(g6697), .Y(n4662));
BUFX1    g6587(.A(g3443), .Y(n4682));
BUFX1    g6588(.A(g3096), .Y(n4717));
BUFX1    g6589(.A(g1227), .Y(n4770));
BUFX1    g6590(.A(g6711), .Y(n4808));
BUFX1    g6591(.A(g194), .Y(n4836));
BUFX1    g6592(.A(g6000), .Y(n4866));
BUFX1    g6593(.A(g3298), .Y(n4906));
BUFX1    g6594(.A(g3649), .Y(n4988));
BUFX1    g6595(.A(g4219), .Y(n5047));
BUFX1    g6596(.A(g6369), .Y(n5111));
BUFX1    g6597(.A(g6365), .Y(n5145));
BUFX1    g6598(.A(g5320), .Y(n5149));
BUFX1    g6599(.A(g4188), .Y(n5162));
BUFX1    g6600(.A(g5290), .Y(n5250));
BUFX1    g6601(.A(g3632), .Y(n5322));
BUFX1    g6602(.A(g4226), .Y(n5330));
BUFX1    g6603(.A(g6346), .Y(n5460));
BUFX1    g6604(.A(g6692), .Y(n5463));
BUFX1    g6605(.A(g4999), .Y(n5511));
BUFX1    g6606(.A(g1459), .Y(n5555));
BUFX1    g6607(.A(g4519), .Y(n5560));
BUFX1    g6608(.A(g4216), .Y(n5564));
BUFX1    g6609(.A(g4027), .Y(n5578));
BUFX1    g6610(.A(g4809), .Y(n5587));
BUFX1    g6611(.A(g4408), .Y(n5611));
BUFX1    g6612(.A(g887), .Y(n5615));
BUFX1    g6613(.A(g344), .Y(n5669));
BUFX1    g6614(.A(g6719), .Y(n5713));
BUFX1    g6615(.A(g3281), .Y(n5787));
BUFX1    g6616(.A(g4287), .Y(n5811));
BUFX1    g6617(.A(g4204), .Y(n5841));
BUFX1    g6618(.A(g215), .Y(n5899));
BUFX1    g6619(.A(g799), .Y(n5996));
BUFX1    g6620(.A(g5976), .Y(n6024));
BUFX1    g6621(.A(g5002), .Y(n6087));
BUFX1    g6622(.A(g6019), .Y(n6096));
BUFX1    g6623(.A(g869), .Y(n6114));
BUFX1    g6624(.A(g1422), .Y(n6132));
AOI22X1  g6625(.A0(n4805), .A1(n4807), .B0(n4804), .B1(n4802), .Y(n6136));
BUFX1    g6626(.A(g4812), .Y(n6170));
BUFX1    g6627(.A(g6322), .Y(n6174));
BUFX1    g6628(.A(g1079), .Y(n6187));
BUFX1    g6629(.A(g3274), .Y(n6351));
BUFX1    g6630(.A(g5005), .Y(n6453));
BUFX1    g6631(.A(g6661), .Y(n6498));
BUFX1    g6632(.A(g4815), .Y(n6526));
BUFX1    g6633(.A(g6675), .Y(n6550));
BUFX1    g6634(.A(g4520), .Y(n6613));
BUFX1    g6635(.A(g4023), .Y(n6662));
AOI22X1  g6636(.A0(n4797), .A1(n4800), .B0(n4796), .B1(n4794), .Y(n6666));
BUFX1    g6637(.A(g4197), .Y(n6685));
BUFX1    g6638(.A(g5105), .Y(n6703));
BUFX1    g6639(.A(g6704), .Y(n6801));
BUFX1    g6640(.A(g5673), .Y(n6868));
BUFX1    g6641(.A(g4185), .Y(n6984));
BUFX1    g6642(.A(g3310), .Y(n7017));
BUFX1    g6643(.A(g3672), .Y(n7051));
BUFX1    g6644(.A(g3325), .Y(n7065));
BUFX1    g6645(.A(g1157), .Y(n7089));
BUFX1    g6646(.A(g5659), .Y(n7221));
BUFX1    g6647(.A(g4229), .Y(n7234));
BUFX1    g6648(.A(g5630), .Y(n7302));
BUFX1    g6649(.A(g3267), .Y(n7310));
BUFX1    g6650(.A(g3321), .Y(n7333));
BUFX1    g6651(.A(g4210), .Y(n7481));
BUFX1    g6652(.A(g5448), .Y(n7515));
BUFX1    g6653(.A(g4200), .Y(n7613));
endmodule
