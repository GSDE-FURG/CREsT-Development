// Benchmark "b15_C" written by ABC on Wed Aug 05 14:41:03 2020

module b15_C ( 
    DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
    DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
    DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
    DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
    DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
    DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
    READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
    M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
    STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
    W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
    BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
    BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
    REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
    REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
    REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
    REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
    REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
    BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
    ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
    ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
    ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
    ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
    ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
    ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
    ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
    ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
    ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
    ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
    ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN,
    ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
    ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN,
    ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN,
    STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
    DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
    DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
    DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
    DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
    DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
    DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
    DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
    DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
    DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
    DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
    DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
    DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
    DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
    DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
    DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
    DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
    STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
    INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
    INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
    INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
    INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
    INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
    INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
    INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
    INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
    INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
    INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
    INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
    INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
    INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
    INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
    INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
    INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
    INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
    INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
    INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
    INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
    INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
    INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
    INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
    INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
    INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
    INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
    INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
    INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
    INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
    INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
    INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
    INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
    INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
    INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
    INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
    INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
    INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
    INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
    INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
    INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
    INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
    INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
    INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
    INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
    INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
    INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
    INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
    INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
    INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
    INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
    INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
    INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
    INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
    INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
    INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
    INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
    INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
    INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
    INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
    INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
    INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
    INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
    INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
    INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
    INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
    INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
    INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
    INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
    INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
    INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
    INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
    INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
    INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
    INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
    INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
    INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
    INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
    INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
    INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
    INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
    INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
    INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
    INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
    INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
    INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
    PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
    PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
    PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
    PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
    PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
    PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
    PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
    PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
    PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
    PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
    PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
    PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
    PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
    PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
    PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
    PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
    LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
    LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
    LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
    LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
    LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
    LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
    UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
    UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
    UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
    UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
    UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
    DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
    DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
    DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
    DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
    DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
    DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
    DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
    DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
    DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
    DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
    EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
    EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
    EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
    EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
    EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
    EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
    EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
    EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
    EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
    EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
    EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
    EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
    EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
    EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
    EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
    EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
    EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
    EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
    EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
    EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
    EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
    EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
    REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
    REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
    REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
    REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
    REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN,
    U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
    U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
    U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
    U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
    U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
    U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
    U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
    U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
    U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
    U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
    U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
    U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
    U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
    U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
    U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
    U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
    U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
    U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
    U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
    U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
    U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
    U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
    U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
    U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
    U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
    U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
    U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
    U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
    U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
    U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
    U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
    U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
    U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
    U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
    U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
    U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
    U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
    U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
    U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
    U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
    U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
    U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
    U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
    U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
    U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788  );
  input  DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_,
    DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_,
    DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_,
    DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_,
    DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_,
    DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N,
    HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN,
    CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN,
    REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN,
    FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
    BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
    BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
    REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
    REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
    REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
    REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
    REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
    BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
    ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
    ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
    ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
    ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
    ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
    ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
    ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
    ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
    ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
    ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
    ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN,
    ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
    ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN,
    ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN,
    STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
    DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
    DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
    DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
    DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
    DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
    DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
    DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
    DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
    DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
    DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
    DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
    DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
    DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
    DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
    DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
    DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
    STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
    INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
    INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
    INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
    INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
    INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
    INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
    INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
    INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
    INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
    INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
    INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
    INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
    INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
    INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
    INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
    INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
    INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
    INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
    INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
    INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
    INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
    INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
    INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
    INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
    INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
    INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
    INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
    INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
    INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
    INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
    INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
    INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
    INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
    INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
    INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
    INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
    INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
    INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
    INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
    INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
    INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
    INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
    INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
    INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
    INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
    INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
    INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
    INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
    INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
    INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
    INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
    INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
    INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
    INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
    INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
    INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
    INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
    INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
    INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
    INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
    INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
    INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
    INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
    INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
    INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
    INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
    INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
    INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
    INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
    INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
    INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
    INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
    INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
    INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
    INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
    INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
    INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
    INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
    INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
    INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
    INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
    INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
    INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
    INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
    INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
    PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
    PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
    PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
    PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
    PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
    PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
    PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
    PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
    PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
    PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
    PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
    PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
    PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
    PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
    PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
    PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
    LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
    LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
    LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
    LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
    LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
    LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
    UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
    UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
    UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
    UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
    UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
    DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
    DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
    DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
    DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
    DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
    DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
    DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
    DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
    DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
    DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
    EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
    EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
    EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
    EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
    EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
    EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
    EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
    EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
    EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
    EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
    EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
    EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
    EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
    EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
    EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
    EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
    EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
    EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
    EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
    EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
    EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
    EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
    REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
    REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
    REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
    REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
    REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
    U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
    U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
    U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
    U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
    U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
    U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
    U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
    U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
    U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
    U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
    U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
    U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
    U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
    U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
    U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
    U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
    U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
    U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
    U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
    U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
    U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
    U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
    U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
    U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
    U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
    U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
    U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
    U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
    U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
    U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
    U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
    U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
    U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
    U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
    U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
    U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
    U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
    U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
    U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
    U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
    U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
    U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
    U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
    U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire n1004, n1005, n1006, n1007, n1009, n1010, n1011, n1012, n1014, n1015,
    n1017, n1018, n1020, n1021, n1022, n1023, n1025, n1026, n1028, n1029,
    n1031, n1032, n1034, n1035, n1037, n1038, n1040, n1041, n1043, n1044,
    n1046, n1047, n1049, n1050, n1052, n1053, n1055, n1056, n1058, n1059,
    n1061, n1062, n1064, n1065, n1067, n1068, n1070, n1071, n1073, n1074,
    n1076, n1077, n1079, n1080, n1082, n1083, n1085, n1086, n1088, n1089,
    n1091, n1092, n1094, n1095, n1097, n1098, n1100, n1101, n1103, n1104,
    n1106, n1107, n1109, n1110, n1112, n1113, n1114, n1115, n1116, n1117,
    n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
    n1128, n1129, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
    n1139, n1141, n1142, n1143, n1144, n1146, n1147, n1148, n1149, n1150,
    n1152, n1153, n1154, n1156, n1158, n1160, n1162, n1164, n1166, n1168,
    n1170, n1172, n1174, n1176, n1178, n1180, n1182, n1184, n1186, n1188,
    n1190, n1192, n1194, n1196, n1198, n1200, n1202, n1204, n1206, n1208,
    n1210, n1212, n1214, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
    n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
    n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
    n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
    n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
    n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
    n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
    n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
    n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
    n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
    n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
    n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
    n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
    n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
    n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
    n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
    n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
    n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
    n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
    n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
    n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
    n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
    n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
    n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
    n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
    n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
    n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
    n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
    n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
    n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
    n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
    n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
    n1533, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
    n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
    n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
    n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
    n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
    n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
    n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
    n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
    n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
    n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
    n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
    n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
    n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
    n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
    n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
    n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
    n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
    n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
    n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
    n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
    n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
    n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
    n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
    n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
    n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
    n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
    n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
    n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
    n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
    n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
    n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
    n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
    n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
    n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
    n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
    n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
    n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
    n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
    n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
    n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
    n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
    n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
    n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
    n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
    n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
    n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
    n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
    n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
    n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
    n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
    n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
    n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
    n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
    n2065, n2066, n2067, n2068, n2070, n2071, n2072, n2073, n2075, n2076,
    n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2086, n2087,
    n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
    n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2108,
    n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
    n2119, n2120, n2121, n2124, n2125, n2127, n2129, n2130, n2131, n2133,
    n2135, n2136, n2138, n2140, n2141, n2142, n2144, n2146, n2147, n2149,
    n2151, n2152, n2153, n2155, n2157, n2158, n2160, n2162, n2163, n2164,
    n2165, n2166, n2167, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
    n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
    n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2195, n2196,
    n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
    n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
    n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
    n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
    n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
    n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
    n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
    n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
    n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
    n2287, n2288, n2289, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
    n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2307, n2308, n2309,
    n2310, n2311, n2312, n2313, n2315, n2316, n2317, n2318, n2319, n2320,
    n2321, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2331, n2332,
    n2333, n2334, n2335, n2336, n2337, n2339, n2340, n2341, n2342, n2343,
    n2344, n2345, n2347, n2348, n2349, n2350, n2353, n2354, n2355, n2358,
    n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
    n2369, n2370, n2371, n2372, n2374, n2375, n2376, n2377, n2379, n2380,
    n2381, n2382, n2384, n2385, n2386, n2387, n2389, n2390, n2391, n2392,
    n2394, n2395, n2396, n2397, n2399, n2400, n2401, n2402, n2404, n2405,
    n2406, n2407, n2409, n2410, n2411, n2412, n2413, n2415, n2416, n2417,
    n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
    n2429, n2430, n2431, n2432, n2434, n2435, n2436, n2437, n2439, n2440,
    n2441, n2442, n2444, n2445, n2446, n2447, n2449, n2450, n2451, n2452,
    n2454, n2455, n2456, n2457, n2459, n2460, n2461, n2462, n2464, n2465,
    n2466, n2467, n2468, n2469, n2470, n2472, n2473, n2474, n2475, n2476,
    n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2486, n2487,
    n2488, n2489, n2491, n2492, n2493, n2494, n2496, n2497, n2498, n2499,
    n2501, n2502, n2503, n2504, n2506, n2507, n2508, n2509, n2511, n2512,
    n2513, n2514, n2516, n2517, n2518, n2519, n2521, n2522, n2523, n2524,
    n2525, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
    n2536, n2537, n2538, n2539, n2541, n2542, n2543, n2544, n2546, n2547,
    n2548, n2549, n2551, n2552, n2553, n2554, n2556, n2557, n2558, n2559,
    n2561, n2562, n2563, n2564, n2566, n2567, n2568, n2569, n2571, n2572,
    n2573, n2574, n2576, n2577, n2578, n2580, n2581, n2582, n2583, n2584,
    n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
    n2596, n2597, n2598, n2599, n2601, n2602, n2603, n2604, n2606, n2607,
    n2608, n2609, n2611, n2612, n2613, n2614, n2616, n2617, n2618, n2619,
    n2621, n2622, n2623, n2624, n2626, n2627, n2628, n2629, n2631, n2632,
    n2633, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
    n2644, n2645, n2646, n2647, n2649, n2650, n2651, n2652, n2654, n2655,
    n2656, n2657, n2659, n2660, n2661, n2662, n2664, n2665, n2666, n2667,
    n2669, n2670, n2671, n2672, n2674, n2675, n2676, n2677, n2679, n2680,
    n2681, n2682, n2684, n2685, n2686, n2687, n2688, n2689, n2691, n2692,
    n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
    n2703, n2704, n2706, n2707, n2708, n2709, n2711, n2712, n2713, n2714,
    n2716, n2717, n2718, n2719, n2721, n2722, n2723, n2724, n2726, n2727,
    n2728, n2729, n2731, n2732, n2733, n2734, n2736, n2737, n2738, n2739,
    n2741, n2742, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
    n2752, n2753, n2754, n2755, n2756, n2757, n2759, n2760, n2761, n2762,
    n2764, n2765, n2766, n2767, n2769, n2770, n2771, n2772, n2774, n2775,
    n2776, n2777, n2779, n2780, n2781, n2782, n2784, n2785, n2786, n2787,
    n2789, n2790, n2791, n2792, n2794, n2795, n2796, n2798, n2799, n2800,
    n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
    n2811, n2813, n2814, n2815, n2816, n2818, n2819, n2820, n2821, n2823,
    n2824, n2825, n2826, n2828, n2829, n2830, n2831, n2833, n2834, n2835,
    n2836, n2838, n2839, n2840, n2841, n2843, n2844, n2845, n2846, n2848,
    n2849, n2850, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
    n2860, n2861, n2862, n2863, n2864, n2866, n2867, n2868, n2869, n2871,
    n2872, n2873, n2874, n2876, n2877, n2878, n2879, n2881, n2882, n2883,
    n2884, n2886, n2887, n2888, n2889, n2891, n2892, n2893, n2894, n2896,
    n2897, n2898, n2899, n2901, n2902, n2903, n2905, n2906, n2907, n2908,
    n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2919,
    n2920, n2921, n2922, n2924, n2925, n2926, n2927, n2929, n2930, n2931,
    n2932, n2934, n2935, n2936, n2937, n2939, n2940, n2941, n2942, n2944,
    n2945, n2946, n2947, n2949, n2950, n2951, n2952, n2954, n2955, n2956,
    n2957, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
    n2968, n2969, n2970, n2971, n2973, n2974, n2975, n2976, n2978, n2979,
    n2980, n2981, n2983, n2984, n2985, n2986, n2988, n2989, n2990, n2991,
    n2993, n2994, n2995, n2996, n2998, n2999, n3000, n3001, n3003, n3004,
    n3005, n3006, n3008, n3009, n3010, n3012, n3013, n3014, n3015, n3016,
    n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3026, n3027,
    n3028, n3029, n3031, n3032, n3033, n3034, n3036, n3037, n3038, n3039,
    n3041, n3042, n3043, n3044, n3046, n3047, n3048, n3049, n3051, n3052,
    n3053, n3054, n3056, n3057, n3058, n3059, n3061, n3062, n3063, n3065,
    n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
    n3076, n3077, n3079, n3080, n3081, n3082, n3084, n3085, n3086, n3087,
    n3089, n3090, n3091, n3092, n3094, n3095, n3096, n3097, n3099, n3100,
    n3101, n3102, n3104, n3105, n3106, n3107, n3109, n3110, n3111, n3112,
    n3114, n3115, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
    n3126, n3127, n3128, n3129, n3130, n3132, n3133, n3134, n3135, n3137,
    n3138, n3139, n3140, n3142, n3143, n3144, n3145, n3147, n3148, n3149,
    n3150, n3152, n3153, n3154, n3155, n3157, n3158, n3159, n3160, n3162,
    n3163, n3164, n3165, n3167, n3168, n3169, n3170, n3171, n3173, n3174,
    n3175, n3177, n3178, n3179, n3180, n3182, n3183, n3184, n3186, n3187,
    n3188, n3189, n3191, n3192, n3193, n3195, n3196, n3197, n3198, n3199,
    n3200, n3201, n3202, n3203, n3204, n3206, n3207, n3208, n3209, n3210,
    n3211, n3215, n3216, n3217, n3219, n3220, n3221, n3222, n3224, n3225,
    n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
    n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
    n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3257,
    n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
    n3268, n3269, n3270, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
    n3279, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
    n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
    n3300, n3301, n3302, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
    n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
    n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
    n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
    n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
    n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3362,
    n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
    n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
    n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
    n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
    n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
    n3413, n3414, n3415, n3416, n3417, n3418, n3420, n3421, n3422, n3423,
    n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
    n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
    n3444, n3445, n3446, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
    n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
    n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
    n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
    n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
    n3496, n3497, n3498, n3499, n3500, n3501, n3503, n3504, n3505, n3506,
    n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
    n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
    n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3539,
    n3540, n3541, n3542, n3543, n3544, n3546, n3547, n3548, n3549, n3550,
    n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
    n3561, n3562, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
    n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
    n3582, n3583, n3584, n3585, n3586, n3588, n3589, n3592, n3595, n3598,
    n3601, n3602, n3605, n3608, n3611, n3614, n3615, n3616, n3617, n3618,
    n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3627, n3628, n3629,
    n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
    n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
    n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
    n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
    n3670, n3671, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
    n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
    n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
    n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
    n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3721,
    n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
    n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
    n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
    n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3762,
    n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
    n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
    n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
    n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3802, n3803,
    n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
    n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
    n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
    n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
    n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
    n3854, n3855, n3856, n3857, n3858, n3859, n3861, n3862, n3863, n3864,
    n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
    n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
    n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
    n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
    n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
    n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
    n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
    n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3946,
    n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
    n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
    n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
    n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
    n3988, n3989, n3990, n3991, n3992, n3996, n3997, n3998, n3999, n4000,
    n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
    n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
    n4021, n4022, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
    n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
    n4042, n4043, n4044, n4045, n4046, n4047, n4049, n4050, n4051, n4052,
    n4053, n4054, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
    n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
    n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4083, n4084, n4086,
    n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
    n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
    n4107, n4109, n4110, n4111, n4112, n4114, n4115, n4116, n4117, n4118,
    n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
    n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
    n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
    n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
    n4161, n4162, n4163, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
    n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
    n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4190, n4191, n4192,
    n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
    n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
    n4213, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
    n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
    n4234, n4235, n4236, n4237, n4238, n4239, n4241, n4242, n4243, n4244,
    n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
    n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
    n4265, n4266, n4267, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
    n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
    n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4296,
    n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
    n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
    n4317, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
    n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
    n4338, n4339, n4340, n4341, n4342, n4344, n4345, n4346, n4347, n4348,
    n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
    n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
    n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
    n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
    n4390, n4391, n4392, n4393, n4395, n4396, n4397, n4398, n4399, n4400,
    n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
    n4411, n4412, n4413, n4414, n4415, n4416, n4418, n4419, n4420, n4421,
    n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
    n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
    n4446, n4447, n4448, n4449, n4450, n4453, n4454, n4455, n4456, n4457,
    n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
    n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4477, n4478,
    n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
    n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
    n4499, n4500, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
    n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4520,
    n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
    n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
    n4541, n4542, n4543, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
    n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
    n4562, n4563, n4564, n4565, n4566, n4567, n4569, n4570, n4571, n4572,
    n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4581, n4582, n4583,
    n4584, n4585, n4586, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
    n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
    n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4613, n4614, n4615,
    n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
    n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
    n4636, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646,
    n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656,
    n4657, n4658, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
    n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
    n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4687, n4688,
    n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
    n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4708, n4709,
    n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
    n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
    n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
    n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
    n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4759, n4760, n4761,
    n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
    n4772, n4773, n4774, n4775, n4777, n4778, n4779, n4780, n4782, n4783,
    n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
    n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
    n4804, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
    n4815, n4816, n4817, n4818, n4823, n4828, n4833, n4838, n4839, n4844,
    n4849, n4854, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866,
    n4867, n4868, n4869, n4870, n4871, n4872, n4874, n4875, n4876, n4877,
    n4878, n4879, n4880, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
    n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
    n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
    n4909, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
    n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
    n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
    n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
    n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
    n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
    n4971, n4972, n4973, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
    n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
    n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
    n5002, n5003, n5005, n5006, n5007, n5008, n5009, n5011, n5012, n5013,
    n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
    n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
    n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
    n5044, n5045, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
    n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
    n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
    n5075, n5076, n5077, n5081, n5084, n5085, n5088, n5091, n5092, n5095,
    n5098, n5101, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
    n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
    n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
    n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
    n5142, n5143, n5144, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
    n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
    n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
    n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5181, n5182, n5183,
    n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
    n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
    n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
    n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5222, n5223, n5224,
    n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
    n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
    n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
    n5255, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
    n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
    n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
    n5286, n5287, n5288, n5289, n5291, n5292, n5293, n5294, n5295, n5296,
    n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306,
    n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
    n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
    n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5336, n5337,
    n5338, n5339, n5340, n5341, n5343, n5344, n5345, n5346, n5347, n5348,
    n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
    n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
    n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5377, n5378, n5379,
    n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
    n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
    n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
    n5410, n5411, n5413, n5414, n5415, n5416, n5419, n5420, n5421, n5422,
    n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
    n5433, n5434, n5435, n5437, n5438, n5439, n5440, n5441, n5442, n5444,
    n5445, n5447, n5448, n5450, n5451, n5453, n5454, n5456, n5457, n5459,
    n5460, n5462, n5463, n5465, n5466, n5468, n5469, n5471, n5472, n5474,
    n5475, n5477, n5478, n5480, n5481, n5483, n5484, n5486, n5487, n5489,
    n5490, n5492, n5493, n5495, n5496, n5498, n5499, n5501, n5502, n5504,
    n5505, n5507, n5508, n5510, n5511, n5513, n5514, n5516, n5517, n5519,
    n5520, n5522, n5523, n5525, n5526, n5528, n5529, n5531, n5532, n5534,
    n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5543, n5545, n5547,
    n5548, n5550, n5552, n5553, n5555, n5556, n5558, n5559, n5561, n5562,
    n5564, n5565, n5567, n5568, n5570, n5571, n5573, n5574, n5576, n5578,
    n5580, n5582, n5583, n5584, n5586, n5587, n5589, n5590, n5592, n5593,
    n5595, n5596, n5598, n5599, n5601, n5602, n5604, n5605, n5607, n5609,
    n5611, n5613, n5614, n5616, n5618, n5620, n5621, n5623, n5625, n5626,
    n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5637,
    n5639, n5641, n5642, n5644, n5646, n5648, n5649, n5651, n5653, n5654,
    n5656, n5658, n5660, n5661, n5663, n5665, n5667, n5668, n5669, n5671,
    n5672, n5673, n5674, n5676, n5677, n5678, n5679, n5680, n5681, n5683,
    n5684, n5685, n5687, n5688, n5690, n5691, n5692, n5694, n5695, n5696,
    n5698, n5699, n5700, n5701, n5703, n5704, n5705, n5707, n5708, n5709,
    n5711, n5712, n5713, n5714, n5716, n5717, n5718, n5719, n5721, n5722,
    n5723, n5725, n5726, n5727, n5728, n5730, n5731, n5732, n5733, n5734,
    n5736, n5737, n5738, n5739, n5740, n5742, n5743, n5744, n5745, n5746,
    n5748, n5749, n5750, n5751, n5753, n5754, n5755, n5756, n5757, n5758,
    n5759, n5760, n5761, n5763, n5765, n5767, n5768, n5770, n5771, n5773,
    n5774, n5776, n5777, n5779, n5780, n5782, n5783, n5785, n5786, n5788,
    n5789, n5791, n5792, n5794, n5795, n5797, n5798, n5800, n5801, n5803,
    n5804, n5806, n5807, n5809, n5810, n5812, n5813, n5815, n5816, n5818,
    n5820, n5821, n5823, n5824, n5826, n5827, n5829, n5830, n5832, n5834,
    n5835, n5837, n5839, n5840, n5841, n5843, n5845, n5846, n5848, n5850,
    n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
    n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
    n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5881,
    n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5892,
    n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5901, n5902, n5903,
    n5904, n5905, n5906, n5907, n5908, n5910, n5911, n5912, n5913, n5914,
    n5915, n5916, n5917, n5918, n5919, n5921, n5922, n5923, n5924, n5925,
    n5926, n5927, n5928, n5929, n5930, n5932, n5933, n5934, n5935, n5936,
    n5937, n5938, n5939, n5940, n5941, n5943, n5944, n5945, n5946, n5947,
    n5948, n5949, n5950, n5951, n5953, n5954, n5955, n5956, n5957, n5958,
    n5959, n5960, n5961, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
    n5970, n5971, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
    n5981, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
    n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6003,
    n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6013, n6014,
    n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6023, n6024, n6025,
    n6026, n6027, n6028, n6029, n6030, n6031, n6033, n6034, n6035, n6036,
    n6037, n6038, n6039, n6040, n6041, n6043, n6044, n6045, n6046, n6047,
    n6048, n6049, n6050, n6051, n6053, n6054, n6055, n6056, n6057, n6058,
    n6059, n6060, n6061, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
    n6070, n6071, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
    n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6091, n6092,
    n6093, n6094, n6095, n6096, n6097, n6098, n6100, n6101, n6102, n6103,
    n6104, n6105, n6106, n6107, n6109, n6110, n6111, n6112, n6113, n6114,
    n6115, n6116, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
    n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6136, n6137,
    n6138, n6139, n6140, n6141, n6142, n6143, n6145, n6146, n6147, n6148,
    n6149, n6150, n6151, n6152, n6153, n6155, n6156, n6157, n6158, n6159,
    n6160, n6161, n6162, n6163, n6165, n6166, n6167, n6168, n6169, n6170,
    n6171, n6172, n6173, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
    n6182, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
    n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6202, n6203,
    n6204, n6205, n6207, n6208, n6210, n6212, n6214, n6216, n6217, n6219,
    n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6229, n6230, n6231,
    n6233, n6234, n6236, n6237, n6239, n6241, n6242, n6243, n6244, n6246,
    n6247, n6248, n6249;
  INVX1   g0000(.A(STATE_REG_0__SCAN_IN), .Y(n1004));
  NAND3X1 g0001(.A(n1004), .B(STATE_REG_1__SCAN_IN), .C(BYTEENABLE_REG_3__SCAN_IN), .Y(n1005));
  INVX1   g0002(.A(STATE_REG_1__SCAN_IN), .Y(n1006));
  OAI21X1 g0003(.A0(STATE_REG_0__SCAN_IN), .A1(n1006), .B0(BE_N_REG_3__SCAN_IN), .Y(n1007));
  NAND2X1 g0004(.A(n1007), .B(n1005), .Y(U3445));
  INVX1   g0005(.A(BYTEENABLE_REG_2__SCAN_IN), .Y(n1009));
  NOR2X1  g0006(.A(STATE_REG_0__SCAN_IN), .B(n1006), .Y(n1010));
  INVX1   g0007(.A(n1010), .Y(n1011));
  OAI21X1 g0008(.A0(STATE_REG_0__SCAN_IN), .A1(n1006), .B0(BE_N_REG_2__SCAN_IN), .Y(n1012));
  OAI21X1 g0009(.A0(n1011), .A1(n1009), .B0(n1012), .Y(U3446));
  NAND3X1 g0010(.A(n1004), .B(STATE_REG_1__SCAN_IN), .C(BYTEENABLE_REG_1__SCAN_IN), .Y(n1014));
  OAI21X1 g0011(.A0(STATE_REG_0__SCAN_IN), .A1(n1006), .B0(BE_N_REG_1__SCAN_IN), .Y(n1015));
  NAND2X1 g0012(.A(n1015), .B(n1014), .Y(U3447));
  INVX1   g0013(.A(BYTEENABLE_REG_0__SCAN_IN), .Y(n1017));
  OAI21X1 g0014(.A0(STATE_REG_0__SCAN_IN), .A1(n1006), .B0(BE_N_REG_0__SCAN_IN), .Y(n1018));
  OAI21X1 g0015(.A0(n1011), .A1(n1017), .B0(n1018), .Y(U3448));
  INVX1   g0016(.A(REIP_REG_30__SCAN_IN), .Y(n1020));
  NAND3X1 g0017(.A(n1004), .B(STATE_REG_1__SCAN_IN), .C(STATE_REG_2__SCAN_IN), .Y(n1021));
  NOR3X1  g0018(.A(STATE_REG_0__SCAN_IN), .B(n1006), .C(STATE_REG_2__SCAN_IN), .Y(n1022));
  AOI22X1 g0019(.A0(n1011), .A1(ADDRESS_REG_29__SCAN_IN), .B0(REIP_REG_31__SCAN_IN), .B1(n1022), .Y(n1023));
  OAI21X1 g0020(.A0(n1021), .A1(n1020), .B0(n1023), .Y(U3213));
  INVX1   g0021(.A(REIP_REG_29__SCAN_IN), .Y(n1025));
  AOI22X1 g0022(.A0(n1011), .A1(ADDRESS_REG_28__SCAN_IN), .B0(REIP_REG_30__SCAN_IN), .B1(n1022), .Y(n1026));
  OAI21X1 g0023(.A0(n1021), .A1(n1025), .B0(n1026), .Y(U3212));
  INVX1   g0024(.A(REIP_REG_28__SCAN_IN), .Y(n1028));
  AOI22X1 g0025(.A0(n1011), .A1(ADDRESS_REG_27__SCAN_IN), .B0(REIP_REG_29__SCAN_IN), .B1(n1022), .Y(n1029));
  OAI21X1 g0026(.A0(n1021), .A1(n1028), .B0(n1029), .Y(U3211));
  INVX1   g0027(.A(REIP_REG_27__SCAN_IN), .Y(n1031));
  AOI22X1 g0028(.A0(n1011), .A1(ADDRESS_REG_26__SCAN_IN), .B0(REIP_REG_28__SCAN_IN), .B1(n1022), .Y(n1032));
  OAI21X1 g0029(.A0(n1021), .A1(n1031), .B0(n1032), .Y(U3210));
  INVX1   g0030(.A(REIP_REG_26__SCAN_IN), .Y(n1034));
  AOI22X1 g0031(.A0(n1011), .A1(ADDRESS_REG_25__SCAN_IN), .B0(REIP_REG_27__SCAN_IN), .B1(n1022), .Y(n1035));
  OAI21X1 g0032(.A0(n1021), .A1(n1034), .B0(n1035), .Y(U3209));
  INVX1   g0033(.A(REIP_REG_25__SCAN_IN), .Y(n1037));
  AOI22X1 g0034(.A0(n1011), .A1(ADDRESS_REG_24__SCAN_IN), .B0(REIP_REG_26__SCAN_IN), .B1(n1022), .Y(n1038));
  OAI21X1 g0035(.A0(n1021), .A1(n1037), .B0(n1038), .Y(U3208));
  INVX1   g0036(.A(REIP_REG_24__SCAN_IN), .Y(n1040));
  AOI22X1 g0037(.A0(n1011), .A1(ADDRESS_REG_23__SCAN_IN), .B0(REIP_REG_25__SCAN_IN), .B1(n1022), .Y(n1041));
  OAI21X1 g0038(.A0(n1021), .A1(n1040), .B0(n1041), .Y(U3207));
  INVX1   g0039(.A(REIP_REG_23__SCAN_IN), .Y(n1043));
  AOI22X1 g0040(.A0(n1011), .A1(ADDRESS_REG_22__SCAN_IN), .B0(REIP_REG_24__SCAN_IN), .B1(n1022), .Y(n1044));
  OAI21X1 g0041(.A0(n1021), .A1(n1043), .B0(n1044), .Y(U3206));
  INVX1   g0042(.A(REIP_REG_22__SCAN_IN), .Y(n1046));
  AOI22X1 g0043(.A0(n1011), .A1(ADDRESS_REG_21__SCAN_IN), .B0(REIP_REG_23__SCAN_IN), .B1(n1022), .Y(n1047));
  OAI21X1 g0044(.A0(n1021), .A1(n1046), .B0(n1047), .Y(U3205));
  INVX1   g0045(.A(REIP_REG_21__SCAN_IN), .Y(n1049));
  AOI22X1 g0046(.A0(n1011), .A1(ADDRESS_REG_20__SCAN_IN), .B0(REIP_REG_22__SCAN_IN), .B1(n1022), .Y(n1050));
  OAI21X1 g0047(.A0(n1021), .A1(n1049), .B0(n1050), .Y(U3204));
  INVX1   g0048(.A(REIP_REG_20__SCAN_IN), .Y(n1052));
  AOI22X1 g0049(.A0(n1011), .A1(ADDRESS_REG_19__SCAN_IN), .B0(REIP_REG_21__SCAN_IN), .B1(n1022), .Y(n1053));
  OAI21X1 g0050(.A0(n1021), .A1(n1052), .B0(n1053), .Y(U3203));
  INVX1   g0051(.A(REIP_REG_19__SCAN_IN), .Y(n1055));
  AOI22X1 g0052(.A0(n1011), .A1(ADDRESS_REG_18__SCAN_IN), .B0(REIP_REG_20__SCAN_IN), .B1(n1022), .Y(n1056));
  OAI21X1 g0053(.A0(n1021), .A1(n1055), .B0(n1056), .Y(U3202));
  INVX1   g0054(.A(REIP_REG_18__SCAN_IN), .Y(n1058));
  AOI22X1 g0055(.A0(n1011), .A1(ADDRESS_REG_17__SCAN_IN), .B0(REIP_REG_19__SCAN_IN), .B1(n1022), .Y(n1059));
  OAI21X1 g0056(.A0(n1021), .A1(n1058), .B0(n1059), .Y(U3201));
  INVX1   g0057(.A(REIP_REG_17__SCAN_IN), .Y(n1061));
  AOI22X1 g0058(.A0(n1011), .A1(ADDRESS_REG_16__SCAN_IN), .B0(REIP_REG_18__SCAN_IN), .B1(n1022), .Y(n1062));
  OAI21X1 g0059(.A0(n1021), .A1(n1061), .B0(n1062), .Y(U3200));
  INVX1   g0060(.A(REIP_REG_16__SCAN_IN), .Y(n1064));
  AOI22X1 g0061(.A0(n1011), .A1(ADDRESS_REG_15__SCAN_IN), .B0(REIP_REG_17__SCAN_IN), .B1(n1022), .Y(n1065));
  OAI21X1 g0062(.A0(n1021), .A1(n1064), .B0(n1065), .Y(U3199));
  INVX1   g0063(.A(REIP_REG_15__SCAN_IN), .Y(n1067));
  AOI22X1 g0064(.A0(n1011), .A1(ADDRESS_REG_14__SCAN_IN), .B0(REIP_REG_16__SCAN_IN), .B1(n1022), .Y(n1068));
  OAI21X1 g0065(.A0(n1021), .A1(n1067), .B0(n1068), .Y(U3198));
  INVX1   g0066(.A(REIP_REG_14__SCAN_IN), .Y(n1070));
  AOI22X1 g0067(.A0(n1011), .A1(ADDRESS_REG_13__SCAN_IN), .B0(REIP_REG_15__SCAN_IN), .B1(n1022), .Y(n1071));
  OAI21X1 g0068(.A0(n1021), .A1(n1070), .B0(n1071), .Y(U3197));
  INVX1   g0069(.A(REIP_REG_13__SCAN_IN), .Y(n1073));
  AOI22X1 g0070(.A0(n1011), .A1(ADDRESS_REG_12__SCAN_IN), .B0(REIP_REG_14__SCAN_IN), .B1(n1022), .Y(n1074));
  OAI21X1 g0071(.A0(n1021), .A1(n1073), .B0(n1074), .Y(U3196));
  INVX1   g0072(.A(REIP_REG_12__SCAN_IN), .Y(n1076));
  AOI22X1 g0073(.A0(n1011), .A1(ADDRESS_REG_11__SCAN_IN), .B0(REIP_REG_13__SCAN_IN), .B1(n1022), .Y(n1077));
  OAI21X1 g0074(.A0(n1021), .A1(n1076), .B0(n1077), .Y(U3195));
  INVX1   g0075(.A(REIP_REG_11__SCAN_IN), .Y(n1079));
  AOI22X1 g0076(.A0(n1011), .A1(ADDRESS_REG_10__SCAN_IN), .B0(REIP_REG_12__SCAN_IN), .B1(n1022), .Y(n1080));
  OAI21X1 g0077(.A0(n1021), .A1(n1079), .B0(n1080), .Y(U3194));
  INVX1   g0078(.A(REIP_REG_10__SCAN_IN), .Y(n1082));
  AOI22X1 g0079(.A0(n1011), .A1(ADDRESS_REG_9__SCAN_IN), .B0(REIP_REG_11__SCAN_IN), .B1(n1022), .Y(n1083));
  OAI21X1 g0080(.A0(n1021), .A1(n1082), .B0(n1083), .Y(U3193));
  INVX1   g0081(.A(REIP_REG_9__SCAN_IN), .Y(n1085));
  AOI22X1 g0082(.A0(n1011), .A1(ADDRESS_REG_8__SCAN_IN), .B0(REIP_REG_10__SCAN_IN), .B1(n1022), .Y(n1086));
  OAI21X1 g0083(.A0(n1021), .A1(n1085), .B0(n1086), .Y(U3192));
  INVX1   g0084(.A(REIP_REG_8__SCAN_IN), .Y(n1088));
  AOI22X1 g0085(.A0(n1011), .A1(ADDRESS_REG_7__SCAN_IN), .B0(REIP_REG_9__SCAN_IN), .B1(n1022), .Y(n1089));
  OAI21X1 g0086(.A0(n1021), .A1(n1088), .B0(n1089), .Y(U3191));
  INVX1   g0087(.A(REIP_REG_7__SCAN_IN), .Y(n1091));
  AOI22X1 g0088(.A0(n1011), .A1(ADDRESS_REG_6__SCAN_IN), .B0(REIP_REG_8__SCAN_IN), .B1(n1022), .Y(n1092));
  OAI21X1 g0089(.A0(n1021), .A1(n1091), .B0(n1092), .Y(U3190));
  INVX1   g0090(.A(REIP_REG_6__SCAN_IN), .Y(n1094));
  AOI22X1 g0091(.A0(n1011), .A1(ADDRESS_REG_5__SCAN_IN), .B0(REIP_REG_7__SCAN_IN), .B1(n1022), .Y(n1095));
  OAI21X1 g0092(.A0(n1021), .A1(n1094), .B0(n1095), .Y(U3189));
  INVX1   g0093(.A(REIP_REG_5__SCAN_IN), .Y(n1097));
  AOI22X1 g0094(.A0(n1011), .A1(ADDRESS_REG_4__SCAN_IN), .B0(REIP_REG_6__SCAN_IN), .B1(n1022), .Y(n1098));
  OAI21X1 g0095(.A0(n1021), .A1(n1097), .B0(n1098), .Y(U3188));
  INVX1   g0096(.A(REIP_REG_4__SCAN_IN), .Y(n1100));
  AOI22X1 g0097(.A0(n1011), .A1(ADDRESS_REG_3__SCAN_IN), .B0(REIP_REG_5__SCAN_IN), .B1(n1022), .Y(n1101));
  OAI21X1 g0098(.A0(n1021), .A1(n1100), .B0(n1101), .Y(U3187));
  INVX1   g0099(.A(REIP_REG_3__SCAN_IN), .Y(n1103));
  AOI22X1 g0100(.A0(n1011), .A1(ADDRESS_REG_2__SCAN_IN), .B0(REIP_REG_4__SCAN_IN), .B1(n1022), .Y(n1104));
  OAI21X1 g0101(.A0(n1021), .A1(n1103), .B0(n1104), .Y(U3186));
  INVX1   g0102(.A(REIP_REG_2__SCAN_IN), .Y(n1106));
  AOI22X1 g0103(.A0(n1011), .A1(ADDRESS_REG_1__SCAN_IN), .B0(REIP_REG_3__SCAN_IN), .B1(n1022), .Y(n1107));
  OAI21X1 g0104(.A0(n1021), .A1(n1106), .B0(n1107), .Y(U3185));
  INVX1   g0105(.A(REIP_REG_1__SCAN_IN), .Y(n1109));
  AOI22X1 g0106(.A0(n1011), .A1(ADDRESS_REG_0__SCAN_IN), .B0(REIP_REG_2__SCAN_IN), .B1(n1022), .Y(n1110));
  OAI21X1 g0107(.A0(n1021), .A1(n1109), .B0(n1110), .Y(U3184));
  INVX1   g0108(.A(STATE_REG_2__SCAN_IN), .Y(n1112));
  INVX1   g0109(.A(READY_N), .Y(n1113));
  NOR2X1  g0110(.A(REQUESTPENDING_REG_SCAN_IN), .B(HOLD), .Y(n1114));
  NAND2X1 g0111(.A(n1114), .B(n1113), .Y(n1115));
  INVX1   g0112(.A(REQUESTPENDING_REG_SCAN_IN), .Y(n1116));
  NOR2X1  g0113(.A(n1116), .B(HOLD), .Y(n1117));
  AOI21X1 g0114(.A0(n1117), .A1(n1113), .B0(n1006), .Y(n1118));
  OAI21X1 g0115(.A0(n1116), .A1(HOLD), .B0(STATE_REG_0__SCAN_IN), .Y(n1119));
  OAI22X1 g0116(.A0(n1114), .A1(n1119), .B0(STATE_REG_0__SCAN_IN), .B1(NA_N), .Y(n1120));
  AOI21X1 g0117(.A0(n1118), .A1(n1115), .B0(n1120), .Y(n1121));
  NAND2X1 g0118(.A(STATE_REG_1__SCAN_IN), .B(READY_N), .Y(n1122));
  NOR2X1  g0119(.A(STATE_REG_1__SCAN_IN), .B(STATE_REG_2__SCAN_IN), .Y(n1123));
  NAND3X1 g0120(.A(n1123), .B(n1116), .C(HOLD), .Y(n1124));
  OAI21X1 g0121(.A0(n1122), .A1(n1114), .B0(n1124), .Y(n1125));
  INVX1   g0122(.A(NA_N), .Y(n1126));
  NOR3X1  g0123(.A(n1006), .B(STATE_REG_2__SCAN_IN), .C(n1126), .Y(n1127));
  NOR2X1  g0124(.A(n1127), .B(n1004), .Y(n1128));
  AOI22X1 g0125(.A0(n1125), .A1(n1128), .B0(n1010), .B1(STATE_REG_2__SCAN_IN), .Y(n1129));
  OAI21X1 g0126(.A0(n1121), .A1(n1112), .B0(n1129), .Y(U3183));
  NAND2X1 g0127(.A(STATE_REG_0__SCAN_IN), .B(REQUESTPENDING_REG_SCAN_IN), .Y(n1131));
  NOR2X1  g0128(.A(n1131), .B(STATE_REG_2__SCAN_IN), .Y(n1132));
  AOI21X1 g0129(.A0(n1119), .A1(STATE_REG_2__SCAN_IN), .B0(n1132), .Y(n1133));
  INVX1   g0130(.A(HOLD), .Y(n1134));
  OAI21X1 g0131(.A0(n1134), .A1(READY_N), .B0(STATE_REG_0__SCAN_IN), .Y(n1135));
  NAND2X1 g0132(.A(n1115), .B(STATE_REG_1__SCAN_IN), .Y(n1136));
  AOI21X1 g0133(.A0(n1135), .A1(STATE_REG_2__SCAN_IN), .B0(n1136), .Y(n1137));
  AOI21X1 g0134(.A0(STATE_REG_2__SCAN_IN), .A1(n1113), .B0(n1011), .Y(n1138));
  NOR2X1  g0135(.A(n1138), .B(n1137), .Y(n1139));
  OAI21X1 g0136(.A0(n1133), .A1(STATE_REG_1__SCAN_IN), .B0(n1139), .Y(U3182));
  OAI21X1 g0137(.A0(n1131), .A1(n1118), .B0(n1112), .Y(n1141));
  OAI22X1 g0138(.A0(STATE_REG_0__SCAN_IN), .A1(n1126), .B0(n1112), .B1(n1117), .Y(n1142));
  NOR3X1  g0139(.A(n1117), .B(n1004), .C(n1112), .Y(n1143));
  AOI21X1 g0140(.A0(n1142), .A1(n1006), .B0(n1143), .Y(n1144));
  NAND2X1 g0141(.A(n1144), .B(n1141), .Y(U3181));
  INVX1   g0142(.A(BS16_N), .Y(n1146));
  OAI21X1 g0143(.A0(STATE_REG_1__SCAN_IN), .A1(STATE_REG_2__SCAN_IN), .B0(n1146), .Y(n1147));
  NOR3X1  g0144(.A(n1004), .B(n1006), .C(STATE_REG_2__SCAN_IN), .Y(n1148));
  AOI21X1 g0145(.A0(n1004), .A1(n1006), .B0(n1148), .Y(n1149));
  NAND2X1 g0146(.A(n1149), .B(DATAWIDTH_REG_0__SCAN_IN), .Y(n1150));
  OAI21X1 g0147(.A0(n1149), .A1(n1147), .B0(n1150), .Y(U3451));
  INVX1   g0148(.A(DATAWIDTH_REG_1__SCAN_IN), .Y(n1152));
  INVX1   g0149(.A(n1149), .Y(n1153));
  NAND2X1 g0150(.A(n1153), .B(n1147), .Y(n1154));
  OAI21X1 g0151(.A0(n1153), .A1(n1152), .B0(n1154), .Y(U3452));
  INVX1   g0152(.A(DATAWIDTH_REG_2__SCAN_IN), .Y(n1156));
  NOR2X1  g0153(.A(n1153), .B(n1156), .Y(U3180));
  INVX1   g0154(.A(DATAWIDTH_REG_3__SCAN_IN), .Y(n1158));
  NOR2X1  g0155(.A(n1153), .B(n1158), .Y(U3179));
  INVX1   g0156(.A(DATAWIDTH_REG_4__SCAN_IN), .Y(n1160));
  NOR2X1  g0157(.A(n1153), .B(n1160), .Y(U3178));
  INVX1   g0158(.A(DATAWIDTH_REG_5__SCAN_IN), .Y(n1162));
  NOR2X1  g0159(.A(n1153), .B(n1162), .Y(U3177));
  INVX1   g0160(.A(DATAWIDTH_REG_6__SCAN_IN), .Y(n1164));
  NOR2X1  g0161(.A(n1153), .B(n1164), .Y(U3176));
  INVX1   g0162(.A(DATAWIDTH_REG_7__SCAN_IN), .Y(n1166));
  NOR2X1  g0163(.A(n1153), .B(n1166), .Y(U3175));
  INVX1   g0164(.A(DATAWIDTH_REG_8__SCAN_IN), .Y(n1168));
  NOR2X1  g0165(.A(n1153), .B(n1168), .Y(U3174));
  INVX1   g0166(.A(DATAWIDTH_REG_9__SCAN_IN), .Y(n1170));
  NOR2X1  g0167(.A(n1153), .B(n1170), .Y(U3173));
  INVX1   g0168(.A(DATAWIDTH_REG_10__SCAN_IN), .Y(n1172));
  NOR2X1  g0169(.A(n1153), .B(n1172), .Y(U3172));
  INVX1   g0170(.A(DATAWIDTH_REG_11__SCAN_IN), .Y(n1174));
  NOR2X1  g0171(.A(n1153), .B(n1174), .Y(U3171));
  INVX1   g0172(.A(DATAWIDTH_REG_12__SCAN_IN), .Y(n1176));
  NOR2X1  g0173(.A(n1153), .B(n1176), .Y(U3170));
  INVX1   g0174(.A(DATAWIDTH_REG_13__SCAN_IN), .Y(n1178));
  NOR2X1  g0175(.A(n1153), .B(n1178), .Y(U3169));
  INVX1   g0176(.A(DATAWIDTH_REG_14__SCAN_IN), .Y(n1180));
  NOR2X1  g0177(.A(n1153), .B(n1180), .Y(U3168));
  INVX1   g0178(.A(DATAWIDTH_REG_15__SCAN_IN), .Y(n1182));
  NOR2X1  g0179(.A(n1153), .B(n1182), .Y(U3167));
  INVX1   g0180(.A(DATAWIDTH_REG_16__SCAN_IN), .Y(n1184));
  NOR2X1  g0181(.A(n1153), .B(n1184), .Y(U3166));
  INVX1   g0182(.A(DATAWIDTH_REG_17__SCAN_IN), .Y(n1186));
  NOR2X1  g0183(.A(n1153), .B(n1186), .Y(U3165));
  INVX1   g0184(.A(DATAWIDTH_REG_18__SCAN_IN), .Y(n1188));
  NOR2X1  g0185(.A(n1153), .B(n1188), .Y(U3164));
  INVX1   g0186(.A(DATAWIDTH_REG_19__SCAN_IN), .Y(n1190));
  NOR2X1  g0187(.A(n1153), .B(n1190), .Y(U3163));
  INVX1   g0188(.A(DATAWIDTH_REG_20__SCAN_IN), .Y(n1192));
  NOR2X1  g0189(.A(n1153), .B(n1192), .Y(U3162));
  INVX1   g0190(.A(DATAWIDTH_REG_21__SCAN_IN), .Y(n1194));
  NOR2X1  g0191(.A(n1153), .B(n1194), .Y(U3161));
  INVX1   g0192(.A(DATAWIDTH_REG_22__SCAN_IN), .Y(n1196));
  NOR2X1  g0193(.A(n1153), .B(n1196), .Y(U3160));
  INVX1   g0194(.A(DATAWIDTH_REG_23__SCAN_IN), .Y(n1198));
  NOR2X1  g0195(.A(n1153), .B(n1198), .Y(U3159));
  INVX1   g0196(.A(DATAWIDTH_REG_24__SCAN_IN), .Y(n1200));
  NOR2X1  g0197(.A(n1153), .B(n1200), .Y(U3158));
  INVX1   g0198(.A(DATAWIDTH_REG_25__SCAN_IN), .Y(n1202));
  NOR2X1  g0199(.A(n1153), .B(n1202), .Y(U3157));
  INVX1   g0200(.A(DATAWIDTH_REG_26__SCAN_IN), .Y(n1204));
  NOR2X1  g0201(.A(n1153), .B(n1204), .Y(U3156));
  INVX1   g0202(.A(DATAWIDTH_REG_27__SCAN_IN), .Y(n1206));
  NOR2X1  g0203(.A(n1153), .B(n1206), .Y(U3155));
  INVX1   g0204(.A(DATAWIDTH_REG_28__SCAN_IN), .Y(n1208));
  NOR2X1  g0205(.A(n1153), .B(n1208), .Y(U3154));
  INVX1   g0206(.A(DATAWIDTH_REG_29__SCAN_IN), .Y(n1210));
  NOR2X1  g0207(.A(n1153), .B(n1210), .Y(U3153));
  INVX1   g0208(.A(DATAWIDTH_REG_30__SCAN_IN), .Y(n1212));
  NOR2X1  g0209(.A(n1153), .B(n1212), .Y(U3152));
  INVX1   g0210(.A(DATAWIDTH_REG_31__SCAN_IN), .Y(n1214));
  NOR2X1  g0211(.A(n1153), .B(n1214), .Y(U3151));
  INVX1   g0212(.A(STATE2_REG_3__SCAN_IN), .Y(n1216));
  INVX1   g0213(.A(STATE2_REG_0__SCAN_IN), .Y(n1217));
  INVX1   g0214(.A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .Y(n1218));
  NOR2X1  g0215(.A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B(n1218), .Y(n1219));
  INVX1   g0216(.A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .Y(n1220));
  NOR2X1  g0217(.A(n1220), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n1221));
  INVX1   g0218(.A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n1222));
  NOR2X1  g0219(.A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n1222), .Y(n1223));
  INVX1   g0220(.A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .Y(n1224));
  NOR2X1  g0221(.A(n1224), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Y(n1225));
  INVX1   g0222(.A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Y(n1226));
  NOR2X1  g0223(.A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n1226), .Y(n1227));
  INVX1   g0224(.A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Y(n1228));
  INVX1   g0225(.A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Y(n1229));
  AOI21X1 g0226(.A0(n1229), .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B0(n1228), .Y(n1230));
  INVX1   g0227(.A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n1231));
  NOR2X1  g0228(.A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n1231), .Y(n1232));
  AOI21X1 g0229(.A0(n1232), .A1(n1228), .B0(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Y(n1233));
  NOR2X1  g0230(.A(n1233), .B(n1230), .Y(n1234));
  NOR2X1  g0231(.A(n1234), .B(n1227), .Y(n1235));
  NOR2X1  g0232(.A(n1235), .B(n1225), .Y(n1236));
  NOR2X1  g0233(.A(n1236), .B(n1223), .Y(n1237));
  INVX1   g0234(.A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .Y(n1238));
  NOR2X1  g0235(.A(n1238), .B(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .Y(n1239));
  NOR3X1  g0236(.A(n1239), .B(n1237), .C(n1221), .Y(n1240));
  NOR2X1  g0237(.A(n1240), .B(n1219), .Y(n1241));
  INVX1   g0238(.A(INSTQUEUE_REG_7__0__SCAN_IN), .Y(n1242));
  NAND4X1 g0239(.A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(n1222), .D(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n1243));
  NOR4X1  g0240(.A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .D(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n1244));
  INVX1   g0241(.A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Y(n1245));
  NOR4X1  g0242(.A(n1245), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .D(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n1246));
  AOI22X1 g0243(.A0(n1244), .A1(INSTQUEUE_REG_0__0__SCAN_IN), .B0(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n1246), .Y(n1247));
  OAI21X1 g0244(.A0(n1243), .A1(n1242), .B0(n1247), .Y(n1248));
  INVX1   g0245(.A(INSTQUEUE_REG_4__0__SCAN_IN), .Y(n1249));
  NOR2X1  g0246(.A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Y(n1250));
  NAND3X1 g0247(.A(n1250), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(n1222), .Y(n1251));
  NAND2X1 g0248(.A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Y(n1252));
  NOR3X1  g0249(.A(n1252), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(n1222), .Y(n1253));
  NAND2X1 g0250(.A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n1254));
  NOR3X1  g0251(.A(n1254), .B(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Y(n1255));
  AOI22X1 g0252(.A0(n1253), .A1(INSTQUEUE_REG_11__0__SCAN_IN), .B0(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n1255), .Y(n1256));
  OAI21X1 g0253(.A0(n1251), .A1(n1249), .B0(n1256), .Y(n1257));
  INVX1   g0254(.A(INSTQUEUE_REG_8__0__SCAN_IN), .Y(n1258));
  INVX1   g0255(.A(INSTQUEUE_REG_1__0__SCAN_IN), .Y(n1259));
  NOR2X1  g0256(.A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n1260));
  NAND3X1 g0257(.A(n1260), .B(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C(n1245), .Y(n1261));
  NOR3X1  g0258(.A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Y(n1262));
  NAND2X1 g0259(.A(n1262), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n1263));
  OAI22X1 g0260(.A0(n1261), .A1(n1259), .B0(n1258), .B1(n1263), .Y(n1264));
  NAND2X1 g0261(.A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Y(n1265));
  NOR3X1  g0262(.A(n1265), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C(n1222), .Y(n1266));
  NAND2X1 g0263(.A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n1267));
  NOR2X1  g0264(.A(n1267), .B(n1252), .Y(n1268));
  AOI22X1 g0265(.A0(n1266), .A1(INSTQUEUE_REG_13__0__SCAN_IN), .B0(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n1268), .Y(n1269));
  NOR3X1  g0266(.A(n1265), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n1270));
  NOR3X1  g0267(.A(n1267), .B(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Y(n1271));
  AOI22X1 g0268(.A0(n1270), .A1(INSTQUEUE_REG_5__0__SCAN_IN), .B0(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n1271), .Y(n1272));
  NOR3X1  g0269(.A(n1252), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n1273));
  NAND2X1 g0270(.A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n1274));
  NOR3X1  g0271(.A(n1274), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Y(n1275));
  AOI22X1 g0272(.A0(n1273), .A1(INSTQUEUE_REG_3__0__SCAN_IN), .B0(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n1275), .Y(n1276));
  NAND2X1 g0273(.A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Y(n1277));
  NOR3X1  g0274(.A(n1277), .B(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n1278));
  NOR3X1  g0275(.A(n1277), .B(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C(n1222), .Y(n1279));
  AOI22X1 g0276(.A0(n1278), .A1(INSTQUEUE_REG_6__0__SCAN_IN), .B0(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n1279), .Y(n1280));
  NAND4X1 g0277(.A(n1276), .B(n1272), .C(n1269), .D(n1280), .Y(n1281));
  NOR4X1  g0278(.A(n1264), .B(n1257), .C(n1248), .D(n1281), .Y(n1282));
  INVX1   g0279(.A(INSTQUEUE_REG_0__4__SCAN_IN), .Y(n1283));
  NAND2X1 g0280(.A(n1262), .B(n1222), .Y(n1284));
  NOR2X1  g0281(.A(n1284), .B(n1283), .Y(n1285));
  NAND4X1 g0282(.A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(n1245), .C(INSTQUEUE_REG_1__4__SCAN_IN), .D(n1260), .Y(n1286));
  NAND3X1 g0283(.A(n1262), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C(INSTQUEUE_REG_8__4__SCAN_IN), .Y(n1287));
  INVX1   g0284(.A(INSTQUEUE_REG_14__4__SCAN_IN), .Y(n1288));
  NOR4X1  g0285(.A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(n1222), .C(n1288), .D(n1277), .Y(n1289));
  NAND3X1 g0286(.A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(INSTQUEUE_REG_15__4__SCAN_IN), .Y(n1290));
  NOR2X1  g0287(.A(n1290), .B(n1274), .Y(n1291));
  NOR2X1  g0288(.A(n1291), .B(n1289), .Y(n1292));
  NAND3X1 g0289(.A(n1292), .B(n1287), .C(n1286), .Y(n1293));
  NAND3X1 g0290(.A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n1222), .C(INSTQUEUE_REG_7__4__SCAN_IN), .Y(n1294));
  NAND2X1 g0291(.A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(INSTQUEUE_REG_2__4__SCAN_IN), .Y(n1295));
  NOR4X1  g0292(.A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .D(n1295), .Y(n1296));
  NAND3X1 g0293(.A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(INSTQUEUE_REG_5__4__SCAN_IN), .Y(n1297));
  NOR3X1  g0294(.A(n1297), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n1298));
  NOR2X1  g0295(.A(n1298), .B(n1296), .Y(n1299));
  OAI21X1 g0296(.A0(n1294), .A1(n1265), .B0(n1299), .Y(n1300));
  NAND3X1 g0297(.A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(INSTQUEUE_REG_6__4__SCAN_IN), .Y(n1301));
  NOR3X1  g0298(.A(n1301), .B(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n1302));
  INVX1   g0299(.A(INSTQUEUE_REG_13__4__SCAN_IN), .Y(n1303));
  NOR4X1  g0300(.A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n1222), .C(n1303), .D(n1265), .Y(n1304));
  NOR2X1  g0301(.A(n1304), .B(n1302), .Y(n1305));
  NAND4X1 g0302(.A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n1222), .C(INSTQUEUE_REG_4__4__SCAN_IN), .D(n1250), .Y(n1306));
  NAND4X1 g0303(.A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C(INSTQUEUE_REG_12__4__SCAN_IN), .D(n1250), .Y(n1307));
  INVX1   g0304(.A(INSTQUEUE_REG_11__4__SCAN_IN), .Y(n1308));
  NOR4X1  g0305(.A(n1245), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(n1308), .D(n1274), .Y(n1309));
  NAND3X1 g0306(.A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C(INSTQUEUE_REG_3__4__SCAN_IN), .Y(n1310));
  NOR3X1  g0307(.A(n1310), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n1311));
  NAND3X1 g0308(.A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C(INSTQUEUE_REG_10__4__SCAN_IN), .Y(n1312));
  NOR3X1  g0309(.A(n1312), .B(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Y(n1313));
  NAND3X1 g0310(.A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C(INSTQUEUE_REG_9__4__SCAN_IN), .Y(n1314));
  NOR3X1  g0311(.A(n1314), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Y(n1315));
  NOR4X1  g0312(.A(n1313), .B(n1311), .C(n1309), .D(n1315), .Y(n1316));
  NAND4X1 g0313(.A(n1307), .B(n1306), .C(n1305), .D(n1316), .Y(n1317));
  NOR4X1  g0314(.A(n1300), .B(n1293), .C(n1285), .D(n1317), .Y(n1318));
  NOR3X1  g0315(.A(n1318), .B(n1282), .C(n1217), .Y(n1319));
  INVX1   g0316(.A(n1319), .Y(n1320));
  NOR2X1  g0317(.A(n1320), .B(n1241), .Y(n1321));
  INVX1   g0318(.A(n1321), .Y(n1322));
  NOR4X1  g0319(.A(n1245), .B(n1226), .C(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .D(n1231), .Y(n1323));
  INVX1   g0320(.A(INSTQUEUE_REG_2__1__SCAN_IN), .Y(n1324));
  INVX1   g0321(.A(INSTQUEUE_REG_0__1__SCAN_IN), .Y(n1325));
  NAND3X1 g0322(.A(n1260), .B(n1231), .C(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Y(n1326));
  OAI22X1 g0323(.A0(n1284), .A1(n1325), .B0(n1324), .B1(n1326), .Y(n1327));
  AOI21X1 g0324(.A0(n1323), .A1(INSTQUEUE_REG_7__1__SCAN_IN), .B0(n1327), .Y(n1328));
  NOR4X1  g0325(.A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n1226), .C(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .D(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n1329));
  INVX1   g0326(.A(INSTQUEUE_REG_11__1__SCAN_IN), .Y(n1330));
  INVX1   g0327(.A(INSTQUEUE_REG_10__1__SCAN_IN), .Y(n1331));
  NAND4X1 g0328(.A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n1226), .C(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .D(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n1332));
  NOR2X1  g0329(.A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Y(n1333));
  NAND3X1 g0330(.A(n1333), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n1334));
  OAI22X1 g0331(.A0(n1332), .A1(n1330), .B0(n1331), .B1(n1334), .Y(n1335));
  AOI21X1 g0332(.A0(n1329), .A1(INSTQUEUE_REG_4__1__SCAN_IN), .B0(n1335), .Y(n1336));
  NOR4X1  g0333(.A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .D(n1231), .Y(n1337));
  NOR4X1  g0334(.A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(n1222), .D(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n1338));
  AOI22X1 g0335(.A0(n1337), .A1(INSTQUEUE_REG_1__1__SCAN_IN), .B0(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n1338), .Y(n1339));
  INVX1   g0336(.A(INSTQUEUE_REG_15__1__SCAN_IN), .Y(n1340));
  INVX1   g0337(.A(INSTQUEUE_REG_13__1__SCAN_IN), .Y(n1341));
  NAND4X1 g0338(.A(n1245), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .D(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n1342));
  NAND4X1 g0339(.A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .D(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n1343));
  OAI22X1 g0340(.A0(n1342), .A1(n1341), .B0(n1340), .B1(n1343), .Y(n1344));
  INVX1   g0341(.A(INSTQUEUE_REG_12__1__SCAN_IN), .Y(n1345));
  INVX1   g0342(.A(INSTQUEUE_REG_5__1__SCAN_IN), .Y(n1346));
  NAND4X1 g0343(.A(n1245), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(n1222), .D(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n1347));
  NAND3X1 g0344(.A(n1250), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n1348));
  OAI22X1 g0345(.A0(n1347), .A1(n1346), .B0(n1345), .B1(n1348), .Y(n1349));
  INVX1   g0346(.A(INSTQUEUE_REG_9__1__SCAN_IN), .Y(n1350));
  INVX1   g0347(.A(INSTQUEUE_REG_3__1__SCAN_IN), .Y(n1351));
  NAND3X1 g0348(.A(n1260), .B(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Y(n1352));
  NOR2X1  g0349(.A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Y(n1353));
  NAND3X1 g0350(.A(n1353), .B(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n1354));
  OAI22X1 g0351(.A0(n1352), .A1(n1351), .B0(n1350), .B1(n1354), .Y(n1355));
  INVX1   g0352(.A(INSTQUEUE_REG_14__1__SCAN_IN), .Y(n1356));
  INVX1   g0353(.A(INSTQUEUE_REG_6__1__SCAN_IN), .Y(n1357));
  NAND4X1 g0354(.A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(n1222), .D(n1231), .Y(n1358));
  NAND4X1 g0355(.A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .D(n1231), .Y(n1359));
  OAI22X1 g0356(.A0(n1358), .A1(n1357), .B0(n1356), .B1(n1359), .Y(n1360));
  NOR4X1  g0357(.A(n1355), .B(n1349), .C(n1344), .D(n1360), .Y(n1361));
  NAND4X1 g0358(.A(n1339), .B(n1336), .C(n1328), .D(n1361), .Y(n1362));
  NAND4X1 g0359(.A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C(INSTQUEUE_REG_12__5__SCAN_IN), .D(n1250), .Y(n1363));
  NAND3X1 g0360(.A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(INSTQUEUE_REG_15__5__SCAN_IN), .Y(n1364));
  OAI21X1 g0361(.A0(n1364), .A1(n1274), .B0(n1363), .Y(n1365));
  NAND2X1 g0362(.A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(n1245), .Y(n1366));
  NAND3X1 g0363(.A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n1226), .C(INSTQUEUE_REG_11__5__SCAN_IN), .Y(n1367));
  NAND3X1 g0364(.A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C(INSTQUEUE_REG_13__5__SCAN_IN), .Y(n1368));
  OAI22X1 g0365(.A0(n1367), .A1(n1274), .B0(n1366), .B1(n1368), .Y(n1369));
  NAND2X1 g0366(.A(n1226), .B(n1222), .Y(n1370));
  NAND4X1 g0367(.A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C(INSTQUEUE_REG_10__5__SCAN_IN), .D(n1333), .Y(n1371));
  NAND3X1 g0368(.A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C(INSTQUEUE_REG_3__5__SCAN_IN), .Y(n1372));
  OAI21X1 g0369(.A0(n1372), .A1(n1370), .B0(n1371), .Y(n1373));
  NAND3X1 g0370(.A(n1231), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(INSTQUEUE_REG_14__5__SCAN_IN), .Y(n1374));
  NAND4X1 g0371(.A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C(INSTQUEUE_REG_9__5__SCAN_IN), .D(n1353), .Y(n1375));
  OAI21X1 g0372(.A0(n1374), .A1(n1254), .B0(n1375), .Y(n1376));
  NOR4X1  g0373(.A(n1373), .B(n1369), .C(n1365), .D(n1376), .Y(n1377));
  NAND2X1 g0374(.A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(INSTQUEUE_REG_2__5__SCAN_IN), .Y(n1378));
  NOR4X1  g0375(.A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .D(n1378), .Y(n1379));
  NAND4X1 g0376(.A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(n1245), .C(INSTQUEUE_REG_1__5__SCAN_IN), .D(n1260), .Y(n1380));
  NAND4X1 g0377(.A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n1222), .C(INSTQUEUE_REG_4__5__SCAN_IN), .D(n1250), .Y(n1381));
  NAND2X1 g0378(.A(n1381), .B(n1380), .Y(n1382));
  NOR2X1  g0379(.A(n1382), .B(n1379), .Y(n1383));
  NAND2X1 g0380(.A(n1244), .B(INSTQUEUE_REG_0__5__SCAN_IN), .Y(n1384));
  INVX1   g0381(.A(INSTQUEUE_REG_7__5__SCAN_IN), .Y(n1385));
  NOR4X1  g0382(.A(n1245), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C(n1385), .D(n1265), .Y(n1386));
  NAND3X1 g0383(.A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(INSTQUEUE_REG_6__5__SCAN_IN), .Y(n1387));
  NOR3X1  g0384(.A(n1387), .B(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n1388));
  NAND3X1 g0385(.A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(INSTQUEUE_REG_5__5__SCAN_IN), .Y(n1389));
  NOR3X1  g0386(.A(n1389), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n1390));
  NAND2X1 g0387(.A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(INSTQUEUE_REG_8__5__SCAN_IN), .Y(n1391));
  NOR4X1  g0388(.A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .D(n1391), .Y(n1392));
  NOR4X1  g0389(.A(n1390), .B(n1388), .C(n1386), .D(n1392), .Y(n1393));
  NAND4X1 g0390(.A(n1384), .B(n1383), .C(n1377), .D(n1393), .Y(n1394));
  NOR3X1  g0391(.A(n1394), .B(n1362), .C(n1217), .Y(n1395));
  NAND2X1 g0392(.A(n1287), .B(n1286), .Y(n1396));
  NOR4X1  g0393(.A(n1289), .B(n1396), .C(n1285), .D(n1291), .Y(n1397));
  INVX1   g0394(.A(INSTQUEUE_REG_7__4__SCAN_IN), .Y(n1398));
  NOR4X1  g0395(.A(n1245), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C(n1398), .D(n1265), .Y(n1399));
  NOR3X1  g0396(.A(n1298), .B(n1296), .C(n1399), .Y(n1400));
  NAND2X1 g0397(.A(n1307), .B(n1306), .Y(n1401));
  NOR3X1  g0398(.A(n1401), .B(n1304), .C(n1302), .Y(n1402));
  NAND4X1 g0399(.A(n1402), .B(n1400), .C(n1397), .D(n1316), .Y(n1403));
  NOR2X1  g0400(.A(n1231), .B(n1222), .Y(n1404));
  NAND4X1 g0401(.A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(INSTQUEUE_REG_15__5__SCAN_IN), .D(n1404), .Y(n1405));
  INVX1   g0402(.A(INSTQUEUE_REG_11__5__SCAN_IN), .Y(n1406));
  NOR4X1  g0403(.A(n1245), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(n1406), .D(n1274), .Y(n1407));
  NOR3X1  g0404(.A(n1368), .B(n1231), .C(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Y(n1408));
  NOR2X1  g0405(.A(n1408), .B(n1407), .Y(n1409));
  NAND3X1 g0406(.A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C(INSTQUEUE_REG_10__5__SCAN_IN), .Y(n1410));
  NOR3X1  g0407(.A(n1410), .B(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Y(n1411));
  NOR3X1  g0408(.A(n1372), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n1412));
  INVX1   g0409(.A(INSTQUEUE_REG_14__5__SCAN_IN), .Y(n1413));
  NOR4X1  g0410(.A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(n1226), .C(n1413), .D(n1254), .Y(n1414));
  NAND3X1 g0411(.A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C(INSTQUEUE_REG_9__5__SCAN_IN), .Y(n1415));
  NOR3X1  g0412(.A(n1415), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Y(n1416));
  NOR4X1  g0413(.A(n1414), .B(n1412), .C(n1411), .D(n1416), .Y(n1417));
  NAND4X1 g0414(.A(n1409), .B(n1405), .C(n1363), .D(n1417), .Y(n1418));
  NAND4X1 g0415(.A(n1231), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C(INSTQUEUE_REG_2__5__SCAN_IN), .D(n1260), .Y(n1419));
  NAND3X1 g0416(.A(n1381), .B(n1380), .C(n1419), .Y(n1420));
  NAND2X1 g0417(.A(n1393), .B(n1384), .Y(n1421));
  NOR3X1  g0418(.A(n1421), .B(n1420), .C(n1418), .Y(n1422));
  NOR3X1  g0419(.A(n1422), .B(n1403), .C(n1217), .Y(n1423));
  INVX1   g0420(.A(n1423), .Y(n1424));
  INVX1   g0421(.A(INSTQUEUE_REG_2__0__SCAN_IN), .Y(n1425));
  INVX1   g0422(.A(INSTQUEUE_REG_0__0__SCAN_IN), .Y(n1426));
  OAI22X1 g0423(.A0(n1284), .A1(n1426), .B0(n1425), .B1(n1326), .Y(n1427));
  AOI21X1 g0424(.A0(n1323), .A1(INSTQUEUE_REG_7__0__SCAN_IN), .B0(n1427), .Y(n1428));
  INVX1   g0425(.A(INSTQUEUE_REG_11__0__SCAN_IN), .Y(n1429));
  INVX1   g0426(.A(INSTQUEUE_REG_10__0__SCAN_IN), .Y(n1430));
  OAI22X1 g0427(.A0(n1332), .A1(n1429), .B0(n1430), .B1(n1334), .Y(n1431));
  AOI21X1 g0428(.A0(n1329), .A1(INSTQUEUE_REG_4__0__SCAN_IN), .B0(n1431), .Y(n1432));
  AOI22X1 g0429(.A0(n1337), .A1(INSTQUEUE_REG_1__0__SCAN_IN), .B0(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n1338), .Y(n1433));
  INVX1   g0430(.A(INSTQUEUE_REG_15__0__SCAN_IN), .Y(n1434));
  INVX1   g0431(.A(INSTQUEUE_REG_13__0__SCAN_IN), .Y(n1435));
  OAI22X1 g0432(.A0(n1342), .A1(n1435), .B0(n1434), .B1(n1343), .Y(n1436));
  INVX1   g0433(.A(INSTQUEUE_REG_12__0__SCAN_IN), .Y(n1437));
  INVX1   g0434(.A(INSTQUEUE_REG_5__0__SCAN_IN), .Y(n1438));
  OAI22X1 g0435(.A0(n1347), .A1(n1438), .B0(n1437), .B1(n1348), .Y(n1439));
  INVX1   g0436(.A(INSTQUEUE_REG_9__0__SCAN_IN), .Y(n1440));
  INVX1   g0437(.A(INSTQUEUE_REG_3__0__SCAN_IN), .Y(n1441));
  OAI22X1 g0438(.A0(n1352), .A1(n1441), .B0(n1440), .B1(n1354), .Y(n1442));
  INVX1   g0439(.A(INSTQUEUE_REG_14__0__SCAN_IN), .Y(n1443));
  INVX1   g0440(.A(INSTQUEUE_REG_6__0__SCAN_IN), .Y(n1444));
  OAI22X1 g0441(.A0(n1358), .A1(n1444), .B0(n1443), .B1(n1359), .Y(n1445));
  NOR4X1  g0442(.A(n1442), .B(n1439), .C(n1436), .D(n1445), .Y(n1446));
  NAND4X1 g0443(.A(n1433), .B(n1432), .C(n1428), .D(n1446), .Y(n1447));
  NAND2X1 g0444(.A(n1362), .B(n1447), .Y(n1448));
  NOR4X1  g0445(.A(n1362), .B(n1282), .C(n1217), .D(n1422), .Y(n1449));
  INVX1   g0446(.A(INSTQUEUE_REG_7__1__SCAN_IN), .Y(n1450));
  AOI22X1 g0447(.A0(n1244), .A1(INSTQUEUE_REG_0__1__SCAN_IN), .B0(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n1246), .Y(n1451));
  OAI21X1 g0448(.A0(n1243), .A1(n1450), .B0(n1451), .Y(n1452));
  INVX1   g0449(.A(INSTQUEUE_REG_4__1__SCAN_IN), .Y(n1453));
  AOI22X1 g0450(.A0(n1253), .A1(INSTQUEUE_REG_11__1__SCAN_IN), .B0(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n1255), .Y(n1454));
  OAI21X1 g0451(.A0(n1251), .A1(n1453), .B0(n1454), .Y(n1455));
  INVX1   g0452(.A(INSTQUEUE_REG_8__1__SCAN_IN), .Y(n1456));
  INVX1   g0453(.A(INSTQUEUE_REG_1__1__SCAN_IN), .Y(n1457));
  OAI22X1 g0454(.A0(n1261), .A1(n1457), .B0(n1456), .B1(n1263), .Y(n1458));
  AOI22X1 g0455(.A0(n1266), .A1(INSTQUEUE_REG_13__1__SCAN_IN), .B0(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n1268), .Y(n1459));
  AOI22X1 g0456(.A0(n1270), .A1(INSTQUEUE_REG_5__1__SCAN_IN), .B0(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n1271), .Y(n1460));
  AOI22X1 g0457(.A0(n1273), .A1(INSTQUEUE_REG_3__1__SCAN_IN), .B0(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n1275), .Y(n1461));
  AOI22X1 g0458(.A0(n1278), .A1(INSTQUEUE_REG_6__1__SCAN_IN), .B0(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n1279), .Y(n1462));
  NAND4X1 g0459(.A(n1461), .B(n1460), .C(n1459), .D(n1462), .Y(n1463));
  NOR4X1  g0460(.A(n1458), .B(n1455), .C(n1452), .D(n1463), .Y(n1464));
  NOR3X1  g0461(.A(n1464), .B(n1447), .C(n1217), .Y(n1465));
  NOR3X1  g0462(.A(n1394), .B(n1464), .C(n1217), .Y(n1466));
  NOR3X1  g0463(.A(n1362), .B(n1447), .C(n1217), .Y(n1467));
  NOR4X1  g0464(.A(n1466), .B(n1465), .C(n1449), .D(n1467), .Y(n1468));
  OAI21X1 g0465(.A0(n1448), .A1(n1424), .B0(n1468), .Y(n1469));
  OAI22X1 g0466(.A0(n1395), .A1(n1469), .B0(n1240), .B1(n1219), .Y(n1470));
  INVX1   g0467(.A(n1470), .Y(n1471));
  NOR2X1  g0468(.A(n1422), .B(n1464), .Y(n1472));
  INVX1   g0469(.A(n1472), .Y(n1473));
  NOR2X1  g0470(.A(n1473), .B(n1320), .Y(n1474));
  NOR2X1  g0471(.A(n1422), .B(n1217), .Y(n1475));
  NOR2X1  g0472(.A(n1447), .B(n1217), .Y(n1476));
  OAI21X1 g0473(.A0(n1476), .A1(n1475), .B0(n1464), .Y(n1477));
  XOR2X1  g0474(.A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n1231), .Y(n1478));
  INVX1   g0475(.A(n1478), .Y(n1479));
  NAND4X1 g0476(.A(n1403), .B(n1447), .C(STATE2_REG_0__SCAN_IN), .D(n1479), .Y(n1480));
  AOI22X1 g0477(.A0(n1447), .A1(n1423), .B0(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(n1217), .Y(n1481));
  NAND3X1 g0478(.A(n1481), .B(n1480), .C(n1477), .Y(n1482));
  INVX1   g0479(.A(n1395), .Y(n1483));
  AOI21X1 g0480(.A0(n1403), .A1(n1447), .B0(n1217), .Y(n1484));
  OAI21X1 g0481(.A0(n1478), .A1(n1483), .B0(n1484), .Y(n1485));
  AOI21X1 g0482(.A0(n1479), .A1(n1469), .B0(n1485), .Y(n1486));
  OAI21X1 g0483(.A0(n1486), .A1(n1482), .B0(n1474), .Y(n1487));
  XOR2X1  g0484(.A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n1245), .Y(n1488));
  XOR2X1  g0485(.A(n1488), .B(n1232), .Y(n1489));
  INVX1   g0486(.A(n1489), .Y(n1490));
  OAI21X1 g0487(.A0(n1489), .A1(n1483), .B0(STATE2_REG_0__SCAN_IN), .Y(n1491));
  AOI21X1 g0488(.A0(n1490), .A1(n1469), .B0(n1491), .Y(n1492));
  NAND3X1 g0489(.A(n1362), .B(n1282), .C(STATE2_REG_0__SCAN_IN), .Y(n1493));
  NAND4X1 g0490(.A(n1403), .B(n1447), .C(STATE2_REG_0__SCAN_IN), .D(n1490), .Y(n1494));
  NAND3X1 g0491(.A(n1362), .B(n1318), .C(STATE2_REG_0__SCAN_IN), .Y(n1495));
  NOR4X1  g0492(.A(n1420), .B(n1418), .C(n1217), .D(n1421), .Y(n1496));
  AOI21X1 g0493(.A0(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A1(n1217), .B0(n1496), .Y(n1497));
  NAND4X1 g0494(.A(n1495), .B(n1494), .C(n1493), .D(n1497), .Y(n1498));
  AOI22X1 g0495(.A0(n1492), .A1(n1498), .B0(n1486), .B1(n1482), .Y(n1499));
  XOR2X1  g0496(.A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n1226), .Y(n1500));
  XOR2X1  g0497(.A(n1500), .B(n1234), .Y(n1501));
  INVX1   g0498(.A(n1501), .Y(n1502));
  AOI22X1 g0499(.A0(n1319), .A1(n1502), .B0(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(n1217), .Y(n1503));
  NAND2X1 g0500(.A(n1503), .B(n1477), .Y(n1504));
  OAI21X1 g0501(.A0(n1501), .A1(n1483), .B0(n1484), .Y(n1505));
  AOI21X1 g0502(.A0(n1502), .A1(n1469), .B0(n1505), .Y(n1506));
  OAI22X1 g0503(.A0(n1504), .A1(n1506), .B0(n1498), .B1(n1492), .Y(n1507));
  AOI21X1 g0504(.A0(n1499), .A1(n1487), .B0(n1507), .Y(n1508));
  NAND2X1 g0505(.A(n1506), .B(n1504), .Y(n1509));
  INVX1   g0506(.A(n1469), .Y(n1510));
  XOR2X1  g0507(.A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n1222), .Y(n1511));
  XOR2X1  g0508(.A(n1511), .B(n1236), .Y(n1512));
  INVX1   g0509(.A(n1512), .Y(n1513));
  AOI21X1 g0510(.A0(n1513), .A1(n1395), .B0(n1217), .Y(n1514));
  OAI21X1 g0511(.A0(n1512), .A1(n1510), .B0(n1514), .Y(n1515));
  AOI22X1 g0512(.A0(n1319), .A1(n1513), .B0(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(n1217), .Y(n1516));
  OAI21X1 g0513(.A0(n1516), .A1(n1515), .B0(n1509), .Y(n1517));
  NOR2X1  g0514(.A(n1237), .B(n1221), .Y(n1518));
  XOR2X1  g0515(.A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B(n1218), .Y(n1519));
  XOR2X1  g0516(.A(n1519), .B(n1518), .Y(n1520));
  INVX1   g0517(.A(n1520), .Y(n1521));
  AOI22X1 g0518(.A0(n1319), .A1(n1521), .B0(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B1(n1217), .Y(n1522));
  AOI21X1 g0519(.A0(n1510), .A1(n1483), .B0(n1520), .Y(n1523));
  AOI22X1 g0520(.A0(n1522), .A1(n1523), .B0(n1516), .B1(n1515), .Y(n1524));
  OAI21X1 g0521(.A0(n1517), .A1(n1508), .B0(n1524), .Y(n1525));
  INVX1   g0522(.A(n1522), .Y(n1526));
  INVX1   g0523(.A(n1523), .Y(n1527));
  AOI22X1 g0524(.A0(n1526), .A1(n1527), .B0(n1470), .B1(n1321), .Y(n1528));
  AOI22X1 g0525(.A0(n1525), .A1(n1528), .B0(n1471), .B1(n1322), .Y(n1529));
  NOR2X1  g0526(.A(n1529), .B(n1470), .Y(n1530));
  AOI21X1 g0527(.A0(n1470), .A1(STATE2_REG_0__SCAN_IN), .B0(n1530), .Y(n1531));
  NAND2X1 g0528(.A(n1527), .B(n1526), .Y(n1532));
  NAND4X1 g0529(.A(n1525), .B(n1470), .C(n1322), .D(n1532), .Y(n1533));
  OAI21X1 g0530(.A0(n1531), .A1(n1322), .B0(n1533), .Y(n1536));
  NAND2X1 g0531(.A(n1244), .B(INSTQUEUE_REG_0__6__SCAN_IN), .Y(n1537));
  NAND3X1 g0532(.A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C(INSTQUEUE_REG_3__6__SCAN_IN), .Y(n1538));
  NOR3X1  g0533(.A(n1538), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n1539));
  NAND3X1 g0534(.A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C(INSTQUEUE_REG_9__6__SCAN_IN), .Y(n1540));
  NOR3X1  g0535(.A(n1540), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Y(n1541));
  NOR2X1  g0536(.A(n1541), .B(n1539), .Y(n1542));
  NOR2X1  g0537(.A(n1226), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n1543));
  NOR2X1  g0538(.A(n1231), .B(n1245), .Y(n1544));
  NAND3X1 g0539(.A(n1544), .B(n1543), .C(INSTQUEUE_REG_7__6__SCAN_IN), .Y(n1545));
  NAND3X1 g0540(.A(n1262), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C(INSTQUEUE_REG_8__6__SCAN_IN), .Y(n1546));
  NAND4X1 g0541(.A(n1545), .B(n1542), .C(n1537), .D(n1546), .Y(n1547));
  NAND3X1 g0542(.A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(n1245), .C(INSTQUEUE_REG_1__6__SCAN_IN), .Y(n1548));
  NOR2X1  g0543(.A(n1548), .B(n1370), .Y(n1549));
  NAND4X1 g0544(.A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n1222), .C(INSTQUEUE_REG_4__6__SCAN_IN), .D(n1250), .Y(n1550));
  NAND4X1 g0545(.A(n1231), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C(INSTQUEUE_REG_2__6__SCAN_IN), .D(n1260), .Y(n1551));
  NAND2X1 g0546(.A(n1551), .B(n1550), .Y(n1552));
  NAND4X1 g0547(.A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(n1245), .C(INSTQUEUE_REG_5__6__SCAN_IN), .D(n1543), .Y(n1553));
  NAND4X1 g0548(.A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C(INSTQUEUE_REG_15__6__SCAN_IN), .D(n1544), .Y(n1554));
  INVX1   g0549(.A(INSTQUEUE_REG_6__6__SCAN_IN), .Y(n1555));
  NOR3X1  g0550(.A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(n1245), .C(n1555), .Y(n1556));
  AOI22X1 g0551(.A0(n1271), .A1(INSTQUEUE_REG_12__6__SCAN_IN), .B0(n1543), .B1(n1556), .Y(n1557));
  NAND3X1 g0552(.A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C(INSTQUEUE_REG_10__6__SCAN_IN), .Y(n1558));
  NOR3X1  g0553(.A(n1558), .B(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Y(n1559));
  INVX1   g0554(.A(INSTQUEUE_REG_11__6__SCAN_IN), .Y(n1560));
  NOR4X1  g0555(.A(n1245), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(n1560), .D(n1274), .Y(n1561));
  INVX1   g0556(.A(INSTQUEUE_REG_14__6__SCAN_IN), .Y(n1562));
  NOR4X1  g0557(.A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(n1245), .C(n1562), .D(n1267), .Y(n1563));
  INVX1   g0558(.A(INSTQUEUE_REG_13__6__SCAN_IN), .Y(n1564));
  NOR4X1  g0559(.A(n1231), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C(n1564), .D(n1267), .Y(n1565));
  NOR4X1  g0560(.A(n1563), .B(n1561), .C(n1559), .D(n1565), .Y(n1566));
  NAND4X1 g0561(.A(n1557), .B(n1554), .C(n1553), .D(n1566), .Y(n1567));
  NOR4X1  g0562(.A(n1552), .B(n1549), .C(n1547), .D(n1567), .Y(n1568));
  NAND2X1 g0563(.A(n1568), .B(n1422), .Y(n1569));
  INVX1   g0564(.A(INSTQUEUE_REG_2__3__SCAN_IN), .Y(n1570));
  INVX1   g0565(.A(INSTQUEUE_REG_0__3__SCAN_IN), .Y(n1571));
  OAI22X1 g0566(.A0(n1284), .A1(n1571), .B0(n1570), .B1(n1326), .Y(n1572));
  AOI21X1 g0567(.A0(n1323), .A1(INSTQUEUE_REG_7__3__SCAN_IN), .B0(n1572), .Y(n1573));
  INVX1   g0568(.A(INSTQUEUE_REG_11__3__SCAN_IN), .Y(n1574));
  INVX1   g0569(.A(INSTQUEUE_REG_10__3__SCAN_IN), .Y(n1575));
  OAI22X1 g0570(.A0(n1332), .A1(n1574), .B0(n1575), .B1(n1334), .Y(n1576));
  AOI21X1 g0571(.A0(n1329), .A1(INSTQUEUE_REG_4__3__SCAN_IN), .B0(n1576), .Y(n1577));
  AOI22X1 g0572(.A0(n1337), .A1(INSTQUEUE_REG_1__3__SCAN_IN), .B0(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n1338), .Y(n1578));
  INVX1   g0573(.A(INSTQUEUE_REG_15__3__SCAN_IN), .Y(n1579));
  INVX1   g0574(.A(INSTQUEUE_REG_13__3__SCAN_IN), .Y(n1580));
  OAI22X1 g0575(.A0(n1342), .A1(n1580), .B0(n1579), .B1(n1343), .Y(n1581));
  INVX1   g0576(.A(INSTQUEUE_REG_12__3__SCAN_IN), .Y(n1582));
  INVX1   g0577(.A(INSTQUEUE_REG_5__3__SCAN_IN), .Y(n1583));
  OAI22X1 g0578(.A0(n1347), .A1(n1583), .B0(n1582), .B1(n1348), .Y(n1584));
  INVX1   g0579(.A(INSTQUEUE_REG_9__3__SCAN_IN), .Y(n1585));
  INVX1   g0580(.A(INSTQUEUE_REG_3__3__SCAN_IN), .Y(n1586));
  OAI22X1 g0581(.A0(n1352), .A1(n1586), .B0(n1585), .B1(n1354), .Y(n1587));
  INVX1   g0582(.A(INSTQUEUE_REG_14__3__SCAN_IN), .Y(n1588));
  INVX1   g0583(.A(INSTQUEUE_REG_6__3__SCAN_IN), .Y(n1589));
  OAI22X1 g0584(.A0(n1358), .A1(n1589), .B0(n1588), .B1(n1359), .Y(n1590));
  NOR4X1  g0585(.A(n1587), .B(n1584), .C(n1581), .D(n1590), .Y(n1591));
  NAND4X1 g0586(.A(n1578), .B(n1577), .C(n1573), .D(n1591), .Y(n1592));
  INVX1   g0587(.A(INSTQUEUE_REG_2__7__SCAN_IN), .Y(n1593));
  INVX1   g0588(.A(INSTQUEUE_REG_0__7__SCAN_IN), .Y(n1594));
  OAI22X1 g0589(.A0(n1284), .A1(n1594), .B0(n1593), .B1(n1326), .Y(n1595));
  AOI21X1 g0590(.A0(n1323), .A1(INSTQUEUE_REG_7__7__SCAN_IN), .B0(n1595), .Y(n1596));
  INVX1   g0591(.A(INSTQUEUE_REG_11__7__SCAN_IN), .Y(n1597));
  INVX1   g0592(.A(INSTQUEUE_REG_10__7__SCAN_IN), .Y(n1598));
  OAI22X1 g0593(.A0(n1332), .A1(n1597), .B0(n1598), .B1(n1334), .Y(n1599));
  AOI21X1 g0594(.A0(n1329), .A1(INSTQUEUE_REG_4__7__SCAN_IN), .B0(n1599), .Y(n1600));
  AOI22X1 g0595(.A0(n1337), .A1(INSTQUEUE_REG_1__7__SCAN_IN), .B0(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n1338), .Y(n1601));
  INVX1   g0596(.A(INSTQUEUE_REG_15__7__SCAN_IN), .Y(n1602));
  INVX1   g0597(.A(INSTQUEUE_REG_13__7__SCAN_IN), .Y(n1603));
  OAI22X1 g0598(.A0(n1342), .A1(n1603), .B0(n1602), .B1(n1343), .Y(n1604));
  INVX1   g0599(.A(INSTQUEUE_REG_12__7__SCAN_IN), .Y(n1605));
  INVX1   g0600(.A(INSTQUEUE_REG_5__7__SCAN_IN), .Y(n1606));
  OAI22X1 g0601(.A0(n1347), .A1(n1606), .B0(n1605), .B1(n1348), .Y(n1607));
  INVX1   g0602(.A(INSTQUEUE_REG_9__7__SCAN_IN), .Y(n1608));
  INVX1   g0603(.A(INSTQUEUE_REG_3__7__SCAN_IN), .Y(n1609));
  OAI22X1 g0604(.A0(n1352), .A1(n1609), .B0(n1608), .B1(n1354), .Y(n1610));
  INVX1   g0605(.A(INSTQUEUE_REG_14__7__SCAN_IN), .Y(n1611));
  INVX1   g0606(.A(INSTQUEUE_REG_6__7__SCAN_IN), .Y(n1612));
  OAI22X1 g0607(.A0(n1358), .A1(n1612), .B0(n1611), .B1(n1359), .Y(n1613));
  NOR4X1  g0608(.A(n1610), .B(n1607), .C(n1604), .D(n1613), .Y(n1614));
  NAND4X1 g0609(.A(n1601), .B(n1600), .C(n1596), .D(n1614), .Y(n1615));
  NAND2X1 g0610(.A(n1615), .B(n1592), .Y(n1616));
  INVX1   g0611(.A(INSTQUEUE_REG_2__2__SCAN_IN), .Y(n1617));
  INVX1   g0612(.A(INSTQUEUE_REG_0__2__SCAN_IN), .Y(n1618));
  OAI22X1 g0613(.A0(n1284), .A1(n1618), .B0(n1617), .B1(n1326), .Y(n1619));
  AOI21X1 g0614(.A0(n1323), .A1(INSTQUEUE_REG_7__2__SCAN_IN), .B0(n1619), .Y(n1620));
  INVX1   g0615(.A(INSTQUEUE_REG_11__2__SCAN_IN), .Y(n1621));
  INVX1   g0616(.A(INSTQUEUE_REG_10__2__SCAN_IN), .Y(n1622));
  OAI22X1 g0617(.A0(n1332), .A1(n1621), .B0(n1622), .B1(n1334), .Y(n1623));
  AOI21X1 g0618(.A0(n1329), .A1(INSTQUEUE_REG_4__2__SCAN_IN), .B0(n1623), .Y(n1624));
  AOI22X1 g0619(.A0(n1337), .A1(INSTQUEUE_REG_1__2__SCAN_IN), .B0(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n1338), .Y(n1625));
  INVX1   g0620(.A(INSTQUEUE_REG_15__2__SCAN_IN), .Y(n1626));
  INVX1   g0621(.A(INSTQUEUE_REG_13__2__SCAN_IN), .Y(n1627));
  OAI22X1 g0622(.A0(n1342), .A1(n1627), .B0(n1626), .B1(n1343), .Y(n1628));
  INVX1   g0623(.A(INSTQUEUE_REG_12__2__SCAN_IN), .Y(n1629));
  INVX1   g0624(.A(INSTQUEUE_REG_5__2__SCAN_IN), .Y(n1630));
  OAI22X1 g0625(.A0(n1347), .A1(n1630), .B0(n1629), .B1(n1348), .Y(n1631));
  INVX1   g0626(.A(INSTQUEUE_REG_9__2__SCAN_IN), .Y(n1632));
  INVX1   g0627(.A(INSTQUEUE_REG_3__2__SCAN_IN), .Y(n1633));
  OAI22X1 g0628(.A0(n1352), .A1(n1633), .B0(n1632), .B1(n1354), .Y(n1634));
  INVX1   g0629(.A(INSTQUEUE_REG_14__2__SCAN_IN), .Y(n1635));
  INVX1   g0630(.A(INSTQUEUE_REG_6__2__SCAN_IN), .Y(n1636));
  OAI22X1 g0631(.A0(n1358), .A1(n1636), .B0(n1635), .B1(n1359), .Y(n1637));
  NOR4X1  g0632(.A(n1634), .B(n1631), .C(n1628), .D(n1637), .Y(n1638));
  NAND4X1 g0633(.A(n1625), .B(n1624), .C(n1620), .D(n1638), .Y(n1639));
  NOR4X1  g0634(.A(n1616), .B(n1569), .C(n1403), .D(n1639), .Y(n1640));
  INVX1   g0635(.A(INSTQUEUE_REG_7__3__SCAN_IN), .Y(n1641));
  AOI22X1 g0636(.A0(n1244), .A1(INSTQUEUE_REG_0__3__SCAN_IN), .B0(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n1246), .Y(n1642));
  OAI21X1 g0637(.A0(n1243), .A1(n1641), .B0(n1642), .Y(n1643));
  INVX1   g0638(.A(INSTQUEUE_REG_4__3__SCAN_IN), .Y(n1644));
  AOI22X1 g0639(.A0(n1253), .A1(INSTQUEUE_REG_11__3__SCAN_IN), .B0(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n1255), .Y(n1645));
  OAI21X1 g0640(.A0(n1251), .A1(n1644), .B0(n1645), .Y(n1646));
  INVX1   g0641(.A(INSTQUEUE_REG_8__3__SCAN_IN), .Y(n1647));
  INVX1   g0642(.A(INSTQUEUE_REG_1__3__SCAN_IN), .Y(n1648));
  OAI22X1 g0643(.A0(n1261), .A1(n1648), .B0(n1647), .B1(n1263), .Y(n1649));
  AOI22X1 g0644(.A0(n1266), .A1(INSTQUEUE_REG_13__3__SCAN_IN), .B0(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n1268), .Y(n1650));
  AOI22X1 g0645(.A0(n1270), .A1(INSTQUEUE_REG_5__3__SCAN_IN), .B0(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n1271), .Y(n1651));
  AOI22X1 g0646(.A0(n1273), .A1(INSTQUEUE_REG_3__3__SCAN_IN), .B0(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n1275), .Y(n1652));
  AOI22X1 g0647(.A0(n1278), .A1(INSTQUEUE_REG_6__3__SCAN_IN), .B0(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n1279), .Y(n1653));
  NAND4X1 g0648(.A(n1652), .B(n1651), .C(n1650), .D(n1653), .Y(n1654));
  NOR4X1  g0649(.A(n1649), .B(n1646), .C(n1643), .D(n1654), .Y(n1655));
  NAND2X1 g0650(.A(n1639), .B(n1655), .Y(n1656));
  INVX1   g0651(.A(INSTQUEUE_REG_0__6__SCAN_IN), .Y(n1657));
  NOR2X1  g0652(.A(n1284), .B(n1657), .Y(n1658));
  NAND3X1 g0653(.A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n1222), .C(INSTQUEUE_REG_7__6__SCAN_IN), .Y(n1659));
  OAI21X1 g0654(.A0(n1659), .A1(n1252), .B0(n1546), .Y(n1660));
  NOR4X1  g0655(.A(n1541), .B(n1539), .C(n1658), .D(n1660), .Y(n1661));
  NOR2X1  g0656(.A(n1552), .B(n1549), .Y(n1662));
  NAND2X1 g0657(.A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n1222), .Y(n1663));
  NAND3X1 g0658(.A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(n1245), .C(INSTQUEUE_REG_5__6__SCAN_IN), .Y(n1664));
  NAND3X1 g0659(.A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C(INSTQUEUE_REG_15__6__SCAN_IN), .Y(n1665));
  OAI22X1 g0660(.A0(n1664), .A1(n1663), .B0(n1267), .B1(n1665), .Y(n1666));
  INVX1   g0661(.A(INSTQUEUE_REG_12__6__SCAN_IN), .Y(n1667));
  NAND3X1 g0662(.A(n1231), .B(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C(INSTQUEUE_REG_6__6__SCAN_IN), .Y(n1668));
  OAI22X1 g0663(.A0(n1348), .A1(n1667), .B0(n1663), .B1(n1668), .Y(n1669));
  NOR2X1  g0664(.A(n1669), .B(n1666), .Y(n1670));
  NAND4X1 g0665(.A(n1670), .B(n1662), .C(n1661), .D(n1566), .Y(n1671));
  NAND4X1 g0666(.A(n1671), .B(n1394), .C(n1318), .D(n1615), .Y(n1672));
  NOR4X1  g0667(.A(n1656), .B(n1464), .C(n1447), .D(n1672), .Y(n1673));
  XOR2X1  g0668(.A(STATE_REG_1__SCAN_IN), .B(n1112), .Y(n1674));
  NOR3X1  g0669(.A(n1674), .B(STATE_REG_0__SCAN_IN), .C(READY_N), .Y(n1675));
  OAI21X1 g0670(.A0(n1673), .A1(n1640), .B0(n1675), .Y(n1676));
  NAND4X1 g0671(.A(n1568), .B(n1394), .C(n1403), .D(n1615), .Y(n1677));
  NAND2X1 g0672(.A(n1464), .B(n1282), .Y(n1678));
  NOR4X1  g0673(.A(n1677), .B(n1639), .C(n1655), .D(n1678), .Y(n1679));
  NOR3X1  g0674(.A(n1464), .B(n1282), .C(READY_N), .Y(n1680));
  AOI21X1 g0675(.A0(n1680), .A1(n1640), .B0(n1679), .Y(n1681));
  NAND2X1 g0676(.A(n1681), .B(n1676), .Y(n1682));
  NAND3X1 g0677(.A(n1592), .B(n1362), .C(n1447), .Y(n1683));
  NOR3X1  g0678(.A(n1683), .B(n1677), .C(n1639), .Y(n1684));
  INVX1   g0679(.A(n1684), .Y(n1685));
  INVX1   g0680(.A(INSTQUEUE_REG_7__7__SCAN_IN), .Y(n1686));
  AOI22X1 g0681(.A0(n1244), .A1(INSTQUEUE_REG_0__7__SCAN_IN), .B0(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n1246), .Y(n1687));
  OAI21X1 g0682(.A0(n1243), .A1(n1686), .B0(n1687), .Y(n1688));
  INVX1   g0683(.A(INSTQUEUE_REG_4__7__SCAN_IN), .Y(n1689));
  AOI22X1 g0684(.A0(n1253), .A1(INSTQUEUE_REG_11__7__SCAN_IN), .B0(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n1255), .Y(n1690));
  OAI21X1 g0685(.A0(n1251), .A1(n1689), .B0(n1690), .Y(n1691));
  INVX1   g0686(.A(INSTQUEUE_REG_8__7__SCAN_IN), .Y(n1692));
  INVX1   g0687(.A(INSTQUEUE_REG_1__7__SCAN_IN), .Y(n1693));
  OAI22X1 g0688(.A0(n1261), .A1(n1693), .B0(n1692), .B1(n1263), .Y(n1694));
  AOI22X1 g0689(.A0(n1266), .A1(INSTQUEUE_REG_13__7__SCAN_IN), .B0(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n1268), .Y(n1695));
  AOI22X1 g0690(.A0(n1270), .A1(INSTQUEUE_REG_5__7__SCAN_IN), .B0(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n1271), .Y(n1696));
  AOI22X1 g0691(.A0(n1273), .A1(INSTQUEUE_REG_3__7__SCAN_IN), .B0(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n1275), .Y(n1697));
  AOI22X1 g0692(.A0(n1278), .A1(INSTQUEUE_REG_6__7__SCAN_IN), .B0(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n1279), .Y(n1698));
  NAND4X1 g0693(.A(n1697), .B(n1696), .C(n1695), .D(n1698), .Y(n1699));
  NOR4X1  g0694(.A(n1694), .B(n1691), .C(n1688), .D(n1699), .Y(n1700));
  AOI21X1 g0695(.A0(n1671), .A1(n1422), .B0(n1700), .Y(n1701));
  NAND3X1 g0696(.A(n1568), .B(n1394), .C(n1318), .Y(n1702));
  NAND3X1 g0697(.A(n1702), .B(n1701), .C(n1592), .Y(n1703));
  AOI21X1 g0698(.A0(n1677), .A1(n1282), .B0(n1703), .Y(n1704));
  NOR2X1  g0699(.A(n1704), .B(n1639), .Y(n1705));
  INVX1   g0700(.A(INSTQUEUE_REG_7__2__SCAN_IN), .Y(n1706));
  AOI22X1 g0701(.A0(n1244), .A1(INSTQUEUE_REG_0__2__SCAN_IN), .B0(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n1246), .Y(n1707));
  OAI21X1 g0702(.A0(n1243), .A1(n1706), .B0(n1707), .Y(n1708));
  INVX1   g0703(.A(INSTQUEUE_REG_4__2__SCAN_IN), .Y(n1709));
  AOI22X1 g0704(.A0(n1253), .A1(INSTQUEUE_REG_11__2__SCAN_IN), .B0(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n1255), .Y(n1710));
  OAI21X1 g0705(.A0(n1251), .A1(n1709), .B0(n1710), .Y(n1711));
  INVX1   g0706(.A(INSTQUEUE_REG_8__2__SCAN_IN), .Y(n1712));
  INVX1   g0707(.A(INSTQUEUE_REG_1__2__SCAN_IN), .Y(n1713));
  OAI22X1 g0708(.A0(n1261), .A1(n1713), .B0(n1712), .B1(n1263), .Y(n1714));
  AOI22X1 g0709(.A0(n1266), .A1(INSTQUEUE_REG_13__2__SCAN_IN), .B0(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n1268), .Y(n1715));
  AOI22X1 g0710(.A0(n1270), .A1(INSTQUEUE_REG_5__2__SCAN_IN), .B0(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n1271), .Y(n1716));
  AOI22X1 g0711(.A0(n1273), .A1(INSTQUEUE_REG_3__2__SCAN_IN), .B0(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n1275), .Y(n1717));
  AOI22X1 g0712(.A0(n1278), .A1(INSTQUEUE_REG_6__2__SCAN_IN), .B0(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n1279), .Y(n1718));
  NAND4X1 g0713(.A(n1717), .B(n1716), .C(n1715), .D(n1718), .Y(n1719));
  NOR4X1  g0714(.A(n1714), .B(n1711), .C(n1708), .D(n1719), .Y(n1720));
  NAND2X1 g0715(.A(n1464), .B(n1447), .Y(n1721));
  NAND2X1 g0716(.A(n1568), .B(n1394), .Y(n1722));
  AOI21X1 g0717(.A0(n1722), .A1(n1701), .B0(n1721), .Y(n1723));
  INVX1   g0718(.A(n1723), .Y(n1724));
  NOR3X1  g0719(.A(n1672), .B(n1592), .C(n1447), .Y(n1725));
  OAI21X1 g0720(.A0(n1725), .A1(n1720), .B0(n1724), .Y(n1726));
  NOR2X1  g0721(.A(n1726), .B(n1705), .Y(n1727));
  INVX1   g0722(.A(n1727), .Y(n1728));
  NOR3X1  g0723(.A(n1678), .B(n1672), .C(n1656), .Y(n1729));
  INVX1   g0724(.A(n1729), .Y(n1730));
  INVX1   g0725(.A(n1241), .Y(n1731));
  NOR3X1  g0726(.A(n1513), .B(n1502), .C(n1490), .Y(n1732));
  AOI21X1 g0727(.A0(n1732), .A1(n1520), .B0(n1731), .Y(n1733));
  INVX1   g0728(.A(n1733), .Y(n1734));
  NOR3X1  g0729(.A(n1734), .B(n1730), .C(READY_N), .Y(n1735));
  NOR2X1  g0730(.A(n1671), .B(n1422), .Y(n1736));
  NOR3X1  g0731(.A(n1736), .B(n1318), .C(n1282), .Y(n1737));
  NOR3X1  g0732(.A(n1639), .B(n1464), .C(n1447), .Y(n1738));
  NOR4X1  g0733(.A(n1737), .B(n1735), .C(n1728), .D(n1738), .Y(n1739));
  OAI21X1 g0734(.A0(n1685), .A1(n1536), .B0(n1739), .Y(n1740));
  AOI21X1 g0735(.A0(n1682), .A1(n1536), .B0(n1740), .Y(n1741));
  INVX1   g0736(.A(n1741), .Y(n1742));
  NAND2X1 g0737(.A(n1671), .B(n1422), .Y(n1743));
  AOI21X1 g0738(.A0(n1568), .A1(n1403), .B0(n1639), .Y(n1744));
  NAND2X1 g0739(.A(n1744), .B(n1743), .Y(n1745));
  AOI21X1 g0740(.A0(n1422), .A1(n1318), .B0(n1615), .Y(n1746));
  AOI21X1 g0741(.A0(n1677), .A1(n1592), .B0(n1746), .Y(n1747));
  NOR2X1  g0742(.A(n1568), .B(n1394), .Y(n1748));
  OAI21X1 g0743(.A0(n1700), .A1(n1671), .B0(n1318), .Y(n1749));
  OAI21X1 g0744(.A0(n1749), .A1(n1748), .B0(n1639), .Y(n1750));
  NAND3X1 g0745(.A(n1750), .B(n1747), .C(n1745), .Y(n1751));
  AOI21X1 g0746(.A0(n1394), .A1(n1318), .B0(n1464), .Y(n1752));
  AOI21X1 g0747(.A0(n1751), .A1(n1464), .B0(n1752), .Y(n1753));
  NOR2X1  g0748(.A(n1753), .B(n1447), .Y(n1754));
  NAND3X1 g0749(.A(n1720), .B(n1655), .C(n1282), .Y(n1755));
  NAND2X1 g0750(.A(n1639), .B(n1568), .Y(n1756));
  AOI21X1 g0751(.A0(n1756), .A1(n1755), .B0(n1464), .Y(n1757));
  NOR2X1  g0752(.A(n1655), .B(n1464), .Y(n1758));
  OAI21X1 g0753(.A0(n1758), .A1(n1447), .B0(n1639), .Y(n1759));
  NOR2X1  g0754(.A(n1592), .B(n1282), .Y(n1760));
  NOR2X1  g0755(.A(n1760), .B(n1737), .Y(n1761));
  NAND2X1 g0756(.A(n1761), .B(n1759), .Y(n1762));
  NAND2X1 g0757(.A(n1592), .B(n1362), .Y(n1763));
  NOR3X1  g0758(.A(n1671), .B(n1422), .C(n1403), .Y(n1764));
  NOR3X1  g0759(.A(n1764), .B(n1748), .C(n1700), .Y(n1765));
  OAI21X1 g0760(.A0(n1765), .A1(n1763), .B0(n1724), .Y(n1766));
  NOR4X1  g0761(.A(n1762), .B(n1757), .C(n1754), .D(n1766), .Y(n1767));
  NOR2X1  g0762(.A(n1763), .B(n1672), .Y(n1768));
  NOR2X1  g0763(.A(n1639), .B(n1592), .Y(n1769));
  NOR3X1  g0764(.A(n1394), .B(n1362), .C(n1447), .Y(n1770));
  NAND2X1 g0765(.A(n1770), .B(n1769), .Y(n1771));
  INVX1   g0766(.A(n1771), .Y(n1772));
  NOR2X1  g0767(.A(n1671), .B(n1394), .Y(n1773));
  NOR2X1  g0768(.A(n1615), .B(n1403), .Y(n1774));
  NAND4X1 g0769(.A(n1639), .B(n1655), .C(n1773), .D(n1774), .Y(n1775));
  INVX1   g0770(.A(n1755), .Y(n1776));
  NAND4X1 g0771(.A(n1671), .B(n1422), .C(n1318), .D(n1700), .Y(n1777));
  INVX1   g0772(.A(n1777), .Y(n1778));
  AOI22X1 g0773(.A0(n1776), .A1(n1778), .B0(n1700), .B1(n1362), .Y(n1779));
  NAND3X1 g0774(.A(n1779), .B(n1775), .C(n1730), .Y(n1780));
  NOR4X1  g0775(.A(n1772), .B(n1768), .C(n1640), .D(n1780), .Y(n1781));
  NAND2X1 g0776(.A(n1781), .B(n1767), .Y(n1782));
  INVX1   g0777(.A(n1782), .Y(n1783));
  AOI21X1 g0778(.A0(n1568), .A1(n1394), .B0(n1318), .Y(n1784));
  NOR4X1  g0779(.A(n1764), .B(n1748), .C(n1700), .D(n1784), .Y(n1785));
  AOI21X1 g0780(.A0(n1720), .A1(n1655), .B0(n1282), .Y(n1786));
  AOI21X1 g0781(.A0(n1786), .A1(n1785), .B0(n1464), .Y(n1787));
  NOR4X1  g0782(.A(n1568), .B(n1422), .C(n1403), .D(n1700), .Y(n1788));
  NOR3X1  g0783(.A(n1217), .B(STATE2_REG_1__SCAN_IN), .C(STATE2_REG_3__SCAN_IN), .Y(n1789));
  OAI21X1 g0784(.A0(n1720), .A1(n1282), .B0(n1789), .Y(n1790));
  AOI21X1 g0785(.A0(n1758), .A1(n1788), .B0(n1790), .Y(n1791));
  NAND2X1 g0786(.A(n1791), .B(n1775), .Y(n1792));
  NAND3X1 g0787(.A(n1615), .B(n1568), .C(n1403), .Y(n1793));
  AOI21X1 g0788(.A0(n1793), .A1(n1777), .B0(n1755), .Y(n1794));
  NOR4X1  g0789(.A(n1748), .B(n1616), .C(n1403), .D(n1736), .Y(n1795));
  NOR2X1  g0790(.A(n1795), .B(n1721), .Y(n1796));
  NOR4X1  g0791(.A(n1794), .B(n1792), .C(n1787), .D(n1796), .Y(n1797));
  OAI21X1 g0792(.A0(n1753), .A1(n1447), .B0(n1797), .Y(n1798));
  NOR3X1  g0793(.A(n1700), .B(n1671), .C(n1318), .Y(n1799));
  NAND2X1 g0794(.A(n1799), .B(n1769), .Y(n1800));
  NAND4X1 g0795(.A(n1750), .B(n1747), .C(n1745), .D(n1800), .Y(n1801));
  NAND2X1 g0796(.A(n1801), .B(n1467), .Y(n1802));
  NOR3X1  g0797(.A(n1785), .B(n1683), .C(n1217), .Y(n1803));
  NAND2X1 g0798(.A(n1615), .B(n1671), .Y(n1804));
  NOR4X1  g0799(.A(n1804), .B(n1403), .C(n1217), .D(n1771), .Y(n1805));
  NOR3X1  g0800(.A(n1777), .B(n1755), .C(n1217), .Y(n1806));
  NAND3X1 g0801(.A(n1655), .B(n1447), .C(STATE2_REG_0__SCAN_IN), .Y(n1807));
  NAND2X1 g0802(.A(n1807), .B(n1493), .Y(n1808));
  NOR4X1  g0803(.A(n1806), .B(n1805), .C(n1803), .D(n1808), .Y(n1809));
  NAND4X1 g0804(.A(n1381), .B(n1380), .C(n1419), .D(n1393), .Y(n1810));
  NOR2X1  g0805(.A(n1810), .B(n1418), .Y(n1811));
  NOR2X1  g0806(.A(n1811), .B(n1671), .Y(n1812));
  NOR4X1  g0807(.A(n1748), .B(n1700), .C(n1403), .D(n1812), .Y(n1813));
  OAI21X1 g0808(.A0(n1813), .A1(n1721), .B0(n1759), .Y(n1814));
  NAND2X1 g0809(.A(n1814), .B(STATE2_REG_0__SCAN_IN), .Y(n1815));
  NAND2X1 g0810(.A(n1720), .B(n1655), .Y(n1816));
  NAND3X1 g0811(.A(n1422), .B(n1464), .C(n1282), .Y(n1817));
  NAND3X1 g0812(.A(n1615), .B(n1671), .C(n1403), .Y(n1818));
  NOR4X1  g0813(.A(n1817), .B(n1816), .C(n1217), .D(n1818), .Y(n1819));
  NAND4X1 g0814(.A(n1639), .B(n1773), .C(STATE2_REG_0__SCAN_IN), .D(n1774), .Y(n1820));
  NAND3X1 g0815(.A(n1758), .B(n1788), .C(STATE2_REG_0__SCAN_IN), .Y(n1821));
  NAND2X1 g0816(.A(n1821), .B(n1820), .Y(n1822));
  NOR2X1  g0817(.A(n1700), .B(n1655), .Y(n1823));
  NOR2X1  g0818(.A(n1639), .B(n1403), .Y(n1824));
  NAND3X1 g0819(.A(n1824), .B(n1823), .C(n1773), .Y(n1825));
  NOR2X1  g0820(.A(n1362), .B(n1447), .Y(n1826));
  NOR3X1  g0821(.A(n1720), .B(n1592), .C(n1217), .Y(n1827));
  NAND3X1 g0822(.A(n1827), .B(n1826), .C(n1788), .Y(n1828));
  NOR2X1  g0823(.A(n1464), .B(n1282), .Y(n1829));
  NOR4X1  g0824(.A(n1362), .B(n1282), .C(n1217), .D(n1674), .Y(n1830));
  AOI21X1 g0825(.A0(n1829), .A1(STATE2_REG_0__SCAN_IN), .B0(n1830), .Y(n1831));
  OAI21X1 g0826(.A0(n1831), .A1(n1825), .B0(n1828), .Y(n1832));
  INVX1   g0827(.A(STATE2_REG_2__SCAN_IN), .Y(n1833));
  NOR2X1  g0828(.A(STATE2_REG_1__SCAN_IN), .B(n1833), .Y(n1834));
  NOR4X1  g0829(.A(STATE2_REG_0__SCAN_IN), .B(STATE2_REG_1__SCAN_IN), .C(STATE2_REG_3__SCAN_IN), .D(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Y(n1835));
  INVX1   g0830(.A(n1835), .Y(n1836));
  OAI21X1 g0831(.A0(n1834), .A1(n1229), .B0(n1836), .Y(n1837));
  NOR4X1  g0832(.A(n1832), .B(n1822), .C(n1819), .D(n1837), .Y(n1838));
  NAND4X1 g0833(.A(n1815), .B(n1809), .C(n1802), .D(n1838), .Y(n1839));
  NOR2X1  g0834(.A(n1837), .B(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n1840));
  INVX1   g0835(.A(n1840), .Y(n1841));
  NAND2X1 g0836(.A(n1841), .B(n1839), .Y(n1842));
  XOR2X1  g0837(.A(n1842), .B(n1798), .Y(n1843));
  NOR3X1  g0838(.A(n1678), .B(n1677), .C(n1639), .Y(n1844));
  NOR2X1  g0839(.A(n1844), .B(n1684), .Y(n1845));
  INVX1   g0840(.A(n1845), .Y(n1846));
  NOR2X1  g0841(.A(n1464), .B(n1447), .Y(n1847));
  INVX1   g0842(.A(n1847), .Y(n1848));
  NOR4X1  g0843(.A(n1656), .B(n1848), .C(n1231), .D(n1672), .Y(n1849));
  AOI21X1 g0844(.A0(n1846), .A1(n1231), .B0(n1849), .Y(n1850));
  OAI21X1 g0845(.A0(n1843), .A1(n1783), .B0(n1850), .Y(n1851));
  NOR2X1  g0846(.A(n1742), .B(n1231), .Y(n1852));
  AOI21X1 g0847(.A0(n1851), .A1(n1742), .B0(n1852), .Y(n1853));
  OAI21X1 g0848(.A0(n1671), .A1(n1318), .B0(n1720), .Y(n1854));
  NOR2X1  g0849(.A(n1854), .B(n1748), .Y(n1855));
  NOR4X1  g0850(.A(n1671), .B(n1422), .C(n1318), .D(n1700), .Y(n1856));
  OAI21X1 g0851(.A0(n1394), .A1(n1403), .B0(n1700), .Y(n1857));
  OAI21X1 g0852(.A0(n1856), .A1(n1655), .B0(n1857), .Y(n1858));
  AOI21X1 g0853(.A0(n1615), .A1(n1568), .B0(n1403), .Y(n1859));
  AOI21X1 g0854(.A0(n1859), .A1(n1743), .B0(n1720), .Y(n1860));
  NOR3X1  g0855(.A(n1860), .B(n1858), .C(n1855), .Y(n1861));
  INVX1   g0856(.A(n1752), .Y(n1862));
  OAI21X1 g0857(.A0(n1861), .A1(n1362), .B0(n1862), .Y(n1863));
  OAI21X1 g0858(.A0(n1671), .A1(n1422), .B0(n1403), .Y(n1864));
  NAND4X1 g0859(.A(n1864), .B(n1702), .C(n1701), .D(n1786), .Y(n1865));
  NAND2X1 g0860(.A(n1865), .B(n1362), .Y(n1866));
  NOR2X1  g0861(.A(n1362), .B(n1282), .Y(n1867));
  NAND4X1 g0862(.A(n1743), .B(n1823), .C(n1318), .D(n1722), .Y(n1868));
  AOI21X1 g0863(.A0(n1868), .A1(n1867), .B0(n1794), .Y(n1869));
  NAND4X1 g0864(.A(n1791), .B(n1866), .C(n1775), .D(n1869), .Y(n1870));
  AOI21X1 g0865(.A0(n1863), .A1(n1282), .B0(n1870), .Y(n1871));
  NAND3X1 g0866(.A(n1464), .B(n1282), .C(STATE2_REG_0__SCAN_IN), .Y(n1872));
  NOR2X1  g0867(.A(n1793), .B(n1816), .Y(n1873));
  NOR4X1  g0868(.A(n1860), .B(n1858), .C(n1855), .D(n1873), .Y(n1874));
  NOR2X1  g0869(.A(n1874), .B(n1872), .Y(n1875));
  NAND3X1 g0870(.A(n1864), .B(n1702), .C(n1701), .Y(n1876));
  NAND4X1 g0871(.A(n1758), .B(n1447), .C(STATE2_REG_0__SCAN_IN), .D(n1876), .Y(n1877));
  NOR4X1  g0872(.A(n1816), .B(n1804), .C(n1403), .D(n1817), .Y(n1878));
  NAND2X1 g0873(.A(n1878), .B(STATE2_REG_0__SCAN_IN), .Y(n1879));
  NOR2X1  g0874(.A(n1808), .B(n1806), .Y(n1880));
  NAND3X1 g0875(.A(n1880), .B(n1879), .C(n1877), .Y(n1881));
  OAI21X1 g0876(.A0(n1810), .A1(n1418), .B0(n1568), .Y(n1882));
  NAND4X1 g0877(.A(n1743), .B(n1615), .C(n1318), .D(n1882), .Y(n1883));
  NAND2X1 g0878(.A(n1883), .B(n1867), .Y(n1884));
  AOI21X1 g0879(.A0(n1884), .A1(n1759), .B0(n1217), .Y(n1885));
  NAND2X1 g0880(.A(n1700), .B(n1318), .Y(n1886));
  NOR4X1  g0881(.A(n1720), .B(n1569), .C(n1217), .D(n1886), .Y(n1887));
  NOR3X1  g0882(.A(n1763), .B(n1672), .C(n1217), .Y(n1888));
  NOR3X1  g0883(.A(n1888), .B(n1887), .C(n1819), .Y(n1889));
  NOR4X1  g0884(.A(n1672), .B(n1656), .C(n1217), .D(n1678), .Y(n1890));
  INVX1   g0885(.A(n1674), .Y(n1891));
  NAND4X1 g0886(.A(n1464), .B(n1447), .C(STATE2_REG_0__SCAN_IN), .D(n1891), .Y(n1892));
  OAI21X1 g0887(.A0(n1448), .A1(n1217), .B0(n1892), .Y(n1893));
  AOI21X1 g0888(.A0(n1893), .A1(n1640), .B0(n1890), .Y(n1894));
  INVX1   g0889(.A(n1837), .Y(n1895));
  NAND3X1 g0890(.A(n1895), .B(n1894), .C(n1889), .Y(n1896));
  NOR4X1  g0891(.A(n1885), .B(n1881), .C(n1875), .D(n1896), .Y(n1897));
  NOR3X1  g0892(.A(n1840), .B(n1897), .C(n1871), .Y(n1898));
  NOR3X1  g0893(.A(n1755), .B(n1804), .C(n1483), .Y(n1899));
  NOR2X1  g0894(.A(n1899), .B(n1832), .Y(n1900));
  AOI21X1 g0895(.A0(n1860), .A1(n1467), .B0(n1819), .Y(n1901));
  NAND3X1 g0896(.A(n1901), .B(n1879), .C(n1877), .Y(n1902));
  NOR3X1  g0897(.A(n1888), .B(n1887), .C(n1806), .Y(n1903));
  NAND3X1 g0898(.A(n1799), .B(n1769), .C(n1467), .Y(n1904));
  NOR3X1  g0899(.A(n1592), .B(n1282), .C(n1217), .Y(n1905));
  NOR3X1  g0900(.A(STATE2_REG_0__SCAN_IN), .B(STATE2_REG_1__SCAN_IN), .C(STATE2_REG_3__SCAN_IN), .Y(n1906));
  INVX1   g0901(.A(n1906), .Y(n1907));
  XOR2X1  g0902(.A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n1228), .Y(n1908));
  NOR2X1  g0903(.A(n1908), .B(n1907), .Y(n1909));
  INVX1   g0904(.A(STATE2_REG_1__SCAN_IN), .Y(n1910));
  AOI21X1 g0905(.A0(n1910), .A1(STATE2_REG_2__SCAN_IN), .B0(n1228), .Y(n1911));
  NOR4X1  g0906(.A(n1909), .B(n1905), .C(n1465), .D(n1911), .Y(n1912));
  NAND4X1 g0907(.A(n1904), .B(n1903), .C(n1894), .D(n1912), .Y(n1913));
  AOI21X1 g0908(.A0(n1747), .A1(n1745), .B0(n1872), .Y(n1914));
  NOR4X1  g0909(.A(n1913), .B(n1902), .C(n1885), .D(n1914), .Y(n1915));
  OAI21X1 g0910(.A0(n1834), .A1(n1228), .B0(n1245), .Y(n1916));
  NOR2X1  g0911(.A(n1916), .B(n1909), .Y(n1917));
  NOR3X1  g0912(.A(n1917), .B(n1915), .C(n1900), .Y(n1918));
  INVX1   g0913(.A(n1804), .Y(n1919));
  NAND3X1 g0914(.A(n1776), .B(n1919), .C(n1395), .Y(n1920));
  NAND2X1 g0915(.A(n1920), .B(n1894), .Y(n1921));
  NOR3X1  g0916(.A(n1700), .B(n1568), .C(n1318), .Y(n1922));
  NAND3X1 g0917(.A(n1922), .B(n1770), .C(n1769), .Y(n1923));
  OAI22X1 g0918(.A0(n1750), .A1(n1872), .B0(n1217), .B1(n1923), .Y(n1924));
  NOR3X1  g0919(.A(n1924), .B(n1805), .C(n1803), .Y(n1925));
  NAND2X1 g0920(.A(n1912), .B(n1904), .Y(n1926));
  NOR2X1  g0921(.A(n1926), .B(n1832), .Y(n1927));
  AOI21X1 g0922(.A0(n1814), .A1(STATE2_REG_0__SCAN_IN), .B0(n1914), .Y(n1928));
  NAND4X1 g0923(.A(n1927), .B(n1903), .C(n1925), .D(n1928), .Y(n1929));
  INVX1   g0924(.A(n1917), .Y(n1930));
  AOI21X1 g0925(.A0(n1930), .A1(n1929), .B0(n1921), .Y(n1931));
  NOR3X1  g0926(.A(n1931), .B(n1918), .C(n1898), .Y(n1932));
  NAND3X1 g0927(.A(n1841), .B(n1839), .C(n1798), .Y(n1933));
  NAND3X1 g0928(.A(n1930), .B(n1929), .C(n1921), .Y(n1934));
  OAI21X1 g0929(.A0(n1917), .A1(n1915), .B0(n1900), .Y(n1935));
  AOI21X1 g0930(.A0(n1935), .A1(n1934), .B0(n1933), .Y(n1936));
  NOR2X1  g0931(.A(n1936), .B(n1932), .Y(n1937));
  NOR3X1  g0932(.A(n1845), .B(n1544), .C(n1250), .Y(n1938));
  AOI21X1 g0933(.A0(n1673), .A1(n1245), .B0(n1938), .Y(n1939));
  OAI21X1 g0934(.A0(n1937), .A1(n1783), .B0(n1939), .Y(n1940));
  INVX1   g0935(.A(n1940), .Y(n1941));
  NOR2X1  g0936(.A(n1941), .B(n1741), .Y(n1942));
  AOI21X1 g0937(.A0(n1741), .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B0(n1942), .Y(n1943));
  NAND3X1 g0938(.A(n1943), .B(n1853), .C(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Y(n1944));
  NOR2X1  g0939(.A(n1229), .B(n1228), .Y(n1945));
  NAND2X1 g0940(.A(n1943), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Y(n1946));
  OAI21X1 g0941(.A0(n1931), .A1(n1933), .B0(n1934), .Y(n1947));
  NOR3X1  g0942(.A(n1832), .B(n1822), .C(n1819), .Y(n1948));
  NAND4X1 g0943(.A(n1815), .B(n1809), .C(n1802), .D(n1948), .Y(n1949));
  INVX1   g0944(.A(n1834), .Y(n1950));
  XOR2X1  g0945(.A(n1945), .B(n1224), .Y(n1951));
  NOR2X1  g0946(.A(n1951), .B(n1907), .Y(n1952));
  AOI21X1 g0947(.A0(n1950), .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B0(n1952), .Y(n1953));
  INVX1   g0948(.A(n1953), .Y(n1954));
  AOI21X1 g0949(.A0(n1950), .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B0(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Y(n1955));
  OAI21X1 g0950(.A0(n1951), .A1(n1907), .B0(n1955), .Y(n1956));
  OAI21X1 g0951(.A0(n1954), .A1(n1949), .B0(n1956), .Y(n1957));
  XOR2X1  g0952(.A(n1957), .B(n1947), .Y(n1958));
  NOR2X1  g0953(.A(n1684), .B(n1679), .Y(n1959));
  INVX1   g0954(.A(n1959), .Y(n1960));
  NOR3X1  g0955(.A(n1231), .B(n1245), .C(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Y(n1961));
  AOI21X1 g0956(.A0(n1252), .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B0(n1961), .Y(n1962));
  INVX1   g0957(.A(n1673), .Y(n1963));
  XOR2X1  g0958(.A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n1226), .Y(n1964));
  NOR3X1  g0959(.A(n1755), .B(n1677), .C(n1362), .Y(n1965));
  INVX1   g0960(.A(n1965), .Y(n1966));
  OAI22X1 g0961(.A0(n1964), .A1(n1963), .B0(n1962), .B1(n1966), .Y(n1967));
  AOI21X1 g0962(.A0(n1962), .A1(n1960), .B0(n1967), .Y(n1968));
  OAI21X1 g0963(.A0(n1958), .A1(n1783), .B0(n1968), .Y(n1969));
  INVX1   g0964(.A(n1969), .Y(n1970));
  NAND2X1 g0965(.A(n1741), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Y(n1971));
  OAI21X1 g0966(.A0(n1970), .A1(n1741), .B0(n1971), .Y(n1972));
  OAI21X1 g0967(.A0(n1972), .A1(n1224), .B0(n1946), .Y(n1973));
  AOI21X1 g0968(.A0(n1945), .A1(n1853), .B0(n1973), .Y(n1974));
  NAND2X1 g0969(.A(n1974), .B(n1944), .Y(n1975));
  INVX1   g0970(.A(n1952), .Y(n1976));
  NOR2X1  g0971(.A(n1954), .B(n1949), .Y(n1977));
  AOI21X1 g0972(.A0(n1955), .A1(n1976), .B0(n1977), .Y(n1978));
  NAND2X1 g0973(.A(n1978), .B(n1947), .Y(n1979));
  AOI21X1 g0974(.A0(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B0(n1220), .Y(n1980));
  NOR4X1  g0975(.A(n1228), .B(n1224), .C(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .D(n1229), .Y(n1981));
  NOR2X1  g0976(.A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n1220), .Y(n1982));
  NOR3X1  g0977(.A(n1982), .B(n1981), .C(n1980), .Y(n1983));
  INVX1   g0978(.A(n1983), .Y(n1984));
  AOI22X1 g0979(.A0(n1906), .A1(n1984), .B0(n1950), .B1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .Y(n1985));
  INVX1   g0980(.A(n1985), .Y(n1986));
  AOI21X1 g0981(.A0(n1949), .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B0(n1986), .Y(n1987));
  XOR2X1  g0982(.A(n1987), .B(n1979), .Y(n1988));
  INVX1   g0983(.A(n1988), .Y(n1989));
  AOI21X1 g0984(.A0(n1252), .A1(n1226), .B0(n1222), .Y(n1990));
  AOI21X1 g0985(.A0(n1252), .A1(n1260), .B0(n1990), .Y(n1991));
  AOI22X1 g0986(.A0(n1543), .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B0(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(n1277), .Y(n1992));
  INVX1   g0987(.A(n1992), .Y(n1993));
  OAI21X1 g0988(.A0(n1252), .A1(n1226), .B0(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n1994));
  NAND2X1 g0989(.A(n1994), .B(n1243), .Y(n1995));
  AOI22X1 g0990(.A0(n1993), .A1(n1673), .B0(n1965), .B1(n1995), .Y(n1996));
  INVX1   g0991(.A(n1996), .Y(n1997));
  AOI21X1 g0992(.A0(n1991), .A1(n1960), .B0(n1997), .Y(n1998));
  OAI21X1 g0993(.A0(n1989), .A1(n1783), .B0(n1998), .Y(n1999));
  NAND2X1 g0994(.A(n1999), .B(n1742), .Y(n2000));
  OAI21X1 g0995(.A0(n1742), .A1(n1222), .B0(n2000), .Y(n2001));
  AOI22X1 g0996(.A0(n1972), .A1(n1224), .B0(n1220), .B1(n2001), .Y(n2002));
  NOR4X1  g0997(.A(n1656), .B(n1848), .C(n1217), .D(n1672), .Y(n2003));
  NOR2X1  g0998(.A(n2003), .B(n1890), .Y(n2004));
  NOR2X1  g0999(.A(n2004), .B(n1218), .Y(n2005));
  NOR2X1  g1000(.A(n1987), .B(n1957), .Y(n2006));
  NAND2X1 g1001(.A(n2006), .B(n1947), .Y(n2007));
  XOR2X1  g1002(.A(n2007), .B(n2005), .Y(n2008));
  NOR2X1  g1003(.A(n2008), .B(n1730), .Y(n2009));
  NAND2X1 g1004(.A(n2009), .B(n1742), .Y(n2010));
  OAI21X1 g1005(.A0(n1742), .A1(n1218), .B0(n2010), .Y(n2011));
  OAI22X1 g1006(.A0(n2001), .A1(n1220), .B0(n1238), .B1(n2011), .Y(n2012));
  AOI21X1 g1007(.A0(n2002), .A1(n1975), .B0(n2012), .Y(n2013));
  NOR2X1  g1008(.A(n1910), .B(FLUSH_REG_SCAN_IN), .Y(n2014));
  INVX1   g1009(.A(FLUSH_REG_SCAN_IN), .Y(n2015));
  INVX1   g1010(.A(INSTADDRPOINTER_REG_0__SCAN_IN), .Y(n2016));
  NOR2X1  g1011(.A(n2016), .B(n1910), .Y(n2017));
  INVX1   g1012(.A(n2017), .Y(n2018));
  XOR2X1  g1013(.A(INSTADDRPOINTER_REG_1__SCAN_IN), .B(n2016), .Y(n2019));
  INVX1   g1014(.A(n2019), .Y(n2020));
  INVX1   g1015(.A(INSTADDRPOINTER_REG_1__SCAN_IN), .Y(n2021));
  NOR2X1  g1016(.A(INSTADDRPOINTER_REG_31__SCAN_IN), .B(n2021), .Y(n2022));
  AOI21X1 g1017(.A0(n2020), .A1(INSTADDRPOINTER_REG_31__SCAN_IN), .B0(n2022), .Y(n2023));
  NOR3X1  g1018(.A(n2023), .B(n2018), .C(n2015), .Y(n2024));
  AOI21X1 g1019(.A0(n2014), .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B0(n2024), .Y(n2025));
  INVX1   g1020(.A(n2025), .Y(n2026));
  AOI21X1 g1021(.A0(n1972), .A1(n1910), .B0(n2026), .Y(n2027));
  AOI22X1 g1022(.A0(n2011), .A1(n1910), .B0(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B1(n2014), .Y(n2028));
  AOI22X1 g1023(.A0(n2001), .A1(n1910), .B0(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(n2014), .Y(n2029));
  OAI21X1 g1024(.A0(n2029), .A1(n2027), .B0(n2028), .Y(n2030));
  NAND2X1 g1025(.A(n2011), .B(n1238), .Y(n2031));
  INVX1   g1026(.A(n1536), .Y(n2032));
  OAI21X1 g1027(.A0(n1825), .A1(n2032), .B0(n1447), .Y(n2033));
  NOR2X1  g1028(.A(n1536), .B(n1464), .Y(n2034));
  INVX1   g1029(.A(n2034), .Y(n2035));
  NOR2X1  g1030(.A(n1672), .B(n1656), .Y(n2036));
  INVX1   g1031(.A(n2036), .Y(n2037));
  NOR2X1  g1032(.A(n1733), .B(n1362), .Y(n2038));
  OAI21X1 g1033(.A0(n2038), .A1(n2037), .B0(n1282), .Y(n2039));
  NAND3X1 g1034(.A(n2039), .B(n2035), .C(n2033), .Y(n2040));
  NOR2X1  g1035(.A(n1674), .B(STATE_REG_0__SCAN_IN), .Y(n2041));
  INVX1   g1036(.A(n2041), .Y(n2042));
  NAND3X1 g1037(.A(n1678), .B(n2042), .C(n1448), .Y(n2043));
  AOI21X1 g1038(.A0(n2043), .A1(n1113), .B0(n2040), .Y(n2044));
  OAI21X1 g1039(.A0(FLUSH_REG_SCAN_IN), .A1(MORE_REG_SCAN_IN), .B0(n2044), .Y(n2045));
  NOR3X1  g1040(.A(n1672), .B(n1639), .C(n1655), .Y(n2046));
  NOR4X1  g1041(.A(n1655), .B(n1403), .C(n1282), .D(n1639), .Y(n2047));
  OAI21X1 g1042(.A0(n2046), .A1(n1773), .B0(n2047), .Y(n2048));
  NOR2X1  g1043(.A(n1679), .B(n1673), .Y(n2049));
  NAND2X1 g1044(.A(n2049), .B(n2048), .Y(n2050));
  NAND2X1 g1045(.A(n2050), .B(n2032), .Y(n2051));
  AOI22X1 g1046(.A0(n1729), .A1(n1734), .B0(n1684), .B1(n1536), .Y(n2052));
  AOI21X1 g1047(.A0(n2052), .A1(n2051), .B0(n1700), .Y(n2053));
  NAND2X1 g1048(.A(n1536), .B(n1447), .Y(n2054));
  NOR4X1  g1049(.A(n1672), .B(n1639), .C(n1655), .D(n2054), .Y(n2055));
  NOR2X1  g1050(.A(n2055), .B(n2053), .Y(n2056));
  NAND3X1 g1051(.A(n2056), .B(n2045), .C(n2031), .Y(n2057));
  NOR4X1  g1052(.A(n2030), .B(n2013), .C(STATE2_REG_1__SCAN_IN), .D(n2057), .Y(n2058));
  NOR2X1  g1053(.A(n2042), .B(n2032), .Y(n2059));
  INVX1   g1054(.A(n2059), .Y(n2060));
  NOR2X1  g1055(.A(STATEBS16_REG_SCAN_IN), .B(READY_N), .Y(n2061));
  INVX1   g1056(.A(n2061), .Y(n2062));
  NOR4X1  g1057(.A(n2060), .B(n1825), .C(n1721), .D(n2062), .Y(n2063));
  AOI21X1 g1058(.A0(STATE2_REG_1__SCAN_IN), .A1(READY_N), .B0(STATE2_REG_0__SCAN_IN), .Y(n2064));
  NOR3X1  g1059(.A(n2064), .B(n2063), .C(n1833), .Y(n2065));
  AOI21X1 g1060(.A0(n2065), .A1(n2058), .B0(n1217), .Y(n2066));
  NOR3X1  g1061(.A(n2057), .B(n2030), .C(n2013), .Y(n2067));
  NAND3X1 g1062(.A(STATE2_REG_0__SCAN_IN), .B(STATE2_REG_1__SCAN_IN), .C(STATE2_REG_2__SCAN_IN), .Y(n2068));
  OAI21X1 g1063(.A0(n2066), .A1(n1216), .B0(n2068), .Y(U3453));
  OAI21X1 g1064(.A0(STATE2_REG_2__SCAN_IN), .A1(READY_N), .B0(STATE2_REG_0__SCAN_IN), .Y(n2070));
  INVX1   g1065(.A(STATEBS16_REG_SCAN_IN), .Y(n2071));
  AOI21X1 g1066(.A0(n1217), .A1(n2071), .B0(n1910), .Y(n2072));
  AOI21X1 g1067(.A0(n2072), .A1(n2070), .B0(n1834), .Y(n2073));
  OAI21X1 g1068(.A0(n2066), .A1(n1833), .B0(n2073), .Y(U3150));
  NOR2X1  g1069(.A(STATE2_REG_1__SCAN_IN), .B(STATE2_REG_3__SCAN_IN), .Y(n2075));
  NAND3X1 g1070(.A(n2066), .B(n2075), .C(n1113), .Y(n2076));
  NOR2X1  g1071(.A(n2058), .B(n1217), .Y(n2077));
  NOR4X1  g1072(.A(n2063), .B(n2077), .C(n1833), .D(n2064), .Y(n2078));
  NOR3X1  g1073(.A(n1217), .B(STATE2_REG_2__SCAN_IN), .C(n1113), .Y(n2079));
  OAI21X1 g1074(.A0(n2079), .A1(n2078), .B0(STATE2_REG_1__SCAN_IN), .Y(n2080));
  OAI21X1 g1075(.A0(n2058), .A1(n1217), .B0(n2065), .Y(n2081));
  NOR4X1  g1076(.A(n1910), .B(STATE2_REG_2__SCAN_IN), .C(STATEBS16_REG_SCAN_IN), .D(STATE2_REG_0__SCAN_IN), .Y(n2082));
  NOR3X1  g1077(.A(n1217), .B(STATE2_REG_1__SCAN_IN), .C(n1833), .Y(n2083));
  AOI21X1 g1078(.A0(n2083), .A1(n2081), .B0(n2082), .Y(n2084));
  NAND3X1 g1079(.A(n2084), .B(n2080), .C(n2076), .Y(U3149));
  NOR2X1  g1080(.A(n1910), .B(n1833), .Y(n2086));
  INVX1   g1081(.A(n2086), .Y(n2087));
  NOR2X1  g1082(.A(n1853), .B(STATE2_REG_1__SCAN_IN), .Y(n2088));
  NAND2X1 g1083(.A(n2023), .B(n2017), .Y(n2089));
  NOR2X1  g1084(.A(n2089), .B(n2015), .Y(n2090));
  NAND3X1 g1085(.A(n2016), .B(STATE2_REG_1__SCAN_IN), .C(FLUSH_REG_SCAN_IN), .Y(n2091));
  OAI21X1 g1086(.A0(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B0(n2014), .Y(n2092));
  NAND2X1 g1087(.A(n2092), .B(n2091), .Y(n2093));
  NOR2X1  g1088(.A(n2093), .B(n2090), .Y(n2094));
  OAI21X1 g1089(.A0(n1943), .A1(STATE2_REG_1__SCAN_IN), .B0(n2094), .Y(n2095));
  NOR2X1  g1090(.A(n2029), .B(n2027), .Y(n2096));
  OAI21X1 g1091(.A0(n2095), .A1(n2088), .B0(n2096), .Y(n2097));
  NAND2X1 g1092(.A(n2097), .B(n2028), .Y(n2098));
  NOR2X1  g1093(.A(n2098), .B(n2087), .Y(n2099));
  OAI21X1 g1094(.A0(n2099), .A1(n2078), .B0(STATE2_REG_0__SCAN_IN), .Y(n2100));
  NAND4X1 g1095(.A(n1910), .B(n1833), .C(STATE2_REG_3__SCAN_IN), .D(n1536), .Y(n2101));
  NAND3X1 g1096(.A(n2101), .B(n2081), .C(n1217), .Y(n2102));
  INVX1   g1097(.A(n2083), .Y(n2103));
  NOR2X1  g1098(.A(n2103), .B(n2067), .Y(n2104));
  NOR4X1  g1099(.A(STATE2_REG_1__SCAN_IN), .B(STATE2_REG_2__SCAN_IN), .C(n1216), .D(n1217), .Y(n2105));
  NOR3X1  g1100(.A(n2105), .B(n2104), .C(n2079), .Y(n2106));
  NAND3X1 g1101(.A(n2106), .B(n2102), .C(n2100), .Y(U3148));
  NOR2X1  g1102(.A(n2032), .B(n1216), .Y(n2108));
  INVX1   g1103(.A(n2108), .Y(n2109));
  XOR2X1  g1104(.A(STATE2_REG_1__SCAN_IN), .B(n1833), .Y(n2110));
  AOI21X1 g1105(.A0(n2110), .A1(n2109), .B0(STATE2_REG_0__SCAN_IN), .Y(n2111));
  NOR4X1  g1106(.A(n1228), .B(n1224), .C(n1220), .D(n1229), .Y(n2112));
  NOR2X1  g1107(.A(n1989), .B(n1958), .Y(n2113));
  NAND3X1 g1108(.A(n1935), .B(n1934), .C(n1933), .Y(n2114));
  OAI21X1 g1109(.A0(n1931), .A1(n1918), .B0(n1898), .Y(n2115));
  AOI21X1 g1110(.A0(n2115), .A1(n2114), .B0(n1843), .Y(n2116));
  AOI21X1 g1111(.A0(n2116), .A1(n2113), .B0(n2112), .Y(n2117));
  NOR3X1  g1112(.A(STATE2_REG_2__SCAN_IN), .B(STATE2_REG_3__SCAN_IN), .C(STATEBS16_REG_SCAN_IN), .Y(n2118));
  NOR3X1  g1113(.A(STATE2_REG_2__SCAN_IN), .B(STATE2_REG_3__SCAN_IN), .C(n2071), .Y(n2119));
  NAND2X1 g1114(.A(n2111), .B(n2119), .Y(n2120));
  NOR2X1  g1115(.A(n1403), .B(n1217), .Y(n2121));
  NAND2X1 g1116(.A(n1244), .B(INSTQUEUE_REG_1__7__SCAN_IN), .Y(n2124));
  OAI21X1 g1117(.A0(n1343), .A1(n1594), .B0(n2124), .Y(n2125));
  NAND2X1 g1118(.A(n1246), .B(INSTQUEUE_REG_3__7__SCAN_IN), .Y(n2127));
  NAND2X1 g1119(.A(n1337), .B(INSTQUEUE_REG_2__7__SCAN_IN), .Y(n2129));
  NAND2X1 g1120(.A(n2129), .B(n2127), .Y(n2130));
  NOR2X1  g1121(.A(n2130), .B(n2125), .Y(n2131));
  NAND2X1 g1122(.A(n1273), .B(INSTQUEUE_REG_4__7__SCAN_IN), .Y(n2133));
  NAND2X1 g1123(.A(n1329), .B(INSTQUEUE_REG_5__7__SCAN_IN), .Y(n2135));
  NAND2X1 g1124(.A(n2135), .B(n2133), .Y(n2136));
  NAND2X1 g1125(.A(n1278), .B(INSTQUEUE_REG_7__7__SCAN_IN), .Y(n2138));
  NAND2X1 g1126(.A(n1270), .B(INSTQUEUE_REG_6__7__SCAN_IN), .Y(n2140));
  NAND2X1 g1127(.A(n2140), .B(n2138), .Y(n2141));
  NOR2X1  g1128(.A(n2141), .B(n2136), .Y(n2142));
  NAND2X1 g1129(.A(n1253), .B(INSTQUEUE_REG_12__7__SCAN_IN), .Y(n2144));
  NAND2X1 g1130(.A(n1271), .B(INSTQUEUE_REG_13__7__SCAN_IN), .Y(n2146));
  NAND2X1 g1131(.A(n2146), .B(n2144), .Y(n2147));
  NAND2X1 g1132(.A(n1279), .B(INSTQUEUE_REG_15__7__SCAN_IN), .Y(n2149));
  NAND2X1 g1133(.A(n1266), .B(INSTQUEUE_REG_14__7__SCAN_IN), .Y(n2151));
  NAND2X1 g1134(.A(n2151), .B(n2149), .Y(n2152));
  NOR2X1  g1135(.A(n2152), .B(n2147), .Y(n2153));
  NAND2X1 g1136(.A(n1323), .B(INSTQUEUE_REG_8__7__SCAN_IN), .Y(n2155));
  NAND2X1 g1137(.A(n1338), .B(INSTQUEUE_REG_9__7__SCAN_IN), .Y(n2157));
  NAND2X1 g1138(.A(n2157), .B(n2155), .Y(n2158));
  NAND2X1 g1139(.A(n1255), .B(INSTQUEUE_REG_11__7__SCAN_IN), .Y(n2160));
  NAND2X1 g1140(.A(n1275), .B(INSTQUEUE_REG_10__7__SCAN_IN), .Y(n2162));
  NAND2X1 g1141(.A(n2162), .B(n2160), .Y(n2163));
  NOR2X1  g1142(.A(n2163), .B(n2158), .Y(n2164));
  NAND4X1 g1143(.A(n2153), .B(n2142), .C(n2131), .D(n2164), .Y(n2165));
  NAND2X1 g1144(.A(n2165), .B(n2121), .Y(n2166));
  INVX1   g1145(.A(n2166), .Y(n2167));
  AOI22X1 g1146(.A0(n1268), .A1(INSTQUEUE_REG_0__0__SCAN_IN), .B0(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n1244), .Y(n2169));
  AOI22X1 g1147(.A0(n1246), .A1(INSTQUEUE_REG_3__0__SCAN_IN), .B0(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n1337), .Y(n2170));
  AOI22X1 g1148(.A0(n1273), .A1(INSTQUEUE_REG_4__0__SCAN_IN), .B0(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n1329), .Y(n2171));
  AOI22X1 g1149(.A0(n1278), .A1(INSTQUEUE_REG_7__0__SCAN_IN), .B0(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n1270), .Y(n2172));
  NAND4X1 g1150(.A(n2171), .B(n2170), .C(n2169), .D(n2172), .Y(n2173));
  AOI22X1 g1151(.A0(n1253), .A1(INSTQUEUE_REG_12__0__SCAN_IN), .B0(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n1271), .Y(n2174));
  AOI22X1 g1152(.A0(n1279), .A1(INSTQUEUE_REG_15__0__SCAN_IN), .B0(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n1266), .Y(n2175));
  AOI22X1 g1153(.A0(n1323), .A1(INSTQUEUE_REG_8__0__SCAN_IN), .B0(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n1338), .Y(n2176));
  AOI22X1 g1154(.A0(n1255), .A1(INSTQUEUE_REG_11__0__SCAN_IN), .B0(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n1275), .Y(n2177));
  NAND4X1 g1155(.A(n2176), .B(n2175), .C(n2174), .D(n2177), .Y(n2178));
  NOR2X1  g1156(.A(n2178), .B(n2173), .Y(n2179));
  NOR3X1  g1157(.A(n2179), .B(n1447), .C(n1217), .Y(n2180));
  INVX1   g1158(.A(n2165), .Y(n2181));
  NOR2X1  g1159(.A(n2181), .B(n1403), .Y(n2182));
  NOR4X1  g1160(.A(n1282), .B(n1426), .C(n1217), .D(n1318), .Y(n2183));
  NOR4X1  g1161(.A(n2182), .B(n2180), .C(n1217), .D(n2183), .Y(n2184));
  XOR2X1  g1162(.A(n1842), .B(n1871), .Y(n2185));
  NOR4X1  g1163(.A(n2165), .B(n1403), .C(n1217), .D(n2179), .Y(n2186));
  AOI21X1 g1164(.A0(n2179), .A1(n2167), .B0(n2186), .Y(n2187));
  INVX1   g1165(.A(n2187), .Y(n2188));
  AOI21X1 g1166(.A0(n2185), .A1(n1217), .B0(n2188), .Y(n2189));
  XOR2X1  g1167(.A(n2189), .B(n2167), .Y(n2190));
  XOR2X1  g1168(.A(n2190), .B(n2184), .Y(n2191));
  XOR2X1  g1169(.A(n2191), .B(n2167), .Y(n2192));
  INVX1   g1170(.A(n2184), .Y(n2193));
  OAI21X1 g1171(.A0(n2190), .A1(n2184), .B0(n2166), .Y(n2195));
  AOI21X1 g1172(.A0(n2115), .A1(n2114), .B0(STATE2_REG_0__SCAN_IN), .Y(n2196));
  AOI22X1 g1173(.A0(n1268), .A1(INSTQUEUE_REG_0__1__SCAN_IN), .B0(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n1244), .Y(n2197));
  AOI22X1 g1174(.A0(n1246), .A1(INSTQUEUE_REG_3__1__SCAN_IN), .B0(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n1337), .Y(n2198));
  AOI22X1 g1175(.A0(n1273), .A1(INSTQUEUE_REG_4__1__SCAN_IN), .B0(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n1329), .Y(n2199));
  AOI22X1 g1176(.A0(n1278), .A1(INSTQUEUE_REG_7__1__SCAN_IN), .B0(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n1270), .Y(n2200));
  NAND4X1 g1177(.A(n2199), .B(n2198), .C(n2197), .D(n2200), .Y(n2201));
  AOI22X1 g1178(.A0(n1253), .A1(INSTQUEUE_REG_12__1__SCAN_IN), .B0(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n1271), .Y(n2202));
  AOI22X1 g1179(.A0(n1279), .A1(INSTQUEUE_REG_15__1__SCAN_IN), .B0(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n1266), .Y(n2203));
  AOI22X1 g1180(.A0(n1323), .A1(INSTQUEUE_REG_8__1__SCAN_IN), .B0(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n1338), .Y(n2204));
  AOI22X1 g1181(.A0(n1255), .A1(INSTQUEUE_REG_11__1__SCAN_IN), .B0(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n1275), .Y(n2205));
  NAND4X1 g1182(.A(n2204), .B(n2203), .C(n2202), .D(n2205), .Y(n2206));
  NOR2X1  g1183(.A(n2206), .B(n2201), .Y(n2207));
  NOR4X1  g1184(.A(n2165), .B(n1403), .C(n1217), .D(n2207), .Y(n2208));
  AOI21X1 g1185(.A0(n2207), .A1(n2167), .B0(n2208), .Y(n2209));
  INVX1   g1186(.A(n2209), .Y(n2210));
  NOR2X1  g1187(.A(n2210), .B(n2196), .Y(n2211));
  XOR2X1  g1188(.A(n2211), .B(n2167), .Y(n2212));
  OAI21X1 g1189(.A0(n2206), .A1(n2201), .B0(n1476), .Y(n2213));
  NOR3X1  g1190(.A(n2165), .B(n1403), .C(n1217), .Y(n2214));
  AOI21X1 g1191(.A0(n1319), .A1(INSTQUEUE_REG_0__1__SCAN_IN), .B0(n2214), .Y(n2215));
  NAND2X1 g1192(.A(n2215), .B(n2213), .Y(n2216));
  XOR2X1  g1193(.A(n2216), .B(n2212), .Y(n2217));
  XOR2X1  g1194(.A(n2217), .B(n2195), .Y(n2218));
  AOI22X1 g1195(.A0(n1268), .A1(INSTQUEUE_REG_0__2__SCAN_IN), .B0(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n1244), .Y(n2219));
  AOI22X1 g1196(.A0(n1246), .A1(INSTQUEUE_REG_3__2__SCAN_IN), .B0(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n1337), .Y(n2220));
  AOI22X1 g1197(.A0(n1273), .A1(INSTQUEUE_REG_4__2__SCAN_IN), .B0(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n1329), .Y(n2221));
  AOI22X1 g1198(.A0(n1278), .A1(INSTQUEUE_REG_7__2__SCAN_IN), .B0(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n1270), .Y(n2222));
  NAND4X1 g1199(.A(n2221), .B(n2220), .C(n2219), .D(n2222), .Y(n2223));
  AOI22X1 g1200(.A0(n1253), .A1(INSTQUEUE_REG_12__2__SCAN_IN), .B0(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n1271), .Y(n2224));
  AOI22X1 g1201(.A0(n1279), .A1(INSTQUEUE_REG_15__2__SCAN_IN), .B0(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n1266), .Y(n2225));
  AOI22X1 g1202(.A0(n1323), .A1(INSTQUEUE_REG_8__2__SCAN_IN), .B0(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n1338), .Y(n2226));
  AOI22X1 g1203(.A0(n1255), .A1(INSTQUEUE_REG_11__2__SCAN_IN), .B0(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n1275), .Y(n2227));
  NAND4X1 g1204(.A(n2226), .B(n2225), .C(n2224), .D(n2227), .Y(n2228));
  NOR2X1  g1205(.A(n2228), .B(n2223), .Y(n2229));
  INVX1   g1206(.A(n2229), .Y(n2230));
  AOI22X1 g1207(.A0(n1476), .A1(n2230), .B0(n1319), .B1(INSTQUEUE_REG_0__2__SCAN_IN), .Y(n2231));
  NOR4X1  g1208(.A(n2165), .B(n1403), .C(n1217), .D(n2229), .Y(n2232));
  AOI21X1 g1209(.A0(n2229), .A1(n2167), .B0(n2232), .Y(n2233));
  OAI21X1 g1210(.A0(n1958), .A1(STATE2_REG_0__SCAN_IN), .B0(n2233), .Y(n2234));
  XOR2X1  g1211(.A(n2234), .B(n2166), .Y(n2235));
  XOR2X1  g1212(.A(n2235), .B(n2231), .Y(n2236));
  OAI21X1 g1213(.A0(n2210), .A1(n2196), .B0(n2166), .Y(n2237));
  OAI21X1 g1214(.A0(n1936), .A1(n1932), .B0(n1217), .Y(n2238));
  NAND3X1 g1215(.A(n2209), .B(n2238), .C(n2167), .Y(n2239));
  INVX1   g1216(.A(n2216), .Y(n2240));
  AOI21X1 g1217(.A0(n2239), .A1(n2237), .B0(n2240), .Y(n2241));
  NAND3X1 g1218(.A(n2240), .B(n2239), .C(n2237), .Y(n2242));
  AOI21X1 g1219(.A0(n2242), .A1(n2195), .B0(n2241), .Y(n2243));
  XOR2X1  g1220(.A(n2243), .B(n2236), .Y(n2244));
  AOI22X1 g1221(.A0(n1268), .A1(INSTQUEUE_REG_0__3__SCAN_IN), .B0(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n1244), .Y(n2245));
  AOI22X1 g1222(.A0(n1246), .A1(INSTQUEUE_REG_3__3__SCAN_IN), .B0(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n1337), .Y(n2246));
  AOI22X1 g1223(.A0(n1273), .A1(INSTQUEUE_REG_4__3__SCAN_IN), .B0(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n1329), .Y(n2247));
  AOI22X1 g1224(.A0(n1278), .A1(INSTQUEUE_REG_7__3__SCAN_IN), .B0(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n1270), .Y(n2248));
  NAND4X1 g1225(.A(n2247), .B(n2246), .C(n2245), .D(n2248), .Y(n2249));
  AOI22X1 g1226(.A0(n1253), .A1(INSTQUEUE_REG_12__3__SCAN_IN), .B0(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n1271), .Y(n2250));
  AOI22X1 g1227(.A0(n1279), .A1(INSTQUEUE_REG_15__3__SCAN_IN), .B0(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n1266), .Y(n2251));
  AOI22X1 g1228(.A0(n1323), .A1(INSTQUEUE_REG_8__3__SCAN_IN), .B0(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n1338), .Y(n2252));
  AOI22X1 g1229(.A0(n1255), .A1(INSTQUEUE_REG_11__3__SCAN_IN), .B0(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n1275), .Y(n2253));
  NAND4X1 g1230(.A(n2252), .B(n2251), .C(n2250), .D(n2253), .Y(n2254));
  NOR2X1  g1231(.A(n2254), .B(n2249), .Y(n2255));
  INVX1   g1232(.A(n2255), .Y(n2256));
  AOI22X1 g1233(.A0(n1476), .A1(n2256), .B0(n1319), .B1(INSTQUEUE_REG_0__3__SCAN_IN), .Y(n2257));
  NAND2X1 g1234(.A(n2256), .B(n2214), .Y(n2258));
  OAI21X1 g1235(.A0(n2256), .A1(n2166), .B0(n2258), .Y(n2259));
  AOI21X1 g1236(.A0(n1988), .A1(n1217), .B0(n2259), .Y(n2260));
  XOR2X1  g1237(.A(n2260), .B(n2166), .Y(n2261));
  XOR2X1  g1238(.A(n2261), .B(n2257), .Y(n2262));
  INVX1   g1239(.A(n2231), .Y(n2263));
  XOR2X1  g1240(.A(n2234), .B(n2167), .Y(n2264));
  NAND2X1 g1241(.A(n2264), .B(n2263), .Y(n2265));
  NOR2X1  g1242(.A(n2264), .B(n2263), .Y(n2266));
  OAI21X1 g1243(.A0(n2243), .A1(n2266), .B0(n2265), .Y(n2267));
  XOR2X1  g1244(.A(n2267), .B(n2262), .Y(n2268));
  NOR4X1  g1245(.A(n2244), .B(n2218), .C(n2192), .D(n2268), .Y(n2269));
  XOR2X1  g1246(.A(n2191), .B(n2166), .Y(n2270));
  NOR4X1  g1247(.A(n2244), .B(n2218), .C(n2270), .D(n2268), .Y(n2271));
  NOR3X1  g1248(.A(n2271), .B(n2269), .C(n2120), .Y(n2272));
  OAI21X1 g1249(.A0(n2272), .A1(n2118), .B0(n2117), .Y(n2273));
  NOR2X1  g1250(.A(n2112), .B(n1216), .Y(n2274));
  NAND3X1 g1251(.A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .Y(n2275));
  AOI21X1 g1252(.A0(n2275), .A1(STATE2_REG_2__SCAN_IN), .B0(n2274), .Y(n2276));
  NAND3X1 g1253(.A(n2276), .B(n2273), .C(n2111), .Y(n2277));
  NAND2X1 g1254(.A(n2277), .B(INSTQUEUE_REG_15__7__SCAN_IN), .Y(n2278));
  INVX1   g1255(.A(n2119), .Y(n2279));
  NOR3X1  g1256(.A(n2271), .B(n2269), .C(n2279), .Y(n2280));
  NOR2X1  g1257(.A(n2280), .B(n2118), .Y(n2281));
  OAI22X1 g1258(.A0(n2275), .A1(n1833), .B0(n2117), .B1(n2281), .Y(n2282));
  NAND3X1 g1259(.A(n2282), .B(n2111), .C(DATAI_7_), .Y(n2283));
  NAND4X1 g1260(.A(n2111), .B(n2119), .C(DATAI_31_), .D(n2269), .Y(n2284));
  INVX1   g1261(.A(DATAI_23_), .Y(n2285));
  NOR2X1  g1262(.A(n2120), .B(n2285), .Y(n2286));
  INVX1   g1263(.A(n2111), .Y(n2287));
  NOR3X1  g1264(.A(n2287), .B(n1700), .C(n1216), .Y(n2288));
  AOI22X1 g1265(.A0(n2286), .A1(n2271), .B0(n2112), .B1(n2288), .Y(n2289));
  NAND4X1 g1266(.A(n2284), .B(n2283), .C(n2278), .D(n2289), .Y(U3147));
  NAND2X1 g1267(.A(n2277), .B(INSTQUEUE_REG_15__6__SCAN_IN), .Y(n2291));
  NAND3X1 g1268(.A(n2282), .B(n2111), .C(DATAI_6_), .Y(n2292));
  NAND4X1 g1269(.A(n2111), .B(n2119), .C(DATAI_30_), .D(n2269), .Y(n2293));
  INVX1   g1270(.A(DATAI_22_), .Y(n2294));
  NOR2X1  g1271(.A(n2120), .B(n2294), .Y(n2295));
  NOR3X1  g1272(.A(n2287), .B(n1568), .C(n1216), .Y(n2296));
  AOI22X1 g1273(.A0(n2295), .A1(n2271), .B0(n2112), .B1(n2296), .Y(n2297));
  NAND4X1 g1274(.A(n2293), .B(n2292), .C(n2291), .D(n2297), .Y(U3146));
  NAND2X1 g1275(.A(n2277), .B(INSTQUEUE_REG_15__5__SCAN_IN), .Y(n2299));
  NAND3X1 g1276(.A(n2282), .B(n2111), .C(DATAI_5_), .Y(n2300));
  NAND4X1 g1277(.A(n2111), .B(n2119), .C(DATAI_29_), .D(n2269), .Y(n2301));
  INVX1   g1278(.A(DATAI_21_), .Y(n2302));
  NOR2X1  g1279(.A(n2120), .B(n2302), .Y(n2303));
  NOR3X1  g1280(.A(n2287), .B(n1422), .C(n1216), .Y(n2304));
  AOI22X1 g1281(.A0(n2303), .A1(n2271), .B0(n2112), .B1(n2304), .Y(n2305));
  NAND4X1 g1282(.A(n2301), .B(n2300), .C(n2299), .D(n2305), .Y(U3145));
  NAND2X1 g1283(.A(n2277), .B(INSTQUEUE_REG_15__4__SCAN_IN), .Y(n2307));
  NAND3X1 g1284(.A(n2282), .B(n2111), .C(DATAI_4_), .Y(n2308));
  NAND4X1 g1285(.A(n2111), .B(n2119), .C(DATAI_28_), .D(n2269), .Y(n2309));
  INVX1   g1286(.A(DATAI_20_), .Y(n2310));
  NOR2X1  g1287(.A(n2120), .B(n2310), .Y(n2311));
  NOR3X1  g1288(.A(n2287), .B(n1318), .C(n1216), .Y(n2312));
  AOI22X1 g1289(.A0(n2311), .A1(n2271), .B0(n2112), .B1(n2312), .Y(n2313));
  NAND4X1 g1290(.A(n2309), .B(n2308), .C(n2307), .D(n2313), .Y(U3144));
  NAND2X1 g1291(.A(n2277), .B(INSTQUEUE_REG_15__3__SCAN_IN), .Y(n2315));
  NAND3X1 g1292(.A(n2282), .B(n2111), .C(DATAI_3_), .Y(n2316));
  NAND4X1 g1293(.A(n2111), .B(n2119), .C(DATAI_27_), .D(n2269), .Y(n2317));
  INVX1   g1294(.A(DATAI_19_), .Y(n2318));
  NOR2X1  g1295(.A(n2120), .B(n2318), .Y(n2319));
  NOR3X1  g1296(.A(n2287), .B(n1655), .C(n1216), .Y(n2320));
  AOI22X1 g1297(.A0(n2319), .A1(n2271), .B0(n2112), .B1(n2320), .Y(n2321));
  NAND4X1 g1298(.A(n2317), .B(n2316), .C(n2315), .D(n2321), .Y(U3143));
  NAND2X1 g1299(.A(n2277), .B(INSTQUEUE_REG_15__2__SCAN_IN), .Y(n2323));
  NAND3X1 g1300(.A(n2282), .B(n2111), .C(DATAI_2_), .Y(n2324));
  NAND4X1 g1301(.A(n2111), .B(n2119), .C(DATAI_26_), .D(n2269), .Y(n2325));
  INVX1   g1302(.A(DATAI_18_), .Y(n2326));
  NOR2X1  g1303(.A(n2120), .B(n2326), .Y(n2327));
  NOR3X1  g1304(.A(n2287), .B(n1720), .C(n1216), .Y(n2328));
  AOI22X1 g1305(.A0(n2327), .A1(n2271), .B0(n2112), .B1(n2328), .Y(n2329));
  NAND4X1 g1306(.A(n2325), .B(n2324), .C(n2323), .D(n2329), .Y(U3142));
  NAND2X1 g1307(.A(n2277), .B(INSTQUEUE_REG_15__1__SCAN_IN), .Y(n2331));
  NAND3X1 g1308(.A(n2282), .B(n2111), .C(DATAI_1_), .Y(n2332));
  NAND4X1 g1309(.A(n2111), .B(n2119), .C(DATAI_25_), .D(n2269), .Y(n2333));
  INVX1   g1310(.A(DATAI_17_), .Y(n2334));
  NOR2X1  g1311(.A(n2120), .B(n2334), .Y(n2335));
  NOR3X1  g1312(.A(n2287), .B(n1464), .C(n1216), .Y(n2336));
  AOI22X1 g1313(.A0(n2335), .A1(n2271), .B0(n2112), .B1(n2336), .Y(n2337));
  NAND4X1 g1314(.A(n2333), .B(n2332), .C(n2331), .D(n2337), .Y(U3141));
  NAND2X1 g1315(.A(n2277), .B(INSTQUEUE_REG_15__0__SCAN_IN), .Y(n2339));
  NAND3X1 g1316(.A(n2282), .B(n2111), .C(DATAI_0_), .Y(n2340));
  NAND4X1 g1317(.A(n2111), .B(n2119), .C(DATAI_24_), .D(n2269), .Y(n2341));
  INVX1   g1318(.A(DATAI_16_), .Y(n2342));
  NOR2X1  g1319(.A(n2120), .B(n2342), .Y(n2343));
  NOR3X1  g1320(.A(n2287), .B(n1282), .C(n1216), .Y(n2344));
  AOI22X1 g1321(.A0(n2343), .A1(n2271), .B0(n2112), .B1(n2344), .Y(n2345));
  NAND4X1 g1322(.A(n2341), .B(n2340), .C(n2339), .D(n2345), .Y(U3140));
  NOR4X1  g1323(.A(n1228), .B(n1224), .C(n1220), .D(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Y(n2347));
  AOI21X1 g1324(.A0(n2115), .A1(n2114), .B0(n2185), .Y(n2348));
  AOI21X1 g1325(.A0(n2348), .A1(n2113), .B0(n2347), .Y(n2349));
  XOR2X1  g1326(.A(n2189), .B(n2166), .Y(n2350));
  AOI21X1 g1327(.A0(n2350), .A1(n2193), .B0(n2167), .Y(n2353));
  XOR2X1  g1328(.A(n2217), .B(n2353), .Y(n2354));
  NOR4X1  g1329(.A(n2244), .B(n2354), .C(n2270), .D(n2268), .Y(n2355));
  NOR3X1  g1330(.A(n2269), .B(n2355), .C(n2120), .Y(n2358));
  OAI21X1 g1331(.A0(n2358), .A1(n2118), .B0(n2349), .Y(n2359));
  NOR2X1  g1332(.A(n2347), .B(n1216), .Y(n2360));
  INVX1   g1333(.A(n1908), .Y(n2361));
  NOR2X1  g1334(.A(n1983), .B(n1951), .Y(n2362));
  NAND2X1 g1335(.A(n2362), .B(n2361), .Y(n2363));
  AOI21X1 g1336(.A0(n2363), .A1(STATE2_REG_2__SCAN_IN), .B0(n2360), .Y(n2364));
  NAND3X1 g1337(.A(n2364), .B(n2359), .C(n2111), .Y(n2365));
  NAND2X1 g1338(.A(n2365), .B(INSTQUEUE_REG_14__7__SCAN_IN), .Y(n2366));
  NOR3X1  g1339(.A(n2269), .B(n2355), .C(n2279), .Y(n2367));
  NOR2X1  g1340(.A(n2367), .B(n2118), .Y(n2368));
  OAI22X1 g1341(.A0(n2363), .A1(n1833), .B0(n2349), .B1(n2368), .Y(n2369));
  NAND3X1 g1342(.A(n2369), .B(n2111), .C(DATAI_7_), .Y(n2370));
  NAND4X1 g1343(.A(n2111), .B(n2119), .C(DATAI_31_), .D(n2355), .Y(n2371));
  AOI22X1 g1344(.A0(n2347), .A1(n2288), .B0(n2286), .B1(n2269), .Y(n2372));
  NAND4X1 g1345(.A(n2371), .B(n2370), .C(n2366), .D(n2372), .Y(U3139));
  NAND2X1 g1346(.A(n2365), .B(INSTQUEUE_REG_14__6__SCAN_IN), .Y(n2374));
  NAND3X1 g1347(.A(n2369), .B(n2111), .C(DATAI_6_), .Y(n2375));
  NAND4X1 g1348(.A(n2111), .B(n2119), .C(DATAI_30_), .D(n2355), .Y(n2376));
  AOI22X1 g1349(.A0(n2347), .A1(n2296), .B0(n2295), .B1(n2269), .Y(n2377));
  NAND4X1 g1350(.A(n2376), .B(n2375), .C(n2374), .D(n2377), .Y(U3138));
  NAND2X1 g1351(.A(n2365), .B(INSTQUEUE_REG_14__5__SCAN_IN), .Y(n2379));
  NAND3X1 g1352(.A(n2369), .B(n2111), .C(DATAI_5_), .Y(n2380));
  NAND4X1 g1353(.A(n2111), .B(n2119), .C(DATAI_29_), .D(n2355), .Y(n2381));
  AOI22X1 g1354(.A0(n2347), .A1(n2304), .B0(n2303), .B1(n2269), .Y(n2382));
  NAND4X1 g1355(.A(n2381), .B(n2380), .C(n2379), .D(n2382), .Y(U3137));
  NAND2X1 g1356(.A(n2365), .B(INSTQUEUE_REG_14__4__SCAN_IN), .Y(n2384));
  NAND3X1 g1357(.A(n2369), .B(n2111), .C(DATAI_4_), .Y(n2385));
  NAND4X1 g1358(.A(n2111), .B(n2119), .C(DATAI_28_), .D(n2355), .Y(n2386));
  AOI22X1 g1359(.A0(n2347), .A1(n2312), .B0(n2311), .B1(n2269), .Y(n2387));
  NAND4X1 g1360(.A(n2386), .B(n2385), .C(n2384), .D(n2387), .Y(U3136));
  NAND2X1 g1361(.A(n2365), .B(INSTQUEUE_REG_14__3__SCAN_IN), .Y(n2389));
  NAND3X1 g1362(.A(n2369), .B(n2111), .C(DATAI_3_), .Y(n2390));
  NAND4X1 g1363(.A(n2111), .B(n2119), .C(DATAI_27_), .D(n2355), .Y(n2391));
  AOI22X1 g1364(.A0(n2347), .A1(n2320), .B0(n2319), .B1(n2269), .Y(n2392));
  NAND4X1 g1365(.A(n2391), .B(n2390), .C(n2389), .D(n2392), .Y(U3135));
  NAND2X1 g1366(.A(n2365), .B(INSTQUEUE_REG_14__2__SCAN_IN), .Y(n2394));
  NAND3X1 g1367(.A(n2369), .B(n2111), .C(DATAI_2_), .Y(n2395));
  NAND4X1 g1368(.A(n2111), .B(n2119), .C(DATAI_26_), .D(n2355), .Y(n2396));
  AOI22X1 g1369(.A0(n2347), .A1(n2328), .B0(n2327), .B1(n2269), .Y(n2397));
  NAND4X1 g1370(.A(n2396), .B(n2395), .C(n2394), .D(n2397), .Y(U3134));
  NAND2X1 g1371(.A(n2365), .B(INSTQUEUE_REG_14__1__SCAN_IN), .Y(n2399));
  NAND3X1 g1372(.A(n2369), .B(n2111), .C(DATAI_1_), .Y(n2400));
  NAND4X1 g1373(.A(n2111), .B(n2119), .C(DATAI_25_), .D(n2355), .Y(n2401));
  AOI22X1 g1374(.A0(n2347), .A1(n2336), .B0(n2335), .B1(n2269), .Y(n2402));
  NAND4X1 g1375(.A(n2401), .B(n2400), .C(n2399), .D(n2402), .Y(U3133));
  NAND2X1 g1376(.A(n2365), .B(INSTQUEUE_REG_14__0__SCAN_IN), .Y(n2404));
  NAND3X1 g1377(.A(n2369), .B(n2111), .C(DATAI_0_), .Y(n2405));
  NAND4X1 g1378(.A(n2111), .B(n2119), .C(DATAI_24_), .D(n2355), .Y(n2406));
  AOI22X1 g1379(.A0(n2347), .A1(n2344), .B0(n2343), .B1(n2269), .Y(n2407));
  NAND4X1 g1380(.A(n2406), .B(n2405), .C(n2404), .D(n2407), .Y(U3132));
  NOR4X1  g1381(.A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n1224), .C(n1220), .D(n1229), .Y(n2409));
  NOR3X1  g1382(.A(n1936), .B(n1932), .C(n1843), .Y(n2410));
  AOI21X1 g1383(.A0(n2410), .A1(n2113), .B0(n2409), .Y(n2411));
  NOR4X1  g1384(.A(n2244), .B(n2354), .C(n2192), .D(n2268), .Y(n2412));
  NAND2X1 g1385(.A(n2218), .B(n2192), .Y(n2413));
  NOR3X1  g1386(.A(n2355), .B(n2412), .C(n2120), .Y(n2415));
  OAI21X1 g1387(.A0(n2415), .A1(n2118), .B0(n2411), .Y(n2416));
  NOR2X1  g1388(.A(n2409), .B(n1216), .Y(n2417));
  NAND3X1 g1389(.A(n1228), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .Y(n2418));
  AOI21X1 g1390(.A0(n2418), .A1(STATE2_REG_2__SCAN_IN), .B0(n2417), .Y(n2419));
  NAND3X1 g1391(.A(n2419), .B(n2416), .C(n2111), .Y(n2420));
  NAND2X1 g1392(.A(n2420), .B(INSTQUEUE_REG_13__7__SCAN_IN), .Y(n2421));
  NOR3X1  g1393(.A(n2355), .B(n2412), .C(n2279), .Y(n2422));
  NOR2X1  g1394(.A(n2422), .B(n2118), .Y(n2423));
  OAI22X1 g1395(.A0(n2418), .A1(n1833), .B0(n2411), .B1(n2423), .Y(n2424));
  NAND3X1 g1396(.A(n2424), .B(n2111), .C(DATAI_7_), .Y(n2425));
  NAND4X1 g1397(.A(n2111), .B(n2119), .C(DATAI_31_), .D(n2412), .Y(n2426));
  AOI22X1 g1398(.A0(n2409), .A1(n2288), .B0(n2286), .B1(n2355), .Y(n2427));
  NAND4X1 g1399(.A(n2426), .B(n2425), .C(n2421), .D(n2427), .Y(U3131));
  NAND2X1 g1400(.A(n2420), .B(INSTQUEUE_REG_13__6__SCAN_IN), .Y(n2429));
  NAND3X1 g1401(.A(n2424), .B(n2111), .C(DATAI_6_), .Y(n2430));
  NAND4X1 g1402(.A(n2111), .B(n2119), .C(DATAI_30_), .D(n2412), .Y(n2431));
  AOI22X1 g1403(.A0(n2409), .A1(n2296), .B0(n2295), .B1(n2355), .Y(n2432));
  NAND4X1 g1404(.A(n2431), .B(n2430), .C(n2429), .D(n2432), .Y(U3130));
  NAND2X1 g1405(.A(n2420), .B(INSTQUEUE_REG_13__5__SCAN_IN), .Y(n2434));
  NAND3X1 g1406(.A(n2424), .B(n2111), .C(DATAI_5_), .Y(n2435));
  NAND4X1 g1407(.A(n2111), .B(n2119), .C(DATAI_29_), .D(n2412), .Y(n2436));
  AOI22X1 g1408(.A0(n2409), .A1(n2304), .B0(n2303), .B1(n2355), .Y(n2437));
  NAND4X1 g1409(.A(n2436), .B(n2435), .C(n2434), .D(n2437), .Y(U3129));
  NAND2X1 g1410(.A(n2420), .B(INSTQUEUE_REG_13__4__SCAN_IN), .Y(n2439));
  NAND3X1 g1411(.A(n2424), .B(n2111), .C(DATAI_4_), .Y(n2440));
  NAND4X1 g1412(.A(n2111), .B(n2119), .C(DATAI_28_), .D(n2412), .Y(n2441));
  AOI22X1 g1413(.A0(n2409), .A1(n2312), .B0(n2311), .B1(n2355), .Y(n2442));
  NAND4X1 g1414(.A(n2441), .B(n2440), .C(n2439), .D(n2442), .Y(U3128));
  NAND2X1 g1415(.A(n2420), .B(INSTQUEUE_REG_13__3__SCAN_IN), .Y(n2444));
  NAND3X1 g1416(.A(n2424), .B(n2111), .C(DATAI_3_), .Y(n2445));
  NAND4X1 g1417(.A(n2111), .B(n2119), .C(DATAI_27_), .D(n2412), .Y(n2446));
  AOI22X1 g1418(.A0(n2409), .A1(n2320), .B0(n2319), .B1(n2355), .Y(n2447));
  NAND4X1 g1419(.A(n2446), .B(n2445), .C(n2444), .D(n2447), .Y(U3127));
  NAND2X1 g1420(.A(n2420), .B(INSTQUEUE_REG_13__2__SCAN_IN), .Y(n2449));
  NAND3X1 g1421(.A(n2424), .B(n2111), .C(DATAI_2_), .Y(n2450));
  NAND4X1 g1422(.A(n2111), .B(n2119), .C(DATAI_26_), .D(n2412), .Y(n2451));
  AOI22X1 g1423(.A0(n2409), .A1(n2328), .B0(n2327), .B1(n2355), .Y(n2452));
  NAND4X1 g1424(.A(n2451), .B(n2450), .C(n2449), .D(n2452), .Y(U3126));
  NAND2X1 g1425(.A(n2420), .B(INSTQUEUE_REG_13__1__SCAN_IN), .Y(n2454));
  NAND3X1 g1426(.A(n2424), .B(n2111), .C(DATAI_1_), .Y(n2455));
  NAND4X1 g1427(.A(n2111), .B(n2119), .C(DATAI_25_), .D(n2412), .Y(n2456));
  AOI22X1 g1428(.A0(n2409), .A1(n2336), .B0(n2335), .B1(n2355), .Y(n2457));
  NAND4X1 g1429(.A(n2456), .B(n2455), .C(n2454), .D(n2457), .Y(U3125));
  NAND2X1 g1430(.A(n2420), .B(INSTQUEUE_REG_13__0__SCAN_IN), .Y(n2459));
  NAND3X1 g1431(.A(n2424), .B(n2111), .C(DATAI_0_), .Y(n2460));
  NAND4X1 g1432(.A(n2111), .B(n2119), .C(DATAI_24_), .D(n2412), .Y(n2461));
  AOI22X1 g1433(.A0(n2409), .A1(n2344), .B0(n2343), .B1(n2355), .Y(n2462));
  NAND4X1 g1434(.A(n2461), .B(n2460), .C(n2459), .D(n2462), .Y(U3124));
  NOR4X1  g1435(.A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n1224), .C(n1220), .D(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Y(n2464));
  NOR3X1  g1436(.A(n1936), .B(n1932), .C(n2185), .Y(n2465));
  AOI21X1 g1437(.A0(n2465), .A1(n2113), .B0(n2464), .Y(n2466));
  XOR2X1  g1438(.A(n2235), .B(n2263), .Y(n2467));
  XOR2X1  g1439(.A(n2243), .B(n2467), .Y(n2468));
  NOR4X1  g1440(.A(n2468), .B(n2218), .C(n2270), .D(n2268), .Y(n2469));
  NAND2X1 g1441(.A(n2218), .B(n2270), .Y(n2470));
  NOR3X1  g1442(.A(n2412), .B(n2469), .C(n2120), .Y(n2472));
  OAI21X1 g1443(.A0(n2472), .A1(n2118), .B0(n2466), .Y(n2473));
  NOR2X1  g1444(.A(n2464), .B(n1216), .Y(n2474));
  NAND2X1 g1445(.A(n2362), .B(n1908), .Y(n2475));
  AOI21X1 g1446(.A0(n2475), .A1(STATE2_REG_2__SCAN_IN), .B0(n2474), .Y(n2476));
  NAND3X1 g1447(.A(n2476), .B(n2473), .C(n2111), .Y(n2477));
  NAND2X1 g1448(.A(n2477), .B(INSTQUEUE_REG_12__7__SCAN_IN), .Y(n2478));
  NOR3X1  g1449(.A(n2412), .B(n2469), .C(n2279), .Y(n2479));
  NOR2X1  g1450(.A(n2479), .B(n2118), .Y(n2480));
  OAI22X1 g1451(.A0(n2475), .A1(n1833), .B0(n2466), .B1(n2480), .Y(n2481));
  NAND3X1 g1452(.A(n2481), .B(n2111), .C(DATAI_7_), .Y(n2482));
  NAND4X1 g1453(.A(n2111), .B(n2119), .C(DATAI_31_), .D(n2469), .Y(n2483));
  AOI22X1 g1454(.A0(n2464), .A1(n2288), .B0(n2286), .B1(n2412), .Y(n2484));
  NAND4X1 g1455(.A(n2483), .B(n2482), .C(n2478), .D(n2484), .Y(U3123));
  NAND2X1 g1456(.A(n2477), .B(INSTQUEUE_REG_12__6__SCAN_IN), .Y(n2486));
  NAND3X1 g1457(.A(n2481), .B(n2111), .C(DATAI_6_), .Y(n2487));
  NAND4X1 g1458(.A(n2111), .B(n2119), .C(DATAI_30_), .D(n2469), .Y(n2488));
  AOI22X1 g1459(.A0(n2464), .A1(n2296), .B0(n2295), .B1(n2412), .Y(n2489));
  NAND4X1 g1460(.A(n2488), .B(n2487), .C(n2486), .D(n2489), .Y(U3122));
  NAND2X1 g1461(.A(n2477), .B(INSTQUEUE_REG_12__5__SCAN_IN), .Y(n2491));
  NAND3X1 g1462(.A(n2481), .B(n2111), .C(DATAI_5_), .Y(n2492));
  NAND4X1 g1463(.A(n2111), .B(n2119), .C(DATAI_29_), .D(n2469), .Y(n2493));
  AOI22X1 g1464(.A0(n2464), .A1(n2304), .B0(n2303), .B1(n2412), .Y(n2494));
  NAND4X1 g1465(.A(n2493), .B(n2492), .C(n2491), .D(n2494), .Y(U3121));
  NAND2X1 g1466(.A(n2477), .B(INSTQUEUE_REG_12__4__SCAN_IN), .Y(n2496));
  NAND3X1 g1467(.A(n2481), .B(n2111), .C(DATAI_4_), .Y(n2497));
  NAND4X1 g1468(.A(n2111), .B(n2119), .C(DATAI_28_), .D(n2469), .Y(n2498));
  AOI22X1 g1469(.A0(n2464), .A1(n2312), .B0(n2311), .B1(n2412), .Y(n2499));
  NAND4X1 g1470(.A(n2498), .B(n2497), .C(n2496), .D(n2499), .Y(U3120));
  NAND2X1 g1471(.A(n2477), .B(INSTQUEUE_REG_12__3__SCAN_IN), .Y(n2501));
  NAND3X1 g1472(.A(n2481), .B(n2111), .C(DATAI_3_), .Y(n2502));
  NAND4X1 g1473(.A(n2111), .B(n2119), .C(DATAI_27_), .D(n2469), .Y(n2503));
  AOI22X1 g1474(.A0(n2464), .A1(n2320), .B0(n2319), .B1(n2412), .Y(n2504));
  NAND4X1 g1475(.A(n2503), .B(n2502), .C(n2501), .D(n2504), .Y(U3119));
  NAND2X1 g1476(.A(n2477), .B(INSTQUEUE_REG_12__2__SCAN_IN), .Y(n2506));
  NAND3X1 g1477(.A(n2481), .B(n2111), .C(DATAI_2_), .Y(n2507));
  NAND4X1 g1478(.A(n2111), .B(n2119), .C(DATAI_26_), .D(n2469), .Y(n2508));
  AOI22X1 g1479(.A0(n2464), .A1(n2328), .B0(n2327), .B1(n2412), .Y(n2509));
  NAND4X1 g1480(.A(n2508), .B(n2507), .C(n2506), .D(n2509), .Y(U3118));
  NAND2X1 g1481(.A(n2477), .B(INSTQUEUE_REG_12__1__SCAN_IN), .Y(n2511));
  NAND3X1 g1482(.A(n2481), .B(n2111), .C(DATAI_1_), .Y(n2512));
  NAND4X1 g1483(.A(n2111), .B(n2119), .C(DATAI_25_), .D(n2469), .Y(n2513));
  AOI22X1 g1484(.A0(n2464), .A1(n2336), .B0(n2335), .B1(n2412), .Y(n2514));
  NAND4X1 g1485(.A(n2513), .B(n2512), .C(n2511), .D(n2514), .Y(U3117));
  NAND2X1 g1486(.A(n2477), .B(INSTQUEUE_REG_12__0__SCAN_IN), .Y(n2516));
  NAND3X1 g1487(.A(n2481), .B(n2111), .C(DATAI_0_), .Y(n2517));
  NAND4X1 g1488(.A(n2111), .B(n2119), .C(DATAI_24_), .D(n2469), .Y(n2518));
  AOI22X1 g1489(.A0(n2464), .A1(n2344), .B0(n2343), .B1(n2412), .Y(n2519));
  NAND4X1 g1490(.A(n2518), .B(n2517), .C(n2516), .D(n2519), .Y(U3116));
  NOR4X1  g1491(.A(n1228), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C(n1220), .D(n1229), .Y(n2521));
  INVX1   g1492(.A(n1958), .Y(n2522));
  NOR2X1  g1493(.A(n1989), .B(n2522), .Y(n2523));
  AOI21X1 g1494(.A0(n2523), .A1(n2116), .B0(n2521), .Y(n2524));
  NOR4X1  g1495(.A(n2468), .B(n2218), .C(n2192), .D(n2268), .Y(n2525));
  NOR3X1  g1496(.A(n2469), .B(n2525), .C(n2120), .Y(n2527));
  OAI21X1 g1497(.A0(n2527), .A1(n2118), .B0(n2524), .Y(n2528));
  NOR2X1  g1498(.A(n2521), .B(n1216), .Y(n2529));
  NAND3X1 g1499(.A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n1224), .C(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .Y(n2530));
  AOI21X1 g1500(.A0(n2530), .A1(STATE2_REG_2__SCAN_IN), .B0(n2529), .Y(n2531));
  NAND3X1 g1501(.A(n2531), .B(n2528), .C(n2111), .Y(n2532));
  NAND2X1 g1502(.A(n2532), .B(INSTQUEUE_REG_11__7__SCAN_IN), .Y(n2533));
  NOR3X1  g1503(.A(n2469), .B(n2525), .C(n2279), .Y(n2534));
  NOR2X1  g1504(.A(n2534), .B(n2118), .Y(n2535));
  OAI22X1 g1505(.A0(n2530), .A1(n1833), .B0(n2524), .B1(n2535), .Y(n2536));
  NAND3X1 g1506(.A(n2536), .B(n2111), .C(DATAI_7_), .Y(n2537));
  NAND4X1 g1507(.A(n2111), .B(n2119), .C(DATAI_31_), .D(n2525), .Y(n2538));
  AOI22X1 g1508(.A0(n2521), .A1(n2288), .B0(n2286), .B1(n2469), .Y(n2539));
  NAND4X1 g1509(.A(n2538), .B(n2537), .C(n2533), .D(n2539), .Y(U3115));
  NAND2X1 g1510(.A(n2532), .B(INSTQUEUE_REG_11__6__SCAN_IN), .Y(n2541));
  NAND3X1 g1511(.A(n2536), .B(n2111), .C(DATAI_6_), .Y(n2542));
  NAND4X1 g1512(.A(n2111), .B(n2119), .C(DATAI_30_), .D(n2525), .Y(n2543));
  AOI22X1 g1513(.A0(n2521), .A1(n2296), .B0(n2295), .B1(n2469), .Y(n2544));
  NAND4X1 g1514(.A(n2543), .B(n2542), .C(n2541), .D(n2544), .Y(U3114));
  NAND2X1 g1515(.A(n2532), .B(INSTQUEUE_REG_11__5__SCAN_IN), .Y(n2546));
  NAND3X1 g1516(.A(n2536), .B(n2111), .C(DATAI_5_), .Y(n2547));
  NAND4X1 g1517(.A(n2111), .B(n2119), .C(DATAI_29_), .D(n2525), .Y(n2548));
  AOI22X1 g1518(.A0(n2521), .A1(n2304), .B0(n2303), .B1(n2469), .Y(n2549));
  NAND4X1 g1519(.A(n2548), .B(n2547), .C(n2546), .D(n2549), .Y(U3113));
  NAND2X1 g1520(.A(n2532), .B(INSTQUEUE_REG_11__4__SCAN_IN), .Y(n2551));
  NAND3X1 g1521(.A(n2536), .B(n2111), .C(DATAI_4_), .Y(n2552));
  NAND4X1 g1522(.A(n2111), .B(n2119), .C(DATAI_28_), .D(n2525), .Y(n2553));
  AOI22X1 g1523(.A0(n2521), .A1(n2312), .B0(n2311), .B1(n2469), .Y(n2554));
  NAND4X1 g1524(.A(n2553), .B(n2552), .C(n2551), .D(n2554), .Y(U3112));
  NAND2X1 g1525(.A(n2532), .B(INSTQUEUE_REG_11__3__SCAN_IN), .Y(n2556));
  NAND3X1 g1526(.A(n2536), .B(n2111), .C(DATAI_3_), .Y(n2557));
  NAND4X1 g1527(.A(n2111), .B(n2119), .C(DATAI_27_), .D(n2525), .Y(n2558));
  AOI22X1 g1528(.A0(n2521), .A1(n2320), .B0(n2319), .B1(n2469), .Y(n2559));
  NAND4X1 g1529(.A(n2558), .B(n2557), .C(n2556), .D(n2559), .Y(U3111));
  NAND2X1 g1530(.A(n2532), .B(INSTQUEUE_REG_11__2__SCAN_IN), .Y(n2561));
  NAND3X1 g1531(.A(n2536), .B(n2111), .C(DATAI_2_), .Y(n2562));
  NAND4X1 g1532(.A(n2111), .B(n2119), .C(DATAI_26_), .D(n2525), .Y(n2563));
  AOI22X1 g1533(.A0(n2521), .A1(n2328), .B0(n2327), .B1(n2469), .Y(n2564));
  NAND4X1 g1534(.A(n2563), .B(n2562), .C(n2561), .D(n2564), .Y(U3110));
  NAND2X1 g1535(.A(n2532), .B(INSTQUEUE_REG_11__1__SCAN_IN), .Y(n2566));
  NAND3X1 g1536(.A(n2536), .B(n2111), .C(DATAI_1_), .Y(n2567));
  NAND4X1 g1537(.A(n2111), .B(n2119), .C(DATAI_25_), .D(n2525), .Y(n2568));
  AOI22X1 g1538(.A0(n2521), .A1(n2336), .B0(n2335), .B1(n2469), .Y(n2569));
  NAND4X1 g1539(.A(n2568), .B(n2567), .C(n2566), .D(n2569), .Y(U3109));
  NAND2X1 g1540(.A(n2532), .B(INSTQUEUE_REG_11__0__SCAN_IN), .Y(n2571));
  NAND3X1 g1541(.A(n2536), .B(n2111), .C(DATAI_0_), .Y(n2572));
  NAND4X1 g1542(.A(n2111), .B(n2119), .C(DATAI_24_), .D(n2525), .Y(n2573));
  AOI22X1 g1543(.A0(n2521), .A1(n2344), .B0(n2343), .B1(n2469), .Y(n2574));
  NAND4X1 g1544(.A(n2573), .B(n2572), .C(n2571), .D(n2574), .Y(U3108));
  NOR4X1  g1545(.A(n1228), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C(n1220), .D(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Y(n2576));
  AOI21X1 g1546(.A0(n2523), .A1(n2348), .B0(n2576), .Y(n2577));
  NOR4X1  g1547(.A(n2468), .B(n2354), .C(n2270), .D(n2268), .Y(n2578));
  NOR3X1  g1548(.A(n2525), .B(n2578), .C(n2120), .Y(n2580));
  OAI21X1 g1549(.A0(n2580), .A1(n2118), .B0(n2577), .Y(n2581));
  INVX1   g1550(.A(n1951), .Y(n2582));
  NOR3X1  g1551(.A(n1983), .B(n2582), .C(n1908), .Y(n2583));
  OAI22X1 g1552(.A0(n2576), .A1(n1216), .B0(n1833), .B1(n2583), .Y(n2584));
  NOR2X1  g1553(.A(n2584), .B(n2287), .Y(n2585));
  NAND2X1 g1554(.A(n2585), .B(n2581), .Y(n2586));
  NAND2X1 g1555(.A(n2586), .B(INSTQUEUE_REG_10__7__SCAN_IN), .Y(n2587));
  NAND4X1 g1556(.A(n1951), .B(n2361), .C(STATE2_REG_2__SCAN_IN), .D(n1984), .Y(n2588));
  NOR3X1  g1557(.A(n2525), .B(n2578), .C(n2279), .Y(n2589));
  NOR2X1  g1558(.A(n2589), .B(n2118), .Y(n2590));
  OAI21X1 g1559(.A0(n2590), .A1(n2577), .B0(n2588), .Y(n2591));
  NAND3X1 g1560(.A(n2591), .B(n2111), .C(DATAI_7_), .Y(n2592));
  NAND4X1 g1561(.A(n2111), .B(n2119), .C(DATAI_31_), .D(n2578), .Y(n2593));
  AOI22X1 g1562(.A0(n2576), .A1(n2288), .B0(n2286), .B1(n2525), .Y(n2594));
  NAND4X1 g1563(.A(n2593), .B(n2592), .C(n2587), .D(n2594), .Y(U3107));
  NAND2X1 g1564(.A(n2586), .B(INSTQUEUE_REG_10__6__SCAN_IN), .Y(n2596));
  NAND3X1 g1565(.A(n2591), .B(n2111), .C(DATAI_6_), .Y(n2597));
  NAND4X1 g1566(.A(n2111), .B(n2119), .C(DATAI_30_), .D(n2578), .Y(n2598));
  AOI22X1 g1567(.A0(n2576), .A1(n2296), .B0(n2295), .B1(n2525), .Y(n2599));
  NAND4X1 g1568(.A(n2598), .B(n2597), .C(n2596), .D(n2599), .Y(U3106));
  NAND2X1 g1569(.A(n2586), .B(INSTQUEUE_REG_10__5__SCAN_IN), .Y(n2601));
  NAND3X1 g1570(.A(n2591), .B(n2111), .C(DATAI_5_), .Y(n2602));
  NAND4X1 g1571(.A(n2111), .B(n2119), .C(DATAI_29_), .D(n2578), .Y(n2603));
  AOI22X1 g1572(.A0(n2576), .A1(n2304), .B0(n2303), .B1(n2525), .Y(n2604));
  NAND4X1 g1573(.A(n2603), .B(n2602), .C(n2601), .D(n2604), .Y(U3105));
  NAND2X1 g1574(.A(n2586), .B(INSTQUEUE_REG_10__4__SCAN_IN), .Y(n2606));
  NAND3X1 g1575(.A(n2591), .B(n2111), .C(DATAI_4_), .Y(n2607));
  NAND4X1 g1576(.A(n2111), .B(n2119), .C(DATAI_28_), .D(n2578), .Y(n2608));
  AOI22X1 g1577(.A0(n2576), .A1(n2312), .B0(n2311), .B1(n2525), .Y(n2609));
  NAND4X1 g1578(.A(n2608), .B(n2607), .C(n2606), .D(n2609), .Y(U3104));
  NAND2X1 g1579(.A(n2586), .B(INSTQUEUE_REG_10__3__SCAN_IN), .Y(n2611));
  NAND3X1 g1580(.A(n2591), .B(n2111), .C(DATAI_3_), .Y(n2612));
  NAND4X1 g1581(.A(n2111), .B(n2119), .C(DATAI_27_), .D(n2578), .Y(n2613));
  AOI22X1 g1582(.A0(n2576), .A1(n2320), .B0(n2319), .B1(n2525), .Y(n2614));
  NAND4X1 g1583(.A(n2613), .B(n2612), .C(n2611), .D(n2614), .Y(U3103));
  NAND2X1 g1584(.A(n2586), .B(INSTQUEUE_REG_10__2__SCAN_IN), .Y(n2616));
  NAND3X1 g1585(.A(n2591), .B(n2111), .C(DATAI_2_), .Y(n2617));
  NAND4X1 g1586(.A(n2111), .B(n2119), .C(DATAI_26_), .D(n2578), .Y(n2618));
  AOI22X1 g1587(.A0(n2576), .A1(n2328), .B0(n2327), .B1(n2525), .Y(n2619));
  NAND4X1 g1588(.A(n2618), .B(n2617), .C(n2616), .D(n2619), .Y(U3102));
  NAND2X1 g1589(.A(n2586), .B(INSTQUEUE_REG_10__1__SCAN_IN), .Y(n2621));
  NAND3X1 g1590(.A(n2591), .B(n2111), .C(DATAI_1_), .Y(n2622));
  NAND4X1 g1591(.A(n2111), .B(n2119), .C(DATAI_25_), .D(n2578), .Y(n2623));
  AOI22X1 g1592(.A0(n2576), .A1(n2336), .B0(n2335), .B1(n2525), .Y(n2624));
  NAND4X1 g1593(.A(n2623), .B(n2622), .C(n2621), .D(n2624), .Y(U3101));
  NAND2X1 g1594(.A(n2586), .B(INSTQUEUE_REG_10__0__SCAN_IN), .Y(n2626));
  NAND3X1 g1595(.A(n2591), .B(n2111), .C(DATAI_0_), .Y(n2627));
  NAND4X1 g1596(.A(n2111), .B(n2119), .C(DATAI_24_), .D(n2578), .Y(n2628));
  AOI22X1 g1597(.A0(n2576), .A1(n2344), .B0(n2343), .B1(n2525), .Y(n2629));
  NAND4X1 g1598(.A(n2628), .B(n2627), .C(n2626), .D(n2629), .Y(U3100));
  NOR4X1  g1599(.A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C(n1220), .D(n1229), .Y(n2631));
  AOI21X1 g1600(.A0(n2523), .A1(n2410), .B0(n2631), .Y(n2632));
  NOR4X1  g1601(.A(n2468), .B(n2354), .C(n2192), .D(n2268), .Y(n2633));
  NOR3X1  g1602(.A(n2578), .B(n2633), .C(n2120), .Y(n2635));
  OAI21X1 g1603(.A0(n2635), .A1(n2118), .B0(n2632), .Y(n2636));
  NOR2X1  g1604(.A(n2631), .B(n1216), .Y(n2637));
  NAND3X1 g1605(.A(n1228), .B(n1224), .C(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .Y(n2638));
  AOI21X1 g1606(.A0(n2638), .A1(STATE2_REG_2__SCAN_IN), .B0(n2637), .Y(n2639));
  NAND3X1 g1607(.A(n2639), .B(n2636), .C(n2111), .Y(n2640));
  NAND2X1 g1608(.A(n2640), .B(INSTQUEUE_REG_9__7__SCAN_IN), .Y(n2641));
  NOR3X1  g1609(.A(n2578), .B(n2633), .C(n2279), .Y(n2642));
  NOR2X1  g1610(.A(n2642), .B(n2118), .Y(n2643));
  OAI22X1 g1611(.A0(n2638), .A1(n1833), .B0(n2632), .B1(n2643), .Y(n2644));
  NAND3X1 g1612(.A(n2644), .B(n2111), .C(DATAI_7_), .Y(n2645));
  NAND4X1 g1613(.A(n2111), .B(n2119), .C(DATAI_31_), .D(n2633), .Y(n2646));
  AOI22X1 g1614(.A0(n2631), .A1(n2288), .B0(n2286), .B1(n2578), .Y(n2647));
  NAND4X1 g1615(.A(n2646), .B(n2645), .C(n2641), .D(n2647), .Y(U3099));
  NAND2X1 g1616(.A(n2640), .B(INSTQUEUE_REG_9__6__SCAN_IN), .Y(n2649));
  NAND3X1 g1617(.A(n2644), .B(n2111), .C(DATAI_6_), .Y(n2650));
  NAND4X1 g1618(.A(n2111), .B(n2119), .C(DATAI_30_), .D(n2633), .Y(n2651));
  AOI22X1 g1619(.A0(n2631), .A1(n2296), .B0(n2295), .B1(n2578), .Y(n2652));
  NAND4X1 g1620(.A(n2651), .B(n2650), .C(n2649), .D(n2652), .Y(U3098));
  NAND2X1 g1621(.A(n2640), .B(INSTQUEUE_REG_9__5__SCAN_IN), .Y(n2654));
  NAND3X1 g1622(.A(n2644), .B(n2111), .C(DATAI_5_), .Y(n2655));
  NAND4X1 g1623(.A(n2111), .B(n2119), .C(DATAI_29_), .D(n2633), .Y(n2656));
  AOI22X1 g1624(.A0(n2631), .A1(n2304), .B0(n2303), .B1(n2578), .Y(n2657));
  NAND4X1 g1625(.A(n2656), .B(n2655), .C(n2654), .D(n2657), .Y(U3097));
  NAND2X1 g1626(.A(n2640), .B(INSTQUEUE_REG_9__4__SCAN_IN), .Y(n2659));
  NAND3X1 g1627(.A(n2644), .B(n2111), .C(DATAI_4_), .Y(n2660));
  NAND4X1 g1628(.A(n2111), .B(n2119), .C(DATAI_28_), .D(n2633), .Y(n2661));
  AOI22X1 g1629(.A0(n2631), .A1(n2312), .B0(n2311), .B1(n2578), .Y(n2662));
  NAND4X1 g1630(.A(n2661), .B(n2660), .C(n2659), .D(n2662), .Y(U3096));
  NAND2X1 g1631(.A(n2640), .B(INSTQUEUE_REG_9__3__SCAN_IN), .Y(n2664));
  NAND3X1 g1632(.A(n2644), .B(n2111), .C(DATAI_3_), .Y(n2665));
  NAND4X1 g1633(.A(n2111), .B(n2119), .C(DATAI_27_), .D(n2633), .Y(n2666));
  AOI22X1 g1634(.A0(n2631), .A1(n2320), .B0(n2319), .B1(n2578), .Y(n2667));
  NAND4X1 g1635(.A(n2666), .B(n2665), .C(n2664), .D(n2667), .Y(U3095));
  NAND2X1 g1636(.A(n2640), .B(INSTQUEUE_REG_9__2__SCAN_IN), .Y(n2669));
  NAND3X1 g1637(.A(n2644), .B(n2111), .C(DATAI_2_), .Y(n2670));
  NAND4X1 g1638(.A(n2111), .B(n2119), .C(DATAI_26_), .D(n2633), .Y(n2671));
  AOI22X1 g1639(.A0(n2631), .A1(n2328), .B0(n2327), .B1(n2578), .Y(n2672));
  NAND4X1 g1640(.A(n2671), .B(n2670), .C(n2669), .D(n2672), .Y(U3094));
  NAND2X1 g1641(.A(n2640), .B(INSTQUEUE_REG_9__1__SCAN_IN), .Y(n2674));
  NAND3X1 g1642(.A(n2644), .B(n2111), .C(DATAI_1_), .Y(n2675));
  NAND4X1 g1643(.A(n2111), .B(n2119), .C(DATAI_25_), .D(n2633), .Y(n2676));
  AOI22X1 g1644(.A0(n2631), .A1(n2336), .B0(n2335), .B1(n2578), .Y(n2677));
  NAND4X1 g1645(.A(n2676), .B(n2675), .C(n2674), .D(n2677), .Y(U3093));
  NAND2X1 g1646(.A(n2640), .B(INSTQUEUE_REG_9__0__SCAN_IN), .Y(n2679));
  NAND3X1 g1647(.A(n2644), .B(n2111), .C(DATAI_0_), .Y(n2680));
  NAND4X1 g1648(.A(n2111), .B(n2119), .C(DATAI_24_), .D(n2633), .Y(n2681));
  AOI22X1 g1649(.A0(n2631), .A1(n2344), .B0(n2343), .B1(n2578), .Y(n2682));
  NAND4X1 g1650(.A(n2681), .B(n2680), .C(n2679), .D(n2682), .Y(U3092));
  NOR4X1  g1651(.A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C(n1220), .D(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Y(n2684));
  AOI21X1 g1652(.A0(n2523), .A1(n2465), .B0(n2684), .Y(n2685));
  XOR2X1  g1653(.A(n2260), .B(n2167), .Y(n2686));
  XOR2X1  g1654(.A(n2686), .B(n2257), .Y(n2687));
  XOR2X1  g1655(.A(n2267), .B(n2687), .Y(n2688));
  NOR4X1  g1656(.A(n2244), .B(n2218), .C(n2270), .D(n2688), .Y(n2689));
  NOR3X1  g1657(.A(n2633), .B(n2689), .C(n2120), .Y(n2691));
  OAI21X1 g1658(.A0(n2691), .A1(n2118), .B0(n2685), .Y(n2692));
  NOR3X1  g1659(.A(n1983), .B(n2582), .C(n2361), .Y(n2693));
  OAI22X1 g1660(.A0(n2684), .A1(n1216), .B0(n1833), .B1(n2693), .Y(n2694));
  NOR2X1  g1661(.A(n2694), .B(n2287), .Y(n2695));
  NAND2X1 g1662(.A(n2695), .B(n2692), .Y(n2696));
  NAND2X1 g1663(.A(n2696), .B(INSTQUEUE_REG_8__7__SCAN_IN), .Y(n2697));
  NAND4X1 g1664(.A(n1951), .B(n1908), .C(STATE2_REG_2__SCAN_IN), .D(n1984), .Y(n2698));
  NOR3X1  g1665(.A(n2633), .B(n2689), .C(n2279), .Y(n2699));
  NOR2X1  g1666(.A(n2699), .B(n2118), .Y(n2700));
  OAI21X1 g1667(.A0(n2700), .A1(n2685), .B0(n2698), .Y(n2701));
  NAND3X1 g1668(.A(n2701), .B(n2111), .C(DATAI_7_), .Y(n2702));
  NAND4X1 g1669(.A(n2111), .B(n2119), .C(DATAI_31_), .D(n2689), .Y(n2703));
  AOI22X1 g1670(.A0(n2684), .A1(n2288), .B0(n2286), .B1(n2633), .Y(n2704));
  NAND4X1 g1671(.A(n2703), .B(n2702), .C(n2697), .D(n2704), .Y(U3091));
  NAND2X1 g1672(.A(n2696), .B(INSTQUEUE_REG_8__6__SCAN_IN), .Y(n2706));
  NAND3X1 g1673(.A(n2701), .B(n2111), .C(DATAI_6_), .Y(n2707));
  NAND4X1 g1674(.A(n2111), .B(n2119), .C(DATAI_30_), .D(n2689), .Y(n2708));
  AOI22X1 g1675(.A0(n2684), .A1(n2296), .B0(n2295), .B1(n2633), .Y(n2709));
  NAND4X1 g1676(.A(n2708), .B(n2707), .C(n2706), .D(n2709), .Y(U3090));
  NAND2X1 g1677(.A(n2696), .B(INSTQUEUE_REG_8__5__SCAN_IN), .Y(n2711));
  NAND3X1 g1678(.A(n2701), .B(n2111), .C(DATAI_5_), .Y(n2712));
  NAND4X1 g1679(.A(n2111), .B(n2119), .C(DATAI_29_), .D(n2689), .Y(n2713));
  AOI22X1 g1680(.A0(n2684), .A1(n2304), .B0(n2303), .B1(n2633), .Y(n2714));
  NAND4X1 g1681(.A(n2713), .B(n2712), .C(n2711), .D(n2714), .Y(U3089));
  NAND2X1 g1682(.A(n2696), .B(INSTQUEUE_REG_8__4__SCAN_IN), .Y(n2716));
  NAND3X1 g1683(.A(n2701), .B(n2111), .C(DATAI_4_), .Y(n2717));
  NAND4X1 g1684(.A(n2111), .B(n2119), .C(DATAI_28_), .D(n2689), .Y(n2718));
  AOI22X1 g1685(.A0(n2684), .A1(n2312), .B0(n2311), .B1(n2633), .Y(n2719));
  NAND4X1 g1686(.A(n2718), .B(n2717), .C(n2716), .D(n2719), .Y(U3088));
  NAND2X1 g1687(.A(n2696), .B(INSTQUEUE_REG_8__3__SCAN_IN), .Y(n2721));
  NAND3X1 g1688(.A(n2701), .B(n2111), .C(DATAI_3_), .Y(n2722));
  NAND4X1 g1689(.A(n2111), .B(n2119), .C(DATAI_27_), .D(n2689), .Y(n2723));
  AOI22X1 g1690(.A0(n2684), .A1(n2320), .B0(n2319), .B1(n2633), .Y(n2724));
  NAND4X1 g1691(.A(n2723), .B(n2722), .C(n2721), .D(n2724), .Y(U3087));
  NAND2X1 g1692(.A(n2696), .B(INSTQUEUE_REG_8__2__SCAN_IN), .Y(n2726));
  NAND3X1 g1693(.A(n2701), .B(n2111), .C(DATAI_2_), .Y(n2727));
  NAND4X1 g1694(.A(n2111), .B(n2119), .C(DATAI_26_), .D(n2689), .Y(n2728));
  AOI22X1 g1695(.A0(n2684), .A1(n2328), .B0(n2327), .B1(n2633), .Y(n2729));
  NAND4X1 g1696(.A(n2728), .B(n2727), .C(n2726), .D(n2729), .Y(U3086));
  NAND2X1 g1697(.A(n2696), .B(INSTQUEUE_REG_8__1__SCAN_IN), .Y(n2731));
  NAND3X1 g1698(.A(n2701), .B(n2111), .C(DATAI_1_), .Y(n2732));
  NAND4X1 g1699(.A(n2111), .B(n2119), .C(DATAI_25_), .D(n2689), .Y(n2733));
  AOI22X1 g1700(.A0(n2684), .A1(n2336), .B0(n2335), .B1(n2633), .Y(n2734));
  NAND4X1 g1701(.A(n2733), .B(n2732), .C(n2731), .D(n2734), .Y(U3085));
  NAND2X1 g1702(.A(n2696), .B(INSTQUEUE_REG_8__0__SCAN_IN), .Y(n2736));
  NAND3X1 g1703(.A(n2701), .B(n2111), .C(DATAI_0_), .Y(n2737));
  NAND4X1 g1704(.A(n2111), .B(n2119), .C(DATAI_24_), .D(n2689), .Y(n2738));
  AOI22X1 g1705(.A0(n2684), .A1(n2344), .B0(n2343), .B1(n2633), .Y(n2739));
  NAND4X1 g1706(.A(n2738), .B(n2737), .C(n2736), .D(n2739), .Y(U3084));
  NOR2X1  g1707(.A(n1988), .B(n1958), .Y(n2741));
  AOI21X1 g1708(.A0(n2741), .A1(n2116), .B0(n1981), .Y(n2742));
  NOR4X1  g1709(.A(n2244), .B(n2218), .C(n2192), .D(n2688), .Y(n2744));
  NOR3X1  g1710(.A(n2744), .B(n2689), .C(n2120), .Y(n2745));
  OAI21X1 g1711(.A0(n2745), .A1(n2118), .B0(n2742), .Y(n2746));
  NOR2X1  g1712(.A(n1981), .B(n1216), .Y(n2747));
  NAND3X1 g1713(.A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C(n1220), .Y(n2748));
  AOI21X1 g1714(.A0(n2748), .A1(STATE2_REG_2__SCAN_IN), .B0(n2747), .Y(n2749));
  NAND3X1 g1715(.A(n2749), .B(n2746), .C(n2111), .Y(n2750));
  NAND2X1 g1716(.A(n2750), .B(INSTQUEUE_REG_7__7__SCAN_IN), .Y(n2751));
  NOR3X1  g1717(.A(n2744), .B(n2689), .C(n2279), .Y(n2752));
  NOR2X1  g1718(.A(n2752), .B(n2118), .Y(n2753));
  OAI22X1 g1719(.A0(n2748), .A1(n1833), .B0(n2742), .B1(n2753), .Y(n2754));
  NAND3X1 g1720(.A(n2754), .B(n2111), .C(DATAI_7_), .Y(n2755));
  NAND4X1 g1721(.A(n2111), .B(n2119), .C(DATAI_31_), .D(n2744), .Y(n2756));
  AOI22X1 g1722(.A0(n2286), .A1(n2689), .B0(n1981), .B1(n2288), .Y(n2757));
  NAND4X1 g1723(.A(n2756), .B(n2755), .C(n2751), .D(n2757), .Y(U3083));
  NAND2X1 g1724(.A(n2750), .B(INSTQUEUE_REG_7__6__SCAN_IN), .Y(n2759));
  NAND3X1 g1725(.A(n2754), .B(n2111), .C(DATAI_6_), .Y(n2760));
  NAND4X1 g1726(.A(n2111), .B(n2119), .C(DATAI_30_), .D(n2744), .Y(n2761));
  AOI22X1 g1727(.A0(n2295), .A1(n2689), .B0(n1981), .B1(n2296), .Y(n2762));
  NAND4X1 g1728(.A(n2761), .B(n2760), .C(n2759), .D(n2762), .Y(U3082));
  NAND2X1 g1729(.A(n2750), .B(INSTQUEUE_REG_7__5__SCAN_IN), .Y(n2764));
  NAND3X1 g1730(.A(n2754), .B(n2111), .C(DATAI_5_), .Y(n2765));
  NAND4X1 g1731(.A(n2111), .B(n2119), .C(DATAI_29_), .D(n2744), .Y(n2766));
  AOI22X1 g1732(.A0(n2303), .A1(n2689), .B0(n1981), .B1(n2304), .Y(n2767));
  NAND4X1 g1733(.A(n2766), .B(n2765), .C(n2764), .D(n2767), .Y(U3081));
  NAND2X1 g1734(.A(n2750), .B(INSTQUEUE_REG_7__4__SCAN_IN), .Y(n2769));
  NAND3X1 g1735(.A(n2754), .B(n2111), .C(DATAI_4_), .Y(n2770));
  NAND4X1 g1736(.A(n2111), .B(n2119), .C(DATAI_28_), .D(n2744), .Y(n2771));
  AOI22X1 g1737(.A0(n2311), .A1(n2689), .B0(n1981), .B1(n2312), .Y(n2772));
  NAND4X1 g1738(.A(n2771), .B(n2770), .C(n2769), .D(n2772), .Y(U3080));
  NAND2X1 g1739(.A(n2750), .B(INSTQUEUE_REG_7__3__SCAN_IN), .Y(n2774));
  NAND3X1 g1740(.A(n2754), .B(n2111), .C(DATAI_3_), .Y(n2775));
  NAND4X1 g1741(.A(n2111), .B(n2119), .C(DATAI_27_), .D(n2744), .Y(n2776));
  AOI22X1 g1742(.A0(n2319), .A1(n2689), .B0(n1981), .B1(n2320), .Y(n2777));
  NAND4X1 g1743(.A(n2776), .B(n2775), .C(n2774), .D(n2777), .Y(U3079));
  NAND2X1 g1744(.A(n2750), .B(INSTQUEUE_REG_7__2__SCAN_IN), .Y(n2779));
  NAND3X1 g1745(.A(n2754), .B(n2111), .C(DATAI_2_), .Y(n2780));
  NAND4X1 g1746(.A(n2111), .B(n2119), .C(DATAI_26_), .D(n2744), .Y(n2781));
  AOI22X1 g1747(.A0(n2327), .A1(n2689), .B0(n1981), .B1(n2328), .Y(n2782));
  NAND4X1 g1748(.A(n2781), .B(n2780), .C(n2779), .D(n2782), .Y(U3078));
  NAND2X1 g1749(.A(n2750), .B(INSTQUEUE_REG_7__1__SCAN_IN), .Y(n2784));
  NAND3X1 g1750(.A(n2754), .B(n2111), .C(DATAI_1_), .Y(n2785));
  NAND4X1 g1751(.A(n2111), .B(n2119), .C(DATAI_25_), .D(n2744), .Y(n2786));
  AOI22X1 g1752(.A0(n2335), .A1(n2689), .B0(n1981), .B1(n2336), .Y(n2787));
  NAND4X1 g1753(.A(n2786), .B(n2785), .C(n2784), .D(n2787), .Y(U3077));
  NAND2X1 g1754(.A(n2750), .B(INSTQUEUE_REG_7__0__SCAN_IN), .Y(n2789));
  NAND3X1 g1755(.A(n2754), .B(n2111), .C(DATAI_0_), .Y(n2790));
  NAND4X1 g1756(.A(n2111), .B(n2119), .C(DATAI_24_), .D(n2744), .Y(n2791));
  AOI22X1 g1757(.A0(n2343), .A1(n2689), .B0(n1981), .B1(n2344), .Y(n2792));
  NAND4X1 g1758(.A(n2791), .B(n2790), .C(n2789), .D(n2792), .Y(U3076));
  NOR4X1  g1759(.A(n1228), .B(n1224), .C(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .D(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Y(n2794));
  AOI21X1 g1760(.A0(n2741), .A1(n2348), .B0(n2794), .Y(n2795));
  NOR4X1  g1761(.A(n2244), .B(n2354), .C(n2270), .D(n2688), .Y(n2796));
  NOR3X1  g1762(.A(n2744), .B(n2796), .C(n2120), .Y(n2798));
  OAI21X1 g1763(.A0(n2798), .A1(n2118), .B0(n2795), .Y(n2799));
  NOR2X1  g1764(.A(n2794), .B(n1216), .Y(n2800));
  NOR4X1  g1765(.A(n1981), .B(n1980), .C(n1951), .D(n1982), .Y(n2801));
  NAND2X1 g1766(.A(n2801), .B(n2361), .Y(n2802));
  AOI21X1 g1767(.A0(n2802), .A1(STATE2_REG_2__SCAN_IN), .B0(n2800), .Y(n2803));
  NAND3X1 g1768(.A(n2803), .B(n2799), .C(n2111), .Y(n2804));
  NAND2X1 g1769(.A(n2804), .B(INSTQUEUE_REG_6__7__SCAN_IN), .Y(n2805));
  NOR3X1  g1770(.A(n2744), .B(n2796), .C(n2279), .Y(n2806));
  NOR2X1  g1771(.A(n2806), .B(n2118), .Y(n2807));
  OAI22X1 g1772(.A0(n2802), .A1(n1833), .B0(n2795), .B1(n2807), .Y(n2808));
  NAND3X1 g1773(.A(n2808), .B(n2111), .C(DATAI_7_), .Y(n2809));
  NAND4X1 g1774(.A(n2111), .B(n2119), .C(DATAI_31_), .D(n2796), .Y(n2810));
  AOI22X1 g1775(.A0(n2794), .A1(n2288), .B0(n2286), .B1(n2744), .Y(n2811));
  NAND4X1 g1776(.A(n2810), .B(n2809), .C(n2805), .D(n2811), .Y(U3075));
  NAND2X1 g1777(.A(n2804), .B(INSTQUEUE_REG_6__6__SCAN_IN), .Y(n2813));
  NAND3X1 g1778(.A(n2808), .B(n2111), .C(DATAI_6_), .Y(n2814));
  NAND4X1 g1779(.A(n2111), .B(n2119), .C(DATAI_30_), .D(n2796), .Y(n2815));
  AOI22X1 g1780(.A0(n2794), .A1(n2296), .B0(n2295), .B1(n2744), .Y(n2816));
  NAND4X1 g1781(.A(n2815), .B(n2814), .C(n2813), .D(n2816), .Y(U3074));
  NAND2X1 g1782(.A(n2804), .B(INSTQUEUE_REG_6__5__SCAN_IN), .Y(n2818));
  NAND3X1 g1783(.A(n2808), .B(n2111), .C(DATAI_5_), .Y(n2819));
  NAND4X1 g1784(.A(n2111), .B(n2119), .C(DATAI_29_), .D(n2796), .Y(n2820));
  AOI22X1 g1785(.A0(n2794), .A1(n2304), .B0(n2303), .B1(n2744), .Y(n2821));
  NAND4X1 g1786(.A(n2820), .B(n2819), .C(n2818), .D(n2821), .Y(U3073));
  NAND2X1 g1787(.A(n2804), .B(INSTQUEUE_REG_6__4__SCAN_IN), .Y(n2823));
  NAND3X1 g1788(.A(n2808), .B(n2111), .C(DATAI_4_), .Y(n2824));
  NAND4X1 g1789(.A(n2111), .B(n2119), .C(DATAI_28_), .D(n2796), .Y(n2825));
  AOI22X1 g1790(.A0(n2794), .A1(n2312), .B0(n2311), .B1(n2744), .Y(n2826));
  NAND4X1 g1791(.A(n2825), .B(n2824), .C(n2823), .D(n2826), .Y(U3072));
  NAND2X1 g1792(.A(n2804), .B(INSTQUEUE_REG_6__3__SCAN_IN), .Y(n2828));
  NAND3X1 g1793(.A(n2808), .B(n2111), .C(DATAI_3_), .Y(n2829));
  NAND4X1 g1794(.A(n2111), .B(n2119), .C(DATAI_27_), .D(n2796), .Y(n2830));
  AOI22X1 g1795(.A0(n2794), .A1(n2320), .B0(n2319), .B1(n2744), .Y(n2831));
  NAND4X1 g1796(.A(n2830), .B(n2829), .C(n2828), .D(n2831), .Y(U3071));
  NAND2X1 g1797(.A(n2804), .B(INSTQUEUE_REG_6__2__SCAN_IN), .Y(n2833));
  NAND3X1 g1798(.A(n2808), .B(n2111), .C(DATAI_2_), .Y(n2834));
  NAND4X1 g1799(.A(n2111), .B(n2119), .C(DATAI_26_), .D(n2796), .Y(n2835));
  AOI22X1 g1800(.A0(n2794), .A1(n2328), .B0(n2327), .B1(n2744), .Y(n2836));
  NAND4X1 g1801(.A(n2835), .B(n2834), .C(n2833), .D(n2836), .Y(U3070));
  NAND2X1 g1802(.A(n2804), .B(INSTQUEUE_REG_6__1__SCAN_IN), .Y(n2838));
  NAND3X1 g1803(.A(n2808), .B(n2111), .C(DATAI_1_), .Y(n2839));
  NAND4X1 g1804(.A(n2111), .B(n2119), .C(DATAI_25_), .D(n2796), .Y(n2840));
  AOI22X1 g1805(.A0(n2794), .A1(n2336), .B0(n2335), .B1(n2744), .Y(n2841));
  NAND4X1 g1806(.A(n2840), .B(n2839), .C(n2838), .D(n2841), .Y(U3069));
  NAND2X1 g1807(.A(n2804), .B(INSTQUEUE_REG_6__0__SCAN_IN), .Y(n2843));
  NAND3X1 g1808(.A(n2808), .B(n2111), .C(DATAI_0_), .Y(n2844));
  NAND4X1 g1809(.A(n2111), .B(n2119), .C(DATAI_24_), .D(n2796), .Y(n2845));
  AOI22X1 g1810(.A0(n2794), .A1(n2344), .B0(n2343), .B1(n2744), .Y(n2846));
  NAND4X1 g1811(.A(n2845), .B(n2844), .C(n2843), .D(n2846), .Y(U3068));
  NOR4X1  g1812(.A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n1224), .C(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .D(n1229), .Y(n2848));
  AOI21X1 g1813(.A0(n2741), .A1(n2410), .B0(n2848), .Y(n2849));
  NOR4X1  g1814(.A(n2244), .B(n2354), .C(n2192), .D(n2688), .Y(n2850));
  NOR3X1  g1815(.A(n2796), .B(n2850), .C(n2120), .Y(n2852));
  OAI21X1 g1816(.A0(n2852), .A1(n2118), .B0(n2849), .Y(n2853));
  NOR2X1  g1817(.A(n2848), .B(n1216), .Y(n2854));
  NAND3X1 g1818(.A(n1228), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C(n1220), .Y(n2855));
  AOI21X1 g1819(.A0(n2855), .A1(STATE2_REG_2__SCAN_IN), .B0(n2854), .Y(n2856));
  NAND3X1 g1820(.A(n2856), .B(n2853), .C(n2111), .Y(n2857));
  NAND2X1 g1821(.A(n2857), .B(INSTQUEUE_REG_5__7__SCAN_IN), .Y(n2858));
  NOR3X1  g1822(.A(n2796), .B(n2850), .C(n2279), .Y(n2859));
  NOR2X1  g1823(.A(n2859), .B(n2118), .Y(n2860));
  OAI22X1 g1824(.A0(n2855), .A1(n1833), .B0(n2849), .B1(n2860), .Y(n2861));
  NAND3X1 g1825(.A(n2861), .B(n2111), .C(DATAI_7_), .Y(n2862));
  NAND4X1 g1826(.A(n2111), .B(n2119), .C(DATAI_31_), .D(n2850), .Y(n2863));
  AOI22X1 g1827(.A0(n2848), .A1(n2288), .B0(n2286), .B1(n2796), .Y(n2864));
  NAND4X1 g1828(.A(n2863), .B(n2862), .C(n2858), .D(n2864), .Y(U3067));
  NAND2X1 g1829(.A(n2857), .B(INSTQUEUE_REG_5__6__SCAN_IN), .Y(n2866));
  NAND3X1 g1830(.A(n2861), .B(n2111), .C(DATAI_6_), .Y(n2867));
  NAND4X1 g1831(.A(n2111), .B(n2119), .C(DATAI_30_), .D(n2850), .Y(n2868));
  AOI22X1 g1832(.A0(n2848), .A1(n2296), .B0(n2295), .B1(n2796), .Y(n2869));
  NAND4X1 g1833(.A(n2868), .B(n2867), .C(n2866), .D(n2869), .Y(U3066));
  NAND2X1 g1834(.A(n2857), .B(INSTQUEUE_REG_5__5__SCAN_IN), .Y(n2871));
  NAND3X1 g1835(.A(n2861), .B(n2111), .C(DATAI_5_), .Y(n2872));
  NAND4X1 g1836(.A(n2111), .B(n2119), .C(DATAI_29_), .D(n2850), .Y(n2873));
  AOI22X1 g1837(.A0(n2848), .A1(n2304), .B0(n2303), .B1(n2796), .Y(n2874));
  NAND4X1 g1838(.A(n2873), .B(n2872), .C(n2871), .D(n2874), .Y(U3065));
  NAND2X1 g1839(.A(n2857), .B(INSTQUEUE_REG_5__4__SCAN_IN), .Y(n2876));
  NAND3X1 g1840(.A(n2861), .B(n2111), .C(DATAI_4_), .Y(n2877));
  NAND4X1 g1841(.A(n2111), .B(n2119), .C(DATAI_28_), .D(n2850), .Y(n2878));
  AOI22X1 g1842(.A0(n2848), .A1(n2312), .B0(n2311), .B1(n2796), .Y(n2879));
  NAND4X1 g1843(.A(n2878), .B(n2877), .C(n2876), .D(n2879), .Y(U3064));
  NAND2X1 g1844(.A(n2857), .B(INSTQUEUE_REG_5__3__SCAN_IN), .Y(n2881));
  NAND3X1 g1845(.A(n2861), .B(n2111), .C(DATAI_3_), .Y(n2882));
  NAND4X1 g1846(.A(n2111), .B(n2119), .C(DATAI_27_), .D(n2850), .Y(n2883));
  AOI22X1 g1847(.A0(n2848), .A1(n2320), .B0(n2319), .B1(n2796), .Y(n2884));
  NAND4X1 g1848(.A(n2883), .B(n2882), .C(n2881), .D(n2884), .Y(U3063));
  NAND2X1 g1849(.A(n2857), .B(INSTQUEUE_REG_5__2__SCAN_IN), .Y(n2886));
  NAND3X1 g1850(.A(n2861), .B(n2111), .C(DATAI_2_), .Y(n2887));
  NAND4X1 g1851(.A(n2111), .B(n2119), .C(DATAI_26_), .D(n2850), .Y(n2888));
  AOI22X1 g1852(.A0(n2848), .A1(n2328), .B0(n2327), .B1(n2796), .Y(n2889));
  NAND4X1 g1853(.A(n2888), .B(n2887), .C(n2886), .D(n2889), .Y(U3062));
  NAND2X1 g1854(.A(n2857), .B(INSTQUEUE_REG_5__1__SCAN_IN), .Y(n2891));
  NAND3X1 g1855(.A(n2861), .B(n2111), .C(DATAI_1_), .Y(n2892));
  NAND4X1 g1856(.A(n2111), .B(n2119), .C(DATAI_25_), .D(n2850), .Y(n2893));
  AOI22X1 g1857(.A0(n2848), .A1(n2336), .B0(n2335), .B1(n2796), .Y(n2894));
  NAND4X1 g1858(.A(n2893), .B(n2892), .C(n2891), .D(n2894), .Y(U3061));
  NAND2X1 g1859(.A(n2857), .B(INSTQUEUE_REG_5__0__SCAN_IN), .Y(n2896));
  NAND3X1 g1860(.A(n2861), .B(n2111), .C(DATAI_0_), .Y(n2897));
  NAND4X1 g1861(.A(n2111), .B(n2119), .C(DATAI_24_), .D(n2850), .Y(n2898));
  AOI22X1 g1862(.A0(n2848), .A1(n2344), .B0(n2343), .B1(n2796), .Y(n2899));
  NAND4X1 g1863(.A(n2898), .B(n2897), .C(n2896), .D(n2899), .Y(U3060));
  NOR4X1  g1864(.A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n1224), .C(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .D(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Y(n2901));
  AOI21X1 g1865(.A0(n2741), .A1(n2465), .B0(n2901), .Y(n2902));
  NOR4X1  g1866(.A(n2468), .B(n2218), .C(n2270), .D(n2688), .Y(n2903));
  NOR3X1  g1867(.A(n2850), .B(n2903), .C(n2120), .Y(n2905));
  OAI21X1 g1868(.A0(n2905), .A1(n2118), .B0(n2902), .Y(n2906));
  NOR2X1  g1869(.A(n2901), .B(n1216), .Y(n2907));
  NAND2X1 g1870(.A(n2801), .B(n1908), .Y(n2908));
  AOI21X1 g1871(.A0(n2908), .A1(STATE2_REG_2__SCAN_IN), .B0(n2907), .Y(n2909));
  NAND3X1 g1872(.A(n2909), .B(n2906), .C(n2111), .Y(n2910));
  NAND2X1 g1873(.A(n2910), .B(INSTQUEUE_REG_4__7__SCAN_IN), .Y(n2911));
  NOR3X1  g1874(.A(n2850), .B(n2903), .C(n2279), .Y(n2912));
  NOR2X1  g1875(.A(n2912), .B(n2118), .Y(n2913));
  OAI22X1 g1876(.A0(n2908), .A1(n1833), .B0(n2902), .B1(n2913), .Y(n2914));
  NAND3X1 g1877(.A(n2914), .B(n2111), .C(DATAI_7_), .Y(n2915));
  NAND4X1 g1878(.A(n2111), .B(n2119), .C(DATAI_31_), .D(n2903), .Y(n2916));
  AOI22X1 g1879(.A0(n2901), .A1(n2288), .B0(n2286), .B1(n2850), .Y(n2917));
  NAND4X1 g1880(.A(n2916), .B(n2915), .C(n2911), .D(n2917), .Y(U3059));
  NAND2X1 g1881(.A(n2910), .B(INSTQUEUE_REG_4__6__SCAN_IN), .Y(n2919));
  NAND3X1 g1882(.A(n2914), .B(n2111), .C(DATAI_6_), .Y(n2920));
  NAND4X1 g1883(.A(n2111), .B(n2119), .C(DATAI_30_), .D(n2903), .Y(n2921));
  AOI22X1 g1884(.A0(n2901), .A1(n2296), .B0(n2295), .B1(n2850), .Y(n2922));
  NAND4X1 g1885(.A(n2921), .B(n2920), .C(n2919), .D(n2922), .Y(U3058));
  NAND2X1 g1886(.A(n2910), .B(INSTQUEUE_REG_4__5__SCAN_IN), .Y(n2924));
  NAND3X1 g1887(.A(n2914), .B(n2111), .C(DATAI_5_), .Y(n2925));
  NAND4X1 g1888(.A(n2111), .B(n2119), .C(DATAI_29_), .D(n2903), .Y(n2926));
  AOI22X1 g1889(.A0(n2901), .A1(n2304), .B0(n2303), .B1(n2850), .Y(n2927));
  NAND4X1 g1890(.A(n2926), .B(n2925), .C(n2924), .D(n2927), .Y(U3057));
  NAND2X1 g1891(.A(n2910), .B(INSTQUEUE_REG_4__4__SCAN_IN), .Y(n2929));
  NAND3X1 g1892(.A(n2914), .B(n2111), .C(DATAI_4_), .Y(n2930));
  NAND4X1 g1893(.A(n2111), .B(n2119), .C(DATAI_28_), .D(n2903), .Y(n2931));
  AOI22X1 g1894(.A0(n2901), .A1(n2312), .B0(n2311), .B1(n2850), .Y(n2932));
  NAND4X1 g1895(.A(n2931), .B(n2930), .C(n2929), .D(n2932), .Y(U3056));
  NAND2X1 g1896(.A(n2910), .B(INSTQUEUE_REG_4__3__SCAN_IN), .Y(n2934));
  NAND3X1 g1897(.A(n2914), .B(n2111), .C(DATAI_3_), .Y(n2935));
  NAND4X1 g1898(.A(n2111), .B(n2119), .C(DATAI_27_), .D(n2903), .Y(n2936));
  AOI22X1 g1899(.A0(n2901), .A1(n2320), .B0(n2319), .B1(n2850), .Y(n2937));
  NAND4X1 g1900(.A(n2936), .B(n2935), .C(n2934), .D(n2937), .Y(U3055));
  NAND2X1 g1901(.A(n2910), .B(INSTQUEUE_REG_4__2__SCAN_IN), .Y(n2939));
  NAND3X1 g1902(.A(n2914), .B(n2111), .C(DATAI_2_), .Y(n2940));
  NAND4X1 g1903(.A(n2111), .B(n2119), .C(DATAI_26_), .D(n2903), .Y(n2941));
  AOI22X1 g1904(.A0(n2901), .A1(n2328), .B0(n2327), .B1(n2850), .Y(n2942));
  NAND4X1 g1905(.A(n2941), .B(n2940), .C(n2939), .D(n2942), .Y(U3054));
  NAND2X1 g1906(.A(n2910), .B(INSTQUEUE_REG_4__1__SCAN_IN), .Y(n2944));
  NAND3X1 g1907(.A(n2914), .B(n2111), .C(DATAI_1_), .Y(n2945));
  NAND4X1 g1908(.A(n2111), .B(n2119), .C(DATAI_25_), .D(n2903), .Y(n2946));
  AOI22X1 g1909(.A0(n2901), .A1(n2336), .B0(n2335), .B1(n2850), .Y(n2947));
  NAND4X1 g1910(.A(n2946), .B(n2945), .C(n2944), .D(n2947), .Y(U3053));
  NAND2X1 g1911(.A(n2910), .B(INSTQUEUE_REG_4__0__SCAN_IN), .Y(n2949));
  NAND3X1 g1912(.A(n2914), .B(n2111), .C(DATAI_0_), .Y(n2950));
  NAND4X1 g1913(.A(n2111), .B(n2119), .C(DATAI_24_), .D(n2903), .Y(n2951));
  AOI22X1 g1914(.A0(n2901), .A1(n2344), .B0(n2343), .B1(n2850), .Y(n2952));
  NAND4X1 g1915(.A(n2951), .B(n2950), .C(n2949), .D(n2952), .Y(U3052));
  NOR4X1  g1916(.A(n1228), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .D(n1229), .Y(n2954));
  NOR2X1  g1917(.A(n1988), .B(n2522), .Y(n2955));
  AOI21X1 g1918(.A0(n2955), .A1(n2116), .B0(n2954), .Y(n2956));
  NOR4X1  g1919(.A(n2468), .B(n2218), .C(n2192), .D(n2688), .Y(n2957));
  NOR3X1  g1920(.A(n2903), .B(n2957), .C(n2120), .Y(n2959));
  OAI21X1 g1921(.A0(n2959), .A1(n2118), .B0(n2956), .Y(n2960));
  NOR2X1  g1922(.A(n2954), .B(n1216), .Y(n2961));
  NAND3X1 g1923(.A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n1224), .C(n1220), .Y(n2962));
  AOI21X1 g1924(.A0(n2962), .A1(STATE2_REG_2__SCAN_IN), .B0(n2961), .Y(n2963));
  NAND3X1 g1925(.A(n2963), .B(n2960), .C(n2111), .Y(n2964));
  NAND2X1 g1926(.A(n2964), .B(INSTQUEUE_REG_3__7__SCAN_IN), .Y(n2965));
  NOR3X1  g1927(.A(n2903), .B(n2957), .C(n2279), .Y(n2966));
  NOR2X1  g1928(.A(n2966), .B(n2118), .Y(n2967));
  OAI22X1 g1929(.A0(n2962), .A1(n1833), .B0(n2956), .B1(n2967), .Y(n2968));
  NAND3X1 g1930(.A(n2968), .B(n2111), .C(DATAI_7_), .Y(n2969));
  NAND4X1 g1931(.A(n2111), .B(n2119), .C(DATAI_31_), .D(n2957), .Y(n2970));
  AOI22X1 g1932(.A0(n2954), .A1(n2288), .B0(n2286), .B1(n2903), .Y(n2971));
  NAND4X1 g1933(.A(n2970), .B(n2969), .C(n2965), .D(n2971), .Y(U3051));
  NAND2X1 g1934(.A(n2964), .B(INSTQUEUE_REG_3__6__SCAN_IN), .Y(n2973));
  NAND3X1 g1935(.A(n2968), .B(n2111), .C(DATAI_6_), .Y(n2974));
  NAND4X1 g1936(.A(n2111), .B(n2119), .C(DATAI_30_), .D(n2957), .Y(n2975));
  AOI22X1 g1937(.A0(n2954), .A1(n2296), .B0(n2295), .B1(n2903), .Y(n2976));
  NAND4X1 g1938(.A(n2975), .B(n2974), .C(n2973), .D(n2976), .Y(U3050));
  NAND2X1 g1939(.A(n2964), .B(INSTQUEUE_REG_3__5__SCAN_IN), .Y(n2978));
  NAND3X1 g1940(.A(n2968), .B(n2111), .C(DATAI_5_), .Y(n2979));
  NAND4X1 g1941(.A(n2111), .B(n2119), .C(DATAI_29_), .D(n2957), .Y(n2980));
  AOI22X1 g1942(.A0(n2954), .A1(n2304), .B0(n2303), .B1(n2903), .Y(n2981));
  NAND4X1 g1943(.A(n2980), .B(n2979), .C(n2978), .D(n2981), .Y(U3049));
  NAND2X1 g1944(.A(n2964), .B(INSTQUEUE_REG_3__4__SCAN_IN), .Y(n2983));
  NAND3X1 g1945(.A(n2968), .B(n2111), .C(DATAI_4_), .Y(n2984));
  NAND4X1 g1946(.A(n2111), .B(n2119), .C(DATAI_28_), .D(n2957), .Y(n2985));
  AOI22X1 g1947(.A0(n2954), .A1(n2312), .B0(n2311), .B1(n2903), .Y(n2986));
  NAND4X1 g1948(.A(n2985), .B(n2984), .C(n2983), .D(n2986), .Y(U3048));
  NAND2X1 g1949(.A(n2964), .B(INSTQUEUE_REG_3__3__SCAN_IN), .Y(n2988));
  NAND3X1 g1950(.A(n2968), .B(n2111), .C(DATAI_3_), .Y(n2989));
  NAND4X1 g1951(.A(n2111), .B(n2119), .C(DATAI_27_), .D(n2957), .Y(n2990));
  AOI22X1 g1952(.A0(n2954), .A1(n2320), .B0(n2319), .B1(n2903), .Y(n2991));
  NAND4X1 g1953(.A(n2990), .B(n2989), .C(n2988), .D(n2991), .Y(U3047));
  NAND2X1 g1954(.A(n2964), .B(INSTQUEUE_REG_3__2__SCAN_IN), .Y(n2993));
  NAND3X1 g1955(.A(n2968), .B(n2111), .C(DATAI_2_), .Y(n2994));
  NAND4X1 g1956(.A(n2111), .B(n2119), .C(DATAI_26_), .D(n2957), .Y(n2995));
  AOI22X1 g1957(.A0(n2954), .A1(n2328), .B0(n2327), .B1(n2903), .Y(n2996));
  NAND4X1 g1958(.A(n2995), .B(n2994), .C(n2993), .D(n2996), .Y(U3046));
  NAND2X1 g1959(.A(n2964), .B(INSTQUEUE_REG_3__1__SCAN_IN), .Y(n2998));
  NAND3X1 g1960(.A(n2968), .B(n2111), .C(DATAI_1_), .Y(n2999));
  NAND4X1 g1961(.A(n2111), .B(n2119), .C(DATAI_25_), .D(n2957), .Y(n3000));
  AOI22X1 g1962(.A0(n2954), .A1(n2336), .B0(n2335), .B1(n2903), .Y(n3001));
  NAND4X1 g1963(.A(n3000), .B(n2999), .C(n2998), .D(n3001), .Y(U3045));
  NAND2X1 g1964(.A(n2964), .B(INSTQUEUE_REG_3__0__SCAN_IN), .Y(n3003));
  NAND3X1 g1965(.A(n2968), .B(n2111), .C(DATAI_0_), .Y(n3004));
  NAND4X1 g1966(.A(n2111), .B(n2119), .C(DATAI_24_), .D(n2957), .Y(n3005));
  AOI22X1 g1967(.A0(n2954), .A1(n2344), .B0(n2343), .B1(n2903), .Y(n3006));
  NAND4X1 g1968(.A(n3005), .B(n3004), .C(n3003), .D(n3006), .Y(U3044));
  NOR4X1  g1969(.A(n1228), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .D(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Y(n3008));
  AOI21X1 g1970(.A0(n2955), .A1(n2348), .B0(n3008), .Y(n3009));
  NOR4X1  g1971(.A(n2468), .B(n2354), .C(n2270), .D(n2688), .Y(n3010));
  NOR3X1  g1972(.A(n2957), .B(n3010), .C(n2120), .Y(n3012));
  OAI21X1 g1973(.A0(n3012), .A1(n2118), .B0(n3009), .Y(n3013));
  NOR2X1  g1974(.A(n3008), .B(n1216), .Y(n3014));
  NAND3X1 g1975(.A(n1983), .B(n1951), .C(n2361), .Y(n3015));
  AOI21X1 g1976(.A0(n3015), .A1(STATE2_REG_2__SCAN_IN), .B0(n3014), .Y(n3016));
  NAND3X1 g1977(.A(n3016), .B(n3013), .C(n2111), .Y(n3017));
  NAND2X1 g1978(.A(n3017), .B(INSTQUEUE_REG_2__7__SCAN_IN), .Y(n3018));
  NOR3X1  g1979(.A(n2957), .B(n3010), .C(n2279), .Y(n3019));
  NOR2X1  g1980(.A(n3019), .B(n2118), .Y(n3020));
  OAI22X1 g1981(.A0(n3015), .A1(n1833), .B0(n3009), .B1(n3020), .Y(n3021));
  NAND3X1 g1982(.A(n3021), .B(n2111), .C(DATAI_7_), .Y(n3022));
  NAND4X1 g1983(.A(n2111), .B(n2119), .C(DATAI_31_), .D(n3010), .Y(n3023));
  AOI22X1 g1984(.A0(n3008), .A1(n2288), .B0(n2286), .B1(n2957), .Y(n3024));
  NAND4X1 g1985(.A(n3023), .B(n3022), .C(n3018), .D(n3024), .Y(U3043));
  NAND2X1 g1986(.A(n3017), .B(INSTQUEUE_REG_2__6__SCAN_IN), .Y(n3026));
  NAND3X1 g1987(.A(n3021), .B(n2111), .C(DATAI_6_), .Y(n3027));
  NAND4X1 g1988(.A(n2111), .B(n2119), .C(DATAI_30_), .D(n3010), .Y(n3028));
  AOI22X1 g1989(.A0(n3008), .A1(n2296), .B0(n2295), .B1(n2957), .Y(n3029));
  NAND4X1 g1990(.A(n3028), .B(n3027), .C(n3026), .D(n3029), .Y(U3042));
  NAND2X1 g1991(.A(n3017), .B(INSTQUEUE_REG_2__5__SCAN_IN), .Y(n3031));
  NAND3X1 g1992(.A(n3021), .B(n2111), .C(DATAI_5_), .Y(n3032));
  NAND4X1 g1993(.A(n2111), .B(n2119), .C(DATAI_29_), .D(n3010), .Y(n3033));
  AOI22X1 g1994(.A0(n3008), .A1(n2304), .B0(n2303), .B1(n2957), .Y(n3034));
  NAND4X1 g1995(.A(n3033), .B(n3032), .C(n3031), .D(n3034), .Y(U3041));
  NAND2X1 g1996(.A(n3017), .B(INSTQUEUE_REG_2__4__SCAN_IN), .Y(n3036));
  NAND3X1 g1997(.A(n3021), .B(n2111), .C(DATAI_4_), .Y(n3037));
  NAND4X1 g1998(.A(n2111), .B(n2119), .C(DATAI_28_), .D(n3010), .Y(n3038));
  AOI22X1 g1999(.A0(n3008), .A1(n2312), .B0(n2311), .B1(n2957), .Y(n3039));
  NAND4X1 g2000(.A(n3038), .B(n3037), .C(n3036), .D(n3039), .Y(U3040));
  NAND2X1 g2001(.A(n3017), .B(INSTQUEUE_REG_2__3__SCAN_IN), .Y(n3041));
  NAND3X1 g2002(.A(n3021), .B(n2111), .C(DATAI_3_), .Y(n3042));
  NAND4X1 g2003(.A(n2111), .B(n2119), .C(DATAI_27_), .D(n3010), .Y(n3043));
  AOI22X1 g2004(.A0(n3008), .A1(n2320), .B0(n2319), .B1(n2957), .Y(n3044));
  NAND4X1 g2005(.A(n3043), .B(n3042), .C(n3041), .D(n3044), .Y(U3039));
  NAND2X1 g2006(.A(n3017), .B(INSTQUEUE_REG_2__2__SCAN_IN), .Y(n3046));
  NAND3X1 g2007(.A(n3021), .B(n2111), .C(DATAI_2_), .Y(n3047));
  NAND4X1 g2008(.A(n2111), .B(n2119), .C(DATAI_26_), .D(n3010), .Y(n3048));
  AOI22X1 g2009(.A0(n3008), .A1(n2328), .B0(n2327), .B1(n2957), .Y(n3049));
  NAND4X1 g2010(.A(n3048), .B(n3047), .C(n3046), .D(n3049), .Y(U3038));
  NAND2X1 g2011(.A(n3017), .B(INSTQUEUE_REG_2__1__SCAN_IN), .Y(n3051));
  NAND3X1 g2012(.A(n3021), .B(n2111), .C(DATAI_1_), .Y(n3052));
  NAND4X1 g2013(.A(n2111), .B(n2119), .C(DATAI_25_), .D(n3010), .Y(n3053));
  AOI22X1 g2014(.A0(n3008), .A1(n2336), .B0(n2335), .B1(n2957), .Y(n3054));
  NAND4X1 g2015(.A(n3053), .B(n3052), .C(n3051), .D(n3054), .Y(U3037));
  NAND2X1 g2016(.A(n3017), .B(INSTQUEUE_REG_2__0__SCAN_IN), .Y(n3056));
  NAND3X1 g2017(.A(n3021), .B(n2111), .C(DATAI_0_), .Y(n3057));
  NAND4X1 g2018(.A(n2111), .B(n2119), .C(DATAI_24_), .D(n3010), .Y(n3058));
  AOI22X1 g2019(.A0(n3008), .A1(n2344), .B0(n2343), .B1(n2957), .Y(n3059));
  NAND4X1 g2020(.A(n3058), .B(n3057), .C(n3056), .D(n3059), .Y(U3036));
  NOR4X1  g2021(.A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .D(n1229), .Y(n3061));
  AOI21X1 g2022(.A0(n2955), .A1(n2410), .B0(n3061), .Y(n3062));
  NOR4X1  g2023(.A(n2468), .B(n2354), .C(n2192), .D(n2688), .Y(n3063));
  NOR3X1  g2024(.A(n3010), .B(n3063), .C(n2120), .Y(n3065));
  OAI21X1 g2025(.A0(n3065), .A1(n2118), .B0(n3062), .Y(n3066));
  NOR2X1  g2026(.A(n3061), .B(n1216), .Y(n3067));
  NAND3X1 g2027(.A(n1228), .B(n1224), .C(n1220), .Y(n3068));
  AOI21X1 g2028(.A0(n3068), .A1(STATE2_REG_2__SCAN_IN), .B0(n3067), .Y(n3069));
  NAND3X1 g2029(.A(n3069), .B(n3066), .C(n2111), .Y(n3070));
  NAND2X1 g2030(.A(n3070), .B(INSTQUEUE_REG_1__7__SCAN_IN), .Y(n3071));
  NOR3X1  g2031(.A(n3010), .B(n3063), .C(n2279), .Y(n3072));
  NOR2X1  g2032(.A(n3072), .B(n2118), .Y(n3073));
  OAI22X1 g2033(.A0(n3068), .A1(n1833), .B0(n3062), .B1(n3073), .Y(n3074));
  NAND3X1 g2034(.A(n3074), .B(n2111), .C(DATAI_7_), .Y(n3075));
  NAND4X1 g2035(.A(n2111), .B(n2119), .C(DATAI_31_), .D(n3063), .Y(n3076));
  AOI22X1 g2036(.A0(n3061), .A1(n2288), .B0(n2286), .B1(n3010), .Y(n3077));
  NAND4X1 g2037(.A(n3076), .B(n3075), .C(n3071), .D(n3077), .Y(U3035));
  NAND2X1 g2038(.A(n3070), .B(INSTQUEUE_REG_1__6__SCAN_IN), .Y(n3079));
  NAND3X1 g2039(.A(n3074), .B(n2111), .C(DATAI_6_), .Y(n3080));
  NAND4X1 g2040(.A(n2111), .B(n2119), .C(DATAI_30_), .D(n3063), .Y(n3081));
  AOI22X1 g2041(.A0(n3061), .A1(n2296), .B0(n2295), .B1(n3010), .Y(n3082));
  NAND4X1 g2042(.A(n3081), .B(n3080), .C(n3079), .D(n3082), .Y(U3034));
  NAND2X1 g2043(.A(n3070), .B(INSTQUEUE_REG_1__5__SCAN_IN), .Y(n3084));
  NAND3X1 g2044(.A(n3074), .B(n2111), .C(DATAI_5_), .Y(n3085));
  NAND4X1 g2045(.A(n2111), .B(n2119), .C(DATAI_29_), .D(n3063), .Y(n3086));
  AOI22X1 g2046(.A0(n3061), .A1(n2304), .B0(n2303), .B1(n3010), .Y(n3087));
  NAND4X1 g2047(.A(n3086), .B(n3085), .C(n3084), .D(n3087), .Y(U3033));
  NAND2X1 g2048(.A(n3070), .B(INSTQUEUE_REG_1__4__SCAN_IN), .Y(n3089));
  NAND3X1 g2049(.A(n3074), .B(n2111), .C(DATAI_4_), .Y(n3090));
  NAND4X1 g2050(.A(n2111), .B(n2119), .C(DATAI_28_), .D(n3063), .Y(n3091));
  AOI22X1 g2051(.A0(n3061), .A1(n2312), .B0(n2311), .B1(n3010), .Y(n3092));
  NAND4X1 g2052(.A(n3091), .B(n3090), .C(n3089), .D(n3092), .Y(U3032));
  NAND2X1 g2053(.A(n3070), .B(INSTQUEUE_REG_1__3__SCAN_IN), .Y(n3094));
  NAND3X1 g2054(.A(n3074), .B(n2111), .C(DATAI_3_), .Y(n3095));
  NAND4X1 g2055(.A(n2111), .B(n2119), .C(DATAI_27_), .D(n3063), .Y(n3096));
  AOI22X1 g2056(.A0(n3061), .A1(n2320), .B0(n2319), .B1(n3010), .Y(n3097));
  NAND4X1 g2057(.A(n3096), .B(n3095), .C(n3094), .D(n3097), .Y(U3031));
  NAND2X1 g2058(.A(n3070), .B(INSTQUEUE_REG_1__2__SCAN_IN), .Y(n3099));
  NAND3X1 g2059(.A(n3074), .B(n2111), .C(DATAI_2_), .Y(n3100));
  NAND4X1 g2060(.A(n2111), .B(n2119), .C(DATAI_26_), .D(n3063), .Y(n3101));
  AOI22X1 g2061(.A0(n3061), .A1(n2328), .B0(n2327), .B1(n3010), .Y(n3102));
  NAND4X1 g2062(.A(n3101), .B(n3100), .C(n3099), .D(n3102), .Y(U3030));
  NAND2X1 g2063(.A(n3070), .B(INSTQUEUE_REG_1__1__SCAN_IN), .Y(n3104));
  NAND3X1 g2064(.A(n3074), .B(n2111), .C(DATAI_1_), .Y(n3105));
  NAND4X1 g2065(.A(n2111), .B(n2119), .C(DATAI_25_), .D(n3063), .Y(n3106));
  AOI22X1 g2066(.A0(n3061), .A1(n2336), .B0(n2335), .B1(n3010), .Y(n3107));
  NAND4X1 g2067(.A(n3106), .B(n3105), .C(n3104), .D(n3107), .Y(U3029));
  NAND2X1 g2068(.A(n3070), .B(INSTQUEUE_REG_1__0__SCAN_IN), .Y(n3109));
  NAND3X1 g2069(.A(n3074), .B(n2111), .C(DATAI_0_), .Y(n3110));
  NAND4X1 g2070(.A(n2111), .B(n2119), .C(DATAI_24_), .D(n3063), .Y(n3111));
  AOI22X1 g2071(.A0(n3061), .A1(n2344), .B0(n2343), .B1(n3010), .Y(n3112));
  NAND4X1 g2072(.A(n3111), .B(n3110), .C(n3109), .D(n3112), .Y(U3028));
  NOR4X1  g2073(.A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .D(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Y(n3114));
  AOI21X1 g2074(.A0(n2955), .A1(n2465), .B0(n3114), .Y(n3115));
  NOR3X1  g2075(.A(n3063), .B(n2271), .C(n2120), .Y(n3118));
  OAI21X1 g2076(.A0(n3118), .A1(n2118), .B0(n3115), .Y(n3119));
  NOR2X1  g2077(.A(n3114), .B(n1216), .Y(n3120));
  NAND3X1 g2078(.A(n1983), .B(n1951), .C(n1908), .Y(n3121));
  AOI21X1 g2079(.A0(n3121), .A1(STATE2_REG_2__SCAN_IN), .B0(n3120), .Y(n3122));
  NAND3X1 g2080(.A(n3122), .B(n3119), .C(n2111), .Y(n3123));
  NAND2X1 g2081(.A(n3123), .B(INSTQUEUE_REG_0__7__SCAN_IN), .Y(n3124));
  NOR3X1  g2082(.A(n3063), .B(n2271), .C(n2279), .Y(n3125));
  NOR2X1  g2083(.A(n3125), .B(n2118), .Y(n3126));
  OAI22X1 g2084(.A0(n3121), .A1(n1833), .B0(n3115), .B1(n3126), .Y(n3127));
  NAND3X1 g2085(.A(n3127), .B(n2111), .C(DATAI_7_), .Y(n3128));
  NAND4X1 g2086(.A(n2111), .B(n2119), .C(DATAI_31_), .D(n2271), .Y(n3129));
  AOI22X1 g2087(.A0(n3114), .A1(n2288), .B0(n2286), .B1(n3063), .Y(n3130));
  NAND4X1 g2088(.A(n3129), .B(n3128), .C(n3124), .D(n3130), .Y(U3027));
  NAND2X1 g2089(.A(n3123), .B(INSTQUEUE_REG_0__6__SCAN_IN), .Y(n3132));
  NAND3X1 g2090(.A(n3127), .B(n2111), .C(DATAI_6_), .Y(n3133));
  NAND4X1 g2091(.A(n2111), .B(n2119), .C(DATAI_30_), .D(n2271), .Y(n3134));
  AOI22X1 g2092(.A0(n3114), .A1(n2296), .B0(n2295), .B1(n3063), .Y(n3135));
  NAND4X1 g2093(.A(n3134), .B(n3133), .C(n3132), .D(n3135), .Y(U3026));
  NAND2X1 g2094(.A(n3123), .B(INSTQUEUE_REG_0__5__SCAN_IN), .Y(n3137));
  NAND3X1 g2095(.A(n3127), .B(n2111), .C(DATAI_5_), .Y(n3138));
  NAND4X1 g2096(.A(n2111), .B(n2119), .C(DATAI_29_), .D(n2271), .Y(n3139));
  AOI22X1 g2097(.A0(n3114), .A1(n2304), .B0(n2303), .B1(n3063), .Y(n3140));
  NAND4X1 g2098(.A(n3139), .B(n3138), .C(n3137), .D(n3140), .Y(U3025));
  NAND2X1 g2099(.A(n3123), .B(INSTQUEUE_REG_0__4__SCAN_IN), .Y(n3142));
  NAND3X1 g2100(.A(n3127), .B(n2111), .C(DATAI_4_), .Y(n3143));
  NAND4X1 g2101(.A(n2111), .B(n2119), .C(DATAI_28_), .D(n2271), .Y(n3144));
  AOI22X1 g2102(.A0(n3114), .A1(n2312), .B0(n2311), .B1(n3063), .Y(n3145));
  NAND4X1 g2103(.A(n3144), .B(n3143), .C(n3142), .D(n3145), .Y(U3024));
  NAND2X1 g2104(.A(n3123), .B(INSTQUEUE_REG_0__3__SCAN_IN), .Y(n3147));
  NAND3X1 g2105(.A(n3127), .B(n2111), .C(DATAI_3_), .Y(n3148));
  NAND4X1 g2106(.A(n2111), .B(n2119), .C(DATAI_27_), .D(n2271), .Y(n3149));
  AOI22X1 g2107(.A0(n3114), .A1(n2320), .B0(n2319), .B1(n3063), .Y(n3150));
  NAND4X1 g2108(.A(n3149), .B(n3148), .C(n3147), .D(n3150), .Y(U3023));
  NAND2X1 g2109(.A(n3123), .B(INSTQUEUE_REG_0__2__SCAN_IN), .Y(n3152));
  NAND3X1 g2110(.A(n3127), .B(n2111), .C(DATAI_2_), .Y(n3153));
  NAND4X1 g2111(.A(n2111), .B(n2119), .C(DATAI_26_), .D(n2271), .Y(n3154));
  AOI22X1 g2112(.A0(n3114), .A1(n2328), .B0(n2327), .B1(n3063), .Y(n3155));
  NAND4X1 g2113(.A(n3154), .B(n3153), .C(n3152), .D(n3155), .Y(U3022));
  NAND2X1 g2114(.A(n3123), .B(INSTQUEUE_REG_0__1__SCAN_IN), .Y(n3157));
  NAND3X1 g2115(.A(n3127), .B(n2111), .C(DATAI_1_), .Y(n3158));
  NAND4X1 g2116(.A(n2111), .B(n2119), .C(DATAI_25_), .D(n2271), .Y(n3159));
  AOI22X1 g2117(.A0(n3114), .A1(n2336), .B0(n2335), .B1(n3063), .Y(n3160));
  NAND4X1 g2118(.A(n3159), .B(n3158), .C(n3157), .D(n3160), .Y(U3021));
  NAND2X1 g2119(.A(n3123), .B(INSTQUEUE_REG_0__0__SCAN_IN), .Y(n3162));
  NAND3X1 g2120(.A(n3127), .B(n2111), .C(DATAI_0_), .Y(n3163));
  NAND4X1 g2121(.A(n2111), .B(n2119), .C(DATAI_24_), .D(n2271), .Y(n3164));
  AOI22X1 g2122(.A0(n3114), .A1(n2344), .B0(n2343), .B1(n3063), .Y(n3165));
  NAND4X1 g2123(.A(n3164), .B(n3163), .C(n3162), .D(n3165), .Y(U3020));
  NOR4X1  g2124(.A(n1910), .B(n1833), .C(n2015), .D(n1217), .Y(n3167));
  AOI21X1 g2125(.A0(n1217), .A1(STATE2_REG_3__SCAN_IN), .B0(n3167), .Y(n3168));
  OAI21X1 g2126(.A0(n2103), .A1(n1741), .B0(n3168), .Y(n3169));
  INVX1   g2127(.A(n2008), .Y(n3170));
  NAND4X1 g2128(.A(n3170), .B(n2075), .C(n1729), .D(n3169), .Y(n3171));
  OAI21X1 g2129(.A0(n3169), .A1(n1218), .B0(n3171), .Y(U3455));
  INVX1   g2130(.A(n3169), .Y(n3173));
  AOI22X1 g2131(.A0(n1999), .A1(n2075), .B0(n1995), .B1(n2108), .Y(n3174));
  NAND2X1 g2132(.A(n3173), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n3175));
  OAI21X1 g2133(.A0(n3174), .A1(n3173), .B0(n3175), .Y(U3456));
  NOR3X1  g2134(.A(n1962), .B(n2032), .C(n1216), .Y(n3177));
  INVX1   g2135(.A(n2075), .Y(n3178));
  OAI22X1 g2136(.A0(n2018), .A1(n2023), .B0(n1970), .B1(n3178), .Y(n3179));
  OAI21X1 g2137(.A0(n3179), .A1(n3177), .B0(n3169), .Y(n3180));
  OAI21X1 g2138(.A0(n3169), .A1(n1226), .B0(n3180), .Y(U3459));
  NOR4X1  g2139(.A(n1544), .B(n1250), .C(n1216), .D(n2032), .Y(n3182));
  OAI21X1 g2140(.A0(n1941), .A1(n3178), .B0(n2089), .Y(n3183));
  OAI21X1 g2141(.A0(n3183), .A1(n3182), .B0(n3169), .Y(n3184));
  OAI21X1 g2142(.A0(n3169), .A1(n1245), .B0(n3184), .Y(U3460));
  NOR2X1  g2143(.A(INSTADDRPOINTER_REG_0__SCAN_IN), .B(n1910), .Y(n3186));
  AOI21X1 g2144(.A0(n1851), .A1(n2075), .B0(n3186), .Y(n3187));
  OAI21X1 g2145(.A0(n2109), .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B0(n3187), .Y(n3188));
  NAND2X1 g2146(.A(n3188), .B(n3169), .Y(n3189));
  OAI21X1 g2147(.A0(n3169), .A1(n1231), .B0(n3189), .Y(U3461));
  NAND3X1 g2148(.A(n2098), .B(n2086), .C(STATE2_REG_0__SCAN_IN), .Y(n3191));
  NOR2X1  g2149(.A(n3167), .B(n2111), .Y(n3192));
  NAND2X1 g2150(.A(n3192), .B(n3191), .Y(n3193));
  NOR2X1  g2151(.A(n3193), .B(n1238), .Y(U3019));
  INVX1   g2152(.A(n2744), .Y(n3195));
  NOR2X1  g2153(.A(n2218), .B(n2270), .Y(n3196));
  AOI21X1 g2154(.A0(n2468), .A1(n3196), .B0(n2268), .Y(n3197));
  NAND3X1 g2155(.A(n2468), .B(n2354), .C(n2270), .Y(n3198));
  OAI21X1 g2156(.A0(n3197), .A1(n2689), .B0(n3198), .Y(n3199));
  AOI21X1 g2157(.A0(n3199), .A1(n3195), .B0(n2279), .Y(n3200));
  INVX1   g2158(.A(n2118), .Y(n3201));
  NOR2X1  g2159(.A(n1910), .B(STATE2_REG_3__SCAN_IN), .Y(n3202));
  OAI22X1 g2160(.A0(n2268), .A1(n3201), .B0(n1989), .B1(n3202), .Y(n3203));
  OAI21X1 g2161(.A0(n3203), .A1(n3200), .B0(n3193), .Y(n3204));
  OAI21X1 g2162(.A0(n3193), .A1(n1220), .B0(n3204), .Y(U3462));
  NOR2X1  g2163(.A(n2218), .B(n2192), .Y(n3206));
  XOR2X1  g2164(.A(n2244), .B(n3196), .Y(n3207));
  XOR2X1  g2165(.A(n3207), .B(n3206), .Y(n3208));
  NOR2X1  g2166(.A(n3208), .B(n2279), .Y(n3209));
  OAI22X1 g2167(.A0(n2244), .A1(n3201), .B0(n1958), .B1(n3202), .Y(n3210));
  OAI21X1 g2168(.A0(n3210), .A1(n3209), .B0(n3193), .Y(n3211));
  OAI21X1 g2169(.A0(n3193), .A1(n1224), .B0(n3211), .Y(U3463));
  AOI21X1 g2170(.A0(n2470), .A1(n2413), .B0(n2279), .Y(n3215));
  OAI22X1 g2171(.A0(n2218), .A1(n3201), .B0(n1937), .B1(n3202), .Y(n3216));
  OAI21X1 g2172(.A0(n3216), .A1(n3215), .B0(n3193), .Y(n3217));
  OAI21X1 g2173(.A0(n3193), .A1(n1228), .B0(n3217), .Y(U3464));
  NOR2X1  g2174(.A(STATE2_REG_2__SCAN_IN), .B(STATE2_REG_3__SCAN_IN), .Y(n3219));
  INVX1   g2175(.A(n3219), .Y(n3220));
  OAI22X1 g2176(.A0(n2270), .A1(n3220), .B0(n1843), .B1(n3202), .Y(n3221));
  OAI21X1 g2177(.A0(n3221), .A1(n2099), .B0(n3193), .Y(n3222));
  OAI21X1 g2178(.A0(n3193), .A1(n1229), .B0(n3222), .Y(U3465));
  AOI22X1 g2179(.A0(n1592), .A1(n1282), .B0(n1867), .B1(n2179), .Y(n3224));
  INVX1   g2180(.A(n3224), .Y(n3225));
  AOI21X1 g2181(.A0(n2192), .A1(n1472), .B0(n3225), .Y(n3226));
  XOR2X1  g2182(.A(n3226), .B(n2016), .Y(n3227));
  OAI21X1 g2183(.A0(n2042), .A1(n2032), .B0(n1362), .Y(n3228));
  NOR3X1  g2184(.A(n2038), .B(n1720), .C(READY_N), .Y(n3229));
  NAND3X1 g2185(.A(n2034), .B(n1856), .C(n1720), .Y(n3230));
  AOI21X1 g2186(.A0(n2042), .A1(n1464), .B0(READY_N), .Y(n3231));
  NAND4X1 g2187(.A(n1824), .B(n1823), .C(n1773), .D(n3231), .Y(n3232));
  AOI21X1 g2188(.A0(n1615), .A1(n1671), .B0(n1282), .Y(n3233));
  AOI21X1 g2189(.A0(n3233), .A1(n3232), .B0(n1639), .Y(n3234));
  AOI21X1 g2190(.A0(n3234), .A1(n1536), .B0(n1728), .Y(n3235));
  NAND2X1 g2191(.A(n3235), .B(n3230), .Y(n3236));
  AOI21X1 g2192(.A0(n3229), .A1(n3228), .B0(n3236), .Y(n3237));
  NOR2X1  g2193(.A(n3237), .B(n2103), .Y(n3238));
  NOR4X1  g2194(.A(STATE2_REG_1__SCAN_IN), .B(STATE2_REG_2__SCAN_IN), .C(STATE2_REG_3__SCAN_IN), .D(STATE2_REG_0__SCAN_IN), .Y(n3239));
  AOI21X1 g2195(.A0(n1568), .A1(n1394), .B0(n1950), .Y(n3240));
  AOI21X1 g2196(.A0(n3240), .A1(n1319), .B0(n3239), .Y(n3241));
  INVX1   g2197(.A(n3241), .Y(n3242));
  NOR3X1  g2198(.A(n1683), .B(n1672), .C(n1639), .Y(n3243));
  NOR4X1  g2199(.A(n1464), .B(n1282), .C(n1833), .D(n1825), .Y(n3244));
  NOR3X1  g2200(.A(n3244), .B(n3243), .C(n1729), .Y(n3245));
  INVX1   g2201(.A(n1923), .Y(n3246));
  NOR4X1  g2202(.A(n1639), .B(n1655), .C(n1721), .D(n1672), .Y(n3247));
  NOR3X1  g2203(.A(n3247), .B(n3246), .C(n1679), .Y(n3248));
  AOI21X1 g2204(.A0(n3248), .A1(n3245), .B0(n1833), .Y(n3249));
  OAI21X1 g2205(.A0(n3242), .A1(n3238), .B0(n3249), .Y(n3250));
  INVX1   g2206(.A(n3250), .Y(n3251));
  INVX1   g2207(.A(REIP_REG_0__SCAN_IN), .Y(n3252));
  NOR2X1  g2208(.A(n3242), .B(n3238), .Y(n3253));
  INVX1   g2209(.A(n3253), .Y(n3254));
  OAI22X1 g2210(.A0(n3254), .A1(n2016), .B0(n3252), .B1(n5914), .Y(n3257));
  AOI21X1 g2211(.A0(n3251), .A1(n3227), .B0(n3257), .Y(n3258));
  NOR3X1  g2212(.A(n3253), .B(n1685), .C(n1833), .Y(n3259));
  NOR2X1  g2213(.A(n3253), .B(n1833), .Y(n3260));
  NOR3X1  g2214(.A(n1886), .B(n1720), .C(n1569), .Y(n3261));
  AOI21X1 g2215(.A0(n1799), .A1(n1772), .B0(n3261), .Y(n3262));
  INVX1   g2216(.A(n1779), .Y(n3263));
  AOI21X1 g2217(.A0(n1768), .A1(n1282), .B0(n3263), .Y(n3264));
  NAND4X1 g2218(.A(n3262), .B(n1966), .C(n1767), .D(n3264), .Y(n3265));
  NAND2X1 g2219(.A(n3265), .B(n3260), .Y(n3266));
  INVX1   g2220(.A(n3266), .Y(n3267));
  OAI21X1 g2221(.A0(n3267), .A1(n3259), .B0(n2016), .Y(n3268));
  NOR3X1  g2222(.A(n3253), .B(n1963), .C(n1833), .Y(n3269));
  XOR2X1  g2223(.A(n1760), .B(n1758), .Y(n3270));
  AOI21X1 g2224(.A0(n1891), .A1(n1464), .B0(n1282), .Y(n3272));
  INVX1   g2225(.A(n3272), .Y(n3273));
  AOI22X1 g2226(.A0(n3270), .A1(EBX_REG_0__SCAN_IN), .B0(INSTADDRPOINTER_REG_0__SCAN_IN), .B1(n3273), .Y(n3274));
  XOR2X1  g2227(.A(n3274), .B(n1763), .Y(n3275));
  XOR2X1  g2228(.A(n3275), .B(n3270), .Y(n3276));
  AOI21X1 g2229(.A0(n1640), .A1(n1867), .B0(n1878), .Y(n3277));
  NOR3X1  g2230(.A(n3277), .B(n3253), .C(n1833), .Y(n3278));
  AOI22X1 g2231(.A0(n3276), .A1(n3278), .B0(n3269), .B1(INSTADDRPOINTER_REG_0__SCAN_IN), .Y(n3279));
  NAND3X1 g2232(.A(n3279), .B(n3268), .C(n3258), .Y(U3018));
  NAND2X1 g2233(.A(n3269), .B(n2021), .Y(n3281));
  NOR3X1  g2234(.A(n1763), .B(n1592), .C(n1282), .Y(n3282));
  AOI21X1 g2235(.A0(n3275), .A1(n3270), .B0(n3282), .Y(n3283));
  AOI22X1 g2236(.A0(n3270), .A1(EBX_REG_1__SCAN_IN), .B0(INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n3273), .Y(n3284));
  XOR2X1  g2237(.A(n3284), .B(n1758), .Y(n3285));
  XOR2X1  g2238(.A(n3285), .B(n3273), .Y(n3286));
  XOR2X1  g2239(.A(n3286), .B(n3283), .Y(n3287));
  AOI22X1 g2240(.A0(n3278), .A1(n3287), .B0(n3259), .B1(n2020), .Y(n3288));
  NOR2X1  g2241(.A(n3226), .B(n2016), .Y(n3289));
  INVX1   g2242(.A(n2179), .Y(n3290));
  XOR2X1  g2243(.A(n2207), .B(n3290), .Y(n3291));
  NAND2X1 g2244(.A(n1720), .B(n1592), .Y(n3292));
  AOI21X1 g2245(.A0(n1422), .A1(n1447), .B0(n3292), .Y(n3293));
  OAI21X1 g2246(.A0(n3291), .A1(n1721), .B0(n3293), .Y(n3294));
  INVX1   g2247(.A(n3294), .Y(n3295));
  OAI21X1 g2248(.A0(n2218), .A1(n1473), .B0(n3295), .Y(n3296));
  XOR2X1  g2249(.A(n3296), .B(n2021), .Y(n3297));
  XOR2X1  g2250(.A(n3297), .B(n3289), .Y(n3298));
  NOR2X1  g2251(.A(n3298), .B(n3250), .Y(n3299));
  AOI22X1 g2252(.A0(n3253), .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .B0(REIP_REG_1__SCAN_IN), .B1(n3239), .Y(n3300));
  OAI21X1 g2253(.A0(n3266), .A1(n2019), .B0(n3300), .Y(n3301));
  NOR2X1  g2254(.A(n3301), .B(n3299), .Y(n3302));
  NAND3X1 g2255(.A(n3302), .B(n3288), .C(n3281), .Y(U3017));
  INVX1   g2256(.A(INSTADDRPOINTER_REG_2__SCAN_IN), .Y(n3304));
  NOR2X1  g2257(.A(n2207), .B(n2179), .Y(n3305));
  XOR2X1  g2258(.A(n3305), .B(n2230), .Y(n3306));
  OAI22X1 g2259(.A0(n1655), .A1(n1447), .B0(n1721), .B1(n3306), .Y(n3307));
  INVX1   g2260(.A(n3307), .Y(n3308));
  OAI21X1 g2261(.A0(n2244), .A1(n1473), .B0(n3308), .Y(n3309));
  XOR2X1  g2262(.A(n3309), .B(n3304), .Y(n3310));
  NAND2X1 g2263(.A(n2354), .B(n1472), .Y(n3311));
  NAND3X1 g2264(.A(n3295), .B(n3311), .C(n2021), .Y(n3312));
  AOI21X1 g2265(.A0(n3295), .A1(n3311), .B0(n2021), .Y(n3313));
  AOI21X1 g2266(.A0(n3312), .A1(n3289), .B0(n3313), .Y(n3314));
  XOR2X1  g2267(.A(n3314), .B(n3310), .Y(n3315));
  NAND2X1 g2268(.A(n3315), .B(n3251), .Y(n3316));
  NAND2X1 g2269(.A(INSTADDRPOINTER_REG_1__SCAN_IN), .B(INSTADDRPOINTER_REG_0__SCAN_IN), .Y(n3317));
  XOR2X1  g2270(.A(n3317), .B(n3304), .Y(n3318));
  OAI22X1 g2271(.A0(n3254), .A1(n3304), .B0(n1106), .B1(n5914), .Y(n3319));
  AOI21X1 g2272(.A0(n3318), .A1(n3267), .B0(n3319), .Y(n3320));
  XOR2X1  g2273(.A(INSTADDRPOINTER_REG_2__SCAN_IN), .B(INSTADDRPOINTER_REG_1__SCAN_IN), .Y(n3321));
  NAND2X1 g2274(.A(n3321), .B(n3269), .Y(n3322));
  XOR2X1  g2275(.A(n3317), .B(INSTADDRPOINTER_REG_2__SCAN_IN), .Y(n3323));
  AOI22X1 g2276(.A0(n3270), .A1(EBX_REG_2__SCAN_IN), .B0(INSTADDRPOINTER_REG_2__SCAN_IN), .B1(n3273), .Y(n3324));
  XOR2X1  g2277(.A(n3324), .B(n1758), .Y(n3325));
  INVX1   g2278(.A(n3285), .Y(n3326));
  AOI21X1 g2279(.A0(n3285), .A1(n3272), .B0(n3283), .Y(n3327));
  AOI21X1 g2280(.A0(n3326), .A1(n3273), .B0(n3327), .Y(n3328));
  XOR2X1  g2281(.A(n3328), .B(n3325), .Y(n3329));
  AOI22X1 g2282(.A0(n3323), .A1(n3259), .B0(n3278), .B1(n3329), .Y(n3330));
  NAND4X1 g2283(.A(n3322), .B(n3320), .C(n3316), .D(n3330), .Y(U3016));
  INVX1   g2284(.A(INSTADDRPOINTER_REG_3__SCAN_IN), .Y(n3332));
  NOR3X1  g2285(.A(n3305), .B(n2256), .C(n2230), .Y(n3333));
  OAI21X1 g2286(.A0(n3305), .A1(n2230), .B0(n2256), .Y(n3334));
  INVX1   g2287(.A(n3334), .Y(n3335));
  NOR3X1  g2288(.A(n3335), .B(n3333), .C(n1721), .Y(n3336));
  AOI21X1 g2289(.A0(n2688), .A1(n1472), .B0(n3336), .Y(n3337));
  XOR2X1  g2290(.A(n3337), .B(n3332), .Y(n3338));
  NOR2X1  g2291(.A(n3309), .B(INSTADDRPOINTER_REG_2__SCAN_IN), .Y(n3339));
  NAND2X1 g2292(.A(n3309), .B(INSTADDRPOINTER_REG_2__SCAN_IN), .Y(n3340));
  OAI21X1 g2293(.A0(n3314), .A1(n3339), .B0(n3340), .Y(n3341));
  XOR2X1  g2294(.A(n3341), .B(n3338), .Y(n3342));
  NAND2X1 g2295(.A(n3342), .B(n3251), .Y(n3343));
  INVX1   g2296(.A(n3259), .Y(n3344));
  AOI21X1 g2297(.A0(INSTADDRPOINTER_REG_1__SCAN_IN), .A1(INSTADDRPOINTER_REG_0__SCAN_IN), .B0(INSTADDRPOINTER_REG_2__SCAN_IN), .Y(n3345));
  XOR2X1  g2298(.A(n3345), .B(INSTADDRPOINTER_REG_3__SCAN_IN), .Y(n3346));
  AOI22X1 g2299(.A0(n3253), .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .B0(REIP_REG_3__SCAN_IN), .B1(n3239), .Y(n3347));
  OAI21X1 g2300(.A0(n3346), .A1(n3344), .B0(n3347), .Y(n3348));
  NOR2X1  g2301(.A(n3328), .B(n3325), .Y(n3349));
  AOI22X1 g2302(.A0(n3270), .A1(EBX_REG_3__SCAN_IN), .B0(INSTADDRPOINTER_REG_3__SCAN_IN), .B1(n3273), .Y(n3350));
  XOR2X1  g2303(.A(n3350), .B(n1758), .Y(n3351));
  XOR2X1  g2304(.A(n3351), .B(n3349), .Y(n3352));
  NOR4X1  g2305(.A(n3277), .B(n3253), .C(n1833), .D(n3352), .Y(n3353));
  INVX1   g2306(.A(n3269), .Y(n3354));
  NOR2X1  g2307(.A(n3317), .B(n3304), .Y(n3355));
  XOR2X1  g2308(.A(n3355), .B(n3332), .Y(n3356));
  NAND2X1 g2309(.A(INSTADDRPOINTER_REG_2__SCAN_IN), .B(INSTADDRPOINTER_REG_1__SCAN_IN), .Y(n3357));
  XOR2X1  g2310(.A(n3357), .B(INSTADDRPOINTER_REG_3__SCAN_IN), .Y(n3358));
  OAI22X1 g2311(.A0(n3356), .A1(n3266), .B0(n3354), .B1(n3358), .Y(n3359));
  NOR3X1  g2312(.A(n3359), .B(n3353), .C(n3348), .Y(n3360));
  NAND2X1 g2313(.A(n3360), .B(n3343), .Y(U3015));
  INVX1   g2314(.A(INSTADDRPOINTER_REG_4__SCAN_IN), .Y(n3362));
  AOI22X1 g2315(.A0(n1268), .A1(INSTQUEUE_REG_0__4__SCAN_IN), .B0(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n1244), .Y(n3363));
  AOI22X1 g2316(.A0(n1246), .A1(INSTQUEUE_REG_3__4__SCAN_IN), .B0(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n1337), .Y(n3364));
  AOI22X1 g2317(.A0(n1273), .A1(INSTQUEUE_REG_4__4__SCAN_IN), .B0(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n1329), .Y(n3365));
  AOI22X1 g2318(.A0(n1278), .A1(INSTQUEUE_REG_7__4__SCAN_IN), .B0(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n1270), .Y(n3366));
  NAND4X1 g2319(.A(n3365), .B(n3364), .C(n3363), .D(n3366), .Y(n3367));
  AOI22X1 g2320(.A0(n1253), .A1(INSTQUEUE_REG_12__4__SCAN_IN), .B0(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n1271), .Y(n3368));
  AOI22X1 g2321(.A0(n1279), .A1(INSTQUEUE_REG_15__4__SCAN_IN), .B0(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n1266), .Y(n3369));
  AOI22X1 g2322(.A0(n1323), .A1(INSTQUEUE_REG_8__4__SCAN_IN), .B0(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n1338), .Y(n3370));
  AOI22X1 g2323(.A0(n1255), .A1(INSTQUEUE_REG_11__4__SCAN_IN), .B0(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n1275), .Y(n3371));
  NAND4X1 g2324(.A(n3370), .B(n3369), .C(n3368), .D(n3371), .Y(n3372));
  NOR2X1  g2325(.A(n3372), .B(n3367), .Y(n3373));
  INVX1   g2326(.A(n3373), .Y(n3374));
  XOR2X1  g2327(.A(n3374), .B(n3334), .Y(n3375));
  NOR2X1  g2328(.A(n3375), .B(n1721), .Y(n3376));
  AOI22X1 g2329(.A0(n1476), .A1(n3374), .B0(n1319), .B1(INSTQUEUE_REG_0__4__SCAN_IN), .Y(n3377));
  NOR4X1  g2330(.A(n2165), .B(n1403), .C(n1217), .D(n3373), .Y(n3378));
  NOR3X1  g2331(.A(n3373), .B(n2214), .C(n2166), .Y(n3379));
  NOR2X1  g2332(.A(n3379), .B(n3378), .Y(n3380));
  XOR2X1  g2333(.A(n3380), .B(n3377), .Y(n3381));
  OAI21X1 g2334(.A0(n2240), .A1(n2212), .B0(n2353), .Y(n3382));
  AOI22X1 g2335(.A0(n2242), .A1(n3382), .B0(n2264), .B1(n2263), .Y(n3383));
  INVX1   g2336(.A(n2257), .Y(n3384));
  OAI22X1 g2337(.A0(n3384), .A1(n2261), .B0(n2264), .B1(n2263), .Y(n3385));
  OAI22X1 g2338(.A0(n3383), .A1(n3385), .B0(n2686), .B1(n2257), .Y(n3386));
  XOR2X1  g2339(.A(n3386), .B(n3381), .Y(n3387));
  AOI21X1 g2340(.A0(n3387), .A1(n1472), .B0(n3376), .Y(n3388));
  XOR2X1  g2341(.A(n3388), .B(n3362), .Y(n3389));
  INVX1   g2342(.A(n3336), .Y(n3390));
  OAI21X1 g2343(.A0(n2268), .A1(n1473), .B0(n3390), .Y(n3391));
  NOR2X1  g2344(.A(n3391), .B(INSTADDRPOINTER_REG_3__SCAN_IN), .Y(n3392));
  NAND2X1 g2345(.A(n3391), .B(INSTADDRPOINTER_REG_3__SCAN_IN), .Y(n3393));
  NAND2X1 g2346(.A(n3296), .B(INSTADDRPOINTER_REG_1__SCAN_IN), .Y(n3394));
  OAI21X1 g2347(.A0(n3296), .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .B0(n3289), .Y(n3395));
  AOI21X1 g2348(.A0(n3395), .A1(n3394), .B0(n3339), .Y(n3396));
  AOI21X1 g2349(.A0(n3309), .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .B0(n3396), .Y(n3397));
  OAI21X1 g2350(.A0(n3397), .A1(n3392), .B0(n3393), .Y(n3398));
  XOR2X1  g2351(.A(n3398), .B(n3389), .Y(n3399));
  NAND2X1 g2352(.A(n3399), .B(n3251), .Y(n3400));
  NOR2X1  g2353(.A(n3345), .B(n3332), .Y(n3401));
  XOR2X1  g2354(.A(n3401), .B(n3362), .Y(n3402));
  AOI22X1 g2355(.A0(n3253), .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .B0(REIP_REG_4__SCAN_IN), .B1(n3239), .Y(n3403));
  OAI21X1 g2356(.A0(n3402), .A1(n3344), .B0(n3403), .Y(n3404));
  NAND4X1 g2357(.A(INSTADDRPOINTER_REG_2__SCAN_IN), .B(INSTADDRPOINTER_REG_1__SCAN_IN), .C(INSTADDRPOINTER_REG_0__SCAN_IN), .D(INSTADDRPOINTER_REG_3__SCAN_IN), .Y(n3405));
  XOR2X1  g2358(.A(n3405), .B(INSTADDRPOINTER_REG_4__SCAN_IN), .Y(n3406));
  NOR2X1  g2359(.A(n3406), .B(n3266), .Y(n3407));
  INVX1   g2360(.A(n3278), .Y(n3408));
  AOI22X1 g2361(.A0(n3270), .A1(EBX_REG_4__SCAN_IN), .B0(INSTADDRPOINTER_REG_4__SCAN_IN), .B1(n3273), .Y(n3409));
  XOR2X1  g2362(.A(n3409), .B(n1763), .Y(n3410));
  INVX1   g2363(.A(n3328), .Y(n3411));
  NOR2X1  g2364(.A(n3351), .B(n3325), .Y(n3412));
  NAND2X1 g2365(.A(n3412), .B(n3411), .Y(n3413));
  XOR2X1  g2366(.A(n3413), .B(n3410), .Y(n3414));
  NAND3X1 g2367(.A(INSTADDRPOINTER_REG_3__SCAN_IN), .B(INSTADDRPOINTER_REG_2__SCAN_IN), .C(INSTADDRPOINTER_REG_1__SCAN_IN), .Y(n3415));
  XOR2X1  g2368(.A(n3415), .B(INSTADDRPOINTER_REG_4__SCAN_IN), .Y(n3416));
  OAI22X1 g2369(.A0(n3414), .A1(n3408), .B0(n3354), .B1(n3416), .Y(n3417));
  NOR3X1  g2370(.A(n3417), .B(n3407), .C(n3404), .Y(n3418));
  NAND2X1 g2371(.A(n3418), .B(n3400), .Y(U3014));
  INVX1   g2372(.A(INSTADDRPOINTER_REG_5__SCAN_IN), .Y(n3420));
  NOR2X1  g2373(.A(n3373), .B(n3334), .Y(n3421));
  AOI22X1 g2374(.A0(n1268), .A1(INSTQUEUE_REG_0__5__SCAN_IN), .B0(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n1244), .Y(n3422));
  AOI22X1 g2375(.A0(n1246), .A1(INSTQUEUE_REG_3__5__SCAN_IN), .B0(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n1337), .Y(n3423));
  AOI22X1 g2376(.A0(n1273), .A1(INSTQUEUE_REG_4__5__SCAN_IN), .B0(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n1329), .Y(n3424));
  AOI22X1 g2377(.A0(n1278), .A1(INSTQUEUE_REG_7__5__SCAN_IN), .B0(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n1270), .Y(n3425));
  NAND4X1 g2378(.A(n3424), .B(n3423), .C(n3422), .D(n3425), .Y(n3426));
  AOI22X1 g2379(.A0(n1253), .A1(INSTQUEUE_REG_12__5__SCAN_IN), .B0(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n1271), .Y(n3427));
  AOI22X1 g2380(.A0(n1279), .A1(INSTQUEUE_REG_15__5__SCAN_IN), .B0(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n1266), .Y(n3428));
  AOI22X1 g2381(.A0(n1323), .A1(INSTQUEUE_REG_8__5__SCAN_IN), .B0(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n1338), .Y(n3429));
  AOI22X1 g2382(.A0(n1255), .A1(INSTQUEUE_REG_11__5__SCAN_IN), .B0(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n1275), .Y(n3430));
  NAND4X1 g2383(.A(n3429), .B(n3428), .C(n3427), .D(n3430), .Y(n3431));
  NOR2X1  g2384(.A(n3431), .B(n3426), .Y(n3432));
  XOR2X1  g2385(.A(n3432), .B(n3421), .Y(n3433));
  NOR2X1  g2386(.A(n3433), .B(n1721), .Y(n3434));
  NOR3X1  g2387(.A(n3432), .B(n1447), .C(n1217), .Y(n3435));
  AOI21X1 g2388(.A0(n1319), .A1(INSTQUEUE_REG_0__5__SCAN_IN), .B0(n3435), .Y(n3436));
  NOR4X1  g2389(.A(n2165), .B(n1403), .C(n1217), .D(n3432), .Y(n3437));
  NOR3X1  g2390(.A(n3432), .B(n2214), .C(n2166), .Y(n3438));
  NOR2X1  g2391(.A(n3438), .B(n3437), .Y(n3439));
  XOR2X1  g2392(.A(n3439), .B(n3436), .Y(n3440));
  NAND2X1 g2393(.A(n3380), .B(n3377), .Y(n3441));
  INVX1   g2394(.A(n3441), .Y(n3442));
  AOI21X1 g2395(.A0(n2235), .A1(n2231), .B0(n3442), .Y(n3443));
  OAI21X1 g2396(.A0(n2261), .A1(n3384), .B0(n3443), .Y(n3444));
  NOR2X1  g2397(.A(n3380), .B(n3377), .Y(n3445));
  AOI21X1 g2398(.A0(n3380), .A1(n3377), .B0(n2257), .Y(n3446));
  OAI21X1 g2399(.A0(n3444), .A1(n3383), .B0(n3506), .Y(n3448));
  XOR2X1  g2400(.A(n3448), .B(n3440), .Y(n3449));
  AOI21X1 g2401(.A0(n3449), .A1(n1472), .B0(n3434), .Y(n3450));
  XOR2X1  g2402(.A(n3450), .B(n3420), .Y(n3451));
  INVX1   g2403(.A(n3451), .Y(n3452));
  NAND2X1 g2404(.A(n3388), .B(n3362), .Y(n3453));
  NOR2X1  g2405(.A(n3388), .B(n3362), .Y(n3454));
  AOI21X1 g2406(.A0(n3398), .A1(n3453), .B0(n3454), .Y(n3455));
  XOR2X1  g2407(.A(n3455), .B(n3452), .Y(n3456));
  NAND2X1 g2408(.A(n3456), .B(n3251), .Y(n3457));
  NOR3X1  g2409(.A(n3345), .B(n3362), .C(n3332), .Y(n3458));
  XOR2X1  g2410(.A(n3458), .B(n3420), .Y(n3459));
  AOI22X1 g2411(.A0(n3253), .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .B0(REIP_REG_5__SCAN_IN), .B1(n3239), .Y(n3460));
  OAI21X1 g2412(.A0(n3459), .A1(n3344), .B0(n3460), .Y(n3461));
  NOR4X1  g2413(.A(n3362), .B(n3332), .C(n3304), .D(n3317), .Y(n3462));
  XOR2X1  g2414(.A(n3462), .B(n3420), .Y(n3463));
  NOR2X1  g2415(.A(n3463), .B(n3266), .Y(n3464));
  AOI22X1 g2416(.A0(n3270), .A1(EBX_REG_5__SCAN_IN), .B0(INSTADDRPOINTER_REG_5__SCAN_IN), .B1(n3273), .Y(n3465));
  XOR2X1  g2417(.A(n3465), .B(n1763), .Y(n3466));
  INVX1   g2418(.A(n3466), .Y(n3467));
  INVX1   g2419(.A(n3410), .Y(n3468));
  NOR4X1  g2420(.A(n3351), .B(n3328), .C(n3325), .D(n3468), .Y(n3469));
  XOR2X1  g2421(.A(n3469), .B(n3467), .Y(n3470));
  NAND4X1 g2422(.A(INSTADDRPOINTER_REG_3__SCAN_IN), .B(INSTADDRPOINTER_REG_2__SCAN_IN), .C(INSTADDRPOINTER_REG_1__SCAN_IN), .D(INSTADDRPOINTER_REG_4__SCAN_IN), .Y(n3471));
  XOR2X1  g2423(.A(n3471), .B(INSTADDRPOINTER_REG_5__SCAN_IN), .Y(n3472));
  OAI22X1 g2424(.A0(n3470), .A1(n3408), .B0(n3354), .B1(n3472), .Y(n3473));
  NOR3X1  g2425(.A(n3473), .B(n3464), .C(n3461), .Y(n3474));
  NAND2X1 g2426(.A(n3474), .B(n3457), .Y(U3013));
  INVX1   g2427(.A(INSTADDRPOINTER_REG_6__SCAN_IN), .Y(n3476));
  NOR3X1  g2428(.A(n3432), .B(n3373), .C(n3334), .Y(n3477));
  AOI22X1 g2429(.A0(n1268), .A1(INSTQUEUE_REG_0__6__SCAN_IN), .B0(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n1244), .Y(n3478));
  AOI22X1 g2430(.A0(n1246), .A1(INSTQUEUE_REG_3__6__SCAN_IN), .B0(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n1337), .Y(n3479));
  AOI22X1 g2431(.A0(n1273), .A1(INSTQUEUE_REG_4__6__SCAN_IN), .B0(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n1329), .Y(n3480));
  AOI22X1 g2432(.A0(n1278), .A1(INSTQUEUE_REG_7__6__SCAN_IN), .B0(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n1270), .Y(n3481));
  NAND4X1 g2433(.A(n3480), .B(n3479), .C(n3478), .D(n3481), .Y(n3482));
  AOI22X1 g2434(.A0(n1253), .A1(INSTQUEUE_REG_12__6__SCAN_IN), .B0(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n1271), .Y(n3483));
  AOI22X1 g2435(.A0(n1279), .A1(INSTQUEUE_REG_15__6__SCAN_IN), .B0(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n1266), .Y(n3484));
  AOI22X1 g2436(.A0(n1323), .A1(INSTQUEUE_REG_8__6__SCAN_IN), .B0(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n1338), .Y(n3485));
  AOI22X1 g2437(.A0(n1255), .A1(INSTQUEUE_REG_11__6__SCAN_IN), .B0(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n1275), .Y(n3486));
  NAND4X1 g2438(.A(n3485), .B(n3484), .C(n3483), .D(n3486), .Y(n3487));
  NOR2X1  g2439(.A(n3487), .B(n3482), .Y(n3488));
  XOR2X1  g2440(.A(n3488), .B(n3477), .Y(n3489));
  NOR2X1  g2441(.A(n3489), .B(n1721), .Y(n3490));
  NOR3X1  g2442(.A(n3488), .B(n1447), .C(n1217), .Y(n3491));
  AOI21X1 g2443(.A0(n1319), .A1(INSTQUEUE_REG_0__6__SCAN_IN), .B0(n3491), .Y(n3492));
  NOR4X1  g2444(.A(n2165), .B(n1403), .C(n1217), .D(n3488), .Y(n3493));
  NOR3X1  g2445(.A(n3488), .B(n2214), .C(n2166), .Y(n3494));
  NOR2X1  g2446(.A(n3494), .B(n3493), .Y(n3495));
  XOR2X1  g2447(.A(n3495), .B(n3492), .Y(n3496));
  NAND2X1 g2448(.A(n3439), .B(n3436), .Y(n3497));
  NAND2X1 g2449(.A(n3448), .B(n3497), .Y(n3498));
  NOR2X1  g2450(.A(n3439), .B(n3436), .Y(n3499));
  INVX1   g2451(.A(n3499), .Y(n3500));
  INVX1   g2452(.A(n3497), .Y(n3501));
  NAND2X1 g2453(.A(n2243), .B(n2265), .Y(n3503));
  OAI21X1 g2454(.A0(n2264), .A1(n2263), .B0(n3441), .Y(n3504));
  AOI21X1 g2455(.A0(n2686), .A1(n2257), .B0(n3504), .Y(n3505));
  INVX1   g2456(.A(n3445), .Y(n3506));
  AOI21X1 g2457(.A0(n3505), .A1(n3503), .B0(n3445), .Y(n3509));
  OAI21X1 g2458(.A0(n3509), .A1(n3501), .B0(n3500), .Y(n3510));
  NOR2X1  g2459(.A(n3496), .B(n3499), .Y(n3511));
  AOI22X1 g2460(.A0(n3510), .A1(n3496), .B0(n3498), .B1(n3511), .Y(n3512));
  AOI21X1 g2461(.A0(n3512), .A1(n1472), .B0(n3490), .Y(n3513));
  XOR2X1  g2462(.A(n3513), .B(n3476), .Y(n3514));
  XOR2X1  g2463(.A(n3509), .B(n3440), .Y(n3515));
  OAI22X1 g2464(.A0(n3433), .A1(n1721), .B0(n1473), .B1(n3515), .Y(n3516));
  NOR2X1  g2465(.A(n3516), .B(INSTADDRPOINTER_REG_5__SCAN_IN), .Y(n3517));
  NAND2X1 g2466(.A(n3516), .B(INSTADDRPOINTER_REG_5__SCAN_IN), .Y(n3518));
  OAI21X1 g2467(.A0(n3455), .A1(n3517), .B0(n3518), .Y(n3519));
  XOR2X1  g2468(.A(n3519), .B(n3514), .Y(n3520));
  NAND2X1 g2469(.A(n3520), .B(n3251), .Y(n3521));
  NOR4X1  g2470(.A(n3420), .B(n3362), .C(n3332), .D(n3345), .Y(n3522));
  XOR2X1  g2471(.A(n3522), .B(n3476), .Y(n3523));
  AOI22X1 g2472(.A0(n3253), .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .B0(REIP_REG_6__SCAN_IN), .B1(n3239), .Y(n3524));
  OAI21X1 g2473(.A0(n3523), .A1(n3344), .B0(n3524), .Y(n3525));
  NAND2X1 g2474(.A(n3462), .B(INSTADDRPOINTER_REG_5__SCAN_IN), .Y(n3526));
  XOR2X1  g2475(.A(n3526), .B(INSTADDRPOINTER_REG_6__SCAN_IN), .Y(n3527));
  NOR2X1  g2476(.A(n3527), .B(n3266), .Y(n3528));
  AOI22X1 g2477(.A0(n3270), .A1(EBX_REG_6__SCAN_IN), .B0(INSTADDRPOINTER_REG_6__SCAN_IN), .B1(n3273), .Y(n3529));
  XOR2X1  g2478(.A(n3529), .B(n1758), .Y(n3530));
  INVX1   g2479(.A(n3530), .Y(n3531));
  NAND4X1 g2480(.A(n3412), .B(n3410), .C(n3411), .D(n3466), .Y(n3532));
  XOR2X1  g2481(.A(n3532), .B(n3531), .Y(n3533));
  NOR2X1  g2482(.A(n3471), .B(n3420), .Y(n3534));
  XOR2X1  g2483(.A(n3534), .B(n3476), .Y(n3535));
  OAI22X1 g2484(.A0(n3533), .A1(n3408), .B0(n3354), .B1(n3535), .Y(n3536));
  NOR3X1  g2485(.A(n3536), .B(n3528), .C(n3525), .Y(n3537));
  NAND2X1 g2486(.A(n3537), .B(n3521), .Y(U3012));
  INVX1   g2487(.A(INSTADDRPOINTER_REG_7__SCAN_IN), .Y(n3539));
  NOR4X1  g2488(.A(n3432), .B(n3373), .C(n3334), .D(n3488), .Y(n3540));
  XOR2X1  g2489(.A(n3540), .B(n2181), .Y(n3541));
  NOR2X1  g2490(.A(n3541), .B(n1721), .Y(n3542));
  NOR2X1  g2491(.A(n3495), .B(n3492), .Y(n3543));
  AOI22X1 g2492(.A0(n1476), .A1(n2165), .B0(n1319), .B1(INSTQUEUE_REG_0__7__SCAN_IN), .Y(n3544));
  XOR2X1  g2493(.A(n2166), .B(n3544), .Y(n3546));
  NOR3X1  g2494(.A(n3546), .B(n3543), .C(n3499), .Y(n3547));
  INVX1   g2495(.A(n3547), .Y(n3548));
  AOI21X1 g2496(.A0(n3448), .A1(n3497), .B0(n3548), .Y(n3549));
  NAND2X1 g2497(.A(n3505), .B(n3503), .Y(n3550));
  OAI22X1 g2498(.A0(n3436), .A1(n3439), .B0(n3380), .B1(n3377), .Y(n3551));
  AOI21X1 g2499(.A0(n3446), .A1(n2261), .B0(n3551), .Y(n3552));
  NAND2X1 g2500(.A(n3495), .B(n3492), .Y(n3553));
  INVX1   g2501(.A(n3553), .Y(n3554));
  INVX1   g2502(.A(n3544), .Y(n3555));
  AOI21X1 g2503(.A0(n2165), .A1(n2121), .B0(n3555), .Y(n3556));
  NOR2X1  g2504(.A(n2166), .B(n3544), .Y(n3557));
  NOR4X1  g2505(.A(n3556), .B(n3554), .C(n3501), .D(n3557), .Y(n3558));
  INVX1   g2506(.A(n3558), .Y(n3559));
  AOI21X1 g2507(.A0(n3552), .A1(n3550), .B0(n3559), .Y(n3560));
  NOR2X1  g2508(.A(n3546), .B(n3553), .Y(n3561));
  AOI21X1 g2509(.A0(n3546), .A1(n3543), .B0(n3561), .Y(n3562));
  NOR4X1  g2510(.A(n3560), .B(n3549), .C(n1473), .D(n3561), .Y(n3564));
  NOR2X1  g2511(.A(n3564), .B(n3542), .Y(n3565));
  XOR2X1  g2512(.A(n3565), .B(n3539), .Y(n3566));
  NOR2X1  g2513(.A(n3513), .B(n3476), .Y(n3567));
  NAND2X1 g2514(.A(n3513), .B(n3476), .Y(n3568));
  AOI21X1 g2515(.A0(n3519), .A1(n3568), .B0(n3567), .Y(n3569));
  XOR2X1  g2516(.A(n3569), .B(n3566), .Y(n3570));
  NAND2X1 g2517(.A(n3522), .B(INSTADDRPOINTER_REG_6__SCAN_IN), .Y(n3571));
  XOR2X1  g2518(.A(n3571), .B(INSTADDRPOINTER_REG_7__SCAN_IN), .Y(n3572));
  AOI22X1 g2519(.A0(n3253), .A1(INSTADDRPOINTER_REG_7__SCAN_IN), .B0(REIP_REG_7__SCAN_IN), .B1(n3239), .Y(n3573));
  OAI21X1 g2520(.A0(n3572), .A1(n3344), .B0(n3573), .Y(n3574));
  INVX1   g2521(.A(n3462), .Y(n3575));
  NOR3X1  g2522(.A(n3575), .B(n3476), .C(n3420), .Y(n3576));
  XOR2X1  g2523(.A(n3576), .B(n3539), .Y(n3577));
  NOR2X1  g2524(.A(n3577), .B(n3266), .Y(n3578));
  AOI22X1 g2525(.A0(n3270), .A1(EBX_REG_7__SCAN_IN), .B0(INSTADDRPOINTER_REG_7__SCAN_IN), .B1(n3273), .Y(n3579));
  XOR2X1  g2526(.A(n3579), .B(n1758), .Y(n3580));
  NOR2X1  g2527(.A(n3532), .B(n3530), .Y(n3581));
  XOR2X1  g2528(.A(n3581), .B(n3580), .Y(n3582));
  NOR3X1  g2529(.A(n3471), .B(n3476), .C(n3420), .Y(n3583));
  XOR2X1  g2530(.A(n3583), .B(n3539), .Y(n3584));
  OAI22X1 g2531(.A0(n3582), .A1(n3408), .B0(n3354), .B1(n3584), .Y(n3585));
  NOR3X1  g2532(.A(n3585), .B(n3578), .C(n3574), .Y(n3586));
  OAI21X1 g2533(.A0(n3570), .A1(n3250), .B0(n3586), .Y(U3011));
  INVX1   g2534(.A(INSTADDRPOINTER_REG_8__SCAN_IN), .Y(n3588));
  NOR3X1  g2535(.A(n3488), .B(n2181), .C(n1721), .Y(n3589));
  AOI22X1 g2536(.A0(n1279), .A1(INSTQUEUE_REG_0__0__SCAN_IN), .B0(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n1268), .Y(n3592));
  AOI22X1 g2537(.A0(n1337), .A1(INSTQUEUE_REG_3__0__SCAN_IN), .B0(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n1244), .Y(n3595));
  AOI22X1 g2538(.A0(n1246), .A1(INSTQUEUE_REG_4__0__SCAN_IN), .B0(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n1273), .Y(n3598));
  AOI22X1 g2539(.A0(n1270), .A1(INSTQUEUE_REG_7__0__SCAN_IN), .B0(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n1329), .Y(n3601));
  NAND4X1 g2540(.A(n3598), .B(n3595), .C(n3592), .D(n3601), .Y(n3602));
  AOI22X1 g2541(.A0(n1255), .A1(INSTQUEUE_REG_12__0__SCAN_IN), .B0(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n1253), .Y(n3605));
  AOI22X1 g2542(.A0(n1266), .A1(INSTQUEUE_REG_15__0__SCAN_IN), .B0(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n1271), .Y(n3608));
  AOI22X1 g2543(.A0(n1278), .A1(INSTQUEUE_REG_8__0__SCAN_IN), .B0(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n1323), .Y(n3611));
  AOI22X1 g2544(.A0(n1275), .A1(INSTQUEUE_REG_11__0__SCAN_IN), .B0(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n1338), .Y(n3614));
  NAND4X1 g2545(.A(n3611), .B(n3608), .C(n3605), .D(n3614), .Y(n3615));
  AOI21X1 g2546(.A0(n1318), .A1(n1447), .B0(n1217), .Y(n3616));
  OAI21X1 g2547(.A0(n3615), .A1(n3602), .B0(n3616), .Y(n3617));
  XOR2X1  g2548(.A(n3617), .B(n2167), .Y(n3618));
  AOI21X1 g2549(.A0(n3495), .A1(n3492), .B0(n3556), .Y(n3619));
  INVX1   g2550(.A(n3619), .Y(n3620));
  NOR3X1  g2551(.A(n3620), .B(n3501), .C(n3442), .Y(n3621));
  NOR2X1  g2552(.A(n3620), .B(n3500), .Y(n3622));
  NOR3X1  g2553(.A(n3556), .B(n3495), .C(n3492), .Y(n3623));
  NOR3X1  g2554(.A(n3620), .B(n3501), .C(n3506), .Y(n3624));
  NOR4X1  g2555(.A(n3623), .B(n3622), .C(n3557), .D(n3624), .Y(n3625));
  AOI21X1 g2556(.A0(n3621), .A1(n3386), .B0(n3557), .Y(n3627));
  XOR2X1  g2557(.A(n3627), .B(n3618), .Y(n3628));
  AOI22X1 g2558(.A0(n3589), .A1(n3477), .B0(n1472), .B1(n3628), .Y(n3629));
  XOR2X1  g2559(.A(n3629), .B(n3588), .Y(n3630));
  NAND2X1 g2560(.A(n3337), .B(n3332), .Y(n3631));
  NOR2X1  g2561(.A(n3337), .B(n3332), .Y(n3632));
  AOI21X1 g2562(.A0(n3341), .A1(n3631), .B0(n3632), .Y(n3633));
  INVX1   g2563(.A(n3496), .Y(n3634));
  AOI21X1 g2564(.A0(n3448), .A1(n3497), .B0(n3499), .Y(n3635));
  OAI21X1 g2565(.A0(n3509), .A1(n3501), .B0(n3511), .Y(n3636));
  OAI21X1 g2566(.A0(n3635), .A1(n3634), .B0(n3636), .Y(n3637));
  OAI22X1 g2567(.A0(n3489), .A1(n1721), .B0(n1473), .B1(n3637), .Y(n3638));
  NOR2X1  g2568(.A(n3638), .B(INSTADDRPOINTER_REG_6__SCAN_IN), .Y(n3639));
  INVX1   g2569(.A(n3542), .Y(n3640));
  OAI21X1 g2570(.A0(n3509), .A1(n3501), .B0(n3547), .Y(n3641));
  OAI21X1 g2571(.A0(n3444), .A1(n3383), .B0(n3552), .Y(n3642));
  NAND2X1 g2572(.A(n3558), .B(n3642), .Y(n3643));
  NAND4X1 g2573(.A(n3643), .B(n3641), .C(n1472), .D(n3562), .Y(n3644));
  NAND3X1 g2574(.A(n3644), .B(n3640), .C(n3539), .Y(n3645));
  AOI22X1 g2575(.A0(n3388), .A1(n3362), .B0(n3420), .B1(n3450), .Y(n3646));
  NAND2X1 g2576(.A(n3646), .B(n3645), .Y(n3647));
  NOR3X1  g2577(.A(n3647), .B(n3639), .C(n3633), .Y(n3648));
  NAND2X1 g2578(.A(n3450), .B(n3420), .Y(n3649));
  NAND3X1 g2579(.A(n3645), .B(n3649), .C(n3454), .Y(n3650));
  OAI22X1 g2580(.A0(n3565), .A1(n3539), .B0(n3639), .B1(n3650), .Y(n3651));
  NAND3X1 g2581(.A(n3645), .B(n3516), .C(INSTADDRPOINTER_REG_5__SCAN_IN), .Y(n3652));
  NAND3X1 g2582(.A(n3645), .B(n3638), .C(INSTADDRPOINTER_REG_6__SCAN_IN), .Y(n3653));
  OAI21X1 g2583(.A0(n3652), .A1(n3639), .B0(n3653), .Y(n3654));
  NOR3X1  g2584(.A(n3654), .B(n3651), .C(n3648), .Y(n3655));
  XOR2X1  g2585(.A(n3655), .B(n3630), .Y(n3656));
  NAND3X1 g2586(.A(n3522), .B(INSTADDRPOINTER_REG_7__SCAN_IN), .C(INSTADDRPOINTER_REG_6__SCAN_IN), .Y(n3657));
  XOR2X1  g2587(.A(n3657), .B(INSTADDRPOINTER_REG_8__SCAN_IN), .Y(n3658));
  AOI22X1 g2588(.A0(n3253), .A1(INSTADDRPOINTER_REG_8__SCAN_IN), .B0(REIP_REG_8__SCAN_IN), .B1(n3239), .Y(n3659));
  OAI21X1 g2589(.A0(n3658), .A1(n3344), .B0(n3659), .Y(n3660));
  NAND4X1 g2590(.A(INSTADDRPOINTER_REG_7__SCAN_IN), .B(INSTADDRPOINTER_REG_6__SCAN_IN), .C(INSTADDRPOINTER_REG_5__SCAN_IN), .D(n3462), .Y(n3661));
  XOR2X1  g2591(.A(n3661), .B(INSTADDRPOINTER_REG_8__SCAN_IN), .Y(n3662));
  NOR2X1  g2592(.A(n3662), .B(n3266), .Y(n3663));
  AOI22X1 g2593(.A0(n3270), .A1(EBX_REG_8__SCAN_IN), .B0(INSTADDRPOINTER_REG_8__SCAN_IN), .B1(n3273), .Y(n3664));
  XOR2X1  g2594(.A(n3664), .B(n1758), .Y(n3665));
  NOR3X1  g2595(.A(n3580), .B(n3532), .C(n3530), .Y(n3666));
  XOR2X1  g2596(.A(n3666), .B(n3665), .Y(n3667));
  NOR4X1  g2597(.A(n3539), .B(n3476), .C(n3420), .D(n3471), .Y(n3668));
  XOR2X1  g2598(.A(n3668), .B(n3588), .Y(n3669));
  OAI22X1 g2599(.A0(n3667), .A1(n3408), .B0(n3354), .B1(n3669), .Y(n3670));
  NOR3X1  g2600(.A(n3670), .B(n3663), .C(n3660), .Y(n3671));
  OAI21X1 g2601(.A0(n3656), .A1(n3250), .B0(n3671), .Y(U3010));
  NOR2X1  g2602(.A(n3627), .B(n3618), .Y(n3673));
  AOI22X1 g2603(.A0(n1279), .A1(INSTQUEUE_REG_0__1__SCAN_IN), .B0(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n1268), .Y(n3674));
  AOI22X1 g2604(.A0(n1337), .A1(INSTQUEUE_REG_3__1__SCAN_IN), .B0(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n1244), .Y(n3675));
  AOI22X1 g2605(.A0(n1246), .A1(INSTQUEUE_REG_4__1__SCAN_IN), .B0(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n1273), .Y(n3676));
  AOI22X1 g2606(.A0(n1270), .A1(INSTQUEUE_REG_7__1__SCAN_IN), .B0(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n1329), .Y(n3677));
  NAND4X1 g2607(.A(n3676), .B(n3675), .C(n3674), .D(n3677), .Y(n3678));
  AOI22X1 g2608(.A0(n1255), .A1(INSTQUEUE_REG_12__1__SCAN_IN), .B0(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n1253), .Y(n3679));
  AOI22X1 g2609(.A0(n1266), .A1(INSTQUEUE_REG_15__1__SCAN_IN), .B0(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n1271), .Y(n3680));
  AOI22X1 g2610(.A0(n1278), .A1(INSTQUEUE_REG_8__1__SCAN_IN), .B0(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n1323), .Y(n3681));
  AOI22X1 g2611(.A0(n1275), .A1(INSTQUEUE_REG_11__1__SCAN_IN), .B0(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n1338), .Y(n3682));
  NAND4X1 g2612(.A(n3681), .B(n3680), .C(n3679), .D(n3682), .Y(n3683));
  OAI21X1 g2613(.A0(n3683), .A1(n3678), .B0(n3616), .Y(n3684));
  XOR2X1  g2614(.A(n3684), .B(n2167), .Y(n3685));
  INVX1   g2615(.A(n3685), .Y(n3686));
  XOR2X1  g2616(.A(n3686), .B(n3673), .Y(n3687));
  AOI21X1 g2617(.A0(n3687), .A1(n1472), .B0(INSTADDRPOINTER_REG_9__SCAN_IN), .Y(n3688));
  INVX1   g2618(.A(INSTADDRPOINTER_REG_9__SCAN_IN), .Y(n3689));
  XOR2X1  g2619(.A(n3685), .B(n3673), .Y(n3690));
  NOR3X1  g2620(.A(n3690), .B(n1473), .C(n3689), .Y(n3691));
  NOR2X1  g2621(.A(n3691), .B(n3688), .Y(n3692));
  NAND2X1 g2622(.A(n3629), .B(n3588), .Y(n3693));
  NOR2X1  g2623(.A(n3629), .B(n3588), .Y(n3694));
  NAND4X1 g2624(.A(n3645), .B(n3568), .C(n3398), .D(n3646), .Y(n3695));
  AOI21X1 g2625(.A0(n3644), .A1(n3640), .B0(n3539), .Y(n3696));
  NOR3X1  g2626(.A(n3564), .B(n3542), .C(INSTADDRPOINTER_REG_7__SCAN_IN), .Y(n3697));
  NOR4X1  g2627(.A(n3517), .B(n3388), .C(n3362), .D(n3697), .Y(n3698));
  AOI21X1 g2628(.A0(n3698), .A1(n3568), .B0(n3696), .Y(n3699));
  NOR2X1  g2629(.A(n3697), .B(n3518), .Y(n3700));
  AOI22X1 g2630(.A0(n3645), .A1(n3567), .B0(n3568), .B1(n3700), .Y(n3701));
  NAND3X1 g2631(.A(n3701), .B(n3699), .C(n3695), .Y(n3702));
  AOI21X1 g2632(.A0(n3702), .A1(n3693), .B0(n3694), .Y(n3703));
  XOR2X1  g2633(.A(n3703), .B(n3692), .Y(n3704));
  NAND4X1 g2634(.A(INSTADDRPOINTER_REG_8__SCAN_IN), .B(INSTADDRPOINTER_REG_7__SCAN_IN), .C(INSTADDRPOINTER_REG_6__SCAN_IN), .D(n3522), .Y(n3705));
  XOR2X1  g2635(.A(n3705), .B(INSTADDRPOINTER_REG_9__SCAN_IN), .Y(n3706));
  AOI22X1 g2636(.A0(n3253), .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .B0(REIP_REG_9__SCAN_IN), .B1(n3239), .Y(n3707));
  OAI21X1 g2637(.A0(n3706), .A1(n3344), .B0(n3707), .Y(n3708));
  NAND3X1 g2638(.A(n3576), .B(INSTADDRPOINTER_REG_8__SCAN_IN), .C(INSTADDRPOINTER_REG_7__SCAN_IN), .Y(n3709));
  XOR2X1  g2639(.A(n3709), .B(INSTADDRPOINTER_REG_9__SCAN_IN), .Y(n3710));
  NOR2X1  g2640(.A(n3710), .B(n3266), .Y(n3711));
  AOI22X1 g2641(.A0(n3270), .A1(EBX_REG_9__SCAN_IN), .B0(INSTADDRPOINTER_REG_9__SCAN_IN), .B1(n3273), .Y(n3712));
  XOR2X1  g2642(.A(n3712), .B(n1758), .Y(n3713));
  NOR4X1  g2643(.A(n3580), .B(n3532), .C(n3530), .D(n3665), .Y(n3714));
  XOR2X1  g2644(.A(n3714), .B(n3713), .Y(n3715));
  NAND2X1 g2645(.A(n3668), .B(INSTADDRPOINTER_REG_8__SCAN_IN), .Y(n3716));
  XOR2X1  g2646(.A(n3716), .B(INSTADDRPOINTER_REG_9__SCAN_IN), .Y(n3717));
  OAI22X1 g2647(.A0(n3715), .A1(n3408), .B0(n3354), .B1(n3717), .Y(n3718));
  NOR3X1  g2648(.A(n3718), .B(n3711), .C(n3708), .Y(n3719));
  OAI21X1 g2649(.A0(n3704), .A1(n3250), .B0(n3719), .Y(U3009));
  INVX1   g2650(.A(INSTADDRPOINTER_REG_10__SCAN_IN), .Y(n3721));
  AOI22X1 g2651(.A0(n1279), .A1(INSTQUEUE_REG_0__2__SCAN_IN), .B0(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n1268), .Y(n3722));
  AOI22X1 g2652(.A0(n1337), .A1(INSTQUEUE_REG_3__2__SCAN_IN), .B0(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n1244), .Y(n3723));
  AOI22X1 g2653(.A0(n1246), .A1(INSTQUEUE_REG_4__2__SCAN_IN), .B0(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n1273), .Y(n3724));
  AOI22X1 g2654(.A0(n1270), .A1(INSTQUEUE_REG_7__2__SCAN_IN), .B0(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n1329), .Y(n3725));
  NAND4X1 g2655(.A(n3724), .B(n3723), .C(n3722), .D(n3725), .Y(n3726));
  AOI22X1 g2656(.A0(n1255), .A1(INSTQUEUE_REG_12__2__SCAN_IN), .B0(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n1253), .Y(n3727));
  AOI22X1 g2657(.A0(n1266), .A1(INSTQUEUE_REG_15__2__SCAN_IN), .B0(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n1271), .Y(n3728));
  AOI22X1 g2658(.A0(n1278), .A1(INSTQUEUE_REG_8__2__SCAN_IN), .B0(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n1323), .Y(n3729));
  AOI22X1 g2659(.A0(n1275), .A1(INSTQUEUE_REG_11__2__SCAN_IN), .B0(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n1338), .Y(n3730));
  NAND4X1 g2660(.A(n3729), .B(n3728), .C(n3727), .D(n3730), .Y(n3731));
  OAI21X1 g2661(.A0(n3731), .A1(n3726), .B0(n3616), .Y(n3732));
  XOR2X1  g2662(.A(n3732), .B(n2167), .Y(n3733));
  INVX1   g2663(.A(n3733), .Y(n3734));
  NOR2X1  g2664(.A(n3685), .B(n3618), .Y(n3735));
  INVX1   g2665(.A(n3735), .Y(n3736));
  NOR2X1  g2666(.A(n3736), .B(n3627), .Y(n3737));
  XOR2X1  g2667(.A(n3737), .B(n3734), .Y(n3738));
  NAND2X1 g2668(.A(n3738), .B(n1472), .Y(n3739));
  XOR2X1  g2669(.A(n3739), .B(n3721), .Y(n3740));
  NOR2X1  g2670(.A(n3703), .B(n3688), .Y(n3741));
  NOR2X1  g2671(.A(n3741), .B(n3691), .Y(n3742));
  XOR2X1  g2672(.A(n3742), .B(n3740), .Y(n3743));
  NOR2X1  g2673(.A(n3705), .B(n3689), .Y(n3744));
  XOR2X1  g2674(.A(n3744), .B(n3721), .Y(n3745));
  AOI22X1 g2675(.A0(n3253), .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .B0(REIP_REG_10__SCAN_IN), .B1(n3239), .Y(n3746));
  OAI21X1 g2676(.A0(n3745), .A1(n3344), .B0(n3746), .Y(n3747));
  NAND4X1 g2677(.A(INSTADDRPOINTER_REG_9__SCAN_IN), .B(INSTADDRPOINTER_REG_8__SCAN_IN), .C(INSTADDRPOINTER_REG_7__SCAN_IN), .D(n3576), .Y(n3748));
  XOR2X1  g2678(.A(n3748), .B(INSTADDRPOINTER_REG_10__SCAN_IN), .Y(n3749));
  NOR2X1  g2679(.A(n3749), .B(n3266), .Y(n3750));
  AOI22X1 g2680(.A0(n3270), .A1(EBX_REG_10__SCAN_IN), .B0(INSTADDRPOINTER_REG_10__SCAN_IN), .B1(n3273), .Y(n3751));
  XOR2X1  g2681(.A(n3751), .B(n1758), .Y(n3752));
  INVX1   g2682(.A(n3752), .Y(n3753));
  NOR2X1  g2683(.A(n3713), .B(n3665), .Y(n3754));
  NAND2X1 g2684(.A(n3754), .B(n3666), .Y(n3755));
  XOR2X1  g2685(.A(n3755), .B(n3753), .Y(n3756));
  NAND3X1 g2686(.A(n3668), .B(INSTADDRPOINTER_REG_9__SCAN_IN), .C(INSTADDRPOINTER_REG_8__SCAN_IN), .Y(n3757));
  XOR2X1  g2687(.A(n3757), .B(INSTADDRPOINTER_REG_10__SCAN_IN), .Y(n3758));
  OAI22X1 g2688(.A0(n3756), .A1(n3408), .B0(n3354), .B1(n3758), .Y(n3759));
  NOR3X1  g2689(.A(n3759), .B(n3750), .C(n3747), .Y(n3760));
  OAI21X1 g2690(.A0(n3743), .A1(n3250), .B0(n3760), .Y(U3008));
  INVX1   g2691(.A(INSTADDRPOINTER_REG_11__SCAN_IN), .Y(n3762));
  AOI22X1 g2692(.A0(n1279), .A1(INSTQUEUE_REG_0__3__SCAN_IN), .B0(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n1268), .Y(n3763));
  AOI22X1 g2693(.A0(n1337), .A1(INSTQUEUE_REG_3__3__SCAN_IN), .B0(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n1244), .Y(n3764));
  AOI22X1 g2694(.A0(n1246), .A1(INSTQUEUE_REG_4__3__SCAN_IN), .B0(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n1273), .Y(n3765));
  AOI22X1 g2695(.A0(n1270), .A1(INSTQUEUE_REG_7__3__SCAN_IN), .B0(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n1329), .Y(n3766));
  NAND4X1 g2696(.A(n3765), .B(n3764), .C(n3763), .D(n3766), .Y(n3767));
  AOI22X1 g2697(.A0(n1255), .A1(INSTQUEUE_REG_12__3__SCAN_IN), .B0(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n1253), .Y(n3768));
  AOI22X1 g2698(.A0(n1266), .A1(INSTQUEUE_REG_15__3__SCAN_IN), .B0(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n1271), .Y(n3769));
  AOI22X1 g2699(.A0(n1278), .A1(INSTQUEUE_REG_8__3__SCAN_IN), .B0(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n1323), .Y(n3770));
  AOI22X1 g2700(.A0(n1275), .A1(INSTQUEUE_REG_11__3__SCAN_IN), .B0(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n1338), .Y(n3771));
  NAND4X1 g2701(.A(n3770), .B(n3769), .C(n3768), .D(n3771), .Y(n3772));
  OAI21X1 g2702(.A0(n3772), .A1(n3767), .B0(n3616), .Y(n3773));
  XOR2X1  g2703(.A(n3773), .B(n2167), .Y(n3774));
  NOR3X1  g2704(.A(n3736), .B(n3733), .C(n3627), .Y(n3775));
  XOR2X1  g2705(.A(n3775), .B(n3774), .Y(n3776));
  OAI21X1 g2706(.A0(n3776), .A1(n1473), .B0(n3762), .Y(n3777));
  INVX1   g2707(.A(n3774), .Y(n3778));
  XOR2X1  g2708(.A(n3775), .B(n3778), .Y(n3779));
  NAND3X1 g2709(.A(n3779), .B(n1472), .C(INSTADDRPOINTER_REG_11__SCAN_IN), .Y(n3780));
  NAND2X1 g2710(.A(n3780), .B(n3777), .Y(n3781));
  NAND3X1 g2711(.A(n3738), .B(n1472), .C(INSTADDRPOINTER_REG_10__SCAN_IN), .Y(n3782));
  AOI21X1 g2712(.A0(n3738), .A1(n1472), .B0(INSTADDRPOINTER_REG_10__SCAN_IN), .Y(n3783));
  OAI21X1 g2713(.A0(n3742), .A1(n3783), .B0(n3782), .Y(n3784));
  XOR2X1  g2714(.A(n3784), .B(n3781), .Y(n3785));
  NOR3X1  g2715(.A(n3705), .B(n3721), .C(n3689), .Y(n3786));
  XOR2X1  g2716(.A(n3786), .B(n3762), .Y(n3787));
  AOI22X1 g2717(.A0(n3253), .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .B0(REIP_REG_11__SCAN_IN), .B1(n3239), .Y(n3788));
  OAI21X1 g2718(.A0(n3787), .A1(n3344), .B0(n3788), .Y(n3789));
  NOR3X1  g2719(.A(n3709), .B(n3721), .C(n3689), .Y(n3790));
  XOR2X1  g2720(.A(n3790), .B(n3762), .Y(n3791));
  NOR2X1  g2721(.A(n3791), .B(n3266), .Y(n3792));
  AOI22X1 g2722(.A0(n3270), .A1(EBX_REG_11__SCAN_IN), .B0(INSTADDRPOINTER_REG_11__SCAN_IN), .B1(n3273), .Y(n3793));
  XOR2X1  g2723(.A(n3793), .B(n1758), .Y(n3794));
  NOR2X1  g2724(.A(n3755), .B(n3752), .Y(n3795));
  XOR2X1  g2725(.A(n3795), .B(n3794), .Y(n3796));
  NAND4X1 g2726(.A(INSTADDRPOINTER_REG_10__SCAN_IN), .B(INSTADDRPOINTER_REG_9__SCAN_IN), .C(INSTADDRPOINTER_REG_8__SCAN_IN), .D(n3668), .Y(n3797));
  XOR2X1  g2727(.A(n3797), .B(INSTADDRPOINTER_REG_11__SCAN_IN), .Y(n3798));
  OAI22X1 g2728(.A0(n3796), .A1(n3408), .B0(n3354), .B1(n3798), .Y(n3799));
  NOR3X1  g2729(.A(n3799), .B(n3792), .C(n3789), .Y(n3800));
  OAI21X1 g2730(.A0(n3785), .A1(n3250), .B0(n3800), .Y(U3007));
  AOI22X1 g2731(.A0(n1279), .A1(INSTQUEUE_REG_0__4__SCAN_IN), .B0(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n1268), .Y(n3802));
  AOI22X1 g2732(.A0(n1337), .A1(INSTQUEUE_REG_3__4__SCAN_IN), .B0(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n1244), .Y(n3803));
  AOI22X1 g2733(.A0(n1246), .A1(INSTQUEUE_REG_4__4__SCAN_IN), .B0(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n1273), .Y(n3804));
  AOI22X1 g2734(.A0(n1270), .A1(INSTQUEUE_REG_7__4__SCAN_IN), .B0(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n1329), .Y(n3805));
  NAND4X1 g2735(.A(n3804), .B(n3803), .C(n3802), .D(n3805), .Y(n3806));
  AOI22X1 g2736(.A0(n1255), .A1(INSTQUEUE_REG_12__4__SCAN_IN), .B0(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n1253), .Y(n3807));
  AOI22X1 g2737(.A0(n1266), .A1(INSTQUEUE_REG_15__4__SCAN_IN), .B0(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n1271), .Y(n3808));
  AOI22X1 g2738(.A0(n1278), .A1(INSTQUEUE_REG_8__4__SCAN_IN), .B0(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n1323), .Y(n3809));
  AOI22X1 g2739(.A0(n1275), .A1(INSTQUEUE_REG_11__4__SCAN_IN), .B0(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n1338), .Y(n3810));
  NAND4X1 g2740(.A(n3809), .B(n3808), .C(n3807), .D(n3810), .Y(n3811));
  OAI21X1 g2741(.A0(n3811), .A1(n3806), .B0(n3616), .Y(n3812));
  XOR2X1  g2742(.A(n3812), .B(n2167), .Y(n3813));
  INVX1   g2743(.A(n3813), .Y(n3814));
  NOR4X1  g2744(.A(n3733), .B(n3685), .C(n3618), .D(n3774), .Y(n3815));
  INVX1   g2745(.A(n3815), .Y(n3816));
  NOR2X1  g2746(.A(n3816), .B(n3627), .Y(n3817));
  XOR2X1  g2747(.A(n3817), .B(n3814), .Y(n3818));
  AOI21X1 g2748(.A0(n3818), .A1(n1472), .B0(INSTADDRPOINTER_REG_12__SCAN_IN), .Y(n3819));
  INVX1   g2749(.A(n3819), .Y(n3820));
  NAND3X1 g2750(.A(n3818), .B(n1472), .C(INSTADDRPOINTER_REG_12__SCAN_IN), .Y(n3821));
  NAND2X1 g2751(.A(n3821), .B(n3820), .Y(n3822));
  OAI21X1 g2752(.A0(n3690), .A1(n1473), .B0(n3689), .Y(n3823));
  XOR2X1  g2753(.A(n3737), .B(n3733), .Y(n3824));
  OAI21X1 g2754(.A0(n3824), .A1(n1473), .B0(n3721), .Y(n3825));
  NAND4X1 g2755(.A(n3825), .B(n3823), .C(n3693), .D(n3777), .Y(n3826));
  NOR3X1  g2756(.A(n3776), .B(n1473), .C(n3762), .Y(n3827));
  NAND3X1 g2757(.A(n3687), .B(n1472), .C(INSTADDRPOINTER_REG_9__SCAN_IN), .Y(n3828));
  AOI21X1 g2758(.A0(n3779), .A1(n1472), .B0(INSTADDRPOINTER_REG_11__SCAN_IN), .Y(n3829));
  NOR3X1  g2759(.A(n3829), .B(n3783), .C(n3828), .Y(n3830));
  NOR3X1  g2760(.A(n3829), .B(n3739), .C(n3721), .Y(n3831));
  NAND2X1 g2761(.A(n3589), .B(n3477), .Y(n3832));
  AOI21X1 g2762(.A0(n2686), .A1(n2257), .B0(n2266), .Y(n3833));
  AOI22X1 g2763(.A0(n3503), .A1(n3833), .B0(n2261), .B1(n3384), .Y(n3834));
  INVX1   g2764(.A(n3621), .Y(n3835));
  OAI21X1 g2765(.A0(n3835), .A1(n3834), .B0(n3625), .Y(n3836));
  XOR2X1  g2766(.A(n3836), .B(n3618), .Y(n3837));
  OAI21X1 g2767(.A0(n3837), .A1(n1473), .B0(n3832), .Y(n3838));
  NAND2X1 g2768(.A(n3838), .B(INSTADDRPOINTER_REG_8__SCAN_IN), .Y(n3839));
  NOR4X1  g2769(.A(n3783), .B(n3688), .C(n3839), .D(n3829), .Y(n3840));
  NOR4X1  g2770(.A(n3831), .B(n3830), .C(n3827), .D(n3840), .Y(n3841));
  OAI21X1 g2771(.A0(n3826), .A1(n3655), .B0(n3841), .Y(n3842));
  XOR2X1  g2772(.A(n3842), .B(n3822), .Y(n3843));
  INVX1   g2773(.A(INSTADDRPOINTER_REG_12__SCAN_IN), .Y(n3844));
  NOR4X1  g2774(.A(n3762), .B(n3721), .C(n3689), .D(n3705), .Y(n3845));
  XOR2X1  g2775(.A(n3845), .B(n3844), .Y(n3846));
  AOI22X1 g2776(.A0(n3253), .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .B0(REIP_REG_12__SCAN_IN), .B1(n3239), .Y(n3847));
  OAI21X1 g2777(.A0(n3846), .A1(n3344), .B0(n3847), .Y(n3848));
  NOR4X1  g2778(.A(n3762), .B(n3721), .C(n3689), .D(n3709), .Y(n3849));
  XOR2X1  g2779(.A(n3849), .B(n3844), .Y(n3850));
  NOR2X1  g2780(.A(n3850), .B(n3266), .Y(n3851));
  AOI22X1 g2781(.A0(n3270), .A1(EBX_REG_12__SCAN_IN), .B0(INSTADDRPOINTER_REG_12__SCAN_IN), .B1(n3273), .Y(n3852));
  XOR2X1  g2782(.A(n3852), .B(n1758), .Y(n3853));
  NOR3X1  g2783(.A(n3794), .B(n3755), .C(n3752), .Y(n3854));
  XOR2X1  g2784(.A(n3854), .B(n3853), .Y(n3855));
  NOR2X1  g2785(.A(n3797), .B(n3762), .Y(n3856));
  XOR2X1  g2786(.A(n3856), .B(n3844), .Y(n3857));
  OAI22X1 g2787(.A0(n3855), .A1(n3408), .B0(n3354), .B1(n3857), .Y(n3858));
  NOR3X1  g2788(.A(n3858), .B(n3851), .C(n3848), .Y(n3859));
  OAI21X1 g2789(.A0(n3843), .A1(n3250), .B0(n3859), .Y(U3006));
  INVX1   g2790(.A(INSTADDRPOINTER_REG_13__SCAN_IN), .Y(n3861));
  AOI22X1 g2791(.A0(n1279), .A1(INSTQUEUE_REG_0__5__SCAN_IN), .B0(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n1268), .Y(n3862));
  AOI22X1 g2792(.A0(n1337), .A1(INSTQUEUE_REG_3__5__SCAN_IN), .B0(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n1244), .Y(n3863));
  AOI22X1 g2793(.A0(n1246), .A1(INSTQUEUE_REG_4__5__SCAN_IN), .B0(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n1273), .Y(n3864));
  AOI22X1 g2794(.A0(n1270), .A1(INSTQUEUE_REG_7__5__SCAN_IN), .B0(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n1329), .Y(n3865));
  NAND4X1 g2795(.A(n3864), .B(n3863), .C(n3862), .D(n3865), .Y(n3866));
  AOI22X1 g2796(.A0(n1255), .A1(INSTQUEUE_REG_12__5__SCAN_IN), .B0(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n1253), .Y(n3867));
  AOI22X1 g2797(.A0(n1266), .A1(INSTQUEUE_REG_15__5__SCAN_IN), .B0(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n1271), .Y(n3868));
  AOI22X1 g2798(.A0(n1278), .A1(INSTQUEUE_REG_8__5__SCAN_IN), .B0(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n1323), .Y(n3869));
  AOI22X1 g2799(.A0(n1275), .A1(INSTQUEUE_REG_11__5__SCAN_IN), .B0(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n1338), .Y(n3870));
  NAND4X1 g2800(.A(n3869), .B(n3868), .C(n3867), .D(n3870), .Y(n3871));
  OAI21X1 g2801(.A0(n3871), .A1(n3866), .B0(n3616), .Y(n3872));
  XOR2X1  g2802(.A(n3872), .B(n2167), .Y(n3873));
  NOR3X1  g2803(.A(n3816), .B(n3813), .C(n3627), .Y(n3874));
  XOR2X1  g2804(.A(n3874), .B(n3873), .Y(n3875));
  OAI21X1 g2805(.A0(n3875), .A1(n1473), .B0(n3861), .Y(n3876));
  INVX1   g2806(.A(n3873), .Y(n3877));
  XOR2X1  g2807(.A(n3874), .B(n3877), .Y(n3878));
  NAND3X1 g2808(.A(n3878), .B(n1472), .C(INSTADDRPOINTER_REG_13__SCAN_IN), .Y(n3879));
  NAND2X1 g2809(.A(n3879), .B(n3876), .Y(n3880));
  NOR2X1  g2810(.A(n3838), .B(INSTADDRPOINTER_REG_8__SCAN_IN), .Y(n3881));
  NOR4X1  g2811(.A(n3783), .B(n3688), .C(n3881), .D(n3829), .Y(n3882));
  NAND3X1 g2812(.A(n3777), .B(n3825), .C(n3691), .Y(n3883));
  NAND4X1 g2813(.A(n3738), .B(n1472), .C(INSTADDRPOINTER_REG_10__SCAN_IN), .D(n3777), .Y(n3884));
  NAND4X1 g2814(.A(n3825), .B(n3823), .C(n3694), .D(n3777), .Y(n3885));
  NAND4X1 g2815(.A(n3884), .B(n3883), .C(n3780), .D(n3885), .Y(n3886));
  AOI21X1 g2816(.A0(n3882), .A1(n3702), .B0(n3886), .Y(n3887));
  OAI21X1 g2817(.A0(n3887), .A1(n3819), .B0(n3821), .Y(n3888));
  XOR2X1  g2818(.A(n3888), .B(n3880), .Y(n3889));
  AOI22X1 g2819(.A0(n3270), .A1(EBX_REG_13__SCAN_IN), .B0(INSTADDRPOINTER_REG_13__SCAN_IN), .B1(n3273), .Y(n3890));
  XOR2X1  g2820(.A(n3890), .B(n1758), .Y(n3891));
  NOR4X1  g2821(.A(n3794), .B(n3755), .C(n3752), .D(n3853), .Y(n3892));
  XOR2X1  g2822(.A(n3892), .B(n3891), .Y(n3893));
  AOI22X1 g2823(.A0(n3253), .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .B0(REIP_REG_13__SCAN_IN), .B1(n3239), .Y(n3894));
  OAI21X1 g2824(.A0(n3893), .A1(n3408), .B0(n3894), .Y(n3895));
  NAND3X1 g2825(.A(n3790), .B(INSTADDRPOINTER_REG_12__SCAN_IN), .C(INSTADDRPOINTER_REG_11__SCAN_IN), .Y(n3896));
  XOR2X1  g2826(.A(n3896), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .Y(n3897));
  NOR2X1  g2827(.A(n3897), .B(n3266), .Y(n3898));
  NOR3X1  g2828(.A(n3797), .B(n3844), .C(n3762), .Y(n3899));
  XOR2X1  g2829(.A(n3899), .B(n3861), .Y(n3900));
  NAND2X1 g2830(.A(n3845), .B(INSTADDRPOINTER_REG_12__SCAN_IN), .Y(n3901));
  XOR2X1  g2831(.A(n3901), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .Y(n3902));
  OAI22X1 g2832(.A0(n3900), .A1(n3354), .B0(n3344), .B1(n3902), .Y(n3903));
  NOR3X1  g2833(.A(n3903), .B(n3898), .C(n3895), .Y(n3904));
  OAI21X1 g2834(.A0(n3889), .A1(n3250), .B0(n3904), .Y(U3005));
  AOI22X1 g2835(.A0(n1279), .A1(INSTQUEUE_REG_0__6__SCAN_IN), .B0(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n1268), .Y(n3906));
  AOI22X1 g2836(.A0(n1337), .A1(INSTQUEUE_REG_3__6__SCAN_IN), .B0(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n1244), .Y(n3907));
  AOI22X1 g2837(.A0(n1246), .A1(INSTQUEUE_REG_4__6__SCAN_IN), .B0(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n1273), .Y(n3908));
  AOI22X1 g2838(.A0(n1270), .A1(INSTQUEUE_REG_7__6__SCAN_IN), .B0(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n1329), .Y(n3909));
  NAND4X1 g2839(.A(n3908), .B(n3907), .C(n3906), .D(n3909), .Y(n3910));
  AOI22X1 g2840(.A0(n1255), .A1(INSTQUEUE_REG_12__6__SCAN_IN), .B0(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n1253), .Y(n3911));
  AOI22X1 g2841(.A0(n1266), .A1(INSTQUEUE_REG_15__6__SCAN_IN), .B0(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n1271), .Y(n3912));
  AOI22X1 g2842(.A0(n1278), .A1(INSTQUEUE_REG_8__6__SCAN_IN), .B0(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n1323), .Y(n3913));
  AOI22X1 g2843(.A0(n1275), .A1(INSTQUEUE_REG_11__6__SCAN_IN), .B0(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n1338), .Y(n3914));
  NAND4X1 g2844(.A(n3913), .B(n3912), .C(n3911), .D(n3914), .Y(n3915));
  OAI21X1 g2845(.A0(n3915), .A1(n3910), .B0(n3616), .Y(n3916));
  XOR2X1  g2846(.A(n3916), .B(n2167), .Y(n3917));
  NOR2X1  g2847(.A(n3873), .B(n3813), .Y(n3918));
  INVX1   g2848(.A(n3918), .Y(n3919));
  NOR3X1  g2849(.A(n3919), .B(n3816), .C(n3627), .Y(n3920));
  XOR2X1  g2850(.A(n3920), .B(n3917), .Y(n3921));
  NOR2X1  g2851(.A(n3921), .B(n1473), .Y(n3922));
  XOR2X1  g2852(.A(n3922), .B(INSTADDRPOINTER_REG_14__SCAN_IN), .Y(n3923));
  INVX1   g2853(.A(n3879), .Y(n3924));
  AOI21X1 g2854(.A0(n3888), .A1(n3876), .B0(n3924), .Y(n3925));
  XOR2X1  g2855(.A(n3925), .B(n3923), .Y(n3926));
  AOI22X1 g2856(.A0(n3270), .A1(EBX_REG_14__SCAN_IN), .B0(INSTADDRPOINTER_REG_14__SCAN_IN), .B1(n3273), .Y(n3927));
  XOR2X1  g2857(.A(n3927), .B(n1758), .Y(n3928));
  INVX1   g2858(.A(n3928), .Y(n3929));
  NOR2X1  g2859(.A(n3891), .B(n3853), .Y(n3930));
  NAND2X1 g2860(.A(n3930), .B(n3854), .Y(n3931));
  XOR2X1  g2861(.A(n3931), .B(n3929), .Y(n3932));
  AOI22X1 g2862(.A0(n3253), .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .B0(REIP_REG_14__SCAN_IN), .B1(n3239), .Y(n3933));
  OAI21X1 g2863(.A0(n3932), .A1(n3408), .B0(n3933), .Y(n3934));
  NAND4X1 g2864(.A(INSTADDRPOINTER_REG_13__SCAN_IN), .B(INSTADDRPOINTER_REG_12__SCAN_IN), .C(INSTADDRPOINTER_REG_11__SCAN_IN), .D(n3790), .Y(n3935));
  XOR2X1  g2865(.A(n3935), .B(INSTADDRPOINTER_REG_14__SCAN_IN), .Y(n3936));
  NOR2X1  g2866(.A(n3936), .B(n3266), .Y(n3937));
  INVX1   g2867(.A(INSTADDRPOINTER_REG_14__SCAN_IN), .Y(n3938));
  NOR4X1  g2868(.A(n3861), .B(n3844), .C(n3762), .D(n3797), .Y(n3939));
  XOR2X1  g2869(.A(n3939), .B(n3938), .Y(n3940));
  NAND3X1 g2870(.A(n3845), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .C(INSTADDRPOINTER_REG_12__SCAN_IN), .Y(n3941));
  XOR2X1  g2871(.A(n3941), .B(INSTADDRPOINTER_REG_14__SCAN_IN), .Y(n3942));
  OAI22X1 g2872(.A0(n3940), .A1(n3354), .B0(n3344), .B1(n3942), .Y(n3943));
  NOR3X1  g2873(.A(n3943), .B(n3937), .C(n3934), .Y(n3944));
  OAI21X1 g2874(.A0(n3926), .A1(n3250), .B0(n3944), .Y(U3004));
  INVX1   g2875(.A(INSTADDRPOINTER_REG_15__SCAN_IN), .Y(n3946));
  AOI22X1 g2876(.A0(n1279), .A1(INSTQUEUE_REG_0__7__SCAN_IN), .B0(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n1268), .Y(n3947));
  AOI22X1 g2877(.A0(n1337), .A1(INSTQUEUE_REG_3__7__SCAN_IN), .B0(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n1244), .Y(n3948));
  AOI22X1 g2878(.A0(n1246), .A1(INSTQUEUE_REG_4__7__SCAN_IN), .B0(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n1273), .Y(n3949));
  AOI22X1 g2879(.A0(n1270), .A1(INSTQUEUE_REG_7__7__SCAN_IN), .B0(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n1329), .Y(n3950));
  NAND4X1 g2880(.A(n3949), .B(n3948), .C(n3947), .D(n3950), .Y(n3951));
  AOI22X1 g2881(.A0(n1255), .A1(INSTQUEUE_REG_12__7__SCAN_IN), .B0(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n1253), .Y(n3952));
  AOI22X1 g2882(.A0(n1266), .A1(INSTQUEUE_REG_15__7__SCAN_IN), .B0(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n1271), .Y(n3953));
  AOI22X1 g2883(.A0(n1278), .A1(INSTQUEUE_REG_8__7__SCAN_IN), .B0(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n1323), .Y(n3954));
  AOI22X1 g2884(.A0(n1275), .A1(INSTQUEUE_REG_11__7__SCAN_IN), .B0(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n1338), .Y(n3955));
  NAND4X1 g2885(.A(n3954), .B(n3953), .C(n3952), .D(n3955), .Y(n3956));
  OAI21X1 g2886(.A0(n3956), .A1(n3951), .B0(n3616), .Y(n3957));
  XOR2X1  g2887(.A(n3957), .B(n2167), .Y(n3958));
  NOR4X1  g2888(.A(n3917), .B(n3816), .C(n3627), .D(n3919), .Y(n3959));
  XOR2X1  g2889(.A(n3959), .B(n3958), .Y(n3960));
  OAI21X1 g2890(.A0(n3960), .A1(n1473), .B0(n3946), .Y(n3961));
  INVX1   g2891(.A(n3958), .Y(n3962));
  XOR2X1  g2892(.A(n3959), .B(n3962), .Y(n3963));
  NAND3X1 g2893(.A(n3963), .B(n1472), .C(INSTADDRPOINTER_REG_15__SCAN_IN), .Y(n3964));
  NAND2X1 g2894(.A(n3964), .B(n3961), .Y(n3965));
  INVX1   g2895(.A(n3917), .Y(n3966));
  XOR2X1  g2896(.A(n3920), .B(n3966), .Y(n3967));
  NAND3X1 g2897(.A(n3967), .B(n1472), .C(INSTADDRPOINTER_REG_14__SCAN_IN), .Y(n3968));
  AOI21X1 g2898(.A0(n3967), .A1(n1472), .B0(INSTADDRPOINTER_REG_14__SCAN_IN), .Y(n3969));
  OAI21X1 g2899(.A0(n3925), .A1(n3969), .B0(n3968), .Y(n3970));
  XOR2X1  g2900(.A(n3970), .B(n3965), .Y(n3971));
  AOI22X1 g2901(.A0(n3270), .A1(EBX_REG_15__SCAN_IN), .B0(INSTADDRPOINTER_REG_15__SCAN_IN), .B1(n3273), .Y(n3972));
  XOR2X1  g2902(.A(n3972), .B(n1758), .Y(n3973));
  NOR2X1  g2903(.A(n3931), .B(n3928), .Y(n3974));
  XOR2X1  g2904(.A(n3974), .B(n3973), .Y(n3975));
  AOI22X1 g2905(.A0(n3253), .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .B0(REIP_REG_15__SCAN_IN), .B1(n3239), .Y(n3976));
  OAI21X1 g2906(.A0(n3975), .A1(n3408), .B0(n3976), .Y(n3977));
  NOR3X1  g2907(.A(n3896), .B(n3938), .C(n3861), .Y(n3978));
  XOR2X1  g2908(.A(n3978), .B(n3946), .Y(n3979));
  NOR2X1  g2909(.A(n3979), .B(n3266), .Y(n3980));
  NAND2X1 g2910(.A(n3939), .B(INSTADDRPOINTER_REG_14__SCAN_IN), .Y(n3981));
  XOR2X1  g2911(.A(n3981), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .Y(n3982));
  NAND4X1 g2912(.A(INSTADDRPOINTER_REG_14__SCAN_IN), .B(INSTADDRPOINTER_REG_13__SCAN_IN), .C(INSTADDRPOINTER_REG_12__SCAN_IN), .D(n3845), .Y(n3983));
  XOR2X1  g2913(.A(n3983), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .Y(n3984));
  OAI22X1 g2914(.A0(n3982), .A1(n3354), .B0(n3344), .B1(n3984), .Y(n3985));
  NOR3X1  g2915(.A(n3985), .B(n3980), .C(n3977), .Y(n3986));
  OAI21X1 g2916(.A0(n3971), .A1(n3250), .B0(n3986), .Y(U3003));
  INVX1   g2917(.A(INSTADDRPOINTER_REG_16__SCAN_IN), .Y(n3988));
  NOR4X1  g2918(.A(n3917), .B(n3873), .C(n3813), .D(n3958), .Y(n3989));
  INVX1   g2919(.A(n3989), .Y(n3990));
  NOR2X1  g2920(.A(n3990), .B(n3816), .Y(n3991));
  INVX1   g2921(.A(n3991), .Y(n3992));
  XOR2X1  g2922(.A(n4084), .B(n3988), .Y(n3996));
  AOI21X1 g2923(.A0(n3878), .A1(n1472), .B0(INSTADDRPOINTER_REG_13__SCAN_IN), .Y(n3997));
  AOI21X1 g2924(.A0(n3963), .A1(n1472), .B0(INSTADDRPOINTER_REG_15__SCAN_IN), .Y(n3998));
  NOR4X1  g2925(.A(n3969), .B(n3997), .C(n3819), .D(n3998), .Y(n3999));
  NOR3X1  g2926(.A(n3969), .B(n3997), .C(n3821), .Y(n4000));
  NAND2X1 g2927(.A(n4000), .B(n3961), .Y(n4001));
  NOR3X1  g2928(.A(n3998), .B(n3969), .C(n3879), .Y(n4002));
  OAI21X1 g2929(.A0(n3998), .A1(n3968), .B0(n3964), .Y(n4003));
  NOR2X1  g2930(.A(n4003), .B(n4002), .Y(n4004));
  NAND2X1 g2931(.A(n4004), .B(n4001), .Y(n4005));
  AOI21X1 g2932(.A0(n3999), .A1(n3842), .B0(n4005), .Y(n4006));
  XOR2X1  g2933(.A(n4006), .B(n3996), .Y(n4007));
  AOI22X1 g2934(.A0(n3270), .A1(EBX_REG_16__SCAN_IN), .B0(INSTADDRPOINTER_REG_16__SCAN_IN), .B1(n3273), .Y(n4008));
  XOR2X1  g2935(.A(n4008), .B(n1758), .Y(n4009));
  NOR3X1  g2936(.A(n3973), .B(n3931), .C(n3928), .Y(n4010));
  XOR2X1  g2937(.A(n4010), .B(n4009), .Y(n4011));
  AOI22X1 g2938(.A0(n3253), .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .B0(REIP_REG_16__SCAN_IN), .B1(n3239), .Y(n4012));
  OAI21X1 g2939(.A0(n4011), .A1(n3408), .B0(n4012), .Y(n4013));
  NOR4X1  g2940(.A(n3946), .B(n3938), .C(n3861), .D(n3896), .Y(n4014));
  XOR2X1  g2941(.A(n4014), .B(n3988), .Y(n4015));
  NOR2X1  g2942(.A(n4015), .B(n3266), .Y(n4016));
  NAND3X1 g2943(.A(n3939), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .C(INSTADDRPOINTER_REG_14__SCAN_IN), .Y(n4017));
  XOR2X1  g2944(.A(n4017), .B(INSTADDRPOINTER_REG_16__SCAN_IN), .Y(n4018));
  NOR2X1  g2945(.A(n3983), .B(n3946), .Y(n4019));
  XOR2X1  g2946(.A(n4019), .B(n3988), .Y(n4020));
  OAI22X1 g2947(.A0(n4018), .A1(n3354), .B0(n3344), .B1(n4020), .Y(n4021));
  NOR3X1  g2948(.A(n4021), .B(n4016), .C(n4013), .Y(n4022));
  OAI21X1 g2949(.A0(n4007), .A1(n3250), .B0(n4022), .Y(U3002));
  AOI21X1 g2950(.A0(n4058), .A1(n1472), .B0(INSTADDRPOINTER_REG_16__SCAN_IN), .Y(n4024));
  NAND3X1 g2951(.A(n4058), .B(n1472), .C(INSTADDRPOINTER_REG_16__SCAN_IN), .Y(n4025));
  OAI21X1 g2952(.A0(n4006), .A1(n4024), .B0(n4025), .Y(n4026));
  INVX1   g2953(.A(INSTADDRPOINTER_REG_17__SCAN_IN), .Y(n4027));
  OAI21X1 g2954(.A0(n3992), .A1(n3627), .B0(n2167), .Y(n4028));
  NOR2X1  g2955(.A(n4028), .B(n1473), .Y(n4029));
  XOR2X1  g2956(.A(n4029), .B(n4027), .Y(n4030));
  XOR2X1  g2957(.A(n4030), .B(n4026), .Y(n4031));
  AOI22X1 g2958(.A0(n3270), .A1(EBX_REG_17__SCAN_IN), .B0(INSTADDRPOINTER_REG_17__SCAN_IN), .B1(n3273), .Y(n4032));
  XOR2X1  g2959(.A(n4032), .B(n1758), .Y(n4033));
  NOR4X1  g2960(.A(n3973), .B(n3931), .C(n3928), .D(n4009), .Y(n4034));
  XOR2X1  g2961(.A(n4034), .B(n4033), .Y(n4035));
  AOI22X1 g2962(.A0(n3253), .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .B0(REIP_REG_17__SCAN_IN), .B1(n3239), .Y(n4036));
  OAI21X1 g2963(.A0(n4035), .A1(n3408), .B0(n4036), .Y(n4037));
  NAND2X1 g2964(.A(INSTADDRPOINTER_REG_16__SCAN_IN), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .Y(n4038));
  NOR4X1  g2965(.A(n3896), .B(n3938), .C(n3861), .D(n4038), .Y(n4039));
  XOR2X1  g2966(.A(n4039), .B(n4027), .Y(n4040));
  NOR2X1  g2967(.A(n4040), .B(n3266), .Y(n4041));
  NAND4X1 g2968(.A(INSTADDRPOINTER_REG_16__SCAN_IN), .B(INSTADDRPOINTER_REG_15__SCAN_IN), .C(INSTADDRPOINTER_REG_14__SCAN_IN), .D(n3939), .Y(n4042));
  XOR2X1  g2969(.A(n4042), .B(INSTADDRPOINTER_REG_17__SCAN_IN), .Y(n4043));
  NOR3X1  g2970(.A(n3983), .B(n3988), .C(n3946), .Y(n4044));
  XOR2X1  g2971(.A(n4044), .B(n4027), .Y(n4045));
  OAI22X1 g2972(.A0(n4043), .A1(n3354), .B0(n3344), .B1(n4045), .Y(n4046));
  NOR3X1  g2973(.A(n4046), .B(n4041), .C(n4037), .Y(n4047));
  OAI21X1 g2974(.A0(n4031), .A1(n3250), .B0(n4047), .Y(U3001));
  INVX1   g2975(.A(n3999), .Y(n4049));
  NOR4X1  g2976(.A(n3969), .B(n3997), .C(n3821), .D(n3998), .Y(n4050));
  NOR3X1  g2977(.A(n4003), .B(n4002), .C(n4050), .Y(n4051));
  OAI21X1 g2978(.A0(n4049), .A1(n3887), .B0(n4051), .Y(n4052));
  NOR3X1  g2979(.A(n4028), .B(n1473), .C(n4027), .Y(n4053));
  INVX1   g2980(.A(n4053), .Y(n4054));
  NAND2X1 g2981(.A(n4025), .B(n4054), .Y(n4057));
  AOI21X1 g2982(.A0(n3991), .A1(n3836), .B0(n2166), .Y(n4058));
  AOI21X1 g2983(.A0(n4058), .A1(n1472), .B0(INSTADDRPOINTER_REG_17__SCAN_IN), .Y(n4059));
  NOR2X1  g2984(.A(n4059), .B(n4024), .Y(n4060));
  AOI21X1 g2985(.A0(n4060), .A1(n4052), .B0(n4057), .Y(n4061));
  XOR2X1  g2986(.A(n4029), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .Y(n4062));
  XOR2X1  g2987(.A(n4062), .B(n4061), .Y(n4063));
  AOI22X1 g2988(.A0(n3270), .A1(EBX_REG_18__SCAN_IN), .B0(INSTADDRPOINTER_REG_18__SCAN_IN), .B1(n3273), .Y(n4064));
  XOR2X1  g2989(.A(n4064), .B(n1758), .Y(n4065));
  INVX1   g2990(.A(n4065), .Y(n4066));
  NOR2X1  g2991(.A(n4033), .B(n4009), .Y(n4067));
  NAND2X1 g2992(.A(n4067), .B(n4010), .Y(n4068));
  XOR2X1  g2993(.A(n4068), .B(n4066), .Y(n4069));
  AOI22X1 g2994(.A0(n3253), .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .B0(REIP_REG_18__SCAN_IN), .B1(n3239), .Y(n4070));
  OAI21X1 g2995(.A0(n4069), .A1(n3408), .B0(n4070), .Y(n4071));
  NAND2X1 g2996(.A(n4039), .B(INSTADDRPOINTER_REG_17__SCAN_IN), .Y(n4072));
  XOR2X1  g2997(.A(n4072), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .Y(n4073));
  NOR2X1  g2998(.A(n4073), .B(n3266), .Y(n4074));
  INVX1   g2999(.A(INSTADDRPOINTER_REG_18__SCAN_IN), .Y(n4075));
  NOR2X1  g3000(.A(n4042), .B(n4027), .Y(n4076));
  XOR2X1  g3001(.A(n4076), .B(n4075), .Y(n4077));
  NOR4X1  g3002(.A(n4027), .B(n3988), .C(n3946), .D(n3983), .Y(n4078));
  XOR2X1  g3003(.A(n4078), .B(n4075), .Y(n4079));
  OAI22X1 g3004(.A0(n4077), .A1(n3354), .B0(n3344), .B1(n4079), .Y(n4080));
  NOR3X1  g3005(.A(n4080), .B(n4074), .C(n4071), .Y(n4081));
  OAI21X1 g3006(.A0(n4063), .A1(n3250), .B0(n4081), .Y(U3000));
  NOR3X1  g3007(.A(n4028), .B(n1473), .C(n4075), .Y(n4083));
  NAND2X1 g3008(.A(n4058), .B(n1472), .Y(n4084));
  NOR2X1  g3009(.A(n4057), .B(n4083), .Y(n4086));
  OAI21X1 g3010(.A0(n4028), .A1(n1473), .B0(n4075), .Y(n4087));
  NAND2X1 g3011(.A(n4087), .B(n4060), .Y(n4088));
  OAI21X1 g3012(.A0(n4088), .A1(n4006), .B0(n4086), .Y(n4089));
  INVX1   g3013(.A(INSTADDRPOINTER_REG_19__SCAN_IN), .Y(n4090));
  XOR2X1  g3014(.A(n4029), .B(n4090), .Y(n4091));
  XOR2X1  g3015(.A(n4091), .B(n4089), .Y(n4092));
  AOI22X1 g3016(.A0(n3270), .A1(EBX_REG_19__SCAN_IN), .B0(INSTADDRPOINTER_REG_19__SCAN_IN), .B1(n3273), .Y(n4093));
  XOR2X1  g3017(.A(n4093), .B(n1758), .Y(n4094));
  NOR2X1  g3018(.A(n4068), .B(n4065), .Y(n4095));
  XOR2X1  g3019(.A(n4095), .B(n4094), .Y(n4096));
  AOI22X1 g3020(.A0(n3253), .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .B0(REIP_REG_19__SCAN_IN), .B1(n3239), .Y(n4097));
  OAI21X1 g3021(.A0(n4096), .A1(n3408), .B0(n4097), .Y(n4098));
  NAND3X1 g3022(.A(n4039), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .C(INSTADDRPOINTER_REG_17__SCAN_IN), .Y(n4099));
  XOR2X1  g3023(.A(n4099), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .Y(n4100));
  NOR2X1  g3024(.A(n4100), .B(n3266), .Y(n4101));
  NOR3X1  g3025(.A(n4042), .B(n4075), .C(n4027), .Y(n4102));
  XOR2X1  g3026(.A(n4102), .B(n4090), .Y(n4103));
  NAND2X1 g3027(.A(n4078), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .Y(n4104));
  XOR2X1  g3028(.A(n4104), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .Y(n4105));
  OAI22X1 g3029(.A0(n4103), .A1(n3354), .B0(n3344), .B1(n4105), .Y(n4106));
  NOR3X1  g3030(.A(n4106), .B(n4101), .C(n4098), .Y(n4107));
  OAI21X1 g3031(.A0(n4092), .A1(n3250), .B0(n4107), .Y(U2999));
  OAI21X1 g3032(.A0(n4028), .A1(n1473), .B0(n4090), .Y(n4109));
  NAND3X1 g3033(.A(n4109), .B(n4087), .C(n4060), .Y(n4110));
  NOR3X1  g3034(.A(n4028), .B(n1473), .C(n4090), .Y(n4111));
  INVX1   g3035(.A(n4083), .Y(n4112));
  NOR4X1  g3036(.A(n4028), .B(n1473), .C(n3988), .D(n4059), .Y(n4114));
  OAI21X1 g3037(.A0(n4114), .A1(n4053), .B0(n4087), .Y(n4115));
  AOI22X1 g3038(.A0(n4112), .A1(n4115), .B0(n4084), .B1(n4090), .Y(n4116));
  NOR2X1  g3039(.A(n4116), .B(n4111), .Y(n4117));
  OAI21X1 g3040(.A0(n4110), .A1(n4006), .B0(n4117), .Y(n4118));
  XOR2X1  g3041(.A(n4029), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .Y(n4119));
  XOR2X1  g3042(.A(n4119), .B(n4118), .Y(n4120));
  NAND2X1 g3043(.A(n4120), .B(n3251), .Y(n4121));
  AOI22X1 g3044(.A0(n3270), .A1(EBX_REG_20__SCAN_IN), .B0(INSTADDRPOINTER_REG_20__SCAN_IN), .B1(n3273), .Y(n4122));
  XOR2X1  g3045(.A(n4122), .B(n1758), .Y(n4123));
  INVX1   g3046(.A(n4094), .Y(n4124));
  NAND4X1 g3047(.A(n4067), .B(n4066), .C(n4010), .D(n4124), .Y(n4125));
  XOR2X1  g3048(.A(n4125), .B(n4123), .Y(n4126));
  INVX1   g3049(.A(INSTADDRPOINTER_REG_20__SCAN_IN), .Y(n4127));
  OAI22X1 g3050(.A0(n3254), .A1(n4127), .B0(n1052), .B1(n5914), .Y(n4128));
  AOI21X1 g3051(.A0(n4126), .A1(n3278), .B0(n4128), .Y(n4129));
  NAND4X1 g3052(.A(INSTADDRPOINTER_REG_19__SCAN_IN), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .C(INSTADDRPOINTER_REG_17__SCAN_IN), .D(n4039), .Y(n4130));
  XOR2X1  g3053(.A(n4130), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .Y(n4131));
  NOR2X1  g3054(.A(n4131), .B(n3266), .Y(n4132));
  NOR4X1  g3055(.A(n4090), .B(n4075), .C(n4027), .D(n4042), .Y(n4133));
  XOR2X1  g3056(.A(n4133), .B(n4127), .Y(n4134));
  NAND3X1 g3057(.A(n4078), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .C(INSTADDRPOINTER_REG_18__SCAN_IN), .Y(n4135));
  XOR2X1  g3058(.A(n4135), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .Y(n4136));
  OAI22X1 g3059(.A0(n4134), .A1(n3354), .B0(n3344), .B1(n4136), .Y(n4137));
  NOR2X1  g3060(.A(n4137), .B(n4132), .Y(n4138));
  NAND3X1 g3061(.A(n4138), .B(n4129), .C(n4121), .Y(U2998));
  INVX1   g3062(.A(INSTADDRPOINTER_REG_21__SCAN_IN), .Y(n4140));
  XOR2X1  g3063(.A(n4029), .B(n4140), .Y(n4141));
  OAI21X1 g3064(.A0(n4029), .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .B0(n4118), .Y(n4142));
  OAI21X1 g3065(.A0(n4084), .A1(n4127), .B0(n4142), .Y(n4143));
  XOR2X1  g3066(.A(n4143), .B(n4141), .Y(n4144));
  AOI22X1 g3067(.A0(n3270), .A1(EBX_REG_21__SCAN_IN), .B0(INSTADDRPOINTER_REG_21__SCAN_IN), .B1(n3273), .Y(n4145));
  XOR2X1  g3068(.A(n4145), .B(n1758), .Y(n4146));
  NOR2X1  g3069(.A(n4125), .B(n4123), .Y(n4147));
  XOR2X1  g3070(.A(n4147), .B(n4146), .Y(n4148));
  AOI22X1 g3071(.A0(n3253), .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .B0(REIP_REG_21__SCAN_IN), .B1(n3239), .Y(n4149));
  OAI21X1 g3072(.A0(n4148), .A1(n3408), .B0(n4149), .Y(n4150));
  NOR3X1  g3073(.A(n4099), .B(n4127), .C(n4090), .Y(n4151));
  XOR2X1  g3074(.A(n4151), .B(n4140), .Y(n4152));
  NOR2X1  g3075(.A(n4152), .B(n3266), .Y(n4153));
  NAND2X1 g3076(.A(n4133), .B(INSTADDRPOINTER_REG_20__SCAN_IN), .Y(n4154));
  XOR2X1  g3077(.A(n4154), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .Y(n4155));
  NAND4X1 g3078(.A(INSTADDRPOINTER_REG_20__SCAN_IN), .B(INSTADDRPOINTER_REG_19__SCAN_IN), .C(INSTADDRPOINTER_REG_18__SCAN_IN), .D(n4078), .Y(n4156));
  XOR2X1  g3079(.A(n4156), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .Y(n4157));
  OAI22X1 g3080(.A0(n4155), .A1(n3354), .B0(n3344), .B1(n4157), .Y(n4158));
  NOR3X1  g3081(.A(n4158), .B(n4153), .C(n4150), .Y(n4159));
  OAI21X1 g3082(.A0(n4144), .A1(n3250), .B0(n4159), .Y(U2997));
  XOR2X1  g3083(.A(n4029), .B(INSTADDRPOINTER_REG_22__SCAN_IN), .Y(n4161));
  INVX1   g3084(.A(n4110), .Y(n4162));
  INVX1   g3085(.A(n4111), .Y(n4163));
  NAND2X1 g3086(.A(n4086), .B(n4163), .Y(n4165));
  AOI21X1 g3087(.A0(n4162), .A1(n4052), .B0(n4165), .Y(n4166));
  AOI21X1 g3088(.A0(n4140), .A1(n4127), .B0(n4084), .Y(n4167));
  INVX1   g3089(.A(n4167), .Y(n4168));
  AOI22X1 g3090(.A0(n1472), .A1(n4058), .B0(INSTADDRPOINTER_REG_21__SCAN_IN), .B1(INSTADDRPOINTER_REG_20__SCAN_IN), .Y(n4169));
  OAI21X1 g3091(.A0(n4169), .A1(n4166), .B0(n4168), .Y(n4170));
  XOR2X1  g3092(.A(n4170), .B(n4161), .Y(n4171));
  NAND2X1 g3093(.A(n4171), .B(n3251), .Y(n4172));
  AOI22X1 g3094(.A0(n3270), .A1(EBX_REG_22__SCAN_IN), .B0(INSTADDRPOINTER_REG_22__SCAN_IN), .B1(n3273), .Y(n4173));
  XOR2X1  g3095(.A(n4173), .B(n1758), .Y(n4174));
  NOR3X1  g3096(.A(n4146), .B(n4125), .C(n4123), .Y(n4175));
  XOR2X1  g3097(.A(n4175), .B(n4174), .Y(n4176));
  AOI22X1 g3098(.A0(n3253), .A1(INSTADDRPOINTER_REG_22__SCAN_IN), .B0(REIP_REG_22__SCAN_IN), .B1(n3239), .Y(n4177));
  OAI21X1 g3099(.A0(n4176), .A1(n3408), .B0(n4177), .Y(n4178));
  INVX1   g3100(.A(INSTADDRPOINTER_REG_22__SCAN_IN), .Y(n4179));
  NOR4X1  g3101(.A(n4140), .B(n4127), .C(n4090), .D(n4099), .Y(n4180));
  XOR2X1  g3102(.A(n4180), .B(n4179), .Y(n4181));
  NOR2X1  g3103(.A(n4181), .B(n3266), .Y(n4182));
  NAND3X1 g3104(.A(n4133), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .C(INSTADDRPOINTER_REG_20__SCAN_IN), .Y(n4183));
  XOR2X1  g3105(.A(n4183), .B(INSTADDRPOINTER_REG_22__SCAN_IN), .Y(n4184));
  NOR2X1  g3106(.A(n4156), .B(n4140), .Y(n4185));
  XOR2X1  g3107(.A(n4185), .B(n4179), .Y(n4186));
  OAI22X1 g3108(.A0(n4184), .A1(n3354), .B0(n3344), .B1(n4186), .Y(n4187));
  NOR3X1  g3109(.A(n4187), .B(n4182), .C(n4178), .Y(n4188));
  NAND2X1 g3110(.A(n4188), .B(n4172), .Y(U2996));
  INVX1   g3111(.A(INSTADDRPOINTER_REG_23__SCAN_IN), .Y(n4190));
  XOR2X1  g3112(.A(n4029), .B(n4190), .Y(n4191));
  NOR3X1  g3113(.A(n4028), .B(n1473), .C(n4179), .Y(n4192));
  OAI21X1 g3114(.A0(n4028), .A1(n1473), .B0(n4179), .Y(n4193));
  AOI21X1 g3115(.A0(n4167), .A1(n4193), .B0(n4192), .Y(n4194));
  OAI22X1 g3116(.A0(n1473), .A1(n4028), .B0(n4140), .B1(n4127), .Y(n4195));
  NAND2X1 g3117(.A(n4195), .B(n4193), .Y(n4196));
  OAI21X1 g3118(.A0(n4196), .A1(n4166), .B0(n4194), .Y(n4197));
  XOR2X1  g3119(.A(n4197), .B(n4191), .Y(n4198));
  AOI22X1 g3120(.A0(n3270), .A1(EBX_REG_23__SCAN_IN), .B0(INSTADDRPOINTER_REG_23__SCAN_IN), .B1(n3273), .Y(n4199));
  XOR2X1  g3121(.A(n4199), .B(n1758), .Y(n4200));
  NOR4X1  g3122(.A(n4146), .B(n4125), .C(n4123), .D(n4174), .Y(n4201));
  XOR2X1  g3123(.A(n4201), .B(n4200), .Y(n4202));
  AOI22X1 g3124(.A0(n3253), .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .B0(REIP_REG_23__SCAN_IN), .B1(n3239), .Y(n4203));
  OAI21X1 g3125(.A0(n4202), .A1(n3408), .B0(n4203), .Y(n4204));
  NAND3X1 g3126(.A(n4151), .B(INSTADDRPOINTER_REG_22__SCAN_IN), .C(INSTADDRPOINTER_REG_21__SCAN_IN), .Y(n4205));
  XOR2X1  g3127(.A(n4205), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .Y(n4206));
  NOR2X1  g3128(.A(n4206), .B(n3266), .Y(n4207));
  NAND4X1 g3129(.A(INSTADDRPOINTER_REG_22__SCAN_IN), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .C(INSTADDRPOINTER_REG_20__SCAN_IN), .D(n4133), .Y(n4208));
  XOR2X1  g3130(.A(n4208), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .Y(n4209));
  NOR3X1  g3131(.A(n4156), .B(n4179), .C(n4140), .Y(n4210));
  XOR2X1  g3132(.A(n4210), .B(n4190), .Y(n4211));
  OAI22X1 g3133(.A0(n4209), .A1(n3354), .B0(n3344), .B1(n4211), .Y(n4212));
  NOR3X1  g3134(.A(n4212), .B(n4207), .C(n4204), .Y(n4213));
  OAI21X1 g3135(.A0(n4198), .A1(n3250), .B0(n4213), .Y(U2995));
  XOR2X1  g3136(.A(n4029), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .Y(n4215));
  NAND3X1 g3137(.A(n4058), .B(n1472), .C(INSTADDRPOINTER_REG_23__SCAN_IN), .Y(n4216));
  AOI21X1 g3138(.A0(n4058), .A1(n1472), .B0(INSTADDRPOINTER_REG_23__SCAN_IN), .Y(n4217));
  OAI21X1 g3139(.A0(n4194), .A1(n4217), .B0(n4216), .Y(n4218));
  AOI21X1 g3140(.A0(n4058), .A1(n1472), .B0(INSTADDRPOINTER_REG_22__SCAN_IN), .Y(n4219));
  NOR3X1  g3141(.A(n4217), .B(n4169), .C(n4219), .Y(n4220));
  AOI21X1 g3142(.A0(n4220), .A1(n4118), .B0(n4218), .Y(n4221));
  XOR2X1  g3143(.A(n4221), .B(n4215), .Y(n4222));
  AOI22X1 g3144(.A0(n3270), .A1(EBX_REG_24__SCAN_IN), .B0(INSTADDRPOINTER_REG_24__SCAN_IN), .B1(n3273), .Y(n4223));
  XOR2X1  g3145(.A(n4223), .B(n1758), .Y(n4224));
  INVX1   g3146(.A(n4201), .Y(n4225));
  NOR2X1  g3147(.A(n4225), .B(n4200), .Y(n4226));
  XOR2X1  g3148(.A(n4226), .B(n4224), .Y(n4227));
  AOI22X1 g3149(.A0(n3253), .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .B0(REIP_REG_24__SCAN_IN), .B1(n3239), .Y(n4228));
  OAI21X1 g3150(.A0(n4227), .A1(n3408), .B0(n4228), .Y(n4229));
  NAND4X1 g3151(.A(INSTADDRPOINTER_REG_23__SCAN_IN), .B(INSTADDRPOINTER_REG_22__SCAN_IN), .C(INSTADDRPOINTER_REG_21__SCAN_IN), .D(n4151), .Y(n4230));
  XOR2X1  g3152(.A(n4230), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .Y(n4231));
  NOR2X1  g3153(.A(n4231), .B(n3266), .Y(n4232));
  INVX1   g3154(.A(INSTADDRPOINTER_REG_24__SCAN_IN), .Y(n4233));
  NOR2X1  g3155(.A(n4208), .B(n4190), .Y(n4234));
  XOR2X1  g3156(.A(n4234), .B(n4233), .Y(n4235));
  NOR4X1  g3157(.A(n4190), .B(n4179), .C(n4140), .D(n4156), .Y(n4236));
  XOR2X1  g3158(.A(n4236), .B(n4233), .Y(n4237));
  OAI22X1 g3159(.A0(n4235), .A1(n3354), .B0(n3344), .B1(n4237), .Y(n4238));
  NOR3X1  g3160(.A(n4238), .B(n4232), .C(n4229), .Y(n4239));
  OAI21X1 g3161(.A0(n4222), .A1(n3250), .B0(n4239), .Y(U2994));
  XOR2X1  g3162(.A(n4029), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .Y(n4241));
  NOR3X1  g3163(.A(n4028), .B(n1473), .C(n4233), .Y(n4242));
  AOI21X1 g3164(.A0(n4058), .A1(n1472), .B0(INSTADDRPOINTER_REG_24__SCAN_IN), .Y(n4243));
  INVX1   g3165(.A(n4243), .Y(n4244));
  AOI21X1 g3166(.A0(n4218), .A1(n4244), .B0(n4242), .Y(n4245));
  INVX1   g3167(.A(n4245), .Y(n4246));
  NOR4X1  g3168(.A(n4217), .B(n4169), .C(n4219), .D(n4243), .Y(n4247));
  AOI21X1 g3169(.A0(n4247), .A1(n4118), .B0(n4246), .Y(n4248));
  XOR2X1  g3170(.A(n4248), .B(n4241), .Y(n4249));
  AOI22X1 g3171(.A0(n3270), .A1(EBX_REG_25__SCAN_IN), .B0(INSTADDRPOINTER_REG_25__SCAN_IN), .B1(n3273), .Y(n4250));
  XOR2X1  g3172(.A(n4250), .B(n1758), .Y(n4251));
  INVX1   g3173(.A(n4251), .Y(n4252));
  NOR3X1  g3174(.A(n4224), .B(n4225), .C(n4200), .Y(n4253));
  XOR2X1  g3175(.A(n4253), .B(n4252), .Y(n4254));
  NAND2X1 g3176(.A(n4254), .B(n3278), .Y(n4255));
  AOI22X1 g3177(.A0(n3253), .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .B0(REIP_REG_25__SCAN_IN), .B1(n3239), .Y(n4256));
  NAND2X1 g3178(.A(n4256), .B(n4255), .Y(n4257));
  INVX1   g3179(.A(INSTADDRPOINTER_REG_25__SCAN_IN), .Y(n4258));
  NOR3X1  g3180(.A(n4205), .B(n4233), .C(n4190), .Y(n4259));
  XOR2X1  g3181(.A(n4259), .B(n4258), .Y(n4260));
  NOR2X1  g3182(.A(n4260), .B(n3266), .Y(n4261));
  NOR3X1  g3183(.A(n4208), .B(n4233), .C(n4190), .Y(n4262));
  XOR2X1  g3184(.A(n4262), .B(n4258), .Y(n4263));
  NAND2X1 g3185(.A(n4236), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .Y(n4264));
  XOR2X1  g3186(.A(n4264), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .Y(n4265));
  OAI22X1 g3187(.A0(n4263), .A1(n3354), .B0(n3344), .B1(n4265), .Y(n4266));
  NOR3X1  g3188(.A(n4266), .B(n4261), .C(n4257), .Y(n4267));
  OAI21X1 g3189(.A0(n4249), .A1(n3250), .B0(n4267), .Y(U2993));
  OAI21X1 g3190(.A0(n4029), .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .B0(n4247), .Y(n4269));
  NOR2X1  g3191(.A(n4269), .B(n4110), .Y(n4270));
  AOI21X1 g3192(.A0(n4058), .A1(n1472), .B0(INSTADDRPOINTER_REG_25__SCAN_IN), .Y(n4271));
  NOR4X1  g3193(.A(n4243), .B(n4196), .C(n4217), .D(n4271), .Y(n4272));
  OAI22X1 g3194(.A0(n4163), .A1(n4269), .B0(n4084), .B1(n4258), .Y(n4273));
  AOI21X1 g3195(.A0(n4272), .A1(n4116), .B0(n4273), .Y(n4274));
  OAI21X1 g3196(.A0(n4245), .A1(n4271), .B0(n4274), .Y(n4275));
  AOI21X1 g3197(.A0(n4270), .A1(n4052), .B0(n4275), .Y(n4276));
  XOR2X1  g3198(.A(n4029), .B(INSTADDRPOINTER_REG_26__SCAN_IN), .Y(n4277));
  XOR2X1  g3199(.A(n4277), .B(n4276), .Y(n4278));
  AOI22X1 g3200(.A0(n3270), .A1(EBX_REG_26__SCAN_IN), .B0(INSTADDRPOINTER_REG_26__SCAN_IN), .B1(n3273), .Y(n4279));
  XOR2X1  g3201(.A(n4279), .B(n1758), .Y(n4280));
  NOR4X1  g3202(.A(n4224), .B(n4225), .C(n4200), .D(n4251), .Y(n4281));
  XOR2X1  g3203(.A(n4281), .B(n4280), .Y(n4282));
  NOR4X1  g3204(.A(n3277), .B(n3253), .C(n1833), .D(n4282), .Y(n4283));
  INVX1   g3205(.A(INSTADDRPOINTER_REG_26__SCAN_IN), .Y(n4284));
  NOR4X1  g3206(.A(n4258), .B(n4233), .C(n4190), .D(n4205), .Y(n4285));
  XOR2X1  g3207(.A(n4285), .B(n4284), .Y(n4286));
  AOI22X1 g3208(.A0(n3253), .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .B0(REIP_REG_26__SCAN_IN), .B1(n3239), .Y(n4287));
  OAI21X1 g3209(.A0(n4286), .A1(n3266), .B0(n4287), .Y(n4288));
  NOR4X1  g3210(.A(n4258), .B(n4233), .C(n4190), .D(n4208), .Y(n4289));
  XOR2X1  g3211(.A(n4289), .B(n4284), .Y(n4290));
  NAND3X1 g3212(.A(n4236), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .C(INSTADDRPOINTER_REG_24__SCAN_IN), .Y(n4291));
  XOR2X1  g3213(.A(n4291), .B(INSTADDRPOINTER_REG_26__SCAN_IN), .Y(n4292));
  OAI22X1 g3214(.A0(n4290), .A1(n3354), .B0(n3344), .B1(n4292), .Y(n4293));
  NOR3X1  g3215(.A(n4293), .B(n4288), .C(n4283), .Y(n4294));
  OAI21X1 g3216(.A0(n4278), .A1(n3250), .B0(n4294), .Y(U2992));
  XOR2X1  g3217(.A(n4029), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .Y(n4296));
  AOI21X1 g3218(.A0(n4058), .A1(n1472), .B0(INSTADDRPOINTER_REG_26__SCAN_IN), .Y(n4297));
  NAND3X1 g3219(.A(n4058), .B(n1472), .C(INSTADDRPOINTER_REG_26__SCAN_IN), .Y(n4298));
  OAI21X1 g3220(.A0(n4297), .A1(n4276), .B0(n4298), .Y(n4299));
  XOR2X1  g3221(.A(n4299), .B(n4296), .Y(n4300));
  NAND2X1 g3222(.A(n4300), .B(n3251), .Y(n4301));
  AOI22X1 g3223(.A0(n3270), .A1(EBX_REG_27__SCAN_IN), .B0(INSTADDRPOINTER_REG_27__SCAN_IN), .B1(n3273), .Y(n4302));
  XOR2X1  g3224(.A(n4302), .B(n1758), .Y(n4303));
  INVX1   g3225(.A(n4280), .Y(n4304));
  NAND2X1 g3226(.A(n4281), .B(n4304), .Y(n4305));
  XOR2X1  g3227(.A(n4305), .B(n4303), .Y(n4306));
  NAND2X1 g3228(.A(n4306), .B(n3278), .Y(n4307));
  NAND3X1 g3229(.A(n4259), .B(INSTADDRPOINTER_REG_26__SCAN_IN), .C(INSTADDRPOINTER_REG_25__SCAN_IN), .Y(n4308));
  XOR2X1  g3230(.A(n4308), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .Y(n4309));
  AOI22X1 g3231(.A0(n3253), .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .B0(REIP_REG_27__SCAN_IN), .B1(n3239), .Y(n4310));
  OAI21X1 g3232(.A0(n4309), .A1(n3266), .B0(n4310), .Y(n4311));
  NAND2X1 g3233(.A(n4289), .B(INSTADDRPOINTER_REG_26__SCAN_IN), .Y(n4312));
  XOR2X1  g3234(.A(n4312), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .Y(n4313));
  NAND4X1 g3235(.A(INSTADDRPOINTER_REG_26__SCAN_IN), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .C(INSTADDRPOINTER_REG_24__SCAN_IN), .D(n4236), .Y(n4314));
  XOR2X1  g3236(.A(n4314), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .Y(n4315));
  OAI22X1 g3237(.A0(n4313), .A1(n3354), .B0(n3344), .B1(n4315), .Y(n4316));
  NOR2X1  g3238(.A(n4316), .B(n4311), .Y(n4317));
  NAND3X1 g3239(.A(n4317), .B(n4307), .C(n4301), .Y(U2991));
  INVX1   g3240(.A(INSTADDRPOINTER_REG_28__SCAN_IN), .Y(n4319));
  XOR2X1  g3241(.A(n4029), .B(n4319), .Y(n4320));
  OAI21X1 g3242(.A0(INSTADDRPOINTER_REG_27__SCAN_IN), .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .B0(n4029), .Y(n4321));
  AOI22X1 g3243(.A0(n1472), .A1(n4058), .B0(INSTADDRPOINTER_REG_27__SCAN_IN), .B1(INSTADDRPOINTER_REG_26__SCAN_IN), .Y(n4322));
  OAI21X1 g3244(.A0(n4322), .A1(n4276), .B0(n4321), .Y(n4323));
  XOR2X1  g3245(.A(n4323), .B(n4320), .Y(n4324));
  AOI22X1 g3246(.A0(n3270), .A1(EBX_REG_28__SCAN_IN), .B0(INSTADDRPOINTER_REG_28__SCAN_IN), .B1(n3273), .Y(n4325));
  XOR2X1  g3247(.A(n4325), .B(n1758), .Y(n4326));
  INVX1   g3248(.A(n4326), .Y(n4327));
  INVX1   g3249(.A(n4303), .Y(n4328));
  NAND3X1 g3250(.A(n4328), .B(n4281), .C(n4304), .Y(n4329));
  XOR2X1  g3251(.A(n4329), .B(n4327), .Y(n4330));
  NOR2X1  g3252(.A(n4330), .B(n3408), .Y(n4331));
  NAND4X1 g3253(.A(INSTADDRPOINTER_REG_27__SCAN_IN), .B(INSTADDRPOINTER_REG_26__SCAN_IN), .C(INSTADDRPOINTER_REG_25__SCAN_IN), .D(n4259), .Y(n4332));
  XOR2X1  g3254(.A(n4332), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .Y(n4333));
  AOI22X1 g3255(.A0(n3253), .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .B0(REIP_REG_28__SCAN_IN), .B1(n3239), .Y(n4334));
  OAI21X1 g3256(.A0(n4333), .A1(n3266), .B0(n4334), .Y(n4335));
  NAND3X1 g3257(.A(n4289), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .C(INSTADDRPOINTER_REG_26__SCAN_IN), .Y(n4336));
  XOR2X1  g3258(.A(n4336), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .Y(n4337));
  INVX1   g3259(.A(INSTADDRPOINTER_REG_27__SCAN_IN), .Y(n4338));
  NOR2X1  g3260(.A(n4314), .B(n4338), .Y(n4339));
  XOR2X1  g3261(.A(n4339), .B(n4319), .Y(n4340));
  OAI22X1 g3262(.A0(n4337), .A1(n3354), .B0(n3344), .B1(n4340), .Y(n4341));
  NOR3X1  g3263(.A(n4341), .B(n4335), .C(n4331), .Y(n4342));
  OAI21X1 g3264(.A0(n4324), .A1(n3250), .B0(n4342), .Y(U2990));
  INVX1   g3265(.A(INSTADDRPOINTER_REG_29__SCAN_IN), .Y(n4344));
  XOR2X1  g3266(.A(n4029), .B(n4344), .Y(n4345));
  AOI21X1 g3267(.A0(n4058), .A1(n1472), .B0(INSTADDRPOINTER_REG_28__SCAN_IN), .Y(n4346));
  NOR2X1  g3268(.A(n4346), .B(n4321), .Y(n4347));
  AOI21X1 g3269(.A0(n4029), .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .B0(n4347), .Y(n4348));
  NOR2X1  g3270(.A(n4346), .B(n4322), .Y(n4349));
  INVX1   g3271(.A(n4349), .Y(n4350));
  OAI21X1 g3272(.A0(n4350), .A1(n4276), .B0(n4348), .Y(n4351));
  XOR2X1  g3273(.A(n4351), .B(n4345), .Y(n4352));
  AOI22X1 g3274(.A0(n3270), .A1(EBX_REG_29__SCAN_IN), .B0(INSTADDRPOINTER_REG_29__SCAN_IN), .B1(n3273), .Y(n4353));
  XOR2X1  g3275(.A(n4353), .B(n1758), .Y(n4354));
  NAND4X1 g3276(.A(n4328), .B(n4281), .C(n4304), .D(n4327), .Y(n4355));
  XOR2X1  g3277(.A(n4355), .B(n4354), .Y(n4356));
  INVX1   g3278(.A(n4356), .Y(n4357));
  NOR2X1  g3279(.A(n4357), .B(n3408), .Y(n4358));
  NOR3X1  g3280(.A(n4308), .B(n4319), .C(n4338), .Y(n4359));
  XOR2X1  g3281(.A(n4359), .B(n4344), .Y(n4360));
  AOI22X1 g3282(.A0(n3253), .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .B0(REIP_REG_29__SCAN_IN), .B1(n3239), .Y(n4361));
  OAI21X1 g3283(.A0(n4360), .A1(n3266), .B0(n4361), .Y(n4362));
  NAND4X1 g3284(.A(INSTADDRPOINTER_REG_28__SCAN_IN), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .C(INSTADDRPOINTER_REG_26__SCAN_IN), .D(n4289), .Y(n4363));
  XOR2X1  g3285(.A(n4363), .B(INSTADDRPOINTER_REG_29__SCAN_IN), .Y(n4364));
  NOR3X1  g3286(.A(n4314), .B(n4319), .C(n4338), .Y(n4365));
  XOR2X1  g3287(.A(n4365), .B(n4344), .Y(n4366));
  OAI22X1 g3288(.A0(n4364), .A1(n3354), .B0(n3344), .B1(n4366), .Y(n4367));
  NOR3X1  g3289(.A(n4367), .B(n4362), .C(n4358), .Y(n4368));
  OAI21X1 g3290(.A0(n4352), .A1(n3250), .B0(n4368), .Y(U2989));
  INVX1   g3291(.A(INSTADDRPOINTER_REG_30__SCAN_IN), .Y(n4370));
  XOR2X1  g3292(.A(n4029), .B(n4370), .Y(n4371));
  AOI21X1 g3293(.A0(n4058), .A1(n1472), .B0(INSTADDRPOINTER_REG_29__SCAN_IN), .Y(n4372));
  NOR2X1  g3294(.A(n4372), .B(n4348), .Y(n4373));
  AOI21X1 g3295(.A0(n4029), .A1(INSTADDRPOINTER_REG_29__SCAN_IN), .B0(n4373), .Y(n4374));
  NOR3X1  g3296(.A(n4372), .B(n4346), .C(n4322), .Y(n4375));
  INVX1   g3297(.A(n4375), .Y(n4376));
  OAI21X1 g3298(.A0(n4376), .A1(n4276), .B0(n4374), .Y(n4377));
  XOR2X1  g3299(.A(n4377), .B(n4371), .Y(n4378));
  AOI22X1 g3300(.A0(n3270), .A1(EBX_REG_30__SCAN_IN), .B0(INSTADDRPOINTER_REG_30__SCAN_IN), .B1(n3273), .Y(n4379));
  XOR2X1  g3301(.A(n4379), .B(n1758), .Y(n4380));
  NOR2X1  g3302(.A(n4355), .B(n4354), .Y(n4381));
  XOR2X1  g3303(.A(n4381), .B(n4380), .Y(n4382));
  NOR2X1  g3304(.A(n4382), .B(n3408), .Y(n4383));
  NOR4X1  g3305(.A(n4344), .B(n4319), .C(n4338), .D(n4308), .Y(n4384));
  XOR2X1  g3306(.A(n4384), .B(n4370), .Y(n4385));
  AOI22X1 g3307(.A0(n3253), .A1(INSTADDRPOINTER_REG_30__SCAN_IN), .B0(REIP_REG_30__SCAN_IN), .B1(n3239), .Y(n4386));
  OAI21X1 g3308(.A0(n4385), .A1(n3266), .B0(n4386), .Y(n4387));
  NOR2X1  g3309(.A(n4363), .B(n4344), .Y(n4388));
  XOR2X1  g3310(.A(n4388), .B(n4370), .Y(n4389));
  NOR4X1  g3311(.A(n4344), .B(n4319), .C(n4338), .D(n4314), .Y(n4390));
  XOR2X1  g3312(.A(n4390), .B(n4370), .Y(n4391));
  OAI22X1 g3313(.A0(n4389), .A1(n3354), .B0(n3344), .B1(n4391), .Y(n4392));
  NOR3X1  g3314(.A(n4392), .B(n4387), .C(n4383), .Y(n4393));
  OAI21X1 g3315(.A0(n4378), .A1(n3250), .B0(n4393), .Y(U2988));
  XOR2X1  g3316(.A(n4029), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .Y(n4395));
  AOI21X1 g3317(.A0(n4058), .A1(n1472), .B0(INSTADDRPOINTER_REG_30__SCAN_IN), .Y(n4396));
  NOR3X1  g3318(.A(n4396), .B(n4376), .C(n4276), .Y(n4397));
  NAND3X1 g3319(.A(n4058), .B(n1472), .C(INSTADDRPOINTER_REG_30__SCAN_IN), .Y(n4398));
  OAI21X1 g3320(.A0(n4396), .A1(n4374), .B0(n4398), .Y(n4399));
  NOR2X1  g3321(.A(n4399), .B(n4397), .Y(n4400));
  XOR2X1  g3322(.A(n4400), .B(n4395), .Y(n4401));
  AOI22X1 g3323(.A0(n3270), .A1(EBX_REG_31__SCAN_IN), .B0(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n3273), .Y(n4402));
  XOR2X1  g3324(.A(n4402), .B(n1758), .Y(n4403));
  NOR3X1  g3325(.A(n4380), .B(n4355), .C(n4354), .Y(n4404));
  XOR2X1  g3326(.A(n4404), .B(n4403), .Y(n4405));
  NOR2X1  g3327(.A(n4405), .B(n3408), .Y(n4406));
  NAND2X1 g3328(.A(n4384), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .Y(n4407));
  XOR2X1  g3329(.A(n4407), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .Y(n4408));
  AOI22X1 g3330(.A0(n3253), .A1(INSTADDRPOINTER_REG_31__SCAN_IN), .B0(REIP_REG_31__SCAN_IN), .B1(n3239), .Y(n4409));
  OAI21X1 g3331(.A0(n4408), .A1(n3266), .B0(n4409), .Y(n4410));
  NAND2X1 g3332(.A(n4388), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .Y(n4411));
  XOR2X1  g3333(.A(n4411), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .Y(n4412));
  NAND2X1 g3334(.A(n4390), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .Y(n4413));
  XOR2X1  g3335(.A(n4413), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .Y(n4414));
  OAI22X1 g3336(.A0(n4412), .A1(n3354), .B0(n3344), .B1(n4414), .Y(n4415));
  NOR3X1  g3337(.A(n4415), .B(n4410), .C(n4406), .Y(n4416));
  OAI21X1 g3338(.A0(n4401), .A1(n3250), .B0(n4416), .Y(U2987));
  NOR2X1  g3339(.A(STATE2_REG_2__SCAN_IN), .B(STATEBS16_REG_SCAN_IN), .Y(n4418));
  INVX1   g3340(.A(n4418), .Y(n4419));
  AOI21X1 g3341(.A0(n1700), .A1(STATE2_REG_2__SCAN_IN), .B0(n1671), .Y(n4420));
  AOI21X1 g3342(.A0(n4420), .A1(n2270), .B0(n1833), .Y(n4421));
  OAI21X1 g3343(.A0(n1568), .A1(n1362), .B0(STATE2_REG_2__SCAN_IN), .Y(n4422));
  NOR3X1  g3344(.A(n1700), .B(n1568), .C(n1833), .Y(n4423));
  INVX1   g3345(.A(EAX_REG_0__SCAN_IN), .Y(n4424));
  NOR2X1  g3346(.A(n1615), .B(n1833), .Y(n4425));
  INVX1   g3347(.A(n4425), .Y(n4426));
  NOR2X1  g3348(.A(STATE2_REG_2__SCAN_IN), .B(n2071), .Y(n4427));
  OAI21X1 g3349(.A0(n4427), .A1(n4418), .B0(PHYADDRPOINTER_REG_0__SCAN_IN), .Y(n4428));
  OAI21X1 g3350(.A0(n4426), .A1(n4424), .B0(n4428), .Y(n4429));
  AOI21X1 g3351(.A0(n4423), .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B0(n4429), .Y(n4430));
  OAI21X1 g3352(.A0(n4422), .A1(n1843), .B0(n4430), .Y(n4431));
  XOR2X1  g3353(.A(n4431), .B(n4418), .Y(n4432));
  XOR2X1  g3354(.A(n4432), .B(n4421), .Y(n4433));
  XOR2X1  g3355(.A(n4433), .B(n4419), .Y(n4434));
  NAND4X1 g3356(.A(n1592), .B(n1423), .C(n1910), .D(n1720), .Y(n4435));
  NOR4X1  g3357(.A(n2054), .B(n1804), .C(n1833), .D(n4435), .Y(n4436));
  INVX1   g3358(.A(n4436), .Y(n4437));
  OAI21X1 g3359(.A0(n3219), .A1(n2075), .B0(n1217), .Y(n4438));
  NAND2X1 g3360(.A(n4438), .B(n4437), .Y(n4439));
  INVX1   g3361(.A(n4439), .Y(n4440));
  NOR3X1  g3362(.A(n4440), .B(n1910), .C(n2071), .Y(n4441));
  AOI22X1 g3363(.A0(STATE2_REG_1__SCAN_IN), .A1(n2071), .B0(STATE2_REG_2__SCAN_IN), .B1(n1217), .Y(n4446));
  AOI21X1 g3364(.A0(n4438), .A1(n4437), .B0(n4446), .Y(n4447));
  OAI21X1 g3365(.A0(n4447), .A1(n4440), .B0(PHYADDRPOINTER_REG_0__SCAN_IN), .Y(n4448));
  OAI21X1 g3366(.A0(n5914), .A1(n3252), .B0(n4448), .Y(n4449));
  AOI21X1 g3367(.A0(n4436), .A1(n3227), .B0(n4449), .Y(n4450));
  OAI21X1 g3368(.A0(n2120), .A1(n4434), .B0(n4450), .Y(U2986));
  INVX1   g3369(.A(EAX_REG_1__SCAN_IN), .Y(n4453));
  INVX1   g3370(.A(PHYADDRPOINTER_REG_1__SCAN_IN), .Y(n4454));
  NOR3X1  g3371(.A(n4454), .B(STATE2_REG_2__SCAN_IN), .C(n2071), .Y(n4455));
  AOI21X1 g3372(.A0(n4418), .A1(n4454), .B0(n4455), .Y(n4456));
  OAI21X1 g3373(.A0(n4426), .A1(n4453), .B0(n4456), .Y(n4457));
  AOI21X1 g3374(.A0(n4423), .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B0(n4457), .Y(n4458));
  OAI21X1 g3375(.A0(n4422), .A1(n1937), .B0(n4458), .Y(n4459));
  XOR2X1  g3376(.A(n4459), .B(n4419), .Y(n4460));
  NOR3X1  g3377(.A(n4460), .B(n4422), .C(n2218), .Y(n4461));
  INVX1   g3378(.A(n4422), .Y(n4462));
  INVX1   g3379(.A(n4460), .Y(n4463));
  AOI21X1 g3380(.A0(n4462), .A1(n2354), .B0(n4463), .Y(n4464));
  NOR2X1  g3381(.A(n4464), .B(n4461), .Y(n4465));
  NAND2X1 g3382(.A(n4432), .B(n4421), .Y(n4466));
  NOR2X1  g3383(.A(n4432), .B(n4421), .Y(n4467));
  OAI21X1 g3384(.A0(n4467), .A1(n4419), .B0(n4466), .Y(n4468));
  INVX1   g3385(.A(n4468), .Y(n4469));
  XOR2X1  g3386(.A(n4469), .B(n4465), .Y(n4470));
  NOR4X1  g3387(.A(n4440), .B(n1910), .C(n2071), .D(n4470), .Y(n4471));
  NOR4X1  g3388(.A(n1109), .B(STATE2_REG_1__SCAN_IN), .C(STATE2_REG_2__SCAN_IN), .D(n4440), .Y(n4472));
  NAND2X1 g3389(.A(n4447), .B(n4454), .Y(n4473));
  OAI21X1 g3390(.A0(n4439), .A1(n4454), .B0(n4473), .Y(n4474));
  NOR3X1  g3391(.A(n4474), .B(n4472), .C(n4471), .Y(n4475));
  OAI21X1 g3392(.A0(n4437), .A1(n3298), .B0(n4475), .Y(U2985));
  INVX1   g3393(.A(n4464), .Y(n4477));
  AOI21X1 g3394(.A0(n4468), .A1(n4477), .B0(n4461), .Y(n4478));
  INVX1   g3395(.A(n4427), .Y(n4479));
  OAI21X1 g3396(.A0(n4422), .A1(n2244), .B0(n4479), .Y(n4480));
  INVX1   g3397(.A(EAX_REG_2__SCAN_IN), .Y(n4481));
  XOR2X1  g3398(.A(PHYADDRPOINTER_REG_2__SCAN_IN), .B(n4454), .Y(n4482));
  INVX1   g3399(.A(n4482), .Y(n4483));
  AOI22X1 g3400(.A0(n4427), .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .B0(n4418), .B1(n4483), .Y(n4484));
  OAI21X1 g3401(.A0(n4426), .A1(n4481), .B0(n4484), .Y(n4485));
  AOI21X1 g3402(.A0(n4423), .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B0(n4485), .Y(n4486));
  OAI21X1 g3403(.A0(n4422), .A1(n1958), .B0(n4486), .Y(n4487));
  XOR2X1  g3404(.A(n4487), .B(n4419), .Y(n4488));
  INVX1   g3405(.A(n4488), .Y(n4489));
  NOR2X1  g3406(.A(n4489), .B(n4480), .Y(n4490));
  NOR2X1  g3407(.A(n4490), .B(n4478), .Y(n4491));
  AOI21X1 g3408(.A0(n4462), .A1(n2468), .B0(n4427), .Y(n4492));
  NOR2X1  g3409(.A(n4488), .B(n4492), .Y(n4493));
  INVX1   g3410(.A(n4493), .Y(n4494));
  XOR2X1  g3411(.A(n4488), .B(n4480), .Y(n4495));
  AOI22X1 g3412(.A0(n4494), .A1(n4491), .B0(n4478), .B1(n4495), .Y(n4496));
  INVX1   g3413(.A(n4496), .Y(n4497));
  AOI22X1 g3414(.A0(n4447), .A1(n4483), .B0(n4440), .B1(PHYADDRPOINTER_REG_2__SCAN_IN), .Y(n4498));
  OAI21X1 g3415(.A0(n5914), .A1(n1106), .B0(n4498), .Y(n4499));
  AOI21X1 g3416(.A0(n4436), .A1(n3315), .B0(n4499), .Y(n4500));
  OAI21X1 g3417(.A0(n4497), .A1(n2120), .B0(n4500), .Y(U2984));
  NAND2X1 g3418(.A(n4436), .B(n3342), .Y(n4502));
  NOR2X1  g3419(.A(n4422), .B(n2268), .Y(n4503));
  NAND4X1 g3420(.A(n1671), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C(STATE2_REG_2__SCAN_IN), .D(n1615), .Y(n4504));
  NAND3X1 g3421(.A(n1700), .B(EAX_REG_3__SCAN_IN), .C(STATE2_REG_2__SCAN_IN), .Y(n4505));
  NAND2X1 g3422(.A(PHYADDRPOINTER_REG_2__SCAN_IN), .B(PHYADDRPOINTER_REG_1__SCAN_IN), .Y(n4506));
  XOR2X1  g3423(.A(n4506), .B(PHYADDRPOINTER_REG_3__SCAN_IN), .Y(n4507));
  INVX1   g3424(.A(n4507), .Y(n4508));
  AOI22X1 g3425(.A0(n4427), .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .B0(n4418), .B1(n4508), .Y(n4509));
  NAND3X1 g3426(.A(n4509), .B(n4505), .C(n4504), .Y(n4510));
  AOI21X1 g3427(.A0(n4462), .A1(n1988), .B0(n4510), .Y(n4511));
  XOR2X1  g3428(.A(n4511), .B(n4419), .Y(n4512));
  XOR2X1  g3429(.A(n4512), .B(n4503), .Y(n4513));
  OAI21X1 g3430(.A0(n4490), .A1(n4478), .B0(n4494), .Y(n4514));
  XOR2X1  g3431(.A(n4514), .B(n4513), .Y(n4515));
  NAND4X1 g3432(.A(n4439), .B(STATE2_REG_1__SCAN_IN), .C(STATEBS16_REG_SCAN_IN), .D(n4515), .Y(n4516));
  NAND4X1 g3433(.A(REIP_REG_3__SCAN_IN), .B(n1910), .C(n1833), .D(n4439), .Y(n4517));
  AOI22X1 g3434(.A0(n4447), .A1(n4508), .B0(n4440), .B1(PHYADDRPOINTER_REG_3__SCAN_IN), .Y(n4518));
  NAND4X1 g3435(.A(n4517), .B(n4516), .C(n4502), .D(n4518), .Y(U2983));
  NAND2X1 g3436(.A(n4436), .B(n3399), .Y(n4520));
  NAND2X1 g3437(.A(n4462), .B(n3387), .Y(n4521));
  INVX1   g3438(.A(EAX_REG_4__SCAN_IN), .Y(n4522));
  INVX1   g3439(.A(PHYADDRPOINTER_REG_4__SCAN_IN), .Y(n4523));
  NAND3X1 g3440(.A(PHYADDRPOINTER_REG_3__SCAN_IN), .B(PHYADDRPOINTER_REG_2__SCAN_IN), .C(PHYADDRPOINTER_REG_1__SCAN_IN), .Y(n4524));
  XOR2X1  g3441(.A(n4524), .B(n4523), .Y(n4525));
  AOI22X1 g3442(.A0(n4427), .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .B0(n4418), .B1(n4525), .Y(n4526));
  OAI21X1 g3443(.A0(n4426), .A1(n4522), .B0(n4526), .Y(n4527));
  AOI21X1 g3444(.A0(n4423), .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B0(n4527), .Y(n4528));
  OAI21X1 g3445(.A0(n4422), .A1(n2008), .B0(n4528), .Y(n4529));
  XOR2X1  g3446(.A(n4529), .B(n4419), .Y(n4530));
  XOR2X1  g3447(.A(n4530), .B(n4521), .Y(n4531));
  NAND3X1 g3448(.A(n4512), .B(n4462), .C(n2688), .Y(n4532));
  AOI21X1 g3449(.A0(n4432), .A1(n4421), .B0(n4418), .Y(n4533));
  NOR3X1  g3450(.A(n4533), .B(n4464), .C(n4467), .Y(n4534));
  NOR3X1  g3451(.A(n4534), .B(n4493), .C(n4461), .Y(n4535));
  OAI22X1 g3452(.A0(n4503), .A1(n4512), .B0(n4489), .B1(n4480), .Y(n4536));
  OAI21X1 g3453(.A0(n4536), .A1(n4535), .B0(n4532), .Y(n4537));
  INVX1   g3454(.A(n4537), .Y(n4538));
  XOR2X1  g3455(.A(n4538), .B(n4531), .Y(n4539));
  INVX1   g3456(.A(n4539), .Y(n4540));
  NAND2X1 g3457(.A(n4540), .B(n4441), .Y(n4541));
  NAND4X1 g3458(.A(REIP_REG_4__SCAN_IN), .B(n1910), .C(n1833), .D(n4439), .Y(n4542));
  AOI22X1 g3459(.A0(n4447), .A1(n4525), .B0(n4440), .B1(PHYADDRPOINTER_REG_4__SCAN_IN), .Y(n4543));
  NAND4X1 g3460(.A(n4542), .B(n4541), .C(n4520), .D(n4543), .Y(U2982));
  NAND2X1 g3461(.A(n4436), .B(n3456), .Y(n4545));
  NAND3X1 g3462(.A(n2006), .B(n2005), .C(n1947), .Y(n4546));
  INVX1   g3463(.A(PHYADDRPOINTER_REG_5__SCAN_IN), .Y(n4547));
  NAND4X1 g3464(.A(PHYADDRPOINTER_REG_3__SCAN_IN), .B(PHYADDRPOINTER_REG_2__SCAN_IN), .C(PHYADDRPOINTER_REG_1__SCAN_IN), .D(PHYADDRPOINTER_REG_4__SCAN_IN), .Y(n4548));
  XOR2X1  g3465(.A(n4548), .B(PHYADDRPOINTER_REG_5__SCAN_IN), .Y(n4549));
  OAI22X1 g3466(.A0(n4479), .A1(n4547), .B0(n4419), .B1(n4549), .Y(n4550));
  AOI21X1 g3467(.A0(n4425), .A1(EAX_REG_5__SCAN_IN), .B0(n4550), .Y(n4551));
  OAI21X1 g3468(.A0(n4546), .A1(n4422), .B0(n4551), .Y(n4552));
  XOR2X1  g3469(.A(n4552), .B(n4419), .Y(n4553));
  NOR3X1  g3470(.A(n4553), .B(n4422), .C(n3515), .Y(n4554));
  INVX1   g3471(.A(n4553), .Y(n4555));
  AOI21X1 g3472(.A0(n4462), .A1(n3449), .B0(n4555), .Y(n4556));
  NOR2X1  g3473(.A(n4556), .B(n4554), .Y(n4557));
  XOR2X1  g3474(.A(n3834), .B(n3381), .Y(n4558));
  NOR3X1  g3475(.A(n4530), .B(n4422), .C(n4558), .Y(n4559));
  OAI21X1 g3476(.A0(n4422), .A1(n4558), .B0(n4530), .Y(n4560));
  AOI21X1 g3477(.A0(n4537), .A1(n4560), .B0(n4559), .Y(n4561));
  XOR2X1  g3478(.A(n4561), .B(n4557), .Y(n4562));
  INVX1   g3479(.A(n4562), .Y(n4563));
  NAND2X1 g3480(.A(n4563), .B(n4441), .Y(n4564));
  NAND4X1 g3481(.A(REIP_REG_5__SCAN_IN), .B(n1910), .C(n1833), .D(n4439), .Y(n4565));
  INVX1   g3482(.A(n4549), .Y(n4566));
  AOI22X1 g3483(.A0(n4447), .A1(n4566), .B0(n4440), .B1(PHYADDRPOINTER_REG_5__SCAN_IN), .Y(n4567));
  NAND4X1 g3484(.A(n4565), .B(n4564), .C(n4545), .D(n4567), .Y(U2981));
  NAND2X1 g3485(.A(n4436), .B(n3520), .Y(n4569));
  INVX1   g3486(.A(PHYADDRPOINTER_REG_6__SCAN_IN), .Y(n4570));
  NOR2X1  g3487(.A(n4548), .B(n4547), .Y(n4571));
  XOR2X1  g3488(.A(n4571), .B(n4570), .Y(n4572));
  OAI22X1 g3489(.A0(n4479), .A1(n4570), .B0(n4419), .B1(n4572), .Y(n4573));
  AOI21X1 g3490(.A0(n4425), .A1(EAX_REG_6__SCAN_IN), .B0(n4573), .Y(n4574));
  XOR2X1  g3491(.A(n4574), .B(n4418), .Y(n4575));
  NOR2X1  g3492(.A(n4422), .B(n3637), .Y(n4576));
  XOR2X1  g3493(.A(n4576), .B(n4575), .Y(n4577));
  INVX1   g3494(.A(n4554), .Y(n4578));
  OAI21X1 g3495(.A0(n4561), .A1(n4556), .B0(n4578), .Y(n4579));
  NAND2X1 g3496(.A(n4577), .B(n4579), .Y(n4581));
  OAI21X1 g3497(.A0(n4579), .A1(n4577), .B0(n4581), .Y(n4582));
  NAND2X1 g3498(.A(n4582), .B(n4441), .Y(n4583));
  NAND4X1 g3499(.A(REIP_REG_6__SCAN_IN), .B(n1910), .C(n1833), .D(n4439), .Y(n4584));
  INVX1   g3500(.A(n4572), .Y(n4585));
  AOI22X1 g3501(.A0(n4447), .A1(n4585), .B0(n4440), .B1(PHYADDRPOINTER_REG_6__SCAN_IN), .Y(n4586));
  NAND4X1 g3502(.A(n4584), .B(n4583), .C(n4569), .D(n4586), .Y(U2980));
  INVX1   g3503(.A(n4575), .Y(n4588));
  OAI21X1 g3504(.A0(n4576), .A1(n4588), .B0(n4579), .Y(n4589));
  NOR3X1  g3505(.A(n4575), .B(n4422), .C(n3637), .Y(n4590));
  NAND4X1 g3506(.A(n3562), .B(n3643), .C(n3641), .D(n4462), .Y(n4591));
  INVX1   g3507(.A(PHYADDRPOINTER_REG_7__SCAN_IN), .Y(n4592));
  NOR3X1  g3508(.A(n4548), .B(n4570), .C(n4547), .Y(n4593));
  XOR2X1  g3509(.A(n4593), .B(n4592), .Y(n4594));
  OAI22X1 g3510(.A0(n4479), .A1(n4592), .B0(n4419), .B1(n4594), .Y(n4595));
  AOI21X1 g3511(.A0(n4425), .A1(EAX_REG_7__SCAN_IN), .B0(n4595), .Y(n4596));
  XOR2X1  g3512(.A(n4596), .B(n4418), .Y(n4597));
  XOR2X1  g3513(.A(n4597), .B(n4591), .Y(n4598));
  NOR2X1  g3514(.A(n4598), .B(n4590), .Y(n4599));
  NAND2X1 g3515(.A(n4599), .B(n4589), .Y(n4600));
  NOR2X1  g3516(.A(n4597), .B(n4591), .Y(n4601));
  NAND2X1 g3517(.A(n4597), .B(n4591), .Y(n4602));
  OAI21X1 g3518(.A0(n4576), .A1(n4588), .B0(n4602), .Y(n4603));
  NOR2X1  g3519(.A(n4603), .B(n4601), .Y(n4604));
  OAI21X1 g3520(.A0(n4590), .A1(n4579), .B0(n4604), .Y(n4605));
  NAND2X1 g3521(.A(n4605), .B(n4600), .Y(n4606));
  NOR2X1  g3522(.A(n4606), .B(n2120), .Y(n4607));
  INVX1   g3523(.A(n4594), .Y(n4608));
  AOI22X1 g3524(.A0(n4447), .A1(n4608), .B0(n4440), .B1(PHYADDRPOINTER_REG_7__SCAN_IN), .Y(n4609));
  OAI21X1 g3525(.A0(n5914), .A1(n1091), .B0(n4609), .Y(n4610));
  NOR2X1  g3526(.A(n4610), .B(n4607), .Y(n4611));
  OAI21X1 g3527(.A0(n4437), .A1(n3570), .B0(n4611), .Y(U2979));
  INVX1   g3528(.A(PHYADDRPOINTER_REG_8__SCAN_IN), .Y(n4613));
  NOR4X1  g3529(.A(n4592), .B(n4570), .C(n4547), .D(n4548), .Y(n4614));
  XOR2X1  g3530(.A(n4614), .B(n4613), .Y(n4615));
  OAI22X1 g3531(.A0(n4479), .A1(n4613), .B0(n4419), .B1(n4615), .Y(n4616));
  AOI21X1 g3532(.A0(n4425), .A1(EAX_REG_8__SCAN_IN), .B0(n4616), .Y(n4617));
  XOR2X1  g3533(.A(n4617), .B(n4418), .Y(n4618));
  NOR3X1  g3534(.A(n4618), .B(n4422), .C(n3837), .Y(n4619));
  INVX1   g3535(.A(n4618), .Y(n4620));
  AOI21X1 g3536(.A0(n4462), .A1(n3628), .B0(n4620), .Y(n4621));
  NOR2X1  g3537(.A(n4621), .B(n4619), .Y(n4622));
  NAND2X1 g3538(.A(n4462), .B(n3512), .Y(n4623));
  AOI22X1 g3539(.A0(n4591), .A1(n4597), .B0(n4623), .B1(n4575), .Y(n4624));
  NOR2X1  g3540(.A(n4554), .B(n4559), .Y(n4625));
  NOR2X1  g3541(.A(n4625), .B(n4556), .Y(n4626));
  NAND2X1 g3542(.A(n4626), .B(n4624), .Y(n4627));
  OAI21X1 g3543(.A0(n4422), .A1(n3515), .B0(n4553), .Y(n4628));
  NAND4X1 g3544(.A(n4628), .B(n4537), .C(n4560), .D(n4624), .Y(n4629));
  AOI21X1 g3545(.A0(n4602), .A1(n4590), .B0(n4601), .Y(n4630));
  NAND3X1 g3546(.A(n4630), .B(n4629), .C(n4627), .Y(n4631));
  XOR2X1  g3547(.A(n4631), .B(n4622), .Y(n4632));
  INVX1   g3548(.A(n4615), .Y(n4633));
  AOI22X1 g3549(.A0(n4447), .A1(n4633), .B0(n4440), .B1(PHYADDRPOINTER_REG_8__SCAN_IN), .Y(n4634));
  OAI21X1 g3550(.A0(n5914), .A1(n1088), .B0(n4634), .Y(n4635));
  AOI21X1 g3551(.A0(n4632), .A1(n4441), .B0(n4635), .Y(n4636));
  OAI21X1 g3552(.A0(n4437), .A1(n3656), .B0(n4636), .Y(U2978));
  NAND3X1 g3553(.A(n4620), .B(n4462), .C(n3628), .Y(n4638));
  NOR3X1  g3554(.A(n4625), .B(n4603), .C(n4556), .Y(n4639));
  NAND3X1 g3555(.A(n4628), .B(n4537), .C(n4560), .Y(n4640));
  OAI21X1 g3556(.A0(n4640), .A1(n4603), .B0(n4630), .Y(n4641));
  NOR2X1  g3557(.A(n4641), .B(n4639), .Y(n4642));
  OAI21X1 g3558(.A0(n4642), .A1(n4621), .B0(n4638), .Y(n4643));
  INVX1   g3559(.A(PHYADDRPOINTER_REG_9__SCAN_IN), .Y(n4644));
  INVX1   g3560(.A(n4614), .Y(n4645));
  NOR2X1  g3561(.A(n4645), .B(n4613), .Y(n4646));
  XOR2X1  g3562(.A(n4646), .B(n4644), .Y(n4647));
  OAI22X1 g3563(.A0(n4479), .A1(n4644), .B0(n4419), .B1(n4647), .Y(n4648));
  AOI21X1 g3564(.A0(n4425), .A1(EAX_REG_9__SCAN_IN), .B0(n4648), .Y(n4649));
  XOR2X1  g3565(.A(n4649), .B(n4418), .Y(n4650));
  NOR2X1  g3566(.A(n4422), .B(n3690), .Y(n4651));
  XOR2X1  g3567(.A(n4651), .B(n4650), .Y(n4652));
  XOR2X1  g3568(.A(n4652), .B(n4643), .Y(n4653));
  NOR2X1  g3569(.A(n4653), .B(n2120), .Y(n4654));
  INVX1   g3570(.A(n4647), .Y(n4655));
  AOI22X1 g3571(.A0(n4447), .A1(n4655), .B0(n4440), .B1(PHYADDRPOINTER_REG_9__SCAN_IN), .Y(n4656));
  OAI21X1 g3572(.A0(n5914), .A1(n1085), .B0(n4656), .Y(n4657));
  NOR2X1  g3573(.A(n4657), .B(n4654), .Y(n4658));
  OAI21X1 g3574(.A0(n4437), .A1(n3704), .B0(n4658), .Y(U2977));
  OAI21X1 g3575(.A0(n4422), .A1(n3690), .B0(n4650), .Y(n4660));
  NOR3X1  g3576(.A(n4650), .B(n4422), .C(n3690), .Y(n4661));
  AOI21X1 g3577(.A0(n4660), .A1(n4619), .B0(n4661), .Y(n4662));
  INVX1   g3578(.A(n4650), .Y(n4663));
  AOI21X1 g3579(.A0(n4462), .A1(n3687), .B0(n4663), .Y(n4664));
  NOR2X1  g3580(.A(n4664), .B(n4621), .Y(n4665));
  OAI21X1 g3581(.A0(n4641), .A1(n4639), .B0(n4665), .Y(n4666));
  NAND2X1 g3582(.A(n4666), .B(n4662), .Y(n4667));
  INVX1   g3583(.A(PHYADDRPOINTER_REG_10__SCAN_IN), .Y(n4668));
  NOR3X1  g3584(.A(n4645), .B(n4644), .C(n4613), .Y(n4669));
  XOR2X1  g3585(.A(n4669), .B(n4668), .Y(n4670));
  OAI22X1 g3586(.A0(n4479), .A1(n4668), .B0(n4419), .B1(n4670), .Y(n4671));
  AOI21X1 g3587(.A0(n4425), .A1(EAX_REG_10__SCAN_IN), .B0(n4671), .Y(n4672));
  XOR2X1  g3588(.A(n4672), .B(n4418), .Y(n4673));
  OAI21X1 g3589(.A0(n4422), .A1(n3824), .B0(n4673), .Y(n4674));
  NAND2X1 g3590(.A(n4674), .B(n4667), .Y(n4675));
  NOR3X1  g3591(.A(n4673), .B(n4422), .C(n3824), .Y(n4676));
  INVX1   g3592(.A(n4673), .Y(n4677));
  AOI21X1 g3593(.A0(n4462), .A1(n3738), .B0(n4677), .Y(n4678));
  NOR2X1  g3594(.A(n4676), .B(n4678), .Y(n4679));
  OAI22X1 g3595(.A0(n4676), .A1(n4675), .B0(n4667), .B1(n4679), .Y(n4680));
  NOR2X1  g3596(.A(n4680), .B(n2120), .Y(n4681));
  INVX1   g3597(.A(n4670), .Y(n4682));
  AOI22X1 g3598(.A0(n4447), .A1(n4682), .B0(n4440), .B1(PHYADDRPOINTER_REG_10__SCAN_IN), .Y(n4683));
  OAI21X1 g3599(.A0(n5914), .A1(n1082), .B0(n4683), .Y(n4684));
  NOR2X1  g3600(.A(n4684), .B(n4681), .Y(n4685));
  OAI21X1 g3601(.A0(n4437), .A1(n3743), .B0(n4685), .Y(U2976));
  NAND4X1 g3602(.A(PHYADDRPOINTER_REG_10__SCAN_IN), .B(PHYADDRPOINTER_REG_9__SCAN_IN), .C(PHYADDRPOINTER_REG_8__SCAN_IN), .D(n4614), .Y(n4687));
  XOR2X1  g3603(.A(n4687), .B(PHYADDRPOINTER_REG_11__SCAN_IN), .Y(n4688));
  NAND3X1 g3604(.A(PHYADDRPOINTER_REG_11__SCAN_IN), .B(n1833), .C(STATEBS16_REG_SCAN_IN), .Y(n4689));
  OAI21X1 g3605(.A0(n4688), .A1(n4419), .B0(n4689), .Y(n4690));
  AOI21X1 g3606(.A0(n4425), .A1(EAX_REG_11__SCAN_IN), .B0(n4690), .Y(n4691));
  XOR2X1  g3607(.A(n4691), .B(n4418), .Y(n4692));
  INVX1   g3608(.A(n4692), .Y(n4693));
  AOI21X1 g3609(.A0(n4462), .A1(n3779), .B0(n4693), .Y(n4694));
  NOR3X1  g3610(.A(n4692), .B(n4422), .C(n3776), .Y(n4695));
  NOR2X1  g3611(.A(n4695), .B(n4694), .Y(n4696));
  OAI21X1 g3612(.A0(n4422), .A1(n3776), .B0(n4692), .Y(n4697));
  NAND3X1 g3613(.A(n4693), .B(n4462), .C(n3779), .Y(n4698));
  AOI21X1 g3614(.A0(n4698), .A1(n4697), .B0(n4676), .Y(n4699));
  NAND3X1 g3615(.A(n4677), .B(n4462), .C(n3738), .Y(n4700));
  NAND2X1 g3616(.A(n4700), .B(n4675), .Y(n4701));
  AOI22X1 g3617(.A0(n4699), .A1(n4675), .B0(n4696), .B1(n4701), .Y(n4702));
  INVX1   g3618(.A(n4688), .Y(n4703));
  AOI22X1 g3619(.A0(n4447), .A1(n4703), .B0(n4440), .B1(PHYADDRPOINTER_REG_11__SCAN_IN), .Y(n4704));
  OAI21X1 g3620(.A0(n5914), .A1(n1079), .B0(n4704), .Y(n4705));
  AOI21X1 g3621(.A0(n4702), .A1(n4441), .B0(n4705), .Y(n4706));
  OAI21X1 g3622(.A0(n4437), .A1(n3785), .B0(n4706), .Y(U2975));
  XOR2X1  g3623(.A(n3817), .B(n3813), .Y(n4708));
  INVX1   g3624(.A(PHYADDRPOINTER_REG_12__SCAN_IN), .Y(n4709));
  NAND3X1 g3625(.A(n4669), .B(PHYADDRPOINTER_REG_11__SCAN_IN), .C(PHYADDRPOINTER_REG_10__SCAN_IN), .Y(n4710));
  XOR2X1  g3626(.A(n4710), .B(PHYADDRPOINTER_REG_12__SCAN_IN), .Y(n4711));
  OAI22X1 g3627(.A0(n4479), .A1(n4709), .B0(n4419), .B1(n4711), .Y(n4712));
  AOI21X1 g3628(.A0(n4425), .A1(EAX_REG_12__SCAN_IN), .B0(n4712), .Y(n4713));
  XOR2X1  g3629(.A(n4713), .B(n4418), .Y(n4714));
  OAI21X1 g3630(.A0(n4422), .A1(n4708), .B0(n4714), .Y(n4715));
  INVX1   g3631(.A(n4715), .Y(n4716));
  NOR3X1  g3632(.A(n4714), .B(n4422), .C(n4708), .Y(n4717));
  NOR2X1  g3633(.A(n4717), .B(n4716), .Y(n4718));
  NOR4X1  g3634(.A(n4678), .B(n4664), .C(n4621), .D(n4694), .Y(n4719));
  NAND2X1 g3635(.A(n4697), .B(n4674), .Y(n4720));
  OAI21X1 g3636(.A0(n4695), .A1(n4676), .B0(n4697), .Y(n4721));
  OAI21X1 g3637(.A0(n4720), .A1(n4662), .B0(n4721), .Y(n4722));
  AOI21X1 g3638(.A0(n4719), .A1(n4631), .B0(n4722), .Y(n4723));
  XOR2X1  g3639(.A(n4723), .B(n4718), .Y(n4724));
  NOR2X1  g3640(.A(n4724), .B(n2120), .Y(n4725));
  INVX1   g3641(.A(n4711), .Y(n4726));
  AOI22X1 g3642(.A0(n4447), .A1(n4726), .B0(n4440), .B1(PHYADDRPOINTER_REG_12__SCAN_IN), .Y(n4727));
  OAI21X1 g3643(.A0(n5914), .A1(n1076), .B0(n4727), .Y(n4728));
  NOR2X1  g3644(.A(n4728), .B(n4725), .Y(n4729));
  OAI21X1 g3645(.A0(n4437), .A1(n3843), .B0(n4729), .Y(U2974));
  OAI21X1 g3646(.A0(n4641), .A1(n4639), .B0(n4719), .Y(n4731));
  NAND3X1 g3647(.A(n4663), .B(n4462), .C(n3687), .Y(n4732));
  OAI21X1 g3648(.A0(n4664), .A1(n4638), .B0(n4732), .Y(n4733));
  NOR2X1  g3649(.A(n4694), .B(n4678), .Y(n4734));
  AOI21X1 g3650(.A0(n4698), .A1(n4700), .B0(n4694), .Y(n4735));
  AOI21X1 g3651(.A0(n4734), .A1(n4733), .B0(n4735), .Y(n4736));
  AOI21X1 g3652(.A0(n4736), .A1(n4731), .B0(n4716), .Y(n4737));
  NOR2X1  g3653(.A(n4737), .B(n4717), .Y(n4738));
  INVX1   g3654(.A(PHYADDRPOINTER_REG_13__SCAN_IN), .Y(n4739));
  NAND4X1 g3655(.A(PHYADDRPOINTER_REG_12__SCAN_IN), .B(PHYADDRPOINTER_REG_11__SCAN_IN), .C(PHYADDRPOINTER_REG_10__SCAN_IN), .D(n4669), .Y(n4740));
  XOR2X1  g3656(.A(n4740), .B(n4739), .Y(n4741));
  INVX1   g3657(.A(EAX_REG_13__SCAN_IN), .Y(n4742));
  OAI22X1 g3658(.A0(n4426), .A1(n4742), .B0(n4739), .B1(n4479), .Y(n4743));
  AOI21X1 g3659(.A0(n4741), .A1(n4418), .B0(n4743), .Y(n4744));
  XOR2X1  g3660(.A(n4744), .B(n4418), .Y(n4745));
  INVX1   g3661(.A(n4745), .Y(n4746));
  NOR2X1  g3662(.A(n4422), .B(n3875), .Y(n4747));
  XOR2X1  g3663(.A(n4747), .B(n4746), .Y(n4748));
  OAI21X1 g3664(.A0(n4422), .A1(n3875), .B0(n4745), .Y(n4749));
  NOR3X1  g3665(.A(n4745), .B(n4422), .C(n3875), .Y(n4750));
  INVX1   g3666(.A(n4750), .Y(n4751));
  AOI21X1 g3667(.A0(n4751), .A1(n4749), .B0(n4738), .Y(n4752));
  AOI21X1 g3668(.A0(n4748), .A1(n4738), .B0(n4752), .Y(n4753));
  NOR2X1  g3669(.A(n4753), .B(n2120), .Y(n4754));
  AOI22X1 g3670(.A0(n4447), .A1(n4741), .B0(n4440), .B1(PHYADDRPOINTER_REG_13__SCAN_IN), .Y(n4755));
  OAI21X1 g3671(.A0(n5914), .A1(n1073), .B0(n4755), .Y(n4756));
  NOR2X1  g3672(.A(n4756), .B(n4754), .Y(n4757));
  OAI21X1 g3673(.A0(n4437), .A1(n3889), .B0(n4757), .Y(U2973));
  INVX1   g3674(.A(n4714), .Y(n4759));
  NAND3X1 g3675(.A(n4759), .B(n4462), .C(n3818), .Y(n4760));
  OAI21X1 g3676(.A0(n4723), .A1(n4716), .B0(n4760), .Y(n4761));
  AOI21X1 g3677(.A0(n4749), .A1(n4761), .B0(n4750), .Y(n4762));
  NOR3X1  g3678(.A(n4710), .B(n4739), .C(n4709), .Y(n4763));
  XOR2X1  g3679(.A(n4763), .B(PHYADDRPOINTER_REG_14__SCAN_IN), .Y(n4764));
  INVX1   g3680(.A(PHYADDRPOINTER_REG_14__SCAN_IN), .Y(n4765));
  INVX1   g3681(.A(EAX_REG_14__SCAN_IN), .Y(n4766));
  OAI22X1 g3682(.A0(n4426), .A1(n4766), .B0(n4765), .B1(n4479), .Y(n4767));
  AOI21X1 g3683(.A0(n4764), .A1(n4418), .B0(n4767), .Y(n4768));
  XOR2X1  g3684(.A(n4768), .B(n4418), .Y(n4769));
  INVX1   g3685(.A(n4769), .Y(n4770));
  NOR2X1  g3686(.A(n4422), .B(n3921), .Y(n4771));
  XOR2X1  g3687(.A(n4771), .B(n4770), .Y(n4772));
  NAND2X1 g3688(.A(n4762), .B(n4772), .Y(n4773));
  NOR3X1  g3689(.A(n4769), .B(n4422), .C(n3921), .Y(n4774));
  AOI21X1 g3690(.A0(n4462), .A1(n3967), .B0(n4770), .Y(n4775));
  OAI21X1 g3691(.A0(n4772), .A1(n4762), .B0(n4773), .Y(n4777));
  AOI22X1 g3692(.A0(n4447), .A1(n4764), .B0(n4440), .B1(PHYADDRPOINTER_REG_14__SCAN_IN), .Y(n4778));
  OAI21X1 g3693(.A0(n5914), .A1(n1070), .B0(n4778), .Y(n4779));
  AOI21X1 g3694(.A0(n4777), .A1(n4441), .B0(n4779), .Y(n4780));
  OAI21X1 g3695(.A0(n4437), .A1(n3926), .B0(n4780), .Y(U2972));
  AOI21X1 g3696(.A0(n4462), .A1(n3878), .B0(n4746), .Y(n4782));
  OAI21X1 g3697(.A0(n4782), .A1(n4738), .B0(n4751), .Y(n4783));
  OAI21X1 g3698(.A0(n4422), .A1(n3921), .B0(n4769), .Y(n4784));
  NAND2X1 g3699(.A(n4784), .B(n4783), .Y(n4785));
  NOR4X1  g3700(.A(n4765), .B(n4739), .C(n4709), .D(n4710), .Y(n4786));
  XOR2X1  g3701(.A(n4786), .B(PHYADDRPOINTER_REG_15__SCAN_IN), .Y(n4787));
  INVX1   g3702(.A(EAX_REG_15__SCAN_IN), .Y(n4788));
  NAND3X1 g3703(.A(PHYADDRPOINTER_REG_15__SCAN_IN), .B(n1833), .C(STATEBS16_REG_SCAN_IN), .Y(n4789));
  OAI21X1 g3704(.A0(n4426), .A1(n4788), .B0(n4789), .Y(n4790));
  AOI21X1 g3705(.A0(n4787), .A1(n4418), .B0(n4790), .Y(n4791));
  XOR2X1  g3706(.A(n4791), .B(n4418), .Y(n4792));
  NOR3X1  g3707(.A(n4792), .B(n4422), .C(n3960), .Y(n4793));
  INVX1   g3708(.A(n4792), .Y(n4794));
  AOI21X1 g3709(.A0(n4462), .A1(n3963), .B0(n4794), .Y(n4795));
  NOR2X1  g3710(.A(n4795), .B(n4793), .Y(n4796));
  NOR2X1  g3711(.A(n4796), .B(n4774), .Y(n4797));
  NAND3X1 g3712(.A(n4770), .B(n4462), .C(n3967), .Y(n4798));
  NAND2X1 g3713(.A(n4798), .B(n4762), .Y(n4799));
  NOR3X1  g3714(.A(n4795), .B(n4793), .C(n4775), .Y(n4800));
  AOI22X1 g3715(.A0(n4799), .A1(n4800), .B0(n4797), .B1(n4785), .Y(n4801));
  AOI22X1 g3716(.A0(n4447), .A1(n4787), .B0(n4440), .B1(PHYADDRPOINTER_REG_15__SCAN_IN), .Y(n4802));
  OAI21X1 g3717(.A0(n5914), .A1(n1067), .B0(n4802), .Y(n4803));
  AOI21X1 g3718(.A0(n4801), .A1(n4441), .B0(n4803), .Y(n4804));
  OAI21X1 g3719(.A0(n4437), .A1(n3971), .B0(n4804), .Y(U2971));
  OAI21X1 g3720(.A0(n4422), .A1(n3960), .B0(n4792), .Y(n4806));
  NAND4X1 g3721(.A(n4784), .B(n4749), .C(n4715), .D(n4806), .Y(n4807));
  AOI21X1 g3722(.A0(n4736), .A1(n4731), .B0(n4807), .Y(n4808));
  NAND4X1 g3723(.A(n4784), .B(n4749), .C(n4717), .D(n4806), .Y(n4809));
  NAND2X1 g3724(.A(n4462), .B(n3963), .Y(n4810));
  OAI21X1 g3725(.A0(n4792), .A1(n4810), .B0(n4798), .Y(n4811));
  NOR4X1  g3726(.A(n4745), .B(n4422), .C(n3875), .D(n4775), .Y(n4812));
  OAI21X1 g3727(.A0(n4812), .A1(n4811), .B0(n4806), .Y(n4813));
  NAND2X1 g3728(.A(n4813), .B(n4809), .Y(n4814));
  NOR2X1  g3729(.A(n4814), .B(n4808), .Y(n4815));
  NOR3X1  g3730(.A(n1677), .B(n1639), .C(n1872), .Y(n4816));
  AOI21X1 g3731(.A0(n1684), .A1(STATE2_REG_0__SCAN_IN), .B0(n4816), .Y(n4817));
  INVX1   g3732(.A(n4817), .Y(n4818));
  OAI22X1 g3733(.A0(n1251), .A1(n1242), .B0(n1444), .B1(n1352), .Y(n4823));
  OAI22X1 g3734(.A0(n1261), .A1(n1249), .B0(n1438), .B1(n1326), .Y(n4828));
  OAI22X1 g3735(.A0(n1284), .A1(n1441), .B0(n1425), .B1(n1343), .Y(n4833));
  OAI22X1 g3736(.A0(n1342), .A1(n1426), .B0(n1259), .B1(n1359), .Y(n4838));
  NOR4X1  g3737(.A(n4833), .B(n4828), .C(n4823), .D(n4838), .Y(n4839));
  OAI22X1 g3738(.A0(n1263), .A1(n1429), .B0(n1430), .B1(n1243), .Y(n4844));
  OAI22X1 g3739(.A0(n1347), .A1(n1258), .B0(n1440), .B1(n1358), .Y(n4849));
  OAI22X1 g3740(.A0(n1348), .A1(n1434), .B0(n1443), .B1(n1332), .Y(n4854));
  OAI22X1 g3741(.A0(n1354), .A1(n1437), .B0(n1435), .B1(n1334), .Y(n4859));
  NOR4X1  g3742(.A(n4854), .B(n4849), .C(n4844), .D(n4859), .Y(n4860));
  AOI21X1 g3743(.A0(n4860), .A1(n4839), .B0(n4422), .Y(n4861));
  NAND3X1 g3744(.A(n4763), .B(PHYADDRPOINTER_REG_15__SCAN_IN), .C(PHYADDRPOINTER_REG_14__SCAN_IN), .Y(n4862));
  XOR2X1  g3745(.A(n4862), .B(PHYADDRPOINTER_REG_16__SCAN_IN), .Y(n4863));
  AOI22X1 g3746(.A0(n4425), .A1(EAX_REG_16__SCAN_IN), .B0(PHYADDRPOINTER_REG_16__SCAN_IN), .B1(n4427), .Y(n4864));
  OAI21X1 g3747(.A0(n4863), .A1(n4419), .B0(n4864), .Y(n4865));
  AOI21X1 g3748(.A0(n4861), .A1(n4818), .B0(n4865), .Y(n4866));
  XOR2X1  g3749(.A(n4866), .B(n4418), .Y(n4867));
  INVX1   g3750(.A(n4867), .Y(n4868));
  AOI21X1 g3751(.A0(n4462), .A1(n4058), .B0(n4868), .Y(n4869));
  INVX1   g3752(.A(n4869), .Y(n4870));
  OAI21X1 g3753(.A0(n4814), .A1(n4808), .B0(n4870), .Y(n4871));
  NAND3X1 g3754(.A(n4868), .B(n4462), .C(n4058), .Y(n4872));
  NOR2X1  g3755(.A(n4964), .B(n4871), .Y(n4874));
  NAND2X1 g3756(.A(n4872), .B(n4870), .Y(n4875));
  AOI21X1 g3757(.A0(n4875), .A1(n4815), .B0(n4874), .Y(n4876));
  INVX1   g3758(.A(n4863), .Y(n4877));
  AOI22X1 g3759(.A0(n4447), .A1(n4877), .B0(n4440), .B1(PHYADDRPOINTER_REG_16__SCAN_IN), .Y(n4878));
  OAI21X1 g3760(.A0(n5914), .A1(n1064), .B0(n4878), .Y(n4879));
  AOI21X1 g3761(.A0(n4876), .A1(n4441), .B0(n4879), .Y(n4880));
  OAI21X1 g3762(.A0(n4437), .A1(n4007), .B0(n4880), .Y(U2970));
  NOR2X1  g3763(.A(n4422), .B(n4028), .Y(n4882));
  OAI22X1 g3764(.A0(n1251), .A1(n1450), .B0(n1357), .B1(n1352), .Y(n4883));
  OAI22X1 g3765(.A0(n1261), .A1(n1453), .B0(n1346), .B1(n1326), .Y(n4884));
  OAI22X1 g3766(.A0(n1284), .A1(n1351), .B0(n1324), .B1(n1343), .Y(n4885));
  OAI22X1 g3767(.A0(n1342), .A1(n1325), .B0(n1457), .B1(n1359), .Y(n4886));
  NOR4X1  g3768(.A(n4885), .B(n4884), .C(n4883), .D(n4886), .Y(n4887));
  OAI22X1 g3769(.A0(n1263), .A1(n1330), .B0(n1331), .B1(n1243), .Y(n4888));
  OAI22X1 g3770(.A0(n1347), .A1(n1456), .B0(n1350), .B1(n1358), .Y(n4889));
  OAI22X1 g3771(.A0(n1348), .A1(n1340), .B0(n1356), .B1(n1332), .Y(n4890));
  OAI22X1 g3772(.A0(n1354), .A1(n1345), .B0(n1341), .B1(n1334), .Y(n4891));
  NOR4X1  g3773(.A(n4890), .B(n4889), .C(n4888), .D(n4891), .Y(n4892));
  AOI21X1 g3774(.A0(n4892), .A1(n4887), .B0(n4422), .Y(n4893));
  INVX1   g3775(.A(PHYADDRPOINTER_REG_17__SCAN_IN), .Y(n4894));
  INVX1   g3776(.A(PHYADDRPOINTER_REG_16__SCAN_IN), .Y(n4895));
  NOR2X1  g3777(.A(n4862), .B(n4895), .Y(n4896));
  XOR2X1  g3778(.A(n4896), .B(n4894), .Y(n4897));
  AOI22X1 g3779(.A0(n4425), .A1(EAX_REG_17__SCAN_IN), .B0(PHYADDRPOINTER_REG_17__SCAN_IN), .B1(n4427), .Y(n4898));
  OAI21X1 g3780(.A0(n4897), .A1(n4419), .B0(n4898), .Y(n4899));
  AOI21X1 g3781(.A0(n4893), .A1(n4818), .B0(n4899), .Y(n4900));
  XOR2X1  g3782(.A(n4900), .B(n4418), .Y(n4901));
  INVX1   g3783(.A(n4901), .Y(n4902));
  XOR2X1  g3784(.A(n4902), .B(n4882), .Y(n4903));
  NAND2X1 g3785(.A(n4872), .B(n4871), .Y(n4904));
  XOR2X1  g3786(.A(n4904), .B(n4903), .Y(n4905));
  INVX1   g3787(.A(n4897), .Y(n4906));
  AOI22X1 g3788(.A0(n4447), .A1(n4906), .B0(n4440), .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .Y(n4907));
  OAI21X1 g3789(.A0(n5914), .A1(n1061), .B0(n4907), .Y(n4908));
  AOI21X1 g3790(.A0(n4905), .A1(n4441), .B0(n4908), .Y(n4909));
  OAI21X1 g3791(.A0(n4437), .A1(n4031), .B0(n4909), .Y(U2969));
  OAI22X1 g3792(.A0(n1251), .A1(n1706), .B0(n1636), .B1(n1352), .Y(n4911));
  OAI22X1 g3793(.A0(n1261), .A1(n1709), .B0(n1630), .B1(n1326), .Y(n4912));
  OAI22X1 g3794(.A0(n1284), .A1(n1633), .B0(n1617), .B1(n1343), .Y(n4913));
  OAI22X1 g3795(.A0(n1342), .A1(n1618), .B0(n1713), .B1(n1359), .Y(n4914));
  NOR4X1  g3796(.A(n4913), .B(n4912), .C(n4911), .D(n4914), .Y(n4915));
  OAI22X1 g3797(.A0(n1263), .A1(n1621), .B0(n1622), .B1(n1243), .Y(n4916));
  OAI22X1 g3798(.A0(n1347), .A1(n1712), .B0(n1632), .B1(n1358), .Y(n4917));
  OAI22X1 g3799(.A0(n1348), .A1(n1626), .B0(n1635), .B1(n1332), .Y(n4918));
  OAI22X1 g3800(.A0(n1354), .A1(n1629), .B0(n1627), .B1(n1334), .Y(n4919));
  NOR4X1  g3801(.A(n4918), .B(n4917), .C(n4916), .D(n4919), .Y(n4920));
  AOI21X1 g3802(.A0(n4920), .A1(n4915), .B0(n4422), .Y(n4921));
  INVX1   g3803(.A(PHYADDRPOINTER_REG_18__SCAN_IN), .Y(n4922));
  NOR3X1  g3804(.A(n4862), .B(n4894), .C(n4895), .Y(n4923));
  XOR2X1  g3805(.A(n4923), .B(n4922), .Y(n4924));
  AOI22X1 g3806(.A0(n4425), .A1(EAX_REG_18__SCAN_IN), .B0(PHYADDRPOINTER_REG_18__SCAN_IN), .B1(n4427), .Y(n4925));
  OAI21X1 g3807(.A0(n4924), .A1(n4419), .B0(n4925), .Y(n4926));
  AOI21X1 g3808(.A0(n4921), .A1(n4818), .B0(n4926), .Y(n4927));
  XOR2X1  g3809(.A(n4927), .B(n4418), .Y(n4928));
  INVX1   g3810(.A(n4928), .Y(n4929));
  XOR2X1  g3811(.A(n4929), .B(n4882), .Y(n4930));
  INVX1   g3812(.A(n4882), .Y(n4931));
  AOI22X1 g3813(.A0(n4931), .A1(n4901), .B0(n4872), .B1(n4871), .Y(n4932));
  AOI21X1 g3814(.A0(n4902), .A1(n4882), .B0(n4932), .Y(n4933));
  XOR2X1  g3815(.A(n4933), .B(n4930), .Y(n4934));
  NOR2X1  g3816(.A(n4437), .B(n4063), .Y(n4935));
  INVX1   g3817(.A(n4924), .Y(n4936));
  AOI22X1 g3818(.A0(n4447), .A1(n4936), .B0(n4440), .B1(PHYADDRPOINTER_REG_18__SCAN_IN), .Y(n4937));
  OAI21X1 g3819(.A0(n5914), .A1(n1058), .B0(n4937), .Y(n4938));
  NOR2X1  g3820(.A(n4938), .B(n4935), .Y(n4939));
  OAI21X1 g3821(.A0(n4934), .A1(n2120), .B0(n4939), .Y(U2968));
  OAI22X1 g3822(.A0(n1251), .A1(n1641), .B0(n1589), .B1(n1352), .Y(n4941));
  OAI22X1 g3823(.A0(n1261), .A1(n1644), .B0(n1583), .B1(n1326), .Y(n4942));
  OAI22X1 g3824(.A0(n1284), .A1(n1586), .B0(n1570), .B1(n1343), .Y(n4943));
  OAI22X1 g3825(.A0(n1342), .A1(n1571), .B0(n1648), .B1(n1359), .Y(n4944));
  NOR4X1  g3826(.A(n4943), .B(n4942), .C(n4941), .D(n4944), .Y(n4945));
  OAI22X1 g3827(.A0(n1263), .A1(n1574), .B0(n1575), .B1(n1243), .Y(n4946));
  OAI22X1 g3828(.A0(n1347), .A1(n1647), .B0(n1585), .B1(n1358), .Y(n4947));
  OAI22X1 g3829(.A0(n1348), .A1(n1579), .B0(n1588), .B1(n1332), .Y(n4948));
  OAI22X1 g3830(.A0(n1354), .A1(n1582), .B0(n1580), .B1(n1334), .Y(n4949));
  NOR4X1  g3831(.A(n4948), .B(n4947), .C(n4946), .D(n4949), .Y(n4950));
  AOI21X1 g3832(.A0(n4950), .A1(n4945), .B0(n4422), .Y(n4951));
  INVX1   g3833(.A(PHYADDRPOINTER_REG_19__SCAN_IN), .Y(n4952));
  NOR4X1  g3834(.A(n4922), .B(n4894), .C(n4895), .D(n4862), .Y(n4953));
  XOR2X1  g3835(.A(n4953), .B(n4952), .Y(n4954));
  AOI22X1 g3836(.A0(n4425), .A1(EAX_REG_19__SCAN_IN), .B0(PHYADDRPOINTER_REG_19__SCAN_IN), .B1(n4427), .Y(n4955));
  OAI21X1 g3837(.A0(n4954), .A1(n4419), .B0(n4955), .Y(n4956));
  AOI21X1 g3838(.A0(n4951), .A1(n4818), .B0(n4956), .Y(n4957));
  XOR2X1  g3839(.A(n4957), .B(n4418), .Y(n4958));
  INVX1   g3840(.A(n4958), .Y(n4959));
  XOR2X1  g3841(.A(n4959), .B(n4882), .Y(n4960));
  NOR3X1  g3842(.A(n4928), .B(n4422), .C(n4028), .Y(n4961));
  NOR3X1  g3843(.A(n4901), .B(n4422), .C(n4028), .Y(n4962));
  AOI22X1 g3844(.A0(n4902), .A1(n4929), .B0(n4462), .B1(n4058), .Y(n4963));
  NOR4X1  g3845(.A(n4867), .B(n4422), .C(n4028), .D(n4963), .Y(n4964));
  NOR3X1  g3846(.A(n4964), .B(n4962), .C(n4961), .Y(n4965));
  INVX1   g3847(.A(n4963), .Y(n4966));
  NAND2X1 g3848(.A(n4966), .B(n4870), .Y(n4967));
  OAI21X1 g3849(.A0(n4967), .A1(n4815), .B0(n4965), .Y(n4968));
  XOR2X1  g3850(.A(n4968), .B(n4960), .Y(n4969));
  INVX1   g3851(.A(n4954), .Y(n4970));
  AOI22X1 g3852(.A0(n4447), .A1(n4970), .B0(n4440), .B1(PHYADDRPOINTER_REG_19__SCAN_IN), .Y(n4971));
  OAI21X1 g3853(.A0(n5914), .A1(n1055), .B0(n4971), .Y(n4972));
  AOI21X1 g3854(.A0(n4969), .A1(n4441), .B0(n4972), .Y(n4973));
  OAI21X1 g3855(.A0(n4437), .A1(n4092), .B0(n4973), .Y(U2967));
  NAND2X1 g3856(.A(n4436), .B(n4120), .Y(n4975));
  AOI22X1 g3857(.A0(n1329), .A1(INSTQUEUE_REG_7__4__SCAN_IN), .B0(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n1266), .Y(n4976));
  AOI22X1 g3858(.A0(n1273), .A1(INSTQUEUE_REG_6__4__SCAN_IN), .B0(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n1246), .Y(n4977));
  AOI22X1 g3859(.A0(n1337), .A1(INSTQUEUE_REG_4__4__SCAN_IN), .B0(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n1244), .Y(n4978));
  AOI22X1 g3860(.A0(n1268), .A1(INSTQUEUE_REG_2__4__SCAN_IN), .B0(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n1279), .Y(n4979));
  NAND4X1 g3861(.A(n4978), .B(n4977), .C(n4976), .D(n4979), .Y(n4980));
  AOI22X1 g3862(.A0(n1338), .A1(INSTQUEUE_REG_11__4__SCAN_IN), .B0(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n1323), .Y(n4981));
  AOI22X1 g3863(.A0(n1270), .A1(INSTQUEUE_REG_8__4__SCAN_IN), .B0(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n1278), .Y(n4982));
  AOI22X1 g3864(.A0(n1271), .A1(INSTQUEUE_REG_15__4__SCAN_IN), .B0(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n1253), .Y(n4983));
  AOI22X1 g3865(.A0(n1275), .A1(INSTQUEUE_REG_12__4__SCAN_IN), .B0(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n1255), .Y(n4984));
  NAND4X1 g3866(.A(n4983), .B(n4982), .C(n4981), .D(n4984), .Y(n4985));
  OAI21X1 g3867(.A0(n4985), .A1(n4980), .B0(n4462), .Y(n4986));
  NOR2X1  g3868(.A(n4986), .B(n4817), .Y(n4987));
  NAND3X1 g3869(.A(n4923), .B(PHYADDRPOINTER_REG_19__SCAN_IN), .C(PHYADDRPOINTER_REG_18__SCAN_IN), .Y(n4988));
  XOR2X1  g3870(.A(n4988), .B(PHYADDRPOINTER_REG_20__SCAN_IN), .Y(n4989));
  AOI22X1 g3871(.A0(n4425), .A1(EAX_REG_20__SCAN_IN), .B0(PHYADDRPOINTER_REG_20__SCAN_IN), .B1(n4427), .Y(n4990));
  OAI21X1 g3872(.A0(n4989), .A1(n4419), .B0(n4990), .Y(n4991));
  NOR2X1  g3873(.A(n4991), .B(n4987), .Y(n4992));
  XOR2X1  g3874(.A(n4992), .B(n4418), .Y(n4993));
  XOR2X1  g3875(.A(n4993), .B(n4882), .Y(n4994));
  AOI21X1 g3876(.A0(n4462), .A1(n4058), .B0(n4959), .Y(n4995));
  NOR2X1  g3877(.A(n4965), .B(n4995), .Y(n4996));
  AOI21X1 g3878(.A0(n4959), .A1(n4882), .B0(n4996), .Y(n4997));
  NOR3X1  g3879(.A(n4963), .B(n4995), .C(n4869), .Y(n4998));
  OAI21X1 g3880(.A0(n4814), .A1(n4808), .B0(n4998), .Y(n4999));
  NAND2X1 g3881(.A(n4999), .B(n4997), .Y(n5000));
  NOR2X1  g3882(.A(n5000), .B(n4994), .Y(n5001));
  OAI21X1 g3883(.A0(n4422), .A1(n4028), .B0(n4993), .Y(n5002));
  NOR3X1  g3884(.A(n4993), .B(n4422), .C(n4028), .Y(n5003));
  AOI22X1 g3885(.A0(n5002), .A1(n5136), .B0(n4999), .B1(n4997), .Y(n5005));
  OAI21X1 g3886(.A0(n5005), .A1(n5001), .B0(n4441), .Y(n5006));
  NAND4X1 g3887(.A(n1910), .B(n1833), .C(REIP_REG_20__SCAN_IN), .D(n4439), .Y(n5007));
  INVX1   g3888(.A(n4989), .Y(n5008));
  AOI22X1 g3889(.A0(n4447), .A1(n5008), .B0(n4440), .B1(PHYADDRPOINTER_REG_20__SCAN_IN), .Y(n5009));
  NAND4X1 g3890(.A(n5007), .B(n5006), .C(n4975), .D(n5009), .Y(U2966));
  NAND3X1 g3891(.A(n4959), .B(n4462), .C(n4058), .Y(n5011));
  OAI21X1 g3892(.A0(n4965), .A1(n4995), .B0(n5011), .Y(n5012));
  NOR2X1  g3893(.A(n5003), .B(n5012), .Y(n5013));
  AOI22X1 g3894(.A0(n4999), .A1(n5013), .B0(n4993), .B1(n4931), .Y(n5014));
  INVX1   g3895(.A(PHYADDRPOINTER_REG_21__SCAN_IN), .Y(n5015));
  INVX1   g3896(.A(PHYADDRPOINTER_REG_20__SCAN_IN), .Y(n5016));
  NOR2X1  g3897(.A(n4988), .B(n5016), .Y(n5017));
  XOR2X1  g3898(.A(n5017), .B(n5015), .Y(n5018));
  INVX1   g3899(.A(n5018), .Y(n5019));
  AOI22X1 g3900(.A0(n1329), .A1(INSTQUEUE_REG_7__5__SCAN_IN), .B0(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n1273), .Y(n5020));
  AOI22X1 g3901(.A0(n1337), .A1(INSTQUEUE_REG_4__5__SCAN_IN), .B0(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n1246), .Y(n5021));
  AOI22X1 g3902(.A0(n1244), .A1(INSTQUEUE_REG_3__5__SCAN_IN), .B0(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n1268), .Y(n5022));
  AOI22X1 g3903(.A0(n1266), .A1(INSTQUEUE_REG_0__5__SCAN_IN), .B0(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n1279), .Y(n5023));
  NAND4X1 g3904(.A(n5022), .B(n5021), .C(n5020), .D(n5023), .Y(n5024));
  AOI22X1 g3905(.A0(n1338), .A1(INSTQUEUE_REG_11__5__SCAN_IN), .B0(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n1323), .Y(n5025));
  AOI22X1 g3906(.A0(n1270), .A1(INSTQUEUE_REG_8__5__SCAN_IN), .B0(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n1278), .Y(n5026));
  AOI22X1 g3907(.A0(n1271), .A1(INSTQUEUE_REG_15__5__SCAN_IN), .B0(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n1253), .Y(n5027));
  AOI22X1 g3908(.A0(n1275), .A1(INSTQUEUE_REG_12__5__SCAN_IN), .B0(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n1255), .Y(n5028));
  NAND4X1 g3909(.A(n5027), .B(n5026), .C(n5025), .D(n5028), .Y(n5029));
  OAI21X1 g3910(.A0(n5029), .A1(n5024), .B0(n4462), .Y(n5030));
  AOI22X1 g3911(.A0(n4425), .A1(EAX_REG_21__SCAN_IN), .B0(PHYADDRPOINTER_REG_21__SCAN_IN), .B1(n4427), .Y(n5031));
  OAI21X1 g3912(.A0(n5030), .A1(n4817), .B0(n5031), .Y(n5032));
  AOI21X1 g3913(.A0(n5019), .A1(n4418), .B0(n5032), .Y(n5033));
  XOR2X1  g3914(.A(n5033), .B(n4418), .Y(n5034));
  INVX1   g3915(.A(n5034), .Y(n5035));
  XOR2X1  g3916(.A(n5035), .B(n4882), .Y(n5036));
  NOR2X1  g3917(.A(n5036), .B(n5014), .Y(n5037));
  NAND3X1 g3918(.A(n5136), .B(n4999), .C(n4997), .Y(n5038));
  INVX1   g3919(.A(n4993), .Y(n5039));
  AOI22X1 g3920(.A0(n5039), .A1(n5035), .B0(n4462), .B1(n4058), .Y(n5040));
  AOI21X1 g3921(.A0(n5035), .A1(n4882), .B0(n5040), .Y(n5041));
  AOI21X1 g3922(.A0(n5041), .A1(n5038), .B0(n5037), .Y(n5042));
  AOI22X1 g3923(.A0(n4447), .A1(n5019), .B0(n4440), .B1(PHYADDRPOINTER_REG_21__SCAN_IN), .Y(n5043));
  OAI21X1 g3924(.A0(n5914), .A1(n1049), .B0(n5043), .Y(n5044));
  AOI21X1 g3925(.A0(n5042), .A1(n4441), .B0(n5044), .Y(n5045));
  OAI21X1 g3926(.A0(n4437), .A1(n4144), .B0(n5045), .Y(U2965));
  NAND2X1 g3927(.A(n4436), .B(n4171), .Y(n5047));
  INVX1   g3928(.A(PHYADDRPOINTER_REG_22__SCAN_IN), .Y(n5048));
  NOR3X1  g3929(.A(n4988), .B(n5015), .C(n5016), .Y(n5049));
  XOR2X1  g3930(.A(n5049), .B(n5048), .Y(n5050));
  INVX1   g3931(.A(n5050), .Y(n5051));
  AOI22X1 g3932(.A0(n1329), .A1(INSTQUEUE_REG_7__6__SCAN_IN), .B0(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n1273), .Y(n5052));
  AOI22X1 g3933(.A0(n1337), .A1(INSTQUEUE_REG_4__6__SCAN_IN), .B0(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n1246), .Y(n5053));
  AOI22X1 g3934(.A0(n1244), .A1(INSTQUEUE_REG_3__6__SCAN_IN), .B0(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n1268), .Y(n5054));
  AOI22X1 g3935(.A0(n1266), .A1(INSTQUEUE_REG_0__6__SCAN_IN), .B0(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n1279), .Y(n5055));
  NAND4X1 g3936(.A(n5054), .B(n5053), .C(n5052), .D(n5055), .Y(n5056));
  AOI22X1 g3937(.A0(n1338), .A1(INSTQUEUE_REG_11__6__SCAN_IN), .B0(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n1323), .Y(n5057));
  AOI22X1 g3938(.A0(n1270), .A1(INSTQUEUE_REG_8__6__SCAN_IN), .B0(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n1278), .Y(n5058));
  AOI22X1 g3939(.A0(n1271), .A1(INSTQUEUE_REG_15__6__SCAN_IN), .B0(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n1253), .Y(n5059));
  AOI22X1 g3940(.A0(n1275), .A1(INSTQUEUE_REG_12__6__SCAN_IN), .B0(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n1255), .Y(n5060));
  NAND4X1 g3941(.A(n5059), .B(n5058), .C(n5057), .D(n5060), .Y(n5061));
  OAI21X1 g3942(.A0(n5061), .A1(n5056), .B0(n4462), .Y(n5062));
  AOI22X1 g3943(.A0(n4425), .A1(EAX_REG_22__SCAN_IN), .B0(PHYADDRPOINTER_REG_22__SCAN_IN), .B1(n4427), .Y(n5063));
  OAI21X1 g3944(.A0(n5062), .A1(n4817), .B0(n5063), .Y(n5064));
  AOI21X1 g3945(.A0(n5051), .A1(n4418), .B0(n5064), .Y(n5065));
  XOR2X1  g3946(.A(n5065), .B(n4418), .Y(n5066));
  INVX1   g3947(.A(n5066), .Y(n5067));
  XOR2X1  g3948(.A(n5067), .B(n4882), .Y(n5068));
  INVX1   g3949(.A(n5068), .Y(n5069));
  NAND3X1 g3950(.A(n5035), .B(n4462), .C(n4058), .Y(n5070));
  INVX1   g3951(.A(n5070), .Y(n5071));
  OAI21X1 g3952(.A0(n4422), .A1(n4028), .B0(n5034), .Y(n5072));
  OAI21X1 g3953(.A0(n5071), .A1(n5014), .B0(n5072), .Y(n5073));
  XOR2X1  g3954(.A(n5073), .B(n5069), .Y(n5074));
  NAND2X1 g3955(.A(n5074), .B(n4441), .Y(n5075));
  NAND4X1 g3956(.A(n1910), .B(n1833), .C(REIP_REG_22__SCAN_IN), .D(n4439), .Y(n5076));
  AOI22X1 g3957(.A0(n4447), .A1(n5051), .B0(n4440), .B1(PHYADDRPOINTER_REG_22__SCAN_IN), .Y(n5077));
  NAND4X1 g3958(.A(n5076), .B(n5075), .C(n5047), .D(n5077), .Y(U2964));
  AOI22X1 g3959(.A0(n1323), .A1(INSTQUEUE_REG_11__0__SCAN_IN), .B0(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n1278), .Y(n5081));
  AOI22X1 g3960(.A0(n1329), .A1(INSTQUEUE_REG_8__0__SCAN_IN), .B0(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n1270), .Y(n5084));
  NAND2X1 g3961(.A(n5084), .B(n5081), .Y(n5085));
  AOI22X1 g3962(.A0(n1271), .A1(INSTQUEUE_REG_0__0__SCAN_IN), .B0(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n1279), .Y(n5088));
  AOI22X1 g3963(.A0(n1266), .A1(INSTQUEUE_REG_1__0__SCAN_IN), .B0(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n1268), .Y(n5091));
  NAND2X1 g3964(.A(n5091), .B(n5088), .Y(n5092));
  AOI22X1 g3965(.A0(n1253), .A1(INSTQUEUE_REG_15__0__SCAN_IN), .B0(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n1246), .Y(n5095));
  AOI22X1 g3966(.A0(n1337), .A1(INSTQUEUE_REG_5__0__SCAN_IN), .B0(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n1273), .Y(n5098));
  AOI22X1 g3967(.A0(n1255), .A1(INSTQUEUE_REG_14__0__SCAN_IN), .B0(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n1244), .Y(n5101));
  AOI22X1 g3968(.A0(n1338), .A1(INSTQUEUE_REG_12__0__SCAN_IN), .B0(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n1275), .Y(n5104));
  NAND4X1 g3969(.A(n5101), .B(n5098), .C(n5095), .D(n5104), .Y(n5105));
  NOR3X1  g3970(.A(n5105), .B(n5092), .C(n5085), .Y(n5106));
  NOR2X1  g3971(.A(n5106), .B(n4817), .Y(n5107));
  INVX1   g3972(.A(n5107), .Y(n5108));
  AOI22X1 g3973(.A0(n1329), .A1(INSTQUEUE_REG_7__7__SCAN_IN), .B0(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n1273), .Y(n5109));
  AOI22X1 g3974(.A0(n1337), .A1(INSTQUEUE_REG_4__7__SCAN_IN), .B0(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n1246), .Y(n5110));
  AOI22X1 g3975(.A0(n1244), .A1(INSTQUEUE_REG_3__7__SCAN_IN), .B0(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n1268), .Y(n5111));
  AOI22X1 g3976(.A0(n1266), .A1(INSTQUEUE_REG_0__7__SCAN_IN), .B0(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n1279), .Y(n5112));
  NAND4X1 g3977(.A(n5111), .B(n5110), .C(n5109), .D(n5112), .Y(n5113));
  AOI22X1 g3978(.A0(n1338), .A1(INSTQUEUE_REG_11__7__SCAN_IN), .B0(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n1323), .Y(n5114));
  AOI22X1 g3979(.A0(n1270), .A1(INSTQUEUE_REG_8__7__SCAN_IN), .B0(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n1278), .Y(n5115));
  AOI22X1 g3980(.A0(n1271), .A1(INSTQUEUE_REG_15__7__SCAN_IN), .B0(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n1253), .Y(n5116));
  AOI22X1 g3981(.A0(n1275), .A1(INSTQUEUE_REG_12__7__SCAN_IN), .B0(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n1255), .Y(n5117));
  NAND4X1 g3982(.A(n5116), .B(n5115), .C(n5114), .D(n5117), .Y(n5118));
  OAI21X1 g3983(.A0(n5118), .A1(n5113), .B0(n4818), .Y(n5119));
  OAI21X1 g3984(.A0(n5119), .A1(n5108), .B0(n4462), .Y(n5120));
  AOI21X1 g3985(.A0(n5119), .A1(n5108), .B0(n5120), .Y(n5121));
  NAND2X1 g3986(.A(n5049), .B(PHYADDRPOINTER_REG_22__SCAN_IN), .Y(n5122));
  XOR2X1  g3987(.A(n5122), .B(PHYADDRPOINTER_REG_23__SCAN_IN), .Y(n5123));
  AOI22X1 g3988(.A0(n4425), .A1(EAX_REG_23__SCAN_IN), .B0(PHYADDRPOINTER_REG_23__SCAN_IN), .B1(n4427), .Y(n5124));
  OAI21X1 g3989(.A0(n5123), .A1(n4419), .B0(n5124), .Y(n5125));
  NOR2X1  g3990(.A(n5125), .B(n5121), .Y(n5126));
  XOR2X1  g3991(.A(n5126), .B(n4418), .Y(n5127));
  INVX1   g3992(.A(n5127), .Y(n5128));
  XOR2X1  g3993(.A(n5128), .B(n4882), .Y(n5129));
  NOR3X1  g3994(.A(n5012), .B(n4814), .C(n4808), .Y(n5130));
  OAI21X1 g3995(.A0(n4422), .A1(n4028), .B0(n5066), .Y(n5131));
  INVX1   g3996(.A(n5131), .Y(n5132));
  NOR2X1  g3997(.A(n5132), .B(n5040), .Y(n5133));
  OAI21X1 g3998(.A0(n4998), .A1(n5012), .B0(n5133), .Y(n5134));
  NAND3X1 g3999(.A(n5067), .B(n4462), .C(n4058), .Y(n5135));
  NAND3X1 g4000(.A(n5039), .B(n4462), .C(n4058), .Y(n5136));
  NAND3X1 g4001(.A(n5136), .B(n5135), .C(n5070), .Y(n5137));
  NAND2X1 g4002(.A(n5137), .B(n5131), .Y(n5138));
  OAI21X1 g4003(.A0(n5134), .A1(n5130), .B0(n5138), .Y(n5139));
  XOR2X1  g4004(.A(n5139), .B(n5129), .Y(n5140));
  INVX1   g4005(.A(n5123), .Y(n5141));
  AOI22X1 g4006(.A0(n4447), .A1(n5141), .B0(n4440), .B1(PHYADDRPOINTER_REG_23__SCAN_IN), .Y(n5142));
  OAI21X1 g4007(.A0(n5914), .A1(n1043), .B0(n5142), .Y(n5143));
  AOI21X1 g4008(.A0(n5140), .A1(n4441), .B0(n5143), .Y(n5144));
  OAI21X1 g4009(.A0(n4437), .A1(n4198), .B0(n5144), .Y(U2963));
  NOR2X1  g4010(.A(n5119), .B(n5108), .Y(n5146));
  AOI22X1 g4011(.A0(n1323), .A1(INSTQUEUE_REG_11__1__SCAN_IN), .B0(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n1278), .Y(n5147));
  AOI22X1 g4012(.A0(n1329), .A1(INSTQUEUE_REG_8__1__SCAN_IN), .B0(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n1270), .Y(n5148));
  NAND2X1 g4013(.A(n5148), .B(n5147), .Y(n5149));
  AOI22X1 g4014(.A0(n1271), .A1(INSTQUEUE_REG_0__1__SCAN_IN), .B0(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n1279), .Y(n5150));
  AOI22X1 g4015(.A0(n1266), .A1(INSTQUEUE_REG_1__1__SCAN_IN), .B0(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n1268), .Y(n5151));
  NAND2X1 g4016(.A(n5151), .B(n5150), .Y(n5152));
  AOI22X1 g4017(.A0(n1253), .A1(INSTQUEUE_REG_15__1__SCAN_IN), .B0(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n1246), .Y(n5153));
  AOI22X1 g4018(.A0(n1337), .A1(INSTQUEUE_REG_5__1__SCAN_IN), .B0(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n1273), .Y(n5154));
  AOI22X1 g4019(.A0(n1255), .A1(INSTQUEUE_REG_14__1__SCAN_IN), .B0(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n1244), .Y(n5155));
  AOI22X1 g4020(.A0(n1338), .A1(INSTQUEUE_REG_12__1__SCAN_IN), .B0(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n1275), .Y(n5156));
  NAND4X1 g4021(.A(n5155), .B(n5154), .C(n5153), .D(n5156), .Y(n5157));
  NOR3X1  g4022(.A(n5157), .B(n5152), .C(n5149), .Y(n5158));
  NOR2X1  g4023(.A(n5158), .B(n4817), .Y(n5159));
  INVX1   g4024(.A(n5159), .Y(n5160));
  XOR2X1  g4025(.A(n5160), .B(n5146), .Y(n5161));
  INVX1   g4026(.A(PHYADDRPOINTER_REG_24__SCAN_IN), .Y(n5162));
  NAND3X1 g4027(.A(n5049), .B(PHYADDRPOINTER_REG_23__SCAN_IN), .C(PHYADDRPOINTER_REG_22__SCAN_IN), .Y(n5163));
  XOR2X1  g4028(.A(n5163), .B(n5162), .Y(n5164));
  INVX1   g4029(.A(EAX_REG_24__SCAN_IN), .Y(n5165));
  OAI22X1 g4030(.A0(n4426), .A1(n5165), .B0(n5162), .B1(n4479), .Y(n5166));
  AOI21X1 g4031(.A0(n5164), .A1(n4418), .B0(n5166), .Y(n5167));
  OAI21X1 g4032(.A0(n5161), .A1(n4422), .B0(n5167), .Y(n5168));
  XOR2X1  g4033(.A(n5168), .B(n4419), .Y(n5169));
  INVX1   g4034(.A(n5169), .Y(n5170));
  XOR2X1  g4035(.A(n5170), .B(n4882), .Y(n5171));
  INVX1   g4036(.A(n5171), .Y(n5172));
  OAI21X1 g4037(.A0(n4422), .A1(n4028), .B0(n5127), .Y(n5173));
  NOR3X1  g4038(.A(n5127), .B(n4422), .C(n4028), .Y(n5174));
  AOI21X1 g4039(.A0(n5139), .A1(n5173), .B0(n5174), .Y(n5175));
  XOR2X1  g4040(.A(n5175), .B(n5172), .Y(n5176));
  AOI22X1 g4041(.A0(n4447), .A1(n5164), .B0(n4440), .B1(PHYADDRPOINTER_REG_24__SCAN_IN), .Y(n5177));
  OAI21X1 g4042(.A0(n5914), .A1(n1040), .B0(n5177), .Y(n5178));
  AOI21X1 g4043(.A0(n5176), .A1(n4441), .B0(n5178), .Y(n5179));
  OAI21X1 g4044(.A0(n4437), .A1(n4222), .B0(n5179), .Y(U2962));
  NOR3X1  g4045(.A(n5160), .B(n5119), .C(n5108), .Y(n5181));
  AOI22X1 g4046(.A0(n1323), .A1(INSTQUEUE_REG_11__2__SCAN_IN), .B0(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n1278), .Y(n5182));
  AOI22X1 g4047(.A0(n1329), .A1(INSTQUEUE_REG_8__2__SCAN_IN), .B0(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n1270), .Y(n5183));
  NAND2X1 g4048(.A(n5183), .B(n5182), .Y(n5184));
  AOI22X1 g4049(.A0(n1271), .A1(INSTQUEUE_REG_0__2__SCAN_IN), .B0(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n1279), .Y(n5185));
  AOI22X1 g4050(.A0(n1266), .A1(INSTQUEUE_REG_1__2__SCAN_IN), .B0(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n1268), .Y(n5186));
  NAND2X1 g4051(.A(n5186), .B(n5185), .Y(n5187));
  AOI22X1 g4052(.A0(n1253), .A1(INSTQUEUE_REG_15__2__SCAN_IN), .B0(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n1246), .Y(n5188));
  AOI22X1 g4053(.A0(n1337), .A1(INSTQUEUE_REG_5__2__SCAN_IN), .B0(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n1273), .Y(n5189));
  AOI22X1 g4054(.A0(n1255), .A1(INSTQUEUE_REG_14__2__SCAN_IN), .B0(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n1244), .Y(n5190));
  AOI22X1 g4055(.A0(n1338), .A1(INSTQUEUE_REG_12__2__SCAN_IN), .B0(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n1275), .Y(n5191));
  NAND4X1 g4056(.A(n5190), .B(n5189), .C(n5188), .D(n5191), .Y(n5192));
  NOR3X1  g4057(.A(n5192), .B(n5187), .C(n5184), .Y(n5193));
  NOR2X1  g4058(.A(n5193), .B(n4817), .Y(n5194));
  INVX1   g4059(.A(n5194), .Y(n5195));
  XOR2X1  g4060(.A(n5195), .B(n5181), .Y(n5196));
  INVX1   g4061(.A(PHYADDRPOINTER_REG_25__SCAN_IN), .Y(n5197));
  NAND4X1 g4062(.A(PHYADDRPOINTER_REG_24__SCAN_IN), .B(PHYADDRPOINTER_REG_23__SCAN_IN), .C(PHYADDRPOINTER_REG_22__SCAN_IN), .D(n5049), .Y(n5198));
  XOR2X1  g4063(.A(n5198), .B(n5197), .Y(n5199));
  INVX1   g4064(.A(EAX_REG_25__SCAN_IN), .Y(n5200));
  OAI22X1 g4065(.A0(n4426), .A1(n5200), .B0(n5197), .B1(n4479), .Y(n5201));
  AOI21X1 g4066(.A0(n5199), .A1(n4418), .B0(n5201), .Y(n5202));
  OAI21X1 g4067(.A0(n5196), .A1(n4422), .B0(n5202), .Y(n5203));
  XOR2X1  g4068(.A(n5203), .B(n4419), .Y(n5204));
  INVX1   g4069(.A(n5204), .Y(n5205));
  XOR2X1  g4070(.A(n5205), .B(n4882), .Y(n5206));
  OAI22X1 g4071(.A0(n5127), .A1(n5169), .B0(n4422), .B1(n4028), .Y(n5207));
  NAND4X1 g4072(.A(n5131), .B(n5072), .C(n5002), .D(n5207), .Y(n5208));
  NOR4X1  g4073(.A(n4963), .B(n4995), .C(n4869), .D(n5208), .Y(n5209));
  OAI21X1 g4074(.A0(n4814), .A1(n4808), .B0(n5209), .Y(n5210));
  INVX1   g4075(.A(n5208), .Y(n5211));
  INVX1   g4076(.A(n5207), .Y(n5212));
  AOI21X1 g4077(.A0(n5137), .A1(n5131), .B0(n5174), .Y(n5213));
  OAI22X1 g4078(.A0(n5212), .A1(n5213), .B0(n5169), .B1(n4931), .Y(n5214));
  AOI21X1 g4079(.A0(n5211), .A1(n5012), .B0(n5214), .Y(n5215));
  NAND2X1 g4080(.A(n5215), .B(n5210), .Y(n5216));
  XOR2X1  g4081(.A(n5216), .B(n5206), .Y(n5217));
  AOI22X1 g4082(.A0(n4447), .A1(n5199), .B0(n4440), .B1(PHYADDRPOINTER_REG_25__SCAN_IN), .Y(n5218));
  OAI21X1 g4083(.A0(n5914), .A1(n1037), .B0(n5218), .Y(n5219));
  AOI21X1 g4084(.A0(n5217), .A1(n4441), .B0(n5219), .Y(n5220));
  OAI21X1 g4085(.A0(n4437), .A1(n4249), .B0(n5220), .Y(U2961));
  AOI22X1 g4086(.A0(n1323), .A1(INSTQUEUE_REG_11__3__SCAN_IN), .B0(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n1278), .Y(n5222));
  AOI22X1 g4087(.A0(n1329), .A1(INSTQUEUE_REG_8__3__SCAN_IN), .B0(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n1270), .Y(n5223));
  NAND2X1 g4088(.A(n5223), .B(n5222), .Y(n5224));
  AOI22X1 g4089(.A0(n1271), .A1(INSTQUEUE_REG_0__3__SCAN_IN), .B0(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n1279), .Y(n5225));
  AOI22X1 g4090(.A0(n1266), .A1(INSTQUEUE_REG_1__3__SCAN_IN), .B0(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n1268), .Y(n5226));
  NAND2X1 g4091(.A(n5226), .B(n5225), .Y(n5227));
  AOI22X1 g4092(.A0(n1253), .A1(INSTQUEUE_REG_15__3__SCAN_IN), .B0(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n1246), .Y(n5228));
  AOI22X1 g4093(.A0(n1337), .A1(INSTQUEUE_REG_5__3__SCAN_IN), .B0(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n1273), .Y(n5229));
  AOI22X1 g4094(.A0(n1255), .A1(INSTQUEUE_REG_14__3__SCAN_IN), .B0(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n1244), .Y(n5230));
  AOI22X1 g4095(.A0(n1338), .A1(INSTQUEUE_REG_12__3__SCAN_IN), .B0(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n1275), .Y(n5231));
  NAND4X1 g4096(.A(n5230), .B(n5229), .C(n5228), .D(n5231), .Y(n5232));
  NOR3X1  g4097(.A(n5232), .B(n5227), .C(n5224), .Y(n5233));
  NOR2X1  g4098(.A(n5233), .B(n4817), .Y(n5234));
  INVX1   g4099(.A(n5234), .Y(n5235));
  NOR4X1  g4100(.A(n5160), .B(n5119), .C(n5108), .D(n5195), .Y(n5236));
  XOR2X1  g4101(.A(n5236), .B(n5235), .Y(n5237));
  NOR3X1  g4102(.A(n5163), .B(n5197), .C(n5162), .Y(n5238));
  XOR2X1  g4103(.A(n5238), .B(PHYADDRPOINTER_REG_26__SCAN_IN), .Y(n5239));
  INVX1   g4104(.A(EAX_REG_26__SCAN_IN), .Y(n5240));
  NAND3X1 g4105(.A(PHYADDRPOINTER_REG_26__SCAN_IN), .B(n1833), .C(STATEBS16_REG_SCAN_IN), .Y(n5241));
  OAI21X1 g4106(.A0(n4426), .A1(n5240), .B0(n5241), .Y(n5242));
  AOI21X1 g4107(.A0(n5239), .A1(n4418), .B0(n5242), .Y(n5243));
  OAI21X1 g4108(.A0(n5237), .A1(n4422), .B0(n5243), .Y(n5244));
  XOR2X1  g4109(.A(n5244), .B(n4419), .Y(n5245));
  INVX1   g4110(.A(n5245), .Y(n5246));
  XOR2X1  g4111(.A(n5246), .B(n4882), .Y(n5247));
  AOI21X1 g4112(.A0(n4462), .A1(n4058), .B0(n5205), .Y(n5248));
  AOI21X1 g4113(.A0(n5215), .A1(n5210), .B0(n5248), .Y(n5249));
  AOI21X1 g4114(.A0(n5205), .A1(n4882), .B0(n5249), .Y(n5250));
  XOR2X1  g4115(.A(n5250), .B(n5247), .Y(n5251));
  NOR2X1  g4116(.A(n4437), .B(n4278), .Y(n5252));
  AOI22X1 g4117(.A0(n4447), .A1(n5239), .B0(n4440), .B1(PHYADDRPOINTER_REG_26__SCAN_IN), .Y(n5253));
  OAI21X1 g4118(.A0(n5914), .A1(n1034), .B0(n5253), .Y(n5254));
  NOR2X1  g4119(.A(n5254), .B(n5252), .Y(n5255));
  OAI21X1 g4120(.A0(n5251), .A1(n2120), .B0(n5255), .Y(U2960));
  NAND2X1 g4121(.A(n4436), .B(n4300), .Y(n5257));
  INVX1   g4122(.A(n5236), .Y(n5258));
  NOR2X1  g4123(.A(n5258), .B(n5235), .Y(n5259));
  AOI22X1 g4124(.A0(n1323), .A1(INSTQUEUE_REG_11__4__SCAN_IN), .B0(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n1278), .Y(n5260));
  AOI22X1 g4125(.A0(n1329), .A1(INSTQUEUE_REG_8__4__SCAN_IN), .B0(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n1270), .Y(n5261));
  NAND2X1 g4126(.A(n5261), .B(n5260), .Y(n5262));
  AOI22X1 g4127(.A0(n1271), .A1(INSTQUEUE_REG_0__4__SCAN_IN), .B0(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n1268), .Y(n5263));
  AOI22X1 g4128(.A0(n1279), .A1(INSTQUEUE_REG_2__4__SCAN_IN), .B0(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n1266), .Y(n5264));
  NAND2X1 g4129(.A(n5264), .B(n5263), .Y(n5265));
  AOI22X1 g4130(.A0(n1273), .A1(INSTQUEUE_REG_7__4__SCAN_IN), .B0(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n1275), .Y(n5266));
  AOI22X1 g4131(.A0(n1253), .A1(INSTQUEUE_REG_15__4__SCAN_IN), .B0(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n1337), .Y(n5267));
  AOI22X1 g4132(.A0(n1246), .A1(INSTQUEUE_REG_6__4__SCAN_IN), .B0(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n1255), .Y(n5268));
  AOI22X1 g4133(.A0(n1244), .A1(INSTQUEUE_REG_4__4__SCAN_IN), .B0(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n1338), .Y(n5269));
  NAND4X1 g4134(.A(n5268), .B(n5267), .C(n5266), .D(n5269), .Y(n5270));
  NOR3X1  g4135(.A(n5270), .B(n5265), .C(n5262), .Y(n5271));
  NOR2X1  g4136(.A(n5271), .B(n4817), .Y(n5272));
  XOR2X1  g4137(.A(n5272), .B(n5259), .Y(n5273));
  NAND2X1 g4138(.A(n5238), .B(PHYADDRPOINTER_REG_26__SCAN_IN), .Y(n5274));
  XOR2X1  g4139(.A(n5274), .B(PHYADDRPOINTER_REG_27__SCAN_IN), .Y(n5275));
  AOI22X1 g4140(.A0(n4425), .A1(EAX_REG_27__SCAN_IN), .B0(PHYADDRPOINTER_REG_27__SCAN_IN), .B1(n4427), .Y(n5276));
  OAI21X1 g4141(.A0(n5275), .A1(n4419), .B0(n5276), .Y(n5277));
  AOI21X1 g4142(.A0(n5273), .A1(n4462), .B0(n5277), .Y(n5278));
  XOR2X1  g4143(.A(n5278), .B(n4418), .Y(n5279));
  XOR2X1  g4144(.A(n5279), .B(n4931), .Y(n5280));
  INVX1   g4145(.A(n5280), .Y(n5281));
  OAI21X1 g4146(.A0(n4422), .A1(n4028), .B0(n5245), .Y(n5282));
  AOI21X1 g4147(.A0(n5245), .A1(n5204), .B0(n4931), .Y(n5283));
  OAI21X1 g4148(.A0(n5283), .A1(n5249), .B0(n5282), .Y(n5284));
  XOR2X1  g4149(.A(n5284), .B(n5281), .Y(n5285));
  NAND2X1 g4150(.A(n5285), .B(n4441), .Y(n5286));
  NAND4X1 g4151(.A(n1910), .B(n1833), .C(REIP_REG_27__SCAN_IN), .D(n4439), .Y(n5287));
  INVX1   g4152(.A(n5275), .Y(n5288));
  AOI22X1 g4153(.A0(n4447), .A1(n5288), .B0(n4440), .B1(PHYADDRPOINTER_REG_27__SCAN_IN), .Y(n5289));
  NAND4X1 g4154(.A(n5287), .B(n5286), .C(n5257), .D(n5289), .Y(U2959));
  AOI22X1 g4155(.A0(n1323), .A1(INSTQUEUE_REG_11__5__SCAN_IN), .B0(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n1278), .Y(n5291));
  AOI22X1 g4156(.A0(n1329), .A1(INSTQUEUE_REG_8__5__SCAN_IN), .B0(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n1270), .Y(n5292));
  NAND2X1 g4157(.A(n5292), .B(n5291), .Y(n5293));
  AOI22X1 g4158(.A0(n1271), .A1(INSTQUEUE_REG_0__5__SCAN_IN), .B0(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n1279), .Y(n5294));
  AOI22X1 g4159(.A0(n1266), .A1(INSTQUEUE_REG_1__5__SCAN_IN), .B0(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n1268), .Y(n5295));
  NAND2X1 g4160(.A(n5295), .B(n5294), .Y(n5296));
  AOI22X1 g4161(.A0(n1253), .A1(INSTQUEUE_REG_15__5__SCAN_IN), .B0(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n1246), .Y(n5297));
  AOI22X1 g4162(.A0(n1337), .A1(INSTQUEUE_REG_5__5__SCAN_IN), .B0(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n1273), .Y(n5298));
  AOI22X1 g4163(.A0(n1255), .A1(INSTQUEUE_REG_14__5__SCAN_IN), .B0(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n1244), .Y(n5299));
  AOI22X1 g4164(.A0(n1338), .A1(INSTQUEUE_REG_12__5__SCAN_IN), .B0(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n1275), .Y(n5300));
  NAND4X1 g4165(.A(n5299), .B(n5298), .C(n5297), .D(n5300), .Y(n5301));
  NOR3X1  g4166(.A(n5301), .B(n5296), .C(n5293), .Y(n5302));
  NOR2X1  g4167(.A(n5302), .B(n4817), .Y(n5303));
  NOR4X1  g4168(.A(n5258), .B(n5235), .C(n4817), .D(n5271), .Y(n5304));
  XOR2X1  g4169(.A(n5304), .B(n5303), .Y(n5305));
  NAND2X1 g4170(.A(n5305), .B(n4462), .Y(n5306));
  INVX1   g4171(.A(PHYADDRPOINTER_REG_28__SCAN_IN), .Y(n5307));
  NAND3X1 g4172(.A(n5238), .B(PHYADDRPOINTER_REG_27__SCAN_IN), .C(PHYADDRPOINTER_REG_26__SCAN_IN), .Y(n5308));
  XOR2X1  g4173(.A(n5308), .B(n5307), .Y(n5309));
  INVX1   g4174(.A(EAX_REG_28__SCAN_IN), .Y(n5310));
  OAI22X1 g4175(.A0(n4426), .A1(n5310), .B0(n5307), .B1(n4479), .Y(n5311));
  AOI21X1 g4176(.A0(n5309), .A1(n4418), .B0(n5311), .Y(n5312));
  NAND2X1 g4177(.A(n5312), .B(n5306), .Y(n5313));
  XOR2X1  g4178(.A(n5313), .B(n4419), .Y(n5314));
  NOR3X1  g4179(.A(n5314), .B(n4422), .C(n4028), .Y(n5315));
  INVX1   g4180(.A(n5314), .Y(n5316));
  AOI21X1 g4181(.A0(n4462), .A1(n4058), .B0(n5316), .Y(n5317));
  NOR2X1  g4182(.A(n5317), .B(n5315), .Y(n5318));
  NOR4X1  g4183(.A(n4775), .B(n4782), .C(n4760), .D(n4795), .Y(n5319));
  NOR2X1  g4184(.A(n4422), .B(n3960), .Y(n5320));
  AOI21X1 g4185(.A0(n4794), .A1(n5320), .B0(n4774), .Y(n5321));
  NAND2X1 g4186(.A(n4784), .B(n4750), .Y(n5322));
  AOI21X1 g4187(.A0(n5322), .A1(n5321), .B0(n4795), .Y(n5323));
  NOR2X1  g4188(.A(n5323), .B(n5319), .Y(n5324));
  OAI21X1 g4189(.A0(n4807), .A1(n4723), .B0(n5324), .Y(n5325));
  NOR2X1  g4190(.A(n5213), .B(n5212), .Y(n5326));
  AOI21X1 g4191(.A0(n5170), .A1(n4882), .B0(n5326), .Y(n5327));
  OAI21X1 g4192(.A0(n5208), .A1(n4997), .B0(n5327), .Y(n5328));
  AOI21X1 g4193(.A0(n5209), .A1(n5325), .B0(n5328), .Y(n5329));
  INVX1   g4194(.A(n5248), .Y(n5330));
  OAI21X1 g4195(.A0(n4422), .A1(n4028), .B0(n5279), .Y(n5331));
  NAND3X1 g4196(.A(n5331), .B(n5282), .C(n5330), .Y(n5332));
  NOR3X1  g4197(.A(n5279), .B(n4422), .C(n4028), .Y(n5333));
  OAI21X1 g4198(.A0(n5246), .A1(n5205), .B0(n4882), .Y(n5334));
  NOR2X1  g4199(.A(n5283), .B(n5333), .Y(n5336));
  OAI21X1 g4200(.A0(n5332), .A1(n5329), .B0(n5336), .Y(n5337));
  XOR2X1  g4201(.A(n5337), .B(n5318), .Y(n5338));
  AOI22X1 g4202(.A0(n4447), .A1(n5309), .B0(n4440), .B1(PHYADDRPOINTER_REG_28__SCAN_IN), .Y(n5339));
  OAI21X1 g4203(.A0(n5914), .A1(n1028), .B0(n5339), .Y(n5340));
  AOI21X1 g4204(.A0(n5338), .A1(n4441), .B0(n5340), .Y(n5341));
  OAI21X1 g4205(.A0(n4437), .A1(n4324), .B0(n5341), .Y(U2958));
  NAND4X1 g4206(.A(n5272), .B(n5236), .C(n5234), .D(n5303), .Y(n5343));
  AOI22X1 g4207(.A0(n1323), .A1(INSTQUEUE_REG_11__6__SCAN_IN), .B0(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n1278), .Y(n5344));
  AOI22X1 g4208(.A0(n1329), .A1(INSTQUEUE_REG_8__6__SCAN_IN), .B0(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n1270), .Y(n5345));
  NAND2X1 g4209(.A(n5345), .B(n5344), .Y(n5346));
  AOI22X1 g4210(.A0(n1271), .A1(INSTQUEUE_REG_0__6__SCAN_IN), .B0(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n1279), .Y(n5347));
  AOI22X1 g4211(.A0(n1266), .A1(INSTQUEUE_REG_1__6__SCAN_IN), .B0(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n1268), .Y(n5348));
  NAND2X1 g4212(.A(n5348), .B(n5347), .Y(n5349));
  AOI22X1 g4213(.A0(n1253), .A1(INSTQUEUE_REG_15__6__SCAN_IN), .B0(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n1246), .Y(n5350));
  AOI22X1 g4214(.A0(n1337), .A1(INSTQUEUE_REG_5__6__SCAN_IN), .B0(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n1273), .Y(n5351));
  AOI22X1 g4215(.A0(n1255), .A1(INSTQUEUE_REG_14__6__SCAN_IN), .B0(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n1244), .Y(n5352));
  AOI22X1 g4216(.A0(n1338), .A1(INSTQUEUE_REG_12__6__SCAN_IN), .B0(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n1275), .Y(n5353));
  NAND4X1 g4217(.A(n5352), .B(n5351), .C(n5350), .D(n5353), .Y(n5354));
  NOR3X1  g4218(.A(n5354), .B(n5349), .C(n5346), .Y(n5355));
  NOR2X1  g4219(.A(n5355), .B(n4817), .Y(n5356));
  XOR2X1  g4220(.A(n5356), .B(n5343), .Y(n5357));
  INVX1   g4221(.A(PHYADDRPOINTER_REG_29__SCAN_IN), .Y(n5358));
  NAND4X1 g4222(.A(PHYADDRPOINTER_REG_28__SCAN_IN), .B(PHYADDRPOINTER_REG_27__SCAN_IN), .C(PHYADDRPOINTER_REG_26__SCAN_IN), .D(n5238), .Y(n5359));
  XOR2X1  g4223(.A(n5359), .B(n5358), .Y(n5360));
  INVX1   g4224(.A(EAX_REG_29__SCAN_IN), .Y(n5361));
  OAI22X1 g4225(.A0(n4426), .A1(n5361), .B0(n5358), .B1(n4479), .Y(n5362));
  AOI21X1 g4226(.A0(n5360), .A1(n4418), .B0(n5362), .Y(n5363));
  OAI21X1 g4227(.A0(n5357), .A1(n4422), .B0(n5363), .Y(n5364));
  XOR2X1  g4228(.A(n5364), .B(n4419), .Y(n5365));
  INVX1   g4229(.A(n5365), .Y(n5366));
  XOR2X1  g4230(.A(n5366), .B(n4882), .Y(n5367));
  OAI22X1 g4231(.A0(n5245), .A1(n5314), .B0(n4422), .B1(n4028), .Y(n5368));
  NAND3X1 g4232(.A(n5368), .B(n5331), .C(n5330), .Y(n5369));
  NOR3X1  g4233(.A(n5283), .B(n5315), .C(n5333), .Y(n5370));
  OAI22X1 g4234(.A0(n5369), .A1(n5329), .B0(n5317), .B1(n5370), .Y(n5371));
  XOR2X1  g4235(.A(n5371), .B(n5367), .Y(n5372));
  AOI22X1 g4236(.A0(n4447), .A1(n5360), .B0(n4440), .B1(PHYADDRPOINTER_REG_29__SCAN_IN), .Y(n5373));
  OAI21X1 g4237(.A0(n5914), .A1(n1025), .B0(n5373), .Y(n5374));
  AOI21X1 g4238(.A0(n5372), .A1(n4441), .B0(n5374), .Y(n5375));
  OAI21X1 g4239(.A0(n4437), .A1(n4352), .B0(n5375), .Y(U2957));
  NOR3X1  g4240(.A(n5355), .B(n5343), .C(n4817), .Y(n5377));
  AOI22X1 g4241(.A0(n1323), .A1(INSTQUEUE_REG_11__7__SCAN_IN), .B0(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n1278), .Y(n5378));
  AOI22X1 g4242(.A0(n1329), .A1(INSTQUEUE_REG_8__7__SCAN_IN), .B0(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n1270), .Y(n5379));
  NAND2X1 g4243(.A(n5379), .B(n5378), .Y(n5380));
  AOI22X1 g4244(.A0(n1271), .A1(INSTQUEUE_REG_0__7__SCAN_IN), .B0(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n1279), .Y(n5381));
  AOI22X1 g4245(.A0(n1266), .A1(INSTQUEUE_REG_1__7__SCAN_IN), .B0(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n1268), .Y(n5382));
  NAND2X1 g4246(.A(n5382), .B(n5381), .Y(n5383));
  AOI22X1 g4247(.A0(n1253), .A1(INSTQUEUE_REG_15__7__SCAN_IN), .B0(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n1246), .Y(n5384));
  AOI22X1 g4248(.A0(n1337), .A1(INSTQUEUE_REG_5__7__SCAN_IN), .B0(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n1273), .Y(n5385));
  AOI22X1 g4249(.A0(n1255), .A1(INSTQUEUE_REG_14__7__SCAN_IN), .B0(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n1244), .Y(n5386));
  AOI22X1 g4250(.A0(n1338), .A1(INSTQUEUE_REG_12__7__SCAN_IN), .B0(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n1275), .Y(n5387));
  NAND4X1 g4251(.A(n5386), .B(n5385), .C(n5384), .D(n5387), .Y(n5388));
  NOR3X1  g4252(.A(n5388), .B(n5383), .C(n5380), .Y(n5389));
  NOR2X1  g4253(.A(n5389), .B(n4817), .Y(n5390));
  XOR2X1  g4254(.A(n5390), .B(n5377), .Y(n5391));
  NOR2X1  g4255(.A(n5359), .B(n5358), .Y(n5392));
  XOR2X1  g4256(.A(n5392), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .Y(n5393));
  INVX1   g4257(.A(n5393), .Y(n5394));
  AOI22X1 g4258(.A0(n4425), .A1(EAX_REG_30__SCAN_IN), .B0(PHYADDRPOINTER_REG_30__SCAN_IN), .B1(n4427), .Y(n5395));
  OAI21X1 g4259(.A0(n5394), .A1(n4419), .B0(n5395), .Y(n5396));
  AOI21X1 g4260(.A0(n5391), .A1(n4462), .B0(n5396), .Y(n5397));
  XOR2X1  g4261(.A(n5397), .B(n4419), .Y(n5398));
  XOR2X1  g4262(.A(n5398), .B(n4882), .Y(n5399));
  NOR2X1  g4263(.A(n5315), .B(n5333), .Y(n5400));
  AOI22X1 g4264(.A0(n5316), .A1(n5366), .B0(n4462), .B1(n4058), .Y(n5401));
  AOI21X1 g4265(.A0(n5400), .A1(n5334), .B0(n5401), .Y(n5402));
  AOI21X1 g4266(.A0(n5366), .A1(n4882), .B0(n5402), .Y(n5403));
  AOI21X1 g4267(.A0(n4462), .A1(n4058), .B0(n5366), .Y(n5404));
  INVX1   g4268(.A(n5404), .Y(n5405));
  NAND4X1 g4269(.A(n5405), .B(n5331), .C(n5330), .D(n5368), .Y(n5406));
  OAI21X1 g4270(.A0(n5406), .A1(n5329), .B0(n5403), .Y(n5407));
  XOR2X1  g4271(.A(n5407), .B(n5399), .Y(n5408));
  AOI22X1 g4272(.A0(n4447), .A1(n5393), .B0(n4440), .B1(PHYADDRPOINTER_REG_30__SCAN_IN), .Y(n5409));
  OAI21X1 g4273(.A0(n5914), .A1(n1020), .B0(n5409), .Y(n5410));
  AOI21X1 g4274(.A0(n5408), .A1(n4441), .B0(n5410), .Y(n5411));
  OAI21X1 g4275(.A0(n4437), .A1(n4378), .B0(n5411), .Y(U2956));
  AOI21X1 g4276(.A0(n4462), .A1(n4058), .B0(n5398), .Y(n5413));
  NOR3X1  g4277(.A(n5413), .B(n5369), .C(n5404), .Y(n5414));
  NAND3X1 g4278(.A(n5414), .B(n5211), .C(n4998), .Y(n5415));
  NOR2X1  g4279(.A(n5415), .B(n4815), .Y(n5416));
  NOR2X1  g4280(.A(n5403), .B(n5413), .Y(n5419));
  AOI21X1 g4281(.A0(n5398), .A1(n4882), .B0(n5419), .Y(n5420));
  NAND3X1 g4282(.A(n5420), .B(n4997), .C(n5327), .Y(n5421));
  NOR2X1  g4283(.A(n5421), .B(n5416), .Y(n5422));
  NAND2X1 g4284(.A(n5392), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .Y(n5423));
  XOR2X1  g4285(.A(n5423), .B(PHYADDRPOINTER_REG_31__SCAN_IN), .Y(n5424));
  INVX1   g4286(.A(n5424), .Y(n5425));
  NAND3X1 g4287(.A(PHYADDRPOINTER_REG_31__SCAN_IN), .B(n1833), .C(STATEBS16_REG_SCAN_IN), .Y(n5426));
  NAND3X1 g4288(.A(n1700), .B(EAX_REG_31__SCAN_IN), .C(STATE2_REG_2__SCAN_IN), .Y(n5427));
  NAND2X1 g4289(.A(n5427), .B(n5426), .Y(n5428));
  AOI21X1 g4290(.A0(n5425), .A1(n4418), .B0(n5428), .Y(n5429));
  XOR2X1  g4291(.A(n5429), .B(n4418), .Y(n5430));
  XOR2X1  g4292(.A(n5430), .B(n5422), .Y(n5431));
  INVX1   g4293(.A(REIP_REG_31__SCAN_IN), .Y(n5432));
  AOI22X1 g4294(.A0(n4447), .A1(n5425), .B0(n4440), .B1(PHYADDRPOINTER_REG_31__SCAN_IN), .Y(n5433));
  OAI21X1 g4295(.A0(n5914), .A1(n5432), .B0(n5433), .Y(n5434));
  AOI21X1 g4296(.A0(n5431), .A1(n4441), .B0(n5434), .Y(n5435));
  OAI21X1 g4297(.A0(n4437), .A1(n4401), .B0(n5435), .Y(U2955));
  OAI21X1 g4298(.A0(n1362), .A1(n1282), .B0(READY_N), .Y(n5437));
  NAND4X1 g4299(.A(n2083), .B(n1536), .C(n1447), .D(n5437), .Y(n5438));
  NOR2X1  g4300(.A(n5438), .B(n1464), .Y(n5439));
  NOR2X1  g4301(.A(n5438), .B(n1362), .Y(n5440));
  AOI22X1 g4302(.A0(n5439), .A1(DATAI_15_), .B0(EAX_REG_15__SCAN_IN), .B1(n5440), .Y(n5441));
  OAI21X1 g4303(.A0(n5438), .A1(n1825), .B0(LWORD_REG_15__SCAN_IN), .Y(n5442));
  OAI21X1 g4304(.A0(n5441), .A1(n1825), .B0(n5442), .Y(U2954));
  AOI22X1 g4305(.A0(n5439), .A1(DATAI_14_), .B0(EAX_REG_14__SCAN_IN), .B1(n5440), .Y(n5444));
  OAI21X1 g4306(.A0(n5438), .A1(n1825), .B0(LWORD_REG_14__SCAN_IN), .Y(n5445));
  OAI21X1 g4307(.A0(n5444), .A1(n1825), .B0(n5445), .Y(U2953));
  AOI22X1 g4308(.A0(n5439), .A1(DATAI_13_), .B0(EAX_REG_13__SCAN_IN), .B1(n5440), .Y(n5447));
  OAI21X1 g4309(.A0(n5438), .A1(n1825), .B0(LWORD_REG_13__SCAN_IN), .Y(n5448));
  OAI21X1 g4310(.A0(n5447), .A1(n1825), .B0(n5448), .Y(U2952));
  AOI22X1 g4311(.A0(n5439), .A1(DATAI_12_), .B0(EAX_REG_12__SCAN_IN), .B1(n5440), .Y(n5450));
  OAI21X1 g4312(.A0(n5438), .A1(n1825), .B0(LWORD_REG_12__SCAN_IN), .Y(n5451));
  OAI21X1 g4313(.A0(n5450), .A1(n1825), .B0(n5451), .Y(U2951));
  AOI22X1 g4314(.A0(n5439), .A1(DATAI_11_), .B0(EAX_REG_11__SCAN_IN), .B1(n5440), .Y(n5453));
  OAI21X1 g4315(.A0(n5438), .A1(n1825), .B0(LWORD_REG_11__SCAN_IN), .Y(n5454));
  OAI21X1 g4316(.A0(n5453), .A1(n1825), .B0(n5454), .Y(U2950));
  AOI22X1 g4317(.A0(n5439), .A1(DATAI_10_), .B0(EAX_REG_10__SCAN_IN), .B1(n5440), .Y(n5456));
  OAI21X1 g4318(.A0(n5438), .A1(n1825), .B0(LWORD_REG_10__SCAN_IN), .Y(n5457));
  OAI21X1 g4319(.A0(n5456), .A1(n1825), .B0(n5457), .Y(U2949));
  AOI22X1 g4320(.A0(n5439), .A1(DATAI_9_), .B0(EAX_REG_9__SCAN_IN), .B1(n5440), .Y(n5459));
  OAI21X1 g4321(.A0(n5438), .A1(n1825), .B0(LWORD_REG_9__SCAN_IN), .Y(n5460));
  OAI21X1 g4322(.A0(n5459), .A1(n1825), .B0(n5460), .Y(U2948));
  AOI22X1 g4323(.A0(n5439), .A1(DATAI_8_), .B0(EAX_REG_8__SCAN_IN), .B1(n5440), .Y(n5462));
  OAI21X1 g4324(.A0(n5438), .A1(n1825), .B0(LWORD_REG_8__SCAN_IN), .Y(n5463));
  OAI21X1 g4325(.A0(n5462), .A1(n1825), .B0(n5463), .Y(U2947));
  AOI22X1 g4326(.A0(n5439), .A1(DATAI_7_), .B0(EAX_REG_7__SCAN_IN), .B1(n5440), .Y(n5465));
  OAI21X1 g4327(.A0(n5438), .A1(n1825), .B0(LWORD_REG_7__SCAN_IN), .Y(n5466));
  OAI21X1 g4328(.A0(n5465), .A1(n1825), .B0(n5466), .Y(U2946));
  AOI22X1 g4329(.A0(n5439), .A1(DATAI_6_), .B0(EAX_REG_6__SCAN_IN), .B1(n5440), .Y(n5468));
  OAI21X1 g4330(.A0(n5438), .A1(n1825), .B0(LWORD_REG_6__SCAN_IN), .Y(n5469));
  OAI21X1 g4331(.A0(n5468), .A1(n1825), .B0(n5469), .Y(U2945));
  AOI22X1 g4332(.A0(n5439), .A1(DATAI_5_), .B0(EAX_REG_5__SCAN_IN), .B1(n5440), .Y(n5471));
  OAI21X1 g4333(.A0(n5438), .A1(n1825), .B0(LWORD_REG_5__SCAN_IN), .Y(n5472));
  OAI21X1 g4334(.A0(n5471), .A1(n1825), .B0(n5472), .Y(U2944));
  AOI22X1 g4335(.A0(n5439), .A1(DATAI_4_), .B0(EAX_REG_4__SCAN_IN), .B1(n5440), .Y(n5474));
  OAI21X1 g4336(.A0(n5438), .A1(n1825), .B0(LWORD_REG_4__SCAN_IN), .Y(n5475));
  OAI21X1 g4337(.A0(n5474), .A1(n1825), .B0(n5475), .Y(U2943));
  AOI22X1 g4338(.A0(n5439), .A1(DATAI_3_), .B0(EAX_REG_3__SCAN_IN), .B1(n5440), .Y(n5477));
  OAI21X1 g4339(.A0(n5438), .A1(n1825), .B0(LWORD_REG_3__SCAN_IN), .Y(n5478));
  OAI21X1 g4340(.A0(n5477), .A1(n1825), .B0(n5478), .Y(U2942));
  AOI22X1 g4341(.A0(n5439), .A1(DATAI_2_), .B0(EAX_REG_2__SCAN_IN), .B1(n5440), .Y(n5480));
  OAI21X1 g4342(.A0(n5438), .A1(n1825), .B0(LWORD_REG_2__SCAN_IN), .Y(n5481));
  OAI21X1 g4343(.A0(n5480), .A1(n1825), .B0(n5481), .Y(U2941));
  AOI22X1 g4344(.A0(n5439), .A1(DATAI_1_), .B0(EAX_REG_1__SCAN_IN), .B1(n5440), .Y(n5483));
  OAI21X1 g4345(.A0(n5438), .A1(n1825), .B0(LWORD_REG_1__SCAN_IN), .Y(n5484));
  OAI21X1 g4346(.A0(n5483), .A1(n1825), .B0(n5484), .Y(U2940));
  AOI22X1 g4347(.A0(n5439), .A1(DATAI_0_), .B0(EAX_REG_0__SCAN_IN), .B1(n5440), .Y(n5486));
  OAI21X1 g4348(.A0(n5438), .A1(n1825), .B0(LWORD_REG_0__SCAN_IN), .Y(n5487));
  OAI21X1 g4349(.A0(n5486), .A1(n1825), .B0(n5487), .Y(U2939));
  AOI22X1 g4350(.A0(n5439), .A1(DATAI_14_), .B0(EAX_REG_30__SCAN_IN), .B1(n5440), .Y(n5489));
  OAI21X1 g4351(.A0(n5438), .A1(n1825), .B0(UWORD_REG_14__SCAN_IN), .Y(n5490));
  OAI21X1 g4352(.A0(n5489), .A1(n1825), .B0(n5490), .Y(U2938));
  AOI22X1 g4353(.A0(n5439), .A1(DATAI_13_), .B0(EAX_REG_29__SCAN_IN), .B1(n5440), .Y(n5492));
  OAI21X1 g4354(.A0(n5438), .A1(n1825), .B0(UWORD_REG_13__SCAN_IN), .Y(n5493));
  OAI21X1 g4355(.A0(n5492), .A1(n1825), .B0(n5493), .Y(U2937));
  AOI22X1 g4356(.A0(n5439), .A1(DATAI_12_), .B0(EAX_REG_28__SCAN_IN), .B1(n5440), .Y(n5495));
  OAI21X1 g4357(.A0(n5438), .A1(n1825), .B0(UWORD_REG_12__SCAN_IN), .Y(n5496));
  OAI21X1 g4358(.A0(n5495), .A1(n1825), .B0(n5496), .Y(U2936));
  AOI22X1 g4359(.A0(n5439), .A1(DATAI_11_), .B0(EAX_REG_27__SCAN_IN), .B1(n5440), .Y(n5498));
  OAI21X1 g4360(.A0(n5438), .A1(n1825), .B0(UWORD_REG_11__SCAN_IN), .Y(n5499));
  OAI21X1 g4361(.A0(n5498), .A1(n1825), .B0(n5499), .Y(U2935));
  AOI22X1 g4362(.A0(n5439), .A1(DATAI_10_), .B0(EAX_REG_26__SCAN_IN), .B1(n5440), .Y(n5501));
  OAI21X1 g4363(.A0(n5438), .A1(n1825), .B0(UWORD_REG_10__SCAN_IN), .Y(n5502));
  OAI21X1 g4364(.A0(n5501), .A1(n1825), .B0(n5502), .Y(U2934));
  AOI22X1 g4365(.A0(n5439), .A1(DATAI_9_), .B0(EAX_REG_25__SCAN_IN), .B1(n5440), .Y(n5504));
  OAI21X1 g4366(.A0(n5438), .A1(n1825), .B0(UWORD_REG_9__SCAN_IN), .Y(n5505));
  OAI21X1 g4367(.A0(n5504), .A1(n1825), .B0(n5505), .Y(U2933));
  AOI22X1 g4368(.A0(n5439), .A1(DATAI_8_), .B0(EAX_REG_24__SCAN_IN), .B1(n5440), .Y(n5507));
  OAI21X1 g4369(.A0(n5438), .A1(n1825), .B0(UWORD_REG_8__SCAN_IN), .Y(n5508));
  OAI21X1 g4370(.A0(n5507), .A1(n1825), .B0(n5508), .Y(U2932));
  AOI22X1 g4371(.A0(n5439), .A1(DATAI_7_), .B0(EAX_REG_23__SCAN_IN), .B1(n5440), .Y(n5510));
  OAI21X1 g4372(.A0(n5438), .A1(n1825), .B0(UWORD_REG_7__SCAN_IN), .Y(n5511));
  OAI21X1 g4373(.A0(n5510), .A1(n1825), .B0(n5511), .Y(U2931));
  AOI22X1 g4374(.A0(n5439), .A1(DATAI_6_), .B0(EAX_REG_22__SCAN_IN), .B1(n5440), .Y(n5513));
  OAI21X1 g4375(.A0(n5438), .A1(n1825), .B0(UWORD_REG_6__SCAN_IN), .Y(n5514));
  OAI21X1 g4376(.A0(n5513), .A1(n1825), .B0(n5514), .Y(U2930));
  AOI22X1 g4377(.A0(n5439), .A1(DATAI_5_), .B0(EAX_REG_21__SCAN_IN), .B1(n5440), .Y(n5516));
  OAI21X1 g4378(.A0(n5438), .A1(n1825), .B0(UWORD_REG_5__SCAN_IN), .Y(n5517));
  OAI21X1 g4379(.A0(n5516), .A1(n1825), .B0(n5517), .Y(U2929));
  AOI22X1 g4380(.A0(n5439), .A1(DATAI_4_), .B0(EAX_REG_20__SCAN_IN), .B1(n5440), .Y(n5519));
  OAI21X1 g4381(.A0(n5438), .A1(n1825), .B0(UWORD_REG_4__SCAN_IN), .Y(n5520));
  OAI21X1 g4382(.A0(n5519), .A1(n1825), .B0(n5520), .Y(U2928));
  AOI22X1 g4383(.A0(n5439), .A1(DATAI_3_), .B0(EAX_REG_19__SCAN_IN), .B1(n5440), .Y(n5522));
  OAI21X1 g4384(.A0(n5438), .A1(n1825), .B0(UWORD_REG_3__SCAN_IN), .Y(n5523));
  OAI21X1 g4385(.A0(n5522), .A1(n1825), .B0(n5523), .Y(U2927));
  AOI22X1 g4386(.A0(n5439), .A1(DATAI_2_), .B0(EAX_REG_18__SCAN_IN), .B1(n5440), .Y(n5525));
  OAI21X1 g4387(.A0(n5438), .A1(n1825), .B0(UWORD_REG_2__SCAN_IN), .Y(n5526));
  OAI21X1 g4388(.A0(n5525), .A1(n1825), .B0(n5526), .Y(U2926));
  AOI22X1 g4389(.A0(n5439), .A1(DATAI_1_), .B0(EAX_REG_17__SCAN_IN), .B1(n5440), .Y(n5528));
  OAI21X1 g4390(.A0(n5438), .A1(n1825), .B0(UWORD_REG_1__SCAN_IN), .Y(n5529));
  OAI21X1 g4391(.A0(n5528), .A1(n1825), .B0(n5529), .Y(U2925));
  AOI22X1 g4392(.A0(n5439), .A1(DATAI_0_), .B0(EAX_REG_16__SCAN_IN), .B1(n5440), .Y(n5531));
  OAI21X1 g4393(.A0(n5438), .A1(n1825), .B0(UWORD_REG_0__SCAN_IN), .Y(n5532));
  OAI21X1 g4394(.A0(n5531), .A1(n1825), .B0(n5532), .Y(U2924));
  NOR3X1  g4395(.A(n2103), .B(n1825), .C(n1721), .Y(n5534));
  OAI21X1 g4396(.A0(n5534), .A1(n2003), .B0(n1834), .Y(n5535));
  OAI22X1 g4397(.A0(n2060), .A1(n5535), .B0(n2087), .B1(STATE2_REG_0__SCAN_IN), .Y(n5536));
  INVX1   g4398(.A(n5536), .Y(n5537));
  NOR2X1  g4399(.A(n5537), .B(n1217), .Y(n5538));
  INVX1   g4400(.A(n5538), .Y(n5539));
  NOR2X1  g4401(.A(n5537), .B(STATE2_REG_0__SCAN_IN), .Y(n5540));
  AOI22X1 g4402(.A0(n5537), .A1(DATAO_REG_0__SCAN_IN), .B0(LWORD_REG_0__SCAN_IN), .B1(n5540), .Y(n5541));
  OAI21X1 g4403(.A0(n5539), .A1(n4424), .B0(n5541), .Y(U2923));
  AOI22X1 g4404(.A0(n5537), .A1(DATAO_REG_1__SCAN_IN), .B0(LWORD_REG_1__SCAN_IN), .B1(n5540), .Y(n5543));
  OAI21X1 g4405(.A0(n5539), .A1(n4453), .B0(n5543), .Y(U2922));
  AOI22X1 g4406(.A0(n5537), .A1(DATAO_REG_2__SCAN_IN), .B0(LWORD_REG_2__SCAN_IN), .B1(n5540), .Y(n5545));
  OAI21X1 g4407(.A0(n5539), .A1(n4481), .B0(n5545), .Y(U2921));
  NAND3X1 g4408(.A(n5536), .B(EAX_REG_3__SCAN_IN), .C(STATE2_REG_0__SCAN_IN), .Y(n5547));
  AOI22X1 g4409(.A0(n5537), .A1(DATAO_REG_3__SCAN_IN), .B0(LWORD_REG_3__SCAN_IN), .B1(n5540), .Y(n5548));
  NAND2X1 g4410(.A(n5548), .B(n5547), .Y(U2920));
  AOI22X1 g4411(.A0(n5537), .A1(DATAO_REG_4__SCAN_IN), .B0(LWORD_REG_4__SCAN_IN), .B1(n5540), .Y(n5550));
  OAI21X1 g4412(.A0(n5539), .A1(n4522), .B0(n5550), .Y(U2919));
  NAND3X1 g4413(.A(n5536), .B(EAX_REG_5__SCAN_IN), .C(STATE2_REG_0__SCAN_IN), .Y(n5552));
  AOI22X1 g4414(.A0(n5537), .A1(DATAO_REG_5__SCAN_IN), .B0(LWORD_REG_5__SCAN_IN), .B1(n5540), .Y(n5553));
  NAND2X1 g4415(.A(n5553), .B(n5552), .Y(U2918));
  NAND3X1 g4416(.A(n5536), .B(EAX_REG_6__SCAN_IN), .C(STATE2_REG_0__SCAN_IN), .Y(n5555));
  AOI22X1 g4417(.A0(n5537), .A1(DATAO_REG_6__SCAN_IN), .B0(LWORD_REG_6__SCAN_IN), .B1(n5540), .Y(n5556));
  NAND2X1 g4418(.A(n5556), .B(n5555), .Y(U2917));
  NAND3X1 g4419(.A(n5536), .B(EAX_REG_7__SCAN_IN), .C(STATE2_REG_0__SCAN_IN), .Y(n5558));
  AOI22X1 g4420(.A0(n5537), .A1(DATAO_REG_7__SCAN_IN), .B0(LWORD_REG_7__SCAN_IN), .B1(n5540), .Y(n5559));
  NAND2X1 g4421(.A(n5559), .B(n5558), .Y(U2916));
  NAND3X1 g4422(.A(n5536), .B(EAX_REG_8__SCAN_IN), .C(STATE2_REG_0__SCAN_IN), .Y(n5561));
  AOI22X1 g4423(.A0(n5537), .A1(DATAO_REG_8__SCAN_IN), .B0(LWORD_REG_8__SCAN_IN), .B1(n5540), .Y(n5562));
  NAND2X1 g4424(.A(n5562), .B(n5561), .Y(U2915));
  NAND3X1 g4425(.A(n5536), .B(EAX_REG_9__SCAN_IN), .C(STATE2_REG_0__SCAN_IN), .Y(n5564));
  AOI22X1 g4426(.A0(n5537), .A1(DATAO_REG_9__SCAN_IN), .B0(LWORD_REG_9__SCAN_IN), .B1(n5540), .Y(n5565));
  NAND2X1 g4427(.A(n5565), .B(n5564), .Y(U2914));
  NAND3X1 g4428(.A(n5536), .B(EAX_REG_10__SCAN_IN), .C(STATE2_REG_0__SCAN_IN), .Y(n5567));
  AOI22X1 g4429(.A0(n5537), .A1(DATAO_REG_10__SCAN_IN), .B0(LWORD_REG_10__SCAN_IN), .B1(n5540), .Y(n5568));
  NAND2X1 g4430(.A(n5568), .B(n5567), .Y(U2913));
  NAND3X1 g4431(.A(n5536), .B(EAX_REG_11__SCAN_IN), .C(STATE2_REG_0__SCAN_IN), .Y(n5570));
  AOI22X1 g4432(.A0(n5537), .A1(DATAO_REG_11__SCAN_IN), .B0(LWORD_REG_11__SCAN_IN), .B1(n5540), .Y(n5571));
  NAND2X1 g4433(.A(n5571), .B(n5570), .Y(U2912));
  NAND3X1 g4434(.A(n5536), .B(EAX_REG_12__SCAN_IN), .C(STATE2_REG_0__SCAN_IN), .Y(n5573));
  AOI22X1 g4435(.A0(n5537), .A1(DATAO_REG_12__SCAN_IN), .B0(LWORD_REG_12__SCAN_IN), .B1(n5540), .Y(n5574));
  NAND2X1 g4436(.A(n5574), .B(n5573), .Y(U2911));
  AOI22X1 g4437(.A0(n5537), .A1(DATAO_REG_13__SCAN_IN), .B0(LWORD_REG_13__SCAN_IN), .B1(n5540), .Y(n5576));
  OAI21X1 g4438(.A0(n5539), .A1(n4742), .B0(n5576), .Y(U2910));
  AOI22X1 g4439(.A0(n5537), .A1(DATAO_REG_14__SCAN_IN), .B0(LWORD_REG_14__SCAN_IN), .B1(n5540), .Y(n5578));
  OAI21X1 g4440(.A0(n5539), .A1(n4766), .B0(n5578), .Y(U2909));
  AOI22X1 g4441(.A0(n5537), .A1(DATAO_REG_15__SCAN_IN), .B0(LWORD_REG_15__SCAN_IN), .B1(n5540), .Y(n5580));
  OAI21X1 g4442(.A0(n5539), .A1(n4788), .B0(n5580), .Y(U2908));
  INVX1   g4443(.A(EAX_REG_16__SCAN_IN), .Y(n5582));
  NAND3X1 g4444(.A(n5536), .B(n1447), .C(STATE2_REG_0__SCAN_IN), .Y(n5583));
  AOI22X1 g4445(.A0(n5537), .A1(DATAO_REG_16__SCAN_IN), .B0(UWORD_REG_0__SCAN_IN), .B1(n5540), .Y(n5584));
  OAI21X1 g4446(.A0(n5583), .A1(n5582), .B0(n5584), .Y(U2907));
  INVX1   g4447(.A(EAX_REG_17__SCAN_IN), .Y(n5586));
  AOI22X1 g4448(.A0(n5537), .A1(DATAO_REG_17__SCAN_IN), .B0(UWORD_REG_1__SCAN_IN), .B1(n5540), .Y(n5587));
  OAI21X1 g4449(.A0(n5583), .A1(n5586), .B0(n5587), .Y(U2906));
  INVX1   g4450(.A(EAX_REG_18__SCAN_IN), .Y(n5589));
  AOI22X1 g4451(.A0(n5537), .A1(DATAO_REG_18__SCAN_IN), .B0(UWORD_REG_2__SCAN_IN), .B1(n5540), .Y(n5590));
  OAI21X1 g4452(.A0(n5583), .A1(n5589), .B0(n5590), .Y(U2905));
  INVX1   g4453(.A(EAX_REG_19__SCAN_IN), .Y(n5592));
  AOI22X1 g4454(.A0(n5537), .A1(DATAO_REG_19__SCAN_IN), .B0(UWORD_REG_3__SCAN_IN), .B1(n5540), .Y(n5593));
  OAI21X1 g4455(.A0(n5583), .A1(n5592), .B0(n5593), .Y(U2904));
  INVX1   g4456(.A(EAX_REG_20__SCAN_IN), .Y(n5595));
  AOI22X1 g4457(.A0(n5537), .A1(DATAO_REG_20__SCAN_IN), .B0(UWORD_REG_4__SCAN_IN), .B1(n5540), .Y(n5596));
  OAI21X1 g4458(.A0(n5583), .A1(n5595), .B0(n5596), .Y(U2903));
  INVX1   g4459(.A(EAX_REG_21__SCAN_IN), .Y(n5598));
  AOI22X1 g4460(.A0(n5537), .A1(DATAO_REG_21__SCAN_IN), .B0(UWORD_REG_5__SCAN_IN), .B1(n5540), .Y(n5599));
  OAI21X1 g4461(.A0(n5583), .A1(n5598), .B0(n5599), .Y(U2902));
  INVX1   g4462(.A(EAX_REG_22__SCAN_IN), .Y(n5601));
  AOI22X1 g4463(.A0(n5537), .A1(DATAO_REG_22__SCAN_IN), .B0(UWORD_REG_6__SCAN_IN), .B1(n5540), .Y(n5602));
  OAI21X1 g4464(.A0(n5583), .A1(n5601), .B0(n5602), .Y(U2901));
  INVX1   g4465(.A(EAX_REG_23__SCAN_IN), .Y(n5604));
  AOI22X1 g4466(.A0(n5537), .A1(DATAO_REG_23__SCAN_IN), .B0(UWORD_REG_7__SCAN_IN), .B1(n5540), .Y(n5605));
  OAI21X1 g4467(.A0(n5583), .A1(n5604), .B0(n5605), .Y(U2900));
  AOI22X1 g4468(.A0(n5537), .A1(DATAO_REG_24__SCAN_IN), .B0(UWORD_REG_8__SCAN_IN), .B1(n5540), .Y(n5607));
  OAI21X1 g4469(.A0(n5583), .A1(n5165), .B0(n5607), .Y(U2899));
  AOI22X1 g4470(.A0(n5537), .A1(DATAO_REG_25__SCAN_IN), .B0(UWORD_REG_9__SCAN_IN), .B1(n5540), .Y(n5609));
  OAI21X1 g4471(.A0(n5583), .A1(n5200), .B0(n5609), .Y(U2898));
  AOI22X1 g4472(.A0(n5537), .A1(DATAO_REG_26__SCAN_IN), .B0(UWORD_REG_10__SCAN_IN), .B1(n5540), .Y(n5611));
  OAI21X1 g4473(.A0(n5583), .A1(n5240), .B0(n5611), .Y(U2897));
  INVX1   g4474(.A(EAX_REG_27__SCAN_IN), .Y(n5613));
  AOI22X1 g4475(.A0(n5537), .A1(DATAO_REG_27__SCAN_IN), .B0(UWORD_REG_11__SCAN_IN), .B1(n5540), .Y(n5614));
  OAI21X1 g4476(.A0(n5583), .A1(n5613), .B0(n5614), .Y(U2896));
  AOI22X1 g4477(.A0(n5537), .A1(DATAO_REG_28__SCAN_IN), .B0(UWORD_REG_12__SCAN_IN), .B1(n5540), .Y(n5616));
  OAI21X1 g4478(.A0(n5583), .A1(n5310), .B0(n5616), .Y(U2895));
  AOI22X1 g4479(.A0(n5537), .A1(DATAO_REG_29__SCAN_IN), .B0(UWORD_REG_13__SCAN_IN), .B1(n5540), .Y(n5618));
  OAI21X1 g4480(.A0(n5583), .A1(n5361), .B0(n5618), .Y(U2894));
  INVX1   g4481(.A(EAX_REG_30__SCAN_IN), .Y(n5620));
  AOI22X1 g4482(.A0(n5537), .A1(DATAO_REG_30__SCAN_IN), .B0(UWORD_REG_14__SCAN_IN), .B1(n5540), .Y(n5621));
  OAI21X1 g4483(.A0(n5583), .A1(n5620), .B0(n5621), .Y(U2893));
  INVX1   g4484(.A(DATAO_REG_31__SCAN_IN), .Y(n5623));
  NOR2X1  g4485(.A(n5536), .B(n5623), .Y(U2892));
  NOR4X1  g4486(.A(n2032), .B(n1448), .C(n1217), .D(n1825), .Y(n5625));
  NOR3X1  g4487(.A(n1734), .B(n2037), .C(n1872), .Y(n5626));
  OAI21X1 g4488(.A0(n5626), .A1(n5625), .B0(n1113), .Y(n5627));
  NOR4X1  g4489(.A(n1639), .B(n1655), .C(n1872), .D(n1677), .Y(n5628));
  NOR3X1  g4490(.A(n1777), .B(n1816), .C(n1872), .Y(n5629));
  AOI21X1 g4491(.A0(n5628), .A1(n1536), .B0(n5629), .Y(n5630));
  AOI21X1 g4492(.A0(n5630), .A1(n5627), .B0(n1950), .Y(n5631));
  OAI21X1 g4493(.A0(n1736), .A1(n1700), .B0(n5631), .Y(n5632));
  INVX1   g4494(.A(n5631), .Y(n5633));
  NOR3X1  g4495(.A(n5633), .B(n1736), .C(n1700), .Y(n5634));
  AOI22X1 g4496(.A0(n5633), .A1(EAX_REG_0__SCAN_IN), .B0(DATAI_0_), .B1(n5634), .Y(n5635));
  OAI21X1 g4497(.A0(n5632), .A1(n4434), .B0(n5635), .Y(U2891));
  AOI22X1 g4498(.A0(n5633), .A1(EAX_REG_1__SCAN_IN), .B0(DATAI_1_), .B1(n5634), .Y(n5637));
  OAI21X1 g4499(.A0(n5632), .A1(n4470), .B0(n5637), .Y(U2890));
  AOI22X1 g4500(.A0(n5633), .A1(EAX_REG_2__SCAN_IN), .B0(DATAI_2_), .B1(n5634), .Y(n5639));
  OAI21X1 g4501(.A0(n5632), .A1(n4497), .B0(n5639), .Y(U2889));
  INVX1   g4502(.A(n4515), .Y(n5641));
  AOI22X1 g4503(.A0(n5633), .A1(EAX_REG_3__SCAN_IN), .B0(DATAI_3_), .B1(n5634), .Y(n5642));
  OAI21X1 g4504(.A0(n5632), .A1(n5641), .B0(n5642), .Y(U2888));
  AOI22X1 g4505(.A0(n5633), .A1(EAX_REG_4__SCAN_IN), .B0(DATAI_4_), .B1(n5634), .Y(n5644));
  OAI21X1 g4506(.A0(n5632), .A1(n4539), .B0(n5644), .Y(U2887));
  AOI22X1 g4507(.A0(n5633), .A1(EAX_REG_5__SCAN_IN), .B0(DATAI_5_), .B1(n5634), .Y(n5646));
  OAI21X1 g4508(.A0(n5632), .A1(n4562), .B0(n5646), .Y(U2886));
  INVX1   g4509(.A(n4582), .Y(n5648));
  AOI22X1 g4510(.A0(n5633), .A1(EAX_REG_6__SCAN_IN), .B0(DATAI_6_), .B1(n5634), .Y(n5649));
  OAI21X1 g4511(.A0(n5632), .A1(n5648), .B0(n5649), .Y(U2885));
  AOI22X1 g4512(.A0(n5633), .A1(EAX_REG_7__SCAN_IN), .B0(DATAI_7_), .B1(n5634), .Y(n5651));
  OAI21X1 g4513(.A0(n5632), .A1(n4606), .B0(n5651), .Y(U2884));
  INVX1   g4514(.A(n4632), .Y(n5653));
  AOI22X1 g4515(.A0(n5633), .A1(EAX_REG_8__SCAN_IN), .B0(DATAI_8_), .B1(n5634), .Y(n5654));
  OAI21X1 g4516(.A0(n5632), .A1(n5653), .B0(n5654), .Y(U2883));
  AOI22X1 g4517(.A0(n5633), .A1(EAX_REG_9__SCAN_IN), .B0(DATAI_9_), .B1(n5634), .Y(n5656));
  OAI21X1 g4518(.A0(n5632), .A1(n4653), .B0(n5656), .Y(U2882));
  AOI22X1 g4519(.A0(n5633), .A1(EAX_REG_10__SCAN_IN), .B0(DATAI_10_), .B1(n5634), .Y(n5658));
  OAI21X1 g4520(.A0(n5632), .A1(n4680), .B0(n5658), .Y(U2881));
  INVX1   g4521(.A(n4702), .Y(n5660));
  AOI22X1 g4522(.A0(n5633), .A1(EAX_REG_11__SCAN_IN), .B0(DATAI_11_), .B1(n5634), .Y(n5661));
  OAI21X1 g4523(.A0(n5632), .A1(n5660), .B0(n5661), .Y(U2880));
  AOI22X1 g4524(.A0(n5633), .A1(EAX_REG_12__SCAN_IN), .B0(DATAI_12_), .B1(n5634), .Y(n5663));
  OAI21X1 g4525(.A0(n5632), .A1(n4724), .B0(n5663), .Y(U2879));
  AOI22X1 g4526(.A0(n5633), .A1(EAX_REG_13__SCAN_IN), .B0(DATAI_13_), .B1(n5634), .Y(n5665));
  OAI21X1 g4527(.A0(n5632), .A1(n4753), .B0(n5665), .Y(U2878));
  NOR2X1  g4528(.A(n4772), .B(n4762), .Y(n5667));
  AOI21X1 g4529(.A0(n4762), .A1(n4772), .B0(n5667), .Y(n5668));
  AOI22X1 g4530(.A0(n5633), .A1(EAX_REG_14__SCAN_IN), .B0(DATAI_14_), .B1(n5634), .Y(n5669));
  OAI21X1 g4531(.A0(n5632), .A1(n5668), .B0(n5669), .Y(U2877));
  OAI21X1 g4532(.A0(n4775), .A1(n4762), .B0(n4797), .Y(n5671));
  OAI21X1 g4533(.A0(n4774), .A1(n4783), .B0(n4800), .Y(n5672));
  NAND2X1 g4534(.A(n5672), .B(n5671), .Y(n5673));
  AOI22X1 g4535(.A0(n5633), .A1(EAX_REG_15__SCAN_IN), .B0(DATAI_15_), .B1(n5634), .Y(n5674));
  OAI21X1 g4536(.A0(n5632), .A1(n5673), .B0(n5674), .Y(U2876));
  INVX1   g4537(.A(n4876), .Y(n5676));
  NOR3X1  g4538(.A(n5633), .B(n1700), .C(n1394), .Y(n5677));
  NOR2X1  g4539(.A(n5633), .B(n1804), .Y(n5678));
  INVX1   g4540(.A(n5678), .Y(n5679));
  OAI22X1 g4541(.A0(n5631), .A1(n5582), .B0(n2342), .B1(n5679), .Y(n5680));
  AOI21X1 g4542(.A0(n5677), .A1(DATAI_0_), .B0(n5680), .Y(n5681));
  OAI21X1 g4543(.A0(n5632), .A1(n5676), .B0(n5681), .Y(U2875));
  INVX1   g4544(.A(n4905), .Y(n5683));
  OAI22X1 g4545(.A0(n5631), .A1(n5586), .B0(n2334), .B1(n5679), .Y(n5684));
  AOI21X1 g4546(.A0(n5677), .A1(DATAI_1_), .B0(n5684), .Y(n5685));
  OAI21X1 g4547(.A0(n5632), .A1(n5683), .B0(n5685), .Y(U2874));
  OAI22X1 g4548(.A0(n5631), .A1(n5589), .B0(n2326), .B1(n5679), .Y(n5687));
  AOI21X1 g4549(.A0(n5677), .A1(DATAI_2_), .B0(n5687), .Y(n5688));
  OAI21X1 g4550(.A0(n5632), .A1(n4934), .B0(n5688), .Y(U2873));
  INVX1   g4551(.A(n4969), .Y(n5690));
  OAI22X1 g4552(.A0(n5631), .A1(n5592), .B0(n2318), .B1(n5679), .Y(n5691));
  AOI21X1 g4553(.A0(n5677), .A1(DATAI_3_), .B0(n5691), .Y(n5692));
  OAI21X1 g4554(.A0(n5632), .A1(n5690), .B0(n5692), .Y(U2872));
  NOR2X1  g4555(.A(n5005), .B(n5001), .Y(n5694));
  OAI22X1 g4556(.A0(n5631), .A1(n5595), .B0(n2310), .B1(n5679), .Y(n5695));
  AOI21X1 g4557(.A0(n5677), .A1(DATAI_4_), .B0(n5695), .Y(n5696));
  OAI21X1 g4558(.A0(n5632), .A1(n5694), .B0(n5696), .Y(U2871));
  NAND2X1 g4559(.A(n5041), .B(n5038), .Y(n5698));
  OAI21X1 g4560(.A0(n5036), .A1(n5014), .B0(n5698), .Y(n5699));
  OAI22X1 g4561(.A0(n5631), .A1(n5598), .B0(n2302), .B1(n5679), .Y(n5700));
  AOI21X1 g4562(.A0(n5677), .A1(DATAI_5_), .B0(n5700), .Y(n5701));
  OAI21X1 g4563(.A0(n5632), .A1(n5699), .B0(n5701), .Y(U2870));
  XOR2X1  g4564(.A(n5073), .B(n5068), .Y(n5703));
  OAI22X1 g4565(.A0(n5631), .A1(n5601), .B0(n2294), .B1(n5679), .Y(n5704));
  AOI21X1 g4566(.A0(n5677), .A1(DATAI_6_), .B0(n5704), .Y(n5705));
  OAI21X1 g4567(.A0(n5632), .A1(n5703), .B0(n5705), .Y(U2869));
  INVX1   g4568(.A(n5140), .Y(n5707));
  OAI22X1 g4569(.A0(n5631), .A1(n5604), .B0(n2285), .B1(n5679), .Y(n5708));
  AOI21X1 g4570(.A0(n5677), .A1(DATAI_7_), .B0(n5708), .Y(n5709));
  OAI21X1 g4571(.A0(n5632), .A1(n5707), .B0(n5709), .Y(U2868));
  XOR2X1  g4572(.A(n5175), .B(n5171), .Y(n5711));
  NAND3X1 g4573(.A(n5631), .B(n1919), .C(DATAI_24_), .Y(n5712));
  OAI21X1 g4574(.A0(n5631), .A1(n5165), .B0(n5712), .Y(n5713));
  AOI21X1 g4575(.A0(n5677), .A1(DATAI_8_), .B0(n5713), .Y(n5714));
  OAI21X1 g4576(.A0(n5632), .A1(n5711), .B0(n5714), .Y(U2867));
  INVX1   g4577(.A(n5217), .Y(n5716));
  NAND3X1 g4578(.A(n5631), .B(n1919), .C(DATAI_25_), .Y(n5717));
  OAI21X1 g4579(.A0(n5631), .A1(n5200), .B0(n5717), .Y(n5718));
  AOI21X1 g4580(.A0(n5677), .A1(DATAI_9_), .B0(n5718), .Y(n5719));
  OAI21X1 g4581(.A0(n5632), .A1(n5716), .B0(n5719), .Y(U2866));
  NAND3X1 g4582(.A(n5631), .B(n1919), .C(DATAI_26_), .Y(n5721));
  OAI21X1 g4583(.A0(n5631), .A1(n5240), .B0(n5721), .Y(n5722));
  AOI21X1 g4584(.A0(n5677), .A1(DATAI_10_), .B0(n5722), .Y(n5723));
  OAI21X1 g4585(.A0(n5632), .A1(n5251), .B0(n5723), .Y(U2865));
  XOR2X1  g4586(.A(n5284), .B(n5280), .Y(n5725));
  NAND3X1 g4587(.A(n5631), .B(n1919), .C(DATAI_27_), .Y(n5726));
  OAI21X1 g4588(.A0(n5631), .A1(n5613), .B0(n5726), .Y(n5727));
  AOI21X1 g4589(.A0(n5677), .A1(DATAI_11_), .B0(n5727), .Y(n5728));
  OAI21X1 g4590(.A0(n5632), .A1(n5725), .B0(n5728), .Y(U2864));
  INVX1   g4591(.A(n5318), .Y(n5730));
  XOR2X1  g4592(.A(n5337), .B(n5730), .Y(n5731));
  NAND3X1 g4593(.A(n5631), .B(n1919), .C(DATAI_28_), .Y(n5732));
  OAI21X1 g4594(.A0(n5631), .A1(n5310), .B0(n5732), .Y(n5733));
  AOI21X1 g4595(.A0(n5677), .A1(DATAI_12_), .B0(n5733), .Y(n5734));
  OAI21X1 g4596(.A0(n5632), .A1(n5731), .B0(n5734), .Y(U2863));
  INVX1   g4597(.A(n5367), .Y(n5736));
  XOR2X1  g4598(.A(n5371), .B(n5736), .Y(n5737));
  NAND3X1 g4599(.A(n5631), .B(n1919), .C(DATAI_29_), .Y(n5738));
  OAI21X1 g4600(.A0(n5631), .A1(n5361), .B0(n5738), .Y(n5739));
  AOI21X1 g4601(.A0(n5677), .A1(DATAI_13_), .B0(n5739), .Y(n5740));
  OAI21X1 g4602(.A0(n5632), .A1(n5737), .B0(n5740), .Y(U2862));
  INVX1   g4603(.A(n5399), .Y(n5742));
  XOR2X1  g4604(.A(n5407), .B(n5742), .Y(n5743));
  NAND3X1 g4605(.A(n5631), .B(n1919), .C(DATAI_30_), .Y(n5744));
  OAI21X1 g4606(.A0(n5631), .A1(n5620), .B0(n5744), .Y(n5745));
  AOI21X1 g4607(.A0(n5677), .A1(DATAI_14_), .B0(n5745), .Y(n5746));
  OAI21X1 g4608(.A0(n5632), .A1(n5743), .B0(n5746), .Y(U2861));
  INVX1   g4609(.A(n5430), .Y(n5748));
  XOR2X1  g4610(.A(n5748), .B(n5422), .Y(n5749));
  NAND2X1 g4611(.A(n5631), .B(n1700), .Y(n5750));
  AOI22X1 g4612(.A0(n5633), .A1(EAX_REG_31__SCAN_IN), .B0(DATAI_31_), .B1(n5678), .Y(n5751));
  OAI21X1 g4613(.A0(n5750), .A1(n5749), .B0(n5751), .Y(U2860));
  NAND2X1 g4614(.A(n1720), .B(STATE2_REG_0__SCAN_IN), .Y(n5753));
  NOR4X1  g4615(.A(n1592), .B(n1464), .C(n1282), .D(n5753), .Y(n5754));
  NOR3X1  g4616(.A(n1685), .B(n1536), .C(n1217), .Y(n5755));
  AOI21X1 g4617(.A0(n5754), .A1(n1778), .B0(n5755), .Y(n5756));
  NOR2X1  g4618(.A(n5756), .B(n1950), .Y(n5757));
  NAND2X1 g4619(.A(n5757), .B(n1615), .Y(n5758));
  INVX1   g4620(.A(n5757), .Y(n5759));
  NOR3X1  g4621(.A(n5756), .B(n1950), .C(n1615), .Y(n5760));
  AOI22X1 g4622(.A0(n5759), .A1(EBX_REG_0__SCAN_IN), .B0(n3276), .B1(n5760), .Y(n5761));
  OAI21X1 g4623(.A0(n5758), .A1(n4434), .B0(n5761), .Y(U2859));
  AOI22X1 g4624(.A0(n5759), .A1(EBX_REG_1__SCAN_IN), .B0(n3287), .B1(n5760), .Y(n5763));
  OAI21X1 g4625(.A0(n5758), .A1(n4470), .B0(n5763), .Y(U2858));
  AOI22X1 g4626(.A0(n5759), .A1(EBX_REG_2__SCAN_IN), .B0(n3329), .B1(n5760), .Y(n5765));
  OAI21X1 g4627(.A0(n5758), .A1(n4497), .B0(n5765), .Y(U2857));
  INVX1   g4628(.A(n3352), .Y(n5767));
  AOI22X1 g4629(.A0(n5759), .A1(EBX_REG_3__SCAN_IN), .B0(n5767), .B1(n5760), .Y(n5768));
  OAI21X1 g4630(.A0(n5758), .A1(n5641), .B0(n5768), .Y(U2856));
  INVX1   g4631(.A(n3414), .Y(n5770));
  AOI22X1 g4632(.A0(n5759), .A1(EBX_REG_4__SCAN_IN), .B0(n5770), .B1(n5760), .Y(n5771));
  OAI21X1 g4633(.A0(n5758), .A1(n4539), .B0(n5771), .Y(U2855));
  INVX1   g4634(.A(n3470), .Y(n5773));
  AOI22X1 g4635(.A0(n5759), .A1(EBX_REG_5__SCAN_IN), .B0(n5773), .B1(n5760), .Y(n5774));
  OAI21X1 g4636(.A0(n5758), .A1(n4562), .B0(n5774), .Y(U2854));
  INVX1   g4637(.A(n3533), .Y(n5776));
  AOI22X1 g4638(.A0(n5759), .A1(EBX_REG_6__SCAN_IN), .B0(n5776), .B1(n5760), .Y(n5777));
  OAI21X1 g4639(.A0(n5758), .A1(n5648), .B0(n5777), .Y(U2853));
  INVX1   g4640(.A(n3582), .Y(n5779));
  AOI22X1 g4641(.A0(n5759), .A1(EBX_REG_7__SCAN_IN), .B0(n5779), .B1(n5760), .Y(n5780));
  OAI21X1 g4642(.A0(n5758), .A1(n4606), .B0(n5780), .Y(U2852));
  INVX1   g4643(.A(n3667), .Y(n5782));
  AOI22X1 g4644(.A0(n5759), .A1(EBX_REG_8__SCAN_IN), .B0(n5782), .B1(n5760), .Y(n5783));
  OAI21X1 g4645(.A0(n5758), .A1(n5653), .B0(n5783), .Y(U2851));
  INVX1   g4646(.A(n3715), .Y(n5785));
  AOI22X1 g4647(.A0(n5759), .A1(EBX_REG_9__SCAN_IN), .B0(n5785), .B1(n5760), .Y(n5786));
  OAI21X1 g4648(.A0(n5758), .A1(n4653), .B0(n5786), .Y(U2850));
  INVX1   g4649(.A(n3756), .Y(n5788));
  AOI22X1 g4650(.A0(n5759), .A1(EBX_REG_10__SCAN_IN), .B0(n5788), .B1(n5760), .Y(n5789));
  OAI21X1 g4651(.A0(n5758), .A1(n4680), .B0(n5789), .Y(U2849));
  INVX1   g4652(.A(n3796), .Y(n5791));
  AOI22X1 g4653(.A0(n5759), .A1(EBX_REG_11__SCAN_IN), .B0(n5791), .B1(n5760), .Y(n5792));
  OAI21X1 g4654(.A0(n5758), .A1(n5660), .B0(n5792), .Y(U2848));
  INVX1   g4655(.A(n3855), .Y(n5794));
  AOI22X1 g4656(.A0(n5759), .A1(EBX_REG_12__SCAN_IN), .B0(n5794), .B1(n5760), .Y(n5795));
  OAI21X1 g4657(.A0(n5758), .A1(n4724), .B0(n5795), .Y(U2847));
  INVX1   g4658(.A(n3893), .Y(n5797));
  AOI22X1 g4659(.A0(n5759), .A1(EBX_REG_13__SCAN_IN), .B0(n5797), .B1(n5760), .Y(n5798));
  OAI21X1 g4660(.A0(n5758), .A1(n4753), .B0(n5798), .Y(U2846));
  INVX1   g4661(.A(n3932), .Y(n5800));
  AOI22X1 g4662(.A0(n5759), .A1(EBX_REG_14__SCAN_IN), .B0(n5800), .B1(n5760), .Y(n5801));
  OAI21X1 g4663(.A0(n5758), .A1(n5668), .B0(n5801), .Y(U2845));
  INVX1   g4664(.A(n3975), .Y(n5803));
  AOI22X1 g4665(.A0(n5759), .A1(EBX_REG_15__SCAN_IN), .B0(n5803), .B1(n5760), .Y(n5804));
  OAI21X1 g4666(.A0(n5758), .A1(n5673), .B0(n5804), .Y(U2844));
  INVX1   g4667(.A(n4011), .Y(n5806));
  AOI22X1 g4668(.A0(n5759), .A1(EBX_REG_16__SCAN_IN), .B0(n5806), .B1(n5760), .Y(n5807));
  OAI21X1 g4669(.A0(n5758), .A1(n5676), .B0(n5807), .Y(U2843));
  INVX1   g4670(.A(n4035), .Y(n5809));
  AOI22X1 g4671(.A0(n5759), .A1(EBX_REG_17__SCAN_IN), .B0(n5809), .B1(n5760), .Y(n5810));
  OAI21X1 g4672(.A0(n5758), .A1(n5683), .B0(n5810), .Y(U2842));
  INVX1   g4673(.A(n4069), .Y(n5812));
  AOI22X1 g4674(.A0(n5759), .A1(EBX_REG_18__SCAN_IN), .B0(n5812), .B1(n5760), .Y(n5813));
  OAI21X1 g4675(.A0(n5758), .A1(n4934), .B0(n5813), .Y(U2841));
  INVX1   g4676(.A(n4096), .Y(n5815));
  AOI22X1 g4677(.A0(n5759), .A1(EBX_REG_19__SCAN_IN), .B0(n5815), .B1(n5760), .Y(n5816));
  OAI21X1 g4678(.A0(n5758), .A1(n5690), .B0(n5816), .Y(U2840));
  AOI22X1 g4679(.A0(n5759), .A1(EBX_REG_20__SCAN_IN), .B0(n4126), .B1(n5760), .Y(n5818));
  OAI21X1 g4680(.A0(n5758), .A1(n5694), .B0(n5818), .Y(U2839));
  INVX1   g4681(.A(n4148), .Y(n5820));
  AOI22X1 g4682(.A0(n5759), .A1(EBX_REG_21__SCAN_IN), .B0(n5820), .B1(n5760), .Y(n5821));
  OAI21X1 g4683(.A0(n5758), .A1(n5699), .B0(n5821), .Y(U2838));
  INVX1   g4684(.A(n4176), .Y(n5823));
  AOI22X1 g4685(.A0(n5759), .A1(EBX_REG_22__SCAN_IN), .B0(n5823), .B1(n5760), .Y(n5824));
  OAI21X1 g4686(.A0(n5758), .A1(n5703), .B0(n5824), .Y(U2837));
  INVX1   g4687(.A(n4202), .Y(n5826));
  AOI22X1 g4688(.A0(n5759), .A1(EBX_REG_23__SCAN_IN), .B0(n5826), .B1(n5760), .Y(n5827));
  OAI21X1 g4689(.A0(n5758), .A1(n5707), .B0(n5827), .Y(U2836));
  INVX1   g4690(.A(n4227), .Y(n5829));
  AOI22X1 g4691(.A0(n5759), .A1(EBX_REG_24__SCAN_IN), .B0(n5829), .B1(n5760), .Y(n5830));
  OAI21X1 g4692(.A0(n5758), .A1(n5711), .B0(n5830), .Y(U2835));
  AOI22X1 g4693(.A0(n5759), .A1(EBX_REG_25__SCAN_IN), .B0(n4254), .B1(n5760), .Y(n5832));
  OAI21X1 g4694(.A0(n5758), .A1(n5716), .B0(n5832), .Y(U2834));
  INVX1   g4695(.A(n4282), .Y(n5834));
  AOI22X1 g4696(.A0(n5759), .A1(EBX_REG_26__SCAN_IN), .B0(n5834), .B1(n5760), .Y(n5835));
  OAI21X1 g4697(.A0(n5758), .A1(n5251), .B0(n5835), .Y(U2833));
  AOI22X1 g4698(.A0(n5759), .A1(EBX_REG_27__SCAN_IN), .B0(n4306), .B1(n5760), .Y(n5837));
  OAI21X1 g4699(.A0(n5758), .A1(n5725), .B0(n5837), .Y(U2832));
  INVX1   g4700(.A(n5760), .Y(n5839));
  NOR2X1  g4701(.A(n5839), .B(n4330), .Y(n5840));
  AOI21X1 g4702(.A0(n5759), .A1(EBX_REG_28__SCAN_IN), .B0(n5840), .Y(n5841));
  OAI21X1 g4703(.A0(n5758), .A1(n5731), .B0(n5841), .Y(U2831));
  AOI22X1 g4704(.A0(n5759), .A1(EBX_REG_29__SCAN_IN), .B0(n4356), .B1(n5760), .Y(n5843));
  OAI21X1 g4705(.A0(n5758), .A1(n5737), .B0(n5843), .Y(U2830));
  NOR2X1  g4706(.A(n5839), .B(n4382), .Y(n5845));
  AOI21X1 g4707(.A0(n5759), .A1(EBX_REG_30__SCAN_IN), .B0(n5845), .Y(n5846));
  OAI21X1 g4708(.A0(n5758), .A1(n5743), .B0(n5846), .Y(U2829));
  INVX1   g4709(.A(EBX_REG_31__SCAN_IN), .Y(n5848));
  OAI22X1 g4710(.A0(n5757), .A1(n5848), .B0(n4405), .B1(n5839), .Y(U2828));
  NOR3X1  g4711(.A(n2103), .B(n2054), .C(n1825), .Y(n5850));
  AOI22X1 g4712(.A0(n1890), .A1(n1733), .B0(n1536), .B1(n2003), .Y(n5851));
  INVX1   g4713(.A(n5851), .Y(n5852));
  OAI21X1 g4714(.A0(n5852), .A1(n5850), .B0(n1834), .Y(n5853));
  NOR3X1  g4715(.A(n3239), .B(n2105), .C(n2082), .Y(n5854));
  NAND2X1 g4716(.A(n5854), .B(n5853), .Y(n5855));
  NAND3X1 g4717(.A(n5855), .B(n1829), .C(STATE2_REG_2__SCAN_IN), .Y(n5856));
  NOR2X1  g4718(.A(n5856), .B(n2061), .Y(n5857));
  NAND3X1 g4719(.A(n5855), .B(n1867), .C(STATE2_REG_2__SCAN_IN), .Y(n5858));
  AOI21X1 g4720(.A0(n2061), .A1(n2041), .B0(n5858), .Y(n5859));
  AOI21X1 g4721(.A0(n5857), .A1(n5848), .B0(n5859), .Y(n5860));
  INVX1   g4722(.A(n5860), .Y(n5861));
  NAND2X1 g4723(.A(n5861), .B(EBX_REG_0__SCAN_IN), .Y(n5862));
  NAND4X1 g4724(.A(n2041), .B(n1867), .C(STATE2_REG_2__SCAN_IN), .D(n5855), .Y(n5863));
  AOI21X1 g4725(.A0(n5863), .A1(n5856), .B0(n2062), .Y(n5864));
  NOR3X1  g4726(.A(n5856), .B(n2061), .C(n5848), .Y(n5865));
  NAND2X1 g4727(.A(n5865), .B(n3276), .Y(n5866));
  INVX1   g4728(.A(n4434), .Y(n5867));
  AOI22X1 g4729(.A0(n1826), .A1(STATE2_REG_2__SCAN_IN), .B0(STATE2_REG_1__SCAN_IN), .B1(n5425), .Y(n5868));
  AOI21X1 g4730(.A0(n5854), .A1(n5853), .B0(n5868), .Y(n5869));
  NAND2X1 g4731(.A(n5869), .B(n5867), .Y(n5870));
  INVX1   g4732(.A(n5855), .Y(n5871));
  NAND3X1 g4733(.A(n5855), .B(n5424), .C(STATE2_REG_1__SCAN_IN), .Y(n5872));
  INVX1   g4734(.A(n5872), .Y(n5873));
  AOI22X1 g4735(.A0(n5871), .A1(REIP_REG_0__SCAN_IN), .B0(PHYADDRPOINTER_REG_0__SCAN_IN), .B1(n5873), .Y(n5874));
  AOI21X1 g4736(.A0(n5854), .A1(n5853), .B0(n1216), .Y(n5875));
  NOR4X1  g4737(.A(n1464), .B(n1447), .C(n1833), .D(n5871), .Y(n5876));
  AOI22X1 g4738(.A0(n5875), .A1(PHYADDRPOINTER_REG_0__SCAN_IN), .B0(n2185), .B1(n5876), .Y(n5877));
  NAND4X1 g4739(.A(n5874), .B(n5870), .C(n5866), .D(n5877), .Y(n5878));
  AOI21X1 g4740(.A0(n5864), .A1(REIP_REG_0__SCAN_IN), .B0(n5878), .Y(n5879));
  NAND2X1 g4741(.A(n5879), .B(n5862), .Y(U2827));
  NAND2X1 g4742(.A(n5861), .B(EBX_REG_1__SCAN_IN), .Y(n5881));
  NAND2X1 g4743(.A(n5864), .B(n1109), .Y(n5882));
  NAND2X1 g4744(.A(n5865), .B(n3287), .Y(n5883));
  INVX1   g4745(.A(n5869), .Y(n5884));
  NOR2X1  g4746(.A(n5884), .B(n4470), .Y(n5885));
  OAI22X1 g4747(.A0(n5855), .A1(n1109), .B0(PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n5872), .Y(n5886));
  INVX1   g4748(.A(n5875), .Y(n5887));
  OAI21X1 g4749(.A0(n1936), .A1(n1932), .B0(n5876), .Y(n5888));
  OAI21X1 g4750(.A0(n5887), .A1(n4454), .B0(n5888), .Y(n5889));
  NOR3X1  g4751(.A(n5889), .B(n5886), .C(n5885), .Y(n5890));
  NAND4X1 g4752(.A(n5883), .B(n5882), .C(n5881), .D(n5890), .Y(U2826));
  NAND2X1 g4753(.A(n5861), .B(EBX_REG_2__SCAN_IN), .Y(n5892));
  NAND2X1 g4754(.A(n5869), .B(n4496), .Y(n5893));
  XOR2X1  g4755(.A(REIP_REG_2__SCAN_IN), .B(REIP_REG_1__SCAN_IN), .Y(n5894));
  NAND2X1 g4756(.A(n5865), .B(n3329), .Y(n5895));
  AOI22X1 g4757(.A0(n5871), .A1(REIP_REG_2__SCAN_IN), .B0(n4483), .B1(n5873), .Y(n5896));
  AOI22X1 g4758(.A0(n5875), .A1(PHYADDRPOINTER_REG_2__SCAN_IN), .B0(n2522), .B1(n5876), .Y(n5897));
  NAND3X1 g4759(.A(n5897), .B(n5896), .C(n5895), .Y(n5898));
  AOI21X1 g4760(.A0(n5894), .A1(n5864), .B0(n5898), .Y(n5899));
  NAND3X1 g4761(.A(n5899), .B(n5893), .C(n5892), .Y(U2825));
  NAND2X1 g4762(.A(REIP_REG_2__SCAN_IN), .B(REIP_REG_1__SCAN_IN), .Y(n5901));
  XOR2X1  g4763(.A(n5901), .B(n1103), .Y(n5902));
  NAND2X1 g4764(.A(n5902), .B(n5864), .Y(n5903));
  NAND2X1 g4765(.A(n5865), .B(n5767), .Y(n5904));
  AOI22X1 g4766(.A0(n5871), .A1(REIP_REG_3__SCAN_IN), .B0(n4508), .B1(n5873), .Y(n5905));
  AOI22X1 g4767(.A0(n5875), .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .B0(n1988), .B1(n5876), .Y(n5906));
  NAND4X1 g4768(.A(n5905), .B(n5904), .C(n5903), .D(n5906), .Y(n5907));
  AOI21X1 g4769(.A0(n5861), .A1(EBX_REG_3__SCAN_IN), .B0(n5907), .Y(n5908));
  OAI21X1 g4770(.A0(n5884), .A1(n5641), .B0(n5908), .Y(U2824));
  NAND3X1 g4771(.A(REIP_REG_3__SCAN_IN), .B(REIP_REG_2__SCAN_IN), .C(REIP_REG_1__SCAN_IN), .Y(n5910));
  XOR2X1  g4772(.A(n5910), .B(n1100), .Y(n5911));
  NAND2X1 g4773(.A(n5911), .B(n5864), .Y(n5912));
  NAND2X1 g4774(.A(n5865), .B(n5770), .Y(n5913));
  NAND3X1 g4775(.A(n5855), .B(n3219), .C(n1910), .Y(n5914));
  OAI21X1 g4776(.A0(n5855), .A1(n1100), .B0(n5914), .Y(n5915));
  AOI21X1 g4777(.A0(n5875), .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .B0(n5915), .Y(n5916));
  AOI22X1 g4778(.A0(n5873), .A1(n4525), .B0(n3170), .B1(n5876), .Y(n5917));
  NAND4X1 g4779(.A(n5916), .B(n5913), .C(n5912), .D(n5917), .Y(n5918));
  AOI21X1 g4780(.A0(n5861), .A1(EBX_REG_4__SCAN_IN), .B0(n5918), .Y(n5919));
  OAI21X1 g4781(.A0(n5884), .A1(n4539), .B0(n5919), .Y(U2823));
  NAND4X1 g4782(.A(REIP_REG_3__SCAN_IN), .B(REIP_REG_2__SCAN_IN), .C(REIP_REG_1__SCAN_IN), .D(REIP_REG_4__SCAN_IN), .Y(n5921));
  XOR2X1  g4783(.A(n5921), .B(n1097), .Y(n5922));
  NAND2X1 g4784(.A(n5922), .B(n5864), .Y(n5923));
  NAND2X1 g4785(.A(n5865), .B(n5773), .Y(n5924));
  OAI21X1 g4786(.A0(n5855), .A1(n1097), .B0(n5914), .Y(n5925));
  AOI21X1 g4787(.A0(n5875), .A1(PHYADDRPOINTER_REG_5__SCAN_IN), .B0(n5925), .Y(n5926));
  INVX1   g4788(.A(n4546), .Y(n5927));
  AOI22X1 g4789(.A0(n5873), .A1(n4566), .B0(n5927), .B1(n5876), .Y(n5928));
  NAND4X1 g4790(.A(n5926), .B(n5924), .C(n5923), .D(n5928), .Y(n5929));
  AOI21X1 g4791(.A0(n5861), .A1(EBX_REG_5__SCAN_IN), .B0(n5929), .Y(n5930));
  OAI21X1 g4792(.A0(n5884), .A1(n4562), .B0(n5930), .Y(U2822));
  NAND3X1 g4793(.A(n5855), .B(n5425), .C(STATE2_REG_1__SCAN_IN), .Y(n5932));
  NOR2X1  g4794(.A(n5921), .B(n1097), .Y(n5933));
  XOR2X1  g4795(.A(n5933), .B(REIP_REG_6__SCAN_IN), .Y(n5934));
  NAND2X1 g4796(.A(n5934), .B(n5864), .Y(n5935));
  NAND2X1 g4797(.A(n5865), .B(n5776), .Y(n5936));
  NAND2X1 g4798(.A(n5875), .B(PHYADDRPOINTER_REG_6__SCAN_IN), .Y(n5937));
  OAI21X1 g4799(.A0(n5855), .A1(n1094), .B0(n5914), .Y(n5938));
  AOI21X1 g4800(.A0(n5873), .A1(n4585), .B0(n5938), .Y(n5939));
  NAND4X1 g4801(.A(n5937), .B(n5936), .C(n5935), .D(n5939), .Y(n5940));
  AOI21X1 g4802(.A0(n5861), .A1(EBX_REG_6__SCAN_IN), .B0(n5940), .Y(n5941));
  OAI21X1 g4803(.A0(n5932), .A1(n5648), .B0(n5941), .Y(U2821));
  NOR3X1  g4804(.A(n5921), .B(n1094), .C(n1097), .Y(n5943));
  XOR2X1  g4805(.A(n5943), .B(REIP_REG_7__SCAN_IN), .Y(n5944));
  NAND2X1 g4806(.A(n5944), .B(n5864), .Y(n5945));
  NAND2X1 g4807(.A(n5865), .B(n5779), .Y(n5946));
  NAND2X1 g4808(.A(n5875), .B(PHYADDRPOINTER_REG_7__SCAN_IN), .Y(n5947));
  OAI21X1 g4809(.A0(n5855), .A1(n1091), .B0(n5914), .Y(n5948));
  AOI21X1 g4810(.A0(n5873), .A1(n4608), .B0(n5948), .Y(n5949));
  NAND4X1 g4811(.A(n5947), .B(n5946), .C(n5945), .D(n5949), .Y(n5950));
  AOI21X1 g4812(.A0(n5861), .A1(EBX_REG_7__SCAN_IN), .B0(n5950), .Y(n5951));
  OAI21X1 g4813(.A0(n5932), .A1(n4606), .B0(n5951), .Y(U2820));
  NOR4X1  g4814(.A(n1091), .B(n1094), .C(n1097), .D(n5921), .Y(n5953));
  XOR2X1  g4815(.A(n5953), .B(REIP_REG_8__SCAN_IN), .Y(n5954));
  NAND2X1 g4816(.A(n5954), .B(n5864), .Y(n5955));
  NAND2X1 g4817(.A(n5865), .B(n5782), .Y(n5956));
  NAND2X1 g4818(.A(n5875), .B(PHYADDRPOINTER_REG_8__SCAN_IN), .Y(n5957));
  OAI21X1 g4819(.A0(n5855), .A1(n1088), .B0(n5914), .Y(n5958));
  AOI21X1 g4820(.A0(n5873), .A1(n4633), .B0(n5958), .Y(n5959));
  NAND4X1 g4821(.A(n5957), .B(n5956), .C(n5955), .D(n5959), .Y(n5960));
  AOI21X1 g4822(.A0(n5861), .A1(EBX_REG_8__SCAN_IN), .B0(n5960), .Y(n5961));
  OAI21X1 g4823(.A0(n5932), .A1(n5653), .B0(n5961), .Y(U2819));
  NAND2X1 g4824(.A(n5953), .B(REIP_REG_8__SCAN_IN), .Y(n5963));
  XOR2X1  g4825(.A(n5963), .B(n1085), .Y(n5964));
  NAND2X1 g4826(.A(n5964), .B(n5864), .Y(n5965));
  NAND2X1 g4827(.A(n5865), .B(n5785), .Y(n5966));
  NAND2X1 g4828(.A(n5875), .B(PHYADDRPOINTER_REG_9__SCAN_IN), .Y(n5967));
  OAI21X1 g4829(.A0(n5855), .A1(n1085), .B0(n5914), .Y(n5968));
  AOI21X1 g4830(.A0(n5873), .A1(n4655), .B0(n5968), .Y(n5969));
  NAND4X1 g4831(.A(n5967), .B(n5966), .C(n5965), .D(n5969), .Y(n5970));
  AOI21X1 g4832(.A0(n5861), .A1(EBX_REG_9__SCAN_IN), .B0(n5970), .Y(n5971));
  OAI21X1 g4833(.A0(n5932), .A1(n4653), .B0(n5971), .Y(U2818));
  NAND3X1 g4834(.A(n5953), .B(REIP_REG_9__SCAN_IN), .C(REIP_REG_8__SCAN_IN), .Y(n5973));
  XOR2X1  g4835(.A(n5973), .B(n1082), .Y(n5974));
  NAND2X1 g4836(.A(n5974), .B(n5864), .Y(n5975));
  NAND2X1 g4837(.A(n5865), .B(n5788), .Y(n5976));
  NAND2X1 g4838(.A(n5875), .B(PHYADDRPOINTER_REG_10__SCAN_IN), .Y(n5977));
  OAI21X1 g4839(.A0(n5855), .A1(n1082), .B0(n5914), .Y(n5978));
  AOI21X1 g4840(.A0(n5873), .A1(n4682), .B0(n5978), .Y(n5979));
  NAND4X1 g4841(.A(n5977), .B(n5976), .C(n5975), .D(n5979), .Y(n5980));
  AOI21X1 g4842(.A0(n5861), .A1(EBX_REG_10__SCAN_IN), .B0(n5980), .Y(n5981));
  OAI21X1 g4843(.A0(n5932), .A1(n4680), .B0(n5981), .Y(U2817));
  NAND4X1 g4844(.A(REIP_REG_10__SCAN_IN), .B(REIP_REG_9__SCAN_IN), .C(REIP_REG_8__SCAN_IN), .D(n5953), .Y(n5983));
  XOR2X1  g4845(.A(n5983), .B(n1079), .Y(n5984));
  NAND2X1 g4846(.A(n5984), .B(n5864), .Y(n5985));
  NAND2X1 g4847(.A(n5865), .B(n5791), .Y(n5986));
  NAND2X1 g4848(.A(n5875), .B(PHYADDRPOINTER_REG_11__SCAN_IN), .Y(n5987));
  OAI21X1 g4849(.A0(n5855), .A1(n1079), .B0(n5914), .Y(n5988));
  AOI21X1 g4850(.A0(n5873), .A1(n4703), .B0(n5988), .Y(n5989));
  NAND4X1 g4851(.A(n5987), .B(n5986), .C(n5985), .D(n5989), .Y(n5990));
  AOI21X1 g4852(.A0(n5861), .A1(EBX_REG_11__SCAN_IN), .B0(n5990), .Y(n5991));
  OAI21X1 g4853(.A0(n5932), .A1(n5660), .B0(n5991), .Y(U2816));
  NOR2X1  g4854(.A(n5983), .B(n1079), .Y(n5993));
  XOR2X1  g4855(.A(n5993), .B(REIP_REG_12__SCAN_IN), .Y(n5994));
  NAND2X1 g4856(.A(n5994), .B(n5864), .Y(n5995));
  NAND2X1 g4857(.A(n5865), .B(n5794), .Y(n5996));
  NAND2X1 g4858(.A(n5875), .B(PHYADDRPOINTER_REG_12__SCAN_IN), .Y(n5997));
  OAI21X1 g4859(.A0(n5855), .A1(n1076), .B0(n5914), .Y(n5998));
  AOI21X1 g4860(.A0(n5873), .A1(n4726), .B0(n5998), .Y(n5999));
  NAND4X1 g4861(.A(n5997), .B(n5996), .C(n5995), .D(n5999), .Y(n6000));
  AOI21X1 g4862(.A0(n5861), .A1(EBX_REG_12__SCAN_IN), .B0(n6000), .Y(n6001));
  OAI21X1 g4863(.A0(n5932), .A1(n4724), .B0(n6001), .Y(U2815));
  NOR3X1  g4864(.A(n5983), .B(n1076), .C(n1079), .Y(n6003));
  XOR2X1  g4865(.A(n6003), .B(REIP_REG_13__SCAN_IN), .Y(n6004));
  NAND2X1 g4866(.A(n6004), .B(n5864), .Y(n6005));
  NAND2X1 g4867(.A(n5865), .B(n5797), .Y(n6006));
  NAND2X1 g4868(.A(n5875), .B(PHYADDRPOINTER_REG_13__SCAN_IN), .Y(n6007));
  OAI21X1 g4869(.A0(n5855), .A1(n1073), .B0(n5914), .Y(n6008));
  AOI21X1 g4870(.A0(n5873), .A1(n4741), .B0(n6008), .Y(n6009));
  NAND4X1 g4871(.A(n6007), .B(n6006), .C(n6005), .D(n6009), .Y(n6010));
  AOI21X1 g4872(.A0(n5861), .A1(EBX_REG_13__SCAN_IN), .B0(n6010), .Y(n6011));
  OAI21X1 g4873(.A0(n5932), .A1(n4753), .B0(n6011), .Y(U2814));
  NOR4X1  g4874(.A(n1073), .B(n1076), .C(n1079), .D(n5983), .Y(n6013));
  XOR2X1  g4875(.A(n6013), .B(REIP_REG_14__SCAN_IN), .Y(n6014));
  NAND2X1 g4876(.A(n6014), .B(n5864), .Y(n6015));
  NAND2X1 g4877(.A(n5865), .B(n5800), .Y(n6016));
  NAND2X1 g4878(.A(n5875), .B(PHYADDRPOINTER_REG_14__SCAN_IN), .Y(n6017));
  OAI21X1 g4879(.A0(n5855), .A1(n1070), .B0(n5914), .Y(n6018));
  AOI21X1 g4880(.A0(n5873), .A1(n4764), .B0(n6018), .Y(n6019));
  NAND4X1 g4881(.A(n6017), .B(n6016), .C(n6015), .D(n6019), .Y(n6020));
  AOI21X1 g4882(.A0(n5861), .A1(EBX_REG_14__SCAN_IN), .B0(n6020), .Y(n6021));
  OAI21X1 g4883(.A0(n5932), .A1(n5668), .B0(n6021), .Y(U2813));
  NAND2X1 g4884(.A(n6013), .B(REIP_REG_14__SCAN_IN), .Y(n6023));
  XOR2X1  g4885(.A(n6023), .B(n1067), .Y(n6024));
  NAND2X1 g4886(.A(n6024), .B(n5864), .Y(n6025));
  NAND2X1 g4887(.A(n5865), .B(n5803), .Y(n6026));
  NAND2X1 g4888(.A(n5875), .B(PHYADDRPOINTER_REG_15__SCAN_IN), .Y(n6027));
  OAI21X1 g4889(.A0(n5855), .A1(n1067), .B0(n5914), .Y(n6028));
  AOI21X1 g4890(.A0(n5873), .A1(n4787), .B0(n6028), .Y(n6029));
  NAND4X1 g4891(.A(n6027), .B(n6026), .C(n6025), .D(n6029), .Y(n6030));
  AOI21X1 g4892(.A0(n5861), .A1(EBX_REG_15__SCAN_IN), .B0(n6030), .Y(n6031));
  OAI21X1 g4893(.A0(n5932), .A1(n5673), .B0(n6031), .Y(U2812));
  NAND3X1 g4894(.A(n6013), .B(REIP_REG_15__SCAN_IN), .C(REIP_REG_14__SCAN_IN), .Y(n6033));
  XOR2X1  g4895(.A(n6033), .B(n1064), .Y(n6034));
  NAND2X1 g4896(.A(n6034), .B(n5864), .Y(n6035));
  NAND2X1 g4897(.A(n5865), .B(n5806), .Y(n6036));
  NAND2X1 g4898(.A(n5875), .B(PHYADDRPOINTER_REG_16__SCAN_IN), .Y(n6037));
  OAI21X1 g4899(.A0(n5855), .A1(n1064), .B0(n5914), .Y(n6038));
  AOI21X1 g4900(.A0(n5873), .A1(n4877), .B0(n6038), .Y(n6039));
  NAND4X1 g4901(.A(n6037), .B(n6036), .C(n6035), .D(n6039), .Y(n6040));
  AOI21X1 g4902(.A0(n5861), .A1(EBX_REG_16__SCAN_IN), .B0(n6040), .Y(n6041));
  OAI21X1 g4903(.A0(n5932), .A1(n5676), .B0(n6041), .Y(U2811));
  NAND4X1 g4904(.A(REIP_REG_15__SCAN_IN), .B(REIP_REG_14__SCAN_IN), .C(REIP_REG_16__SCAN_IN), .D(n6013), .Y(n6043));
  XOR2X1  g4905(.A(n6043), .B(n1061), .Y(n6044));
  NAND2X1 g4906(.A(n6044), .B(n5864), .Y(n6045));
  NAND2X1 g4907(.A(n5865), .B(n5809), .Y(n6046));
  NAND2X1 g4908(.A(n5875), .B(PHYADDRPOINTER_REG_17__SCAN_IN), .Y(n6047));
  OAI21X1 g4909(.A0(n5855), .A1(n1061), .B0(n5914), .Y(n6048));
  AOI21X1 g4910(.A0(n5873), .A1(n4906), .B0(n6048), .Y(n6049));
  NAND4X1 g4911(.A(n6047), .B(n6046), .C(n6045), .D(n6049), .Y(n6050));
  AOI21X1 g4912(.A0(n5861), .A1(EBX_REG_17__SCAN_IN), .B0(n6050), .Y(n6051));
  OAI21X1 g4913(.A0(n5932), .A1(n5683), .B0(n6051), .Y(U2810));
  NOR2X1  g4914(.A(n6043), .B(n1061), .Y(n6053));
  XOR2X1  g4915(.A(n6053), .B(REIP_REG_18__SCAN_IN), .Y(n6054));
  NAND2X1 g4916(.A(n6054), .B(n5864), .Y(n6055));
  NAND2X1 g4917(.A(n5865), .B(n5812), .Y(n6056));
  NAND2X1 g4918(.A(n5875), .B(PHYADDRPOINTER_REG_18__SCAN_IN), .Y(n6057));
  OAI21X1 g4919(.A0(n5855), .A1(n1058), .B0(n5914), .Y(n6058));
  AOI21X1 g4920(.A0(n5873), .A1(n4936), .B0(n6058), .Y(n6059));
  NAND4X1 g4921(.A(n6057), .B(n6056), .C(n6055), .D(n6059), .Y(n6060));
  AOI21X1 g4922(.A0(n5861), .A1(EBX_REG_18__SCAN_IN), .B0(n6060), .Y(n6061));
  OAI21X1 g4923(.A0(n5932), .A1(n4934), .B0(n6061), .Y(U2809));
  NOR3X1  g4924(.A(n6043), .B(n1061), .C(n1058), .Y(n6063));
  XOR2X1  g4925(.A(n6063), .B(REIP_REG_19__SCAN_IN), .Y(n6064));
  NAND2X1 g4926(.A(n6064), .B(n5864), .Y(n6065));
  NAND2X1 g4927(.A(n5865), .B(n5815), .Y(n6066));
  NAND2X1 g4928(.A(n5875), .B(PHYADDRPOINTER_REG_19__SCAN_IN), .Y(n6067));
  OAI21X1 g4929(.A0(n5855), .A1(n1055), .B0(n5914), .Y(n6068));
  AOI21X1 g4930(.A0(n5873), .A1(n4970), .B0(n6068), .Y(n6069));
  NAND4X1 g4931(.A(n6067), .B(n6066), .C(n6065), .D(n6069), .Y(n6070));
  AOI21X1 g4932(.A0(n5861), .A1(EBX_REG_19__SCAN_IN), .B0(n6070), .Y(n6071));
  OAI21X1 g4933(.A0(n5932), .A1(n5690), .B0(n6071), .Y(U2808));
  INVX1   g4934(.A(n5864), .Y(n6073));
  NOR4X1  g4935(.A(n1061), .B(n1058), .C(n1055), .D(n6043), .Y(n6074));
  XOR2X1  g4936(.A(n6074), .B(n1052), .Y(n6075));
  AOI22X1 g4937(.A0(n5871), .A1(REIP_REG_20__SCAN_IN), .B0(n5008), .B1(n5873), .Y(n6076));
  OAI21X1 g4938(.A0(n5887), .A1(n5016), .B0(n6076), .Y(n6077));
  AOI21X1 g4939(.A0(n5865), .A1(n4126), .B0(n6077), .Y(n6078));
  OAI21X1 g4940(.A0(n6075), .A1(n6073), .B0(n6078), .Y(n6079));
  AOI21X1 g4941(.A0(n5861), .A1(EBX_REG_20__SCAN_IN), .B0(n6079), .Y(n6080));
  OAI21X1 g4942(.A0(n5932), .A1(n5694), .B0(n6080), .Y(U2807));
  NAND2X1 g4943(.A(n6074), .B(REIP_REG_20__SCAN_IN), .Y(n6082));
  XOR2X1  g4944(.A(n6082), .B(n1049), .Y(n6083));
  NAND2X1 g4945(.A(n6083), .B(n5864), .Y(n6084));
  NAND2X1 g4946(.A(n5865), .B(n5820), .Y(n6085));
  OAI22X1 g4947(.A0(n5855), .A1(n1049), .B0(n5018), .B1(n5872), .Y(n6086));
  AOI21X1 g4948(.A0(n5875), .A1(PHYADDRPOINTER_REG_21__SCAN_IN), .B0(n6086), .Y(n6087));
  NAND3X1 g4949(.A(n6087), .B(n6085), .C(n6084), .Y(n6088));
  AOI21X1 g4950(.A0(n5861), .A1(EBX_REG_21__SCAN_IN), .B0(n6088), .Y(n6089));
  OAI21X1 g4951(.A0(n5932), .A1(n5699), .B0(n6089), .Y(U2806));
  NAND3X1 g4952(.A(n6074), .B(REIP_REG_20__SCAN_IN), .C(REIP_REG_21__SCAN_IN), .Y(n6091));
  XOR2X1  g4953(.A(n6091), .B(n1046), .Y(n6092));
  NAND2X1 g4954(.A(n6092), .B(n5864), .Y(n6093));
  NAND2X1 g4955(.A(n5865), .B(n5823), .Y(n6094));
  OAI22X1 g4956(.A0(n5855), .A1(n1046), .B0(n5050), .B1(n5872), .Y(n6095));
  AOI21X1 g4957(.A0(n5875), .A1(PHYADDRPOINTER_REG_22__SCAN_IN), .B0(n6095), .Y(n6096));
  NAND3X1 g4958(.A(n6096), .B(n6094), .C(n6093), .Y(n6097));
  AOI21X1 g4959(.A0(n5861), .A1(EBX_REG_22__SCAN_IN), .B0(n6097), .Y(n6098));
  OAI21X1 g4960(.A0(n5932), .A1(n5703), .B0(n6098), .Y(U2805));
  NAND4X1 g4961(.A(REIP_REG_20__SCAN_IN), .B(REIP_REG_21__SCAN_IN), .C(REIP_REG_22__SCAN_IN), .D(n6074), .Y(n6100));
  XOR2X1  g4962(.A(n6100), .B(n1043), .Y(n6101));
  NAND2X1 g4963(.A(n6101), .B(n5864), .Y(n6102));
  NAND2X1 g4964(.A(n5865), .B(n5826), .Y(n6103));
  OAI22X1 g4965(.A0(n5855), .A1(n1043), .B0(n5123), .B1(n5872), .Y(n6104));
  AOI21X1 g4966(.A0(n5875), .A1(PHYADDRPOINTER_REG_23__SCAN_IN), .B0(n6104), .Y(n6105));
  NAND3X1 g4967(.A(n6105), .B(n6103), .C(n6102), .Y(n6106));
  AOI21X1 g4968(.A0(n5861), .A1(EBX_REG_23__SCAN_IN), .B0(n6106), .Y(n6107));
  OAI21X1 g4969(.A0(n5932), .A1(n5707), .B0(n6107), .Y(U2804));
  NOR2X1  g4970(.A(n6100), .B(n1043), .Y(n6109));
  XOR2X1  g4971(.A(n6109), .B(n1040), .Y(n6110));
  NAND2X1 g4972(.A(n5875), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .Y(n6111));
  AOI22X1 g4973(.A0(n5871), .A1(REIP_REG_24__SCAN_IN), .B0(n5164), .B1(n5873), .Y(n6112));
  NAND2X1 g4974(.A(n6112), .B(n6111), .Y(n6113));
  AOI21X1 g4975(.A0(n5865), .A1(n5829), .B0(n6113), .Y(n6114));
  OAI21X1 g4976(.A0(n6110), .A1(n6073), .B0(n6114), .Y(n6115));
  AOI21X1 g4977(.A0(n5861), .A1(EBX_REG_24__SCAN_IN), .B0(n6115), .Y(n6116));
  OAI21X1 g4978(.A0(n5932), .A1(n5711), .B0(n6116), .Y(U2803));
  NOR3X1  g4979(.A(n6100), .B(n1043), .C(n1040), .Y(n6118));
  XOR2X1  g4980(.A(n6118), .B(REIP_REG_25__SCAN_IN), .Y(n6119));
  NAND2X1 g4981(.A(n6119), .B(n5864), .Y(n6120));
  NAND2X1 g4982(.A(n5865), .B(n4254), .Y(n6121));
  NAND2X1 g4983(.A(n5875), .B(PHYADDRPOINTER_REG_25__SCAN_IN), .Y(n6122));
  AOI22X1 g4984(.A0(n5871), .A1(REIP_REG_25__SCAN_IN), .B0(n5199), .B1(n5873), .Y(n6123));
  NAND4X1 g4985(.A(n6122), .B(n6121), .C(n6120), .D(n6123), .Y(n6124));
  AOI21X1 g4986(.A0(n5861), .A1(EBX_REG_25__SCAN_IN), .B0(n6124), .Y(n6125));
  OAI21X1 g4987(.A0(n5932), .A1(n5716), .B0(n6125), .Y(U2802));
  NOR4X1  g4988(.A(n1043), .B(n1040), .C(n1037), .D(n6100), .Y(n6127));
  XOR2X1  g4989(.A(n6127), .B(n1034), .Y(n6128));
  NAND2X1 g4990(.A(n5875), .B(PHYADDRPOINTER_REG_26__SCAN_IN), .Y(n6129));
  AOI22X1 g4991(.A0(n5871), .A1(REIP_REG_26__SCAN_IN), .B0(n5239), .B1(n5873), .Y(n6130));
  NAND2X1 g4992(.A(n6130), .B(n6129), .Y(n6131));
  AOI21X1 g4993(.A0(n5865), .A1(n5834), .B0(n6131), .Y(n6132));
  OAI21X1 g4994(.A0(n6128), .A1(n6073), .B0(n6132), .Y(n6133));
  AOI21X1 g4995(.A0(n5861), .A1(EBX_REG_26__SCAN_IN), .B0(n6133), .Y(n6134));
  OAI21X1 g4996(.A0(n5932), .A1(n5251), .B0(n6134), .Y(U2801));
  NAND2X1 g4997(.A(n6127), .B(REIP_REG_26__SCAN_IN), .Y(n6136));
  XOR2X1  g4998(.A(n6136), .B(n1031), .Y(n6137));
  NAND2X1 g4999(.A(n6137), .B(n5864), .Y(n6138));
  NAND2X1 g5000(.A(n5865), .B(n4306), .Y(n6139));
  OAI22X1 g5001(.A0(n5855), .A1(n1031), .B0(n5275), .B1(n5872), .Y(n6140));
  AOI21X1 g5002(.A0(n5875), .A1(PHYADDRPOINTER_REG_27__SCAN_IN), .B0(n6140), .Y(n6141));
  NAND3X1 g5003(.A(n6141), .B(n6139), .C(n6138), .Y(n6142));
  AOI21X1 g5004(.A0(n5861), .A1(EBX_REG_27__SCAN_IN), .B0(n6142), .Y(n6143));
  OAI21X1 g5005(.A0(n5932), .A1(n5725), .B0(n6143), .Y(U2800));
  INVX1   g5006(.A(n5865), .Y(n6145));
  NAND3X1 g5007(.A(n6127), .B(REIP_REG_26__SCAN_IN), .C(REIP_REG_27__SCAN_IN), .Y(n6146));
  XOR2X1  g5008(.A(n6146), .B(REIP_REG_28__SCAN_IN), .Y(n6147));
  NOR2X1  g5009(.A(n6147), .B(n6073), .Y(n6148));
  AOI22X1 g5010(.A0(n5871), .A1(REIP_REG_28__SCAN_IN), .B0(n5309), .B1(n5873), .Y(n6149));
  OAI21X1 g5011(.A0(n5887), .A1(n5307), .B0(n6149), .Y(n6150));
  NOR2X1  g5012(.A(n6150), .B(n6148), .Y(n6151));
  OAI21X1 g5013(.A0(n6145), .A1(n4330), .B0(n6151), .Y(n6152));
  AOI21X1 g5014(.A0(n5861), .A1(EBX_REG_28__SCAN_IN), .B0(n6152), .Y(n6153));
  OAI21X1 g5015(.A0(n5932), .A1(n5731), .B0(n6153), .Y(U2799));
  INVX1   g5016(.A(EBX_REG_29__SCAN_IN), .Y(n6155));
  NAND4X1 g5017(.A(REIP_REG_26__SCAN_IN), .B(REIP_REG_27__SCAN_IN), .C(REIP_REG_28__SCAN_IN), .D(n6127), .Y(n6156));
  XOR2X1  g5018(.A(n6156), .B(REIP_REG_29__SCAN_IN), .Y(n6157));
  NOR2X1  g5019(.A(n6157), .B(n6073), .Y(n6158));
  AOI22X1 g5020(.A0(n5871), .A1(REIP_REG_29__SCAN_IN), .B0(n5360), .B1(n5873), .Y(n6159));
  OAI21X1 g5021(.A0(n5887), .A1(n5358), .B0(n6159), .Y(n6160));
  NOR2X1  g5022(.A(n6160), .B(n6158), .Y(n6161));
  OAI21X1 g5023(.A0(n5860), .A1(n6155), .B0(n6161), .Y(n6162));
  AOI21X1 g5024(.A0(n5865), .A1(n4356), .B0(n6162), .Y(n6163));
  OAI21X1 g5025(.A0(n5932), .A1(n5737), .B0(n6163), .Y(U2798));
  NOR2X1  g5026(.A(n6145), .B(n4382), .Y(n6165));
  NAND2X1 g5027(.A(n5861), .B(EBX_REG_30__SCAN_IN), .Y(n6166));
  NOR2X1  g5028(.A(n6156), .B(n1025), .Y(n6167));
  XOR2X1  g5029(.A(n6167), .B(REIP_REG_30__SCAN_IN), .Y(n6168));
  NAND2X1 g5030(.A(n6168), .B(n5864), .Y(n6169));
  OAI22X1 g5031(.A0(n5855), .A1(n1020), .B0(n5394), .B1(n5872), .Y(n6170));
  AOI21X1 g5032(.A0(n5875), .A1(PHYADDRPOINTER_REG_30__SCAN_IN), .B0(n6170), .Y(n6171));
  NAND3X1 g5033(.A(n6171), .B(n6169), .C(n6166), .Y(n6172));
  NOR2X1  g5034(.A(n6172), .B(n6165), .Y(n6173));
  OAI21X1 g5035(.A0(n5932), .A1(n5743), .B0(n6173), .Y(U2797));
  NOR2X1  g5036(.A(n6145), .B(n4405), .Y(n6175));
  NOR2X1  g5037(.A(n5860), .B(n5848), .Y(n6176));
  NOR3X1  g5038(.A(n6156), .B(n1025), .C(n1020), .Y(n6177));
  XOR2X1  g5039(.A(n6177), .B(n5432), .Y(n6178));
  OAI22X1 g5040(.A0(n5855), .A1(n5432), .B0(n5424), .B1(n5872), .Y(n6179));
  AOI21X1 g5041(.A0(n5875), .A1(PHYADDRPOINTER_REG_31__SCAN_IN), .B0(n6179), .Y(n6180));
  OAI21X1 g5042(.A0(n6178), .A1(n6073), .B0(n6180), .Y(n6181));
  NOR3X1  g5043(.A(n6181), .B(n6176), .C(n6175), .Y(n6182));
  OAI21X1 g5044(.A0(n5932), .A1(n5749), .B0(n6182), .Y(U2796));
  NOR4X1  g5045(.A(DATAWIDTH_REG_15__SCAN_IN), .B(DATAWIDTH_REG_14__SCAN_IN), .C(DATAWIDTH_REG_13__SCAN_IN), .D(DATAWIDTH_REG_16__SCAN_IN), .Y(n6184));
  NOR4X1  g5046(.A(DATAWIDTH_REG_12__SCAN_IN), .B(DATAWIDTH_REG_11__SCAN_IN), .C(DATAWIDTH_REG_10__SCAN_IN), .D(DATAWIDTH_REG_26__SCAN_IN), .Y(n6185));
  NOR4X1  g5047(.A(DATAWIDTH_REG_7__SCAN_IN), .B(DATAWIDTH_REG_6__SCAN_IN), .C(DATAWIDTH_REG_5__SCAN_IN), .D(DATAWIDTH_REG_8__SCAN_IN), .Y(n6186));
  NOR4X1  g5048(.A(DATAWIDTH_REG_4__SCAN_IN), .B(DATAWIDTH_REG_3__SCAN_IN), .C(DATAWIDTH_REG_2__SCAN_IN), .D(DATAWIDTH_REG_17__SCAN_IN), .Y(n6187));
  NAND4X1 g5049(.A(n6186), .B(n6185), .C(n6184), .D(n6187), .Y(n6188));
  NOR4X1  g5050(.A(DATAWIDTH_REG_22__SCAN_IN), .B(DATAWIDTH_REG_21__SCAN_IN), .C(DATAWIDTH_REG_20__SCAN_IN), .D(DATAWIDTH_REG_23__SCAN_IN), .Y(n6189));
  INVX1   g5051(.A(DATAWIDTH_REG_0__SCAN_IN), .Y(n6190));
  NOR2X1  g5052(.A(n1152), .B(n6190), .Y(n6191));
  NOR3X1  g5053(.A(n6191), .B(DATAWIDTH_REG_19__SCAN_IN), .C(DATAWIDTH_REG_18__SCAN_IN), .Y(n6192));
  NOR4X1  g5054(.A(DATAWIDTH_REG_29__SCAN_IN), .B(DATAWIDTH_REG_28__SCAN_IN), .C(DATAWIDTH_REG_27__SCAN_IN), .D(DATAWIDTH_REG_30__SCAN_IN), .Y(n6193));
  NOR4X1  g5055(.A(DATAWIDTH_REG_25__SCAN_IN), .B(DATAWIDTH_REG_24__SCAN_IN), .C(DATAWIDTH_REG_9__SCAN_IN), .D(DATAWIDTH_REG_31__SCAN_IN), .Y(n6194));
  NAND4X1 g5056(.A(n6193), .B(n6192), .C(n6189), .D(n6194), .Y(n6195));
  NOR2X1  g5057(.A(n6195), .B(n6188), .Y(n6196));
  NAND3X1 g5058(.A(n6196), .B(n1109), .C(n1152), .Y(n6197));
  NOR2X1  g5059(.A(DATAWIDTH_REG_1__SCAN_IN), .B(DATAWIDTH_REG_0__SCAN_IN), .Y(n6198));
  NAND3X1 g5060(.A(n6198), .B(n6196), .C(n3252), .Y(n6199));
  OAI21X1 g5061(.A0(n6195), .A1(n6188), .B0(BYTEENABLE_REG_3__SCAN_IN), .Y(n6200));
  NAND3X1 g5062(.A(n6200), .B(n6199), .C(n6197), .Y(U2795));
  NAND2X1 g5063(.A(REIP_REG_1__SCAN_IN), .B(REIP_REG_0__SCAN_IN), .Y(n6202));
  AOI21X1 g5064(.A0(n3252), .A1(DATAWIDTH_REG_0__SCAN_IN), .B0(n6198), .Y(n6203));
  OAI21X1 g5065(.A0(n6203), .A1(REIP_REG_1__SCAN_IN), .B0(n6202), .Y(n6204));
  NAND2X1 g5066(.A(n6204), .B(n6196), .Y(n6205));
  OAI21X1 g5067(.A0(n6196), .A1(n1009), .B0(n6205), .Y(U3468));
  NAND2X1 g5068(.A(n6196), .B(REIP_REG_1__SCAN_IN), .Y(n6207));
  OAI21X1 g5069(.A0(n6195), .A1(n6188), .B0(BYTEENABLE_REG_1__SCAN_IN), .Y(n6208));
  NAND3X1 g5070(.A(n6208), .B(n6207), .C(n6199), .Y(U2794));
  OAI21X1 g5071(.A0(REIP_REG_1__SCAN_IN), .A1(REIP_REG_0__SCAN_IN), .B0(n6196), .Y(n6210));
  OAI21X1 g5072(.A0(n6196), .A1(n1017), .B0(n6210), .Y(U3469));
  OAI21X1 g5073(.A0(STATE_REG_0__SCAN_IN), .A1(n1006), .B0(W_R_N_REG_SCAN_IN), .Y(n6212));
  OAI21X1 g5074(.A0(n1011), .A1(READREQUEST_REG_SCAN_IN), .B0(n6212), .Y(U3470));
  NOR2X1  g5075(.A(n2103), .B(n2044), .Y(n6214));
  OAI21X1 g5076(.A0(n6214), .A1(n2015), .B0(n4437), .Y(U2793));
  NAND2X1 g5077(.A(n6214), .B(n2053), .Y(n6216));
  OAI21X1 g5078(.A0(n2103), .A1(n2044), .B0(MORE_REG_SCAN_IN), .Y(n6217));
  NAND2X1 g5079(.A(n6217), .B(n6216), .Y(U3471));
  AOI22X1 g5080(.A0(n1123), .A1(n1004), .B0(STATEBS16_REG_SCAN_IN), .B1(n1149), .Y(n6219));
  OAI21X1 g5081(.A0(n1149), .A1(n1146), .B0(n6219), .Y(U2792));
  NAND4X1 g5082(.A(STATE2_REG_1__SCAN_IN), .B(STATE2_REG_2__SCAN_IN), .C(n1113), .D(n1217), .Y(n6221));
  NAND4X1 g5083(.A(n5853), .B(n3220), .C(n1907), .D(n6221), .Y(n6222));
  AOI21X1 g5084(.A0(n2041), .A1(STATEBS16_REG_SCAN_IN), .B0(n1721), .Y(n6223));
  NOR3X1  g5085(.A(n6223), .B(n1833), .C(READY_N), .Y(n6224));
  AOI22X1 g5086(.A0(n1465), .A1(n2042), .B0(n1910), .B1(n1833), .Y(n6225));
  OAI21X1 g5087(.A0(n6224), .A1(n1217), .B0(n6225), .Y(n6226));
  NAND2X1 g5088(.A(n6222), .B(n6226), .Y(n6227));
  OAI21X1 g5089(.A0(n6222), .A1(n1116), .B0(n6227), .Y(U3472));
  OAI21X1 g5090(.A0(STATE_REG_0__SCAN_IN), .A1(n1006), .B0(D_C_N_REG_SCAN_IN), .Y(n6229));
  NOR3X1  g5091(.A(STATE_REG_0__SCAN_IN), .B(n1006), .C(CODEFETCH_REG_SCAN_IN), .Y(n6230));
  AOI21X1 g5092(.A0(n1123), .A1(n1004), .B0(n6230), .Y(n6231));
  NAND2X1 g5093(.A(n6231), .B(n6229), .Y(U2791));
  NAND3X1 g5094(.A(n1004), .B(STATE_REG_1__SCAN_IN), .C(MEMORYFETCH_REG_SCAN_IN), .Y(n6233));
  OAI21X1 g5095(.A0(STATE_REG_0__SCAN_IN), .A1(n1006), .B0(M_IO_N_REG_SCAN_IN), .Y(n6234));
  NAND2X1 g5096(.A(n6234), .B(n6233), .Y(U3473));
  NAND2X1 g5097(.A(n3219), .B(n1910), .Y(n6236));
  OAI21X1 g5098(.A0(n2103), .A1(n2040), .B0(CODEFETCH_REG_SCAN_IN), .Y(n6237));
  OAI21X1 g5099(.A0(n6236), .A1(n1217), .B0(n6237), .Y(U2790));
  NAND2X1 g5100(.A(STATE_REG_0__SCAN_IN), .B(ADS_N_REG_SCAN_IN), .Y(n6239));
  NAND2X1 g5101(.A(n6239), .B(n1149), .Y(U2789));
  NAND3X1 g5102(.A(n1683), .B(n1678), .C(STATE2_REG_2__SCAN_IN), .Y(n6241));
  NAND2X1 g5103(.A(n6236), .B(n5853), .Y(n6242));
  NAND2X1 g5104(.A(n6242), .B(n6241), .Y(n6243));
  NAND3X1 g5105(.A(n6236), .B(n5853), .C(READREQUEST_REG_SCAN_IN), .Y(n6244));
  NAND2X1 g5106(.A(n6244), .B(n6243), .Y(U3474));
  NOR2X1  g5107(.A(n2038), .B(n2037), .Y(n6246));
  NAND3X1 g5108(.A(n6246), .B(n1834), .C(n1476), .Y(n6247));
  OAI21X1 g5109(.A0(n6247), .A1(n2034), .B0(MEMORYFETCH_REG_SCAN_IN), .Y(n6248));
  AOI21X1 g5110(.A0(n3219), .A1(n1910), .B0(n5850), .Y(n6249));
  NAND2X1 g5111(.A(n6249), .B(n6248), .Y(U2788));
endmodule


