//Converted to Combinational (Partial output: n55) , Module name: s1488_n55 , Timestamp: 2018-12-03T15:51:02.596895 
module s1488_n55 ( v1, CLR, v7, v2, v10, v8, v9, v11, v12, v3, v0, v5, v4, v6, n55 );
input v1, CLR, v7, v2, v10, v8, v9, v11, v12, v3, v0, v5, v4, v6;
output n55;
wire n267, n283, n291, n45, n271, n282, n290, n285, n72, n268, n270, n281, n68, n275, n289, n66, n196, n284, n184, n241, n82, n63, n269, n277, n280, n279, n272, n116, n274, n286, n287, n288, n217, n109, n103, n54, n276, n142, n278, n49, n53, n111, n273, n47, n48, n259, n98, n104, n91;
AOI21X1  g247(.A0(n291), .A1(n283), .B0(n267), .Y(n55));
INVX1    g222(.A(CLR), .Y(n267));
OAI21X1  g238(.A0(n282), .A1(n271), .B0(n45), .Y(n283));
AOI21X1  g246(.A0(n285), .A1(v7), .B0(n290), .Y(n291));
INVX1    g000(.A(v7), .Y(n45));
AOI21X1  g226(.A0(n270), .A1(n268), .B0(n72), .Y(n271));
OAI21X1  g237(.A0(n275), .A1(n68), .B0(n281), .Y(n282));
OAI22X1  g245(.A0(n196), .A1(n66), .B0(v2), .B1(n289), .Y(n290));
OAI22X1  g240(.A0(n241), .A1(n184), .B0(v10), .B1(n284), .Y(n285));
INVX1    g027(.A(v8), .Y(n72));
NAND4X1  g223(.A(n68), .B(v11), .C(n82), .D(v9), .Y(n268));
OAI21X1  g225(.A0(n269), .A1(n63), .B0(v10), .Y(n270));
AOI22X1  g236(.A0(n279), .A1(n280), .B0(n277), .B1(n72), .Y(n281));
INVX1    g023(.A(v10), .Y(n68));
AOI21X1  g230(.A0(n274), .A1(n116), .B0(n272), .Y(n275));
AOI21X1  g244(.A0(n288), .A1(n287), .B0(n286), .Y(n289));
NAND2X1  g021(.A(v8), .B(v10), .Y(n66));
OR2X1    g151(.A(v9), .B(v12), .Y(n196));
AOI22X1  g239(.A0(n109), .A1(n72), .B0(n217), .B1(n196), .Y(n284));
NAND2X1  g139(.A(v11), .B(n82), .Y(n184));
NAND2X1  g196(.A(v9), .B(v10), .Y(n241));
INVX1    g037(.A(v12), .Y(n82));
INVX1    g018(.A(v9), .Y(n63));
AOI21X1  g224(.A0(n54), .A1(n103), .B0(n184), .Y(n269));
OAI21X1  g232(.A0(n142), .A1(n63), .B0(n276), .Y(n277));
AND2X1   g235(.A(v12), .B(v3), .Y(n280));
OAI22X1  g234(.A0(n111), .A1(n53), .B0(n49), .B1(n278), .Y(n279));
NOR3X1   g227(.A(v9), .B(v11), .C(v12), .Y(n272));
INVX1    g071(.A(v0), .Y(n116));
OAI22X1  g229(.A0(n196), .A1(n54), .B0(n47), .B1(n273), .Y(n274));
NOR3X1   g241(.A(n142), .B(n72), .C(v9), .Y(n286));
NOR3X1   g242(.A(n98), .B(n259), .C(n48), .Y(n287));
NOR3X1   g243(.A(n111), .B(v8), .C(n63), .Y(n288));
NOR2X1   g172(.A(n72), .B(v11), .Y(n217));
NOR2X1   g064(.A(n104), .B(v12), .Y(n109));
INVX1    g058(.A(v2), .Y(n103));
NAND2X1  g009(.A(v4), .B(v5), .Y(n54));
NAND4X1  g231(.A(n63), .B(v12), .C(v6), .D(n91), .Y(n276));
NAND2X1  g097(.A(v10), .B(v11), .Y(n142));
NAND4X1  g233(.A(v10), .B(v11), .C(v0), .D(v8), .Y(n278));
NOR2X1   g004(.A(v1), .B(n48), .Y(n49));
OR2X1    g008(.A(v8), .B(v9), .Y(n53));
OR2X1    g066(.A(v10), .B(v11), .Y(n111));
NAND4X1  g228(.A(n259), .B(v3), .C(v6), .D(v8), .Y(n273));
NAND2X1  g002(.A(v11), .B(v12), .Y(n47));
INVX1    g003(.A(v6), .Y(n48));
INVX1    g214(.A(v1), .Y(n259));
OR2X1    g053(.A(v7), .B(v12), .Y(n98));
INVX1    g059(.A(v11), .Y(n104));
NOR2X1   g046(.A(v10), .B(v11), .Y(n91));

endmodule
