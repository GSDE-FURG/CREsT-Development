//Converted to Combinational (Partial output: n3126) , Module name: s38584_n3126 , Timestamp: 2018-12-03T15:51:16.919647 
module s38584_n3126 ( g35, g6311, g4826, g4688, g4801, g4793, g4776, g4653, g4669, g4659, g4709, g4785, g4765, g6381, g6315, g6336, g6307, g6255, g6351, g6377, g6259, g6299, g6329, g6267, g6395, g6322, g6251, g6239, g6271, g6365, g6247, g6346, g6279, g6263, g6373, g6295, g6235, g6287, g6369, g6303, g6243, g6275, g6358, g6291, g6283, n3126 );
input g35, g6311, g4826, g4688, g4801, g4793, g4776, g4653, g4669, g4659, g4709, g4785, g4765, g6381, g6315, g6336, g6307, g6255, g6351, g6377, g6259, g6299, g6329, g6267, g6395, g6322, g6251, g6239, g6271, g6365, g6247, g6346, g6279, g6263, g6373, g6295, g6235, g6287, g6369, g6303, g6243, g6275, g6358, g6291, g6283;
output n3126;
wire n7920, n5907, n6569, n4967, n4721, n5906, n6568, n6535, n6550_1, n6558, n4720, n4723, n4815, n4818, n5905, n6560_1, n6563, n6567, n6530, n6534, n6543, n6546_1, n6549, n6557, n6552, n6554, n6559, n6561, n6532, n6562, n6564, n6565_1, n6566, n6526_1, n6528, n6529, n6531_1, n6533, n6542, n6537, n6538, n6540, n6544, n6545, n6547, n6548, n6555_1, n6556, n6551, n5196_1, n6553, n6277, n6527, n6539, n6279, n6541_1, n6536_1;
MX2X1    g3274(.A(g6311), .B(n7920), .S0(g35), .Y(n3126));
MX2X1    g3273(.A(g4826), .B(n6569), .S0(n5907), .Y(n7920));
AOI21X1  g1267(.A0(n5906), .A1(n4721), .B0(n4967), .Y(n5907));
NAND4X1  g1929(.A(n6558), .B(n6550_1), .C(n6535), .D(n6568), .Y(n6569));
INVX1    g0347(.A(g4688), .Y(n4967));
NOR3X1   g0101(.A(g4793), .B(g4801), .C(n4720), .Y(n4721));
NOR4X1   g1266(.A(n5905), .B(n4818), .C(n4815), .D(n4723), .Y(n5906));
NOR3X1   g1928(.A(n6567), .B(n6563), .C(n6560_1), .Y(n6568));
NOR2X1   g1895(.A(n6534), .B(n6530), .Y(n6535));
NOR3X1   g1910(.A(n6549), .B(n6546_1), .C(n6543), .Y(n6550_1));
AOI21X1  g1918(.A0(n6554), .A1(n6552), .B0(n6557), .Y(n6558));
INVX1    g0100(.A(g4776), .Y(n4720));
NAND3X1  g0103(.A(g4659), .B(g4669), .C(g4653), .Y(n4723));
INVX1    g0195(.A(g4709), .Y(n4815));
INVX1    g0198(.A(g4785), .Y(n4818));
INVX1    g1265(.A(g4765), .Y(n5905));
NOR2X1   g1920(.A(n6559), .B(n6552), .Y(n6560_1));
OAI21X1  g1923(.A0(n6562), .A1(n6532), .B0(n6561), .Y(n6563));
AOI21X1  g1927(.A0(n6566), .A1(n6565_1), .B0(n6564), .Y(n6567));
AOI21X1  g1890(.A0(n6529), .A1(n6528), .B0(n6526_1), .Y(n6530));
OAI21X1  g1894(.A0(n6533), .A1(n6532), .B0(n6531_1), .Y(n6534));
NAND4X1  g1903(.A(n6540), .B(n6538), .C(n6537), .D(n6542), .Y(n6543));
OAI21X1  g1906(.A0(n6545), .A1(n6526_1), .B0(n6544), .Y(n6546_1));
NAND2X1  g1909(.A(n6548), .B(n6547), .Y(n6549));
AOI21X1  g1917(.A0(n6556), .A1(n6555_1), .B0(n6552), .Y(n6557));
XOR2X1   g1912(.A(g6381), .B(n6551), .Y(n6552));
AND2X1   g1914(.A(n6553), .B(n5196_1), .Y(n6554));
NAND4X1  g1919(.A(g6307), .B(n6277), .C(g6336), .D(g6315), .Y(n6559));
NAND4X1  g1921(.A(n6527), .B(g6351), .C(g6255), .D(n5196_1), .Y(n6561));
NAND2X1  g1892(.A(n6277), .B(g6336), .Y(n6532));
NAND3X1  g1922(.A(n6527), .B(g6259), .C(g6377), .Y(n6562));
INVX1    g1924(.A(n6552), .Y(n6564));
NAND3X1  g1925(.A(n6539), .B(g6299), .C(g6315), .Y(n6565_1));
NAND4X1  g1926(.A(g6267), .B(n6277), .C(g6336), .D(g6329), .Y(n6566));
NAND2X1  g1886(.A(g6395), .B(n6279), .Y(n6526_1));
NAND3X1  g1888(.A(n6527), .B(g6251), .C(g6322), .Y(n6528));
NAND3X1  g1889(.A(g6381), .B(g6351), .C(g6239), .Y(n6529));
NAND4X1  g1891(.A(n6527), .B(g6365), .C(g6271), .D(n5196_1), .Y(n6531_1));
NAND3X1  g1893(.A(g6346), .B(n6527), .C(g6247), .Y(n6533));
NAND4X1  g1902(.A(g6279), .B(n6277), .C(g6336), .D(n6541_1), .Y(n6542));
NAND4X1  g1897(.A(g6263), .B(g6395), .C(n6279), .D(n6536_1), .Y(n6537));
NAND4X1  g1898(.A(g6295), .B(g6381), .C(g6373), .D(n5196_1), .Y(n6538));
NAND4X1  g1900(.A(g6346), .B(g6381), .C(g6235), .D(n6539), .Y(n6540));
NAND4X1  g1904(.A(n6527), .B(g6369), .C(g6287), .D(n6539), .Y(n6544));
NAND3X1  g1905(.A(g6303), .B(n6527), .C(g6373), .Y(n6545));
NAND4X1  g1907(.A(g6381), .B(g6243), .C(g6377), .D(n6539), .Y(n6547));
NAND4X1  g1908(.A(g6381), .B(g6311), .C(g6322), .D(n5196_1), .Y(n6548));
NAND3X1  g1915(.A(n6539), .B(g6275), .C(g6329), .Y(n6555_1));
NAND4X1  g1916(.A(g6395), .B(n6279), .C(g6291), .D(g6358), .Y(n6556));
INVX1    g1911(.A(g6351), .Y(n6551));
AND2X1   g0563(.A(g6395), .B(g6336), .Y(n5196_1));
AND2X1   g1913(.A(g6283), .B(g6358), .Y(n6553));
INVX1    g1637(.A(g6395), .Y(n6277));
INVX1    g1887(.A(g6381), .Y(n6527));
NOR2X1   g1899(.A(g6395), .B(g6336), .Y(n6539));
INVX1    g1639(.A(g6336), .Y(n6279));
AND2X1   g1901(.A(g6381), .B(g6369), .Y(n6541_1));
AND2X1   g1896(.A(g6381), .B(g6365), .Y(n6536_1));

endmodule
