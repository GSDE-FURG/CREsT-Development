// Benchmark "b04_C" written by ABC on Wed Aug 05 14:36:50 2020

module b04_C ( 
    RESTART, AVERAGE, ENABLE, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_,
    DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_,
    STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN,
    DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_2__SCAN_IN,
    DATA_OUT_REG_3__SCAN_IN, DATA_OUT_REG_4__SCAN_IN,
    DATA_OUT_REG_5__SCAN_IN, DATA_OUT_REG_6__SCAN_IN,
    DATA_OUT_REG_7__SCAN_IN, REG4_REG_0__SCAN_IN, REG4_REG_1__SCAN_IN,
    REG4_REG_2__SCAN_IN, RMAX_REG_7__SCAN_IN, RMAX_REG_6__SCAN_IN,
    RMAX_REG_5__SCAN_IN, RMAX_REG_4__SCAN_IN, RMAX_REG_3__SCAN_IN,
    RMAX_REG_2__SCAN_IN, RMAX_REG_1__SCAN_IN, RMAX_REG_0__SCAN_IN,
    RMIN_REG_7__SCAN_IN, RMIN_REG_6__SCAN_IN, RMIN_REG_5__SCAN_IN,
    RMIN_REG_4__SCAN_IN, RMIN_REG_3__SCAN_IN, RMIN_REG_2__SCAN_IN,
    RMIN_REG_1__SCAN_IN, RMIN_REG_0__SCAN_IN, RLAST_REG_7__SCAN_IN,
    RLAST_REG_6__SCAN_IN, RLAST_REG_5__SCAN_IN, RLAST_REG_4__SCAN_IN,
    RLAST_REG_3__SCAN_IN, RLAST_REG_2__SCAN_IN, RLAST_REG_1__SCAN_IN,
    RLAST_REG_0__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_6__SCAN_IN,
    REG1_REG_5__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_3__SCAN_IN,
    REG1_REG_2__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_0__SCAN_IN,
    REG2_REG_7__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_5__SCAN_IN,
    REG2_REG_4__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_2__SCAN_IN,
    REG2_REG_1__SCAN_IN, REG2_REG_0__SCAN_IN, REG3_REG_7__SCAN_IN,
    REG3_REG_6__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_4__SCAN_IN,
    REG3_REG_3__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_1__SCAN_IN,
    REG3_REG_0__SCAN_IN, REG4_REG_7__SCAN_IN, REG4_REG_6__SCAN_IN,
    REG4_REG_5__SCAN_IN, REG4_REG_4__SCAN_IN, REG4_REG_3__SCAN_IN,
    U344, U343, U342, U341, U340, U339, U338, U337, U336, U335, U334, U333,
    U332, U331, U330, U329, U328, U327, U326, U325, U324, U323, U322, U321,
    U320, U319, U318, U317, U316, U315, U314, U313, U312, U311, U310, U309,
    U308, U307, U306, U305, U304, U303, U302, U301, U300, U299, U298, U297,
    U296, U295, U294, U293, U292, U291, U290, U289, U288, U287, U286, U285,
    U284, U283, U282, U281, U280, U375  );
  input  RESTART, AVERAGE, ENABLE, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_,
    DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_,
    STATO_REG_0__SCAN_IN, STATO_REG_1__SCAN_IN, DATA_OUT_REG_0__SCAN_IN,
    DATA_OUT_REG_1__SCAN_IN, DATA_OUT_REG_2__SCAN_IN,
    DATA_OUT_REG_3__SCAN_IN, DATA_OUT_REG_4__SCAN_IN,
    DATA_OUT_REG_5__SCAN_IN, DATA_OUT_REG_6__SCAN_IN,
    DATA_OUT_REG_7__SCAN_IN, REG4_REG_0__SCAN_IN, REG4_REG_1__SCAN_IN,
    REG4_REG_2__SCAN_IN, RMAX_REG_7__SCAN_IN, RMAX_REG_6__SCAN_IN,
    RMAX_REG_5__SCAN_IN, RMAX_REG_4__SCAN_IN, RMAX_REG_3__SCAN_IN,
    RMAX_REG_2__SCAN_IN, RMAX_REG_1__SCAN_IN, RMAX_REG_0__SCAN_IN,
    RMIN_REG_7__SCAN_IN, RMIN_REG_6__SCAN_IN, RMIN_REG_5__SCAN_IN,
    RMIN_REG_4__SCAN_IN, RMIN_REG_3__SCAN_IN, RMIN_REG_2__SCAN_IN,
    RMIN_REG_1__SCAN_IN, RMIN_REG_0__SCAN_IN, RLAST_REG_7__SCAN_IN,
    RLAST_REG_6__SCAN_IN, RLAST_REG_5__SCAN_IN, RLAST_REG_4__SCAN_IN,
    RLAST_REG_3__SCAN_IN, RLAST_REG_2__SCAN_IN, RLAST_REG_1__SCAN_IN,
    RLAST_REG_0__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_6__SCAN_IN,
    REG1_REG_5__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_3__SCAN_IN,
    REG1_REG_2__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_0__SCAN_IN,
    REG2_REG_7__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_5__SCAN_IN,
    REG2_REG_4__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_2__SCAN_IN,
    REG2_REG_1__SCAN_IN, REG2_REG_0__SCAN_IN, REG3_REG_7__SCAN_IN,
    REG3_REG_6__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_4__SCAN_IN,
    REG3_REG_3__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_1__SCAN_IN,
    REG3_REG_0__SCAN_IN, REG4_REG_7__SCAN_IN, REG4_REG_6__SCAN_IN,
    REG4_REG_5__SCAN_IN, REG4_REG_4__SCAN_IN, REG4_REG_3__SCAN_IN;
  output U344, U343, U342, U341, U340, U339, U338, U337, U336, U335, U334,
    U333, U332, U331, U330, U329, U328, U327, U326, U325, U324, U323, U322,
    U321, U320, U319, U318, U317, U316, U315, U314, U313, U312, U311, U310,
    U309, U308, U307, U306, U305, U304, U303, U302, U301, U300, U299, U298,
    U297, U296, U295, U294, U293, U292, U291, U290, U289, U288, U287, U286,
    U285, U284, U283, U282, U281, U280, U375;
  wire n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
    n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
    n174, n175, n176, n177, n178, n179, n180, n181, n187, n189, n191, n193,
    n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
    n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
    n226, n228, n229, n230, n231, n233, n235, n237, n239, n241, n243, n245,
    n247, n248, n249, n252, n254, n256, n258, n260, n262, n264, n266, n268,
    n270, n272, n274, n276, n278, n280, n282, n284, n286, n288, n290, n292,
    n294, n296, n298, n300, n302, n304, n306, n308, n310, n312, n314, n315,
    n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
    n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
    n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
    n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
    n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
    n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
    n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
    n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
    n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
    n424, n425, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
    n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
    n449, n450, n452, n453, n454, n455, n456, n457, n458, n459, n461, n462,
    n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n474, n475,
    n476, n477, n478, n479, n481, n482, n483, n484, n485, n486, n487, n488,
    n490, n491, n492, n493, n494, n495, n497, n498, n499, n500, n501, n502,
    n504, n505, n506, n507, n508, n509;
  INVX1   g000(.A(DATA_IN_7_), .Y(n151));
  INVX1   g001(.A(RMAX_REG_7__SCAN_IN), .Y(n152));
  INVX1   g002(.A(DATA_IN_1_), .Y(n153));
  INVX1   g003(.A(RMAX_REG_0__SCAN_IN), .Y(n154));
  NAND2X1 g004(.A(n154), .B(DATA_IN_0_), .Y(n155));
  AOI21X1 g005(.A0(RMAX_REG_1__SCAN_IN), .A1(n153), .B0(n155), .Y(n156));
  INVX1   g006(.A(DATA_IN_2_), .Y(n157));
  OAI22X1 g007(.A0(RMAX_REG_2__SCAN_IN), .A1(n157), .B0(n153), .B1(RMAX_REG_1__SCAN_IN), .Y(n158));
  INVX1   g008(.A(DATA_IN_3_), .Y(n159));
  AOI22X1 g009(.A0(RMAX_REG_3__SCAN_IN), .A1(n159), .B0(n157), .B1(RMAX_REG_2__SCAN_IN), .Y(n160));
  OAI21X1 g010(.A0(n158), .A1(n156), .B0(n160), .Y(n161));
  INVX1   g011(.A(RMAX_REG_4__SCAN_IN), .Y(n162));
  INVX1   g012(.A(RMAX_REG_3__SCAN_IN), .Y(n163));
  AOI22X1 g013(.A0(n162), .A1(DATA_IN_4_), .B0(DATA_IN_3_), .B1(n163), .Y(n164));
  NAND2X1 g014(.A(n164), .B(n161), .Y(n165));
  INVX1   g015(.A(DATA_IN_5_), .Y(n166));
  INVX1   g016(.A(DATA_IN_4_), .Y(n167));
  AOI22X1 g017(.A0(RMAX_REG_5__SCAN_IN), .A1(n166), .B0(n167), .B1(RMAX_REG_4__SCAN_IN), .Y(n168));
  NAND2X1 g018(.A(n168), .B(n165), .Y(n169));
  INVX1   g019(.A(RMAX_REG_6__SCAN_IN), .Y(n170));
  INVX1   g020(.A(RMAX_REG_5__SCAN_IN), .Y(n171));
  AOI22X1 g021(.A0(n170), .A1(DATA_IN_6_), .B0(DATA_IN_5_), .B1(n171), .Y(n172));
  NAND2X1 g022(.A(n172), .B(n169), .Y(n173));
  INVX1   g023(.A(DATA_IN_6_), .Y(n174));
  AOI22X1 g024(.A0(n152), .A1(DATA_IN_7_), .B0(n174), .B1(RMAX_REG_6__SCAN_IN), .Y(n175));
  AOI22X1 g025(.A0(n173), .A1(n175), .B0(RMAX_REG_7__SCAN_IN), .B1(n151), .Y(n176));
  INVX1   g026(.A(n176), .Y(n177));
  AOI21X1 g027(.A0(n177), .A1(STATO_REG_1__SCAN_IN), .B0(STATO_REG_0__SCAN_IN), .Y(n178));
  INVX1   g028(.A(STATO_REG_0__SCAN_IN), .Y(n179));
  INVX1   g029(.A(STATO_REG_1__SCAN_IN), .Y(n180));
  OAI21X1 g030(.A0(n176), .A1(n180), .B0(n179), .Y(n181));
  OAI22X1 g031(.A0(n178), .A1(n151), .B0(n152), .B1(n181), .Y(U344));
  OAI22X1 g032(.A0(n178), .A1(n174), .B0(n170), .B1(n181), .Y(U343));
  OAI22X1 g033(.A0(n178), .A1(n166), .B0(n171), .B1(n181), .Y(U342));
  OAI22X1 g034(.A0(n178), .A1(n167), .B0(n162), .B1(n181), .Y(U341));
  OAI22X1 g035(.A0(n178), .A1(n159), .B0(n163), .B1(n181), .Y(U340));
  INVX1   g036(.A(RMAX_REG_2__SCAN_IN), .Y(n187));
  OAI22X1 g037(.A0(n178), .A1(n157), .B0(n187), .B1(n181), .Y(U339));
  INVX1   g038(.A(RMAX_REG_1__SCAN_IN), .Y(n189));
  OAI22X1 g039(.A0(n178), .A1(n153), .B0(n189), .B1(n181), .Y(U338));
  INVX1   g040(.A(DATA_IN_0_), .Y(n191));
  OAI22X1 g041(.A0(n178), .A1(n191), .B0(n154), .B1(n181), .Y(U337));
  INVX1   g042(.A(RMIN_REG_7__SCAN_IN), .Y(n193));
  NOR2X1  g043(.A(STATO_REG_1__SCAN_IN), .B(STATO_REG_0__SCAN_IN), .Y(U375));
  INVX1   g044(.A(RMIN_REG_1__SCAN_IN), .Y(n195));
  NAND2X1 g045(.A(RMIN_REG_0__SCAN_IN), .B(n191), .Y(n196));
  AOI21X1 g046(.A0(n195), .A1(DATA_IN_1_), .B0(n196), .Y(n197));
  INVX1   g047(.A(RMIN_REG_2__SCAN_IN), .Y(n198));
  OAI22X1 g048(.A0(n198), .A1(DATA_IN_2_), .B0(DATA_IN_1_), .B1(n195), .Y(n199));
  INVX1   g049(.A(RMIN_REG_3__SCAN_IN), .Y(n200));
  AOI22X1 g050(.A0(n200), .A1(DATA_IN_3_), .B0(DATA_IN_2_), .B1(n198), .Y(n201));
  OAI21X1 g051(.A0(n199), .A1(n197), .B0(n201), .Y(n202));
  AOI22X1 g052(.A0(RMIN_REG_4__SCAN_IN), .A1(n167), .B0(n159), .B1(RMIN_REG_3__SCAN_IN), .Y(n203));
  NAND2X1 g053(.A(n203), .B(n202), .Y(n204));
  INVX1   g054(.A(RMIN_REG_5__SCAN_IN), .Y(n205));
  INVX1   g055(.A(RMIN_REG_4__SCAN_IN), .Y(n206));
  AOI22X1 g056(.A0(n205), .A1(DATA_IN_5_), .B0(DATA_IN_4_), .B1(n206), .Y(n207));
  NAND2X1 g057(.A(n207), .B(n204), .Y(n208));
  AOI22X1 g058(.A0(RMIN_REG_6__SCAN_IN), .A1(n174), .B0(n166), .B1(RMIN_REG_5__SCAN_IN), .Y(n209));
  NAND2X1 g059(.A(n209), .B(n208), .Y(n210));
  INVX1   g060(.A(RMIN_REG_6__SCAN_IN), .Y(n211));
  AOI22X1 g061(.A0(RMIN_REG_7__SCAN_IN), .A1(n151), .B0(DATA_IN_6_), .B1(n211), .Y(n212));
  AOI22X1 g062(.A0(n210), .A1(n212), .B0(n193), .B1(DATA_IN_7_), .Y(n213));
  INVX1   g063(.A(n213), .Y(n214));
  AOI21X1 g064(.A0(n214), .A1(n176), .B0(STATO_REG_0__SCAN_IN), .Y(n215));
  NOR2X1  g065(.A(n215), .B(U375), .Y(n216));
  NOR3X1  g066(.A(n213), .B(n177), .C(n180), .Y(n217));
  NOR2X1  g067(.A(n217), .B(STATO_REG_0__SCAN_IN), .Y(n218));
  OAI22X1 g068(.A0(n216), .A1(n193), .B0(n151), .B1(n218), .Y(U336));
  OAI22X1 g069(.A0(n216), .A1(n211), .B0(n174), .B1(n218), .Y(U335));
  OAI22X1 g070(.A0(n216), .A1(n205), .B0(n166), .B1(n218), .Y(U334));
  OAI22X1 g071(.A0(n216), .A1(n206), .B0(n167), .B1(n218), .Y(U333));
  OAI22X1 g072(.A0(n216), .A1(n200), .B0(n159), .B1(n218), .Y(U332));
  OAI22X1 g073(.A0(n216), .A1(n198), .B0(n157), .B1(n218), .Y(U331));
  OAI22X1 g074(.A0(n216), .A1(n195), .B0(n153), .B1(n218), .Y(U330));
  OAI21X1 g075(.A0(n215), .A1(U375), .B0(RMIN_REG_0__SCAN_IN), .Y(n226));
  OAI21X1 g076(.A0(n218), .A1(n191), .B0(n226), .Y(U329));
  INVX1   g077(.A(RLAST_REG_7__SCAN_IN), .Y(n228));
  INVX1   g078(.A(ENABLE), .Y(n229));
  OAI21X1 g079(.A0(n180), .A1(n229), .B0(n179), .Y(n230));
  OAI21X1 g080(.A0(STATO_REG_0__SCAN_IN), .A1(ENABLE), .B0(STATO_REG_1__SCAN_IN), .Y(n231));
  OAI22X1 g081(.A0(n230), .A1(n228), .B0(n151), .B1(n231), .Y(U328));
  INVX1   g082(.A(RLAST_REG_6__SCAN_IN), .Y(n233));
  OAI22X1 g083(.A0(n230), .A1(n233), .B0(n174), .B1(n231), .Y(U327));
  INVX1   g084(.A(RLAST_REG_5__SCAN_IN), .Y(n235));
  OAI22X1 g085(.A0(n230), .A1(n235), .B0(n166), .B1(n231), .Y(U326));
  INVX1   g086(.A(RLAST_REG_4__SCAN_IN), .Y(n237));
  OAI22X1 g087(.A0(n230), .A1(n237), .B0(n167), .B1(n231), .Y(U325));
  INVX1   g088(.A(RLAST_REG_3__SCAN_IN), .Y(n239));
  OAI22X1 g089(.A0(n230), .A1(n239), .B0(n159), .B1(n231), .Y(U324));
  INVX1   g090(.A(RLAST_REG_2__SCAN_IN), .Y(n241));
  OAI22X1 g091(.A0(n230), .A1(n241), .B0(n157), .B1(n231), .Y(U323));
  INVX1   g092(.A(RLAST_REG_1__SCAN_IN), .Y(n243));
  OAI22X1 g093(.A0(n230), .A1(n243), .B0(n153), .B1(n231), .Y(U322));
  INVX1   g094(.A(RLAST_REG_0__SCAN_IN), .Y(n245));
  OAI22X1 g095(.A0(n230), .A1(n245), .B0(n191), .B1(n231), .Y(U321));
  INVX1   g096(.A(REG1_REG_7__SCAN_IN), .Y(n247));
  NAND2X1 g097(.A(STATO_REG_1__SCAN_IN), .B(n179), .Y(n248));
  XOR2X1  g098(.A(STATO_REG_1__SCAN_IN), .B(n179), .Y(n249));
  INVX1   g099(.A(n249), .Y(U280));
  OAI22X1 g100(.A0(n248), .A1(n151), .B0(n247), .B1(U280), .Y(U320));
  INVX1   g101(.A(REG1_REG_6__SCAN_IN), .Y(n252));
  OAI22X1 g102(.A0(n248), .A1(n174), .B0(n252), .B1(U280), .Y(U319));
  INVX1   g103(.A(REG1_REG_5__SCAN_IN), .Y(n254));
  OAI22X1 g104(.A0(n248), .A1(n166), .B0(n254), .B1(U280), .Y(U318));
  INVX1   g105(.A(REG1_REG_4__SCAN_IN), .Y(n256));
  OAI22X1 g106(.A0(n248), .A1(n167), .B0(n256), .B1(U280), .Y(U317));
  INVX1   g107(.A(REG1_REG_3__SCAN_IN), .Y(n258));
  OAI22X1 g108(.A0(n248), .A1(n159), .B0(n258), .B1(U280), .Y(U316));
  INVX1   g109(.A(REG1_REG_2__SCAN_IN), .Y(n260));
  OAI22X1 g110(.A0(n248), .A1(n157), .B0(n260), .B1(U280), .Y(U315));
  INVX1   g111(.A(REG1_REG_1__SCAN_IN), .Y(n262));
  OAI22X1 g112(.A0(n248), .A1(n153), .B0(n262), .B1(U280), .Y(U314));
  INVX1   g113(.A(REG1_REG_0__SCAN_IN), .Y(n264));
  OAI22X1 g114(.A0(n248), .A1(n191), .B0(n264), .B1(U280), .Y(U313));
  INVX1   g115(.A(REG2_REG_7__SCAN_IN), .Y(n266));
  OAI22X1 g116(.A0(n248), .A1(n247), .B0(n266), .B1(U280), .Y(U312));
  INVX1   g117(.A(REG2_REG_6__SCAN_IN), .Y(n268));
  OAI22X1 g118(.A0(n248), .A1(n252), .B0(n268), .B1(U280), .Y(U311));
  INVX1   g119(.A(REG2_REG_5__SCAN_IN), .Y(n270));
  OAI22X1 g120(.A0(n248), .A1(n254), .B0(n270), .B1(U280), .Y(U310));
  INVX1   g121(.A(REG2_REG_4__SCAN_IN), .Y(n272));
  OAI22X1 g122(.A0(n248), .A1(n256), .B0(n272), .B1(U280), .Y(U309));
  INVX1   g123(.A(REG2_REG_3__SCAN_IN), .Y(n274));
  OAI22X1 g124(.A0(n248), .A1(n258), .B0(n274), .B1(U280), .Y(U308));
  INVX1   g125(.A(REG2_REG_2__SCAN_IN), .Y(n276));
  OAI22X1 g126(.A0(n248), .A1(n260), .B0(n276), .B1(U280), .Y(U307));
  INVX1   g127(.A(REG2_REG_1__SCAN_IN), .Y(n278));
  OAI22X1 g128(.A0(n248), .A1(n262), .B0(n278), .B1(U280), .Y(U306));
  INVX1   g129(.A(REG2_REG_0__SCAN_IN), .Y(n280));
  OAI22X1 g130(.A0(n248), .A1(n264), .B0(n280), .B1(U280), .Y(U305));
  INVX1   g131(.A(REG3_REG_7__SCAN_IN), .Y(n282));
  OAI22X1 g132(.A0(n248), .A1(n266), .B0(n282), .B1(U280), .Y(U304));
  INVX1   g133(.A(REG3_REG_6__SCAN_IN), .Y(n284));
  OAI22X1 g134(.A0(n248), .A1(n268), .B0(n284), .B1(U280), .Y(U303));
  INVX1   g135(.A(REG3_REG_5__SCAN_IN), .Y(n286));
  OAI22X1 g136(.A0(n248), .A1(n270), .B0(n286), .B1(U280), .Y(U302));
  INVX1   g137(.A(REG3_REG_4__SCAN_IN), .Y(n288));
  OAI22X1 g138(.A0(n248), .A1(n272), .B0(n288), .B1(U280), .Y(U301));
  INVX1   g139(.A(REG3_REG_3__SCAN_IN), .Y(n290));
  OAI22X1 g140(.A0(n248), .A1(n274), .B0(n290), .B1(U280), .Y(U300));
  INVX1   g141(.A(REG3_REG_2__SCAN_IN), .Y(n292));
  OAI22X1 g142(.A0(n248), .A1(n276), .B0(n292), .B1(U280), .Y(U299));
  INVX1   g143(.A(REG3_REG_1__SCAN_IN), .Y(n294));
  OAI22X1 g144(.A0(n248), .A1(n278), .B0(n294), .B1(U280), .Y(U298));
  INVX1   g145(.A(REG3_REG_0__SCAN_IN), .Y(n296));
  OAI22X1 g146(.A0(n248), .A1(n280), .B0(n296), .B1(U280), .Y(U297));
  INVX1   g147(.A(REG4_REG_7__SCAN_IN), .Y(n298));
  OAI22X1 g148(.A0(n248), .A1(n282), .B0(n298), .B1(U280), .Y(U296));
  INVX1   g149(.A(REG4_REG_6__SCAN_IN), .Y(n300));
  OAI22X1 g150(.A0(n248), .A1(n284), .B0(n300), .B1(U280), .Y(U295));
  INVX1   g151(.A(REG4_REG_5__SCAN_IN), .Y(n302));
  OAI22X1 g152(.A0(n248), .A1(n286), .B0(n302), .B1(U280), .Y(U294));
  INVX1   g153(.A(REG4_REG_4__SCAN_IN), .Y(n304));
  OAI22X1 g154(.A0(n248), .A1(n288), .B0(n304), .B1(U280), .Y(U293));
  INVX1   g155(.A(REG4_REG_3__SCAN_IN), .Y(n306));
  OAI22X1 g156(.A0(n248), .A1(n290), .B0(n306), .B1(U280), .Y(U292));
  INVX1   g157(.A(REG4_REG_2__SCAN_IN), .Y(n308));
  OAI22X1 g158(.A0(n248), .A1(n292), .B0(n308), .B1(U280), .Y(U291));
  INVX1   g159(.A(REG4_REG_1__SCAN_IN), .Y(n310));
  OAI22X1 g160(.A0(n248), .A1(n294), .B0(n310), .B1(U280), .Y(U290));
  INVX1   g161(.A(REG4_REG_0__SCAN_IN), .Y(n312));
  OAI22X1 g162(.A0(n248), .A1(n296), .B0(n312), .B1(U280), .Y(U289));
  NAND2X1 g163(.A(RMAX_REG_1__SCAN_IN), .B(RESTART), .Y(n314));
  OAI21X1 g164(.A0(n153), .A1(RESTART), .B0(n314), .Y(n315));
  NAND2X1 g165(.A(RMIN_REG_0__SCAN_IN), .B(RESTART), .Y(n316));
  OAI21X1 g166(.A0(n312), .A1(RESTART), .B0(n316), .Y(n317));
  NAND2X1 g167(.A(RMAX_REG_0__SCAN_IN), .B(RESTART), .Y(n318));
  OAI21X1 g168(.A0(n191), .A1(RESTART), .B0(n318), .Y(n319));
  NAND3X1 g169(.A(n319), .B(n317), .C(n315), .Y(n320));
  NOR2X1  g170(.A(n310), .B(RESTART), .Y(n321));
  AOI21X1 g171(.A0(RMIN_REG_1__SCAN_IN), .A1(RESTART), .B0(n321), .Y(n322));
  AOI21X1 g172(.A0(n319), .A1(n317), .B0(n315), .Y(n323));
  OAI21X1 g173(.A0(n323), .A1(n322), .B0(n320), .Y(n324));
  NAND2X1 g174(.A(RMAX_REG_2__SCAN_IN), .B(RESTART), .Y(n325));
  OAI21X1 g175(.A0(n157), .A1(RESTART), .B0(n325), .Y(n326));
  NOR2X1  g176(.A(n308), .B(RESTART), .Y(n327));
  AOI21X1 g177(.A0(RMIN_REG_2__SCAN_IN), .A1(RESTART), .B0(n327), .Y(n328));
  XOR2X1  g178(.A(n328), .B(n326), .Y(n329));
  XOR2X1  g179(.A(n329), .B(n324), .Y(n330));
  INVX1   g180(.A(n315), .Y(n331));
  INVX1   g181(.A(RESTART), .Y(n332));
  NAND2X1 g182(.A(REG4_REG_0__SCAN_IN), .B(n332), .Y(n333));
  NAND2X1 g183(.A(DATA_IN_0_), .B(n332), .Y(n334));
  AOI22X1 g184(.A0(n318), .A1(n334), .B0(n333), .B1(n316), .Y(n335));
  NAND2X1 g185(.A(RMIN_REG_1__SCAN_IN), .B(RESTART), .Y(n336));
  OAI21X1 g186(.A0(n310), .A1(RESTART), .B0(n336), .Y(n337));
  XOR2X1  g187(.A(n337), .B(n335), .Y(n338));
  NAND2X1 g188(.A(REG4_REG_1__SCAN_IN), .B(n332), .Y(n339));
  NAND3X1 g189(.A(n339), .B(n336), .C(n315), .Y(n340));
  OAI22X1 g190(.A0(n322), .A1(n320), .B0(n335), .B1(n340), .Y(n341));
  AOI21X1 g191(.A0(n338), .A1(n331), .B0(n341), .Y(n342));
  INVX1   g192(.A(n319), .Y(n343));
  XOR2X1  g193(.A(n343), .B(n317), .Y(n344));
  NAND3X1 g194(.A(n344), .B(n342), .C(n330), .Y(n345));
  NOR2X1  g195(.A(n157), .B(RESTART), .Y(n346));
  AOI21X1 g196(.A0(RMAX_REG_2__SCAN_IN), .A1(RESTART), .B0(n346), .Y(n347));
  NOR2X1  g197(.A(n328), .B(n347), .Y(n348));
  NAND2X1 g198(.A(n328), .B(n347), .Y(n349));
  AOI21X1 g199(.A0(n349), .A1(n324), .B0(n348), .Y(n350));
  NAND2X1 g200(.A(RMAX_REG_3__SCAN_IN), .B(RESTART), .Y(n351));
  OAI21X1 g201(.A0(n159), .A1(RESTART), .B0(n351), .Y(n352));
  NAND2X1 g202(.A(RMIN_REG_3__SCAN_IN), .B(RESTART), .Y(n353));
  OAI21X1 g203(.A0(n306), .A1(RESTART), .B0(n353), .Y(n354));
  INVX1   g204(.A(n354), .Y(n355));
  XOR2X1  g205(.A(n355), .B(n352), .Y(n356));
  XOR2X1  g206(.A(n356), .B(n350), .Y(n357));
  NOR2X1  g207(.A(n357), .B(n345), .Y(n358));
  NAND2X1 g208(.A(n354), .B(n352), .Y(n359));
  NOR2X1  g209(.A(n354), .B(n352), .Y(n360));
  OAI21X1 g210(.A0(n360), .A1(n350), .B0(n359), .Y(n361));
  NOR2X1  g211(.A(n167), .B(RESTART), .Y(n362));
  AOI21X1 g212(.A0(RMAX_REG_4__SCAN_IN), .A1(RESTART), .B0(n362), .Y(n363));
  NOR2X1  g213(.A(n304), .B(RESTART), .Y(n364));
  AOI21X1 g214(.A0(RMIN_REG_4__SCAN_IN), .A1(RESTART), .B0(n364), .Y(n365));
  XOR2X1  g215(.A(n365), .B(n363), .Y(n366));
  INVX1   g216(.A(n366), .Y(n367));
  XOR2X1  g217(.A(n367), .B(n361), .Y(n368));
  NAND2X1 g218(.A(n368), .B(n358), .Y(n369));
  NAND2X1 g219(.A(RMAX_REG_5__SCAN_IN), .B(RESTART), .Y(n370));
  OAI21X1 g220(.A0(n166), .A1(RESTART), .B0(n370), .Y(n371));
  NOR2X1  g221(.A(n302), .B(RESTART), .Y(n372));
  AOI21X1 g222(.A0(RMIN_REG_5__SCAN_IN), .A1(RESTART), .B0(n372), .Y(n373));
  XOR2X1  g223(.A(n373), .B(n371), .Y(n374));
  NOR2X1  g224(.A(n365), .B(n363), .Y(n375));
  NAND2X1 g225(.A(n365), .B(n363), .Y(n376));
  AOI21X1 g226(.A0(n376), .A1(n361), .B0(n375), .Y(n377));
  XOR2X1  g227(.A(n377), .B(n374), .Y(n378));
  INVX1   g228(.A(n373), .Y(n379));
  NAND2X1 g229(.A(n379), .B(n371), .Y(n380));
  NAND2X1 g230(.A(RMAX_REG_6__SCAN_IN), .B(RESTART), .Y(n381));
  OAI21X1 g231(.A0(n174), .A1(RESTART), .B0(n381), .Y(n382));
  NAND2X1 g232(.A(RMIN_REG_6__SCAN_IN), .B(RESTART), .Y(n383));
  OAI21X1 g233(.A0(n300), .A1(RESTART), .B0(n383), .Y(n384));
  XOR2X1  g234(.A(n384), .B(n382), .Y(n385));
  OAI21X1 g235(.A0(n379), .A1(n371), .B0(n385), .Y(n386));
  AOI21X1 g236(.A0(n380), .A1(n377), .B0(n386), .Y(n387));
  OAI21X1 g237(.A0(n335), .A1(n315), .B0(n337), .Y(n388));
  AOI22X1 g238(.A0(n347), .A1(n328), .B0(n388), .B1(n320), .Y(n389));
  OAI22X1 g239(.A0(n352), .A1(n354), .B0(n389), .B1(n348), .Y(n390));
  AOI22X1 g240(.A0(n363), .A1(n365), .B0(n390), .B1(n359), .Y(n391));
  OAI22X1 g241(.A0(n375), .A1(n391), .B0(n379), .B1(n371), .Y(n392));
  NAND2X1 g242(.A(DATA_IN_5_), .B(n332), .Y(n393));
  AOI21X1 g243(.A0(n393), .A1(n370), .B0(n373), .Y(n394));
  NOR2X1  g244(.A(n385), .B(n394), .Y(n395));
  AOI21X1 g245(.A0(n395), .A1(n392), .B0(n387), .Y(n396));
  XOR2X1  g246(.A(n378), .B(n369), .Y(n397));
  XOR2X1  g247(.A(n328), .B(n347), .Y(n398));
  XOR2X1  g248(.A(n398), .B(n324), .Y(n399));
  NAND2X1 g249(.A(n344), .B(n342), .Y(n400));
  NOR2X1  g250(.A(n400), .B(n399), .Y(n401));
  XOR2X1  g251(.A(n357), .B(n401), .Y(n402));
  XOR2X1  g252(.A(n400), .B(n330), .Y(n403));
  INVX1   g253(.A(n342), .Y(n404));
  XOR2X1  g254(.A(n344), .B(n404), .Y(n405));
  XOR2X1  g255(.A(n366), .B(n361), .Y(n406));
  XOR2X1  g256(.A(n406), .B(n358), .Y(n407));
  NAND4X1 g257(.A(n405), .B(n403), .C(n402), .D(n407), .Y(n408));
  NOR2X1  g258(.A(n408), .B(n397), .Y(n409));
  NOR4X1  g259(.A(n396), .B(n378), .C(n369), .D(n409), .Y(n410));
  NAND2X1 g260(.A(RMIN_REG_5__SCAN_IN), .B(RMAX_REG_5__SCAN_IN), .Y(n411));
  AOI22X1 g261(.A0(RMIN_REG_1__SCAN_IN), .A1(RMAX_REG_1__SCAN_IN), .B0(RMAX_REG_0__SCAN_IN), .B1(RMIN_REG_0__SCAN_IN), .Y(n412));
  OAI22X1 g262(.A0(RMIN_REG_2__SCAN_IN), .A1(RMAX_REG_2__SCAN_IN), .B0(RMAX_REG_1__SCAN_IN), .B1(RMIN_REG_1__SCAN_IN), .Y(n413));
  AOI22X1 g263(.A0(RMIN_REG_3__SCAN_IN), .A1(RMAX_REG_3__SCAN_IN), .B0(RMAX_REG_2__SCAN_IN), .B1(RMIN_REG_2__SCAN_IN), .Y(n414));
  OAI21X1 g264(.A0(n413), .A1(n412), .B0(n414), .Y(n415));
  AOI22X1 g265(.A0(n206), .A1(n162), .B0(n163), .B1(n200), .Y(n416));
  AOI22X1 g266(.A0(n415), .A1(n416), .B0(RMIN_REG_4__SCAN_IN), .B1(RMAX_REG_4__SCAN_IN), .Y(n417));
  NOR2X1  g267(.A(RMIN_REG_5__SCAN_IN), .B(RMAX_REG_5__SCAN_IN), .Y(n418));
  OAI21X1 g268(.A0(n418), .A1(n417), .B0(n411), .Y(n419));
  NOR2X1  g269(.A(n419), .B(RMAX_REG_6__SCAN_IN), .Y(n420));
  AOI21X1 g270(.A0(n419), .A1(RMAX_REG_6__SCAN_IN), .B0(RMIN_REG_6__SCAN_IN), .Y(n421));
  NOR2X1  g271(.A(n421), .B(n420), .Y(n422));
  AOI21X1 g272(.A0(n193), .A1(n152), .B0(n422), .Y(n423));
  AOI21X1 g273(.A0(RMIN_REG_7__SCAN_IN), .A1(RMAX_REG_7__SCAN_IN), .B0(n423), .Y(n424));
  NOR2X1  g274(.A(n180), .B(STATO_REG_0__SCAN_IN), .Y(n425));
  NOR3X1  g275(.A(n248), .B(n424), .C(n332), .Y(n427));
  NAND2X1 g276(.A(n427), .B(n410), .Y(n428));
  NAND2X1 g277(.A(REG4_REG_5__SCAN_IN), .B(DATA_IN_5_), .Y(n429));
  AOI22X1 g278(.A0(REG4_REG_0__SCAN_IN), .A1(DATA_IN_0_), .B0(DATA_IN_1_), .B1(REG4_REG_1__SCAN_IN), .Y(n430));
  OAI22X1 g279(.A0(REG4_REG_1__SCAN_IN), .A1(DATA_IN_1_), .B0(DATA_IN_2_), .B1(REG4_REG_2__SCAN_IN), .Y(n431));
  AOI22X1 g280(.A0(REG4_REG_2__SCAN_IN), .A1(DATA_IN_2_), .B0(DATA_IN_3_), .B1(REG4_REG_3__SCAN_IN), .Y(n432));
  OAI21X1 g281(.A0(n431), .A1(n430), .B0(n432), .Y(n433));
  AOI22X1 g282(.A0(n304), .A1(n167), .B0(n159), .B1(n306), .Y(n434));
  AOI22X1 g283(.A0(n433), .A1(n434), .B0(REG4_REG_4__SCAN_IN), .B1(DATA_IN_4_), .Y(n435));
  NOR2X1  g284(.A(REG4_REG_5__SCAN_IN), .B(DATA_IN_5_), .Y(n436));
  OAI21X1 g285(.A0(n436), .A1(n435), .B0(n429), .Y(n437));
  NOR2X1  g286(.A(n437), .B(DATA_IN_6_), .Y(n438));
  AOI21X1 g287(.A0(n437), .A1(DATA_IN_6_), .B0(REG4_REG_6__SCAN_IN), .Y(n439));
  NOR2X1  g288(.A(n439), .B(n438), .Y(n440));
  AOI21X1 g289(.A0(n298), .A1(n151), .B0(n440), .Y(n441));
  AOI21X1 g290(.A0(REG4_REG_7__SCAN_IN), .A1(DATA_IN_7_), .B0(n441), .Y(n442));
  NOR2X1  g291(.A(n229), .B(AVERAGE), .Y(n443));
  NAND3X1 g292(.A(n443), .B(n425), .C(n332), .Y(n444));
  NOR2X1  g293(.A(n444), .B(n442), .Y(n445));
  NAND4X1 g294(.A(ENABLE), .B(AVERAGE), .C(n332), .D(n425), .Y(n446));
  NOR4X1  g295(.A(STATO_REG_0__SCAN_IN), .B(ENABLE), .C(RESTART), .D(n180), .Y(n447));
  AOI22X1 g296(.A0(n249), .A1(DATA_OUT_REG_7__SCAN_IN), .B0(RLAST_REG_7__SCAN_IN), .B1(n447), .Y(n448));
  OAI21X1 g297(.A0(n446), .A1(n298), .B0(n448), .Y(n449));
  AOI21X1 g298(.A0(n445), .A1(n410), .B0(n449), .Y(n450));
  NAND2X1 g299(.A(n450), .B(n428), .Y(U288));
  NOR3X1  g300(.A(n396), .B(n378), .C(n369), .Y(n452));
  OAI21X1 g301(.A0(n378), .A1(n369), .B0(n396), .Y(n453));
  NOR4X1  g302(.A(n408), .B(n397), .C(n452), .D(n453), .Y(n454));
  OAI21X1 g303(.A0(n454), .A1(n410), .B0(n427), .Y(n455));
  OAI21X1 g304(.A0(n454), .A1(n410), .B0(n445), .Y(n456));
  INVX1   g305(.A(n446), .Y(n457));
  NAND2X1 g306(.A(n457), .B(REG4_REG_6__SCAN_IN), .Y(n458));
  AOI22X1 g307(.A0(n249), .A1(DATA_OUT_REG_6__SCAN_IN), .B0(RLAST_REG_6__SCAN_IN), .B1(n447), .Y(n459));
  NAND4X1 g308(.A(n458), .B(n456), .C(n455), .D(n459), .Y(U287));
  NOR2X1  g309(.A(n378), .B(n369), .Y(n461));
  XOR2X1  g310(.A(n396), .B(n461), .Y(n462));
  XOR2X1  g311(.A(n462), .B(n409), .Y(n463));
  NAND2X1 g312(.A(n463), .B(n445), .Y(n464));
  NAND2X1 g313(.A(n463), .B(n427), .Y(n465));
  AOI21X1 g314(.A0(n443), .A1(n442), .B0(RESTART), .Y(n466));
  OAI21X1 g315(.A0(n424), .A1(n332), .B0(n425), .Y(n467));
  NOR2X1  g316(.A(n467), .B(n466), .Y(n468));
  INVX1   g317(.A(n447), .Y(n469));
  AOI22X1 g318(.A0(n249), .A1(DATA_OUT_REG_5__SCAN_IN), .B0(REG4_REG_5__SCAN_IN), .B1(n457), .Y(n470));
  OAI21X1 g319(.A0(n469), .A1(n235), .B0(n470), .Y(n471));
  AOI21X1 g320(.A0(n468), .A1(n396), .B0(n471), .Y(n472));
  NAND3X1 g321(.A(n472), .B(n465), .C(n464), .Y(U286));
  XOR2X1  g322(.A(n408), .B(n397), .Y(n474));
  NAND2X1 g323(.A(n474), .B(n445), .Y(n475));
  NAND2X1 g324(.A(n474), .B(n427), .Y(n476));
  AOI22X1 g325(.A0(n249), .A1(DATA_OUT_REG_4__SCAN_IN), .B0(REG4_REG_4__SCAN_IN), .B1(n457), .Y(n477));
  OAI21X1 g326(.A0(n469), .A1(n237), .B0(n477), .Y(n478));
  AOI21X1 g327(.A0(n468), .A1(n378), .B0(n478), .Y(n479));
  NAND3X1 g328(.A(n479), .B(n476), .C(n475), .Y(U285));
  NAND2X1 g329(.A(n468), .B(n406), .Y(n481));
  NAND2X1 g330(.A(n447), .B(RLAST_REG_3__SCAN_IN), .Y(n482));
  AOI22X1 g331(.A0(n249), .A1(DATA_OUT_REG_3__SCAN_IN), .B0(REG4_REG_3__SCAN_IN), .B1(n457), .Y(n483));
  XOR2X1  g332(.A(n357), .B(n345), .Y(n484));
  NAND2X1 g333(.A(n405), .B(n403), .Y(n485));
  NOR2X1  g334(.A(n485), .B(n484), .Y(n486));
  XOR2X1  g335(.A(n407), .B(n486), .Y(n487));
  OAI21X1 g336(.A0(n445), .A1(n427), .B0(n487), .Y(n488));
  NAND4X1 g337(.A(n483), .B(n482), .C(n481), .D(n488), .Y(U284));
  NAND2X1 g338(.A(n468), .B(n357), .Y(n490));
  XOR2X1  g339(.A(n485), .B(n484), .Y(n491));
  NAND2X1 g340(.A(n491), .B(n427), .Y(n492));
  AOI22X1 g341(.A0(n249), .A1(DATA_OUT_REG_2__SCAN_IN), .B0(REG4_REG_2__SCAN_IN), .B1(n457), .Y(n493));
  OAI21X1 g342(.A0(n469), .A1(n241), .B0(n493), .Y(n494));
  AOI21X1 g343(.A0(n491), .A1(n445), .B0(n494), .Y(n495));
  NAND3X1 g344(.A(n495), .B(n492), .C(n490), .Y(U283));
  NAND2X1 g345(.A(n468), .B(n399), .Y(n497));
  XOR2X1  g346(.A(n405), .B(n403), .Y(n498));
  NAND2X1 g347(.A(n498), .B(n427), .Y(n499));
  AOI22X1 g348(.A0(n249), .A1(DATA_OUT_REG_1__SCAN_IN), .B0(REG4_REG_1__SCAN_IN), .B1(n457), .Y(n500));
  OAI21X1 g349(.A0(n469), .A1(n243), .B0(n500), .Y(n501));
  AOI21X1 g350(.A0(n498), .A1(n445), .B0(n501), .Y(n502));
  NAND3X1 g351(.A(n502), .B(n499), .C(n497), .Y(U282));
  NAND2X1 g352(.A(n468), .B(n404), .Y(n504));
  NOR4X1  g353(.A(n424), .B(n405), .C(n332), .D(n248), .Y(n505));
  NOR3X1  g354(.A(n444), .B(n442), .C(n405), .Y(n506));
  AOI22X1 g355(.A0(n249), .A1(DATA_OUT_REG_0__SCAN_IN), .B0(REG4_REG_0__SCAN_IN), .B1(n457), .Y(n507));
  OAI21X1 g356(.A0(n469), .A1(n245), .B0(n507), .Y(n508));
  NOR3X1  g357(.A(n508), .B(n506), .C(n505), .Y(n509));
  NAND2X1 g358(.A(n509), .B(n504), .Y(U281));
endmodule


