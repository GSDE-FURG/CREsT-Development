// Benchmark "top" written by ABC on Tue Sep 21 20:59:18 2021

module top ( 
    \priority[0] , \priority[1] , \priority[2] , \priority[3] ,
    \priority[4] , \priority[5] , \priority[6] , \priority[7] ,
    \priority[8] , \priority[9] , \priority[10] , \priority[11] ,
    \priority[12] , \priority[13] , \priority[14] , \priority[15] ,
    \priority[16] , \priority[17] , \priority[18] , \priority[19] ,
    \priority[20] , \priority[21] , \priority[22] , \priority[23] ,
    \priority[24] , \priority[25] , \priority[26] , \priority[27] ,
    \priority[28] , \priority[29] , \priority[30] , \priority[31] ,
    \priority[32] , \priority[33] , \priority[34] , \priority[35] ,
    \priority[36] , \priority[37] , \priority[38] , \priority[39] ,
    \priority[40] , \priority[41] , \priority[42] , \priority[43] ,
    \priority[44] , \priority[45] , \priority[46] , \priority[47] ,
    \priority[48] , \priority[49] , \priority[50] , \priority[51] ,
    \priority[52] , \priority[53] , \priority[54] , \priority[55] ,
    \priority[56] , \priority[57] , \priority[58] , \priority[59] ,
    \priority[60] , \priority[61] , \priority[62] , \priority[63] ,
    \priority[64] , \priority[65] , \priority[66] , \priority[67] ,
    \priority[68] , \priority[69] , \priority[70] , \priority[71] ,
    \priority[72] , \priority[73] , \priority[74] , \priority[75] ,
    \priority[76] , \priority[77] , \priority[78] , \priority[79] ,
    \priority[80] , \priority[81] , \priority[82] , \priority[83] ,
    \priority[84] , \priority[85] , \priority[86] , \priority[87] ,
    \priority[88] , \priority[89] , \priority[90] , \priority[91] ,
    \priority[92] , \priority[93] , \priority[94] , \priority[95] ,
    \priority[96] , \priority[97] , \priority[98] , \priority[99] ,
    \priority[100] , \priority[101] , \priority[102] , \priority[103] ,
    \priority[104] , \priority[105] , \priority[106] , \priority[107] ,
    \priority[108] , \priority[109] , \priority[110] , \priority[111] ,
    \priority[112] , \priority[113] , \priority[114] , \priority[115] ,
    \priority[116] , \priority[117] , \priority[118] , \priority[119] ,
    \priority[120] , \priority[121] , \priority[122] , \priority[123] ,
    \priority[124] , \priority[125] , \priority[126] , \priority[127] ,
    \req[0] , \req[1] , \req[2] , \req[3] , \req[4] , \req[5] , \req[6] ,
    \req[7] , \req[8] , \req[9] , \req[10] , \req[11] , \req[12] ,
    \req[13] , \req[14] , \req[15] , \req[16] , \req[17] , \req[18] ,
    \req[19] , \req[20] , \req[21] , \req[22] , \req[23] , \req[24] ,
    \req[25] , \req[26] , \req[27] , \req[28] , \req[29] , \req[30] ,
    \req[31] , \req[32] , \req[33] , \req[34] , \req[35] , \req[36] ,
    \req[37] , \req[38] , \req[39] , \req[40] , \req[41] , \req[42] ,
    \req[43] , \req[44] , \req[45] , \req[46] , \req[47] , \req[48] ,
    \req[49] , \req[50] , \req[51] , \req[52] , \req[53] , \req[54] ,
    \req[55] , \req[56] , \req[57] , \req[58] , \req[59] , \req[60] ,
    \req[61] , \req[62] , \req[63] , \req[64] , \req[65] , \req[66] ,
    \req[67] , \req[68] , \req[69] , \req[70] , \req[71] , \req[72] ,
    \req[73] , \req[74] , \req[75] , \req[76] , \req[77] , \req[78] ,
    \req[79] , \req[80] , \req[81] , \req[82] , \req[83] , \req[84] ,
    \req[85] , \req[86] , \req[87] , \req[88] , \req[89] , \req[90] ,
    \req[91] , \req[92] , \req[93] , \req[94] , \req[95] , \req[96] ,
    \req[97] , \req[98] , \req[99] , \req[100] , \req[101] , \req[102] ,
    \req[103] , \req[104] , \req[105] , \req[106] , \req[107] , \req[108] ,
    \req[109] , \req[110] , \req[111] , \req[112] , \req[113] , \req[114] ,
    \req[115] , \req[116] , \req[117] , \req[118] , \req[119] , \req[120] ,
    \req[121] , \req[122] , \req[123] , \req[124] , \req[125] , \req[126] ,
    \req[127] ,
    \grant[0] , \grant[1] , \grant[2] , \grant[3] , \grant[4] , \grant[5] ,
    \grant[6] , \grant[7] , \grant[8] , \grant[9] , \grant[10] ,
    \grant[11] , \grant[12] , \grant[13] , \grant[14] , \grant[15] ,
    \grant[16] , \grant[17] , \grant[18] , \grant[19] , \grant[20] ,
    \grant[21] , \grant[22] , \grant[23] , \grant[24] , \grant[25] ,
    \grant[26] , \grant[27] , \grant[28] , \grant[29] , \grant[30] ,
    \grant[31] , \grant[32] , \grant[33] , \grant[34] , \grant[35] ,
    \grant[36] , \grant[37] , \grant[38] , \grant[39] , \grant[40] ,
    \grant[41] , \grant[42] , \grant[43] , \grant[44] , \grant[45] ,
    \grant[46] , \grant[47] , \grant[48] , \grant[49] , \grant[50] ,
    \grant[51] , \grant[52] , \grant[53] , \grant[54] , \grant[55] ,
    \grant[56] , \grant[57] , \grant[58] , \grant[59] , \grant[60] ,
    \grant[61] , \grant[62] , \grant[63] , \grant[64] , \grant[65] ,
    \grant[66] , \grant[67] , \grant[68] , \grant[69] , \grant[70] ,
    \grant[71] , \grant[72] , \grant[73] , \grant[74] , \grant[75] ,
    \grant[76] , \grant[77] , \grant[78] , \grant[79] , \grant[80] ,
    \grant[81] , \grant[82] , \grant[83] , \grant[84] , \grant[85] ,
    \grant[86] , \grant[87] , \grant[88] , \grant[89] , \grant[90] ,
    \grant[91] , \grant[92] , \grant[93] , \grant[94] , \grant[95] ,
    \grant[96] , \grant[97] , \grant[98] , \grant[99] , \grant[100] ,
    \grant[101] , \grant[102] , \grant[103] , \grant[104] , \grant[105] ,
    \grant[106] , \grant[107] , \grant[108] , \grant[109] , \grant[110] ,
    \grant[111] , \grant[112] , \grant[113] , \grant[114] , \grant[115] ,
    \grant[116] , \grant[117] , \grant[118] , \grant[119] , \grant[120] ,
    \grant[121] , \grant[122] , \grant[123] , \grant[124] , \grant[125] ,
    \grant[126] , \grant[127] , anyGrant  );
  input  \priority[0] , \priority[1] , \priority[2] , \priority[3] ,
    \priority[4] , \priority[5] , \priority[6] , \priority[7] ,
    \priority[8] , \priority[9] , \priority[10] , \priority[11] ,
    \priority[12] , \priority[13] , \priority[14] , \priority[15] ,
    \priority[16] , \priority[17] , \priority[18] , \priority[19] ,
    \priority[20] , \priority[21] , \priority[22] , \priority[23] ,
    \priority[24] , \priority[25] , \priority[26] , \priority[27] ,
    \priority[28] , \priority[29] , \priority[30] , \priority[31] ,
    \priority[32] , \priority[33] , \priority[34] , \priority[35] ,
    \priority[36] , \priority[37] , \priority[38] , \priority[39] ,
    \priority[40] , \priority[41] , \priority[42] , \priority[43] ,
    \priority[44] , \priority[45] , \priority[46] , \priority[47] ,
    \priority[48] , \priority[49] , \priority[50] , \priority[51] ,
    \priority[52] , \priority[53] , \priority[54] , \priority[55] ,
    \priority[56] , \priority[57] , \priority[58] , \priority[59] ,
    \priority[60] , \priority[61] , \priority[62] , \priority[63] ,
    \priority[64] , \priority[65] , \priority[66] , \priority[67] ,
    \priority[68] , \priority[69] , \priority[70] , \priority[71] ,
    \priority[72] , \priority[73] , \priority[74] , \priority[75] ,
    \priority[76] , \priority[77] , \priority[78] , \priority[79] ,
    \priority[80] , \priority[81] , \priority[82] , \priority[83] ,
    \priority[84] , \priority[85] , \priority[86] , \priority[87] ,
    \priority[88] , \priority[89] , \priority[90] , \priority[91] ,
    \priority[92] , \priority[93] , \priority[94] , \priority[95] ,
    \priority[96] , \priority[97] , \priority[98] , \priority[99] ,
    \priority[100] , \priority[101] , \priority[102] , \priority[103] ,
    \priority[104] , \priority[105] , \priority[106] , \priority[107] ,
    \priority[108] , \priority[109] , \priority[110] , \priority[111] ,
    \priority[112] , \priority[113] , \priority[114] , \priority[115] ,
    \priority[116] , \priority[117] , \priority[118] , \priority[119] ,
    \priority[120] , \priority[121] , \priority[122] , \priority[123] ,
    \priority[124] , \priority[125] , \priority[126] , \priority[127] ,
    \req[0] , \req[1] , \req[2] , \req[3] , \req[4] , \req[5] , \req[6] ,
    \req[7] , \req[8] , \req[9] , \req[10] , \req[11] , \req[12] ,
    \req[13] , \req[14] , \req[15] , \req[16] , \req[17] , \req[18] ,
    \req[19] , \req[20] , \req[21] , \req[22] , \req[23] , \req[24] ,
    \req[25] , \req[26] , \req[27] , \req[28] , \req[29] , \req[30] ,
    \req[31] , \req[32] , \req[33] , \req[34] , \req[35] , \req[36] ,
    \req[37] , \req[38] , \req[39] , \req[40] , \req[41] , \req[42] ,
    \req[43] , \req[44] , \req[45] , \req[46] , \req[47] , \req[48] ,
    \req[49] , \req[50] , \req[51] , \req[52] , \req[53] , \req[54] ,
    \req[55] , \req[56] , \req[57] , \req[58] , \req[59] , \req[60] ,
    \req[61] , \req[62] , \req[63] , \req[64] , \req[65] , \req[66] ,
    \req[67] , \req[68] , \req[69] , \req[70] , \req[71] , \req[72] ,
    \req[73] , \req[74] , \req[75] , \req[76] , \req[77] , \req[78] ,
    \req[79] , \req[80] , \req[81] , \req[82] , \req[83] , \req[84] ,
    \req[85] , \req[86] , \req[87] , \req[88] , \req[89] , \req[90] ,
    \req[91] , \req[92] , \req[93] , \req[94] , \req[95] , \req[96] ,
    \req[97] , \req[98] , \req[99] , \req[100] , \req[101] , \req[102] ,
    \req[103] , \req[104] , \req[105] , \req[106] , \req[107] , \req[108] ,
    \req[109] , \req[110] , \req[111] , \req[112] , \req[113] , \req[114] ,
    \req[115] , \req[116] , \req[117] , \req[118] , \req[119] , \req[120] ,
    \req[121] , \req[122] , \req[123] , \req[124] , \req[125] , \req[126] ,
    \req[127] ;
  output \grant[0] , \grant[1] , \grant[2] , \grant[3] , \grant[4] ,
    \grant[5] , \grant[6] , \grant[7] , \grant[8] , \grant[9] ,
    \grant[10] , \grant[11] , \grant[12] , \grant[13] , \grant[14] ,
    \grant[15] , \grant[16] , \grant[17] , \grant[18] , \grant[19] ,
    \grant[20] , \grant[21] , \grant[22] , \grant[23] , \grant[24] ,
    \grant[25] , \grant[26] , \grant[27] , \grant[28] , \grant[29] ,
    \grant[30] , \grant[31] , \grant[32] , \grant[33] , \grant[34] ,
    \grant[35] , \grant[36] , \grant[37] , \grant[38] , \grant[39] ,
    \grant[40] , \grant[41] , \grant[42] , \grant[43] , \grant[44] ,
    \grant[45] , \grant[46] , \grant[47] , \grant[48] , \grant[49] ,
    \grant[50] , \grant[51] , \grant[52] , \grant[53] , \grant[54] ,
    \grant[55] , \grant[56] , \grant[57] , \grant[58] , \grant[59] ,
    \grant[60] , \grant[61] , \grant[62] , \grant[63] , \grant[64] ,
    \grant[65] , \grant[66] , \grant[67] , \grant[68] , \grant[69] ,
    \grant[70] , \grant[71] , \grant[72] , \grant[73] , \grant[74] ,
    \grant[75] , \grant[76] , \grant[77] , \grant[78] , \grant[79] ,
    \grant[80] , \grant[81] , \grant[82] , \grant[83] , \grant[84] ,
    \grant[85] , \grant[86] , \grant[87] , \grant[88] , \grant[89] ,
    \grant[90] , \grant[91] , \grant[92] , \grant[93] , \grant[94] ,
    \grant[95] , \grant[96] , \grant[97] , \grant[98] , \grant[99] ,
    \grant[100] , \grant[101] , \grant[102] , \grant[103] , \grant[104] ,
    \grant[105] , \grant[106] , \grant[107] , \grant[108] , \grant[109] ,
    \grant[110] , \grant[111] , \grant[112] , \grant[113] , \grant[114] ,
    \grant[115] , \grant[116] , \grant[117] , \grant[118] , \grant[119] ,
    \grant[120] , \grant[121] , \grant[122] , \grant[123] , \grant[124] ,
    \grant[125] , \grant[126] , \grant[127] , anyGrant;
  wire new_n386_, new_n387_, new_n388_, new_n389_, new_n390_, new_n391_,
    new_n392_, new_n393_, new_n394_, new_n395_, new_n396_, new_n397_,
    new_n398_, new_n399_, new_n400_, new_n401_, new_n402_, new_n403_,
    new_n404_, new_n405_, new_n406_, new_n407_, new_n408_, new_n409_,
    new_n410_, new_n411_, new_n412_, new_n413_, new_n414_, new_n415_,
    new_n416_, new_n417_, new_n418_, new_n419_, new_n420_, new_n421_,
    new_n422_, new_n423_, new_n424_, new_n425_, new_n426_, new_n427_,
    new_n428_, new_n429_, new_n430_, new_n431_, new_n432_, new_n433_,
    new_n434_, new_n435_, new_n436_, new_n437_, new_n438_, new_n439_,
    new_n440_, new_n441_, new_n442_, new_n443_, new_n444_, new_n445_,
    new_n446_, new_n447_, new_n448_, new_n449_, new_n450_, new_n451_,
    new_n452_, new_n453_, new_n454_, new_n455_, new_n456_, new_n457_,
    new_n458_, new_n459_, new_n460_, new_n461_, new_n462_, new_n463_,
    new_n464_, new_n465_, new_n466_, new_n467_, new_n468_, new_n469_,
    new_n470_, new_n471_, new_n472_, new_n473_, new_n474_, new_n475_,
    new_n476_, new_n477_, new_n478_, new_n479_, new_n480_, new_n481_,
    new_n482_, new_n483_, new_n484_, new_n485_, new_n486_, new_n487_,
    new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n493_,
    new_n494_, new_n495_, new_n496_, new_n497_, new_n498_, new_n499_,
    new_n500_, new_n501_, new_n502_, new_n503_, new_n504_, new_n505_,
    new_n506_, new_n507_, new_n508_, new_n509_, new_n510_, new_n511_,
    new_n512_, new_n513_, new_n514_, new_n515_, new_n516_, new_n517_,
    new_n518_, new_n519_, new_n520_, new_n521_, new_n522_, new_n523_,
    new_n524_, new_n525_, new_n526_, new_n527_, new_n528_, new_n529_,
    new_n530_, new_n531_, new_n532_, new_n533_, new_n534_, new_n535_,
    new_n536_, new_n537_, new_n538_, new_n539_, new_n540_, new_n541_,
    new_n542_, new_n543_, new_n544_, new_n545_, new_n546_, new_n547_,
    new_n548_, new_n549_, new_n550_, new_n551_, new_n552_, new_n553_,
    new_n554_, new_n555_, new_n556_, new_n557_, new_n558_, new_n559_,
    new_n560_, new_n561_, new_n562_, new_n563_, new_n564_, new_n565_,
    new_n566_, new_n567_, new_n568_, new_n569_, new_n570_, new_n571_,
    new_n572_, new_n573_, new_n574_, new_n575_, new_n576_, new_n577_,
    new_n578_, new_n579_, new_n580_, new_n581_, new_n582_, new_n583_,
    new_n584_, new_n585_, new_n586_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n636_, new_n637_,
    new_n638_, new_n639_, new_n640_, new_n641_, new_n642_, new_n643_,
    new_n644_, new_n645_, new_n646_, new_n647_, new_n648_, new_n649_,
    new_n650_, new_n651_, new_n652_, new_n653_, new_n654_, new_n655_,
    new_n656_, new_n657_, new_n658_, new_n659_, new_n660_, new_n661_,
    new_n662_, new_n663_, new_n664_, new_n665_, new_n666_, new_n667_,
    new_n668_, new_n669_, new_n670_, new_n671_, new_n672_, new_n673_,
    new_n674_, new_n675_, new_n676_, new_n677_, new_n678_, new_n679_,
    new_n680_, new_n681_, new_n682_, new_n683_, new_n684_, new_n685_,
    new_n686_, new_n687_, new_n688_, new_n689_, new_n690_, new_n691_,
    new_n692_, new_n693_, new_n694_, new_n695_, new_n696_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n706_, new_n707_, new_n708_, new_n709_,
    new_n710_, new_n711_, new_n712_, new_n713_, new_n714_, new_n715_,
    new_n716_, new_n717_, new_n718_, new_n719_, new_n720_, new_n721_,
    new_n722_, new_n723_, new_n724_, new_n725_, new_n726_, new_n727_,
    new_n728_, new_n729_, new_n730_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n944_,
    new_n945_, new_n946_, new_n947_, new_n948_, new_n949_, new_n950_,
    new_n951_, new_n952_, new_n953_, new_n954_, new_n955_, new_n956_,
    new_n957_, new_n958_, new_n959_, new_n960_, new_n961_, new_n962_,
    new_n963_, new_n964_, new_n965_, new_n966_, new_n967_, new_n968_,
    new_n969_, new_n970_, new_n971_, new_n972_, new_n973_, new_n974_,
    new_n975_, new_n976_, new_n977_, new_n978_, new_n979_, new_n980_,
    new_n981_, new_n982_, new_n983_, new_n984_, new_n985_, new_n986_,
    new_n987_, new_n988_, new_n989_, new_n990_, new_n991_, new_n992_,
    new_n993_, new_n994_, new_n995_, new_n996_, new_n997_, new_n998_,
    new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_,
    new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_,
    new_n1011_, new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_,
    new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_,
    new_n1023_, new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_,
    new_n1029_, new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_,
    new_n1035_, new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_,
    new_n1041_, new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_,
    new_n1047_, new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_,
    new_n1053_, new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_,
    new_n1059_, new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_,
    new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_,
    new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_,
    new_n1077_, new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_,
    new_n1083_, new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_,
    new_n1089_, new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_,
    new_n1095_, new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_,
    new_n1101_, new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_,
    new_n1107_, new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_,
    new_n1113_, new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_,
    new_n1119_, new_n1120_, new_n1121_, new_n1122_, new_n1123_, new_n1124_,
    new_n1125_, new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_,
    new_n1131_, new_n1132_, new_n1133_, new_n1134_, new_n1135_, new_n1136_,
    new_n1137_, new_n1138_, new_n1139_, new_n1140_, new_n1141_, new_n1142_,
    new_n1143_, new_n1144_, new_n1145_, new_n1146_, new_n1147_, new_n1148_,
    new_n1149_, new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1154_,
    new_n1155_, new_n1156_, new_n1157_, new_n1158_, new_n1159_, new_n1160_,
    new_n1161_, new_n1162_, new_n1163_, new_n1164_, new_n1165_, new_n1166_,
    new_n1167_, new_n1168_, new_n1169_, new_n1170_, new_n1171_, new_n1172_,
    new_n1173_, new_n1174_, new_n1175_, new_n1176_, new_n1177_, new_n1178_,
    new_n1179_, new_n1180_, new_n1181_, new_n1182_, new_n1183_, new_n1184_,
    new_n1185_, new_n1186_, new_n1187_, new_n1188_, new_n1189_, new_n1190_,
    new_n1191_, new_n1192_, new_n1194_, new_n1195_, new_n1196_, new_n1197_,
    new_n1198_, new_n1199_, new_n1200_, new_n1201_, new_n1202_, new_n1203_,
    new_n1204_, new_n1205_, new_n1206_, new_n1207_, new_n1208_, new_n1209_,
    new_n1210_, new_n1211_, new_n1212_, new_n1213_, new_n1214_, new_n1215_,
    new_n1216_, new_n1217_, new_n1218_, new_n1219_, new_n1220_, new_n1221_,
    new_n1222_, new_n1223_, new_n1224_, new_n1225_, new_n1226_, new_n1227_,
    new_n1228_, new_n1229_, new_n1230_, new_n1231_, new_n1232_, new_n1233_,
    new_n1234_, new_n1235_, new_n1236_, new_n1237_, new_n1238_, new_n1239_,
    new_n1240_, new_n1241_, new_n1242_, new_n1243_, new_n1244_, new_n1245_,
    new_n1246_, new_n1247_, new_n1248_, new_n1249_, new_n1250_, new_n1251_,
    new_n1252_, new_n1253_, new_n1254_, new_n1255_, new_n1256_, new_n1257_,
    new_n1258_, new_n1259_, new_n1260_, new_n1261_, new_n1262_, new_n1263_,
    new_n1264_, new_n1265_, new_n1266_, new_n1267_, new_n1268_, new_n1269_,
    new_n1270_, new_n1271_, new_n1272_, new_n1273_, new_n1274_, new_n1275_,
    new_n1276_, new_n1277_, new_n1278_, new_n1279_, new_n1280_, new_n1281_,
    new_n1282_, new_n1283_, new_n1284_, new_n1285_, new_n1286_, new_n1287_,
    new_n1288_, new_n1289_, new_n1290_, new_n1291_, new_n1292_, new_n1293_,
    new_n1294_, new_n1295_, new_n1296_, new_n1297_, new_n1298_, new_n1299_,
    new_n1300_, new_n1301_, new_n1302_, new_n1303_, new_n1304_, new_n1305_,
    new_n1306_, new_n1307_, new_n1308_, new_n1309_, new_n1310_, new_n1311_,
    new_n1312_, new_n1313_, new_n1314_, new_n1315_, new_n1316_, new_n1317_,
    new_n1318_, new_n1319_, new_n1320_, new_n1321_, new_n1322_, new_n1323_,
    new_n1324_, new_n1325_, new_n1326_, new_n1327_, new_n1328_, new_n1329_,
    new_n1330_, new_n1331_, new_n1332_, new_n1333_, new_n1334_, new_n1335_,
    new_n1336_, new_n1337_, new_n1338_, new_n1339_, new_n1340_, new_n1341_,
    new_n1342_, new_n1343_, new_n1344_, new_n1345_, new_n1346_, new_n1347_,
    new_n1348_, new_n1349_, new_n1350_, new_n1351_, new_n1352_, new_n1353_,
    new_n1354_, new_n1355_, new_n1356_, new_n1357_, new_n1358_, new_n1359_,
    new_n1360_, new_n1361_, new_n1362_, new_n1363_, new_n1364_, new_n1365_,
    new_n1366_, new_n1367_, new_n1368_, new_n1369_, new_n1370_, new_n1371_,
    new_n1372_, new_n1373_, new_n1374_, new_n1375_, new_n1376_, new_n1377_,
    new_n1378_, new_n1379_, new_n1380_, new_n1381_, new_n1382_, new_n1383_,
    new_n1384_, new_n1385_, new_n1386_, new_n1387_, new_n1388_, new_n1389_,
    new_n1390_, new_n1391_, new_n1392_, new_n1393_, new_n1394_, new_n1395_,
    new_n1396_, new_n1397_, new_n1398_, new_n1399_, new_n1400_, new_n1401_,
    new_n1402_, new_n1403_, new_n1404_, new_n1405_, new_n1406_, new_n1407_,
    new_n1408_, new_n1409_, new_n1410_, new_n1411_, new_n1412_, new_n1413_,
    new_n1414_, new_n1415_, new_n1416_, new_n1417_, new_n1418_, new_n1419_,
    new_n1420_, new_n1421_, new_n1422_, new_n1423_, new_n1424_, new_n1425_,
    new_n1426_, new_n1427_, new_n1428_, new_n1429_, new_n1430_, new_n1431_,
    new_n1432_, new_n1433_, new_n1434_, new_n1435_, new_n1436_, new_n1437_,
    new_n1438_, new_n1439_, new_n1440_, new_n1441_, new_n1442_, new_n1443_,
    new_n1444_, new_n1445_, new_n1446_, new_n1447_, new_n1448_, new_n1449_,
    new_n1450_, new_n1451_, new_n1452_, new_n1453_, new_n1454_, new_n1455_,
    new_n1456_, new_n1457_, new_n1458_, new_n1459_, new_n1460_, new_n1461_,
    new_n1462_, new_n1463_, new_n1464_, new_n1465_, new_n1466_, new_n1467_,
    new_n1468_, new_n1469_, new_n1470_, new_n1471_, new_n1472_, new_n1473_,
    new_n1474_, new_n1475_, new_n1476_, new_n1477_, new_n1478_, new_n1479_,
    new_n1480_, new_n1481_, new_n1482_, new_n1483_, new_n1484_, new_n1485_,
    new_n1486_, new_n1487_, new_n1488_, new_n1489_, new_n1490_, new_n1491_,
    new_n1492_, new_n1493_, new_n1494_, new_n1495_, new_n1496_, new_n1497_,
    new_n1498_, new_n1499_, new_n1500_, new_n1501_, new_n1502_, new_n1503_,
    new_n1504_, new_n1505_, new_n1506_, new_n1507_, new_n1508_, new_n1509_,
    new_n1510_, new_n1511_, new_n1512_, new_n1513_, new_n1514_, new_n1515_,
    new_n1516_, new_n1517_, new_n1518_, new_n1519_, new_n1520_, new_n1521_,
    new_n1522_, new_n1523_, new_n1524_, new_n1525_, new_n1526_, new_n1527_,
    new_n1528_, new_n1529_, new_n1530_, new_n1532_, new_n1533_, new_n1534_,
    new_n1535_, new_n1536_, new_n1537_, new_n1538_, new_n1539_, new_n1540_,
    new_n1541_, new_n1542_, new_n1543_, new_n1544_, new_n1545_, new_n1546_,
    new_n1547_, new_n1548_, new_n1549_, new_n1550_, new_n1551_, new_n1552_,
    new_n1553_, new_n1554_, new_n1555_, new_n1556_, new_n1557_, new_n1558_,
    new_n1559_, new_n1560_, new_n1561_, new_n1562_, new_n1563_, new_n1564_,
    new_n1565_, new_n1566_, new_n1567_, new_n1568_, new_n1569_, new_n1570_,
    new_n1571_, new_n1572_, new_n1573_, new_n1574_, new_n1575_, new_n1576_,
    new_n1577_, new_n1578_, new_n1579_, new_n1580_, new_n1581_, new_n1582_,
    new_n1583_, new_n1584_, new_n1585_, new_n1586_, new_n1587_, new_n1588_,
    new_n1589_, new_n1590_, new_n1591_, new_n1592_, new_n1593_, new_n1594_,
    new_n1595_, new_n1596_, new_n1597_, new_n1598_, new_n1599_, new_n1600_,
    new_n1601_, new_n1602_, new_n1603_, new_n1604_, new_n1605_, new_n1606_,
    new_n1607_, new_n1608_, new_n1609_, new_n1610_, new_n1611_, new_n1612_,
    new_n1613_, new_n1614_, new_n1615_, new_n1616_, new_n1617_, new_n1618_,
    new_n1619_, new_n1620_, new_n1621_, new_n1623_, new_n1624_, new_n1625_,
    new_n1626_, new_n1627_, new_n1628_, new_n1629_, new_n1630_, new_n1631_,
    new_n1632_, new_n1633_, new_n1634_, new_n1635_, new_n1636_, new_n1637_,
    new_n1638_, new_n1639_, new_n1640_, new_n1641_, new_n1642_, new_n1643_,
    new_n1644_, new_n1645_, new_n1646_, new_n1647_, new_n1648_, new_n1649_,
    new_n1650_, new_n1651_, new_n1652_, new_n1653_, new_n1654_, new_n1655_,
    new_n1656_, new_n1657_, new_n1658_, new_n1659_, new_n1660_, new_n1661_,
    new_n1662_, new_n1663_, new_n1664_, new_n1665_, new_n1666_, new_n1667_,
    new_n1668_, new_n1669_, new_n1670_, new_n1671_, new_n1672_, new_n1673_,
    new_n1674_, new_n1675_, new_n1676_, new_n1677_, new_n1678_, new_n1679_,
    new_n1680_, new_n1681_, new_n1682_, new_n1683_, new_n1684_, new_n1685_,
    new_n1686_, new_n1687_, new_n1688_, new_n1689_, new_n1690_, new_n1691_,
    new_n1692_, new_n1693_, new_n1694_, new_n1695_, new_n1696_, new_n1697_,
    new_n1698_, new_n1699_, new_n1700_, new_n1701_, new_n1702_, new_n1703_,
    new_n1704_, new_n1705_, new_n1706_, new_n1707_, new_n1708_, new_n1709_,
    new_n1710_, new_n1711_, new_n1712_, new_n1714_, new_n1715_, new_n1716_,
    new_n1717_, new_n1718_, new_n1719_, new_n1720_, new_n1721_, new_n1722_,
    new_n1723_, new_n1724_, new_n1725_, new_n1726_, new_n1727_, new_n1728_,
    new_n1729_, new_n1730_, new_n1731_, new_n1732_, new_n1733_, new_n1734_,
    new_n1735_, new_n1736_, new_n1737_, new_n1738_, new_n1739_, new_n1740_,
    new_n1741_, new_n1742_, new_n1743_, new_n1744_, new_n1745_, new_n1746_,
    new_n1747_, new_n1748_, new_n1749_, new_n1750_, new_n1751_, new_n1752_,
    new_n1753_, new_n1754_, new_n1755_, new_n1756_, new_n1757_, new_n1758_,
    new_n1759_, new_n1760_, new_n1761_, new_n1762_, new_n1763_, new_n1764_,
    new_n1765_, new_n1766_, new_n1767_, new_n1768_, new_n1769_, new_n1770_,
    new_n1771_, new_n1772_, new_n1773_, new_n1774_, new_n1775_, new_n1776_,
    new_n1777_, new_n1778_, new_n1779_, new_n1780_, new_n1781_, new_n1782_,
    new_n1783_, new_n1784_, new_n1785_, new_n1786_, new_n1787_, new_n1788_,
    new_n1789_, new_n1790_, new_n1791_, new_n1792_, new_n1793_, new_n1794_,
    new_n1795_, new_n1796_, new_n1797_, new_n1798_, new_n1799_, new_n1800_,
    new_n1802_, new_n1803_, new_n1804_, new_n1805_, new_n1806_, new_n1807_,
    new_n1808_, new_n1809_, new_n1810_, new_n1811_, new_n1812_, new_n1813_,
    new_n1814_, new_n1815_, new_n1816_, new_n1817_, new_n1818_, new_n1819_,
    new_n1820_, new_n1821_, new_n1822_, new_n1823_, new_n1824_, new_n1825_,
    new_n1826_, new_n1827_, new_n1828_, new_n1829_, new_n1830_, new_n1831_,
    new_n1832_, new_n1833_, new_n1834_, new_n1835_, new_n1836_, new_n1837_,
    new_n1838_, new_n1839_, new_n1840_, new_n1841_, new_n1842_, new_n1843_,
    new_n1844_, new_n1845_, new_n1846_, new_n1847_, new_n1848_, new_n1849_,
    new_n1850_, new_n1851_, new_n1852_, new_n1853_, new_n1854_, new_n1855_,
    new_n1856_, new_n1857_, new_n1858_, new_n1859_, new_n1860_, new_n1861_,
    new_n1862_, new_n1863_, new_n1864_, new_n1865_, new_n1866_, new_n1867_,
    new_n1868_, new_n1869_, new_n1870_, new_n1871_, new_n1872_, new_n1873_,
    new_n1874_, new_n1875_, new_n1876_, new_n1877_, new_n1878_, new_n1879_,
    new_n1880_, new_n1881_, new_n1882_, new_n1883_, new_n1884_, new_n1885_,
    new_n1886_, new_n1887_, new_n1888_, new_n1890_, new_n1891_, new_n1892_,
    new_n1893_, new_n1894_, new_n1895_, new_n1896_, new_n1897_, new_n1898_,
    new_n1899_, new_n1900_, new_n1901_, new_n1902_, new_n1903_, new_n1904_,
    new_n1905_, new_n1906_, new_n1907_, new_n1908_, new_n1909_, new_n1910_,
    new_n1911_, new_n1912_, new_n1913_, new_n1914_, new_n1915_, new_n1916_,
    new_n1917_, new_n1918_, new_n1919_, new_n1920_, new_n1921_, new_n1922_,
    new_n1923_, new_n1924_, new_n1925_, new_n1926_, new_n1927_, new_n1928_,
    new_n1929_, new_n1930_, new_n1931_, new_n1932_, new_n1933_, new_n1934_,
    new_n1935_, new_n1936_, new_n1937_, new_n1938_, new_n1939_, new_n1940_,
    new_n1941_, new_n1942_, new_n1943_, new_n1944_, new_n1945_, new_n1946_,
    new_n1947_, new_n1948_, new_n1949_, new_n1950_, new_n1951_, new_n1952_,
    new_n1953_, new_n1954_, new_n1955_, new_n1956_, new_n1957_, new_n1958_,
    new_n1959_, new_n1960_, new_n1961_, new_n1962_, new_n1963_, new_n1964_,
    new_n1965_, new_n1966_, new_n1967_, new_n1968_, new_n1969_, new_n1970_,
    new_n1971_, new_n1972_, new_n1973_, new_n1974_, new_n1975_, new_n1976_,
    new_n1978_, new_n1979_, new_n1980_, new_n1981_, new_n1982_, new_n1983_,
    new_n1984_, new_n1985_, new_n1986_, new_n1987_, new_n1988_, new_n1989_,
    new_n1990_, new_n1991_, new_n1992_, new_n1993_, new_n1994_, new_n1995_,
    new_n1996_, new_n1997_, new_n1998_, new_n1999_, new_n2000_, new_n2001_,
    new_n2002_, new_n2003_, new_n2004_, new_n2005_, new_n2006_, new_n2007_,
    new_n2008_, new_n2009_, new_n2010_, new_n2011_, new_n2012_, new_n2013_,
    new_n2014_, new_n2015_, new_n2016_, new_n2017_, new_n2018_, new_n2019_,
    new_n2020_, new_n2021_, new_n2022_, new_n2023_, new_n2024_, new_n2025_,
    new_n2026_, new_n2027_, new_n2028_, new_n2029_, new_n2030_, new_n2031_,
    new_n2032_, new_n2033_, new_n2034_, new_n2035_, new_n2036_, new_n2037_,
    new_n2038_, new_n2039_, new_n2040_, new_n2041_, new_n2042_, new_n2043_,
    new_n2044_, new_n2045_, new_n2046_, new_n2047_, new_n2048_, new_n2049_,
    new_n2050_, new_n2051_, new_n2052_, new_n2053_, new_n2054_, new_n2055_,
    new_n2056_, new_n2057_, new_n2058_, new_n2059_, new_n2060_, new_n2061_,
    new_n2062_, new_n2063_, new_n2065_, new_n2066_, new_n2067_, new_n2068_,
    new_n2069_, new_n2070_, new_n2071_, new_n2072_, new_n2073_, new_n2074_,
    new_n2075_, new_n2076_, new_n2077_, new_n2078_, new_n2079_, new_n2080_,
    new_n2081_, new_n2082_, new_n2083_, new_n2084_, new_n2085_, new_n2086_,
    new_n2087_, new_n2088_, new_n2089_, new_n2090_, new_n2091_, new_n2092_,
    new_n2093_, new_n2094_, new_n2095_, new_n2096_, new_n2097_, new_n2098_,
    new_n2099_, new_n2100_, new_n2101_, new_n2102_, new_n2103_, new_n2104_,
    new_n2105_, new_n2106_, new_n2107_, new_n2108_, new_n2109_, new_n2110_,
    new_n2111_, new_n2112_, new_n2113_, new_n2114_, new_n2115_, new_n2116_,
    new_n2117_, new_n2118_, new_n2119_, new_n2120_, new_n2121_, new_n2122_,
    new_n2123_, new_n2124_, new_n2125_, new_n2126_, new_n2127_, new_n2128_,
    new_n2129_, new_n2130_, new_n2131_, new_n2132_, new_n2133_, new_n2134_,
    new_n2135_, new_n2136_, new_n2137_, new_n2138_, new_n2139_, new_n2140_,
    new_n2141_, new_n2142_, new_n2143_, new_n2144_, new_n2145_, new_n2146_,
    new_n2147_, new_n2148_, new_n2149_, new_n2150_, new_n2152_, new_n2153_,
    new_n2154_, new_n2155_, new_n2156_, new_n2157_, new_n2158_, new_n2159_,
    new_n2160_, new_n2161_, new_n2162_, new_n2163_, new_n2164_, new_n2165_,
    new_n2166_, new_n2167_, new_n2168_, new_n2169_, new_n2170_, new_n2171_,
    new_n2172_, new_n2173_, new_n2174_, new_n2175_, new_n2176_, new_n2177_,
    new_n2178_, new_n2179_, new_n2180_, new_n2181_, new_n2182_, new_n2183_,
    new_n2184_, new_n2185_, new_n2186_, new_n2187_, new_n2188_, new_n2189_,
    new_n2190_, new_n2191_, new_n2192_, new_n2193_, new_n2194_, new_n2195_,
    new_n2196_, new_n2197_, new_n2198_, new_n2199_, new_n2200_, new_n2201_,
    new_n2202_, new_n2203_, new_n2204_, new_n2205_, new_n2206_, new_n2207_,
    new_n2208_, new_n2209_, new_n2210_, new_n2211_, new_n2212_, new_n2213_,
    new_n2214_, new_n2215_, new_n2216_, new_n2217_, new_n2218_, new_n2219_,
    new_n2220_, new_n2221_, new_n2222_, new_n2223_, new_n2224_, new_n2225_,
    new_n2226_, new_n2227_, new_n2228_, new_n2229_, new_n2230_, new_n2231_,
    new_n2232_, new_n2233_, new_n2234_, new_n2235_, new_n2236_, new_n2237_,
    new_n2239_, new_n2240_, new_n2241_, new_n2242_, new_n2243_, new_n2244_,
    new_n2245_, new_n2246_, new_n2247_, new_n2248_, new_n2249_, new_n2250_,
    new_n2251_, new_n2252_, new_n2253_, new_n2254_, new_n2255_, new_n2256_,
    new_n2257_, new_n2258_, new_n2259_, new_n2260_, new_n2261_, new_n2262_,
    new_n2263_, new_n2264_, new_n2265_, new_n2266_, new_n2267_, new_n2268_,
    new_n2269_, new_n2270_, new_n2271_, new_n2272_, new_n2273_, new_n2274_,
    new_n2275_, new_n2276_, new_n2277_, new_n2278_, new_n2279_, new_n2280_,
    new_n2281_, new_n2282_, new_n2283_, new_n2284_, new_n2285_, new_n2286_,
    new_n2287_, new_n2288_, new_n2289_, new_n2290_, new_n2291_, new_n2292_,
    new_n2293_, new_n2294_, new_n2295_, new_n2296_, new_n2297_, new_n2298_,
    new_n2299_, new_n2300_, new_n2301_, new_n2302_, new_n2303_, new_n2304_,
    new_n2305_, new_n2306_, new_n2307_, new_n2308_, new_n2309_, new_n2310_,
    new_n2311_, new_n2312_, new_n2313_, new_n2314_, new_n2315_, new_n2316_,
    new_n2317_, new_n2318_, new_n2319_, new_n2320_, new_n2321_, new_n2322_,
    new_n2323_, new_n2324_, new_n2326_, new_n2327_, new_n2328_, new_n2329_,
    new_n2330_, new_n2331_, new_n2332_, new_n2333_, new_n2334_, new_n2335_,
    new_n2336_, new_n2337_, new_n2338_, new_n2339_, new_n2340_, new_n2341_,
    new_n2342_, new_n2343_, new_n2344_, new_n2345_, new_n2346_, new_n2347_,
    new_n2348_, new_n2349_, new_n2350_, new_n2351_, new_n2352_, new_n2353_,
    new_n2354_, new_n2355_, new_n2356_, new_n2357_, new_n2358_, new_n2359_,
    new_n2360_, new_n2361_, new_n2362_, new_n2363_, new_n2364_, new_n2365_,
    new_n2366_, new_n2367_, new_n2368_, new_n2369_, new_n2370_, new_n2371_,
    new_n2372_, new_n2373_, new_n2374_, new_n2375_, new_n2376_, new_n2377_,
    new_n2378_, new_n2379_, new_n2380_, new_n2381_, new_n2382_, new_n2383_,
    new_n2384_, new_n2385_, new_n2386_, new_n2387_, new_n2388_, new_n2389_,
    new_n2390_, new_n2391_, new_n2392_, new_n2393_, new_n2394_, new_n2395_,
    new_n2396_, new_n2397_, new_n2398_, new_n2399_, new_n2400_, new_n2401_,
    new_n2402_, new_n2403_, new_n2404_, new_n2405_, new_n2406_, new_n2407_,
    new_n2408_, new_n2409_, new_n2410_, new_n2411_, new_n2413_, new_n2414_,
    new_n2415_, new_n2416_, new_n2417_, new_n2418_, new_n2419_, new_n2420_,
    new_n2421_, new_n2422_, new_n2423_, new_n2424_, new_n2425_, new_n2426_,
    new_n2427_, new_n2428_, new_n2429_, new_n2430_, new_n2431_, new_n2432_,
    new_n2433_, new_n2434_, new_n2435_, new_n2436_, new_n2437_, new_n2438_,
    new_n2439_, new_n2440_, new_n2441_, new_n2442_, new_n2443_, new_n2444_,
    new_n2445_, new_n2446_, new_n2447_, new_n2448_, new_n2449_, new_n2450_,
    new_n2451_, new_n2452_, new_n2453_, new_n2454_, new_n2455_, new_n2456_,
    new_n2457_, new_n2458_, new_n2459_, new_n2460_, new_n2461_, new_n2462_,
    new_n2463_, new_n2464_, new_n2465_, new_n2466_, new_n2467_, new_n2468_,
    new_n2469_, new_n2470_, new_n2471_, new_n2472_, new_n2473_, new_n2474_,
    new_n2475_, new_n2476_, new_n2477_, new_n2478_, new_n2479_, new_n2480_,
    new_n2481_, new_n2482_, new_n2483_, new_n2484_, new_n2485_, new_n2486_,
    new_n2487_, new_n2488_, new_n2489_, new_n2490_, new_n2491_, new_n2492_,
    new_n2493_, new_n2494_, new_n2495_, new_n2496_, new_n2497_, new_n2498_,
    new_n2500_, new_n2501_, new_n2502_, new_n2503_, new_n2504_, new_n2505_,
    new_n2506_, new_n2507_, new_n2508_, new_n2509_, new_n2510_, new_n2511_,
    new_n2512_, new_n2513_, new_n2514_, new_n2515_, new_n2516_, new_n2517_,
    new_n2518_, new_n2519_, new_n2520_, new_n2521_, new_n2522_, new_n2523_,
    new_n2524_, new_n2525_, new_n2526_, new_n2527_, new_n2528_, new_n2529_,
    new_n2530_, new_n2531_, new_n2532_, new_n2533_, new_n2534_, new_n2535_,
    new_n2536_, new_n2537_, new_n2538_, new_n2539_, new_n2540_, new_n2541_,
    new_n2542_, new_n2543_, new_n2544_, new_n2545_, new_n2546_, new_n2547_,
    new_n2548_, new_n2549_, new_n2550_, new_n2551_, new_n2552_, new_n2553_,
    new_n2554_, new_n2555_, new_n2556_, new_n2557_, new_n2558_, new_n2559_,
    new_n2560_, new_n2561_, new_n2562_, new_n2563_, new_n2564_, new_n2565_,
    new_n2566_, new_n2567_, new_n2568_, new_n2569_, new_n2570_, new_n2571_,
    new_n2572_, new_n2573_, new_n2574_, new_n2575_, new_n2576_, new_n2577_,
    new_n2578_, new_n2579_, new_n2580_, new_n2581_, new_n2582_, new_n2583_,
    new_n2584_, new_n2585_, new_n2587_, new_n2588_, new_n2589_, new_n2590_,
    new_n2591_, new_n2592_, new_n2593_, new_n2594_, new_n2595_, new_n2596_,
    new_n2597_, new_n2598_, new_n2599_, new_n2600_, new_n2601_, new_n2602_,
    new_n2603_, new_n2604_, new_n2605_, new_n2606_, new_n2607_, new_n2608_,
    new_n2609_, new_n2610_, new_n2611_, new_n2612_, new_n2613_, new_n2614_,
    new_n2615_, new_n2616_, new_n2617_, new_n2618_, new_n2619_, new_n2620_,
    new_n2621_, new_n2622_, new_n2623_, new_n2624_, new_n2625_, new_n2626_,
    new_n2627_, new_n2628_, new_n2629_, new_n2630_, new_n2631_, new_n2632_,
    new_n2633_, new_n2634_, new_n2635_, new_n2636_, new_n2637_, new_n2638_,
    new_n2639_, new_n2640_, new_n2641_, new_n2642_, new_n2643_, new_n2644_,
    new_n2645_, new_n2646_, new_n2647_, new_n2648_, new_n2649_, new_n2650_,
    new_n2651_, new_n2652_, new_n2653_, new_n2654_, new_n2655_, new_n2656_,
    new_n2657_, new_n2658_, new_n2659_, new_n2660_, new_n2661_, new_n2662_,
    new_n2663_, new_n2664_, new_n2665_, new_n2666_, new_n2667_, new_n2668_,
    new_n2669_, new_n2670_, new_n2671_, new_n2672_, new_n2674_, new_n2675_,
    new_n2676_, new_n2677_, new_n2678_, new_n2679_, new_n2680_, new_n2681_,
    new_n2682_, new_n2683_, new_n2684_, new_n2685_, new_n2686_, new_n2687_,
    new_n2688_, new_n2689_, new_n2690_, new_n2691_, new_n2692_, new_n2693_,
    new_n2694_, new_n2695_, new_n2696_, new_n2697_, new_n2698_, new_n2699_,
    new_n2700_, new_n2701_, new_n2702_, new_n2703_, new_n2704_, new_n2705_,
    new_n2706_, new_n2707_, new_n2708_, new_n2709_, new_n2710_, new_n2711_,
    new_n2712_, new_n2713_, new_n2714_, new_n2715_, new_n2716_, new_n2717_,
    new_n2718_, new_n2719_, new_n2720_, new_n2721_, new_n2722_, new_n2723_,
    new_n2724_, new_n2725_, new_n2726_, new_n2727_, new_n2728_, new_n2729_,
    new_n2730_, new_n2731_, new_n2732_, new_n2733_, new_n2734_, new_n2735_,
    new_n2736_, new_n2737_, new_n2738_, new_n2739_, new_n2740_, new_n2741_,
    new_n2742_, new_n2743_, new_n2744_, new_n2745_, new_n2746_, new_n2747_,
    new_n2748_, new_n2749_, new_n2750_, new_n2751_, new_n2752_, new_n2753_,
    new_n2754_, new_n2755_, new_n2756_, new_n2757_, new_n2758_, new_n2759_,
    new_n2761_, new_n2762_, new_n2763_, new_n2764_, new_n2765_, new_n2766_,
    new_n2767_, new_n2768_, new_n2769_, new_n2770_, new_n2771_, new_n2772_,
    new_n2773_, new_n2774_, new_n2775_, new_n2776_, new_n2777_, new_n2778_,
    new_n2779_, new_n2780_, new_n2781_, new_n2782_, new_n2783_, new_n2784_,
    new_n2785_, new_n2786_, new_n2787_, new_n2788_, new_n2789_, new_n2790_,
    new_n2791_, new_n2792_, new_n2793_, new_n2794_, new_n2795_, new_n2796_,
    new_n2797_, new_n2798_, new_n2799_, new_n2800_, new_n2801_, new_n2802_,
    new_n2803_, new_n2804_, new_n2805_, new_n2806_, new_n2807_, new_n2808_,
    new_n2809_, new_n2810_, new_n2811_, new_n2812_, new_n2813_, new_n2814_,
    new_n2815_, new_n2816_, new_n2817_, new_n2818_, new_n2819_, new_n2820_,
    new_n2821_, new_n2822_, new_n2823_, new_n2824_, new_n2825_, new_n2826_,
    new_n2827_, new_n2828_, new_n2829_, new_n2830_, new_n2831_, new_n2832_,
    new_n2833_, new_n2834_, new_n2835_, new_n2836_, new_n2837_, new_n2838_,
    new_n2839_, new_n2840_, new_n2841_, new_n2842_, new_n2843_, new_n2844_,
    new_n2845_, new_n2846_, new_n2848_, new_n2849_, new_n2850_, new_n2851_,
    new_n2852_, new_n2853_, new_n2854_, new_n2855_, new_n2856_, new_n2857_,
    new_n2858_, new_n2859_, new_n2860_, new_n2861_, new_n2862_, new_n2863_,
    new_n2864_, new_n2865_, new_n2866_, new_n2867_, new_n2868_, new_n2869_,
    new_n2870_, new_n2871_, new_n2872_, new_n2873_, new_n2874_, new_n2875_,
    new_n2876_, new_n2877_, new_n2878_, new_n2879_, new_n2880_, new_n2881_,
    new_n2882_, new_n2883_, new_n2884_, new_n2885_, new_n2886_, new_n2887_,
    new_n2888_, new_n2889_, new_n2890_, new_n2891_, new_n2892_, new_n2893_,
    new_n2894_, new_n2895_, new_n2896_, new_n2897_, new_n2898_, new_n2899_,
    new_n2900_, new_n2901_, new_n2902_, new_n2903_, new_n2904_, new_n2905_,
    new_n2906_, new_n2907_, new_n2908_, new_n2909_, new_n2910_, new_n2911_,
    new_n2912_, new_n2913_, new_n2914_, new_n2915_, new_n2916_, new_n2917_,
    new_n2918_, new_n2919_, new_n2920_, new_n2921_, new_n2922_, new_n2923_,
    new_n2924_, new_n2925_, new_n2926_, new_n2927_, new_n2928_, new_n2929_,
    new_n2930_, new_n2931_, new_n2932_, new_n2933_, new_n2935_, new_n2936_,
    new_n2937_, new_n2938_, new_n2939_, new_n2940_, new_n2941_, new_n2942_,
    new_n2943_, new_n2944_, new_n2945_, new_n2946_, new_n2947_, new_n2948_,
    new_n2949_, new_n2950_, new_n2951_, new_n2952_, new_n2953_, new_n2954_,
    new_n2955_, new_n2956_, new_n2957_, new_n2958_, new_n2959_, new_n2960_,
    new_n2961_, new_n2962_, new_n2963_, new_n2964_, new_n2965_, new_n2966_,
    new_n2967_, new_n2968_, new_n2969_, new_n2970_, new_n2971_, new_n2972_,
    new_n2973_, new_n2974_, new_n2975_, new_n2976_, new_n2977_, new_n2978_,
    new_n2979_, new_n2980_, new_n2981_, new_n2982_, new_n2983_, new_n2984_,
    new_n2985_, new_n2986_, new_n2987_, new_n2988_, new_n2989_, new_n2990_,
    new_n2991_, new_n2992_, new_n2993_, new_n2994_, new_n2995_, new_n2996_,
    new_n2997_, new_n2998_, new_n2999_, new_n3000_, new_n3001_, new_n3002_,
    new_n3003_, new_n3004_, new_n3005_, new_n3006_, new_n3007_, new_n3008_,
    new_n3009_, new_n3010_, new_n3011_, new_n3012_, new_n3013_, new_n3014_,
    new_n3015_, new_n3016_, new_n3017_, new_n3018_, new_n3019_, new_n3020_,
    new_n3022_, new_n3023_, new_n3024_, new_n3025_, new_n3026_, new_n3027_,
    new_n3028_, new_n3029_, new_n3030_, new_n3031_, new_n3032_, new_n3033_,
    new_n3034_, new_n3035_, new_n3036_, new_n3037_, new_n3038_, new_n3039_,
    new_n3040_, new_n3041_, new_n3042_, new_n3043_, new_n3044_, new_n3045_,
    new_n3046_, new_n3047_, new_n3048_, new_n3049_, new_n3050_, new_n3051_,
    new_n3052_, new_n3053_, new_n3054_, new_n3055_, new_n3056_, new_n3057_,
    new_n3058_, new_n3059_, new_n3060_, new_n3061_, new_n3062_, new_n3063_,
    new_n3064_, new_n3065_, new_n3066_, new_n3067_, new_n3068_, new_n3069_,
    new_n3070_, new_n3071_, new_n3072_, new_n3073_, new_n3074_, new_n3075_,
    new_n3076_, new_n3077_, new_n3078_, new_n3079_, new_n3080_, new_n3081_,
    new_n3082_, new_n3083_, new_n3084_, new_n3085_, new_n3086_, new_n3087_,
    new_n3088_, new_n3089_, new_n3090_, new_n3091_, new_n3092_, new_n3093_,
    new_n3094_, new_n3095_, new_n3096_, new_n3097_, new_n3098_, new_n3099_,
    new_n3100_, new_n3101_, new_n3102_, new_n3103_, new_n3104_, new_n3105_,
    new_n3106_, new_n3107_, new_n3109_, new_n3110_, new_n3111_, new_n3112_,
    new_n3113_, new_n3114_, new_n3115_, new_n3116_, new_n3117_, new_n3118_,
    new_n3119_, new_n3120_, new_n3121_, new_n3122_, new_n3123_, new_n3124_,
    new_n3125_, new_n3126_, new_n3127_, new_n3128_, new_n3129_, new_n3130_,
    new_n3131_, new_n3132_, new_n3133_, new_n3134_, new_n3135_, new_n3136_,
    new_n3137_, new_n3138_, new_n3139_, new_n3140_, new_n3141_, new_n3142_,
    new_n3143_, new_n3144_, new_n3145_, new_n3146_, new_n3147_, new_n3148_,
    new_n3149_, new_n3150_, new_n3151_, new_n3152_, new_n3153_, new_n3154_,
    new_n3155_, new_n3156_, new_n3157_, new_n3158_, new_n3159_, new_n3160_,
    new_n3161_, new_n3162_, new_n3163_, new_n3164_, new_n3165_, new_n3166_,
    new_n3167_, new_n3168_, new_n3169_, new_n3170_, new_n3171_, new_n3172_,
    new_n3173_, new_n3174_, new_n3175_, new_n3176_, new_n3177_, new_n3178_,
    new_n3179_, new_n3180_, new_n3181_, new_n3182_, new_n3183_, new_n3184_,
    new_n3185_, new_n3186_, new_n3187_, new_n3188_, new_n3189_, new_n3190_,
    new_n3191_, new_n3192_, new_n3193_, new_n3194_, new_n3196_, new_n3197_,
    new_n3198_, new_n3199_, new_n3200_, new_n3201_, new_n3202_, new_n3203_,
    new_n3204_, new_n3205_, new_n3206_, new_n3207_, new_n3208_, new_n3209_,
    new_n3210_, new_n3211_, new_n3212_, new_n3213_, new_n3214_, new_n3215_,
    new_n3216_, new_n3217_, new_n3218_, new_n3219_, new_n3220_, new_n3221_,
    new_n3222_, new_n3223_, new_n3224_, new_n3225_, new_n3226_, new_n3227_,
    new_n3228_, new_n3229_, new_n3230_, new_n3231_, new_n3232_, new_n3233_,
    new_n3234_, new_n3235_, new_n3236_, new_n3237_, new_n3238_, new_n3239_,
    new_n3240_, new_n3241_, new_n3242_, new_n3243_, new_n3244_, new_n3245_,
    new_n3246_, new_n3247_, new_n3248_, new_n3249_, new_n3250_, new_n3251_,
    new_n3252_, new_n3253_, new_n3254_, new_n3255_, new_n3256_, new_n3257_,
    new_n3258_, new_n3259_, new_n3260_, new_n3261_, new_n3262_, new_n3263_,
    new_n3264_, new_n3265_, new_n3266_, new_n3267_, new_n3268_, new_n3269_,
    new_n3270_, new_n3271_, new_n3272_, new_n3273_, new_n3274_, new_n3275_,
    new_n3276_, new_n3277_, new_n3278_, new_n3279_, new_n3280_, new_n3281_,
    new_n3283_, new_n3284_, new_n3285_, new_n3286_, new_n3287_, new_n3288_,
    new_n3289_, new_n3290_, new_n3291_, new_n3292_, new_n3293_, new_n3294_,
    new_n3295_, new_n3296_, new_n3297_, new_n3298_, new_n3299_, new_n3300_,
    new_n3301_, new_n3302_, new_n3303_, new_n3304_, new_n3305_, new_n3306_,
    new_n3307_, new_n3308_, new_n3309_, new_n3310_, new_n3311_, new_n3312_,
    new_n3313_, new_n3314_, new_n3315_, new_n3316_, new_n3317_, new_n3318_,
    new_n3319_, new_n3320_, new_n3321_, new_n3322_, new_n3323_, new_n3324_,
    new_n3325_, new_n3326_, new_n3327_, new_n3328_, new_n3329_, new_n3330_,
    new_n3331_, new_n3332_, new_n3333_, new_n3334_, new_n3335_, new_n3336_,
    new_n3337_, new_n3338_, new_n3339_, new_n3340_, new_n3341_, new_n3342_,
    new_n3343_, new_n3344_, new_n3345_, new_n3346_, new_n3347_, new_n3348_,
    new_n3349_, new_n3350_, new_n3351_, new_n3352_, new_n3353_, new_n3354_,
    new_n3355_, new_n3356_, new_n3357_, new_n3358_, new_n3359_, new_n3360_,
    new_n3361_, new_n3362_, new_n3363_, new_n3364_, new_n3365_, new_n3366_,
    new_n3367_, new_n3368_, new_n3370_, new_n3371_, new_n3372_, new_n3373_,
    new_n3374_, new_n3375_, new_n3376_, new_n3377_, new_n3378_, new_n3379_,
    new_n3380_, new_n3381_, new_n3382_, new_n3383_, new_n3384_, new_n3385_,
    new_n3386_, new_n3387_, new_n3388_, new_n3389_, new_n3390_, new_n3391_,
    new_n3392_, new_n3393_, new_n3394_, new_n3395_, new_n3396_, new_n3397_,
    new_n3398_, new_n3399_, new_n3400_, new_n3401_, new_n3402_, new_n3403_,
    new_n3404_, new_n3405_, new_n3406_, new_n3407_, new_n3408_, new_n3409_,
    new_n3410_, new_n3411_, new_n3412_, new_n3413_, new_n3414_, new_n3415_,
    new_n3416_, new_n3417_, new_n3418_, new_n3419_, new_n3420_, new_n3421_,
    new_n3422_, new_n3423_, new_n3424_, new_n3425_, new_n3426_, new_n3427_,
    new_n3428_, new_n3429_, new_n3430_, new_n3431_, new_n3432_, new_n3433_,
    new_n3434_, new_n3435_, new_n3436_, new_n3437_, new_n3438_, new_n3439_,
    new_n3440_, new_n3441_, new_n3442_, new_n3443_, new_n3444_, new_n3445_,
    new_n3446_, new_n3447_, new_n3448_, new_n3449_, new_n3450_, new_n3451_,
    new_n3452_, new_n3453_, new_n3454_, new_n3455_, new_n3457_, new_n3458_,
    new_n3459_, new_n3460_, new_n3461_, new_n3462_, new_n3463_, new_n3464_,
    new_n3465_, new_n3466_, new_n3467_, new_n3468_, new_n3469_, new_n3470_,
    new_n3471_, new_n3472_, new_n3473_, new_n3474_, new_n3475_, new_n3476_,
    new_n3477_, new_n3478_, new_n3479_, new_n3480_, new_n3481_, new_n3482_,
    new_n3483_, new_n3484_, new_n3485_, new_n3486_, new_n3487_, new_n3488_,
    new_n3489_, new_n3490_, new_n3491_, new_n3492_, new_n3493_, new_n3494_,
    new_n3495_, new_n3496_, new_n3497_, new_n3498_, new_n3499_, new_n3500_,
    new_n3501_, new_n3502_, new_n3503_, new_n3504_, new_n3505_, new_n3506_,
    new_n3507_, new_n3508_, new_n3509_, new_n3510_, new_n3511_, new_n3512_,
    new_n3513_, new_n3514_, new_n3515_, new_n3516_, new_n3517_, new_n3518_,
    new_n3519_, new_n3520_, new_n3521_, new_n3522_, new_n3523_, new_n3524_,
    new_n3525_, new_n3526_, new_n3527_, new_n3528_, new_n3529_, new_n3530_,
    new_n3531_, new_n3532_, new_n3533_, new_n3534_, new_n3535_, new_n3536_,
    new_n3537_, new_n3538_, new_n3539_, new_n3540_, new_n3541_, new_n3542_,
    new_n3544_, new_n3545_, new_n3546_, new_n3547_, new_n3548_, new_n3549_,
    new_n3550_, new_n3551_, new_n3552_, new_n3553_, new_n3554_, new_n3555_,
    new_n3556_, new_n3557_, new_n3558_, new_n3559_, new_n3560_, new_n3561_,
    new_n3562_, new_n3563_, new_n3564_, new_n3565_, new_n3566_, new_n3567_,
    new_n3568_, new_n3569_, new_n3570_, new_n3571_, new_n3572_, new_n3573_,
    new_n3574_, new_n3575_, new_n3576_, new_n3577_, new_n3578_, new_n3579_,
    new_n3580_, new_n3581_, new_n3582_, new_n3583_, new_n3584_, new_n3585_,
    new_n3586_, new_n3587_, new_n3588_, new_n3589_, new_n3590_, new_n3591_,
    new_n3592_, new_n3593_, new_n3594_, new_n3595_, new_n3596_, new_n3597_,
    new_n3598_, new_n3599_, new_n3600_, new_n3601_, new_n3602_, new_n3603_,
    new_n3604_, new_n3605_, new_n3606_, new_n3607_, new_n3608_, new_n3609_,
    new_n3610_, new_n3611_, new_n3612_, new_n3613_, new_n3614_, new_n3615_,
    new_n3616_, new_n3617_, new_n3618_, new_n3619_, new_n3620_, new_n3621_,
    new_n3622_, new_n3623_, new_n3624_, new_n3625_, new_n3626_, new_n3627_,
    new_n3628_, new_n3629_, new_n3631_, new_n3632_, new_n3633_, new_n3634_,
    new_n3635_, new_n3636_, new_n3637_, new_n3638_, new_n3639_, new_n3640_,
    new_n3641_, new_n3642_, new_n3643_, new_n3644_, new_n3645_, new_n3646_,
    new_n3647_, new_n3648_, new_n3649_, new_n3650_, new_n3651_, new_n3652_,
    new_n3653_, new_n3654_, new_n3655_, new_n3656_, new_n3657_, new_n3658_,
    new_n3659_, new_n3660_, new_n3661_, new_n3662_, new_n3663_, new_n3664_,
    new_n3665_, new_n3666_, new_n3667_, new_n3668_, new_n3669_, new_n3670_,
    new_n3671_, new_n3672_, new_n3673_, new_n3674_, new_n3675_, new_n3676_,
    new_n3677_, new_n3678_, new_n3679_, new_n3680_, new_n3681_, new_n3682_,
    new_n3683_, new_n3684_, new_n3685_, new_n3686_, new_n3687_, new_n3688_,
    new_n3689_, new_n3690_, new_n3691_, new_n3692_, new_n3693_, new_n3694_,
    new_n3695_, new_n3696_, new_n3697_, new_n3698_, new_n3699_, new_n3700_,
    new_n3701_, new_n3702_, new_n3703_, new_n3704_, new_n3705_, new_n3706_,
    new_n3707_, new_n3708_, new_n3709_, new_n3710_, new_n3711_, new_n3712_,
    new_n3713_, new_n3714_, new_n3715_, new_n3716_, new_n3718_, new_n3719_,
    new_n3720_, new_n3721_, new_n3722_, new_n3723_, new_n3724_, new_n3725_,
    new_n3726_, new_n3727_, new_n3728_, new_n3729_, new_n3730_, new_n3731_,
    new_n3732_, new_n3733_, new_n3734_, new_n3735_, new_n3736_, new_n3737_,
    new_n3738_, new_n3739_, new_n3740_, new_n3741_, new_n3742_, new_n3743_,
    new_n3744_, new_n3745_, new_n3746_, new_n3747_, new_n3748_, new_n3749_,
    new_n3750_, new_n3751_, new_n3752_, new_n3753_, new_n3754_, new_n3755_,
    new_n3756_, new_n3757_, new_n3758_, new_n3759_, new_n3760_, new_n3761_,
    new_n3762_, new_n3763_, new_n3764_, new_n3765_, new_n3766_, new_n3767_,
    new_n3768_, new_n3769_, new_n3770_, new_n3771_, new_n3772_, new_n3773_,
    new_n3774_, new_n3775_, new_n3776_, new_n3777_, new_n3778_, new_n3779_,
    new_n3780_, new_n3781_, new_n3782_, new_n3783_, new_n3784_, new_n3785_,
    new_n3786_, new_n3787_, new_n3788_, new_n3789_, new_n3790_, new_n3791_,
    new_n3792_, new_n3793_, new_n3794_, new_n3795_, new_n3796_, new_n3797_,
    new_n3798_, new_n3799_, new_n3800_, new_n3801_, new_n3802_, new_n3803_,
    new_n3805_, new_n3806_, new_n3807_, new_n3808_, new_n3809_, new_n3810_,
    new_n3811_, new_n3812_, new_n3813_, new_n3814_, new_n3815_, new_n3816_,
    new_n3817_, new_n3818_, new_n3819_, new_n3820_, new_n3821_, new_n3822_,
    new_n3823_, new_n3824_, new_n3825_, new_n3826_, new_n3827_, new_n3828_,
    new_n3829_, new_n3830_, new_n3831_, new_n3832_, new_n3833_, new_n3834_,
    new_n3835_, new_n3836_, new_n3837_, new_n3838_, new_n3839_, new_n3840_,
    new_n3841_, new_n3842_, new_n3843_, new_n3844_, new_n3845_, new_n3846_,
    new_n3847_, new_n3848_, new_n3849_, new_n3850_, new_n3851_, new_n3852_,
    new_n3853_, new_n3854_, new_n3855_, new_n3856_, new_n3857_, new_n3858_,
    new_n3859_, new_n3860_, new_n3861_, new_n3862_, new_n3863_, new_n3864_,
    new_n3865_, new_n3866_, new_n3867_, new_n3868_, new_n3869_, new_n3870_,
    new_n3871_, new_n3872_, new_n3873_, new_n3874_, new_n3875_, new_n3876_,
    new_n3877_, new_n3878_, new_n3879_, new_n3880_, new_n3881_, new_n3882_,
    new_n3883_, new_n3884_, new_n3885_, new_n3886_, new_n3887_, new_n3888_,
    new_n3889_, new_n3890_, new_n3892_, new_n3893_, new_n3894_, new_n3895_,
    new_n3896_, new_n3897_, new_n3898_, new_n3899_, new_n3900_, new_n3901_,
    new_n3902_, new_n3903_, new_n3904_, new_n3905_, new_n3906_, new_n3907_,
    new_n3908_, new_n3909_, new_n3910_, new_n3911_, new_n3912_, new_n3913_,
    new_n3914_, new_n3915_, new_n3916_, new_n3917_, new_n3918_, new_n3919_,
    new_n3920_, new_n3921_, new_n3922_, new_n3923_, new_n3924_, new_n3925_,
    new_n3926_, new_n3927_, new_n3928_, new_n3929_, new_n3930_, new_n3931_,
    new_n3932_, new_n3933_, new_n3934_, new_n3935_, new_n3936_, new_n3937_,
    new_n3938_, new_n3939_, new_n3940_, new_n3941_, new_n3942_, new_n3943_,
    new_n3944_, new_n3945_, new_n3946_, new_n3947_, new_n3948_, new_n3949_,
    new_n3950_, new_n3951_, new_n3952_, new_n3953_, new_n3954_, new_n3955_,
    new_n3956_, new_n3957_, new_n3958_, new_n3959_, new_n3960_, new_n3961_,
    new_n3962_, new_n3963_, new_n3964_, new_n3965_, new_n3966_, new_n3967_,
    new_n3968_, new_n3969_, new_n3970_, new_n3971_, new_n3972_, new_n3973_,
    new_n3974_, new_n3975_, new_n3976_, new_n3977_, new_n3979_, new_n3980_,
    new_n3981_, new_n3982_, new_n3983_, new_n3984_, new_n3985_, new_n3986_,
    new_n3987_, new_n3988_, new_n3989_, new_n3990_, new_n3991_, new_n3992_,
    new_n3993_, new_n3994_, new_n3995_, new_n3996_, new_n3997_, new_n3998_,
    new_n3999_, new_n4000_, new_n4001_, new_n4002_, new_n4003_, new_n4004_,
    new_n4005_, new_n4006_, new_n4007_, new_n4008_, new_n4009_, new_n4010_,
    new_n4011_, new_n4012_, new_n4013_, new_n4014_, new_n4015_, new_n4016_,
    new_n4017_, new_n4018_, new_n4019_, new_n4020_, new_n4021_, new_n4022_,
    new_n4023_, new_n4024_, new_n4025_, new_n4026_, new_n4027_, new_n4028_,
    new_n4029_, new_n4030_, new_n4031_, new_n4032_, new_n4033_, new_n4034_,
    new_n4035_, new_n4036_, new_n4037_, new_n4038_, new_n4039_, new_n4040_,
    new_n4041_, new_n4042_, new_n4043_, new_n4044_, new_n4045_, new_n4046_,
    new_n4047_, new_n4048_, new_n4049_, new_n4050_, new_n4051_, new_n4052_,
    new_n4053_, new_n4054_, new_n4055_, new_n4056_, new_n4057_, new_n4058_,
    new_n4059_, new_n4060_, new_n4061_, new_n4062_, new_n4063_, new_n4064_,
    new_n4066_, new_n4067_, new_n4068_, new_n4069_, new_n4070_, new_n4071_,
    new_n4072_, new_n4073_, new_n4074_, new_n4075_, new_n4076_, new_n4077_,
    new_n4078_, new_n4079_, new_n4080_, new_n4081_, new_n4082_, new_n4083_,
    new_n4084_, new_n4085_, new_n4086_, new_n4087_, new_n4088_, new_n4089_,
    new_n4090_, new_n4091_, new_n4092_, new_n4093_, new_n4094_, new_n4095_,
    new_n4096_, new_n4097_, new_n4098_, new_n4099_, new_n4100_, new_n4101_,
    new_n4102_, new_n4103_, new_n4104_, new_n4105_, new_n4106_, new_n4107_,
    new_n4108_, new_n4109_, new_n4110_, new_n4111_, new_n4112_, new_n4113_,
    new_n4114_, new_n4115_, new_n4116_, new_n4117_, new_n4118_, new_n4119_,
    new_n4120_, new_n4121_, new_n4122_, new_n4123_, new_n4124_, new_n4125_,
    new_n4126_, new_n4127_, new_n4128_, new_n4129_, new_n4130_, new_n4131_,
    new_n4132_, new_n4133_, new_n4134_, new_n4135_, new_n4136_, new_n4137_,
    new_n4138_, new_n4139_, new_n4140_, new_n4141_, new_n4142_, new_n4143_,
    new_n4144_, new_n4145_, new_n4146_, new_n4147_, new_n4148_, new_n4149_,
    new_n4150_, new_n4151_, new_n4153_, new_n4154_, new_n4155_, new_n4156_,
    new_n4157_, new_n4158_, new_n4159_, new_n4160_, new_n4161_, new_n4162_,
    new_n4163_, new_n4164_, new_n4165_, new_n4166_, new_n4167_, new_n4168_,
    new_n4169_, new_n4170_, new_n4171_, new_n4172_, new_n4173_, new_n4174_,
    new_n4175_, new_n4176_, new_n4177_, new_n4178_, new_n4179_, new_n4180_,
    new_n4181_, new_n4182_, new_n4183_, new_n4184_, new_n4185_, new_n4186_,
    new_n4187_, new_n4188_, new_n4189_, new_n4190_, new_n4191_, new_n4192_,
    new_n4193_, new_n4194_, new_n4195_, new_n4196_, new_n4197_, new_n4198_,
    new_n4199_, new_n4200_, new_n4201_, new_n4202_, new_n4203_, new_n4204_,
    new_n4205_, new_n4206_, new_n4207_, new_n4208_, new_n4209_, new_n4210_,
    new_n4211_, new_n4212_, new_n4213_, new_n4214_, new_n4215_, new_n4216_,
    new_n4217_, new_n4218_, new_n4219_, new_n4220_, new_n4221_, new_n4222_,
    new_n4223_, new_n4224_, new_n4225_, new_n4226_, new_n4227_, new_n4228_,
    new_n4229_, new_n4230_, new_n4231_, new_n4232_, new_n4233_, new_n4234_,
    new_n4235_, new_n4236_, new_n4237_, new_n4238_, new_n4240_, new_n4241_,
    new_n4242_, new_n4243_, new_n4244_, new_n4245_, new_n4246_, new_n4247_,
    new_n4248_, new_n4249_, new_n4250_, new_n4251_, new_n4252_, new_n4253_,
    new_n4254_, new_n4255_, new_n4256_, new_n4257_, new_n4258_, new_n4259_,
    new_n4260_, new_n4261_, new_n4262_, new_n4263_, new_n4264_, new_n4265_,
    new_n4266_, new_n4267_, new_n4268_, new_n4269_, new_n4270_, new_n4271_,
    new_n4272_, new_n4273_, new_n4274_, new_n4275_, new_n4276_, new_n4277_,
    new_n4278_, new_n4279_, new_n4280_, new_n4281_, new_n4282_, new_n4283_,
    new_n4284_, new_n4285_, new_n4286_, new_n4287_, new_n4288_, new_n4289_,
    new_n4290_, new_n4291_, new_n4292_, new_n4293_, new_n4294_, new_n4295_,
    new_n4296_, new_n4297_, new_n4298_, new_n4299_, new_n4300_, new_n4301_,
    new_n4302_, new_n4303_, new_n4304_, new_n4305_, new_n4306_, new_n4307_,
    new_n4308_, new_n4309_, new_n4310_, new_n4311_, new_n4312_, new_n4313_,
    new_n4314_, new_n4315_, new_n4316_, new_n4317_, new_n4318_, new_n4319_,
    new_n4320_, new_n4321_, new_n4322_, new_n4323_, new_n4324_, new_n4325_,
    new_n4327_, new_n4328_, new_n4329_, new_n4330_, new_n4331_, new_n4332_,
    new_n4333_, new_n4334_, new_n4335_, new_n4336_, new_n4337_, new_n4338_,
    new_n4339_, new_n4340_, new_n4341_, new_n4342_, new_n4343_, new_n4344_,
    new_n4345_, new_n4346_, new_n4347_, new_n4348_, new_n4349_, new_n4350_,
    new_n4351_, new_n4352_, new_n4353_, new_n4354_, new_n4355_, new_n4356_,
    new_n4357_, new_n4358_, new_n4359_, new_n4360_, new_n4361_, new_n4362_,
    new_n4363_, new_n4364_, new_n4365_, new_n4366_, new_n4367_, new_n4368_,
    new_n4369_, new_n4370_, new_n4371_, new_n4372_, new_n4373_, new_n4374_,
    new_n4375_, new_n4376_, new_n4377_, new_n4378_, new_n4379_, new_n4380_,
    new_n4381_, new_n4382_, new_n4383_, new_n4384_, new_n4385_, new_n4386_,
    new_n4387_, new_n4388_, new_n4389_, new_n4390_, new_n4391_, new_n4392_,
    new_n4393_, new_n4394_, new_n4395_, new_n4396_, new_n4397_, new_n4398_,
    new_n4399_, new_n4400_, new_n4401_, new_n4402_, new_n4403_, new_n4404_,
    new_n4405_, new_n4406_, new_n4407_, new_n4408_, new_n4409_, new_n4410_,
    new_n4411_, new_n4412_, new_n4414_, new_n4415_, new_n4416_, new_n4417_,
    new_n4418_, new_n4419_, new_n4420_, new_n4421_, new_n4422_, new_n4423_,
    new_n4424_, new_n4425_, new_n4426_, new_n4427_, new_n4428_, new_n4429_,
    new_n4430_, new_n4431_, new_n4432_, new_n4433_, new_n4434_, new_n4435_,
    new_n4436_, new_n4437_, new_n4438_, new_n4439_, new_n4440_, new_n4441_,
    new_n4442_, new_n4443_, new_n4444_, new_n4445_, new_n4446_, new_n4447_,
    new_n4448_, new_n4449_, new_n4450_, new_n4451_, new_n4452_, new_n4453_,
    new_n4454_, new_n4455_, new_n4456_, new_n4457_, new_n4458_, new_n4459_,
    new_n4460_, new_n4461_, new_n4462_, new_n4463_, new_n4464_, new_n4465_,
    new_n4466_, new_n4467_, new_n4468_, new_n4469_, new_n4470_, new_n4471_,
    new_n4472_, new_n4473_, new_n4474_, new_n4475_, new_n4476_, new_n4477_,
    new_n4478_, new_n4479_, new_n4480_, new_n4481_, new_n4482_, new_n4483_,
    new_n4484_, new_n4485_, new_n4486_, new_n4487_, new_n4488_, new_n4489_,
    new_n4490_, new_n4491_, new_n4492_, new_n4493_, new_n4494_, new_n4495_,
    new_n4496_, new_n4497_, new_n4498_, new_n4499_, new_n4501_, new_n4502_,
    new_n4503_, new_n4504_, new_n4505_, new_n4506_, new_n4507_, new_n4508_,
    new_n4509_, new_n4510_, new_n4511_, new_n4512_, new_n4513_, new_n4514_,
    new_n4515_, new_n4516_, new_n4517_, new_n4518_, new_n4519_, new_n4520_,
    new_n4521_, new_n4522_, new_n4523_, new_n4524_, new_n4525_, new_n4526_,
    new_n4527_, new_n4528_, new_n4529_, new_n4530_, new_n4531_, new_n4532_,
    new_n4533_, new_n4534_, new_n4535_, new_n4536_, new_n4537_, new_n4538_,
    new_n4539_, new_n4540_, new_n4541_, new_n4542_, new_n4543_, new_n4544_,
    new_n4545_, new_n4546_, new_n4547_, new_n4548_, new_n4549_, new_n4550_,
    new_n4551_, new_n4552_, new_n4553_, new_n4554_, new_n4555_, new_n4556_,
    new_n4557_, new_n4558_, new_n4559_, new_n4560_, new_n4561_, new_n4562_,
    new_n4563_, new_n4564_, new_n4565_, new_n4566_, new_n4567_, new_n4568_,
    new_n4569_, new_n4570_, new_n4571_, new_n4572_, new_n4573_, new_n4574_,
    new_n4575_, new_n4576_, new_n4577_, new_n4578_, new_n4579_, new_n4580_,
    new_n4581_, new_n4582_, new_n4583_, new_n4584_, new_n4585_, new_n4586_,
    new_n4588_, new_n4589_, new_n4590_, new_n4591_, new_n4592_, new_n4593_,
    new_n4594_, new_n4595_, new_n4596_, new_n4597_, new_n4598_, new_n4599_,
    new_n4600_, new_n4601_, new_n4602_, new_n4603_, new_n4604_, new_n4605_,
    new_n4606_, new_n4607_, new_n4608_, new_n4609_, new_n4610_, new_n4611_,
    new_n4612_, new_n4613_, new_n4614_, new_n4615_, new_n4616_, new_n4617_,
    new_n4618_, new_n4619_, new_n4620_, new_n4621_, new_n4622_, new_n4623_,
    new_n4624_, new_n4625_, new_n4626_, new_n4627_, new_n4628_, new_n4629_,
    new_n4630_, new_n4631_, new_n4632_, new_n4633_, new_n4634_, new_n4635_,
    new_n4636_, new_n4637_, new_n4638_, new_n4639_, new_n4640_, new_n4641_,
    new_n4642_, new_n4643_, new_n4644_, new_n4645_, new_n4646_, new_n4647_,
    new_n4648_, new_n4649_, new_n4650_, new_n4651_, new_n4652_, new_n4653_,
    new_n4654_, new_n4655_, new_n4656_, new_n4657_, new_n4658_, new_n4659_,
    new_n4660_, new_n4661_, new_n4662_, new_n4663_, new_n4664_, new_n4665_,
    new_n4666_, new_n4667_, new_n4668_, new_n4669_, new_n4670_, new_n4671_,
    new_n4672_, new_n4673_, new_n4675_, new_n4676_, new_n4677_, new_n4678_,
    new_n4679_, new_n4680_, new_n4681_, new_n4682_, new_n4683_, new_n4684_,
    new_n4685_, new_n4686_, new_n4687_, new_n4688_, new_n4689_, new_n4690_,
    new_n4691_, new_n4692_, new_n4693_, new_n4694_, new_n4695_, new_n4696_,
    new_n4697_, new_n4698_, new_n4699_, new_n4700_, new_n4701_, new_n4702_,
    new_n4703_, new_n4704_, new_n4705_, new_n4706_, new_n4707_, new_n4708_,
    new_n4709_, new_n4710_, new_n4711_, new_n4712_, new_n4713_, new_n4714_,
    new_n4715_, new_n4716_, new_n4717_, new_n4718_, new_n4719_, new_n4720_,
    new_n4721_, new_n4722_, new_n4723_, new_n4724_, new_n4725_, new_n4726_,
    new_n4727_, new_n4728_, new_n4729_, new_n4730_, new_n4731_, new_n4732_,
    new_n4733_, new_n4734_, new_n4735_, new_n4736_, new_n4737_, new_n4738_,
    new_n4739_, new_n4740_, new_n4741_, new_n4742_, new_n4743_, new_n4744_,
    new_n4745_, new_n4746_, new_n4747_, new_n4748_, new_n4749_, new_n4750_,
    new_n4751_, new_n4752_, new_n4753_, new_n4754_, new_n4755_, new_n4756_,
    new_n4757_, new_n4758_, new_n4759_, new_n4760_, new_n4762_, new_n4763_,
    new_n4764_, new_n4765_, new_n4766_, new_n4767_, new_n4768_, new_n4769_,
    new_n4770_, new_n4771_, new_n4772_, new_n4773_, new_n4774_, new_n4775_,
    new_n4776_, new_n4777_, new_n4778_, new_n4779_, new_n4780_, new_n4781_,
    new_n4782_, new_n4783_, new_n4784_, new_n4785_, new_n4786_, new_n4787_,
    new_n4788_, new_n4789_, new_n4790_, new_n4791_, new_n4792_, new_n4793_,
    new_n4794_, new_n4795_, new_n4796_, new_n4797_, new_n4798_, new_n4799_,
    new_n4800_, new_n4801_, new_n4802_, new_n4803_, new_n4804_, new_n4805_,
    new_n4806_, new_n4807_, new_n4808_, new_n4809_, new_n4810_, new_n4811_,
    new_n4812_, new_n4813_, new_n4814_, new_n4815_, new_n4816_, new_n4817_,
    new_n4818_, new_n4819_, new_n4820_, new_n4821_, new_n4822_, new_n4823_,
    new_n4824_, new_n4825_, new_n4826_, new_n4827_, new_n4828_, new_n4829_,
    new_n4830_, new_n4831_, new_n4832_, new_n4833_, new_n4834_, new_n4835_,
    new_n4836_, new_n4837_, new_n4838_, new_n4839_, new_n4840_, new_n4841_,
    new_n4842_, new_n4843_, new_n4844_, new_n4845_, new_n4846_, new_n4847_,
    new_n4849_, new_n4850_, new_n4851_, new_n4852_, new_n4853_, new_n4854_,
    new_n4855_, new_n4856_, new_n4857_, new_n4858_, new_n4859_, new_n4860_,
    new_n4861_, new_n4862_, new_n4863_, new_n4864_, new_n4865_, new_n4866_,
    new_n4867_, new_n4868_, new_n4869_, new_n4870_, new_n4871_, new_n4872_,
    new_n4873_, new_n4874_, new_n4875_, new_n4876_, new_n4877_, new_n4878_,
    new_n4879_, new_n4880_, new_n4881_, new_n4882_, new_n4883_, new_n4884_,
    new_n4885_, new_n4886_, new_n4887_, new_n4888_, new_n4889_, new_n4890_,
    new_n4891_, new_n4892_, new_n4893_, new_n4894_, new_n4895_, new_n4896_,
    new_n4897_, new_n4898_, new_n4899_, new_n4900_, new_n4901_, new_n4902_,
    new_n4903_, new_n4904_, new_n4905_, new_n4906_, new_n4907_, new_n4908_,
    new_n4909_, new_n4910_, new_n4911_, new_n4912_, new_n4913_, new_n4914_,
    new_n4915_, new_n4916_, new_n4917_, new_n4918_, new_n4919_, new_n4920_,
    new_n4921_, new_n4922_, new_n4923_, new_n4924_, new_n4925_, new_n4926_,
    new_n4927_, new_n4928_, new_n4929_, new_n4930_, new_n4931_, new_n4932_,
    new_n4933_, new_n4934_, new_n4936_, new_n4937_, new_n4938_, new_n4939_,
    new_n4940_, new_n4941_, new_n4942_, new_n4943_, new_n4944_, new_n4945_,
    new_n4946_, new_n4947_, new_n4948_, new_n4949_, new_n4950_, new_n4951_,
    new_n4952_, new_n4953_, new_n4954_, new_n4955_, new_n4956_, new_n4957_,
    new_n4958_, new_n4959_, new_n4960_, new_n4961_, new_n4962_, new_n4963_,
    new_n4964_, new_n4965_, new_n4966_, new_n4967_, new_n4968_, new_n4969_,
    new_n4970_, new_n4971_, new_n4972_, new_n4973_, new_n4974_, new_n4975_,
    new_n4976_, new_n4977_, new_n4978_, new_n4979_, new_n4980_, new_n4981_,
    new_n4982_, new_n4983_, new_n4984_, new_n4985_, new_n4986_, new_n4987_,
    new_n4988_, new_n4989_, new_n4990_, new_n4991_, new_n4992_, new_n4993_,
    new_n4994_, new_n4995_, new_n4996_, new_n4997_, new_n4998_, new_n4999_,
    new_n5000_, new_n5001_, new_n5002_, new_n5003_, new_n5004_, new_n5005_,
    new_n5006_, new_n5007_, new_n5008_, new_n5009_, new_n5010_, new_n5011_,
    new_n5012_, new_n5013_, new_n5014_, new_n5015_, new_n5016_, new_n5017_,
    new_n5018_, new_n5019_, new_n5020_, new_n5021_, new_n5023_, new_n5024_,
    new_n5025_, new_n5026_, new_n5027_, new_n5028_, new_n5029_, new_n5030_,
    new_n5031_, new_n5032_, new_n5033_, new_n5034_, new_n5035_, new_n5036_,
    new_n5037_, new_n5038_, new_n5039_, new_n5040_, new_n5041_, new_n5042_,
    new_n5043_, new_n5044_, new_n5045_, new_n5046_, new_n5047_, new_n5048_,
    new_n5049_, new_n5050_, new_n5051_, new_n5052_, new_n5053_, new_n5054_,
    new_n5055_, new_n5056_, new_n5057_, new_n5058_, new_n5059_, new_n5060_,
    new_n5061_, new_n5062_, new_n5063_, new_n5064_, new_n5065_, new_n5066_,
    new_n5067_, new_n5068_, new_n5069_, new_n5070_, new_n5071_, new_n5072_,
    new_n5073_, new_n5074_, new_n5075_, new_n5076_, new_n5077_, new_n5078_,
    new_n5079_, new_n5080_, new_n5081_, new_n5082_, new_n5083_, new_n5084_,
    new_n5085_, new_n5086_, new_n5087_, new_n5088_, new_n5089_, new_n5090_,
    new_n5091_, new_n5092_, new_n5093_, new_n5094_, new_n5095_, new_n5096_,
    new_n5097_, new_n5098_, new_n5099_, new_n5100_, new_n5101_, new_n5102_,
    new_n5103_, new_n5104_, new_n5105_, new_n5106_, new_n5107_, new_n5108_,
    new_n5110_, new_n5111_, new_n5112_, new_n5113_, new_n5114_, new_n5115_,
    new_n5116_, new_n5117_, new_n5118_, new_n5119_, new_n5120_, new_n5121_,
    new_n5122_, new_n5123_, new_n5124_, new_n5125_, new_n5126_, new_n5127_,
    new_n5128_, new_n5129_, new_n5130_, new_n5131_, new_n5132_, new_n5133_,
    new_n5134_, new_n5135_, new_n5136_, new_n5137_, new_n5138_, new_n5139_,
    new_n5140_, new_n5141_, new_n5142_, new_n5143_, new_n5144_, new_n5145_,
    new_n5146_, new_n5147_, new_n5148_, new_n5149_, new_n5150_, new_n5151_,
    new_n5152_, new_n5153_, new_n5154_, new_n5155_, new_n5156_, new_n5157_,
    new_n5158_, new_n5159_, new_n5160_, new_n5161_, new_n5162_, new_n5163_,
    new_n5164_, new_n5165_, new_n5166_, new_n5167_, new_n5168_, new_n5169_,
    new_n5170_, new_n5171_, new_n5172_, new_n5173_, new_n5174_, new_n5175_,
    new_n5176_, new_n5177_, new_n5178_, new_n5179_, new_n5180_, new_n5181_,
    new_n5182_, new_n5183_, new_n5184_, new_n5185_, new_n5186_, new_n5187_,
    new_n5188_, new_n5189_, new_n5190_, new_n5191_, new_n5192_, new_n5193_,
    new_n5194_, new_n5195_, new_n5197_, new_n5198_, new_n5199_, new_n5200_,
    new_n5201_, new_n5202_, new_n5203_, new_n5204_, new_n5205_, new_n5206_,
    new_n5207_, new_n5208_, new_n5209_, new_n5210_, new_n5211_, new_n5212_,
    new_n5213_, new_n5214_, new_n5215_, new_n5216_, new_n5217_, new_n5218_,
    new_n5219_, new_n5220_, new_n5221_, new_n5222_, new_n5223_, new_n5224_,
    new_n5225_, new_n5226_, new_n5227_, new_n5228_, new_n5229_, new_n5230_,
    new_n5231_, new_n5232_, new_n5233_, new_n5234_, new_n5235_, new_n5236_,
    new_n5237_, new_n5238_, new_n5239_, new_n5240_, new_n5241_, new_n5242_,
    new_n5243_, new_n5244_, new_n5245_, new_n5246_, new_n5247_, new_n5248_,
    new_n5249_, new_n5250_, new_n5251_, new_n5252_, new_n5253_, new_n5254_,
    new_n5255_, new_n5256_, new_n5257_, new_n5258_, new_n5259_, new_n5260_,
    new_n5261_, new_n5262_, new_n5263_, new_n5264_, new_n5265_, new_n5266_,
    new_n5267_, new_n5268_, new_n5269_, new_n5270_, new_n5271_, new_n5272_,
    new_n5273_, new_n5274_, new_n5275_, new_n5276_, new_n5277_, new_n5278_,
    new_n5279_, new_n5280_, new_n5281_, new_n5282_, new_n5284_, new_n5285_,
    new_n5286_, new_n5287_, new_n5288_, new_n5289_, new_n5290_, new_n5291_,
    new_n5292_, new_n5293_, new_n5294_, new_n5295_, new_n5296_, new_n5297_,
    new_n5298_, new_n5299_, new_n5300_, new_n5301_, new_n5302_, new_n5303_,
    new_n5304_, new_n5305_, new_n5306_, new_n5307_, new_n5308_, new_n5309_,
    new_n5310_, new_n5311_, new_n5312_, new_n5313_, new_n5314_, new_n5315_,
    new_n5316_, new_n5317_, new_n5318_, new_n5319_, new_n5320_, new_n5321_,
    new_n5322_, new_n5323_, new_n5324_, new_n5325_, new_n5326_, new_n5327_,
    new_n5328_, new_n5329_, new_n5330_, new_n5331_, new_n5332_, new_n5333_,
    new_n5334_, new_n5335_, new_n5336_, new_n5337_, new_n5338_, new_n5339_,
    new_n5340_, new_n5341_, new_n5342_, new_n5343_, new_n5344_, new_n5345_,
    new_n5346_, new_n5347_, new_n5348_, new_n5349_, new_n5350_, new_n5351_,
    new_n5352_, new_n5353_, new_n5354_, new_n5355_, new_n5356_, new_n5357_,
    new_n5358_, new_n5359_, new_n5360_, new_n5361_, new_n5362_, new_n5363_,
    new_n5364_, new_n5365_, new_n5366_, new_n5367_, new_n5368_, new_n5369_,
    new_n5371_, new_n5372_, new_n5373_, new_n5374_, new_n5375_, new_n5376_,
    new_n5377_, new_n5378_, new_n5379_, new_n5380_, new_n5381_, new_n5382_,
    new_n5383_, new_n5384_, new_n5385_, new_n5386_, new_n5387_, new_n5388_,
    new_n5389_, new_n5390_, new_n5391_, new_n5392_, new_n5393_, new_n5394_,
    new_n5395_, new_n5396_, new_n5397_, new_n5398_, new_n5399_, new_n5400_,
    new_n5401_, new_n5402_, new_n5403_, new_n5404_, new_n5405_, new_n5406_,
    new_n5407_, new_n5408_, new_n5409_, new_n5410_, new_n5411_, new_n5412_,
    new_n5413_, new_n5414_, new_n5415_, new_n5416_, new_n5417_, new_n5418_,
    new_n5419_, new_n5420_, new_n5421_, new_n5422_, new_n5423_, new_n5424_,
    new_n5425_, new_n5426_, new_n5427_, new_n5428_, new_n5429_, new_n5430_,
    new_n5431_, new_n5432_, new_n5433_, new_n5434_, new_n5435_, new_n5436_,
    new_n5437_, new_n5438_, new_n5439_, new_n5440_, new_n5441_, new_n5442_,
    new_n5443_, new_n5444_, new_n5445_, new_n5446_, new_n5447_, new_n5448_,
    new_n5449_, new_n5450_, new_n5451_, new_n5452_, new_n5453_, new_n5454_,
    new_n5455_, new_n5456_, new_n5458_, new_n5459_, new_n5460_, new_n5461_,
    new_n5462_, new_n5463_, new_n5464_, new_n5465_, new_n5466_, new_n5467_,
    new_n5468_, new_n5469_, new_n5470_, new_n5471_, new_n5472_, new_n5473_,
    new_n5474_, new_n5475_, new_n5476_, new_n5477_, new_n5478_, new_n5479_,
    new_n5480_, new_n5481_, new_n5482_, new_n5483_, new_n5484_, new_n5485_,
    new_n5486_, new_n5487_, new_n5488_, new_n5489_, new_n5490_, new_n5491_,
    new_n5492_, new_n5493_, new_n5494_, new_n5495_, new_n5496_, new_n5497_,
    new_n5498_, new_n5499_, new_n5500_, new_n5501_, new_n5502_, new_n5503_,
    new_n5504_, new_n5505_, new_n5506_, new_n5507_, new_n5508_, new_n5509_,
    new_n5510_, new_n5511_, new_n5512_, new_n5513_, new_n5514_, new_n5515_,
    new_n5516_, new_n5517_, new_n5518_, new_n5519_, new_n5520_, new_n5521_,
    new_n5522_, new_n5523_, new_n5524_, new_n5525_, new_n5526_, new_n5527_,
    new_n5528_, new_n5529_, new_n5530_, new_n5531_, new_n5532_, new_n5533_,
    new_n5534_, new_n5535_, new_n5536_, new_n5537_, new_n5538_, new_n5539_,
    new_n5540_, new_n5541_, new_n5542_, new_n5543_, new_n5545_, new_n5546_,
    new_n5547_, new_n5548_, new_n5549_, new_n5550_, new_n5551_, new_n5552_,
    new_n5553_, new_n5554_, new_n5555_, new_n5556_, new_n5557_, new_n5558_,
    new_n5559_, new_n5560_, new_n5561_, new_n5562_, new_n5563_, new_n5564_,
    new_n5565_, new_n5566_, new_n5567_, new_n5568_, new_n5569_, new_n5570_,
    new_n5571_, new_n5572_, new_n5573_, new_n5574_, new_n5575_, new_n5576_,
    new_n5577_, new_n5578_, new_n5579_, new_n5580_, new_n5581_, new_n5582_,
    new_n5583_, new_n5584_, new_n5585_, new_n5586_, new_n5587_, new_n5588_,
    new_n5589_, new_n5590_, new_n5591_, new_n5592_, new_n5593_, new_n5594_,
    new_n5595_, new_n5596_, new_n5597_, new_n5598_, new_n5599_, new_n5600_,
    new_n5601_, new_n5602_, new_n5603_, new_n5604_, new_n5605_, new_n5606_,
    new_n5607_, new_n5608_, new_n5609_, new_n5610_, new_n5611_, new_n5612_,
    new_n5613_, new_n5614_, new_n5615_, new_n5616_, new_n5617_, new_n5618_,
    new_n5619_, new_n5620_, new_n5621_, new_n5622_, new_n5623_, new_n5624_,
    new_n5625_, new_n5626_, new_n5627_, new_n5628_, new_n5629_, new_n5630_,
    new_n5632_, new_n5633_, new_n5634_, new_n5635_, new_n5636_, new_n5637_,
    new_n5638_, new_n5639_, new_n5640_, new_n5641_, new_n5642_, new_n5643_,
    new_n5644_, new_n5645_, new_n5646_, new_n5647_, new_n5648_, new_n5649_,
    new_n5650_, new_n5651_, new_n5652_, new_n5653_, new_n5654_, new_n5655_,
    new_n5656_, new_n5657_, new_n5658_, new_n5659_, new_n5660_, new_n5661_,
    new_n5662_, new_n5663_, new_n5664_, new_n5665_, new_n5666_, new_n5667_,
    new_n5668_, new_n5669_, new_n5670_, new_n5671_, new_n5672_, new_n5673_,
    new_n5674_, new_n5675_, new_n5676_, new_n5677_, new_n5678_, new_n5679_,
    new_n5680_, new_n5681_, new_n5682_, new_n5683_, new_n5684_, new_n5685_,
    new_n5686_, new_n5687_, new_n5688_, new_n5689_, new_n5690_, new_n5691_,
    new_n5692_, new_n5693_, new_n5694_, new_n5695_, new_n5696_, new_n5697_,
    new_n5698_, new_n5699_, new_n5700_, new_n5701_, new_n5702_, new_n5703_,
    new_n5704_, new_n5705_, new_n5706_, new_n5707_, new_n5708_, new_n5709_,
    new_n5710_, new_n5711_, new_n5712_, new_n5713_, new_n5714_, new_n5715_,
    new_n5716_, new_n5717_, new_n5719_, new_n5720_, new_n5721_, new_n5722_,
    new_n5723_, new_n5724_, new_n5725_, new_n5726_, new_n5727_, new_n5728_,
    new_n5729_, new_n5730_, new_n5731_, new_n5732_, new_n5733_, new_n5734_,
    new_n5735_, new_n5736_, new_n5737_, new_n5738_, new_n5739_, new_n5740_,
    new_n5741_, new_n5742_, new_n5743_, new_n5744_, new_n5745_, new_n5746_,
    new_n5747_, new_n5748_, new_n5749_, new_n5750_, new_n5751_, new_n5752_,
    new_n5753_, new_n5754_, new_n5755_, new_n5756_, new_n5757_, new_n5758_,
    new_n5759_, new_n5760_, new_n5761_, new_n5762_, new_n5763_, new_n5764_,
    new_n5765_, new_n5766_, new_n5767_, new_n5768_, new_n5769_, new_n5770_,
    new_n5771_, new_n5772_, new_n5773_, new_n5774_, new_n5775_, new_n5776_,
    new_n5777_, new_n5778_, new_n5779_, new_n5780_, new_n5781_, new_n5782_,
    new_n5783_, new_n5784_, new_n5785_, new_n5786_, new_n5787_, new_n5788_,
    new_n5789_, new_n5790_, new_n5791_, new_n5792_, new_n5793_, new_n5794_,
    new_n5795_, new_n5796_, new_n5797_, new_n5798_, new_n5799_, new_n5800_,
    new_n5801_, new_n5802_, new_n5803_, new_n5804_, new_n5806_, new_n5807_,
    new_n5808_, new_n5809_, new_n5810_, new_n5811_, new_n5812_, new_n5813_,
    new_n5814_, new_n5815_, new_n5816_, new_n5817_, new_n5818_, new_n5819_,
    new_n5820_, new_n5821_, new_n5822_, new_n5823_, new_n5824_, new_n5825_,
    new_n5826_, new_n5827_, new_n5828_, new_n5829_, new_n5830_, new_n5831_,
    new_n5832_, new_n5833_, new_n5834_, new_n5835_, new_n5836_, new_n5837_,
    new_n5838_, new_n5839_, new_n5840_, new_n5841_, new_n5842_, new_n5843_,
    new_n5844_, new_n5845_, new_n5846_, new_n5847_, new_n5848_, new_n5849_,
    new_n5850_, new_n5851_, new_n5852_, new_n5853_, new_n5854_, new_n5855_,
    new_n5856_, new_n5857_, new_n5858_, new_n5859_, new_n5860_, new_n5861_,
    new_n5862_, new_n5863_, new_n5864_, new_n5865_, new_n5866_, new_n5867_,
    new_n5868_, new_n5869_, new_n5870_, new_n5871_, new_n5872_, new_n5873_,
    new_n5874_, new_n5875_, new_n5876_, new_n5877_, new_n5878_, new_n5879_,
    new_n5880_, new_n5881_, new_n5882_, new_n5883_, new_n5884_, new_n5885_,
    new_n5886_, new_n5887_, new_n5888_, new_n5889_, new_n5890_, new_n5891_,
    new_n5893_, new_n5894_, new_n5895_, new_n5896_, new_n5897_, new_n5898_,
    new_n5899_, new_n5900_, new_n5901_, new_n5902_, new_n5903_, new_n5904_,
    new_n5905_, new_n5906_, new_n5907_, new_n5908_, new_n5909_, new_n5910_,
    new_n5911_, new_n5912_, new_n5913_, new_n5914_, new_n5915_, new_n5916_,
    new_n5917_, new_n5918_, new_n5919_, new_n5920_, new_n5921_, new_n5922_,
    new_n5923_, new_n5924_, new_n5925_, new_n5926_, new_n5927_, new_n5928_,
    new_n5929_, new_n5930_, new_n5931_, new_n5932_, new_n5933_, new_n5934_,
    new_n5935_, new_n5936_, new_n5937_, new_n5938_, new_n5939_, new_n5940_,
    new_n5941_, new_n5942_, new_n5943_, new_n5944_, new_n5945_, new_n5946_,
    new_n5947_, new_n5948_, new_n5949_, new_n5950_, new_n5951_, new_n5952_,
    new_n5953_, new_n5954_, new_n5955_, new_n5956_, new_n5957_, new_n5958_,
    new_n5959_, new_n5960_, new_n5961_, new_n5962_, new_n5963_, new_n5964_,
    new_n5965_, new_n5966_, new_n5967_, new_n5968_, new_n5969_, new_n5970_,
    new_n5971_, new_n5972_, new_n5973_, new_n5974_, new_n5975_, new_n5976_,
    new_n5977_, new_n5978_, new_n5980_, new_n5981_, new_n5982_, new_n5983_,
    new_n5984_, new_n5985_, new_n5986_, new_n5987_, new_n5988_, new_n5989_,
    new_n5990_, new_n5991_, new_n5992_, new_n5993_, new_n5994_, new_n5995_,
    new_n5996_, new_n5997_, new_n5998_, new_n5999_, new_n6000_, new_n6001_,
    new_n6002_, new_n6003_, new_n6004_, new_n6005_, new_n6006_, new_n6007_,
    new_n6008_, new_n6009_, new_n6010_, new_n6011_, new_n6012_, new_n6013_,
    new_n6014_, new_n6015_, new_n6016_, new_n6017_, new_n6018_, new_n6019_,
    new_n6020_, new_n6021_, new_n6022_, new_n6023_, new_n6024_, new_n6025_,
    new_n6026_, new_n6027_, new_n6028_, new_n6029_, new_n6030_, new_n6031_,
    new_n6032_, new_n6033_, new_n6034_, new_n6035_, new_n6036_, new_n6037_,
    new_n6038_, new_n6039_, new_n6040_, new_n6041_, new_n6042_, new_n6043_,
    new_n6044_, new_n6045_, new_n6046_, new_n6047_, new_n6048_, new_n6049_,
    new_n6050_, new_n6051_, new_n6052_, new_n6053_, new_n6054_, new_n6055_,
    new_n6056_, new_n6057_, new_n6058_, new_n6059_, new_n6060_, new_n6061_,
    new_n6062_, new_n6063_, new_n6064_, new_n6065_, new_n6067_, new_n6068_,
    new_n6069_, new_n6070_, new_n6071_, new_n6072_, new_n6073_, new_n6074_,
    new_n6075_, new_n6076_, new_n6077_, new_n6078_, new_n6079_, new_n6080_,
    new_n6081_, new_n6082_, new_n6083_, new_n6084_, new_n6085_, new_n6086_,
    new_n6087_, new_n6088_, new_n6089_, new_n6090_, new_n6091_, new_n6092_,
    new_n6093_, new_n6094_, new_n6095_, new_n6096_, new_n6097_, new_n6098_,
    new_n6099_, new_n6100_, new_n6101_, new_n6102_, new_n6103_, new_n6104_,
    new_n6105_, new_n6106_, new_n6107_, new_n6108_, new_n6109_, new_n6110_,
    new_n6111_, new_n6112_, new_n6113_, new_n6114_, new_n6115_, new_n6116_,
    new_n6117_, new_n6118_, new_n6119_, new_n6120_, new_n6121_, new_n6122_,
    new_n6123_, new_n6124_, new_n6125_, new_n6126_, new_n6127_, new_n6128_,
    new_n6129_, new_n6130_, new_n6131_, new_n6132_, new_n6133_, new_n6134_,
    new_n6135_, new_n6136_, new_n6137_, new_n6138_, new_n6139_, new_n6140_,
    new_n6141_, new_n6142_, new_n6143_, new_n6144_, new_n6145_, new_n6146_,
    new_n6147_, new_n6148_, new_n6149_, new_n6150_, new_n6151_, new_n6152_,
    new_n6154_, new_n6155_, new_n6156_, new_n6157_, new_n6158_, new_n6159_,
    new_n6160_, new_n6161_, new_n6162_, new_n6163_, new_n6164_, new_n6165_,
    new_n6166_, new_n6167_, new_n6168_, new_n6169_, new_n6170_, new_n6171_,
    new_n6172_, new_n6173_, new_n6174_, new_n6175_, new_n6176_, new_n6177_,
    new_n6178_, new_n6179_, new_n6180_, new_n6181_, new_n6182_, new_n6183_,
    new_n6184_, new_n6185_, new_n6186_, new_n6187_, new_n6188_, new_n6189_,
    new_n6190_, new_n6191_, new_n6192_, new_n6193_, new_n6194_, new_n6195_,
    new_n6196_, new_n6197_, new_n6198_, new_n6199_, new_n6200_, new_n6201_,
    new_n6202_, new_n6203_, new_n6204_, new_n6205_, new_n6206_, new_n6207_,
    new_n6208_, new_n6209_, new_n6210_, new_n6211_, new_n6212_, new_n6213_,
    new_n6214_, new_n6215_, new_n6216_, new_n6217_, new_n6218_, new_n6219_,
    new_n6220_, new_n6221_, new_n6222_, new_n6223_, new_n6224_, new_n6225_,
    new_n6226_, new_n6227_, new_n6228_, new_n6229_, new_n6230_, new_n6231_,
    new_n6232_, new_n6233_, new_n6234_, new_n6235_, new_n6236_, new_n6237_,
    new_n6238_, new_n6239_, new_n6241_, new_n6242_, new_n6243_, new_n6244_,
    new_n6245_, new_n6246_, new_n6247_, new_n6248_, new_n6249_, new_n6250_,
    new_n6251_, new_n6252_, new_n6253_, new_n6254_, new_n6255_, new_n6256_,
    new_n6257_, new_n6258_, new_n6259_, new_n6260_, new_n6261_, new_n6262_,
    new_n6263_, new_n6264_, new_n6265_, new_n6266_, new_n6267_, new_n6268_,
    new_n6269_, new_n6270_, new_n6271_, new_n6272_, new_n6273_, new_n6274_,
    new_n6275_, new_n6276_, new_n6277_, new_n6278_, new_n6279_, new_n6280_,
    new_n6281_, new_n6282_, new_n6283_, new_n6284_, new_n6285_, new_n6286_,
    new_n6287_, new_n6288_, new_n6289_, new_n6290_, new_n6291_, new_n6292_,
    new_n6293_, new_n6294_, new_n6295_, new_n6296_, new_n6297_, new_n6298_,
    new_n6299_, new_n6300_, new_n6301_, new_n6302_, new_n6303_, new_n6304_,
    new_n6305_, new_n6306_, new_n6307_, new_n6308_, new_n6309_, new_n6310_,
    new_n6311_, new_n6312_, new_n6313_, new_n6314_, new_n6315_, new_n6316_,
    new_n6317_, new_n6318_, new_n6319_, new_n6320_, new_n6321_, new_n6322_,
    new_n6323_, new_n6324_, new_n6325_, new_n6326_, new_n6328_, new_n6329_,
    new_n6330_, new_n6331_, new_n6332_, new_n6333_, new_n6334_, new_n6335_,
    new_n6336_, new_n6337_, new_n6338_, new_n6339_, new_n6340_, new_n6341_,
    new_n6342_, new_n6343_, new_n6344_, new_n6345_, new_n6346_, new_n6347_,
    new_n6348_, new_n6349_, new_n6350_, new_n6351_, new_n6352_, new_n6353_,
    new_n6354_, new_n6355_, new_n6356_, new_n6357_, new_n6358_, new_n6359_,
    new_n6360_, new_n6361_, new_n6362_, new_n6363_, new_n6364_, new_n6365_,
    new_n6366_, new_n6367_, new_n6368_, new_n6369_, new_n6370_, new_n6371_,
    new_n6372_, new_n6373_, new_n6374_, new_n6375_, new_n6376_, new_n6377_,
    new_n6378_, new_n6379_, new_n6380_, new_n6381_, new_n6382_, new_n6383_,
    new_n6384_, new_n6385_, new_n6386_, new_n6387_, new_n6388_, new_n6389_,
    new_n6390_, new_n6391_, new_n6392_, new_n6393_, new_n6394_, new_n6395_,
    new_n6396_, new_n6397_, new_n6398_, new_n6399_, new_n6400_, new_n6401_,
    new_n6402_, new_n6403_, new_n6404_, new_n6405_, new_n6406_, new_n6407_,
    new_n6408_, new_n6409_, new_n6410_, new_n6411_, new_n6412_, new_n6413_,
    new_n6415_, new_n6416_, new_n6417_, new_n6418_, new_n6419_, new_n6420_,
    new_n6421_, new_n6422_, new_n6423_, new_n6424_, new_n6425_, new_n6426_,
    new_n6427_, new_n6428_, new_n6429_, new_n6430_, new_n6431_, new_n6432_,
    new_n6433_, new_n6434_, new_n6435_, new_n6436_, new_n6437_, new_n6438_,
    new_n6439_, new_n6440_, new_n6441_, new_n6442_, new_n6443_, new_n6444_,
    new_n6445_, new_n6446_, new_n6447_, new_n6448_, new_n6449_, new_n6450_,
    new_n6451_, new_n6452_, new_n6453_, new_n6454_, new_n6455_, new_n6456_,
    new_n6457_, new_n6458_, new_n6459_, new_n6460_, new_n6461_, new_n6462_,
    new_n6463_, new_n6464_, new_n6465_, new_n6466_, new_n6467_, new_n6468_,
    new_n6469_, new_n6470_, new_n6471_, new_n6472_, new_n6473_, new_n6474_,
    new_n6475_, new_n6476_, new_n6477_, new_n6478_, new_n6479_, new_n6480_,
    new_n6481_, new_n6482_, new_n6483_, new_n6484_, new_n6485_, new_n6486_,
    new_n6487_, new_n6488_, new_n6489_, new_n6490_, new_n6491_, new_n6492_,
    new_n6493_, new_n6494_, new_n6495_, new_n6496_, new_n6497_, new_n6498_,
    new_n6499_, new_n6500_, new_n6502_, new_n6503_, new_n6504_, new_n6505_,
    new_n6506_, new_n6507_, new_n6508_, new_n6509_, new_n6510_, new_n6511_,
    new_n6512_, new_n6513_, new_n6514_, new_n6515_, new_n6516_, new_n6517_,
    new_n6518_, new_n6519_, new_n6520_, new_n6521_, new_n6522_, new_n6523_,
    new_n6524_, new_n6525_, new_n6526_, new_n6527_, new_n6528_, new_n6529_,
    new_n6530_, new_n6531_, new_n6532_, new_n6533_, new_n6534_, new_n6535_,
    new_n6536_, new_n6537_, new_n6538_, new_n6539_, new_n6540_, new_n6541_,
    new_n6542_, new_n6543_, new_n6544_, new_n6545_, new_n6546_, new_n6547_,
    new_n6548_, new_n6549_, new_n6550_, new_n6551_, new_n6552_, new_n6553_,
    new_n6554_, new_n6555_, new_n6556_, new_n6557_, new_n6558_, new_n6559_,
    new_n6560_, new_n6561_, new_n6562_, new_n6563_, new_n6564_, new_n6565_,
    new_n6566_, new_n6567_, new_n6568_, new_n6569_, new_n6570_, new_n6571_,
    new_n6572_, new_n6573_, new_n6574_, new_n6575_, new_n6576_, new_n6577_,
    new_n6578_, new_n6579_, new_n6580_, new_n6581_, new_n6582_, new_n6583_,
    new_n6584_, new_n6585_, new_n6586_, new_n6587_, new_n6589_, new_n6590_,
    new_n6591_, new_n6592_, new_n6593_, new_n6594_, new_n6595_, new_n6596_,
    new_n6597_, new_n6598_, new_n6599_, new_n6600_, new_n6601_, new_n6602_,
    new_n6603_, new_n6604_, new_n6605_, new_n6606_, new_n6607_, new_n6608_,
    new_n6609_, new_n6610_, new_n6611_, new_n6612_, new_n6613_, new_n6614_,
    new_n6615_, new_n6616_, new_n6617_, new_n6618_, new_n6619_, new_n6620_,
    new_n6621_, new_n6622_, new_n6623_, new_n6624_, new_n6625_, new_n6626_,
    new_n6627_, new_n6628_, new_n6629_, new_n6630_, new_n6631_, new_n6632_,
    new_n6633_, new_n6634_, new_n6635_, new_n6636_, new_n6637_, new_n6638_,
    new_n6639_, new_n6640_, new_n6641_, new_n6642_, new_n6643_, new_n6644_,
    new_n6645_, new_n6646_, new_n6647_, new_n6648_, new_n6649_, new_n6650_,
    new_n6651_, new_n6652_, new_n6653_, new_n6654_, new_n6655_, new_n6656_,
    new_n6657_, new_n6658_, new_n6659_, new_n6660_, new_n6661_, new_n6662_,
    new_n6663_, new_n6664_, new_n6665_, new_n6666_, new_n6667_, new_n6668_,
    new_n6669_, new_n6670_, new_n6671_, new_n6672_, new_n6673_, new_n6674_,
    new_n6676_, new_n6677_, new_n6678_, new_n6679_, new_n6680_, new_n6681_,
    new_n6682_, new_n6683_, new_n6684_, new_n6685_, new_n6686_, new_n6687_,
    new_n6688_, new_n6689_, new_n6690_, new_n6691_, new_n6692_, new_n6693_,
    new_n6694_, new_n6695_, new_n6696_, new_n6697_, new_n6698_, new_n6699_,
    new_n6700_, new_n6701_, new_n6702_, new_n6703_, new_n6704_, new_n6705_,
    new_n6706_, new_n6707_, new_n6708_, new_n6709_, new_n6710_, new_n6711_,
    new_n6712_, new_n6713_, new_n6714_, new_n6715_, new_n6716_, new_n6717_,
    new_n6718_, new_n6719_, new_n6720_, new_n6721_, new_n6722_, new_n6723_,
    new_n6724_, new_n6725_, new_n6726_, new_n6727_, new_n6728_, new_n6729_,
    new_n6730_, new_n6731_, new_n6732_, new_n6733_, new_n6734_, new_n6735_,
    new_n6736_, new_n6737_, new_n6738_, new_n6739_, new_n6740_, new_n6741_,
    new_n6742_, new_n6743_, new_n6744_, new_n6745_, new_n6746_, new_n6747_,
    new_n6748_, new_n6749_, new_n6750_, new_n6751_, new_n6752_, new_n6753_,
    new_n6754_, new_n6755_, new_n6756_, new_n6757_, new_n6758_, new_n6759_,
    new_n6760_, new_n6761_, new_n6763_, new_n6764_, new_n6765_, new_n6766_,
    new_n6767_, new_n6768_, new_n6769_, new_n6770_, new_n6771_, new_n6772_,
    new_n6773_, new_n6774_, new_n6775_, new_n6776_, new_n6777_, new_n6778_,
    new_n6779_, new_n6780_, new_n6781_, new_n6782_, new_n6783_, new_n6784_,
    new_n6785_, new_n6786_, new_n6787_, new_n6788_, new_n6789_, new_n6790_,
    new_n6791_, new_n6792_, new_n6793_, new_n6794_, new_n6795_, new_n6796_,
    new_n6797_, new_n6798_, new_n6799_, new_n6800_, new_n6801_, new_n6802_,
    new_n6803_, new_n6804_, new_n6805_, new_n6806_, new_n6807_, new_n6808_,
    new_n6809_, new_n6810_, new_n6811_, new_n6812_, new_n6813_, new_n6814_,
    new_n6815_, new_n6816_, new_n6817_, new_n6818_, new_n6819_, new_n6820_,
    new_n6821_, new_n6822_, new_n6823_, new_n6824_, new_n6825_, new_n6826_,
    new_n6827_, new_n6828_, new_n6829_, new_n6830_, new_n6831_, new_n6832_,
    new_n6833_, new_n6834_, new_n6835_, new_n6836_, new_n6837_, new_n6838_,
    new_n6839_, new_n6840_, new_n6841_, new_n6842_, new_n6843_, new_n6844_,
    new_n6845_, new_n6846_, new_n6847_, new_n6848_, new_n6850_, new_n6851_,
    new_n6852_, new_n6853_, new_n6854_, new_n6855_, new_n6856_, new_n6857_,
    new_n6858_, new_n6859_, new_n6860_, new_n6861_, new_n6862_, new_n6863_,
    new_n6864_, new_n6865_, new_n6866_, new_n6867_, new_n6868_, new_n6869_,
    new_n6870_, new_n6871_, new_n6872_, new_n6873_, new_n6874_, new_n6875_,
    new_n6876_, new_n6877_, new_n6878_, new_n6879_, new_n6880_, new_n6881_,
    new_n6882_, new_n6883_, new_n6884_, new_n6885_, new_n6886_, new_n6887_,
    new_n6888_, new_n6889_, new_n6890_, new_n6891_, new_n6892_, new_n6893_,
    new_n6894_, new_n6895_, new_n6896_, new_n6897_, new_n6898_, new_n6899_,
    new_n6900_, new_n6901_, new_n6902_, new_n6903_, new_n6904_, new_n6905_,
    new_n6906_, new_n6907_, new_n6908_, new_n6909_, new_n6910_, new_n6911_,
    new_n6912_, new_n6913_, new_n6914_, new_n6915_, new_n6916_, new_n6917_,
    new_n6918_, new_n6919_, new_n6920_, new_n6921_, new_n6922_, new_n6923_,
    new_n6924_, new_n6925_, new_n6926_, new_n6927_, new_n6928_, new_n6929_,
    new_n6930_, new_n6931_, new_n6932_, new_n6933_, new_n6934_, new_n6935_,
    new_n6937_, new_n6938_, new_n6939_, new_n6940_, new_n6941_, new_n6942_,
    new_n6943_, new_n6944_, new_n6945_, new_n6946_, new_n6947_, new_n6948_,
    new_n6949_, new_n6950_, new_n6951_, new_n6952_, new_n6953_, new_n6954_,
    new_n6955_, new_n6956_, new_n6957_, new_n6958_, new_n6959_, new_n6960_,
    new_n6961_, new_n6962_, new_n6963_, new_n6964_, new_n6965_, new_n6966_,
    new_n6967_, new_n6968_, new_n6969_, new_n6970_, new_n6971_, new_n6972_,
    new_n6973_, new_n6974_, new_n6975_, new_n6976_, new_n6977_, new_n6978_,
    new_n6979_, new_n6980_, new_n6981_, new_n6982_, new_n6983_, new_n6984_,
    new_n6985_, new_n6986_, new_n6987_, new_n6988_, new_n6989_, new_n6990_,
    new_n6991_, new_n6992_, new_n6993_, new_n6994_, new_n6995_, new_n6996_,
    new_n6997_, new_n6998_, new_n6999_, new_n7000_, new_n7001_, new_n7002_,
    new_n7003_, new_n7004_, new_n7005_, new_n7006_, new_n7007_, new_n7008_,
    new_n7009_, new_n7010_, new_n7011_, new_n7012_, new_n7013_, new_n7014_,
    new_n7015_, new_n7016_, new_n7017_, new_n7018_, new_n7019_, new_n7020_,
    new_n7021_, new_n7022_, new_n7024_, new_n7025_, new_n7026_, new_n7027_,
    new_n7028_, new_n7029_, new_n7030_, new_n7031_, new_n7032_, new_n7033_,
    new_n7034_, new_n7035_, new_n7036_, new_n7037_, new_n7038_, new_n7039_,
    new_n7040_, new_n7041_, new_n7042_, new_n7043_, new_n7044_, new_n7045_,
    new_n7046_, new_n7047_, new_n7048_, new_n7049_, new_n7050_, new_n7051_,
    new_n7052_, new_n7053_, new_n7054_, new_n7055_, new_n7056_, new_n7057_,
    new_n7058_, new_n7059_, new_n7060_, new_n7061_, new_n7062_, new_n7063_,
    new_n7064_, new_n7065_, new_n7066_, new_n7067_, new_n7068_, new_n7069_,
    new_n7070_, new_n7071_, new_n7072_, new_n7073_, new_n7074_, new_n7075_,
    new_n7076_, new_n7077_, new_n7078_, new_n7079_, new_n7080_, new_n7081_,
    new_n7082_, new_n7083_, new_n7084_, new_n7085_, new_n7086_, new_n7087_,
    new_n7088_, new_n7089_, new_n7090_, new_n7091_, new_n7092_, new_n7093_,
    new_n7094_, new_n7095_, new_n7096_, new_n7097_, new_n7098_, new_n7099_,
    new_n7100_, new_n7101_, new_n7102_, new_n7103_, new_n7104_, new_n7105_,
    new_n7106_, new_n7107_, new_n7108_, new_n7109_, new_n7111_, new_n7112_,
    new_n7113_, new_n7114_, new_n7115_, new_n7116_, new_n7117_, new_n7118_,
    new_n7119_, new_n7120_, new_n7121_, new_n7122_, new_n7123_, new_n7124_,
    new_n7125_, new_n7126_, new_n7127_, new_n7128_, new_n7129_, new_n7130_,
    new_n7131_, new_n7132_, new_n7133_, new_n7134_, new_n7135_, new_n7136_,
    new_n7137_, new_n7138_, new_n7139_, new_n7140_, new_n7141_, new_n7142_,
    new_n7143_, new_n7144_, new_n7145_, new_n7146_, new_n7147_, new_n7148_,
    new_n7149_, new_n7150_, new_n7151_, new_n7152_, new_n7153_, new_n7154_,
    new_n7155_, new_n7156_, new_n7157_, new_n7158_, new_n7159_, new_n7160_,
    new_n7161_, new_n7162_, new_n7163_, new_n7164_, new_n7165_, new_n7166_,
    new_n7167_, new_n7168_, new_n7169_, new_n7170_, new_n7171_, new_n7172_,
    new_n7173_, new_n7174_, new_n7175_, new_n7176_, new_n7177_, new_n7178_,
    new_n7179_, new_n7180_, new_n7181_, new_n7182_, new_n7183_, new_n7184_,
    new_n7185_, new_n7186_, new_n7187_, new_n7188_, new_n7189_, new_n7190_,
    new_n7191_, new_n7192_, new_n7193_, new_n7194_, new_n7195_, new_n7196_,
    new_n7198_, new_n7199_, new_n7200_, new_n7201_, new_n7202_, new_n7203_,
    new_n7204_, new_n7205_, new_n7206_, new_n7207_, new_n7208_, new_n7209_,
    new_n7210_, new_n7211_, new_n7212_, new_n7213_, new_n7214_, new_n7215_,
    new_n7216_, new_n7217_, new_n7218_, new_n7219_, new_n7220_, new_n7221_,
    new_n7222_, new_n7223_, new_n7224_, new_n7225_, new_n7226_, new_n7227_,
    new_n7228_, new_n7229_, new_n7230_, new_n7231_, new_n7232_, new_n7233_,
    new_n7234_, new_n7235_, new_n7236_, new_n7237_, new_n7238_, new_n7239_,
    new_n7240_, new_n7241_, new_n7242_, new_n7243_, new_n7244_, new_n7245_,
    new_n7246_, new_n7247_, new_n7248_, new_n7249_, new_n7250_, new_n7251_,
    new_n7252_, new_n7253_, new_n7254_, new_n7255_, new_n7256_, new_n7257_,
    new_n7258_, new_n7259_, new_n7260_, new_n7261_, new_n7262_, new_n7263_,
    new_n7264_, new_n7265_, new_n7266_, new_n7267_, new_n7268_, new_n7269_,
    new_n7270_, new_n7271_, new_n7272_, new_n7273_, new_n7274_, new_n7275_,
    new_n7276_, new_n7277_, new_n7278_, new_n7279_, new_n7280_, new_n7281_,
    new_n7282_, new_n7283_, new_n7285_, new_n7286_, new_n7287_, new_n7288_,
    new_n7289_, new_n7290_, new_n7291_, new_n7292_, new_n7293_, new_n7294_,
    new_n7295_, new_n7296_, new_n7297_, new_n7298_, new_n7299_, new_n7300_,
    new_n7301_, new_n7302_, new_n7303_, new_n7304_, new_n7305_, new_n7306_,
    new_n7307_, new_n7308_, new_n7309_, new_n7310_, new_n7311_, new_n7312_,
    new_n7313_, new_n7314_, new_n7315_, new_n7316_, new_n7317_, new_n7318_,
    new_n7319_, new_n7320_, new_n7321_, new_n7322_, new_n7323_, new_n7324_,
    new_n7325_, new_n7326_, new_n7327_, new_n7328_, new_n7329_, new_n7330_,
    new_n7331_, new_n7332_, new_n7333_, new_n7334_, new_n7335_, new_n7336_,
    new_n7337_, new_n7338_, new_n7339_, new_n7340_, new_n7341_, new_n7342_,
    new_n7343_, new_n7344_, new_n7345_, new_n7346_, new_n7347_, new_n7348_,
    new_n7349_, new_n7350_, new_n7351_, new_n7352_, new_n7353_, new_n7354_,
    new_n7355_, new_n7356_, new_n7357_, new_n7358_, new_n7359_, new_n7360_,
    new_n7361_, new_n7362_, new_n7363_, new_n7364_, new_n7365_, new_n7366_,
    new_n7367_, new_n7368_, new_n7369_, new_n7370_, new_n7372_, new_n7373_,
    new_n7374_, new_n7375_, new_n7376_, new_n7377_, new_n7378_, new_n7379_,
    new_n7380_, new_n7381_, new_n7382_, new_n7383_, new_n7384_, new_n7385_,
    new_n7386_, new_n7387_, new_n7388_, new_n7389_, new_n7390_, new_n7391_,
    new_n7392_, new_n7393_, new_n7394_, new_n7395_, new_n7396_, new_n7397_,
    new_n7398_, new_n7399_, new_n7400_, new_n7401_, new_n7402_, new_n7403_,
    new_n7404_, new_n7405_, new_n7406_, new_n7407_, new_n7408_, new_n7409_,
    new_n7410_, new_n7411_, new_n7412_, new_n7413_, new_n7414_, new_n7415_,
    new_n7416_, new_n7417_, new_n7418_, new_n7419_, new_n7420_, new_n7421_,
    new_n7422_, new_n7423_, new_n7424_, new_n7425_, new_n7426_, new_n7427_,
    new_n7428_, new_n7429_, new_n7430_, new_n7431_, new_n7432_, new_n7433_,
    new_n7434_, new_n7435_, new_n7436_, new_n7437_, new_n7438_, new_n7439_,
    new_n7440_, new_n7441_, new_n7442_, new_n7443_, new_n7444_, new_n7445_,
    new_n7446_, new_n7447_, new_n7448_, new_n7449_, new_n7450_, new_n7451_,
    new_n7452_, new_n7453_, new_n7454_, new_n7455_, new_n7456_, new_n7457_,
    new_n7459_, new_n7460_, new_n7461_, new_n7462_, new_n7463_, new_n7464_,
    new_n7465_, new_n7466_, new_n7467_, new_n7468_, new_n7469_, new_n7470_,
    new_n7471_, new_n7472_, new_n7473_, new_n7474_, new_n7475_, new_n7476_,
    new_n7477_, new_n7478_, new_n7479_, new_n7480_, new_n7481_, new_n7482_,
    new_n7483_, new_n7484_, new_n7485_, new_n7486_, new_n7487_, new_n7488_,
    new_n7489_, new_n7490_, new_n7491_, new_n7492_, new_n7493_, new_n7494_,
    new_n7495_, new_n7496_, new_n7497_, new_n7498_, new_n7499_, new_n7500_,
    new_n7501_, new_n7502_, new_n7503_, new_n7504_, new_n7505_, new_n7506_,
    new_n7507_, new_n7508_, new_n7509_, new_n7510_, new_n7511_, new_n7512_,
    new_n7513_, new_n7514_, new_n7515_, new_n7516_, new_n7517_, new_n7518_,
    new_n7519_, new_n7520_, new_n7521_, new_n7522_, new_n7523_, new_n7524_,
    new_n7525_, new_n7526_, new_n7527_, new_n7528_, new_n7529_, new_n7530_,
    new_n7531_, new_n7532_, new_n7533_, new_n7534_, new_n7535_, new_n7536_,
    new_n7537_, new_n7538_, new_n7539_, new_n7540_, new_n7541_, new_n7542_,
    new_n7543_, new_n7544_, new_n7546_, new_n7547_, new_n7548_, new_n7549_,
    new_n7550_, new_n7551_, new_n7552_, new_n7553_, new_n7554_, new_n7555_,
    new_n7556_, new_n7557_, new_n7558_, new_n7559_, new_n7560_, new_n7561_,
    new_n7562_, new_n7563_, new_n7564_, new_n7565_, new_n7566_, new_n7567_,
    new_n7568_, new_n7569_, new_n7570_, new_n7571_, new_n7572_, new_n7573_,
    new_n7574_, new_n7575_, new_n7576_, new_n7577_, new_n7578_, new_n7579_,
    new_n7580_, new_n7581_, new_n7582_, new_n7583_, new_n7584_, new_n7585_,
    new_n7586_, new_n7587_, new_n7588_, new_n7589_, new_n7590_, new_n7591_,
    new_n7592_, new_n7593_, new_n7594_, new_n7595_, new_n7596_, new_n7597_,
    new_n7598_, new_n7599_, new_n7600_, new_n7601_, new_n7602_, new_n7603_,
    new_n7604_, new_n7605_, new_n7606_, new_n7607_, new_n7608_, new_n7609_,
    new_n7610_, new_n7611_, new_n7612_, new_n7613_, new_n7614_, new_n7615_,
    new_n7616_, new_n7617_, new_n7618_, new_n7619_, new_n7620_, new_n7621_,
    new_n7622_, new_n7623_, new_n7624_, new_n7625_, new_n7626_, new_n7627_,
    new_n7628_, new_n7629_, new_n7630_, new_n7631_, new_n7633_, new_n7634_,
    new_n7635_, new_n7636_, new_n7637_, new_n7638_, new_n7639_, new_n7640_,
    new_n7641_, new_n7642_, new_n7643_, new_n7644_, new_n7645_, new_n7646_,
    new_n7647_, new_n7648_, new_n7649_, new_n7650_, new_n7651_, new_n7652_,
    new_n7653_, new_n7654_, new_n7655_, new_n7656_, new_n7657_, new_n7658_,
    new_n7659_, new_n7660_, new_n7661_, new_n7662_, new_n7663_, new_n7664_,
    new_n7665_, new_n7666_, new_n7667_, new_n7668_, new_n7669_, new_n7670_,
    new_n7671_, new_n7672_, new_n7673_, new_n7674_, new_n7675_, new_n7676_,
    new_n7677_, new_n7678_, new_n7679_, new_n7680_, new_n7681_, new_n7682_,
    new_n7683_, new_n7684_, new_n7685_, new_n7686_, new_n7687_, new_n7688_,
    new_n7689_, new_n7690_, new_n7691_, new_n7692_, new_n7693_, new_n7694_,
    new_n7695_, new_n7696_, new_n7697_, new_n7698_, new_n7699_, new_n7700_,
    new_n7701_, new_n7702_, new_n7703_, new_n7704_, new_n7705_, new_n7706_,
    new_n7707_, new_n7708_, new_n7709_, new_n7710_, new_n7711_, new_n7712_,
    new_n7713_, new_n7714_, new_n7715_, new_n7716_, new_n7717_, new_n7718_,
    new_n7720_, new_n7721_, new_n7722_, new_n7723_, new_n7724_, new_n7725_,
    new_n7726_, new_n7727_, new_n7728_, new_n7729_, new_n7730_, new_n7731_,
    new_n7732_, new_n7733_, new_n7734_, new_n7735_, new_n7736_, new_n7737_,
    new_n7738_, new_n7739_, new_n7740_, new_n7741_, new_n7742_, new_n7743_,
    new_n7744_, new_n7745_, new_n7746_, new_n7747_, new_n7748_, new_n7749_,
    new_n7750_, new_n7751_, new_n7752_, new_n7753_, new_n7754_, new_n7755_,
    new_n7756_, new_n7757_, new_n7758_, new_n7759_, new_n7760_, new_n7761_,
    new_n7762_, new_n7763_, new_n7764_, new_n7765_, new_n7766_, new_n7767_,
    new_n7768_, new_n7769_, new_n7770_, new_n7771_, new_n7772_, new_n7773_,
    new_n7774_, new_n7775_, new_n7776_, new_n7777_, new_n7778_, new_n7779_,
    new_n7780_, new_n7781_, new_n7782_, new_n7783_, new_n7784_, new_n7785_,
    new_n7786_, new_n7787_, new_n7788_, new_n7789_, new_n7790_, new_n7791_,
    new_n7792_, new_n7793_, new_n7794_, new_n7795_, new_n7796_, new_n7797_,
    new_n7798_, new_n7799_, new_n7800_, new_n7801_, new_n7802_, new_n7803_,
    new_n7804_, new_n7805_, new_n7807_, new_n7808_, new_n7809_, new_n7810_,
    new_n7811_, new_n7812_, new_n7813_, new_n7814_, new_n7815_, new_n7816_,
    new_n7817_, new_n7818_, new_n7819_, new_n7820_, new_n7821_, new_n7822_,
    new_n7823_, new_n7824_, new_n7825_, new_n7826_, new_n7827_, new_n7828_,
    new_n7829_, new_n7830_, new_n7831_, new_n7832_, new_n7833_, new_n7834_,
    new_n7835_, new_n7836_, new_n7837_, new_n7838_, new_n7839_, new_n7840_,
    new_n7841_, new_n7842_, new_n7843_, new_n7844_, new_n7845_, new_n7846_,
    new_n7847_, new_n7848_, new_n7849_, new_n7850_, new_n7851_, new_n7852_,
    new_n7853_, new_n7854_, new_n7855_, new_n7856_, new_n7857_, new_n7858_,
    new_n7859_, new_n7860_, new_n7861_, new_n7862_, new_n7863_, new_n7864_,
    new_n7865_, new_n7866_, new_n7867_, new_n7868_, new_n7869_, new_n7870_,
    new_n7871_, new_n7872_, new_n7873_, new_n7874_, new_n7875_, new_n7876_,
    new_n7877_, new_n7878_, new_n7879_, new_n7880_, new_n7881_, new_n7882_,
    new_n7883_, new_n7884_, new_n7885_, new_n7886_, new_n7887_, new_n7888_,
    new_n7889_, new_n7890_, new_n7891_, new_n7892_, new_n7894_, new_n7895_,
    new_n7896_, new_n7897_, new_n7898_, new_n7899_, new_n7900_, new_n7901_,
    new_n7902_, new_n7903_, new_n7904_, new_n7905_, new_n7906_, new_n7907_,
    new_n7908_, new_n7909_, new_n7910_, new_n7911_, new_n7912_, new_n7913_,
    new_n7914_, new_n7915_, new_n7916_, new_n7917_, new_n7918_, new_n7919_,
    new_n7920_, new_n7921_, new_n7922_, new_n7923_, new_n7924_, new_n7925_,
    new_n7926_, new_n7927_, new_n7928_, new_n7929_, new_n7930_, new_n7931_,
    new_n7932_, new_n7933_, new_n7934_, new_n7935_, new_n7936_, new_n7937_,
    new_n7938_, new_n7939_, new_n7940_, new_n7941_, new_n7942_, new_n7943_,
    new_n7944_, new_n7945_, new_n7946_, new_n7947_, new_n7948_, new_n7949_,
    new_n7950_, new_n7951_, new_n7952_, new_n7953_, new_n7954_, new_n7955_,
    new_n7956_, new_n7957_, new_n7958_, new_n7959_, new_n7960_, new_n7961_,
    new_n7962_, new_n7963_, new_n7964_, new_n7965_, new_n7966_, new_n7967_,
    new_n7968_, new_n7969_, new_n7970_, new_n7971_, new_n7972_, new_n7973_,
    new_n7974_, new_n7975_, new_n7976_, new_n7977_, new_n7978_, new_n7979_,
    new_n7981_, new_n7982_, new_n7983_, new_n7984_, new_n7985_, new_n7986_,
    new_n7987_, new_n7988_, new_n7989_, new_n7990_, new_n7991_, new_n7992_,
    new_n7993_, new_n7994_, new_n7995_, new_n7996_, new_n7997_, new_n7998_,
    new_n7999_, new_n8000_, new_n8001_, new_n8002_, new_n8003_, new_n8004_,
    new_n8005_, new_n8006_, new_n8007_, new_n8008_, new_n8009_, new_n8010_,
    new_n8011_, new_n8012_, new_n8013_, new_n8014_, new_n8015_, new_n8016_,
    new_n8017_, new_n8018_, new_n8019_, new_n8020_, new_n8021_, new_n8022_,
    new_n8023_, new_n8024_, new_n8025_, new_n8026_, new_n8027_, new_n8028_,
    new_n8029_, new_n8030_, new_n8031_, new_n8032_, new_n8033_, new_n8034_,
    new_n8035_, new_n8036_, new_n8037_, new_n8038_, new_n8039_, new_n8040_,
    new_n8041_, new_n8042_, new_n8043_, new_n8044_, new_n8045_, new_n8046_,
    new_n8047_, new_n8048_, new_n8049_, new_n8050_, new_n8051_, new_n8052_,
    new_n8053_, new_n8054_, new_n8055_, new_n8056_, new_n8057_, new_n8058_,
    new_n8059_, new_n8060_, new_n8061_, new_n8062_, new_n8063_, new_n8064_,
    new_n8065_, new_n8066_, new_n8068_, new_n8069_, new_n8070_, new_n8071_,
    new_n8072_, new_n8073_, new_n8074_, new_n8075_, new_n8076_, new_n8077_,
    new_n8078_, new_n8079_, new_n8080_, new_n8081_, new_n8082_, new_n8083_,
    new_n8084_, new_n8085_, new_n8086_, new_n8087_, new_n8088_, new_n8089_,
    new_n8090_, new_n8091_, new_n8092_, new_n8093_, new_n8094_, new_n8095_,
    new_n8096_, new_n8097_, new_n8098_, new_n8099_, new_n8100_, new_n8101_,
    new_n8102_, new_n8103_, new_n8104_, new_n8105_, new_n8106_, new_n8107_,
    new_n8108_, new_n8109_, new_n8110_, new_n8111_, new_n8112_, new_n8113_,
    new_n8114_, new_n8115_, new_n8116_, new_n8117_, new_n8118_, new_n8119_,
    new_n8120_, new_n8121_, new_n8122_, new_n8123_, new_n8124_, new_n8125_,
    new_n8126_, new_n8127_, new_n8128_, new_n8129_, new_n8130_, new_n8131_,
    new_n8132_, new_n8133_, new_n8134_, new_n8135_, new_n8136_, new_n8137_,
    new_n8138_, new_n8139_, new_n8140_, new_n8141_, new_n8142_, new_n8143_,
    new_n8144_, new_n8145_, new_n8146_, new_n8147_, new_n8148_, new_n8149_,
    new_n8150_, new_n8151_, new_n8152_, new_n8153_, new_n8155_, new_n8156_,
    new_n8157_, new_n8158_, new_n8159_, new_n8160_, new_n8161_, new_n8162_,
    new_n8163_, new_n8164_, new_n8165_, new_n8166_, new_n8167_, new_n8168_,
    new_n8169_, new_n8170_, new_n8171_, new_n8172_, new_n8173_, new_n8174_,
    new_n8175_, new_n8176_, new_n8177_, new_n8178_, new_n8179_, new_n8180_,
    new_n8181_, new_n8182_, new_n8183_, new_n8184_, new_n8185_, new_n8186_,
    new_n8187_, new_n8188_, new_n8189_, new_n8190_, new_n8191_, new_n8192_,
    new_n8193_, new_n8194_, new_n8195_, new_n8196_, new_n8197_, new_n8198_,
    new_n8199_, new_n8200_, new_n8201_, new_n8202_, new_n8203_, new_n8204_,
    new_n8205_, new_n8206_, new_n8207_, new_n8208_, new_n8209_, new_n8210_,
    new_n8211_, new_n8212_, new_n8213_, new_n8214_, new_n8215_, new_n8216_,
    new_n8217_, new_n8218_, new_n8219_, new_n8220_, new_n8221_, new_n8222_,
    new_n8223_, new_n8224_, new_n8225_, new_n8226_, new_n8227_, new_n8228_,
    new_n8229_, new_n8230_, new_n8231_, new_n8232_, new_n8233_, new_n8234_,
    new_n8235_, new_n8236_, new_n8237_, new_n8238_, new_n8239_, new_n8240_,
    new_n8242_, new_n8243_, new_n8244_, new_n8245_, new_n8246_, new_n8247_,
    new_n8248_, new_n8249_, new_n8250_, new_n8251_, new_n8252_, new_n8253_,
    new_n8254_, new_n8255_, new_n8256_, new_n8257_, new_n8258_, new_n8259_,
    new_n8260_, new_n8261_, new_n8262_, new_n8263_, new_n8264_, new_n8265_,
    new_n8266_, new_n8267_, new_n8268_, new_n8269_, new_n8270_, new_n8271_,
    new_n8272_, new_n8273_, new_n8274_, new_n8275_, new_n8276_, new_n8277_,
    new_n8278_, new_n8279_, new_n8280_, new_n8281_, new_n8282_, new_n8283_,
    new_n8284_, new_n8285_, new_n8286_, new_n8287_, new_n8288_, new_n8289_,
    new_n8290_, new_n8291_, new_n8292_, new_n8293_, new_n8294_, new_n8295_,
    new_n8296_, new_n8297_, new_n8298_, new_n8299_, new_n8300_, new_n8301_,
    new_n8302_, new_n8303_, new_n8304_, new_n8305_, new_n8306_, new_n8307_,
    new_n8308_, new_n8309_, new_n8310_, new_n8311_, new_n8312_, new_n8313_,
    new_n8314_, new_n8315_, new_n8316_, new_n8317_, new_n8318_, new_n8319_,
    new_n8320_, new_n8321_, new_n8322_, new_n8323_, new_n8324_, new_n8325_,
    new_n8326_, new_n8327_, new_n8329_, new_n8330_, new_n8331_, new_n8332_,
    new_n8333_, new_n8334_, new_n8335_, new_n8336_, new_n8337_, new_n8338_,
    new_n8339_, new_n8340_, new_n8341_, new_n8342_, new_n8343_, new_n8344_,
    new_n8345_, new_n8346_, new_n8347_, new_n8348_, new_n8349_, new_n8350_,
    new_n8351_, new_n8352_, new_n8353_, new_n8354_, new_n8355_, new_n8356_,
    new_n8357_, new_n8358_, new_n8359_, new_n8360_, new_n8361_, new_n8362_,
    new_n8363_, new_n8364_, new_n8365_, new_n8366_, new_n8367_, new_n8368_,
    new_n8369_, new_n8370_, new_n8371_, new_n8372_, new_n8373_, new_n8374_,
    new_n8375_, new_n8376_, new_n8377_, new_n8378_, new_n8379_, new_n8380_,
    new_n8381_, new_n8382_, new_n8383_, new_n8384_, new_n8385_, new_n8386_,
    new_n8387_, new_n8388_, new_n8389_, new_n8390_, new_n8391_, new_n8392_,
    new_n8393_, new_n8394_, new_n8395_, new_n8396_, new_n8397_, new_n8398_,
    new_n8399_, new_n8400_, new_n8401_, new_n8402_, new_n8403_, new_n8404_,
    new_n8405_, new_n8406_, new_n8407_, new_n8408_, new_n8409_, new_n8410_,
    new_n8411_, new_n8412_, new_n8413_, new_n8414_, new_n8416_, new_n8417_,
    new_n8418_, new_n8419_, new_n8420_, new_n8421_, new_n8422_, new_n8423_,
    new_n8424_, new_n8425_, new_n8426_, new_n8427_, new_n8428_, new_n8429_,
    new_n8430_, new_n8431_, new_n8432_, new_n8433_, new_n8434_, new_n8435_,
    new_n8436_, new_n8437_, new_n8438_, new_n8439_, new_n8440_, new_n8441_,
    new_n8442_, new_n8443_, new_n8444_, new_n8445_, new_n8446_, new_n8447_,
    new_n8448_, new_n8449_, new_n8450_, new_n8451_, new_n8452_, new_n8453_,
    new_n8454_, new_n8455_, new_n8456_, new_n8457_, new_n8458_, new_n8459_,
    new_n8460_, new_n8461_, new_n8462_, new_n8463_, new_n8464_, new_n8465_,
    new_n8466_, new_n8467_, new_n8468_, new_n8469_, new_n8470_, new_n8471_,
    new_n8472_, new_n8473_, new_n8474_, new_n8475_, new_n8476_, new_n8477_,
    new_n8478_, new_n8479_, new_n8480_, new_n8481_, new_n8482_, new_n8483_,
    new_n8484_, new_n8485_, new_n8486_, new_n8487_, new_n8488_, new_n8489_,
    new_n8490_, new_n8491_, new_n8492_, new_n8493_, new_n8494_, new_n8495_,
    new_n8496_, new_n8497_, new_n8498_, new_n8499_, new_n8500_, new_n8501_,
    new_n8503_, new_n8504_, new_n8505_, new_n8506_, new_n8507_, new_n8508_,
    new_n8509_, new_n8510_, new_n8511_, new_n8512_, new_n8513_, new_n8514_,
    new_n8515_, new_n8516_, new_n8517_, new_n8518_, new_n8519_, new_n8520_,
    new_n8521_, new_n8522_, new_n8523_, new_n8524_, new_n8525_, new_n8526_,
    new_n8527_, new_n8528_, new_n8529_, new_n8530_, new_n8531_, new_n8532_,
    new_n8533_, new_n8534_, new_n8535_, new_n8536_, new_n8537_, new_n8538_,
    new_n8539_, new_n8540_, new_n8541_, new_n8542_, new_n8543_, new_n8544_,
    new_n8545_, new_n8546_, new_n8547_, new_n8548_, new_n8549_, new_n8550_,
    new_n8551_, new_n8552_, new_n8553_, new_n8554_, new_n8555_, new_n8556_,
    new_n8557_, new_n8558_, new_n8559_, new_n8560_, new_n8561_, new_n8562_,
    new_n8563_, new_n8564_, new_n8565_, new_n8566_, new_n8567_, new_n8568_,
    new_n8569_, new_n8570_, new_n8571_, new_n8572_, new_n8573_, new_n8574_,
    new_n8575_, new_n8576_, new_n8577_, new_n8578_, new_n8579_, new_n8580_,
    new_n8581_, new_n8582_, new_n8583_, new_n8584_, new_n8585_, new_n8586_,
    new_n8587_, new_n8588_, new_n8590_, new_n8591_, new_n8592_, new_n8593_,
    new_n8594_, new_n8595_, new_n8596_, new_n8597_, new_n8598_, new_n8599_,
    new_n8600_, new_n8601_, new_n8602_, new_n8603_, new_n8604_, new_n8605_,
    new_n8606_, new_n8607_, new_n8608_, new_n8609_, new_n8610_, new_n8611_,
    new_n8612_, new_n8613_, new_n8614_, new_n8615_, new_n8616_, new_n8617_,
    new_n8618_, new_n8619_, new_n8620_, new_n8621_, new_n8622_, new_n8623_,
    new_n8624_, new_n8625_, new_n8626_, new_n8627_, new_n8628_, new_n8629_,
    new_n8630_, new_n8631_, new_n8632_, new_n8633_, new_n8634_, new_n8635_,
    new_n8636_, new_n8637_, new_n8638_, new_n8639_, new_n8640_, new_n8641_,
    new_n8642_, new_n8643_, new_n8644_, new_n8645_, new_n8646_, new_n8647_,
    new_n8648_, new_n8649_, new_n8650_, new_n8651_, new_n8652_, new_n8653_,
    new_n8654_, new_n8655_, new_n8656_, new_n8657_, new_n8658_, new_n8659_,
    new_n8660_, new_n8661_, new_n8662_, new_n8663_, new_n8664_, new_n8665_,
    new_n8666_, new_n8667_, new_n8668_, new_n8669_, new_n8670_, new_n8671_,
    new_n8672_, new_n8673_, new_n8674_, new_n8675_, new_n8677_, new_n8678_,
    new_n8679_, new_n8680_, new_n8681_, new_n8682_, new_n8683_, new_n8684_,
    new_n8685_, new_n8686_, new_n8687_, new_n8688_, new_n8689_, new_n8690_,
    new_n8691_, new_n8692_, new_n8693_, new_n8694_, new_n8695_, new_n8696_,
    new_n8697_, new_n8698_, new_n8699_, new_n8700_, new_n8701_, new_n8702_,
    new_n8703_, new_n8704_, new_n8705_, new_n8706_, new_n8707_, new_n8708_,
    new_n8709_, new_n8710_, new_n8711_, new_n8712_, new_n8713_, new_n8714_,
    new_n8715_, new_n8716_, new_n8717_, new_n8718_, new_n8719_, new_n8720_,
    new_n8721_, new_n8722_, new_n8723_, new_n8724_, new_n8725_, new_n8726_,
    new_n8727_, new_n8728_, new_n8729_, new_n8730_, new_n8731_, new_n8732_,
    new_n8733_, new_n8734_, new_n8735_, new_n8736_, new_n8737_, new_n8738_,
    new_n8739_, new_n8740_, new_n8741_, new_n8742_, new_n8743_, new_n8744_,
    new_n8745_, new_n8746_, new_n8747_, new_n8748_, new_n8749_, new_n8750_,
    new_n8751_, new_n8752_, new_n8753_, new_n8754_, new_n8755_, new_n8756_,
    new_n8757_, new_n8758_, new_n8759_, new_n8760_, new_n8761_, new_n8762_,
    new_n8764_, new_n8765_, new_n8766_, new_n8767_, new_n8768_, new_n8769_,
    new_n8770_, new_n8771_, new_n8772_, new_n8773_, new_n8774_, new_n8775_,
    new_n8776_, new_n8777_, new_n8778_, new_n8779_, new_n8780_, new_n8781_,
    new_n8782_, new_n8783_, new_n8784_, new_n8785_, new_n8786_, new_n8787_,
    new_n8788_, new_n8789_, new_n8790_, new_n8791_, new_n8792_, new_n8793_,
    new_n8794_, new_n8795_, new_n8796_, new_n8797_, new_n8798_, new_n8799_,
    new_n8800_, new_n8801_, new_n8802_, new_n8803_, new_n8804_, new_n8805_,
    new_n8806_, new_n8807_, new_n8808_, new_n8809_, new_n8810_, new_n8811_,
    new_n8812_, new_n8813_, new_n8814_, new_n8815_, new_n8816_, new_n8817_,
    new_n8818_, new_n8819_, new_n8820_, new_n8821_, new_n8822_, new_n8823_,
    new_n8824_, new_n8825_, new_n8826_, new_n8827_, new_n8828_, new_n8829_,
    new_n8830_, new_n8831_, new_n8832_, new_n8833_, new_n8834_, new_n8835_,
    new_n8836_, new_n8837_, new_n8838_, new_n8839_, new_n8840_, new_n8841_,
    new_n8842_, new_n8843_, new_n8844_, new_n8845_, new_n8846_, new_n8847_,
    new_n8848_, new_n8849_, new_n8851_, new_n8852_, new_n8853_, new_n8854_,
    new_n8855_, new_n8856_, new_n8857_, new_n8858_, new_n8859_, new_n8860_,
    new_n8861_, new_n8862_, new_n8863_, new_n8864_, new_n8865_, new_n8866_,
    new_n8867_, new_n8868_, new_n8869_, new_n8870_, new_n8871_, new_n8872_,
    new_n8873_, new_n8874_, new_n8875_, new_n8876_, new_n8877_, new_n8878_,
    new_n8879_, new_n8880_, new_n8881_, new_n8882_, new_n8883_, new_n8884_,
    new_n8885_, new_n8886_, new_n8887_, new_n8888_, new_n8889_, new_n8890_,
    new_n8891_, new_n8892_, new_n8893_, new_n8894_, new_n8895_, new_n8896_,
    new_n8897_, new_n8898_, new_n8899_, new_n8900_, new_n8901_, new_n8902_,
    new_n8903_, new_n8904_, new_n8905_, new_n8906_, new_n8907_, new_n8908_,
    new_n8909_, new_n8910_, new_n8911_, new_n8912_, new_n8913_, new_n8914_,
    new_n8915_, new_n8916_, new_n8917_, new_n8918_, new_n8919_, new_n8920_,
    new_n8921_, new_n8922_, new_n8923_, new_n8924_, new_n8925_, new_n8926_,
    new_n8927_, new_n8928_, new_n8929_, new_n8930_, new_n8931_, new_n8932_,
    new_n8933_, new_n8934_, new_n8935_, new_n8936_, new_n8938_, new_n8939_,
    new_n8940_, new_n8941_, new_n8942_, new_n8943_, new_n8944_, new_n8945_,
    new_n8946_, new_n8947_, new_n8948_, new_n8949_, new_n8950_, new_n8951_,
    new_n8952_, new_n8953_, new_n8954_, new_n8955_, new_n8956_, new_n8957_,
    new_n8958_, new_n8959_, new_n8960_, new_n8961_, new_n8962_, new_n8963_,
    new_n8964_, new_n8965_, new_n8966_, new_n8967_, new_n8968_, new_n8969_,
    new_n8970_, new_n8971_, new_n8972_, new_n8973_, new_n8974_, new_n8975_,
    new_n8976_, new_n8977_, new_n8978_, new_n8979_, new_n8980_, new_n8981_,
    new_n8982_, new_n8983_, new_n8984_, new_n8985_, new_n8986_, new_n8987_,
    new_n8988_, new_n8989_, new_n8990_, new_n8991_, new_n8992_, new_n8993_,
    new_n8994_, new_n8995_, new_n8996_, new_n8997_, new_n8998_, new_n8999_,
    new_n9000_, new_n9001_, new_n9002_, new_n9003_, new_n9004_, new_n9005_,
    new_n9006_, new_n9007_, new_n9008_, new_n9009_, new_n9010_, new_n9011_,
    new_n9012_, new_n9013_, new_n9014_, new_n9015_, new_n9016_, new_n9017_,
    new_n9018_, new_n9019_, new_n9020_, new_n9021_, new_n9022_, new_n9023_,
    new_n9025_, new_n9026_, new_n9027_, new_n9028_, new_n9029_, new_n9030_,
    new_n9031_, new_n9032_, new_n9033_, new_n9034_, new_n9035_, new_n9036_,
    new_n9037_, new_n9038_, new_n9039_, new_n9040_, new_n9041_, new_n9042_,
    new_n9043_, new_n9044_, new_n9045_, new_n9046_, new_n9047_, new_n9048_,
    new_n9049_, new_n9050_, new_n9051_, new_n9052_, new_n9053_, new_n9054_,
    new_n9055_, new_n9056_, new_n9057_, new_n9058_, new_n9059_, new_n9060_,
    new_n9061_, new_n9062_, new_n9063_, new_n9064_, new_n9065_, new_n9066_,
    new_n9067_, new_n9068_, new_n9069_, new_n9070_, new_n9071_, new_n9072_,
    new_n9073_, new_n9074_, new_n9075_, new_n9076_, new_n9077_, new_n9078_,
    new_n9079_, new_n9080_, new_n9081_, new_n9082_, new_n9083_, new_n9084_,
    new_n9085_, new_n9086_, new_n9087_, new_n9088_, new_n9089_, new_n9090_,
    new_n9091_, new_n9092_, new_n9093_, new_n9094_, new_n9095_, new_n9096_,
    new_n9097_, new_n9098_, new_n9099_, new_n9100_, new_n9101_, new_n9102_,
    new_n9103_, new_n9104_, new_n9105_, new_n9106_, new_n9107_, new_n9108_,
    new_n9109_, new_n9110_, new_n9112_, new_n9113_, new_n9114_, new_n9115_,
    new_n9116_, new_n9117_, new_n9118_, new_n9119_, new_n9120_, new_n9121_,
    new_n9122_, new_n9123_, new_n9124_, new_n9125_, new_n9126_, new_n9127_,
    new_n9128_, new_n9129_, new_n9130_, new_n9131_, new_n9132_, new_n9133_,
    new_n9134_, new_n9135_, new_n9136_, new_n9137_, new_n9138_, new_n9139_,
    new_n9140_, new_n9141_, new_n9142_, new_n9143_, new_n9144_, new_n9145_,
    new_n9146_, new_n9147_, new_n9148_, new_n9149_, new_n9150_, new_n9151_,
    new_n9152_, new_n9153_, new_n9154_, new_n9155_, new_n9156_, new_n9157_,
    new_n9158_, new_n9159_, new_n9160_, new_n9161_, new_n9162_, new_n9163_,
    new_n9164_, new_n9165_, new_n9166_, new_n9167_, new_n9168_, new_n9169_,
    new_n9170_, new_n9171_, new_n9172_, new_n9173_, new_n9174_, new_n9175_,
    new_n9176_, new_n9177_, new_n9178_, new_n9179_, new_n9180_, new_n9181_,
    new_n9182_, new_n9183_, new_n9184_, new_n9185_, new_n9186_, new_n9187_,
    new_n9188_, new_n9189_, new_n9190_, new_n9191_, new_n9192_, new_n9193_,
    new_n9194_, new_n9195_, new_n9196_, new_n9197_, new_n9199_, new_n9200_,
    new_n9201_, new_n9202_, new_n9203_, new_n9204_, new_n9205_, new_n9206_,
    new_n9207_, new_n9208_, new_n9209_, new_n9210_, new_n9211_, new_n9212_,
    new_n9213_, new_n9214_, new_n9215_, new_n9216_, new_n9217_, new_n9218_,
    new_n9219_, new_n9220_, new_n9221_, new_n9222_, new_n9223_, new_n9224_,
    new_n9225_, new_n9226_, new_n9227_, new_n9228_, new_n9229_, new_n9230_,
    new_n9231_, new_n9232_, new_n9233_, new_n9234_, new_n9235_, new_n9236_,
    new_n9237_, new_n9238_, new_n9239_, new_n9240_, new_n9241_, new_n9242_,
    new_n9243_, new_n9244_, new_n9245_, new_n9246_, new_n9247_, new_n9248_,
    new_n9249_, new_n9250_, new_n9251_, new_n9252_, new_n9253_, new_n9254_,
    new_n9255_, new_n9256_, new_n9257_, new_n9258_, new_n9259_, new_n9260_,
    new_n9261_, new_n9262_, new_n9263_, new_n9264_, new_n9265_, new_n9266_,
    new_n9267_, new_n9268_, new_n9269_, new_n9270_, new_n9271_, new_n9272_,
    new_n9273_, new_n9274_, new_n9275_, new_n9276_, new_n9277_, new_n9278_,
    new_n9279_, new_n9280_, new_n9281_, new_n9282_, new_n9283_, new_n9284_,
    new_n9286_, new_n9287_, new_n9288_, new_n9289_, new_n9290_, new_n9291_,
    new_n9292_, new_n9293_, new_n9294_, new_n9295_, new_n9296_, new_n9297_,
    new_n9298_, new_n9299_, new_n9300_, new_n9301_, new_n9302_, new_n9303_,
    new_n9304_, new_n9305_, new_n9306_, new_n9307_, new_n9308_, new_n9309_,
    new_n9310_, new_n9311_, new_n9312_, new_n9313_, new_n9314_, new_n9315_,
    new_n9316_, new_n9317_, new_n9318_, new_n9319_, new_n9320_, new_n9321_,
    new_n9322_, new_n9323_, new_n9324_, new_n9325_, new_n9326_, new_n9327_,
    new_n9328_, new_n9329_, new_n9330_, new_n9331_, new_n9332_, new_n9333_,
    new_n9334_, new_n9335_, new_n9336_, new_n9337_, new_n9338_, new_n9339_,
    new_n9340_, new_n9341_, new_n9342_, new_n9343_, new_n9344_, new_n9345_,
    new_n9346_, new_n9347_, new_n9348_, new_n9349_, new_n9350_, new_n9351_,
    new_n9352_, new_n9353_, new_n9354_, new_n9355_, new_n9356_, new_n9357_,
    new_n9358_, new_n9359_, new_n9360_, new_n9361_, new_n9362_, new_n9363_,
    new_n9364_, new_n9365_, new_n9366_, new_n9367_, new_n9368_, new_n9369_,
    new_n9370_, new_n9371_, new_n9373_, new_n9374_, new_n9375_, new_n9376_,
    new_n9377_, new_n9378_, new_n9379_, new_n9380_, new_n9381_, new_n9382_,
    new_n9383_, new_n9384_, new_n9385_, new_n9386_, new_n9387_, new_n9388_,
    new_n9389_, new_n9390_, new_n9391_, new_n9392_, new_n9393_, new_n9394_,
    new_n9395_, new_n9396_, new_n9397_, new_n9398_, new_n9399_, new_n9400_,
    new_n9401_, new_n9402_, new_n9403_, new_n9404_, new_n9405_, new_n9406_,
    new_n9407_, new_n9408_, new_n9409_, new_n9410_, new_n9411_, new_n9412_,
    new_n9413_, new_n9414_, new_n9415_, new_n9416_, new_n9417_, new_n9418_,
    new_n9419_, new_n9420_, new_n9421_, new_n9422_, new_n9423_, new_n9424_,
    new_n9425_, new_n9426_, new_n9427_, new_n9428_, new_n9429_, new_n9430_,
    new_n9431_, new_n9432_, new_n9433_, new_n9434_, new_n9435_, new_n9436_,
    new_n9437_, new_n9438_, new_n9439_, new_n9440_, new_n9441_, new_n9442_,
    new_n9443_, new_n9444_, new_n9445_, new_n9446_, new_n9447_, new_n9448_,
    new_n9449_, new_n9450_, new_n9451_, new_n9452_, new_n9453_, new_n9454_,
    new_n9455_, new_n9456_, new_n9457_, new_n9458_, new_n9460_, new_n9461_,
    new_n9462_, new_n9463_, new_n9464_, new_n9465_, new_n9466_, new_n9467_,
    new_n9468_, new_n9469_, new_n9470_, new_n9471_, new_n9472_, new_n9473_,
    new_n9474_, new_n9475_, new_n9476_, new_n9477_, new_n9478_, new_n9479_,
    new_n9480_, new_n9481_, new_n9482_, new_n9483_, new_n9484_, new_n9485_,
    new_n9486_, new_n9487_, new_n9488_, new_n9489_, new_n9490_, new_n9491_,
    new_n9492_, new_n9493_, new_n9494_, new_n9495_, new_n9496_, new_n9497_,
    new_n9498_, new_n9499_, new_n9500_, new_n9501_, new_n9502_, new_n9503_,
    new_n9504_, new_n9505_, new_n9506_, new_n9507_, new_n9508_, new_n9509_,
    new_n9510_, new_n9511_, new_n9512_, new_n9513_, new_n9514_, new_n9515_,
    new_n9516_, new_n9517_, new_n9518_, new_n9519_, new_n9520_, new_n9521_,
    new_n9522_, new_n9523_, new_n9524_, new_n9525_, new_n9526_, new_n9527_,
    new_n9528_, new_n9529_, new_n9530_, new_n9531_, new_n9532_, new_n9533_,
    new_n9534_, new_n9535_, new_n9536_, new_n9537_, new_n9538_, new_n9539_,
    new_n9540_, new_n9541_, new_n9542_, new_n9543_, new_n9544_, new_n9545_,
    new_n9547_, new_n9548_, new_n9549_, new_n9550_, new_n9551_, new_n9552_,
    new_n9553_, new_n9554_, new_n9555_, new_n9556_, new_n9557_, new_n9558_,
    new_n9559_, new_n9560_, new_n9561_, new_n9562_, new_n9563_, new_n9564_,
    new_n9565_, new_n9566_, new_n9567_, new_n9568_, new_n9569_, new_n9570_,
    new_n9571_, new_n9572_, new_n9573_, new_n9574_, new_n9575_, new_n9576_,
    new_n9577_, new_n9578_, new_n9579_, new_n9580_, new_n9581_, new_n9582_,
    new_n9583_, new_n9584_, new_n9585_, new_n9586_, new_n9587_, new_n9588_,
    new_n9589_, new_n9590_, new_n9591_, new_n9592_, new_n9593_, new_n9594_,
    new_n9595_, new_n9596_, new_n9597_, new_n9598_, new_n9599_, new_n9600_,
    new_n9601_, new_n9602_, new_n9603_, new_n9604_, new_n9605_, new_n9606_,
    new_n9607_, new_n9608_, new_n9609_, new_n9610_, new_n9611_, new_n9612_,
    new_n9613_, new_n9614_, new_n9615_, new_n9616_, new_n9617_, new_n9618_,
    new_n9619_, new_n9620_, new_n9621_, new_n9622_, new_n9623_, new_n9624_,
    new_n9625_, new_n9626_, new_n9627_, new_n9628_, new_n9629_, new_n9630_,
    new_n9631_, new_n9632_, new_n9634_, new_n9635_, new_n9636_, new_n9637_,
    new_n9638_, new_n9639_, new_n9640_, new_n9641_, new_n9642_, new_n9643_,
    new_n9644_, new_n9645_, new_n9646_, new_n9647_, new_n9648_, new_n9649_,
    new_n9650_, new_n9651_, new_n9652_, new_n9653_, new_n9654_, new_n9655_,
    new_n9656_, new_n9657_, new_n9658_, new_n9659_, new_n9660_, new_n9661_,
    new_n9662_, new_n9663_, new_n9664_, new_n9665_, new_n9666_, new_n9667_,
    new_n9668_, new_n9669_, new_n9670_, new_n9671_, new_n9672_, new_n9673_,
    new_n9674_, new_n9675_, new_n9676_, new_n9677_, new_n9678_, new_n9679_,
    new_n9680_, new_n9681_, new_n9682_, new_n9683_, new_n9684_, new_n9685_,
    new_n9686_, new_n9687_, new_n9688_, new_n9689_, new_n9690_, new_n9691_,
    new_n9692_, new_n9693_, new_n9694_, new_n9695_, new_n9696_, new_n9697_,
    new_n9698_, new_n9699_, new_n9700_, new_n9701_, new_n9702_, new_n9703_,
    new_n9704_, new_n9705_, new_n9706_, new_n9707_, new_n9708_, new_n9709_,
    new_n9710_, new_n9711_, new_n9712_, new_n9713_, new_n9714_, new_n9715_,
    new_n9716_, new_n9717_, new_n9718_, new_n9719_, new_n9721_, new_n9722_,
    new_n9723_, new_n9724_, new_n9725_, new_n9726_, new_n9727_, new_n9728_,
    new_n9729_, new_n9730_, new_n9731_, new_n9732_, new_n9733_, new_n9734_,
    new_n9735_, new_n9736_, new_n9737_, new_n9738_, new_n9739_, new_n9740_,
    new_n9741_, new_n9742_, new_n9743_, new_n9744_, new_n9745_, new_n9746_,
    new_n9747_, new_n9748_, new_n9749_, new_n9750_, new_n9751_, new_n9752_,
    new_n9753_, new_n9754_, new_n9755_, new_n9756_, new_n9757_, new_n9758_,
    new_n9759_, new_n9760_, new_n9761_, new_n9762_, new_n9763_, new_n9764_,
    new_n9765_, new_n9766_, new_n9767_, new_n9768_, new_n9769_, new_n9770_,
    new_n9771_, new_n9772_, new_n9773_, new_n9774_, new_n9775_, new_n9776_,
    new_n9777_, new_n9778_, new_n9779_, new_n9780_, new_n9781_, new_n9782_,
    new_n9783_, new_n9784_, new_n9785_, new_n9786_, new_n9787_, new_n9788_,
    new_n9789_, new_n9790_, new_n9791_, new_n9792_, new_n9793_, new_n9794_,
    new_n9795_, new_n9796_, new_n9797_, new_n9798_, new_n9799_, new_n9800_,
    new_n9801_, new_n9802_, new_n9803_, new_n9804_, new_n9805_, new_n9806_,
    new_n9808_, new_n9809_, new_n9810_, new_n9811_, new_n9812_, new_n9813_,
    new_n9814_, new_n9815_, new_n9816_, new_n9817_, new_n9818_, new_n9819_,
    new_n9820_, new_n9821_, new_n9822_, new_n9823_, new_n9824_, new_n9825_,
    new_n9826_, new_n9827_, new_n9828_, new_n9829_, new_n9830_, new_n9831_,
    new_n9832_, new_n9833_, new_n9834_, new_n9835_, new_n9836_, new_n9837_,
    new_n9838_, new_n9839_, new_n9840_, new_n9841_, new_n9842_, new_n9843_,
    new_n9844_, new_n9845_, new_n9846_, new_n9847_, new_n9848_, new_n9849_,
    new_n9850_, new_n9851_, new_n9852_, new_n9853_, new_n9854_, new_n9855_,
    new_n9856_, new_n9857_, new_n9858_, new_n9859_, new_n9860_, new_n9861_,
    new_n9862_, new_n9863_, new_n9864_, new_n9865_, new_n9866_, new_n9867_,
    new_n9868_, new_n9869_, new_n9870_, new_n9871_, new_n9872_, new_n9873_,
    new_n9874_, new_n9875_, new_n9876_, new_n9877_, new_n9878_, new_n9879_,
    new_n9880_, new_n9881_, new_n9882_, new_n9883_, new_n9884_, new_n9885_,
    new_n9886_, new_n9887_, new_n9888_, new_n9889_, new_n9890_, new_n9891_,
    new_n9892_, new_n9893_, new_n9895_, new_n9896_, new_n9897_, new_n9898_,
    new_n9899_, new_n9900_, new_n9901_, new_n9902_, new_n9903_, new_n9904_,
    new_n9905_, new_n9906_, new_n9907_, new_n9908_, new_n9909_, new_n9910_,
    new_n9911_, new_n9912_, new_n9913_, new_n9914_, new_n9915_, new_n9916_,
    new_n9917_, new_n9918_, new_n9919_, new_n9920_, new_n9921_, new_n9922_,
    new_n9923_, new_n9924_, new_n9925_, new_n9926_, new_n9927_, new_n9928_,
    new_n9929_, new_n9930_, new_n9931_, new_n9932_, new_n9933_, new_n9934_,
    new_n9935_, new_n9936_, new_n9937_, new_n9938_, new_n9939_, new_n9940_,
    new_n9941_, new_n9942_, new_n9943_, new_n9944_, new_n9945_, new_n9946_,
    new_n9947_, new_n9948_, new_n9949_, new_n9950_, new_n9951_, new_n9952_,
    new_n9953_, new_n9954_, new_n9955_, new_n9956_, new_n9957_, new_n9958_,
    new_n9959_, new_n9960_, new_n9961_, new_n9962_, new_n9963_, new_n9964_,
    new_n9965_, new_n9966_, new_n9967_, new_n9968_, new_n9969_, new_n9970_,
    new_n9971_, new_n9972_, new_n9973_, new_n9974_, new_n9975_, new_n9976_,
    new_n9977_, new_n9978_, new_n9979_, new_n9980_, new_n9982_, new_n9983_,
    new_n9984_, new_n9985_, new_n9986_, new_n9987_, new_n9988_, new_n9989_,
    new_n9990_, new_n9991_, new_n9992_, new_n9993_, new_n9994_, new_n9995_,
    new_n9996_, new_n9997_, new_n9998_, new_n9999_, new_n10000_,
    new_n10001_, new_n10002_, new_n10003_, new_n10004_, new_n10005_,
    new_n10006_, new_n10007_, new_n10008_, new_n10009_, new_n10010_,
    new_n10011_, new_n10012_, new_n10013_, new_n10014_, new_n10015_,
    new_n10016_, new_n10017_, new_n10018_, new_n10019_, new_n10020_,
    new_n10021_, new_n10022_, new_n10023_, new_n10024_, new_n10025_,
    new_n10026_, new_n10027_, new_n10028_, new_n10029_, new_n10030_,
    new_n10031_, new_n10032_, new_n10033_, new_n10034_, new_n10035_,
    new_n10036_, new_n10037_, new_n10038_, new_n10039_, new_n10040_,
    new_n10041_, new_n10042_, new_n10043_, new_n10044_, new_n10045_,
    new_n10046_, new_n10047_, new_n10048_, new_n10049_, new_n10050_,
    new_n10051_, new_n10052_, new_n10053_, new_n10054_, new_n10055_,
    new_n10056_, new_n10057_, new_n10058_, new_n10059_, new_n10060_,
    new_n10061_, new_n10062_, new_n10063_, new_n10064_, new_n10065_,
    new_n10066_, new_n10067_, new_n10069_, new_n10070_, new_n10071_,
    new_n10072_, new_n10073_, new_n10074_, new_n10075_, new_n10076_,
    new_n10077_, new_n10078_, new_n10079_, new_n10080_, new_n10081_,
    new_n10082_, new_n10083_, new_n10084_, new_n10085_, new_n10086_,
    new_n10087_, new_n10088_, new_n10089_, new_n10090_, new_n10091_,
    new_n10092_, new_n10093_, new_n10094_, new_n10095_, new_n10096_,
    new_n10097_, new_n10098_, new_n10099_, new_n10100_, new_n10101_,
    new_n10102_, new_n10103_, new_n10104_, new_n10105_, new_n10106_,
    new_n10107_, new_n10108_, new_n10109_, new_n10110_, new_n10111_,
    new_n10112_, new_n10113_, new_n10114_, new_n10115_, new_n10116_,
    new_n10117_, new_n10118_, new_n10119_, new_n10120_, new_n10121_,
    new_n10122_, new_n10123_, new_n10124_, new_n10125_, new_n10126_,
    new_n10127_, new_n10128_, new_n10129_, new_n10130_, new_n10131_,
    new_n10132_, new_n10133_, new_n10134_, new_n10135_, new_n10136_,
    new_n10137_, new_n10138_, new_n10139_, new_n10140_, new_n10141_,
    new_n10142_, new_n10143_, new_n10144_, new_n10145_, new_n10146_,
    new_n10147_, new_n10148_, new_n10149_, new_n10150_, new_n10151_,
    new_n10152_, new_n10153_, new_n10154_, new_n10156_, new_n10157_,
    new_n10158_, new_n10159_, new_n10160_, new_n10161_, new_n10162_,
    new_n10163_, new_n10164_, new_n10165_, new_n10166_, new_n10167_,
    new_n10168_, new_n10169_, new_n10170_, new_n10171_, new_n10172_,
    new_n10173_, new_n10174_, new_n10175_, new_n10176_, new_n10177_,
    new_n10178_, new_n10179_, new_n10180_, new_n10181_, new_n10182_,
    new_n10183_, new_n10184_, new_n10185_, new_n10186_, new_n10187_,
    new_n10188_, new_n10189_, new_n10190_, new_n10191_, new_n10192_,
    new_n10193_, new_n10194_, new_n10195_, new_n10196_, new_n10197_,
    new_n10198_, new_n10199_, new_n10200_, new_n10201_, new_n10202_,
    new_n10203_, new_n10204_, new_n10205_, new_n10206_, new_n10207_,
    new_n10208_, new_n10209_, new_n10210_, new_n10211_, new_n10212_,
    new_n10213_, new_n10214_, new_n10215_, new_n10216_, new_n10217_,
    new_n10218_, new_n10219_, new_n10220_, new_n10221_, new_n10222_,
    new_n10223_, new_n10224_, new_n10225_, new_n10226_, new_n10227_,
    new_n10228_, new_n10229_, new_n10230_, new_n10231_, new_n10232_,
    new_n10233_, new_n10234_, new_n10235_, new_n10236_, new_n10237_,
    new_n10238_, new_n10239_, new_n10240_, new_n10241_, new_n10243_,
    new_n10244_, new_n10245_, new_n10246_, new_n10247_, new_n10248_,
    new_n10249_, new_n10250_, new_n10251_, new_n10252_, new_n10253_,
    new_n10254_, new_n10255_, new_n10256_, new_n10257_, new_n10258_,
    new_n10259_, new_n10260_, new_n10261_, new_n10262_, new_n10263_,
    new_n10264_, new_n10265_, new_n10266_, new_n10267_, new_n10268_,
    new_n10269_, new_n10270_, new_n10271_, new_n10272_, new_n10273_,
    new_n10274_, new_n10275_, new_n10276_, new_n10277_, new_n10278_,
    new_n10279_, new_n10280_, new_n10281_, new_n10282_, new_n10283_,
    new_n10284_, new_n10285_, new_n10286_, new_n10287_, new_n10288_,
    new_n10289_, new_n10290_, new_n10291_, new_n10292_, new_n10293_,
    new_n10294_, new_n10295_, new_n10296_, new_n10297_, new_n10298_,
    new_n10299_, new_n10300_, new_n10301_, new_n10302_, new_n10303_,
    new_n10304_, new_n10305_, new_n10306_, new_n10307_, new_n10308_,
    new_n10309_, new_n10310_, new_n10311_, new_n10312_, new_n10313_,
    new_n10314_, new_n10315_, new_n10316_, new_n10317_, new_n10318_,
    new_n10319_, new_n10320_, new_n10321_, new_n10322_, new_n10323_,
    new_n10324_, new_n10325_, new_n10326_, new_n10327_, new_n10328_,
    new_n10330_, new_n10331_, new_n10332_, new_n10333_, new_n10334_,
    new_n10335_, new_n10336_, new_n10337_, new_n10338_, new_n10339_,
    new_n10340_, new_n10341_, new_n10342_, new_n10343_, new_n10344_,
    new_n10345_, new_n10346_, new_n10347_, new_n10348_, new_n10349_,
    new_n10350_, new_n10351_, new_n10352_, new_n10353_, new_n10354_,
    new_n10355_, new_n10356_, new_n10357_, new_n10358_, new_n10359_,
    new_n10360_, new_n10361_, new_n10362_, new_n10363_, new_n10364_,
    new_n10365_, new_n10366_, new_n10367_, new_n10368_, new_n10369_,
    new_n10370_, new_n10371_, new_n10372_, new_n10373_, new_n10374_,
    new_n10375_, new_n10376_, new_n10377_, new_n10378_, new_n10379_,
    new_n10380_, new_n10381_, new_n10382_, new_n10383_, new_n10384_,
    new_n10385_, new_n10386_, new_n10387_, new_n10388_, new_n10389_,
    new_n10390_, new_n10391_, new_n10392_, new_n10393_, new_n10394_,
    new_n10395_, new_n10396_, new_n10397_, new_n10398_, new_n10399_,
    new_n10400_, new_n10401_, new_n10402_, new_n10403_, new_n10404_,
    new_n10405_, new_n10406_, new_n10407_, new_n10408_, new_n10409_,
    new_n10410_, new_n10411_, new_n10412_, new_n10413_, new_n10414_,
    new_n10415_, new_n10417_, new_n10418_, new_n10419_, new_n10420_,
    new_n10421_, new_n10422_, new_n10423_, new_n10424_, new_n10425_,
    new_n10426_, new_n10427_, new_n10428_, new_n10429_, new_n10430_,
    new_n10431_, new_n10432_, new_n10433_, new_n10434_, new_n10435_,
    new_n10436_, new_n10437_, new_n10438_, new_n10439_, new_n10440_,
    new_n10441_, new_n10442_, new_n10443_, new_n10444_, new_n10445_,
    new_n10446_, new_n10447_, new_n10448_, new_n10449_, new_n10450_,
    new_n10451_, new_n10452_, new_n10453_, new_n10454_, new_n10455_,
    new_n10456_, new_n10457_, new_n10458_, new_n10459_, new_n10460_,
    new_n10461_, new_n10462_, new_n10463_, new_n10464_, new_n10465_,
    new_n10466_, new_n10467_, new_n10468_, new_n10469_, new_n10470_,
    new_n10471_, new_n10472_, new_n10473_, new_n10474_, new_n10475_,
    new_n10476_, new_n10477_, new_n10478_, new_n10479_, new_n10480_,
    new_n10481_, new_n10482_, new_n10483_, new_n10484_, new_n10485_,
    new_n10486_, new_n10487_, new_n10488_, new_n10489_, new_n10490_,
    new_n10491_, new_n10492_, new_n10493_, new_n10494_, new_n10495_,
    new_n10496_, new_n10497_, new_n10498_, new_n10499_, new_n10500_,
    new_n10501_, new_n10502_, new_n10504_, new_n10505_, new_n10506_,
    new_n10507_, new_n10508_, new_n10509_, new_n10510_, new_n10511_,
    new_n10512_, new_n10513_, new_n10514_, new_n10515_, new_n10516_,
    new_n10517_, new_n10518_, new_n10519_, new_n10520_, new_n10521_,
    new_n10522_, new_n10523_, new_n10524_, new_n10525_, new_n10526_,
    new_n10527_, new_n10528_, new_n10529_, new_n10530_, new_n10531_,
    new_n10532_, new_n10533_, new_n10534_, new_n10535_, new_n10536_,
    new_n10537_, new_n10538_, new_n10539_, new_n10540_, new_n10541_,
    new_n10542_, new_n10543_, new_n10544_, new_n10545_, new_n10546_,
    new_n10547_, new_n10548_, new_n10549_, new_n10550_, new_n10551_,
    new_n10552_, new_n10553_, new_n10554_, new_n10555_, new_n10556_,
    new_n10557_, new_n10558_, new_n10559_, new_n10560_, new_n10561_,
    new_n10562_, new_n10563_, new_n10564_, new_n10565_, new_n10566_,
    new_n10567_, new_n10568_, new_n10569_, new_n10570_, new_n10571_,
    new_n10572_, new_n10573_, new_n10574_, new_n10575_, new_n10576_,
    new_n10577_, new_n10578_, new_n10579_, new_n10580_, new_n10581_,
    new_n10582_, new_n10583_, new_n10584_, new_n10585_, new_n10586_,
    new_n10587_, new_n10588_, new_n10589_, new_n10591_, new_n10592_,
    new_n10593_, new_n10594_, new_n10595_, new_n10596_, new_n10597_,
    new_n10598_, new_n10599_, new_n10600_, new_n10601_, new_n10602_,
    new_n10603_, new_n10604_, new_n10605_, new_n10606_, new_n10607_,
    new_n10608_, new_n10609_, new_n10610_, new_n10611_, new_n10612_,
    new_n10613_, new_n10614_, new_n10615_, new_n10616_, new_n10617_,
    new_n10618_, new_n10619_, new_n10620_, new_n10621_, new_n10622_,
    new_n10623_, new_n10624_, new_n10625_, new_n10626_, new_n10627_,
    new_n10628_, new_n10629_, new_n10630_, new_n10631_, new_n10632_,
    new_n10633_, new_n10634_, new_n10635_, new_n10636_, new_n10637_,
    new_n10638_, new_n10639_, new_n10640_, new_n10641_, new_n10642_,
    new_n10643_, new_n10644_, new_n10645_, new_n10646_, new_n10647_,
    new_n10648_, new_n10649_, new_n10650_, new_n10651_, new_n10652_,
    new_n10653_, new_n10654_, new_n10655_, new_n10656_, new_n10657_,
    new_n10658_, new_n10659_, new_n10660_, new_n10661_, new_n10662_,
    new_n10663_, new_n10664_, new_n10665_, new_n10666_, new_n10667_,
    new_n10668_, new_n10669_, new_n10670_, new_n10671_, new_n10672_,
    new_n10673_, new_n10674_, new_n10675_, new_n10676_, new_n10678_,
    new_n10679_, new_n10680_, new_n10681_, new_n10682_, new_n10683_,
    new_n10684_, new_n10685_, new_n10686_, new_n10687_, new_n10688_,
    new_n10689_, new_n10690_, new_n10691_, new_n10692_, new_n10693_,
    new_n10694_, new_n10695_, new_n10696_, new_n10697_, new_n10698_,
    new_n10699_, new_n10700_, new_n10701_, new_n10702_, new_n10703_,
    new_n10704_, new_n10705_, new_n10706_, new_n10707_, new_n10708_,
    new_n10709_, new_n10710_, new_n10711_, new_n10712_, new_n10713_,
    new_n10714_, new_n10715_, new_n10716_, new_n10717_, new_n10718_,
    new_n10719_, new_n10720_, new_n10721_, new_n10722_, new_n10723_,
    new_n10724_, new_n10725_, new_n10726_, new_n10727_, new_n10728_,
    new_n10729_, new_n10730_, new_n10731_, new_n10732_, new_n10733_,
    new_n10734_, new_n10735_, new_n10736_, new_n10737_, new_n10738_,
    new_n10739_, new_n10740_, new_n10741_, new_n10742_, new_n10743_,
    new_n10744_, new_n10745_, new_n10746_, new_n10747_, new_n10748_,
    new_n10749_, new_n10750_, new_n10751_, new_n10752_, new_n10753_,
    new_n10754_, new_n10755_, new_n10756_, new_n10757_, new_n10758_,
    new_n10759_, new_n10760_, new_n10761_, new_n10762_, new_n10763_,
    new_n10765_, new_n10766_, new_n10767_, new_n10768_, new_n10769_,
    new_n10770_, new_n10771_, new_n10772_, new_n10773_, new_n10774_,
    new_n10775_, new_n10776_, new_n10777_, new_n10778_, new_n10779_,
    new_n10780_, new_n10781_, new_n10782_, new_n10783_, new_n10784_,
    new_n10785_, new_n10786_, new_n10787_, new_n10788_, new_n10789_,
    new_n10790_, new_n10791_, new_n10792_, new_n10793_, new_n10794_,
    new_n10795_, new_n10796_, new_n10797_, new_n10798_, new_n10799_,
    new_n10800_, new_n10801_, new_n10802_, new_n10803_, new_n10804_,
    new_n10805_, new_n10806_, new_n10807_, new_n10808_, new_n10809_,
    new_n10810_, new_n10811_, new_n10812_, new_n10813_, new_n10814_,
    new_n10815_, new_n10816_, new_n10817_, new_n10818_, new_n10819_,
    new_n10820_, new_n10821_, new_n10822_, new_n10823_, new_n10824_,
    new_n10825_, new_n10826_, new_n10827_, new_n10828_, new_n10829_,
    new_n10830_, new_n10831_, new_n10832_, new_n10833_, new_n10834_,
    new_n10835_, new_n10836_, new_n10837_, new_n10838_, new_n10839_,
    new_n10840_, new_n10841_, new_n10842_, new_n10843_, new_n10844_,
    new_n10845_, new_n10846_, new_n10847_, new_n10848_, new_n10849_,
    new_n10850_, new_n10852_, new_n10853_, new_n10854_, new_n10855_,
    new_n10856_, new_n10857_, new_n10858_, new_n10859_, new_n10860_,
    new_n10861_, new_n10862_, new_n10863_, new_n10864_, new_n10865_,
    new_n10866_, new_n10867_, new_n10868_, new_n10869_, new_n10870_,
    new_n10871_, new_n10872_, new_n10873_, new_n10874_, new_n10875_,
    new_n10876_, new_n10877_, new_n10878_, new_n10879_, new_n10880_,
    new_n10881_, new_n10882_, new_n10883_, new_n10884_, new_n10885_,
    new_n10886_, new_n10887_, new_n10888_, new_n10889_, new_n10890_,
    new_n10891_, new_n10892_, new_n10893_, new_n10894_, new_n10895_,
    new_n10896_, new_n10897_, new_n10898_, new_n10899_, new_n10900_,
    new_n10901_, new_n10902_, new_n10903_, new_n10904_, new_n10905_,
    new_n10906_, new_n10907_, new_n10908_, new_n10909_, new_n10910_,
    new_n10911_, new_n10912_, new_n10913_, new_n10914_, new_n10915_,
    new_n10916_, new_n10917_, new_n10918_, new_n10919_, new_n10920_,
    new_n10921_, new_n10922_, new_n10923_, new_n10924_, new_n10925_,
    new_n10926_, new_n10927_, new_n10928_, new_n10929_, new_n10930_,
    new_n10931_, new_n10932_, new_n10933_, new_n10934_, new_n10935_,
    new_n10936_, new_n10937_, new_n10939_, new_n10940_, new_n10941_,
    new_n10942_, new_n10943_, new_n10944_, new_n10945_, new_n10946_,
    new_n10947_, new_n10948_, new_n10949_, new_n10950_, new_n10951_,
    new_n10952_, new_n10953_, new_n10954_, new_n10955_, new_n10956_,
    new_n10957_, new_n10958_, new_n10959_, new_n10960_, new_n10961_,
    new_n10962_, new_n10963_, new_n10964_, new_n10965_, new_n10966_,
    new_n10967_, new_n10968_, new_n10969_, new_n10970_, new_n10971_,
    new_n10972_, new_n10973_, new_n10974_, new_n10975_, new_n10976_,
    new_n10977_, new_n10978_, new_n10979_, new_n10980_, new_n10981_,
    new_n10982_, new_n10983_, new_n10984_, new_n10985_, new_n10986_,
    new_n10987_, new_n10988_, new_n10989_, new_n10990_, new_n10991_,
    new_n10992_, new_n10993_, new_n10994_, new_n10995_, new_n10996_,
    new_n10997_, new_n10998_, new_n10999_, new_n11000_, new_n11001_,
    new_n11002_, new_n11003_, new_n11004_, new_n11005_, new_n11006_,
    new_n11007_, new_n11008_, new_n11009_, new_n11010_, new_n11011_,
    new_n11012_, new_n11013_, new_n11014_, new_n11015_, new_n11016_,
    new_n11017_, new_n11018_, new_n11019_, new_n11020_, new_n11021_,
    new_n11022_, new_n11023_, new_n11024_, new_n11026_, new_n11027_,
    new_n11028_, new_n11029_, new_n11030_, new_n11031_, new_n11032_,
    new_n11033_, new_n11034_, new_n11035_, new_n11036_, new_n11037_,
    new_n11038_, new_n11039_, new_n11040_, new_n11041_, new_n11042_,
    new_n11043_, new_n11044_, new_n11045_, new_n11046_, new_n11047_,
    new_n11048_, new_n11049_, new_n11050_, new_n11051_, new_n11052_,
    new_n11053_, new_n11054_, new_n11055_, new_n11056_, new_n11057_,
    new_n11058_, new_n11059_, new_n11060_, new_n11061_, new_n11062_,
    new_n11063_, new_n11064_, new_n11065_, new_n11066_, new_n11067_,
    new_n11068_, new_n11069_, new_n11070_, new_n11071_, new_n11072_,
    new_n11073_, new_n11074_, new_n11075_, new_n11076_, new_n11077_,
    new_n11078_, new_n11079_, new_n11080_, new_n11081_, new_n11082_,
    new_n11083_, new_n11084_, new_n11085_, new_n11086_, new_n11087_,
    new_n11088_, new_n11089_, new_n11090_, new_n11091_, new_n11092_,
    new_n11093_, new_n11094_, new_n11095_, new_n11096_, new_n11097_,
    new_n11098_, new_n11099_, new_n11100_, new_n11101_, new_n11102_,
    new_n11103_, new_n11104_, new_n11105_, new_n11106_, new_n11107_,
    new_n11108_, new_n11109_, new_n11110_, new_n11111_, new_n11113_,
    new_n11114_, new_n11115_, new_n11116_, new_n11117_, new_n11118_,
    new_n11119_, new_n11120_, new_n11121_, new_n11122_, new_n11123_,
    new_n11124_, new_n11125_, new_n11126_, new_n11127_, new_n11128_,
    new_n11129_, new_n11130_, new_n11131_, new_n11132_, new_n11133_,
    new_n11134_, new_n11135_, new_n11136_, new_n11137_, new_n11138_,
    new_n11139_, new_n11140_, new_n11141_, new_n11142_, new_n11143_,
    new_n11144_, new_n11145_, new_n11146_, new_n11147_, new_n11148_,
    new_n11149_, new_n11150_, new_n11151_, new_n11152_, new_n11153_,
    new_n11154_, new_n11155_, new_n11156_, new_n11157_, new_n11158_,
    new_n11159_, new_n11160_, new_n11161_, new_n11162_, new_n11163_,
    new_n11164_, new_n11165_, new_n11166_, new_n11167_, new_n11168_,
    new_n11169_, new_n11170_, new_n11171_, new_n11172_, new_n11173_,
    new_n11174_, new_n11175_, new_n11176_, new_n11177_, new_n11178_,
    new_n11179_, new_n11180_, new_n11181_, new_n11182_, new_n11183_,
    new_n11184_, new_n11185_, new_n11186_, new_n11187_, new_n11188_,
    new_n11189_, new_n11190_, new_n11191_, new_n11192_, new_n11193_,
    new_n11194_, new_n11195_, new_n11196_, new_n11197_, new_n11198_,
    new_n11200_, new_n11201_, new_n11202_, new_n11203_, new_n11204_,
    new_n11205_, new_n11206_, new_n11207_, new_n11208_, new_n11209_,
    new_n11210_, new_n11211_, new_n11212_, new_n11213_, new_n11214_,
    new_n11215_, new_n11216_, new_n11217_, new_n11218_, new_n11219_,
    new_n11220_, new_n11221_, new_n11222_, new_n11223_, new_n11224_,
    new_n11225_, new_n11226_, new_n11227_, new_n11228_, new_n11229_,
    new_n11230_, new_n11231_, new_n11232_, new_n11233_, new_n11234_,
    new_n11235_, new_n11236_, new_n11237_, new_n11238_, new_n11239_,
    new_n11240_, new_n11241_, new_n11242_, new_n11243_, new_n11244_,
    new_n11245_, new_n11246_, new_n11247_, new_n11248_, new_n11249_,
    new_n11250_, new_n11251_, new_n11252_, new_n11253_, new_n11254_,
    new_n11255_, new_n11256_, new_n11257_, new_n11258_, new_n11259_,
    new_n11260_, new_n11261_, new_n11262_, new_n11263_, new_n11264_,
    new_n11265_, new_n11266_, new_n11267_, new_n11268_, new_n11269_,
    new_n11270_, new_n11271_, new_n11272_, new_n11273_, new_n11274_,
    new_n11275_, new_n11276_, new_n11277_, new_n11278_, new_n11279_,
    new_n11280_, new_n11281_, new_n11282_, new_n11283_, new_n11284_,
    new_n11285_, new_n11287_, new_n11288_, new_n11289_, new_n11290_,
    new_n11291_, new_n11292_, new_n11293_, new_n11294_, new_n11295_,
    new_n11296_, new_n11297_, new_n11298_, new_n11299_, new_n11300_,
    new_n11301_, new_n11302_, new_n11303_, new_n11304_, new_n11305_,
    new_n11306_, new_n11307_, new_n11308_, new_n11309_, new_n11310_,
    new_n11311_, new_n11312_, new_n11313_, new_n11314_, new_n11315_,
    new_n11316_, new_n11317_, new_n11318_, new_n11319_, new_n11320_,
    new_n11321_, new_n11322_, new_n11323_, new_n11324_, new_n11325_,
    new_n11326_, new_n11327_, new_n11328_, new_n11329_, new_n11330_,
    new_n11331_, new_n11332_, new_n11333_, new_n11334_, new_n11335_,
    new_n11336_, new_n11337_, new_n11338_, new_n11339_, new_n11340_,
    new_n11341_, new_n11342_, new_n11343_, new_n11344_, new_n11345_,
    new_n11346_, new_n11347_, new_n11348_, new_n11349_, new_n11350_,
    new_n11351_, new_n11352_, new_n11353_, new_n11354_, new_n11355_,
    new_n11356_, new_n11357_, new_n11358_, new_n11359_, new_n11360_,
    new_n11361_, new_n11362_, new_n11363_, new_n11364_, new_n11365_,
    new_n11366_, new_n11367_, new_n11368_, new_n11369_, new_n11370_,
    new_n11371_, new_n11372_, new_n11374_, new_n11375_, new_n11376_,
    new_n11377_, new_n11378_, new_n11379_, new_n11380_, new_n11381_,
    new_n11382_, new_n11383_, new_n11384_, new_n11385_, new_n11386_,
    new_n11387_, new_n11388_, new_n11389_, new_n11390_, new_n11391_,
    new_n11392_, new_n11393_, new_n11394_, new_n11395_, new_n11396_,
    new_n11397_, new_n11398_, new_n11399_, new_n11400_, new_n11401_,
    new_n11402_, new_n11403_, new_n11404_, new_n11405_, new_n11406_,
    new_n11407_, new_n11408_, new_n11409_, new_n11410_, new_n11411_,
    new_n11412_, new_n11413_, new_n11414_, new_n11415_, new_n11416_,
    new_n11417_, new_n11418_, new_n11419_, new_n11420_, new_n11421_,
    new_n11422_, new_n11423_, new_n11424_, new_n11425_, new_n11426_,
    new_n11427_, new_n11428_, new_n11429_, new_n11430_, new_n11431_,
    new_n11432_, new_n11433_, new_n11434_, new_n11435_, new_n11436_,
    new_n11437_, new_n11438_, new_n11439_, new_n11440_, new_n11441_,
    new_n11442_, new_n11443_, new_n11444_, new_n11445_, new_n11446_,
    new_n11447_, new_n11448_, new_n11449_, new_n11450_, new_n11451_,
    new_n11452_, new_n11453_, new_n11454_, new_n11455_, new_n11456_,
    new_n11457_, new_n11458_, new_n11459_, new_n11461_, new_n11462_,
    new_n11463_, new_n11464_, new_n11465_, new_n11466_, new_n11467_,
    new_n11468_, new_n11469_, new_n11470_, new_n11471_, new_n11472_,
    new_n11473_, new_n11474_, new_n11475_, new_n11476_, new_n11477_,
    new_n11478_, new_n11479_, new_n11480_, new_n11481_, new_n11482_,
    new_n11483_, new_n11484_, new_n11485_, new_n11486_, new_n11487_,
    new_n11488_, new_n11489_, new_n11490_, new_n11491_, new_n11492_,
    new_n11493_, new_n11494_, new_n11495_, new_n11496_, new_n11497_,
    new_n11498_, new_n11499_, new_n11500_, new_n11501_, new_n11502_,
    new_n11503_, new_n11504_, new_n11505_, new_n11506_, new_n11507_,
    new_n11508_, new_n11509_, new_n11510_, new_n11511_, new_n11512_,
    new_n11513_, new_n11514_, new_n11515_, new_n11516_, new_n11517_,
    new_n11518_, new_n11519_, new_n11520_, new_n11521_, new_n11522_,
    new_n11523_, new_n11524_, new_n11525_, new_n11526_, new_n11527_,
    new_n11528_, new_n11529_, new_n11530_, new_n11531_, new_n11532_,
    new_n11533_, new_n11534_, new_n11535_, new_n11536_, new_n11537_,
    new_n11538_, new_n11539_, new_n11540_, new_n11541_, new_n11542_,
    new_n11543_, new_n11544_, new_n11545_, new_n11546_, new_n11548_,
    new_n11549_, new_n11550_, new_n11551_, new_n11552_, new_n11553_,
    new_n11554_, new_n11555_, new_n11556_, new_n11557_, new_n11558_,
    new_n11559_, new_n11560_, new_n11561_, new_n11562_, new_n11563_,
    new_n11564_, new_n11565_, new_n11566_, new_n11567_, new_n11568_,
    new_n11569_, new_n11570_, new_n11571_, new_n11572_, new_n11573_,
    new_n11574_, new_n11575_, new_n11576_, new_n11577_, new_n11578_,
    new_n11579_, new_n11580_, new_n11581_, new_n11582_, new_n11583_,
    new_n11584_, new_n11585_, new_n11586_, new_n11587_, new_n11588_,
    new_n11589_, new_n11590_, new_n11591_, new_n11592_, new_n11593_,
    new_n11594_, new_n11595_, new_n11596_, new_n11597_, new_n11598_,
    new_n11599_, new_n11600_, new_n11601_, new_n11602_, new_n11603_,
    new_n11604_, new_n11605_, new_n11606_, new_n11607_, new_n11608_,
    new_n11609_, new_n11610_, new_n11611_, new_n11612_, new_n11613_,
    new_n11614_, new_n11615_, new_n11616_, new_n11617_, new_n11618_,
    new_n11619_, new_n11620_, new_n11621_, new_n11622_, new_n11623_,
    new_n11624_, new_n11625_, new_n11626_, new_n11627_, new_n11628_,
    new_n11629_, new_n11630_, new_n11631_, new_n11632_, new_n11633_,
    new_n11635_, new_n11636_, new_n11637_, new_n11638_, new_n11639_,
    new_n11640_, new_n11641_, new_n11642_, new_n11643_, new_n11644_,
    new_n11645_, new_n11646_, new_n11647_, new_n11648_, new_n11649_,
    new_n11650_, new_n11651_, new_n11652_, new_n11653_, new_n11654_,
    new_n11655_, new_n11656_, new_n11657_, new_n11658_, new_n11659_,
    new_n11660_, new_n11661_, new_n11662_, new_n11663_, new_n11664_,
    new_n11665_, new_n11666_, new_n11667_, new_n11668_, new_n11669_,
    new_n11670_, new_n11671_, new_n11672_, new_n11673_, new_n11674_,
    new_n11675_, new_n11676_, new_n11677_, new_n11678_, new_n11679_,
    new_n11680_, new_n11681_, new_n11682_, new_n11683_, new_n11684_,
    new_n11685_, new_n11686_, new_n11687_, new_n11688_, new_n11689_,
    new_n11690_, new_n11691_, new_n11692_, new_n11693_, new_n11694_,
    new_n11695_, new_n11696_, new_n11697_, new_n11698_, new_n11699_,
    new_n11700_, new_n11701_, new_n11702_, new_n11703_, new_n11704_,
    new_n11705_, new_n11706_, new_n11707_, new_n11708_, new_n11709_,
    new_n11710_, new_n11711_, new_n11712_, new_n11713_, new_n11714_,
    new_n11715_, new_n11716_, new_n11717_, new_n11718_, new_n11719_,
    new_n11720_, new_n11722_, new_n11723_, new_n11724_, new_n11725_,
    new_n11726_, new_n11727_, new_n11728_, new_n11729_, new_n11730_,
    new_n11731_, new_n11732_, new_n11733_, new_n11734_, new_n11735_,
    new_n11736_, new_n11737_, new_n11738_, new_n11739_, new_n11740_,
    new_n11741_, new_n11742_, new_n11743_, new_n11744_, new_n11745_,
    new_n11746_, new_n11747_, new_n11748_, new_n11749_, new_n11750_,
    new_n11751_, new_n11752_, new_n11753_, new_n11754_, new_n11755_,
    new_n11756_, new_n11757_, new_n11758_, new_n11759_, new_n11760_,
    new_n11761_, new_n11762_, new_n11763_, new_n11764_, new_n11765_,
    new_n11766_, new_n11767_, new_n11768_, new_n11769_, new_n11770_,
    new_n11771_, new_n11772_, new_n11773_, new_n11774_, new_n11775_,
    new_n11776_, new_n11777_, new_n11778_, new_n11779_, new_n11780_,
    new_n11781_, new_n11782_, new_n11783_, new_n11784_, new_n11785_,
    new_n11786_, new_n11787_, new_n11788_, new_n11789_, new_n11790_,
    new_n11791_, new_n11792_, new_n11793_, new_n11794_, new_n11795_,
    new_n11796_, new_n11797_, new_n11798_, new_n11799_, new_n11800_,
    new_n11801_, new_n11802_, new_n11803_, new_n11804_, new_n11805_,
    new_n11806_, new_n11807_, new_n11809_, new_n11810_, new_n11811_,
    new_n11812_, new_n11813_, new_n11814_, new_n11815_, new_n11816_,
    new_n11817_, new_n11818_, new_n11819_, new_n11820_, new_n11821_,
    new_n11822_, new_n11823_, new_n11824_, new_n11825_, new_n11826_,
    new_n11827_, new_n11828_, new_n11829_, new_n11830_, new_n11831_,
    new_n11832_, new_n11833_, new_n11834_, new_n11835_, new_n11836_,
    new_n11837_, new_n11838_, new_n11839_, new_n11840_, new_n11841_,
    new_n11842_, new_n11843_, new_n11844_, new_n11845_, new_n11846_,
    new_n11847_, new_n11848_, new_n11849_, new_n11850_, new_n11851_,
    new_n11852_, new_n11853_, new_n11854_, new_n11855_, new_n11856_,
    new_n11857_, new_n11858_, new_n11859_, new_n11860_, new_n11861_,
    new_n11862_, new_n11863_, new_n11864_, new_n11865_, new_n11866_,
    new_n11867_, new_n11868_, new_n11869_, new_n11870_, new_n11871_,
    new_n11872_, new_n11873_, new_n11874_, new_n11875_, new_n11876_,
    new_n11877_, new_n11878_, new_n11879_, new_n11880_, new_n11881_,
    new_n11882_, new_n11883_, new_n11884_, new_n11885_, new_n11886_,
    new_n11887_, new_n11888_, new_n11889_, new_n11890_, new_n11891_,
    new_n11892_, new_n11893_, new_n11894_, new_n11896_, new_n11897_,
    new_n11898_, new_n11899_, new_n11900_, new_n11901_, new_n11902_,
    new_n11903_, new_n11904_, new_n11905_, new_n11906_, new_n11907_,
    new_n11908_, new_n11909_, new_n11910_, new_n11911_, new_n11912_,
    new_n11913_, new_n11914_, new_n11915_, new_n11916_, new_n11917_,
    new_n11918_, new_n11919_, new_n11920_, new_n11921_, new_n11922_,
    new_n11923_, new_n11924_, new_n11925_, new_n11926_, new_n11927_,
    new_n11928_, new_n11929_, new_n11930_, new_n11931_, new_n11932_,
    new_n11933_, new_n11934_, new_n11935_, new_n11936_, new_n11937_,
    new_n11938_, new_n11939_, new_n11940_, new_n11941_, new_n11942_,
    new_n11943_, new_n11944_, new_n11945_, new_n11946_, new_n11947_,
    new_n11948_, new_n11949_, new_n11950_, new_n11951_, new_n11952_,
    new_n11953_, new_n11954_, new_n11955_, new_n11956_, new_n11957_,
    new_n11958_, new_n11959_, new_n11960_, new_n11961_, new_n11962_,
    new_n11963_, new_n11964_, new_n11965_, new_n11966_, new_n11967_,
    new_n11968_, new_n11969_, new_n11970_, new_n11971_, new_n11972_,
    new_n11973_, new_n11974_, new_n11975_, new_n11976_, new_n11977_,
    new_n11978_, new_n11979_, new_n11980_, new_n11981_, new_n11983_,
    new_n11984_, new_n11985_, new_n11986_, new_n11987_, new_n11988_,
    new_n11989_, new_n11990_, new_n11991_, new_n11992_, new_n11993_,
    new_n11994_, new_n11995_, new_n11996_, new_n11997_, new_n11998_,
    new_n11999_, new_n12000_, new_n12001_, new_n12002_, new_n12003_,
    new_n12004_, new_n12005_, new_n12006_, new_n12007_, new_n12008_,
    new_n12009_, new_n12010_, new_n12011_, new_n12012_, new_n12013_,
    new_n12014_, new_n12015_, new_n12016_, new_n12017_, new_n12018_,
    new_n12019_, new_n12020_, new_n12021_, new_n12022_, new_n12023_,
    new_n12024_, new_n12025_, new_n12026_, new_n12027_, new_n12028_,
    new_n12029_, new_n12030_, new_n12031_, new_n12032_, new_n12033_,
    new_n12034_, new_n12035_, new_n12036_, new_n12037_, new_n12038_,
    new_n12039_, new_n12040_, new_n12041_, new_n12042_, new_n12043_,
    new_n12044_, new_n12045_, new_n12046_, new_n12047_, new_n12048_,
    new_n12049_, new_n12050_, new_n12051_, new_n12052_, new_n12053_,
    new_n12054_, new_n12055_, new_n12056_, new_n12057_, new_n12058_,
    new_n12059_, new_n12060_, new_n12061_, new_n12062_, new_n12063_,
    new_n12064_, new_n12065_, new_n12066_, new_n12067_, new_n12068_,
    new_n12070_, new_n12071_, new_n12072_, new_n12073_, new_n12074_,
    new_n12075_, new_n12076_, new_n12077_, new_n12078_, new_n12079_,
    new_n12080_, new_n12081_, new_n12082_, new_n12083_, new_n12084_,
    new_n12085_, new_n12086_, new_n12087_, new_n12088_, new_n12089_,
    new_n12090_, new_n12091_, new_n12092_, new_n12093_, new_n12094_,
    new_n12095_, new_n12096_, new_n12097_, new_n12098_, new_n12099_,
    new_n12100_, new_n12101_, new_n12102_, new_n12103_, new_n12104_,
    new_n12105_, new_n12106_, new_n12107_, new_n12108_, new_n12109_,
    new_n12110_, new_n12111_, new_n12112_, new_n12113_, new_n12114_,
    new_n12115_, new_n12116_, new_n12117_, new_n12118_, new_n12119_,
    new_n12120_, new_n12121_, new_n12122_, new_n12123_, new_n12124_,
    new_n12125_, new_n12126_, new_n12127_, new_n12128_, new_n12129_,
    new_n12130_, new_n12131_, new_n12132_, new_n12133_, new_n12134_,
    new_n12135_, new_n12136_, new_n12137_, new_n12138_, new_n12139_,
    new_n12140_, new_n12141_, new_n12142_, new_n12143_, new_n12144_,
    new_n12145_, new_n12146_, new_n12147_, new_n12148_, new_n12149_,
    new_n12150_, new_n12151_, new_n12152_, new_n12153_, new_n12154_,
    new_n12155_, new_n12157_, new_n12158_, new_n12159_, new_n12160_,
    new_n12161_, new_n12162_, new_n12163_, new_n12164_, new_n12165_,
    new_n12166_, new_n12167_, new_n12168_, new_n12169_, new_n12170_,
    new_n12171_, new_n12172_, new_n12173_, new_n12174_, new_n12175_,
    new_n12176_, new_n12177_, new_n12178_, new_n12179_, new_n12180_,
    new_n12181_, new_n12182_, new_n12183_, new_n12184_, new_n12185_,
    new_n12186_, new_n12187_, new_n12188_, new_n12189_, new_n12190_,
    new_n12191_, new_n12192_, new_n12193_, new_n12194_, new_n12195_,
    new_n12196_, new_n12197_, new_n12198_, new_n12199_, new_n12200_,
    new_n12201_, new_n12202_, new_n12203_, new_n12204_, new_n12205_,
    new_n12206_, new_n12207_, new_n12208_, new_n12209_, new_n12210_,
    new_n12211_, new_n12212_, new_n12213_, new_n12214_, new_n12215_,
    new_n12216_, new_n12217_, new_n12218_, new_n12219_, new_n12220_,
    new_n12221_, new_n12222_, new_n12223_, new_n12224_, new_n12225_,
    new_n12226_, new_n12227_, new_n12228_, new_n12229_, new_n12230_,
    new_n12231_, new_n12232_, new_n12233_, new_n12234_, new_n12235_,
    new_n12236_, new_n12237_, new_n12238_, new_n12239_, new_n12240_,
    new_n12241_, new_n12242_, new_n12244_, new_n12245_, new_n12246_,
    new_n12247_, new_n12248_, new_n12249_, new_n12250_, new_n12251_,
    new_n12252_, new_n12253_, new_n12254_, new_n12255_, new_n12256_,
    new_n12257_, new_n12258_, new_n12259_, new_n12260_, new_n12261_,
    new_n12262_, new_n12263_, new_n12264_, new_n12265_, new_n12266_,
    new_n12267_, new_n12268_, new_n12269_, new_n12270_, new_n12271_,
    new_n12272_, new_n12273_, new_n12274_, new_n12275_, new_n12276_,
    new_n12277_, new_n12278_, new_n12279_, new_n12280_, new_n12281_,
    new_n12282_, new_n12283_, new_n12284_, new_n12285_, new_n12286_,
    new_n12287_, new_n12288_, new_n12289_, new_n12290_, new_n12291_,
    new_n12292_, new_n12293_, new_n12294_, new_n12295_, new_n12296_,
    new_n12297_, new_n12298_, new_n12299_, new_n12300_, new_n12301_,
    new_n12302_, new_n12303_, new_n12304_, new_n12305_, new_n12306_,
    new_n12307_, new_n12308_, new_n12309_, new_n12310_, new_n12311_,
    new_n12312_, new_n12313_, new_n12314_, new_n12315_, new_n12316_,
    new_n12317_, new_n12318_, new_n12319_, new_n12320_, new_n12321_,
    new_n12322_, new_n12323_, new_n12324_, new_n12325_, new_n12326_,
    new_n12327_, new_n12328_, new_n12329_, new_n12331_, new_n12332_,
    new_n12333_, new_n12334_, new_n12335_, new_n12336_, new_n12337_,
    new_n12338_, new_n12339_, new_n12340_, new_n12341_, new_n12342_,
    new_n12343_, new_n12344_, new_n12345_, new_n12346_, new_n12347_,
    new_n12348_, new_n12349_, new_n12350_, new_n12351_, new_n12352_,
    new_n12353_, new_n12354_, new_n12355_, new_n12356_, new_n12357_,
    new_n12358_, new_n12359_, new_n12360_, new_n12361_, new_n12362_,
    new_n12363_, new_n12364_, new_n12365_, new_n12366_, new_n12367_,
    new_n12368_, new_n12369_, new_n12370_, new_n12371_, new_n12372_,
    new_n12373_, new_n12374_, new_n12375_, new_n12376_, new_n12377_,
    new_n12378_, new_n12379_, new_n12380_, new_n12381_, new_n12382_,
    new_n12383_, new_n12384_, new_n12385_, new_n12386_, new_n12387_,
    new_n12388_, new_n12389_, new_n12390_, new_n12391_, new_n12392_,
    new_n12393_, new_n12394_, new_n12395_, new_n12396_, new_n12397_,
    new_n12398_, new_n12399_, new_n12400_, new_n12401_, new_n12402_,
    new_n12403_, new_n12404_, new_n12405_, new_n12406_, new_n12407_,
    new_n12408_, new_n12409_, new_n12410_, new_n12411_, new_n12412_,
    new_n12413_, new_n12414_, new_n12415_, new_n12416_, new_n12418_,
    new_n12419_, new_n12420_, new_n12421_, new_n12422_, new_n12423_,
    new_n12424_, new_n12425_, new_n12426_, new_n12427_, new_n12428_,
    new_n12429_, new_n12430_, new_n12431_, new_n12432_, new_n12433_,
    new_n12434_, new_n12435_, new_n12436_, new_n12437_, new_n12438_,
    new_n12439_, new_n12440_, new_n12441_, new_n12442_, new_n12443_,
    new_n12444_, new_n12445_, new_n12446_, new_n12447_, new_n12448_,
    new_n12449_, new_n12450_, new_n12451_, new_n12452_, new_n12453_,
    new_n12454_, new_n12455_, new_n12456_, new_n12457_, new_n12458_,
    new_n12459_, new_n12460_, new_n12461_, new_n12462_, new_n12463_,
    new_n12464_, new_n12465_, new_n12466_, new_n12467_, new_n12468_,
    new_n12469_, new_n12470_, new_n12471_, new_n12472_, new_n12473_,
    new_n12474_, new_n12475_, new_n12476_, new_n12477_, new_n12478_,
    new_n12479_;
  INV   g00000(.A(\priority[1] ), .Y(new_n386_));
  NOR2  g00001(.A(\req[1] ), .B(new_n386_), .Y(new_n387_));
  NOR2  g00002(.A(new_n387_), .B(\priority[2] ), .Y(new_n388_));
  NOR2  g00003(.A(\req[3] ), .B(\req[2] ), .Y(new_n389_));
  INV   g00004(.A(new_n389_), .Y(new_n390_));
  NOR2  g00005(.A(new_n390_), .B(new_n388_), .Y(new_n391_));
  INV   g00006(.A(\priority[5] ), .Y(new_n392_));
  INV   g00007(.A(\priority[3] ), .Y(new_n393_));
  NOR2  g00008(.A(\req[3] ), .B(new_n393_), .Y(new_n394_));
  NOR2  g00009(.A(new_n394_), .B(\priority[4] ), .Y(new_n395_));
  NAND2 g00010(.A(new_n395_), .B(new_n392_), .Y(new_n396_));
  NOR2  g00011(.A(new_n396_), .B(new_n391_), .Y(new_n397_));
  NAND2 g00012(.A(\req[4] ), .B(new_n392_), .Y(new_n398_));
  NOR2  g00013(.A(\req[6] ), .B(\req[5] ), .Y(new_n399_));
  NAND2 g00014(.A(new_n399_), .B(new_n398_), .Y(new_n400_));
  NOR2  g00015(.A(new_n400_), .B(new_n397_), .Y(new_n401_));
  INV   g00016(.A(\priority[8] ), .Y(new_n402_));
  INV   g00017(.A(\priority[6] ), .Y(new_n403_));
  NOR2  g00018(.A(\req[6] ), .B(new_n403_), .Y(new_n404_));
  NOR2  g00019(.A(new_n404_), .B(\priority[7] ), .Y(new_n405_));
  NAND2 g00020(.A(new_n405_), .B(new_n402_), .Y(new_n406_));
  NOR2  g00021(.A(new_n406_), .B(new_n401_), .Y(new_n407_));
  NAND2 g00022(.A(\req[7] ), .B(new_n402_), .Y(new_n408_));
  NOR2  g00023(.A(\req[9] ), .B(\req[8] ), .Y(new_n409_));
  NAND2 g00024(.A(new_n409_), .B(new_n408_), .Y(new_n410_));
  NOR2  g00025(.A(new_n410_), .B(new_n407_), .Y(new_n411_));
  INV   g00026(.A(\priority[11] ), .Y(new_n412_));
  INV   g00027(.A(\priority[9] ), .Y(new_n413_));
  NOR2  g00028(.A(\req[9] ), .B(new_n413_), .Y(new_n414_));
  NOR2  g00029(.A(new_n414_), .B(\priority[10] ), .Y(new_n415_));
  NAND2 g00030(.A(new_n415_), .B(new_n412_), .Y(new_n416_));
  NOR2  g00031(.A(new_n416_), .B(new_n411_), .Y(new_n417_));
  NAND2 g00032(.A(\req[10] ), .B(new_n412_), .Y(new_n418_));
  NOR2  g00033(.A(\req[12] ), .B(\req[11] ), .Y(new_n419_));
  NAND2 g00034(.A(new_n419_), .B(new_n418_), .Y(new_n420_));
  NOR2  g00035(.A(new_n420_), .B(new_n417_), .Y(new_n421_));
  INV   g00036(.A(\priority[14] ), .Y(new_n422_));
  INV   g00037(.A(\priority[12] ), .Y(new_n423_));
  NOR2  g00038(.A(\req[12] ), .B(new_n423_), .Y(new_n424_));
  NOR2  g00039(.A(new_n424_), .B(\priority[13] ), .Y(new_n425_));
  NAND2 g00040(.A(new_n425_), .B(new_n422_), .Y(new_n426_));
  NOR2  g00041(.A(new_n426_), .B(new_n421_), .Y(new_n427_));
  NAND2 g00042(.A(\req[13] ), .B(new_n422_), .Y(new_n428_));
  NOR2  g00043(.A(\req[15] ), .B(\req[14] ), .Y(new_n429_));
  NAND2 g00044(.A(new_n429_), .B(new_n428_), .Y(new_n430_));
  NOR2  g00045(.A(new_n430_), .B(new_n427_), .Y(new_n431_));
  INV   g00046(.A(\priority[17] ), .Y(new_n432_));
  INV   g00047(.A(\priority[15] ), .Y(new_n433_));
  NOR2  g00048(.A(\req[15] ), .B(new_n433_), .Y(new_n434_));
  NOR2  g00049(.A(new_n434_), .B(\priority[16] ), .Y(new_n435_));
  NAND2 g00050(.A(new_n435_), .B(new_n432_), .Y(new_n436_));
  NOR2  g00051(.A(new_n436_), .B(new_n431_), .Y(new_n437_));
  NAND2 g00052(.A(\req[16] ), .B(new_n432_), .Y(new_n438_));
  NOR2  g00053(.A(\req[18] ), .B(\req[17] ), .Y(new_n439_));
  NAND2 g00054(.A(new_n439_), .B(new_n438_), .Y(new_n440_));
  NOR2  g00055(.A(new_n440_), .B(new_n437_), .Y(new_n441_));
  INV   g00056(.A(\priority[20] ), .Y(new_n442_));
  INV   g00057(.A(\priority[18] ), .Y(new_n443_));
  NOR2  g00058(.A(\req[18] ), .B(new_n443_), .Y(new_n444_));
  NOR2  g00059(.A(new_n444_), .B(\priority[19] ), .Y(new_n445_));
  NAND2 g00060(.A(new_n445_), .B(new_n442_), .Y(new_n446_));
  NOR2  g00061(.A(new_n446_), .B(new_n441_), .Y(new_n447_));
  NAND2 g00062(.A(\req[19] ), .B(new_n442_), .Y(new_n448_));
  NOR2  g00063(.A(\req[21] ), .B(\req[20] ), .Y(new_n449_));
  NAND2 g00064(.A(new_n449_), .B(new_n448_), .Y(new_n450_));
  NOR2  g00065(.A(new_n450_), .B(new_n447_), .Y(new_n451_));
  INV   g00066(.A(\priority[23] ), .Y(new_n452_));
  INV   g00067(.A(\priority[21] ), .Y(new_n453_));
  NOR2  g00068(.A(\req[21] ), .B(new_n453_), .Y(new_n454_));
  NOR2  g00069(.A(new_n454_), .B(\priority[22] ), .Y(new_n455_));
  NAND2 g00070(.A(new_n455_), .B(new_n452_), .Y(new_n456_));
  NOR2  g00071(.A(new_n456_), .B(new_n451_), .Y(new_n457_));
  NAND2 g00072(.A(\req[22] ), .B(new_n452_), .Y(new_n458_));
  NOR2  g00073(.A(\req[24] ), .B(\req[23] ), .Y(new_n459_));
  NAND2 g00074(.A(new_n459_), .B(new_n458_), .Y(new_n460_));
  NOR2  g00075(.A(new_n460_), .B(new_n457_), .Y(new_n461_));
  INV   g00076(.A(\priority[26] ), .Y(new_n462_));
  INV   g00077(.A(\priority[24] ), .Y(new_n463_));
  NOR2  g00078(.A(\req[24] ), .B(new_n463_), .Y(new_n464_));
  NOR2  g00079(.A(new_n464_), .B(\priority[25] ), .Y(new_n465_));
  NAND2 g00080(.A(new_n465_), .B(new_n462_), .Y(new_n466_));
  NOR2  g00081(.A(new_n466_), .B(new_n461_), .Y(new_n467_));
  NAND2 g00082(.A(\req[25] ), .B(new_n462_), .Y(new_n468_));
  NOR2  g00083(.A(\req[27] ), .B(\req[26] ), .Y(new_n469_));
  NAND2 g00084(.A(new_n469_), .B(new_n468_), .Y(new_n470_));
  NOR2  g00085(.A(new_n470_), .B(new_n467_), .Y(new_n471_));
  INV   g00086(.A(\priority[29] ), .Y(new_n472_));
  INV   g00087(.A(\priority[27] ), .Y(new_n473_));
  NOR2  g00088(.A(\req[27] ), .B(new_n473_), .Y(new_n474_));
  NOR2  g00089(.A(new_n474_), .B(\priority[28] ), .Y(new_n475_));
  NAND2 g00090(.A(new_n475_), .B(new_n472_), .Y(new_n476_));
  NOR2  g00091(.A(new_n476_), .B(new_n471_), .Y(new_n477_));
  NAND2 g00092(.A(\req[28] ), .B(new_n472_), .Y(new_n478_));
  NOR2  g00093(.A(\req[30] ), .B(\req[29] ), .Y(new_n479_));
  NAND2 g00094(.A(new_n479_), .B(new_n478_), .Y(new_n480_));
  NOR2  g00095(.A(new_n480_), .B(new_n477_), .Y(new_n481_));
  INV   g00096(.A(\priority[32] ), .Y(new_n482_));
  INV   g00097(.A(\priority[30] ), .Y(new_n483_));
  NOR2  g00098(.A(\req[30] ), .B(new_n483_), .Y(new_n484_));
  NOR2  g00099(.A(new_n484_), .B(\priority[31] ), .Y(new_n485_));
  NAND2 g00100(.A(new_n485_), .B(new_n482_), .Y(new_n486_));
  NOR2  g00101(.A(new_n486_), .B(new_n481_), .Y(new_n487_));
  NAND2 g00102(.A(\req[31] ), .B(new_n482_), .Y(new_n488_));
  NOR2  g00103(.A(\req[33] ), .B(\req[32] ), .Y(new_n489_));
  NAND2 g00104(.A(new_n489_), .B(new_n488_), .Y(new_n490_));
  NOR2  g00105(.A(new_n490_), .B(new_n487_), .Y(new_n491_));
  INV   g00106(.A(\priority[35] ), .Y(new_n492_));
  INV   g00107(.A(\priority[33] ), .Y(new_n493_));
  NOR2  g00108(.A(\req[33] ), .B(new_n493_), .Y(new_n494_));
  NOR2  g00109(.A(new_n494_), .B(\priority[34] ), .Y(new_n495_));
  NAND2 g00110(.A(new_n495_), .B(new_n492_), .Y(new_n496_));
  NOR2  g00111(.A(new_n496_), .B(new_n491_), .Y(new_n497_));
  NAND2 g00112(.A(\req[34] ), .B(new_n492_), .Y(new_n498_));
  NOR2  g00113(.A(\req[36] ), .B(\req[35] ), .Y(new_n499_));
  NAND2 g00114(.A(new_n499_), .B(new_n498_), .Y(new_n500_));
  NOR2  g00115(.A(new_n500_), .B(new_n497_), .Y(new_n501_));
  INV   g00116(.A(\priority[38] ), .Y(new_n502_));
  INV   g00117(.A(\priority[36] ), .Y(new_n503_));
  NOR2  g00118(.A(\req[36] ), .B(new_n503_), .Y(new_n504_));
  NOR2  g00119(.A(new_n504_), .B(\priority[37] ), .Y(new_n505_));
  NAND2 g00120(.A(new_n505_), .B(new_n502_), .Y(new_n506_));
  NOR2  g00121(.A(new_n506_), .B(new_n501_), .Y(new_n507_));
  NAND2 g00122(.A(\req[37] ), .B(new_n502_), .Y(new_n508_));
  NOR2  g00123(.A(\req[39] ), .B(\req[38] ), .Y(new_n509_));
  NAND2 g00124(.A(new_n509_), .B(new_n508_), .Y(new_n510_));
  NOR2  g00125(.A(new_n510_), .B(new_n507_), .Y(new_n511_));
  INV   g00126(.A(\priority[41] ), .Y(new_n512_));
  INV   g00127(.A(\priority[39] ), .Y(new_n513_));
  NOR2  g00128(.A(\req[39] ), .B(new_n513_), .Y(new_n514_));
  NOR2  g00129(.A(new_n514_), .B(\priority[40] ), .Y(new_n515_));
  NAND2 g00130(.A(new_n515_), .B(new_n512_), .Y(new_n516_));
  NOR2  g00131(.A(new_n516_), .B(new_n511_), .Y(new_n517_));
  NAND2 g00132(.A(\req[40] ), .B(new_n512_), .Y(new_n518_));
  NOR2  g00133(.A(\req[42] ), .B(\req[41] ), .Y(new_n519_));
  NAND2 g00134(.A(new_n519_), .B(new_n518_), .Y(new_n520_));
  NOR2  g00135(.A(new_n520_), .B(new_n517_), .Y(new_n521_));
  INV   g00136(.A(\priority[44] ), .Y(new_n522_));
  INV   g00137(.A(\priority[42] ), .Y(new_n523_));
  NOR2  g00138(.A(\req[42] ), .B(new_n523_), .Y(new_n524_));
  NOR2  g00139(.A(new_n524_), .B(\priority[43] ), .Y(new_n525_));
  NAND2 g00140(.A(new_n525_), .B(new_n522_), .Y(new_n526_));
  NOR2  g00141(.A(new_n526_), .B(new_n521_), .Y(new_n527_));
  NAND2 g00142(.A(\req[43] ), .B(new_n522_), .Y(new_n528_));
  NOR2  g00143(.A(\req[45] ), .B(\req[44] ), .Y(new_n529_));
  NAND2 g00144(.A(new_n529_), .B(new_n528_), .Y(new_n530_));
  NOR2  g00145(.A(new_n530_), .B(new_n527_), .Y(new_n531_));
  INV   g00146(.A(\priority[47] ), .Y(new_n532_));
  INV   g00147(.A(\priority[45] ), .Y(new_n533_));
  NOR2  g00148(.A(\req[45] ), .B(new_n533_), .Y(new_n534_));
  NOR2  g00149(.A(new_n534_), .B(\priority[46] ), .Y(new_n535_));
  NAND2 g00150(.A(new_n535_), .B(new_n532_), .Y(new_n536_));
  NOR2  g00151(.A(new_n536_), .B(new_n531_), .Y(new_n537_));
  NAND2 g00152(.A(\req[46] ), .B(new_n532_), .Y(new_n538_));
  NOR2  g00153(.A(\req[48] ), .B(\req[47] ), .Y(new_n539_));
  NAND2 g00154(.A(new_n539_), .B(new_n538_), .Y(new_n540_));
  NOR2  g00155(.A(new_n540_), .B(new_n537_), .Y(new_n541_));
  INV   g00156(.A(\priority[50] ), .Y(new_n542_));
  INV   g00157(.A(\priority[48] ), .Y(new_n543_));
  NOR2  g00158(.A(\req[48] ), .B(new_n543_), .Y(new_n544_));
  NOR2  g00159(.A(new_n544_), .B(\priority[49] ), .Y(new_n545_));
  NAND2 g00160(.A(new_n545_), .B(new_n542_), .Y(new_n546_));
  NOR2  g00161(.A(new_n546_), .B(new_n541_), .Y(new_n547_));
  NAND2 g00162(.A(\req[49] ), .B(new_n542_), .Y(new_n548_));
  NOR2  g00163(.A(\req[51] ), .B(\req[50] ), .Y(new_n549_));
  NAND2 g00164(.A(new_n549_), .B(new_n548_), .Y(new_n550_));
  NOR2  g00165(.A(new_n550_), .B(new_n547_), .Y(new_n551_));
  INV   g00166(.A(\priority[53] ), .Y(new_n552_));
  INV   g00167(.A(\priority[51] ), .Y(new_n553_));
  NOR2  g00168(.A(\req[51] ), .B(new_n553_), .Y(new_n554_));
  NOR2  g00169(.A(new_n554_), .B(\priority[52] ), .Y(new_n555_));
  NAND2 g00170(.A(new_n555_), .B(new_n552_), .Y(new_n556_));
  NOR2  g00171(.A(new_n556_), .B(new_n551_), .Y(new_n557_));
  NAND2 g00172(.A(\req[52] ), .B(new_n552_), .Y(new_n558_));
  NOR2  g00173(.A(\req[54] ), .B(\req[53] ), .Y(new_n559_));
  NAND2 g00174(.A(new_n559_), .B(new_n558_), .Y(new_n560_));
  NOR2  g00175(.A(new_n560_), .B(new_n557_), .Y(new_n561_));
  INV   g00176(.A(\priority[56] ), .Y(new_n562_));
  INV   g00177(.A(\priority[54] ), .Y(new_n563_));
  NOR2  g00178(.A(\req[54] ), .B(new_n563_), .Y(new_n564_));
  NOR2  g00179(.A(new_n564_), .B(\priority[55] ), .Y(new_n565_));
  NAND2 g00180(.A(new_n565_), .B(new_n562_), .Y(new_n566_));
  NOR2  g00181(.A(new_n566_), .B(new_n561_), .Y(new_n567_));
  NAND2 g00182(.A(\req[55] ), .B(new_n562_), .Y(new_n568_));
  NOR2  g00183(.A(\req[57] ), .B(\req[56] ), .Y(new_n569_));
  NAND2 g00184(.A(new_n569_), .B(new_n568_), .Y(new_n570_));
  NOR2  g00185(.A(new_n570_), .B(new_n567_), .Y(new_n571_));
  INV   g00186(.A(\priority[59] ), .Y(new_n572_));
  INV   g00187(.A(\priority[57] ), .Y(new_n573_));
  NOR2  g00188(.A(\req[57] ), .B(new_n573_), .Y(new_n574_));
  NOR2  g00189(.A(new_n574_), .B(\priority[58] ), .Y(new_n575_));
  NAND2 g00190(.A(new_n575_), .B(new_n572_), .Y(new_n576_));
  NOR2  g00191(.A(new_n576_), .B(new_n571_), .Y(new_n577_));
  NAND2 g00192(.A(\req[58] ), .B(new_n572_), .Y(new_n578_));
  NOR2  g00193(.A(\req[60] ), .B(\req[59] ), .Y(new_n579_));
  NAND2 g00194(.A(new_n579_), .B(new_n578_), .Y(new_n580_));
  NOR2  g00195(.A(new_n580_), .B(new_n577_), .Y(new_n581_));
  INV   g00196(.A(\priority[62] ), .Y(new_n582_));
  INV   g00197(.A(\priority[60] ), .Y(new_n583_));
  NOR2  g00198(.A(\req[60] ), .B(new_n583_), .Y(new_n584_));
  NOR2  g00199(.A(new_n584_), .B(\priority[61] ), .Y(new_n585_));
  NAND2 g00200(.A(new_n585_), .B(new_n582_), .Y(new_n586_));
  NOR2  g00201(.A(new_n586_), .B(new_n581_), .Y(new_n587_));
  NAND2 g00202(.A(\req[61] ), .B(new_n582_), .Y(new_n588_));
  NOR2  g00203(.A(\req[63] ), .B(\req[62] ), .Y(new_n589_));
  NAND2 g00204(.A(new_n589_), .B(new_n588_), .Y(new_n590_));
  NOR2  g00205(.A(new_n590_), .B(new_n587_), .Y(new_n591_));
  INV   g00206(.A(\priority[65] ), .Y(new_n592_));
  INV   g00207(.A(\priority[63] ), .Y(new_n593_));
  NOR2  g00208(.A(\req[63] ), .B(new_n593_), .Y(new_n594_));
  NOR2  g00209(.A(new_n594_), .B(\priority[64] ), .Y(new_n595_));
  NAND2 g00210(.A(new_n595_), .B(new_n592_), .Y(new_n596_));
  NOR2  g00211(.A(new_n596_), .B(new_n591_), .Y(new_n597_));
  NAND2 g00212(.A(\req[64] ), .B(new_n592_), .Y(new_n598_));
  NOR2  g00213(.A(\req[66] ), .B(\req[65] ), .Y(new_n599_));
  NAND2 g00214(.A(new_n599_), .B(new_n598_), .Y(new_n600_));
  NOR2  g00215(.A(new_n600_), .B(new_n597_), .Y(new_n601_));
  INV   g00216(.A(\priority[68] ), .Y(new_n602_));
  INV   g00217(.A(\priority[66] ), .Y(new_n603_));
  NOR2  g00218(.A(\req[66] ), .B(new_n603_), .Y(new_n604_));
  NOR2  g00219(.A(new_n604_), .B(\priority[67] ), .Y(new_n605_));
  NAND2 g00220(.A(new_n605_), .B(new_n602_), .Y(new_n606_));
  NOR2  g00221(.A(new_n606_), .B(new_n601_), .Y(new_n607_));
  NAND2 g00222(.A(\req[67] ), .B(new_n602_), .Y(new_n608_));
  NOR2  g00223(.A(\req[69] ), .B(\req[68] ), .Y(new_n609_));
  NAND2 g00224(.A(new_n609_), .B(new_n608_), .Y(new_n610_));
  NOR2  g00225(.A(new_n610_), .B(new_n607_), .Y(new_n611_));
  INV   g00226(.A(\priority[71] ), .Y(new_n612_));
  INV   g00227(.A(\priority[69] ), .Y(new_n613_));
  NOR2  g00228(.A(\req[69] ), .B(new_n613_), .Y(new_n614_));
  NOR2  g00229(.A(new_n614_), .B(\priority[70] ), .Y(new_n615_));
  NAND2 g00230(.A(new_n615_), .B(new_n612_), .Y(new_n616_));
  NOR2  g00231(.A(new_n616_), .B(new_n611_), .Y(new_n617_));
  NAND2 g00232(.A(\req[70] ), .B(new_n612_), .Y(new_n618_));
  NOR2  g00233(.A(\req[72] ), .B(\req[71] ), .Y(new_n619_));
  NAND2 g00234(.A(new_n619_), .B(new_n618_), .Y(new_n620_));
  NOR2  g00235(.A(new_n620_), .B(new_n617_), .Y(new_n621_));
  INV   g00236(.A(\priority[74] ), .Y(new_n622_));
  INV   g00237(.A(\priority[72] ), .Y(new_n623_));
  NOR2  g00238(.A(\req[72] ), .B(new_n623_), .Y(new_n624_));
  NOR2  g00239(.A(new_n624_), .B(\priority[73] ), .Y(new_n625_));
  NAND2 g00240(.A(new_n625_), .B(new_n622_), .Y(new_n626_));
  NOR2  g00241(.A(new_n626_), .B(new_n621_), .Y(new_n627_));
  NAND2 g00242(.A(\req[73] ), .B(new_n622_), .Y(new_n628_));
  NOR2  g00243(.A(\req[75] ), .B(\req[74] ), .Y(new_n629_));
  NAND2 g00244(.A(new_n629_), .B(new_n628_), .Y(new_n630_));
  NOR2  g00245(.A(new_n630_), .B(new_n627_), .Y(new_n631_));
  INV   g00246(.A(\priority[77] ), .Y(new_n632_));
  INV   g00247(.A(\priority[75] ), .Y(new_n633_));
  NOR2  g00248(.A(\req[75] ), .B(new_n633_), .Y(new_n634_));
  NOR2  g00249(.A(new_n634_), .B(\priority[76] ), .Y(new_n635_));
  NAND2 g00250(.A(new_n635_), .B(new_n632_), .Y(new_n636_));
  NOR2  g00251(.A(new_n636_), .B(new_n631_), .Y(new_n637_));
  NAND2 g00252(.A(\req[76] ), .B(new_n632_), .Y(new_n638_));
  NOR2  g00253(.A(\req[78] ), .B(\req[77] ), .Y(new_n639_));
  NAND2 g00254(.A(new_n639_), .B(new_n638_), .Y(new_n640_));
  NOR2  g00255(.A(new_n640_), .B(new_n637_), .Y(new_n641_));
  INV   g00256(.A(\priority[80] ), .Y(new_n642_));
  INV   g00257(.A(\priority[78] ), .Y(new_n643_));
  NOR2  g00258(.A(\req[78] ), .B(new_n643_), .Y(new_n644_));
  NOR2  g00259(.A(new_n644_), .B(\priority[79] ), .Y(new_n645_));
  NAND2 g00260(.A(new_n645_), .B(new_n642_), .Y(new_n646_));
  NOR2  g00261(.A(new_n646_), .B(new_n641_), .Y(new_n647_));
  NAND2 g00262(.A(\req[79] ), .B(new_n642_), .Y(new_n648_));
  NOR2  g00263(.A(\req[81] ), .B(\req[80] ), .Y(new_n649_));
  NAND2 g00264(.A(new_n649_), .B(new_n648_), .Y(new_n650_));
  NOR2  g00265(.A(new_n650_), .B(new_n647_), .Y(new_n651_));
  INV   g00266(.A(\priority[83] ), .Y(new_n652_));
  INV   g00267(.A(\priority[81] ), .Y(new_n653_));
  NOR2  g00268(.A(\req[81] ), .B(new_n653_), .Y(new_n654_));
  NOR2  g00269(.A(new_n654_), .B(\priority[82] ), .Y(new_n655_));
  NAND2 g00270(.A(new_n655_), .B(new_n652_), .Y(new_n656_));
  NOR2  g00271(.A(new_n656_), .B(new_n651_), .Y(new_n657_));
  NAND2 g00272(.A(\req[82] ), .B(new_n652_), .Y(new_n658_));
  NOR2  g00273(.A(\req[84] ), .B(\req[83] ), .Y(new_n659_));
  NAND2 g00274(.A(new_n659_), .B(new_n658_), .Y(new_n660_));
  NOR2  g00275(.A(new_n660_), .B(new_n657_), .Y(new_n661_));
  INV   g00276(.A(\priority[86] ), .Y(new_n662_));
  INV   g00277(.A(\priority[84] ), .Y(new_n663_));
  NOR2  g00278(.A(\req[84] ), .B(new_n663_), .Y(new_n664_));
  NOR2  g00279(.A(new_n664_), .B(\priority[85] ), .Y(new_n665_));
  NAND2 g00280(.A(new_n665_), .B(new_n662_), .Y(new_n666_));
  NOR2  g00281(.A(new_n666_), .B(new_n661_), .Y(new_n667_));
  NAND2 g00282(.A(\req[85] ), .B(new_n662_), .Y(new_n668_));
  NOR2  g00283(.A(\req[87] ), .B(\req[86] ), .Y(new_n669_));
  NAND2 g00284(.A(new_n669_), .B(new_n668_), .Y(new_n670_));
  NOR2  g00285(.A(new_n670_), .B(new_n667_), .Y(new_n671_));
  INV   g00286(.A(\priority[89] ), .Y(new_n672_));
  INV   g00287(.A(\priority[87] ), .Y(new_n673_));
  NOR2  g00288(.A(\req[87] ), .B(new_n673_), .Y(new_n674_));
  NOR2  g00289(.A(new_n674_), .B(\priority[88] ), .Y(new_n675_));
  NAND2 g00290(.A(new_n675_), .B(new_n672_), .Y(new_n676_));
  NOR2  g00291(.A(new_n676_), .B(new_n671_), .Y(new_n677_));
  NAND2 g00292(.A(\req[88] ), .B(new_n672_), .Y(new_n678_));
  NOR2  g00293(.A(\req[90] ), .B(\req[89] ), .Y(new_n679_));
  NAND2 g00294(.A(new_n679_), .B(new_n678_), .Y(new_n680_));
  NOR2  g00295(.A(new_n680_), .B(new_n677_), .Y(new_n681_));
  INV   g00296(.A(\priority[92] ), .Y(new_n682_));
  INV   g00297(.A(\priority[90] ), .Y(new_n683_));
  NOR2  g00298(.A(\req[90] ), .B(new_n683_), .Y(new_n684_));
  NOR2  g00299(.A(new_n684_), .B(\priority[91] ), .Y(new_n685_));
  NAND2 g00300(.A(new_n685_), .B(new_n682_), .Y(new_n686_));
  NOR2  g00301(.A(new_n686_), .B(new_n681_), .Y(new_n687_));
  NAND2 g00302(.A(\req[91] ), .B(new_n682_), .Y(new_n688_));
  NOR2  g00303(.A(\req[93] ), .B(\req[92] ), .Y(new_n689_));
  NAND2 g00304(.A(new_n689_), .B(new_n688_), .Y(new_n690_));
  NOR2  g00305(.A(new_n690_), .B(new_n687_), .Y(new_n691_));
  INV   g00306(.A(\priority[95] ), .Y(new_n692_));
  INV   g00307(.A(\priority[93] ), .Y(new_n693_));
  NOR2  g00308(.A(\req[93] ), .B(new_n693_), .Y(new_n694_));
  NOR2  g00309(.A(new_n694_), .B(\priority[94] ), .Y(new_n695_));
  NAND2 g00310(.A(new_n695_), .B(new_n692_), .Y(new_n696_));
  NOR2  g00311(.A(new_n696_), .B(new_n691_), .Y(new_n697_));
  NAND2 g00312(.A(\req[94] ), .B(new_n692_), .Y(new_n698_));
  NOR2  g00313(.A(\req[96] ), .B(\req[95] ), .Y(new_n699_));
  NAND2 g00314(.A(new_n699_), .B(new_n698_), .Y(new_n700_));
  NOR2  g00315(.A(new_n700_), .B(new_n697_), .Y(new_n701_));
  INV   g00316(.A(\priority[98] ), .Y(new_n702_));
  INV   g00317(.A(\priority[96] ), .Y(new_n703_));
  NOR2  g00318(.A(\req[96] ), .B(new_n703_), .Y(new_n704_));
  NOR2  g00319(.A(new_n704_), .B(\priority[97] ), .Y(new_n705_));
  NAND2 g00320(.A(new_n705_), .B(new_n702_), .Y(new_n706_));
  NOR2  g00321(.A(new_n706_), .B(new_n701_), .Y(new_n707_));
  NAND2 g00322(.A(\req[97] ), .B(new_n702_), .Y(new_n708_));
  NOR2  g00323(.A(\req[99] ), .B(\req[98] ), .Y(new_n709_));
  NAND2 g00324(.A(new_n709_), .B(new_n708_), .Y(new_n710_));
  NOR2  g00325(.A(new_n710_), .B(new_n707_), .Y(new_n711_));
  INV   g00326(.A(\priority[101] ), .Y(new_n712_));
  INV   g00327(.A(\priority[99] ), .Y(new_n713_));
  NOR2  g00328(.A(\req[99] ), .B(new_n713_), .Y(new_n714_));
  NOR2  g00329(.A(new_n714_), .B(\priority[100] ), .Y(new_n715_));
  NAND2 g00330(.A(new_n715_), .B(new_n712_), .Y(new_n716_));
  NOR2  g00331(.A(new_n716_), .B(new_n711_), .Y(new_n717_));
  NAND2 g00332(.A(\req[100] ), .B(new_n712_), .Y(new_n718_));
  NOR2  g00333(.A(\req[102] ), .B(\req[101] ), .Y(new_n719_));
  NAND2 g00334(.A(new_n719_), .B(new_n718_), .Y(new_n720_));
  NOR2  g00335(.A(new_n720_), .B(new_n717_), .Y(new_n721_));
  INV   g00336(.A(\priority[104] ), .Y(new_n722_));
  INV   g00337(.A(\priority[102] ), .Y(new_n723_));
  NOR2  g00338(.A(\req[102] ), .B(new_n723_), .Y(new_n724_));
  NOR2  g00339(.A(new_n724_), .B(\priority[103] ), .Y(new_n725_));
  NAND2 g00340(.A(new_n725_), .B(new_n722_), .Y(new_n726_));
  NOR2  g00341(.A(new_n726_), .B(new_n721_), .Y(new_n727_));
  NAND2 g00342(.A(\req[103] ), .B(new_n722_), .Y(new_n728_));
  NOR2  g00343(.A(\req[105] ), .B(\req[104] ), .Y(new_n729_));
  NAND2 g00344(.A(new_n729_), .B(new_n728_), .Y(new_n730_));
  NOR2  g00345(.A(new_n730_), .B(new_n727_), .Y(new_n731_));
  INV   g00346(.A(\priority[107] ), .Y(new_n732_));
  INV   g00347(.A(\priority[105] ), .Y(new_n733_));
  NOR2  g00348(.A(\req[105] ), .B(new_n733_), .Y(new_n734_));
  NOR2  g00349(.A(new_n734_), .B(\priority[106] ), .Y(new_n735_));
  NAND2 g00350(.A(new_n735_), .B(new_n732_), .Y(new_n736_));
  NOR2  g00351(.A(new_n736_), .B(new_n731_), .Y(new_n737_));
  NAND2 g00352(.A(\req[106] ), .B(new_n732_), .Y(new_n738_));
  NOR2  g00353(.A(\req[108] ), .B(\req[107] ), .Y(new_n739_));
  NAND2 g00354(.A(new_n739_), .B(new_n738_), .Y(new_n740_));
  NOR2  g00355(.A(new_n740_), .B(new_n737_), .Y(new_n741_));
  INV   g00356(.A(\priority[110] ), .Y(new_n742_));
  INV   g00357(.A(\priority[108] ), .Y(new_n743_));
  NOR2  g00358(.A(\req[108] ), .B(new_n743_), .Y(new_n744_));
  NOR2  g00359(.A(new_n744_), .B(\priority[109] ), .Y(new_n745_));
  NAND2 g00360(.A(new_n745_), .B(new_n742_), .Y(new_n746_));
  NOR2  g00361(.A(new_n746_), .B(new_n741_), .Y(new_n747_));
  NAND2 g00362(.A(\req[109] ), .B(new_n742_), .Y(new_n748_));
  NOR2  g00363(.A(\req[111] ), .B(\req[110] ), .Y(new_n749_));
  NAND2 g00364(.A(new_n749_), .B(new_n748_), .Y(new_n750_));
  NOR2  g00365(.A(new_n750_), .B(new_n747_), .Y(new_n751_));
  INV   g00366(.A(\priority[113] ), .Y(new_n752_));
  INV   g00367(.A(\priority[111] ), .Y(new_n753_));
  NOR2  g00368(.A(\req[111] ), .B(new_n753_), .Y(new_n754_));
  NOR2  g00369(.A(new_n754_), .B(\priority[112] ), .Y(new_n755_));
  NAND2 g00370(.A(new_n755_), .B(new_n752_), .Y(new_n756_));
  NOR2  g00371(.A(new_n756_), .B(new_n751_), .Y(new_n757_));
  NAND2 g00372(.A(\req[112] ), .B(new_n752_), .Y(new_n758_));
  NOR2  g00373(.A(\req[114] ), .B(\req[113] ), .Y(new_n759_));
  NAND2 g00374(.A(new_n759_), .B(new_n758_), .Y(new_n760_));
  NOR2  g00375(.A(new_n760_), .B(new_n757_), .Y(new_n761_));
  INV   g00376(.A(\priority[116] ), .Y(new_n762_));
  INV   g00377(.A(\priority[114] ), .Y(new_n763_));
  NOR2  g00378(.A(\req[114] ), .B(new_n763_), .Y(new_n764_));
  NOR2  g00379(.A(new_n764_), .B(\priority[115] ), .Y(new_n765_));
  NAND2 g00380(.A(new_n765_), .B(new_n762_), .Y(new_n766_));
  NOR2  g00381(.A(new_n766_), .B(new_n761_), .Y(new_n767_));
  NAND2 g00382(.A(\req[115] ), .B(new_n762_), .Y(new_n768_));
  NOR2  g00383(.A(\req[117] ), .B(\req[116] ), .Y(new_n769_));
  NAND2 g00384(.A(new_n769_), .B(new_n768_), .Y(new_n770_));
  NOR2  g00385(.A(new_n770_), .B(new_n767_), .Y(new_n771_));
  INV   g00386(.A(\priority[119] ), .Y(new_n772_));
  INV   g00387(.A(\priority[117] ), .Y(new_n773_));
  NOR2  g00388(.A(\req[117] ), .B(new_n773_), .Y(new_n774_));
  NOR2  g00389(.A(new_n774_), .B(\priority[118] ), .Y(new_n775_));
  NAND2 g00390(.A(new_n775_), .B(new_n772_), .Y(new_n776_));
  NOR2  g00391(.A(new_n776_), .B(new_n771_), .Y(new_n777_));
  NAND2 g00392(.A(\req[118] ), .B(new_n772_), .Y(new_n778_));
  NOR2  g00393(.A(\req[120] ), .B(\req[119] ), .Y(new_n779_));
  NAND2 g00394(.A(new_n779_), .B(new_n778_), .Y(new_n780_));
  NOR2  g00395(.A(new_n780_), .B(new_n777_), .Y(new_n781_));
  INV   g00396(.A(\priority[122] ), .Y(new_n782_));
  INV   g00397(.A(\priority[120] ), .Y(new_n783_));
  NOR2  g00398(.A(\req[120] ), .B(new_n783_), .Y(new_n784_));
  NOR2  g00399(.A(new_n784_), .B(\priority[121] ), .Y(new_n785_));
  NAND2 g00400(.A(new_n785_), .B(new_n782_), .Y(new_n786_));
  NOR2  g00401(.A(new_n786_), .B(new_n781_), .Y(new_n787_));
  NAND2 g00402(.A(\req[121] ), .B(new_n782_), .Y(new_n788_));
  NOR2  g00403(.A(\req[123] ), .B(\req[122] ), .Y(new_n789_));
  NAND2 g00404(.A(new_n789_), .B(new_n788_), .Y(new_n790_));
  NOR2  g00405(.A(new_n790_), .B(new_n787_), .Y(new_n791_));
  INV   g00406(.A(\priority[125] ), .Y(new_n792_));
  INV   g00407(.A(\priority[123] ), .Y(new_n793_));
  NOR2  g00408(.A(\req[123] ), .B(new_n793_), .Y(new_n794_));
  NOR2  g00409(.A(new_n794_), .B(\priority[124] ), .Y(new_n795_));
  NAND2 g00410(.A(new_n795_), .B(new_n792_), .Y(new_n796_));
  NOR2  g00411(.A(new_n796_), .B(new_n791_), .Y(new_n797_));
  NAND2 g00412(.A(\req[124] ), .B(new_n792_), .Y(new_n798_));
  NOR2  g00413(.A(\req[126] ), .B(\req[125] ), .Y(new_n799_));
  NAND2 g00414(.A(new_n799_), .B(new_n798_), .Y(new_n800_));
  NOR2  g00415(.A(new_n800_), .B(new_n797_), .Y(new_n801_));
  INV   g00416(.A(\priority[0] ), .Y(new_n802_));
  INV   g00417(.A(\priority[126] ), .Y(new_n803_));
  NOR2  g00418(.A(\req[126] ), .B(new_n803_), .Y(new_n804_));
  NOR2  g00419(.A(new_n804_), .B(\priority[127] ), .Y(new_n805_));
  NAND2 g00420(.A(new_n805_), .B(new_n802_), .Y(new_n806_));
  NOR2  g00421(.A(new_n806_), .B(new_n801_), .Y(new_n807_));
  NAND2 g00422(.A(\req[127] ), .B(new_n802_), .Y(new_n808_));
  NAND2 g00423(.A(new_n808_), .B(\req[0] ), .Y(new_n809_));
  NOR2  g00424(.A(new_n809_), .B(new_n807_), .Y(\grant[0] ));
  INV   g00425(.A(\priority[2] ), .Y(new_n811_));
  NOR2  g00426(.A(\req[2] ), .B(new_n811_), .Y(new_n812_));
  NOR2  g00427(.A(new_n812_), .B(\priority[3] ), .Y(new_n813_));
  NOR2  g00428(.A(\req[4] ), .B(\req[3] ), .Y(new_n814_));
  INV   g00429(.A(new_n814_), .Y(new_n815_));
  NOR2  g00430(.A(new_n815_), .B(new_n813_), .Y(new_n816_));
  INV   g00431(.A(\priority[4] ), .Y(new_n817_));
  NOR2  g00432(.A(\req[4] ), .B(new_n817_), .Y(new_n818_));
  NOR2  g00433(.A(new_n818_), .B(\priority[5] ), .Y(new_n819_));
  NAND2 g00434(.A(new_n819_), .B(new_n403_), .Y(new_n820_));
  NOR2  g00435(.A(new_n820_), .B(new_n816_), .Y(new_n821_));
  NAND2 g00436(.A(\req[5] ), .B(new_n403_), .Y(new_n822_));
  NOR2  g00437(.A(\req[7] ), .B(\req[6] ), .Y(new_n823_));
  NAND2 g00438(.A(new_n823_), .B(new_n822_), .Y(new_n824_));
  NOR2  g00439(.A(new_n824_), .B(new_n821_), .Y(new_n825_));
  INV   g00440(.A(\priority[7] ), .Y(new_n826_));
  NOR2  g00441(.A(\req[7] ), .B(new_n826_), .Y(new_n827_));
  NOR2  g00442(.A(new_n827_), .B(\priority[8] ), .Y(new_n828_));
  NAND2 g00443(.A(new_n828_), .B(new_n413_), .Y(new_n829_));
  NOR2  g00444(.A(new_n829_), .B(new_n825_), .Y(new_n830_));
  NAND2 g00445(.A(\req[8] ), .B(new_n413_), .Y(new_n831_));
  NOR2  g00446(.A(\req[10] ), .B(\req[9] ), .Y(new_n832_));
  NAND2 g00447(.A(new_n832_), .B(new_n831_), .Y(new_n833_));
  NOR2  g00448(.A(new_n833_), .B(new_n830_), .Y(new_n834_));
  INV   g00449(.A(\priority[10] ), .Y(new_n835_));
  NOR2  g00450(.A(\req[10] ), .B(new_n835_), .Y(new_n836_));
  NOR2  g00451(.A(new_n836_), .B(\priority[11] ), .Y(new_n837_));
  NAND2 g00452(.A(new_n837_), .B(new_n423_), .Y(new_n838_));
  NOR2  g00453(.A(new_n838_), .B(new_n834_), .Y(new_n839_));
  NAND2 g00454(.A(\req[11] ), .B(new_n423_), .Y(new_n840_));
  NOR2  g00455(.A(\req[13] ), .B(\req[12] ), .Y(new_n841_));
  NAND2 g00456(.A(new_n841_), .B(new_n840_), .Y(new_n842_));
  NOR2  g00457(.A(new_n842_), .B(new_n839_), .Y(new_n843_));
  INV   g00458(.A(\priority[13] ), .Y(new_n844_));
  NOR2  g00459(.A(\req[13] ), .B(new_n844_), .Y(new_n845_));
  NOR2  g00460(.A(new_n845_), .B(\priority[14] ), .Y(new_n846_));
  NAND2 g00461(.A(new_n846_), .B(new_n433_), .Y(new_n847_));
  NOR2  g00462(.A(new_n847_), .B(new_n843_), .Y(new_n848_));
  NAND2 g00463(.A(\req[14] ), .B(new_n433_), .Y(new_n849_));
  NOR2  g00464(.A(\req[16] ), .B(\req[15] ), .Y(new_n850_));
  NAND2 g00465(.A(new_n850_), .B(new_n849_), .Y(new_n851_));
  NOR2  g00466(.A(new_n851_), .B(new_n848_), .Y(new_n852_));
  INV   g00467(.A(\priority[16] ), .Y(new_n853_));
  NOR2  g00468(.A(\req[16] ), .B(new_n853_), .Y(new_n854_));
  NOR2  g00469(.A(new_n854_), .B(\priority[17] ), .Y(new_n855_));
  NAND2 g00470(.A(new_n855_), .B(new_n443_), .Y(new_n856_));
  NOR2  g00471(.A(new_n856_), .B(new_n852_), .Y(new_n857_));
  NAND2 g00472(.A(\req[17] ), .B(new_n443_), .Y(new_n858_));
  NOR2  g00473(.A(\req[19] ), .B(\req[18] ), .Y(new_n859_));
  NAND2 g00474(.A(new_n859_), .B(new_n858_), .Y(new_n860_));
  NOR2  g00475(.A(new_n860_), .B(new_n857_), .Y(new_n861_));
  INV   g00476(.A(\priority[19] ), .Y(new_n862_));
  NOR2  g00477(.A(\req[19] ), .B(new_n862_), .Y(new_n863_));
  NOR2  g00478(.A(new_n863_), .B(\priority[20] ), .Y(new_n864_));
  NAND2 g00479(.A(new_n864_), .B(new_n453_), .Y(new_n865_));
  NOR2  g00480(.A(new_n865_), .B(new_n861_), .Y(new_n866_));
  NAND2 g00481(.A(\req[20] ), .B(new_n453_), .Y(new_n867_));
  NOR2  g00482(.A(\req[22] ), .B(\req[21] ), .Y(new_n868_));
  NAND2 g00483(.A(new_n868_), .B(new_n867_), .Y(new_n869_));
  NOR2  g00484(.A(new_n869_), .B(new_n866_), .Y(new_n870_));
  INV   g00485(.A(\priority[22] ), .Y(new_n871_));
  NOR2  g00486(.A(\req[22] ), .B(new_n871_), .Y(new_n872_));
  NOR2  g00487(.A(new_n872_), .B(\priority[23] ), .Y(new_n873_));
  NAND2 g00488(.A(new_n873_), .B(new_n463_), .Y(new_n874_));
  NOR2  g00489(.A(new_n874_), .B(new_n870_), .Y(new_n875_));
  NAND2 g00490(.A(\req[23] ), .B(new_n463_), .Y(new_n876_));
  NOR2  g00491(.A(\req[25] ), .B(\req[24] ), .Y(new_n877_));
  NAND2 g00492(.A(new_n877_), .B(new_n876_), .Y(new_n878_));
  NOR2  g00493(.A(new_n878_), .B(new_n875_), .Y(new_n879_));
  INV   g00494(.A(\priority[25] ), .Y(new_n880_));
  NOR2  g00495(.A(\req[25] ), .B(new_n880_), .Y(new_n881_));
  NOR2  g00496(.A(new_n881_), .B(\priority[26] ), .Y(new_n882_));
  NAND2 g00497(.A(new_n882_), .B(new_n473_), .Y(new_n883_));
  NOR2  g00498(.A(new_n883_), .B(new_n879_), .Y(new_n884_));
  NAND2 g00499(.A(\req[26] ), .B(new_n473_), .Y(new_n885_));
  NOR2  g00500(.A(\req[28] ), .B(\req[27] ), .Y(new_n886_));
  NAND2 g00501(.A(new_n886_), .B(new_n885_), .Y(new_n887_));
  NOR2  g00502(.A(new_n887_), .B(new_n884_), .Y(new_n888_));
  INV   g00503(.A(\priority[28] ), .Y(new_n889_));
  NOR2  g00504(.A(\req[28] ), .B(new_n889_), .Y(new_n890_));
  NOR2  g00505(.A(new_n890_), .B(\priority[29] ), .Y(new_n891_));
  NAND2 g00506(.A(new_n891_), .B(new_n483_), .Y(new_n892_));
  NOR2  g00507(.A(new_n892_), .B(new_n888_), .Y(new_n893_));
  NAND2 g00508(.A(\req[29] ), .B(new_n483_), .Y(new_n894_));
  NOR2  g00509(.A(\req[31] ), .B(\req[30] ), .Y(new_n895_));
  NAND2 g00510(.A(new_n895_), .B(new_n894_), .Y(new_n896_));
  NOR2  g00511(.A(new_n896_), .B(new_n893_), .Y(new_n897_));
  INV   g00512(.A(\priority[31] ), .Y(new_n898_));
  NOR2  g00513(.A(\req[31] ), .B(new_n898_), .Y(new_n899_));
  NOR2  g00514(.A(new_n899_), .B(\priority[32] ), .Y(new_n900_));
  NAND2 g00515(.A(new_n900_), .B(new_n493_), .Y(new_n901_));
  NOR2  g00516(.A(new_n901_), .B(new_n897_), .Y(new_n902_));
  NAND2 g00517(.A(\req[32] ), .B(new_n493_), .Y(new_n903_));
  NOR2  g00518(.A(\req[34] ), .B(\req[33] ), .Y(new_n904_));
  NAND2 g00519(.A(new_n904_), .B(new_n903_), .Y(new_n905_));
  NOR2  g00520(.A(new_n905_), .B(new_n902_), .Y(new_n906_));
  INV   g00521(.A(\priority[34] ), .Y(new_n907_));
  NOR2  g00522(.A(\req[34] ), .B(new_n907_), .Y(new_n908_));
  NOR2  g00523(.A(new_n908_), .B(\priority[35] ), .Y(new_n909_));
  NAND2 g00524(.A(new_n909_), .B(new_n503_), .Y(new_n910_));
  NOR2  g00525(.A(new_n910_), .B(new_n906_), .Y(new_n911_));
  NAND2 g00526(.A(\req[35] ), .B(new_n503_), .Y(new_n912_));
  NOR2  g00527(.A(\req[37] ), .B(\req[36] ), .Y(new_n913_));
  NAND2 g00528(.A(new_n913_), .B(new_n912_), .Y(new_n914_));
  NOR2  g00529(.A(new_n914_), .B(new_n911_), .Y(new_n915_));
  INV   g00530(.A(\priority[37] ), .Y(new_n916_));
  NOR2  g00531(.A(\req[37] ), .B(new_n916_), .Y(new_n917_));
  NOR2  g00532(.A(new_n917_), .B(\priority[38] ), .Y(new_n918_));
  NAND2 g00533(.A(new_n918_), .B(new_n513_), .Y(new_n919_));
  NOR2  g00534(.A(new_n919_), .B(new_n915_), .Y(new_n920_));
  NAND2 g00535(.A(\req[38] ), .B(new_n513_), .Y(new_n921_));
  NOR2  g00536(.A(\req[40] ), .B(\req[39] ), .Y(new_n922_));
  NAND2 g00537(.A(new_n922_), .B(new_n921_), .Y(new_n923_));
  NOR2  g00538(.A(new_n923_), .B(new_n920_), .Y(new_n924_));
  INV   g00539(.A(\priority[40] ), .Y(new_n925_));
  NOR2  g00540(.A(\req[40] ), .B(new_n925_), .Y(new_n926_));
  NOR2  g00541(.A(new_n926_), .B(\priority[41] ), .Y(new_n927_));
  NAND2 g00542(.A(new_n927_), .B(new_n523_), .Y(new_n928_));
  NOR2  g00543(.A(new_n928_), .B(new_n924_), .Y(new_n929_));
  NAND2 g00544(.A(\req[41] ), .B(new_n523_), .Y(new_n930_));
  NOR2  g00545(.A(\req[43] ), .B(\req[42] ), .Y(new_n931_));
  NAND2 g00546(.A(new_n931_), .B(new_n930_), .Y(new_n932_));
  NOR2  g00547(.A(new_n932_), .B(new_n929_), .Y(new_n933_));
  INV   g00548(.A(\priority[43] ), .Y(new_n934_));
  NOR2  g00549(.A(\req[43] ), .B(new_n934_), .Y(new_n935_));
  NOR2  g00550(.A(new_n935_), .B(\priority[44] ), .Y(new_n936_));
  NAND2 g00551(.A(new_n936_), .B(new_n533_), .Y(new_n937_));
  NOR2  g00552(.A(new_n937_), .B(new_n933_), .Y(new_n938_));
  NAND2 g00553(.A(\req[44] ), .B(new_n533_), .Y(new_n939_));
  NOR2  g00554(.A(\req[46] ), .B(\req[45] ), .Y(new_n940_));
  NAND2 g00555(.A(new_n940_), .B(new_n939_), .Y(new_n941_));
  NOR2  g00556(.A(new_n941_), .B(new_n938_), .Y(new_n942_));
  INV   g00557(.A(\priority[46] ), .Y(new_n943_));
  NOR2  g00558(.A(\req[46] ), .B(new_n943_), .Y(new_n944_));
  NOR2  g00559(.A(new_n944_), .B(\priority[47] ), .Y(new_n945_));
  NAND2 g00560(.A(new_n945_), .B(new_n543_), .Y(new_n946_));
  NOR2  g00561(.A(new_n946_), .B(new_n942_), .Y(new_n947_));
  NAND2 g00562(.A(\req[47] ), .B(new_n543_), .Y(new_n948_));
  NOR2  g00563(.A(\req[49] ), .B(\req[48] ), .Y(new_n949_));
  NAND2 g00564(.A(new_n949_), .B(new_n948_), .Y(new_n950_));
  NOR2  g00565(.A(new_n950_), .B(new_n947_), .Y(new_n951_));
  INV   g00566(.A(\priority[49] ), .Y(new_n952_));
  NOR2  g00567(.A(\req[49] ), .B(new_n952_), .Y(new_n953_));
  NOR2  g00568(.A(new_n953_), .B(\priority[50] ), .Y(new_n954_));
  NAND2 g00569(.A(new_n954_), .B(new_n553_), .Y(new_n955_));
  NOR2  g00570(.A(new_n955_), .B(new_n951_), .Y(new_n956_));
  NAND2 g00571(.A(\req[50] ), .B(new_n553_), .Y(new_n957_));
  NOR2  g00572(.A(\req[52] ), .B(\req[51] ), .Y(new_n958_));
  NAND2 g00573(.A(new_n958_), .B(new_n957_), .Y(new_n959_));
  NOR2  g00574(.A(new_n959_), .B(new_n956_), .Y(new_n960_));
  INV   g00575(.A(\priority[52] ), .Y(new_n961_));
  NOR2  g00576(.A(\req[52] ), .B(new_n961_), .Y(new_n962_));
  NOR2  g00577(.A(new_n962_), .B(\priority[53] ), .Y(new_n963_));
  NAND2 g00578(.A(new_n963_), .B(new_n563_), .Y(new_n964_));
  NOR2  g00579(.A(new_n964_), .B(new_n960_), .Y(new_n965_));
  NAND2 g00580(.A(\req[53] ), .B(new_n563_), .Y(new_n966_));
  NOR2  g00581(.A(\req[55] ), .B(\req[54] ), .Y(new_n967_));
  NAND2 g00582(.A(new_n967_), .B(new_n966_), .Y(new_n968_));
  NOR2  g00583(.A(new_n968_), .B(new_n965_), .Y(new_n969_));
  INV   g00584(.A(\priority[55] ), .Y(new_n970_));
  NOR2  g00585(.A(\req[55] ), .B(new_n970_), .Y(new_n971_));
  NOR2  g00586(.A(new_n971_), .B(\priority[56] ), .Y(new_n972_));
  NAND2 g00587(.A(new_n972_), .B(new_n573_), .Y(new_n973_));
  NOR2  g00588(.A(new_n973_), .B(new_n969_), .Y(new_n974_));
  NAND2 g00589(.A(\req[56] ), .B(new_n573_), .Y(new_n975_));
  NOR2  g00590(.A(\req[58] ), .B(\req[57] ), .Y(new_n976_));
  NAND2 g00591(.A(new_n976_), .B(new_n975_), .Y(new_n977_));
  NOR2  g00592(.A(new_n977_), .B(new_n974_), .Y(new_n978_));
  INV   g00593(.A(\priority[58] ), .Y(new_n979_));
  NOR2  g00594(.A(\req[58] ), .B(new_n979_), .Y(new_n980_));
  NOR2  g00595(.A(new_n980_), .B(\priority[59] ), .Y(new_n981_));
  NAND2 g00596(.A(new_n981_), .B(new_n583_), .Y(new_n982_));
  NOR2  g00597(.A(new_n982_), .B(new_n978_), .Y(new_n983_));
  NAND2 g00598(.A(\req[59] ), .B(new_n583_), .Y(new_n984_));
  NOR2  g00599(.A(\req[61] ), .B(\req[60] ), .Y(new_n985_));
  NAND2 g00600(.A(new_n985_), .B(new_n984_), .Y(new_n986_));
  NOR2  g00601(.A(new_n986_), .B(new_n983_), .Y(new_n987_));
  INV   g00602(.A(\priority[61] ), .Y(new_n988_));
  NOR2  g00603(.A(\req[61] ), .B(new_n988_), .Y(new_n989_));
  NOR2  g00604(.A(new_n989_), .B(\priority[62] ), .Y(new_n990_));
  NAND2 g00605(.A(new_n990_), .B(new_n593_), .Y(new_n991_));
  NOR2  g00606(.A(new_n991_), .B(new_n987_), .Y(new_n992_));
  NAND2 g00607(.A(\req[62] ), .B(new_n593_), .Y(new_n993_));
  NOR2  g00608(.A(\req[64] ), .B(\req[63] ), .Y(new_n994_));
  NAND2 g00609(.A(new_n994_), .B(new_n993_), .Y(new_n995_));
  NOR2  g00610(.A(new_n995_), .B(new_n992_), .Y(new_n996_));
  INV   g00611(.A(\priority[64] ), .Y(new_n997_));
  NOR2  g00612(.A(\req[64] ), .B(new_n997_), .Y(new_n998_));
  NOR2  g00613(.A(new_n998_), .B(\priority[65] ), .Y(new_n999_));
  NAND2 g00614(.A(new_n999_), .B(new_n603_), .Y(new_n1000_));
  NOR2  g00615(.A(new_n1000_), .B(new_n996_), .Y(new_n1001_));
  NAND2 g00616(.A(\req[65] ), .B(new_n603_), .Y(new_n1002_));
  NOR2  g00617(.A(\req[67] ), .B(\req[66] ), .Y(new_n1003_));
  NAND2 g00618(.A(new_n1003_), .B(new_n1002_), .Y(new_n1004_));
  NOR2  g00619(.A(new_n1004_), .B(new_n1001_), .Y(new_n1005_));
  INV   g00620(.A(\priority[67] ), .Y(new_n1006_));
  NOR2  g00621(.A(\req[67] ), .B(new_n1006_), .Y(new_n1007_));
  NOR2  g00622(.A(new_n1007_), .B(\priority[68] ), .Y(new_n1008_));
  NAND2 g00623(.A(new_n1008_), .B(new_n613_), .Y(new_n1009_));
  NOR2  g00624(.A(new_n1009_), .B(new_n1005_), .Y(new_n1010_));
  NAND2 g00625(.A(\req[68] ), .B(new_n613_), .Y(new_n1011_));
  NOR2  g00626(.A(\req[70] ), .B(\req[69] ), .Y(new_n1012_));
  NAND2 g00627(.A(new_n1012_), .B(new_n1011_), .Y(new_n1013_));
  NOR2  g00628(.A(new_n1013_), .B(new_n1010_), .Y(new_n1014_));
  INV   g00629(.A(\priority[70] ), .Y(new_n1015_));
  NOR2  g00630(.A(\req[70] ), .B(new_n1015_), .Y(new_n1016_));
  NOR2  g00631(.A(new_n1016_), .B(\priority[71] ), .Y(new_n1017_));
  NAND2 g00632(.A(new_n1017_), .B(new_n623_), .Y(new_n1018_));
  NOR2  g00633(.A(new_n1018_), .B(new_n1014_), .Y(new_n1019_));
  NAND2 g00634(.A(\req[71] ), .B(new_n623_), .Y(new_n1020_));
  NOR2  g00635(.A(\req[73] ), .B(\req[72] ), .Y(new_n1021_));
  NAND2 g00636(.A(new_n1021_), .B(new_n1020_), .Y(new_n1022_));
  NOR2  g00637(.A(new_n1022_), .B(new_n1019_), .Y(new_n1023_));
  INV   g00638(.A(\priority[73] ), .Y(new_n1024_));
  NOR2  g00639(.A(\req[73] ), .B(new_n1024_), .Y(new_n1025_));
  NOR2  g00640(.A(new_n1025_), .B(\priority[74] ), .Y(new_n1026_));
  NAND2 g00641(.A(new_n1026_), .B(new_n633_), .Y(new_n1027_));
  NOR2  g00642(.A(new_n1027_), .B(new_n1023_), .Y(new_n1028_));
  NAND2 g00643(.A(\req[74] ), .B(new_n633_), .Y(new_n1029_));
  NOR2  g00644(.A(\req[76] ), .B(\req[75] ), .Y(new_n1030_));
  NAND2 g00645(.A(new_n1030_), .B(new_n1029_), .Y(new_n1031_));
  NOR2  g00646(.A(new_n1031_), .B(new_n1028_), .Y(new_n1032_));
  INV   g00647(.A(\priority[76] ), .Y(new_n1033_));
  NOR2  g00648(.A(\req[76] ), .B(new_n1033_), .Y(new_n1034_));
  NOR2  g00649(.A(new_n1034_), .B(\priority[77] ), .Y(new_n1035_));
  NAND2 g00650(.A(new_n1035_), .B(new_n643_), .Y(new_n1036_));
  NOR2  g00651(.A(new_n1036_), .B(new_n1032_), .Y(new_n1037_));
  NAND2 g00652(.A(\req[77] ), .B(new_n643_), .Y(new_n1038_));
  NOR2  g00653(.A(\req[79] ), .B(\req[78] ), .Y(new_n1039_));
  NAND2 g00654(.A(new_n1039_), .B(new_n1038_), .Y(new_n1040_));
  NOR2  g00655(.A(new_n1040_), .B(new_n1037_), .Y(new_n1041_));
  INV   g00656(.A(\priority[79] ), .Y(new_n1042_));
  NOR2  g00657(.A(\req[79] ), .B(new_n1042_), .Y(new_n1043_));
  NOR2  g00658(.A(new_n1043_), .B(\priority[80] ), .Y(new_n1044_));
  NAND2 g00659(.A(new_n1044_), .B(new_n653_), .Y(new_n1045_));
  NOR2  g00660(.A(new_n1045_), .B(new_n1041_), .Y(new_n1046_));
  NAND2 g00661(.A(\req[80] ), .B(new_n653_), .Y(new_n1047_));
  NOR2  g00662(.A(\req[82] ), .B(\req[81] ), .Y(new_n1048_));
  NAND2 g00663(.A(new_n1048_), .B(new_n1047_), .Y(new_n1049_));
  NOR2  g00664(.A(new_n1049_), .B(new_n1046_), .Y(new_n1050_));
  INV   g00665(.A(\priority[82] ), .Y(new_n1051_));
  NOR2  g00666(.A(\req[82] ), .B(new_n1051_), .Y(new_n1052_));
  NOR2  g00667(.A(new_n1052_), .B(\priority[83] ), .Y(new_n1053_));
  NAND2 g00668(.A(new_n1053_), .B(new_n663_), .Y(new_n1054_));
  NOR2  g00669(.A(new_n1054_), .B(new_n1050_), .Y(new_n1055_));
  NAND2 g00670(.A(\req[83] ), .B(new_n663_), .Y(new_n1056_));
  NOR2  g00671(.A(\req[85] ), .B(\req[84] ), .Y(new_n1057_));
  NAND2 g00672(.A(new_n1057_), .B(new_n1056_), .Y(new_n1058_));
  NOR2  g00673(.A(new_n1058_), .B(new_n1055_), .Y(new_n1059_));
  INV   g00674(.A(\priority[85] ), .Y(new_n1060_));
  NOR2  g00675(.A(\req[85] ), .B(new_n1060_), .Y(new_n1061_));
  NOR2  g00676(.A(new_n1061_), .B(\priority[86] ), .Y(new_n1062_));
  NAND2 g00677(.A(new_n1062_), .B(new_n673_), .Y(new_n1063_));
  NOR2  g00678(.A(new_n1063_), .B(new_n1059_), .Y(new_n1064_));
  NAND2 g00679(.A(\req[86] ), .B(new_n673_), .Y(new_n1065_));
  NOR2  g00680(.A(\req[88] ), .B(\req[87] ), .Y(new_n1066_));
  NAND2 g00681(.A(new_n1066_), .B(new_n1065_), .Y(new_n1067_));
  NOR2  g00682(.A(new_n1067_), .B(new_n1064_), .Y(new_n1068_));
  INV   g00683(.A(\priority[88] ), .Y(new_n1069_));
  NOR2  g00684(.A(\req[88] ), .B(new_n1069_), .Y(new_n1070_));
  NOR2  g00685(.A(new_n1070_), .B(\priority[89] ), .Y(new_n1071_));
  NAND2 g00686(.A(new_n1071_), .B(new_n683_), .Y(new_n1072_));
  NOR2  g00687(.A(new_n1072_), .B(new_n1068_), .Y(new_n1073_));
  NAND2 g00688(.A(\req[89] ), .B(new_n683_), .Y(new_n1074_));
  NOR2  g00689(.A(\req[91] ), .B(\req[90] ), .Y(new_n1075_));
  NAND2 g00690(.A(new_n1075_), .B(new_n1074_), .Y(new_n1076_));
  NOR2  g00691(.A(new_n1076_), .B(new_n1073_), .Y(new_n1077_));
  INV   g00692(.A(\priority[91] ), .Y(new_n1078_));
  NOR2  g00693(.A(\req[91] ), .B(new_n1078_), .Y(new_n1079_));
  NOR2  g00694(.A(new_n1079_), .B(\priority[92] ), .Y(new_n1080_));
  NAND2 g00695(.A(new_n1080_), .B(new_n693_), .Y(new_n1081_));
  NOR2  g00696(.A(new_n1081_), .B(new_n1077_), .Y(new_n1082_));
  NAND2 g00697(.A(\req[92] ), .B(new_n693_), .Y(new_n1083_));
  NOR2  g00698(.A(\req[94] ), .B(\req[93] ), .Y(new_n1084_));
  NAND2 g00699(.A(new_n1084_), .B(new_n1083_), .Y(new_n1085_));
  NOR2  g00700(.A(new_n1085_), .B(new_n1082_), .Y(new_n1086_));
  INV   g00701(.A(\priority[94] ), .Y(new_n1087_));
  NOR2  g00702(.A(\req[94] ), .B(new_n1087_), .Y(new_n1088_));
  NOR2  g00703(.A(new_n1088_), .B(\priority[95] ), .Y(new_n1089_));
  NAND2 g00704(.A(new_n1089_), .B(new_n703_), .Y(new_n1090_));
  NOR2  g00705(.A(new_n1090_), .B(new_n1086_), .Y(new_n1091_));
  NAND2 g00706(.A(\req[95] ), .B(new_n703_), .Y(new_n1092_));
  NOR2  g00707(.A(\req[97] ), .B(\req[96] ), .Y(new_n1093_));
  NAND2 g00708(.A(new_n1093_), .B(new_n1092_), .Y(new_n1094_));
  NOR2  g00709(.A(new_n1094_), .B(new_n1091_), .Y(new_n1095_));
  INV   g00710(.A(\priority[97] ), .Y(new_n1096_));
  NOR2  g00711(.A(\req[97] ), .B(new_n1096_), .Y(new_n1097_));
  NOR2  g00712(.A(new_n1097_), .B(\priority[98] ), .Y(new_n1098_));
  NAND2 g00713(.A(new_n1098_), .B(new_n713_), .Y(new_n1099_));
  NOR2  g00714(.A(new_n1099_), .B(new_n1095_), .Y(new_n1100_));
  NAND2 g00715(.A(\req[98] ), .B(new_n713_), .Y(new_n1101_));
  NOR2  g00716(.A(\req[100] ), .B(\req[99] ), .Y(new_n1102_));
  NAND2 g00717(.A(new_n1102_), .B(new_n1101_), .Y(new_n1103_));
  NOR2  g00718(.A(new_n1103_), .B(new_n1100_), .Y(new_n1104_));
  INV   g00719(.A(\priority[100] ), .Y(new_n1105_));
  NOR2  g00720(.A(\req[100] ), .B(new_n1105_), .Y(new_n1106_));
  NOR2  g00721(.A(new_n1106_), .B(\priority[101] ), .Y(new_n1107_));
  NAND2 g00722(.A(new_n1107_), .B(new_n723_), .Y(new_n1108_));
  NOR2  g00723(.A(new_n1108_), .B(new_n1104_), .Y(new_n1109_));
  NAND2 g00724(.A(\req[101] ), .B(new_n723_), .Y(new_n1110_));
  NOR2  g00725(.A(\req[103] ), .B(\req[102] ), .Y(new_n1111_));
  NAND2 g00726(.A(new_n1111_), .B(new_n1110_), .Y(new_n1112_));
  NOR2  g00727(.A(new_n1112_), .B(new_n1109_), .Y(new_n1113_));
  INV   g00728(.A(\priority[103] ), .Y(new_n1114_));
  NOR2  g00729(.A(\req[103] ), .B(new_n1114_), .Y(new_n1115_));
  NOR2  g00730(.A(new_n1115_), .B(\priority[104] ), .Y(new_n1116_));
  NAND2 g00731(.A(new_n1116_), .B(new_n733_), .Y(new_n1117_));
  NOR2  g00732(.A(new_n1117_), .B(new_n1113_), .Y(new_n1118_));
  NAND2 g00733(.A(\req[104] ), .B(new_n733_), .Y(new_n1119_));
  NOR2  g00734(.A(\req[106] ), .B(\req[105] ), .Y(new_n1120_));
  NAND2 g00735(.A(new_n1120_), .B(new_n1119_), .Y(new_n1121_));
  NOR2  g00736(.A(new_n1121_), .B(new_n1118_), .Y(new_n1122_));
  INV   g00737(.A(\priority[106] ), .Y(new_n1123_));
  NOR2  g00738(.A(\req[106] ), .B(new_n1123_), .Y(new_n1124_));
  NOR2  g00739(.A(new_n1124_), .B(\priority[107] ), .Y(new_n1125_));
  NAND2 g00740(.A(new_n1125_), .B(new_n743_), .Y(new_n1126_));
  NOR2  g00741(.A(new_n1126_), .B(new_n1122_), .Y(new_n1127_));
  NAND2 g00742(.A(\req[107] ), .B(new_n743_), .Y(new_n1128_));
  NOR2  g00743(.A(\req[109] ), .B(\req[108] ), .Y(new_n1129_));
  NAND2 g00744(.A(new_n1129_), .B(new_n1128_), .Y(new_n1130_));
  NOR2  g00745(.A(new_n1130_), .B(new_n1127_), .Y(new_n1131_));
  INV   g00746(.A(\priority[109] ), .Y(new_n1132_));
  NOR2  g00747(.A(\req[109] ), .B(new_n1132_), .Y(new_n1133_));
  NOR2  g00748(.A(new_n1133_), .B(\priority[110] ), .Y(new_n1134_));
  NAND2 g00749(.A(new_n1134_), .B(new_n753_), .Y(new_n1135_));
  NOR2  g00750(.A(new_n1135_), .B(new_n1131_), .Y(new_n1136_));
  NAND2 g00751(.A(\req[110] ), .B(new_n753_), .Y(new_n1137_));
  NOR2  g00752(.A(\req[112] ), .B(\req[111] ), .Y(new_n1138_));
  NAND2 g00753(.A(new_n1138_), .B(new_n1137_), .Y(new_n1139_));
  NOR2  g00754(.A(new_n1139_), .B(new_n1136_), .Y(new_n1140_));
  INV   g00755(.A(\priority[112] ), .Y(new_n1141_));
  NOR2  g00756(.A(\req[112] ), .B(new_n1141_), .Y(new_n1142_));
  NOR2  g00757(.A(new_n1142_), .B(\priority[113] ), .Y(new_n1143_));
  NAND2 g00758(.A(new_n1143_), .B(new_n763_), .Y(new_n1144_));
  NOR2  g00759(.A(new_n1144_), .B(new_n1140_), .Y(new_n1145_));
  NAND2 g00760(.A(\req[113] ), .B(new_n763_), .Y(new_n1146_));
  NOR2  g00761(.A(\req[115] ), .B(\req[114] ), .Y(new_n1147_));
  NAND2 g00762(.A(new_n1147_), .B(new_n1146_), .Y(new_n1148_));
  NOR2  g00763(.A(new_n1148_), .B(new_n1145_), .Y(new_n1149_));
  INV   g00764(.A(\priority[115] ), .Y(new_n1150_));
  NOR2  g00765(.A(\req[115] ), .B(new_n1150_), .Y(new_n1151_));
  NOR2  g00766(.A(new_n1151_), .B(\priority[116] ), .Y(new_n1152_));
  NAND2 g00767(.A(new_n1152_), .B(new_n773_), .Y(new_n1153_));
  NOR2  g00768(.A(new_n1153_), .B(new_n1149_), .Y(new_n1154_));
  NAND2 g00769(.A(\req[116] ), .B(new_n773_), .Y(new_n1155_));
  NOR2  g00770(.A(\req[118] ), .B(\req[117] ), .Y(new_n1156_));
  NAND2 g00771(.A(new_n1156_), .B(new_n1155_), .Y(new_n1157_));
  NOR2  g00772(.A(new_n1157_), .B(new_n1154_), .Y(new_n1158_));
  INV   g00773(.A(\priority[118] ), .Y(new_n1159_));
  NOR2  g00774(.A(\req[118] ), .B(new_n1159_), .Y(new_n1160_));
  NOR2  g00775(.A(new_n1160_), .B(\priority[119] ), .Y(new_n1161_));
  NAND2 g00776(.A(new_n1161_), .B(new_n783_), .Y(new_n1162_));
  NOR2  g00777(.A(new_n1162_), .B(new_n1158_), .Y(new_n1163_));
  NAND2 g00778(.A(\req[119] ), .B(new_n783_), .Y(new_n1164_));
  NOR2  g00779(.A(\req[121] ), .B(\req[120] ), .Y(new_n1165_));
  NAND2 g00780(.A(new_n1165_), .B(new_n1164_), .Y(new_n1166_));
  NOR2  g00781(.A(new_n1166_), .B(new_n1163_), .Y(new_n1167_));
  INV   g00782(.A(\priority[121] ), .Y(new_n1168_));
  NOR2  g00783(.A(\req[121] ), .B(new_n1168_), .Y(new_n1169_));
  NOR2  g00784(.A(new_n1169_), .B(\priority[122] ), .Y(new_n1170_));
  NAND2 g00785(.A(new_n1170_), .B(new_n793_), .Y(new_n1171_));
  NOR2  g00786(.A(new_n1171_), .B(new_n1167_), .Y(new_n1172_));
  NAND2 g00787(.A(\req[122] ), .B(new_n793_), .Y(new_n1173_));
  NOR2  g00788(.A(\req[124] ), .B(\req[123] ), .Y(new_n1174_));
  NAND2 g00789(.A(new_n1174_), .B(new_n1173_), .Y(new_n1175_));
  NOR2  g00790(.A(new_n1175_), .B(new_n1172_), .Y(new_n1176_));
  INV   g00791(.A(\priority[124] ), .Y(new_n1177_));
  NOR2  g00792(.A(\req[124] ), .B(new_n1177_), .Y(new_n1178_));
  NOR2  g00793(.A(new_n1178_), .B(\priority[125] ), .Y(new_n1179_));
  NAND2 g00794(.A(new_n1179_), .B(new_n803_), .Y(new_n1180_));
  NOR2  g00795(.A(new_n1180_), .B(new_n1176_), .Y(new_n1181_));
  NAND2 g00796(.A(\req[125] ), .B(new_n803_), .Y(new_n1182_));
  NOR2  g00797(.A(\req[127] ), .B(\req[126] ), .Y(new_n1183_));
  NAND2 g00798(.A(new_n1183_), .B(new_n1182_), .Y(new_n1184_));
  NOR2  g00799(.A(new_n1184_), .B(new_n1181_), .Y(new_n1185_));
  INV   g00800(.A(\priority[127] ), .Y(new_n1186_));
  NOR2  g00801(.A(\req[127] ), .B(new_n1186_), .Y(new_n1187_));
  NOR2  g00802(.A(new_n1187_), .B(\priority[0] ), .Y(new_n1188_));
  NAND2 g00803(.A(new_n1188_), .B(new_n386_), .Y(new_n1189_));
  NOR2  g00804(.A(new_n1189_), .B(new_n1185_), .Y(new_n1190_));
  NAND2 g00805(.A(\req[0] ), .B(new_n386_), .Y(new_n1191_));
  NAND2 g00806(.A(new_n1191_), .B(\req[1] ), .Y(new_n1192_));
  NOR2  g00807(.A(new_n1192_), .B(new_n1190_), .Y(\grant[1] ));
  NOR2  g00808(.A(\req[5] ), .B(\req[4] ), .Y(new_n1194_));
  INV   g00809(.A(new_n1194_), .Y(new_n1195_));
  NOR2  g00810(.A(new_n1195_), .B(new_n395_), .Y(new_n1196_));
  NOR2  g00811(.A(\req[5] ), .B(new_n392_), .Y(new_n1197_));
  NOR2  g00812(.A(new_n1197_), .B(\priority[6] ), .Y(new_n1198_));
  NAND2 g00813(.A(new_n1198_), .B(new_n826_), .Y(new_n1199_));
  NOR2  g00814(.A(new_n1199_), .B(new_n1196_), .Y(new_n1200_));
  NAND2 g00815(.A(\req[6] ), .B(new_n826_), .Y(new_n1201_));
  NOR2  g00816(.A(\req[8] ), .B(\req[7] ), .Y(new_n1202_));
  NAND2 g00817(.A(new_n1202_), .B(new_n1201_), .Y(new_n1203_));
  NOR2  g00818(.A(new_n1203_), .B(new_n1200_), .Y(new_n1204_));
  NOR2  g00819(.A(\req[8] ), .B(new_n402_), .Y(new_n1205_));
  NOR2  g00820(.A(new_n1205_), .B(\priority[9] ), .Y(new_n1206_));
  NAND2 g00821(.A(new_n1206_), .B(new_n835_), .Y(new_n1207_));
  NOR2  g00822(.A(new_n1207_), .B(new_n1204_), .Y(new_n1208_));
  NAND2 g00823(.A(\req[9] ), .B(new_n835_), .Y(new_n1209_));
  NOR2  g00824(.A(\req[11] ), .B(\req[10] ), .Y(new_n1210_));
  NAND2 g00825(.A(new_n1210_), .B(new_n1209_), .Y(new_n1211_));
  NOR2  g00826(.A(new_n1211_), .B(new_n1208_), .Y(new_n1212_));
  NOR2  g00827(.A(\req[11] ), .B(new_n412_), .Y(new_n1213_));
  NOR2  g00828(.A(new_n1213_), .B(\priority[12] ), .Y(new_n1214_));
  NAND2 g00829(.A(new_n1214_), .B(new_n844_), .Y(new_n1215_));
  NOR2  g00830(.A(new_n1215_), .B(new_n1212_), .Y(new_n1216_));
  NAND2 g00831(.A(\req[12] ), .B(new_n844_), .Y(new_n1217_));
  NOR2  g00832(.A(\req[14] ), .B(\req[13] ), .Y(new_n1218_));
  NAND2 g00833(.A(new_n1218_), .B(new_n1217_), .Y(new_n1219_));
  NOR2  g00834(.A(new_n1219_), .B(new_n1216_), .Y(new_n1220_));
  NOR2  g00835(.A(\req[14] ), .B(new_n422_), .Y(new_n1221_));
  NOR2  g00836(.A(new_n1221_), .B(\priority[15] ), .Y(new_n1222_));
  NAND2 g00837(.A(new_n1222_), .B(new_n853_), .Y(new_n1223_));
  NOR2  g00838(.A(new_n1223_), .B(new_n1220_), .Y(new_n1224_));
  NAND2 g00839(.A(\req[15] ), .B(new_n853_), .Y(new_n1225_));
  NOR2  g00840(.A(\req[17] ), .B(\req[16] ), .Y(new_n1226_));
  NAND2 g00841(.A(new_n1226_), .B(new_n1225_), .Y(new_n1227_));
  NOR2  g00842(.A(new_n1227_), .B(new_n1224_), .Y(new_n1228_));
  NOR2  g00843(.A(\req[17] ), .B(new_n432_), .Y(new_n1229_));
  NOR2  g00844(.A(new_n1229_), .B(\priority[18] ), .Y(new_n1230_));
  NAND2 g00845(.A(new_n1230_), .B(new_n862_), .Y(new_n1231_));
  NOR2  g00846(.A(new_n1231_), .B(new_n1228_), .Y(new_n1232_));
  NAND2 g00847(.A(\req[18] ), .B(new_n862_), .Y(new_n1233_));
  NOR2  g00848(.A(\req[20] ), .B(\req[19] ), .Y(new_n1234_));
  NAND2 g00849(.A(new_n1234_), .B(new_n1233_), .Y(new_n1235_));
  NOR2  g00850(.A(new_n1235_), .B(new_n1232_), .Y(new_n1236_));
  NOR2  g00851(.A(\req[20] ), .B(new_n442_), .Y(new_n1237_));
  NOR2  g00852(.A(new_n1237_), .B(\priority[21] ), .Y(new_n1238_));
  NAND2 g00853(.A(new_n1238_), .B(new_n871_), .Y(new_n1239_));
  NOR2  g00854(.A(new_n1239_), .B(new_n1236_), .Y(new_n1240_));
  NAND2 g00855(.A(\req[21] ), .B(new_n871_), .Y(new_n1241_));
  NOR2  g00856(.A(\req[23] ), .B(\req[22] ), .Y(new_n1242_));
  NAND2 g00857(.A(new_n1242_), .B(new_n1241_), .Y(new_n1243_));
  NOR2  g00858(.A(new_n1243_), .B(new_n1240_), .Y(new_n1244_));
  NOR2  g00859(.A(\req[23] ), .B(new_n452_), .Y(new_n1245_));
  NOR2  g00860(.A(new_n1245_), .B(\priority[24] ), .Y(new_n1246_));
  NAND2 g00861(.A(new_n1246_), .B(new_n880_), .Y(new_n1247_));
  NOR2  g00862(.A(new_n1247_), .B(new_n1244_), .Y(new_n1248_));
  NAND2 g00863(.A(\req[24] ), .B(new_n880_), .Y(new_n1249_));
  NOR2  g00864(.A(\req[26] ), .B(\req[25] ), .Y(new_n1250_));
  NAND2 g00865(.A(new_n1250_), .B(new_n1249_), .Y(new_n1251_));
  NOR2  g00866(.A(new_n1251_), .B(new_n1248_), .Y(new_n1252_));
  NOR2  g00867(.A(\req[26] ), .B(new_n462_), .Y(new_n1253_));
  NOR2  g00868(.A(new_n1253_), .B(\priority[27] ), .Y(new_n1254_));
  NAND2 g00869(.A(new_n1254_), .B(new_n889_), .Y(new_n1255_));
  NOR2  g00870(.A(new_n1255_), .B(new_n1252_), .Y(new_n1256_));
  NAND2 g00871(.A(\req[27] ), .B(new_n889_), .Y(new_n1257_));
  NOR2  g00872(.A(\req[29] ), .B(\req[28] ), .Y(new_n1258_));
  NAND2 g00873(.A(new_n1258_), .B(new_n1257_), .Y(new_n1259_));
  NOR2  g00874(.A(new_n1259_), .B(new_n1256_), .Y(new_n1260_));
  NOR2  g00875(.A(\req[29] ), .B(new_n472_), .Y(new_n1261_));
  NOR2  g00876(.A(new_n1261_), .B(\priority[30] ), .Y(new_n1262_));
  NAND2 g00877(.A(new_n1262_), .B(new_n898_), .Y(new_n1263_));
  NOR2  g00878(.A(new_n1263_), .B(new_n1260_), .Y(new_n1264_));
  NAND2 g00879(.A(\req[30] ), .B(new_n898_), .Y(new_n1265_));
  NOR2  g00880(.A(\req[32] ), .B(\req[31] ), .Y(new_n1266_));
  NAND2 g00881(.A(new_n1266_), .B(new_n1265_), .Y(new_n1267_));
  NOR2  g00882(.A(new_n1267_), .B(new_n1264_), .Y(new_n1268_));
  NOR2  g00883(.A(\req[32] ), .B(new_n482_), .Y(new_n1269_));
  NOR2  g00884(.A(new_n1269_), .B(\priority[33] ), .Y(new_n1270_));
  NAND2 g00885(.A(new_n1270_), .B(new_n907_), .Y(new_n1271_));
  NOR2  g00886(.A(new_n1271_), .B(new_n1268_), .Y(new_n1272_));
  NAND2 g00887(.A(\req[33] ), .B(new_n907_), .Y(new_n1273_));
  NOR2  g00888(.A(\req[35] ), .B(\req[34] ), .Y(new_n1274_));
  NAND2 g00889(.A(new_n1274_), .B(new_n1273_), .Y(new_n1275_));
  NOR2  g00890(.A(new_n1275_), .B(new_n1272_), .Y(new_n1276_));
  NOR2  g00891(.A(\req[35] ), .B(new_n492_), .Y(new_n1277_));
  NOR2  g00892(.A(new_n1277_), .B(\priority[36] ), .Y(new_n1278_));
  NAND2 g00893(.A(new_n1278_), .B(new_n916_), .Y(new_n1279_));
  NOR2  g00894(.A(new_n1279_), .B(new_n1276_), .Y(new_n1280_));
  NAND2 g00895(.A(\req[36] ), .B(new_n916_), .Y(new_n1281_));
  NOR2  g00896(.A(\req[38] ), .B(\req[37] ), .Y(new_n1282_));
  NAND2 g00897(.A(new_n1282_), .B(new_n1281_), .Y(new_n1283_));
  NOR2  g00898(.A(new_n1283_), .B(new_n1280_), .Y(new_n1284_));
  NOR2  g00899(.A(\req[38] ), .B(new_n502_), .Y(new_n1285_));
  NOR2  g00900(.A(new_n1285_), .B(\priority[39] ), .Y(new_n1286_));
  NAND2 g00901(.A(new_n1286_), .B(new_n925_), .Y(new_n1287_));
  NOR2  g00902(.A(new_n1287_), .B(new_n1284_), .Y(new_n1288_));
  NAND2 g00903(.A(\req[39] ), .B(new_n925_), .Y(new_n1289_));
  NOR2  g00904(.A(\req[41] ), .B(\req[40] ), .Y(new_n1290_));
  NAND2 g00905(.A(new_n1290_), .B(new_n1289_), .Y(new_n1291_));
  NOR2  g00906(.A(new_n1291_), .B(new_n1288_), .Y(new_n1292_));
  NOR2  g00907(.A(\req[41] ), .B(new_n512_), .Y(new_n1293_));
  NOR2  g00908(.A(new_n1293_), .B(\priority[42] ), .Y(new_n1294_));
  NAND2 g00909(.A(new_n1294_), .B(new_n934_), .Y(new_n1295_));
  NOR2  g00910(.A(new_n1295_), .B(new_n1292_), .Y(new_n1296_));
  NAND2 g00911(.A(\req[42] ), .B(new_n934_), .Y(new_n1297_));
  NOR2  g00912(.A(\req[44] ), .B(\req[43] ), .Y(new_n1298_));
  NAND2 g00913(.A(new_n1298_), .B(new_n1297_), .Y(new_n1299_));
  NOR2  g00914(.A(new_n1299_), .B(new_n1296_), .Y(new_n1300_));
  NOR2  g00915(.A(\req[44] ), .B(new_n522_), .Y(new_n1301_));
  NOR2  g00916(.A(new_n1301_), .B(\priority[45] ), .Y(new_n1302_));
  NAND2 g00917(.A(new_n1302_), .B(new_n943_), .Y(new_n1303_));
  NOR2  g00918(.A(new_n1303_), .B(new_n1300_), .Y(new_n1304_));
  NAND2 g00919(.A(\req[45] ), .B(new_n943_), .Y(new_n1305_));
  NOR2  g00920(.A(\req[47] ), .B(\req[46] ), .Y(new_n1306_));
  NAND2 g00921(.A(new_n1306_), .B(new_n1305_), .Y(new_n1307_));
  NOR2  g00922(.A(new_n1307_), .B(new_n1304_), .Y(new_n1308_));
  NOR2  g00923(.A(\req[47] ), .B(new_n532_), .Y(new_n1309_));
  NOR2  g00924(.A(new_n1309_), .B(\priority[48] ), .Y(new_n1310_));
  NAND2 g00925(.A(new_n1310_), .B(new_n952_), .Y(new_n1311_));
  NOR2  g00926(.A(new_n1311_), .B(new_n1308_), .Y(new_n1312_));
  NAND2 g00927(.A(\req[48] ), .B(new_n952_), .Y(new_n1313_));
  NOR2  g00928(.A(\req[50] ), .B(\req[49] ), .Y(new_n1314_));
  NAND2 g00929(.A(new_n1314_), .B(new_n1313_), .Y(new_n1315_));
  NOR2  g00930(.A(new_n1315_), .B(new_n1312_), .Y(new_n1316_));
  NOR2  g00931(.A(\req[50] ), .B(new_n542_), .Y(new_n1317_));
  NOR2  g00932(.A(new_n1317_), .B(\priority[51] ), .Y(new_n1318_));
  NAND2 g00933(.A(new_n1318_), .B(new_n961_), .Y(new_n1319_));
  NOR2  g00934(.A(new_n1319_), .B(new_n1316_), .Y(new_n1320_));
  NAND2 g00935(.A(\req[51] ), .B(new_n961_), .Y(new_n1321_));
  NOR2  g00936(.A(\req[53] ), .B(\req[52] ), .Y(new_n1322_));
  NAND2 g00937(.A(new_n1322_), .B(new_n1321_), .Y(new_n1323_));
  NOR2  g00938(.A(new_n1323_), .B(new_n1320_), .Y(new_n1324_));
  NOR2  g00939(.A(\req[53] ), .B(new_n552_), .Y(new_n1325_));
  NOR2  g00940(.A(new_n1325_), .B(\priority[54] ), .Y(new_n1326_));
  NAND2 g00941(.A(new_n1326_), .B(new_n970_), .Y(new_n1327_));
  NOR2  g00942(.A(new_n1327_), .B(new_n1324_), .Y(new_n1328_));
  NAND2 g00943(.A(\req[54] ), .B(new_n970_), .Y(new_n1329_));
  NOR2  g00944(.A(\req[56] ), .B(\req[55] ), .Y(new_n1330_));
  NAND2 g00945(.A(new_n1330_), .B(new_n1329_), .Y(new_n1331_));
  NOR2  g00946(.A(new_n1331_), .B(new_n1328_), .Y(new_n1332_));
  NOR2  g00947(.A(\req[56] ), .B(new_n562_), .Y(new_n1333_));
  NOR2  g00948(.A(new_n1333_), .B(\priority[57] ), .Y(new_n1334_));
  NAND2 g00949(.A(new_n1334_), .B(new_n979_), .Y(new_n1335_));
  NOR2  g00950(.A(new_n1335_), .B(new_n1332_), .Y(new_n1336_));
  NAND2 g00951(.A(\req[57] ), .B(new_n979_), .Y(new_n1337_));
  NOR2  g00952(.A(\req[59] ), .B(\req[58] ), .Y(new_n1338_));
  NAND2 g00953(.A(new_n1338_), .B(new_n1337_), .Y(new_n1339_));
  NOR2  g00954(.A(new_n1339_), .B(new_n1336_), .Y(new_n1340_));
  NOR2  g00955(.A(\req[59] ), .B(new_n572_), .Y(new_n1341_));
  NOR2  g00956(.A(new_n1341_), .B(\priority[60] ), .Y(new_n1342_));
  NAND2 g00957(.A(new_n1342_), .B(new_n988_), .Y(new_n1343_));
  NOR2  g00958(.A(new_n1343_), .B(new_n1340_), .Y(new_n1344_));
  NAND2 g00959(.A(\req[60] ), .B(new_n988_), .Y(new_n1345_));
  NOR2  g00960(.A(\req[62] ), .B(\req[61] ), .Y(new_n1346_));
  NAND2 g00961(.A(new_n1346_), .B(new_n1345_), .Y(new_n1347_));
  NOR2  g00962(.A(new_n1347_), .B(new_n1344_), .Y(new_n1348_));
  NOR2  g00963(.A(\req[62] ), .B(new_n582_), .Y(new_n1349_));
  NOR2  g00964(.A(new_n1349_), .B(\priority[63] ), .Y(new_n1350_));
  NAND2 g00965(.A(new_n1350_), .B(new_n997_), .Y(new_n1351_));
  NOR2  g00966(.A(new_n1351_), .B(new_n1348_), .Y(new_n1352_));
  NAND2 g00967(.A(\req[63] ), .B(new_n997_), .Y(new_n1353_));
  NOR2  g00968(.A(\req[65] ), .B(\req[64] ), .Y(new_n1354_));
  NAND2 g00969(.A(new_n1354_), .B(new_n1353_), .Y(new_n1355_));
  NOR2  g00970(.A(new_n1355_), .B(new_n1352_), .Y(new_n1356_));
  NOR2  g00971(.A(\req[65] ), .B(new_n592_), .Y(new_n1357_));
  NOR2  g00972(.A(new_n1357_), .B(\priority[66] ), .Y(new_n1358_));
  NAND2 g00973(.A(new_n1358_), .B(new_n1006_), .Y(new_n1359_));
  NOR2  g00974(.A(new_n1359_), .B(new_n1356_), .Y(new_n1360_));
  NAND2 g00975(.A(\req[66] ), .B(new_n1006_), .Y(new_n1361_));
  NOR2  g00976(.A(\req[68] ), .B(\req[67] ), .Y(new_n1362_));
  NAND2 g00977(.A(new_n1362_), .B(new_n1361_), .Y(new_n1363_));
  NOR2  g00978(.A(new_n1363_), .B(new_n1360_), .Y(new_n1364_));
  NOR2  g00979(.A(\req[68] ), .B(new_n602_), .Y(new_n1365_));
  NOR2  g00980(.A(new_n1365_), .B(\priority[69] ), .Y(new_n1366_));
  NAND2 g00981(.A(new_n1366_), .B(new_n1015_), .Y(new_n1367_));
  NOR2  g00982(.A(new_n1367_), .B(new_n1364_), .Y(new_n1368_));
  NAND2 g00983(.A(\req[69] ), .B(new_n1015_), .Y(new_n1369_));
  NOR2  g00984(.A(\req[71] ), .B(\req[70] ), .Y(new_n1370_));
  NAND2 g00985(.A(new_n1370_), .B(new_n1369_), .Y(new_n1371_));
  NOR2  g00986(.A(new_n1371_), .B(new_n1368_), .Y(new_n1372_));
  NOR2  g00987(.A(\req[71] ), .B(new_n612_), .Y(new_n1373_));
  NOR2  g00988(.A(new_n1373_), .B(\priority[72] ), .Y(new_n1374_));
  NAND2 g00989(.A(new_n1374_), .B(new_n1024_), .Y(new_n1375_));
  NOR2  g00990(.A(new_n1375_), .B(new_n1372_), .Y(new_n1376_));
  NAND2 g00991(.A(\req[72] ), .B(new_n1024_), .Y(new_n1377_));
  NOR2  g00992(.A(\req[74] ), .B(\req[73] ), .Y(new_n1378_));
  NAND2 g00993(.A(new_n1378_), .B(new_n1377_), .Y(new_n1379_));
  NOR2  g00994(.A(new_n1379_), .B(new_n1376_), .Y(new_n1380_));
  NOR2  g00995(.A(\req[74] ), .B(new_n622_), .Y(new_n1381_));
  NOR2  g00996(.A(new_n1381_), .B(\priority[75] ), .Y(new_n1382_));
  NAND2 g00997(.A(new_n1382_), .B(new_n1033_), .Y(new_n1383_));
  NOR2  g00998(.A(new_n1383_), .B(new_n1380_), .Y(new_n1384_));
  NAND2 g00999(.A(\req[75] ), .B(new_n1033_), .Y(new_n1385_));
  NOR2  g01000(.A(\req[77] ), .B(\req[76] ), .Y(new_n1386_));
  NAND2 g01001(.A(new_n1386_), .B(new_n1385_), .Y(new_n1387_));
  NOR2  g01002(.A(new_n1387_), .B(new_n1384_), .Y(new_n1388_));
  NOR2  g01003(.A(\req[77] ), .B(new_n632_), .Y(new_n1389_));
  NOR2  g01004(.A(new_n1389_), .B(\priority[78] ), .Y(new_n1390_));
  NAND2 g01005(.A(new_n1390_), .B(new_n1042_), .Y(new_n1391_));
  NOR2  g01006(.A(new_n1391_), .B(new_n1388_), .Y(new_n1392_));
  NAND2 g01007(.A(\req[78] ), .B(new_n1042_), .Y(new_n1393_));
  NOR2  g01008(.A(\req[80] ), .B(\req[79] ), .Y(new_n1394_));
  NAND2 g01009(.A(new_n1394_), .B(new_n1393_), .Y(new_n1395_));
  NOR2  g01010(.A(new_n1395_), .B(new_n1392_), .Y(new_n1396_));
  NOR2  g01011(.A(\req[80] ), .B(new_n642_), .Y(new_n1397_));
  NOR2  g01012(.A(new_n1397_), .B(\priority[81] ), .Y(new_n1398_));
  NAND2 g01013(.A(new_n1398_), .B(new_n1051_), .Y(new_n1399_));
  NOR2  g01014(.A(new_n1399_), .B(new_n1396_), .Y(new_n1400_));
  NAND2 g01015(.A(\req[81] ), .B(new_n1051_), .Y(new_n1401_));
  NOR2  g01016(.A(\req[83] ), .B(\req[82] ), .Y(new_n1402_));
  NAND2 g01017(.A(new_n1402_), .B(new_n1401_), .Y(new_n1403_));
  NOR2  g01018(.A(new_n1403_), .B(new_n1400_), .Y(new_n1404_));
  NOR2  g01019(.A(\req[83] ), .B(new_n652_), .Y(new_n1405_));
  NOR2  g01020(.A(new_n1405_), .B(\priority[84] ), .Y(new_n1406_));
  NAND2 g01021(.A(new_n1406_), .B(new_n1060_), .Y(new_n1407_));
  NOR2  g01022(.A(new_n1407_), .B(new_n1404_), .Y(new_n1408_));
  NAND2 g01023(.A(\req[84] ), .B(new_n1060_), .Y(new_n1409_));
  NOR2  g01024(.A(\req[86] ), .B(\req[85] ), .Y(new_n1410_));
  NAND2 g01025(.A(new_n1410_), .B(new_n1409_), .Y(new_n1411_));
  NOR2  g01026(.A(new_n1411_), .B(new_n1408_), .Y(new_n1412_));
  NOR2  g01027(.A(\req[86] ), .B(new_n662_), .Y(new_n1413_));
  NOR2  g01028(.A(new_n1413_), .B(\priority[87] ), .Y(new_n1414_));
  NAND2 g01029(.A(new_n1414_), .B(new_n1069_), .Y(new_n1415_));
  NOR2  g01030(.A(new_n1415_), .B(new_n1412_), .Y(new_n1416_));
  NAND2 g01031(.A(\req[87] ), .B(new_n1069_), .Y(new_n1417_));
  NOR2  g01032(.A(\req[89] ), .B(\req[88] ), .Y(new_n1418_));
  NAND2 g01033(.A(new_n1418_), .B(new_n1417_), .Y(new_n1419_));
  NOR2  g01034(.A(new_n1419_), .B(new_n1416_), .Y(new_n1420_));
  NOR2  g01035(.A(\req[89] ), .B(new_n672_), .Y(new_n1421_));
  NOR2  g01036(.A(new_n1421_), .B(\priority[90] ), .Y(new_n1422_));
  NAND2 g01037(.A(new_n1422_), .B(new_n1078_), .Y(new_n1423_));
  NOR2  g01038(.A(new_n1423_), .B(new_n1420_), .Y(new_n1424_));
  NAND2 g01039(.A(\req[90] ), .B(new_n1078_), .Y(new_n1425_));
  NOR2  g01040(.A(\req[92] ), .B(\req[91] ), .Y(new_n1426_));
  NAND2 g01041(.A(new_n1426_), .B(new_n1425_), .Y(new_n1427_));
  NOR2  g01042(.A(new_n1427_), .B(new_n1424_), .Y(new_n1428_));
  NOR2  g01043(.A(\req[92] ), .B(new_n682_), .Y(new_n1429_));
  NOR2  g01044(.A(new_n1429_), .B(\priority[93] ), .Y(new_n1430_));
  NAND2 g01045(.A(new_n1430_), .B(new_n1087_), .Y(new_n1431_));
  NOR2  g01046(.A(new_n1431_), .B(new_n1428_), .Y(new_n1432_));
  NAND2 g01047(.A(\req[93] ), .B(new_n1087_), .Y(new_n1433_));
  NOR2  g01048(.A(\req[95] ), .B(\req[94] ), .Y(new_n1434_));
  NAND2 g01049(.A(new_n1434_), .B(new_n1433_), .Y(new_n1435_));
  NOR2  g01050(.A(new_n1435_), .B(new_n1432_), .Y(new_n1436_));
  NOR2  g01051(.A(\req[95] ), .B(new_n692_), .Y(new_n1437_));
  NOR2  g01052(.A(new_n1437_), .B(\priority[96] ), .Y(new_n1438_));
  NAND2 g01053(.A(new_n1438_), .B(new_n1096_), .Y(new_n1439_));
  NOR2  g01054(.A(new_n1439_), .B(new_n1436_), .Y(new_n1440_));
  NAND2 g01055(.A(\req[96] ), .B(new_n1096_), .Y(new_n1441_));
  NOR2  g01056(.A(\req[98] ), .B(\req[97] ), .Y(new_n1442_));
  NAND2 g01057(.A(new_n1442_), .B(new_n1441_), .Y(new_n1443_));
  NOR2  g01058(.A(new_n1443_), .B(new_n1440_), .Y(new_n1444_));
  NOR2  g01059(.A(\req[98] ), .B(new_n702_), .Y(new_n1445_));
  NOR2  g01060(.A(new_n1445_), .B(\priority[99] ), .Y(new_n1446_));
  NAND2 g01061(.A(new_n1446_), .B(new_n1105_), .Y(new_n1447_));
  NOR2  g01062(.A(new_n1447_), .B(new_n1444_), .Y(new_n1448_));
  NAND2 g01063(.A(\req[99] ), .B(new_n1105_), .Y(new_n1449_));
  NOR2  g01064(.A(\req[101] ), .B(\req[100] ), .Y(new_n1450_));
  NAND2 g01065(.A(new_n1450_), .B(new_n1449_), .Y(new_n1451_));
  NOR2  g01066(.A(new_n1451_), .B(new_n1448_), .Y(new_n1452_));
  NOR2  g01067(.A(\req[101] ), .B(new_n712_), .Y(new_n1453_));
  NOR2  g01068(.A(new_n1453_), .B(\priority[102] ), .Y(new_n1454_));
  NAND2 g01069(.A(new_n1454_), .B(new_n1114_), .Y(new_n1455_));
  NOR2  g01070(.A(new_n1455_), .B(new_n1452_), .Y(new_n1456_));
  NAND2 g01071(.A(\req[102] ), .B(new_n1114_), .Y(new_n1457_));
  NOR2  g01072(.A(\req[104] ), .B(\req[103] ), .Y(new_n1458_));
  NAND2 g01073(.A(new_n1458_), .B(new_n1457_), .Y(new_n1459_));
  NOR2  g01074(.A(new_n1459_), .B(new_n1456_), .Y(new_n1460_));
  NOR2  g01075(.A(\req[104] ), .B(new_n722_), .Y(new_n1461_));
  NOR2  g01076(.A(new_n1461_), .B(\priority[105] ), .Y(new_n1462_));
  NAND2 g01077(.A(new_n1462_), .B(new_n1123_), .Y(new_n1463_));
  NOR2  g01078(.A(new_n1463_), .B(new_n1460_), .Y(new_n1464_));
  NAND2 g01079(.A(\req[105] ), .B(new_n1123_), .Y(new_n1465_));
  NOR2  g01080(.A(\req[107] ), .B(\req[106] ), .Y(new_n1466_));
  NAND2 g01081(.A(new_n1466_), .B(new_n1465_), .Y(new_n1467_));
  NOR2  g01082(.A(new_n1467_), .B(new_n1464_), .Y(new_n1468_));
  NOR2  g01083(.A(\req[107] ), .B(new_n732_), .Y(new_n1469_));
  NOR2  g01084(.A(new_n1469_), .B(\priority[108] ), .Y(new_n1470_));
  NAND2 g01085(.A(new_n1470_), .B(new_n1132_), .Y(new_n1471_));
  NOR2  g01086(.A(new_n1471_), .B(new_n1468_), .Y(new_n1472_));
  NAND2 g01087(.A(\req[108] ), .B(new_n1132_), .Y(new_n1473_));
  NOR2  g01088(.A(\req[110] ), .B(\req[109] ), .Y(new_n1474_));
  NAND2 g01089(.A(new_n1474_), .B(new_n1473_), .Y(new_n1475_));
  NOR2  g01090(.A(new_n1475_), .B(new_n1472_), .Y(new_n1476_));
  NOR2  g01091(.A(\req[110] ), .B(new_n742_), .Y(new_n1477_));
  NOR2  g01092(.A(new_n1477_), .B(\priority[111] ), .Y(new_n1478_));
  NAND2 g01093(.A(new_n1478_), .B(new_n1141_), .Y(new_n1479_));
  NOR2  g01094(.A(new_n1479_), .B(new_n1476_), .Y(new_n1480_));
  NAND2 g01095(.A(\req[111] ), .B(new_n1141_), .Y(new_n1481_));
  NOR2  g01096(.A(\req[113] ), .B(\req[112] ), .Y(new_n1482_));
  NAND2 g01097(.A(new_n1482_), .B(new_n1481_), .Y(new_n1483_));
  NOR2  g01098(.A(new_n1483_), .B(new_n1480_), .Y(new_n1484_));
  NOR2  g01099(.A(\req[113] ), .B(new_n752_), .Y(new_n1485_));
  NOR2  g01100(.A(new_n1485_), .B(\priority[114] ), .Y(new_n1486_));
  NAND2 g01101(.A(new_n1486_), .B(new_n1150_), .Y(new_n1487_));
  NOR2  g01102(.A(new_n1487_), .B(new_n1484_), .Y(new_n1488_));
  NAND2 g01103(.A(\req[114] ), .B(new_n1150_), .Y(new_n1489_));
  NOR2  g01104(.A(\req[116] ), .B(\req[115] ), .Y(new_n1490_));
  NAND2 g01105(.A(new_n1490_), .B(new_n1489_), .Y(new_n1491_));
  NOR2  g01106(.A(new_n1491_), .B(new_n1488_), .Y(new_n1492_));
  NOR2  g01107(.A(\req[116] ), .B(new_n762_), .Y(new_n1493_));
  NOR2  g01108(.A(new_n1493_), .B(\priority[117] ), .Y(new_n1494_));
  NAND2 g01109(.A(new_n1494_), .B(new_n1159_), .Y(new_n1495_));
  NOR2  g01110(.A(new_n1495_), .B(new_n1492_), .Y(new_n1496_));
  NAND2 g01111(.A(\req[117] ), .B(new_n1159_), .Y(new_n1497_));
  NOR2  g01112(.A(\req[119] ), .B(\req[118] ), .Y(new_n1498_));
  NAND2 g01113(.A(new_n1498_), .B(new_n1497_), .Y(new_n1499_));
  NOR2  g01114(.A(new_n1499_), .B(new_n1496_), .Y(new_n1500_));
  NOR2  g01115(.A(\req[119] ), .B(new_n772_), .Y(new_n1501_));
  NOR2  g01116(.A(new_n1501_), .B(\priority[120] ), .Y(new_n1502_));
  NAND2 g01117(.A(new_n1502_), .B(new_n1168_), .Y(new_n1503_));
  NOR2  g01118(.A(new_n1503_), .B(new_n1500_), .Y(new_n1504_));
  NAND2 g01119(.A(\req[120] ), .B(new_n1168_), .Y(new_n1505_));
  NOR2  g01120(.A(\req[122] ), .B(\req[121] ), .Y(new_n1506_));
  NAND2 g01121(.A(new_n1506_), .B(new_n1505_), .Y(new_n1507_));
  NOR2  g01122(.A(new_n1507_), .B(new_n1504_), .Y(new_n1508_));
  NOR2  g01123(.A(\req[122] ), .B(new_n782_), .Y(new_n1509_));
  NOR2  g01124(.A(new_n1509_), .B(\priority[123] ), .Y(new_n1510_));
  NAND2 g01125(.A(new_n1510_), .B(new_n1177_), .Y(new_n1511_));
  NOR2  g01126(.A(new_n1511_), .B(new_n1508_), .Y(new_n1512_));
  NAND2 g01127(.A(\req[123] ), .B(new_n1177_), .Y(new_n1513_));
  NOR2  g01128(.A(\req[125] ), .B(\req[124] ), .Y(new_n1514_));
  NAND2 g01129(.A(new_n1514_), .B(new_n1513_), .Y(new_n1515_));
  NOR2  g01130(.A(new_n1515_), .B(new_n1512_), .Y(new_n1516_));
  NOR2  g01131(.A(\req[125] ), .B(new_n792_), .Y(new_n1517_));
  NOR2  g01132(.A(new_n1517_), .B(\priority[126] ), .Y(new_n1518_));
  NAND2 g01133(.A(new_n1518_), .B(new_n1186_), .Y(new_n1519_));
  NOR2  g01134(.A(new_n1519_), .B(new_n1516_), .Y(new_n1520_));
  NAND2 g01135(.A(\req[126] ), .B(new_n1186_), .Y(new_n1521_));
  NOR2  g01136(.A(\req[127] ), .B(\req[0] ), .Y(new_n1522_));
  NAND2 g01137(.A(new_n1522_), .B(new_n1521_), .Y(new_n1523_));
  NOR2  g01138(.A(new_n1523_), .B(new_n1520_), .Y(new_n1524_));
  NOR2  g01139(.A(\req[0] ), .B(new_n802_), .Y(new_n1525_));
  NOR2  g01140(.A(new_n1525_), .B(\priority[1] ), .Y(new_n1526_));
  NAND2 g01141(.A(new_n1526_), .B(new_n811_), .Y(new_n1527_));
  NOR2  g01142(.A(new_n1527_), .B(new_n1524_), .Y(new_n1528_));
  NAND2 g01143(.A(\req[1] ), .B(new_n811_), .Y(new_n1529_));
  NAND2 g01144(.A(new_n1529_), .B(\req[2] ), .Y(new_n1530_));
  NOR2  g01145(.A(new_n1530_), .B(new_n1528_), .Y(\grant[2] ));
  INV   g01146(.A(new_n399_), .Y(new_n1532_));
  NOR2  g01147(.A(new_n819_), .B(new_n1532_), .Y(new_n1533_));
  NOR2  g01148(.A(new_n1533_), .B(new_n406_), .Y(new_n1534_));
  NOR2  g01149(.A(new_n1534_), .B(new_n410_), .Y(new_n1535_));
  NOR2  g01150(.A(new_n1535_), .B(new_n416_), .Y(new_n1536_));
  NOR2  g01151(.A(new_n1536_), .B(new_n420_), .Y(new_n1537_));
  NOR2  g01152(.A(new_n1537_), .B(new_n426_), .Y(new_n1538_));
  NOR2  g01153(.A(new_n1538_), .B(new_n430_), .Y(new_n1539_));
  NOR2  g01154(.A(new_n1539_), .B(new_n436_), .Y(new_n1540_));
  NOR2  g01155(.A(new_n1540_), .B(new_n440_), .Y(new_n1541_));
  NOR2  g01156(.A(new_n1541_), .B(new_n446_), .Y(new_n1542_));
  NOR2  g01157(.A(new_n1542_), .B(new_n450_), .Y(new_n1543_));
  NOR2  g01158(.A(new_n1543_), .B(new_n456_), .Y(new_n1544_));
  NOR2  g01159(.A(new_n1544_), .B(new_n460_), .Y(new_n1545_));
  NOR2  g01160(.A(new_n1545_), .B(new_n466_), .Y(new_n1546_));
  NOR2  g01161(.A(new_n1546_), .B(new_n470_), .Y(new_n1547_));
  NOR2  g01162(.A(new_n1547_), .B(new_n476_), .Y(new_n1548_));
  NOR2  g01163(.A(new_n1548_), .B(new_n480_), .Y(new_n1549_));
  NOR2  g01164(.A(new_n1549_), .B(new_n486_), .Y(new_n1550_));
  NOR2  g01165(.A(new_n1550_), .B(new_n490_), .Y(new_n1551_));
  NOR2  g01166(.A(new_n1551_), .B(new_n496_), .Y(new_n1552_));
  NOR2  g01167(.A(new_n1552_), .B(new_n500_), .Y(new_n1553_));
  NOR2  g01168(.A(new_n1553_), .B(new_n506_), .Y(new_n1554_));
  NOR2  g01169(.A(new_n1554_), .B(new_n510_), .Y(new_n1555_));
  NOR2  g01170(.A(new_n1555_), .B(new_n516_), .Y(new_n1556_));
  NOR2  g01171(.A(new_n1556_), .B(new_n520_), .Y(new_n1557_));
  NOR2  g01172(.A(new_n1557_), .B(new_n526_), .Y(new_n1558_));
  NOR2  g01173(.A(new_n1558_), .B(new_n530_), .Y(new_n1559_));
  NOR2  g01174(.A(new_n1559_), .B(new_n536_), .Y(new_n1560_));
  NOR2  g01175(.A(new_n1560_), .B(new_n540_), .Y(new_n1561_));
  NOR2  g01176(.A(new_n1561_), .B(new_n546_), .Y(new_n1562_));
  NOR2  g01177(.A(new_n1562_), .B(new_n550_), .Y(new_n1563_));
  NOR2  g01178(.A(new_n1563_), .B(new_n556_), .Y(new_n1564_));
  NOR2  g01179(.A(new_n1564_), .B(new_n560_), .Y(new_n1565_));
  NOR2  g01180(.A(new_n1565_), .B(new_n566_), .Y(new_n1566_));
  NOR2  g01181(.A(new_n1566_), .B(new_n570_), .Y(new_n1567_));
  NOR2  g01182(.A(new_n1567_), .B(new_n576_), .Y(new_n1568_));
  NOR2  g01183(.A(new_n1568_), .B(new_n580_), .Y(new_n1569_));
  NOR2  g01184(.A(new_n1569_), .B(new_n586_), .Y(new_n1570_));
  NOR2  g01185(.A(new_n1570_), .B(new_n590_), .Y(new_n1571_));
  NOR2  g01186(.A(new_n1571_), .B(new_n596_), .Y(new_n1572_));
  NOR2  g01187(.A(new_n1572_), .B(new_n600_), .Y(new_n1573_));
  NOR2  g01188(.A(new_n1573_), .B(new_n606_), .Y(new_n1574_));
  NOR2  g01189(.A(new_n1574_), .B(new_n610_), .Y(new_n1575_));
  NOR2  g01190(.A(new_n1575_), .B(new_n616_), .Y(new_n1576_));
  NOR2  g01191(.A(new_n1576_), .B(new_n620_), .Y(new_n1577_));
  NOR2  g01192(.A(new_n1577_), .B(new_n626_), .Y(new_n1578_));
  NOR2  g01193(.A(new_n1578_), .B(new_n630_), .Y(new_n1579_));
  NOR2  g01194(.A(new_n1579_), .B(new_n636_), .Y(new_n1580_));
  NOR2  g01195(.A(new_n1580_), .B(new_n640_), .Y(new_n1581_));
  NOR2  g01196(.A(new_n1581_), .B(new_n646_), .Y(new_n1582_));
  NOR2  g01197(.A(new_n1582_), .B(new_n650_), .Y(new_n1583_));
  NOR2  g01198(.A(new_n1583_), .B(new_n656_), .Y(new_n1584_));
  NOR2  g01199(.A(new_n1584_), .B(new_n660_), .Y(new_n1585_));
  NOR2  g01200(.A(new_n1585_), .B(new_n666_), .Y(new_n1586_));
  NOR2  g01201(.A(new_n1586_), .B(new_n670_), .Y(new_n1587_));
  NOR2  g01202(.A(new_n1587_), .B(new_n676_), .Y(new_n1588_));
  NOR2  g01203(.A(new_n1588_), .B(new_n680_), .Y(new_n1589_));
  NOR2  g01204(.A(new_n1589_), .B(new_n686_), .Y(new_n1590_));
  NOR2  g01205(.A(new_n1590_), .B(new_n690_), .Y(new_n1591_));
  NOR2  g01206(.A(new_n1591_), .B(new_n696_), .Y(new_n1592_));
  NOR2  g01207(.A(new_n1592_), .B(new_n700_), .Y(new_n1593_));
  NOR2  g01208(.A(new_n1593_), .B(new_n706_), .Y(new_n1594_));
  NOR2  g01209(.A(new_n1594_), .B(new_n710_), .Y(new_n1595_));
  NOR2  g01210(.A(new_n1595_), .B(new_n716_), .Y(new_n1596_));
  NOR2  g01211(.A(new_n1596_), .B(new_n720_), .Y(new_n1597_));
  NOR2  g01212(.A(new_n1597_), .B(new_n726_), .Y(new_n1598_));
  NOR2  g01213(.A(new_n1598_), .B(new_n730_), .Y(new_n1599_));
  NOR2  g01214(.A(new_n1599_), .B(new_n736_), .Y(new_n1600_));
  NOR2  g01215(.A(new_n1600_), .B(new_n740_), .Y(new_n1601_));
  NOR2  g01216(.A(new_n1601_), .B(new_n746_), .Y(new_n1602_));
  NOR2  g01217(.A(new_n1602_), .B(new_n750_), .Y(new_n1603_));
  NOR2  g01218(.A(new_n1603_), .B(new_n756_), .Y(new_n1604_));
  NOR2  g01219(.A(new_n1604_), .B(new_n760_), .Y(new_n1605_));
  NOR2  g01220(.A(new_n1605_), .B(new_n766_), .Y(new_n1606_));
  NOR2  g01221(.A(new_n1606_), .B(new_n770_), .Y(new_n1607_));
  NOR2  g01222(.A(new_n1607_), .B(new_n776_), .Y(new_n1608_));
  NOR2  g01223(.A(new_n1608_), .B(new_n780_), .Y(new_n1609_));
  NOR2  g01224(.A(new_n1609_), .B(new_n786_), .Y(new_n1610_));
  NOR2  g01225(.A(new_n1610_), .B(new_n790_), .Y(new_n1611_));
  NOR2  g01226(.A(new_n1611_), .B(new_n796_), .Y(new_n1612_));
  NOR2  g01227(.A(new_n1612_), .B(new_n800_), .Y(new_n1613_));
  NOR2  g01228(.A(new_n1613_), .B(new_n806_), .Y(new_n1614_));
  NOR2  g01229(.A(\req[1] ), .B(\req[0] ), .Y(new_n1615_));
  NAND2 g01230(.A(new_n1615_), .B(new_n808_), .Y(new_n1616_));
  NOR2  g01231(.A(new_n1616_), .B(new_n1614_), .Y(new_n1617_));
  NAND2 g01232(.A(new_n388_), .B(new_n393_), .Y(new_n1618_));
  NOR2  g01233(.A(new_n1618_), .B(new_n1617_), .Y(new_n1619_));
  NAND2 g01234(.A(\req[2] ), .B(new_n393_), .Y(new_n1620_));
  NAND2 g01235(.A(new_n1620_), .B(\req[3] ), .Y(new_n1621_));
  NOR2  g01236(.A(new_n1621_), .B(new_n1619_), .Y(\grant[3] ));
  INV   g01237(.A(new_n823_), .Y(new_n1623_));
  NOR2  g01238(.A(new_n1198_), .B(new_n1623_), .Y(new_n1624_));
  NOR2  g01239(.A(new_n1624_), .B(new_n829_), .Y(new_n1625_));
  NOR2  g01240(.A(new_n1625_), .B(new_n833_), .Y(new_n1626_));
  NOR2  g01241(.A(new_n1626_), .B(new_n838_), .Y(new_n1627_));
  NOR2  g01242(.A(new_n1627_), .B(new_n842_), .Y(new_n1628_));
  NOR2  g01243(.A(new_n1628_), .B(new_n847_), .Y(new_n1629_));
  NOR2  g01244(.A(new_n1629_), .B(new_n851_), .Y(new_n1630_));
  NOR2  g01245(.A(new_n1630_), .B(new_n856_), .Y(new_n1631_));
  NOR2  g01246(.A(new_n1631_), .B(new_n860_), .Y(new_n1632_));
  NOR2  g01247(.A(new_n1632_), .B(new_n865_), .Y(new_n1633_));
  NOR2  g01248(.A(new_n1633_), .B(new_n869_), .Y(new_n1634_));
  NOR2  g01249(.A(new_n1634_), .B(new_n874_), .Y(new_n1635_));
  NOR2  g01250(.A(new_n1635_), .B(new_n878_), .Y(new_n1636_));
  NOR2  g01251(.A(new_n1636_), .B(new_n883_), .Y(new_n1637_));
  NOR2  g01252(.A(new_n1637_), .B(new_n887_), .Y(new_n1638_));
  NOR2  g01253(.A(new_n1638_), .B(new_n892_), .Y(new_n1639_));
  NOR2  g01254(.A(new_n1639_), .B(new_n896_), .Y(new_n1640_));
  NOR2  g01255(.A(new_n1640_), .B(new_n901_), .Y(new_n1641_));
  NOR2  g01256(.A(new_n1641_), .B(new_n905_), .Y(new_n1642_));
  NOR2  g01257(.A(new_n1642_), .B(new_n910_), .Y(new_n1643_));
  NOR2  g01258(.A(new_n1643_), .B(new_n914_), .Y(new_n1644_));
  NOR2  g01259(.A(new_n1644_), .B(new_n919_), .Y(new_n1645_));
  NOR2  g01260(.A(new_n1645_), .B(new_n923_), .Y(new_n1646_));
  NOR2  g01261(.A(new_n1646_), .B(new_n928_), .Y(new_n1647_));
  NOR2  g01262(.A(new_n1647_), .B(new_n932_), .Y(new_n1648_));
  NOR2  g01263(.A(new_n1648_), .B(new_n937_), .Y(new_n1649_));
  NOR2  g01264(.A(new_n1649_), .B(new_n941_), .Y(new_n1650_));
  NOR2  g01265(.A(new_n1650_), .B(new_n946_), .Y(new_n1651_));
  NOR2  g01266(.A(new_n1651_), .B(new_n950_), .Y(new_n1652_));
  NOR2  g01267(.A(new_n1652_), .B(new_n955_), .Y(new_n1653_));
  NOR2  g01268(.A(new_n1653_), .B(new_n959_), .Y(new_n1654_));
  NOR2  g01269(.A(new_n1654_), .B(new_n964_), .Y(new_n1655_));
  NOR2  g01270(.A(new_n1655_), .B(new_n968_), .Y(new_n1656_));
  NOR2  g01271(.A(new_n1656_), .B(new_n973_), .Y(new_n1657_));
  NOR2  g01272(.A(new_n1657_), .B(new_n977_), .Y(new_n1658_));
  NOR2  g01273(.A(new_n1658_), .B(new_n982_), .Y(new_n1659_));
  NOR2  g01274(.A(new_n1659_), .B(new_n986_), .Y(new_n1660_));
  NOR2  g01275(.A(new_n1660_), .B(new_n991_), .Y(new_n1661_));
  NOR2  g01276(.A(new_n1661_), .B(new_n995_), .Y(new_n1662_));
  NOR2  g01277(.A(new_n1662_), .B(new_n1000_), .Y(new_n1663_));
  NOR2  g01278(.A(new_n1663_), .B(new_n1004_), .Y(new_n1664_));
  NOR2  g01279(.A(new_n1664_), .B(new_n1009_), .Y(new_n1665_));
  NOR2  g01280(.A(new_n1665_), .B(new_n1013_), .Y(new_n1666_));
  NOR2  g01281(.A(new_n1666_), .B(new_n1018_), .Y(new_n1667_));
  NOR2  g01282(.A(new_n1667_), .B(new_n1022_), .Y(new_n1668_));
  NOR2  g01283(.A(new_n1668_), .B(new_n1027_), .Y(new_n1669_));
  NOR2  g01284(.A(new_n1669_), .B(new_n1031_), .Y(new_n1670_));
  NOR2  g01285(.A(new_n1670_), .B(new_n1036_), .Y(new_n1671_));
  NOR2  g01286(.A(new_n1671_), .B(new_n1040_), .Y(new_n1672_));
  NOR2  g01287(.A(new_n1672_), .B(new_n1045_), .Y(new_n1673_));
  NOR2  g01288(.A(new_n1673_), .B(new_n1049_), .Y(new_n1674_));
  NOR2  g01289(.A(new_n1674_), .B(new_n1054_), .Y(new_n1675_));
  NOR2  g01290(.A(new_n1675_), .B(new_n1058_), .Y(new_n1676_));
  NOR2  g01291(.A(new_n1676_), .B(new_n1063_), .Y(new_n1677_));
  NOR2  g01292(.A(new_n1677_), .B(new_n1067_), .Y(new_n1678_));
  NOR2  g01293(.A(new_n1678_), .B(new_n1072_), .Y(new_n1679_));
  NOR2  g01294(.A(new_n1679_), .B(new_n1076_), .Y(new_n1680_));
  NOR2  g01295(.A(new_n1680_), .B(new_n1081_), .Y(new_n1681_));
  NOR2  g01296(.A(new_n1681_), .B(new_n1085_), .Y(new_n1682_));
  NOR2  g01297(.A(new_n1682_), .B(new_n1090_), .Y(new_n1683_));
  NOR2  g01298(.A(new_n1683_), .B(new_n1094_), .Y(new_n1684_));
  NOR2  g01299(.A(new_n1684_), .B(new_n1099_), .Y(new_n1685_));
  NOR2  g01300(.A(new_n1685_), .B(new_n1103_), .Y(new_n1686_));
  NOR2  g01301(.A(new_n1686_), .B(new_n1108_), .Y(new_n1687_));
  NOR2  g01302(.A(new_n1687_), .B(new_n1112_), .Y(new_n1688_));
  NOR2  g01303(.A(new_n1688_), .B(new_n1117_), .Y(new_n1689_));
  NOR2  g01304(.A(new_n1689_), .B(new_n1121_), .Y(new_n1690_));
  NOR2  g01305(.A(new_n1690_), .B(new_n1126_), .Y(new_n1691_));
  NOR2  g01306(.A(new_n1691_), .B(new_n1130_), .Y(new_n1692_));
  NOR2  g01307(.A(new_n1692_), .B(new_n1135_), .Y(new_n1693_));
  NOR2  g01308(.A(new_n1693_), .B(new_n1139_), .Y(new_n1694_));
  NOR2  g01309(.A(new_n1694_), .B(new_n1144_), .Y(new_n1695_));
  NOR2  g01310(.A(new_n1695_), .B(new_n1148_), .Y(new_n1696_));
  NOR2  g01311(.A(new_n1696_), .B(new_n1153_), .Y(new_n1697_));
  NOR2  g01312(.A(new_n1697_), .B(new_n1157_), .Y(new_n1698_));
  NOR2  g01313(.A(new_n1698_), .B(new_n1162_), .Y(new_n1699_));
  NOR2  g01314(.A(new_n1699_), .B(new_n1166_), .Y(new_n1700_));
  NOR2  g01315(.A(new_n1700_), .B(new_n1171_), .Y(new_n1701_));
  NOR2  g01316(.A(new_n1701_), .B(new_n1175_), .Y(new_n1702_));
  NOR2  g01317(.A(new_n1702_), .B(new_n1180_), .Y(new_n1703_));
  NOR2  g01318(.A(new_n1703_), .B(new_n1184_), .Y(new_n1704_));
  NOR2  g01319(.A(new_n1704_), .B(new_n1189_), .Y(new_n1705_));
  NOR2  g01320(.A(\req[2] ), .B(\req[1] ), .Y(new_n1706_));
  NAND2 g01321(.A(new_n1706_), .B(new_n1191_), .Y(new_n1707_));
  NOR2  g01322(.A(new_n1707_), .B(new_n1705_), .Y(new_n1708_));
  NAND2 g01323(.A(new_n813_), .B(new_n817_), .Y(new_n1709_));
  NOR2  g01324(.A(new_n1709_), .B(new_n1708_), .Y(new_n1710_));
  NAND2 g01325(.A(\req[3] ), .B(new_n817_), .Y(new_n1711_));
  NAND2 g01326(.A(new_n1711_), .B(\req[4] ), .Y(new_n1712_));
  NOR2  g01327(.A(new_n1712_), .B(new_n1710_), .Y(\grant[4] ));
  INV   g01328(.A(new_n1202_), .Y(new_n1714_));
  NOR2  g01329(.A(new_n1714_), .B(new_n405_), .Y(new_n1715_));
  NOR2  g01330(.A(new_n1715_), .B(new_n1207_), .Y(new_n1716_));
  NOR2  g01331(.A(new_n1716_), .B(new_n1211_), .Y(new_n1717_));
  NOR2  g01332(.A(new_n1717_), .B(new_n1215_), .Y(new_n1718_));
  NOR2  g01333(.A(new_n1718_), .B(new_n1219_), .Y(new_n1719_));
  NOR2  g01334(.A(new_n1719_), .B(new_n1223_), .Y(new_n1720_));
  NOR2  g01335(.A(new_n1720_), .B(new_n1227_), .Y(new_n1721_));
  NOR2  g01336(.A(new_n1721_), .B(new_n1231_), .Y(new_n1722_));
  NOR2  g01337(.A(new_n1722_), .B(new_n1235_), .Y(new_n1723_));
  NOR2  g01338(.A(new_n1723_), .B(new_n1239_), .Y(new_n1724_));
  NOR2  g01339(.A(new_n1724_), .B(new_n1243_), .Y(new_n1725_));
  NOR2  g01340(.A(new_n1725_), .B(new_n1247_), .Y(new_n1726_));
  NOR2  g01341(.A(new_n1726_), .B(new_n1251_), .Y(new_n1727_));
  NOR2  g01342(.A(new_n1727_), .B(new_n1255_), .Y(new_n1728_));
  NOR2  g01343(.A(new_n1728_), .B(new_n1259_), .Y(new_n1729_));
  NOR2  g01344(.A(new_n1729_), .B(new_n1263_), .Y(new_n1730_));
  NOR2  g01345(.A(new_n1730_), .B(new_n1267_), .Y(new_n1731_));
  NOR2  g01346(.A(new_n1731_), .B(new_n1271_), .Y(new_n1732_));
  NOR2  g01347(.A(new_n1732_), .B(new_n1275_), .Y(new_n1733_));
  NOR2  g01348(.A(new_n1733_), .B(new_n1279_), .Y(new_n1734_));
  NOR2  g01349(.A(new_n1734_), .B(new_n1283_), .Y(new_n1735_));
  NOR2  g01350(.A(new_n1735_), .B(new_n1287_), .Y(new_n1736_));
  NOR2  g01351(.A(new_n1736_), .B(new_n1291_), .Y(new_n1737_));
  NOR2  g01352(.A(new_n1737_), .B(new_n1295_), .Y(new_n1738_));
  NOR2  g01353(.A(new_n1738_), .B(new_n1299_), .Y(new_n1739_));
  NOR2  g01354(.A(new_n1739_), .B(new_n1303_), .Y(new_n1740_));
  NOR2  g01355(.A(new_n1740_), .B(new_n1307_), .Y(new_n1741_));
  NOR2  g01356(.A(new_n1741_), .B(new_n1311_), .Y(new_n1742_));
  NOR2  g01357(.A(new_n1742_), .B(new_n1315_), .Y(new_n1743_));
  NOR2  g01358(.A(new_n1743_), .B(new_n1319_), .Y(new_n1744_));
  NOR2  g01359(.A(new_n1744_), .B(new_n1323_), .Y(new_n1745_));
  NOR2  g01360(.A(new_n1745_), .B(new_n1327_), .Y(new_n1746_));
  NOR2  g01361(.A(new_n1746_), .B(new_n1331_), .Y(new_n1747_));
  NOR2  g01362(.A(new_n1747_), .B(new_n1335_), .Y(new_n1748_));
  NOR2  g01363(.A(new_n1748_), .B(new_n1339_), .Y(new_n1749_));
  NOR2  g01364(.A(new_n1749_), .B(new_n1343_), .Y(new_n1750_));
  NOR2  g01365(.A(new_n1750_), .B(new_n1347_), .Y(new_n1751_));
  NOR2  g01366(.A(new_n1751_), .B(new_n1351_), .Y(new_n1752_));
  NOR2  g01367(.A(new_n1752_), .B(new_n1355_), .Y(new_n1753_));
  NOR2  g01368(.A(new_n1753_), .B(new_n1359_), .Y(new_n1754_));
  NOR2  g01369(.A(new_n1754_), .B(new_n1363_), .Y(new_n1755_));
  NOR2  g01370(.A(new_n1755_), .B(new_n1367_), .Y(new_n1756_));
  NOR2  g01371(.A(new_n1756_), .B(new_n1371_), .Y(new_n1757_));
  NOR2  g01372(.A(new_n1757_), .B(new_n1375_), .Y(new_n1758_));
  NOR2  g01373(.A(new_n1758_), .B(new_n1379_), .Y(new_n1759_));
  NOR2  g01374(.A(new_n1759_), .B(new_n1383_), .Y(new_n1760_));
  NOR2  g01375(.A(new_n1760_), .B(new_n1387_), .Y(new_n1761_));
  NOR2  g01376(.A(new_n1761_), .B(new_n1391_), .Y(new_n1762_));
  NOR2  g01377(.A(new_n1762_), .B(new_n1395_), .Y(new_n1763_));
  NOR2  g01378(.A(new_n1763_), .B(new_n1399_), .Y(new_n1764_));
  NOR2  g01379(.A(new_n1764_), .B(new_n1403_), .Y(new_n1765_));
  NOR2  g01380(.A(new_n1765_), .B(new_n1407_), .Y(new_n1766_));
  NOR2  g01381(.A(new_n1766_), .B(new_n1411_), .Y(new_n1767_));
  NOR2  g01382(.A(new_n1767_), .B(new_n1415_), .Y(new_n1768_));
  NOR2  g01383(.A(new_n1768_), .B(new_n1419_), .Y(new_n1769_));
  NOR2  g01384(.A(new_n1769_), .B(new_n1423_), .Y(new_n1770_));
  NOR2  g01385(.A(new_n1770_), .B(new_n1427_), .Y(new_n1771_));
  NOR2  g01386(.A(new_n1771_), .B(new_n1431_), .Y(new_n1772_));
  NOR2  g01387(.A(new_n1772_), .B(new_n1435_), .Y(new_n1773_));
  NOR2  g01388(.A(new_n1773_), .B(new_n1439_), .Y(new_n1774_));
  NOR2  g01389(.A(new_n1774_), .B(new_n1443_), .Y(new_n1775_));
  NOR2  g01390(.A(new_n1775_), .B(new_n1447_), .Y(new_n1776_));
  NOR2  g01391(.A(new_n1776_), .B(new_n1451_), .Y(new_n1777_));
  NOR2  g01392(.A(new_n1777_), .B(new_n1455_), .Y(new_n1778_));
  NOR2  g01393(.A(new_n1778_), .B(new_n1459_), .Y(new_n1779_));
  NOR2  g01394(.A(new_n1779_), .B(new_n1463_), .Y(new_n1780_));
  NOR2  g01395(.A(new_n1780_), .B(new_n1467_), .Y(new_n1781_));
  NOR2  g01396(.A(new_n1781_), .B(new_n1471_), .Y(new_n1782_));
  NOR2  g01397(.A(new_n1782_), .B(new_n1475_), .Y(new_n1783_));
  NOR2  g01398(.A(new_n1783_), .B(new_n1479_), .Y(new_n1784_));
  NOR2  g01399(.A(new_n1784_), .B(new_n1483_), .Y(new_n1785_));
  NOR2  g01400(.A(new_n1785_), .B(new_n1487_), .Y(new_n1786_));
  NOR2  g01401(.A(new_n1786_), .B(new_n1491_), .Y(new_n1787_));
  NOR2  g01402(.A(new_n1787_), .B(new_n1495_), .Y(new_n1788_));
  NOR2  g01403(.A(new_n1788_), .B(new_n1499_), .Y(new_n1789_));
  NOR2  g01404(.A(new_n1789_), .B(new_n1503_), .Y(new_n1790_));
  NOR2  g01405(.A(new_n1790_), .B(new_n1507_), .Y(new_n1791_));
  NOR2  g01406(.A(new_n1791_), .B(new_n1511_), .Y(new_n1792_));
  NOR2  g01407(.A(new_n1792_), .B(new_n1515_), .Y(new_n1793_));
  NOR2  g01408(.A(new_n1793_), .B(new_n1519_), .Y(new_n1794_));
  NOR2  g01409(.A(new_n1794_), .B(new_n1523_), .Y(new_n1795_));
  NOR2  g01410(.A(new_n1795_), .B(new_n1527_), .Y(new_n1796_));
  NAND2 g01411(.A(new_n1529_), .B(new_n389_), .Y(new_n1797_));
  NOR2  g01412(.A(new_n1797_), .B(new_n1796_), .Y(new_n1798_));
  NOR2  g01413(.A(new_n1798_), .B(new_n396_), .Y(new_n1799_));
  NAND2 g01414(.A(new_n398_), .B(\req[5] ), .Y(new_n1800_));
  NOR2  g01415(.A(new_n1800_), .B(new_n1799_), .Y(\grant[5] ));
  INV   g01416(.A(new_n409_), .Y(new_n1802_));
  NOR2  g01417(.A(new_n828_), .B(new_n1802_), .Y(new_n1803_));
  NOR2  g01418(.A(new_n1803_), .B(new_n416_), .Y(new_n1804_));
  NOR2  g01419(.A(new_n1804_), .B(new_n420_), .Y(new_n1805_));
  NOR2  g01420(.A(new_n1805_), .B(new_n426_), .Y(new_n1806_));
  NOR2  g01421(.A(new_n1806_), .B(new_n430_), .Y(new_n1807_));
  NOR2  g01422(.A(new_n1807_), .B(new_n436_), .Y(new_n1808_));
  NOR2  g01423(.A(new_n1808_), .B(new_n440_), .Y(new_n1809_));
  NOR2  g01424(.A(new_n1809_), .B(new_n446_), .Y(new_n1810_));
  NOR2  g01425(.A(new_n1810_), .B(new_n450_), .Y(new_n1811_));
  NOR2  g01426(.A(new_n1811_), .B(new_n456_), .Y(new_n1812_));
  NOR2  g01427(.A(new_n1812_), .B(new_n460_), .Y(new_n1813_));
  NOR2  g01428(.A(new_n1813_), .B(new_n466_), .Y(new_n1814_));
  NOR2  g01429(.A(new_n1814_), .B(new_n470_), .Y(new_n1815_));
  NOR2  g01430(.A(new_n1815_), .B(new_n476_), .Y(new_n1816_));
  NOR2  g01431(.A(new_n1816_), .B(new_n480_), .Y(new_n1817_));
  NOR2  g01432(.A(new_n1817_), .B(new_n486_), .Y(new_n1818_));
  NOR2  g01433(.A(new_n1818_), .B(new_n490_), .Y(new_n1819_));
  NOR2  g01434(.A(new_n1819_), .B(new_n496_), .Y(new_n1820_));
  NOR2  g01435(.A(new_n1820_), .B(new_n500_), .Y(new_n1821_));
  NOR2  g01436(.A(new_n1821_), .B(new_n506_), .Y(new_n1822_));
  NOR2  g01437(.A(new_n1822_), .B(new_n510_), .Y(new_n1823_));
  NOR2  g01438(.A(new_n1823_), .B(new_n516_), .Y(new_n1824_));
  NOR2  g01439(.A(new_n1824_), .B(new_n520_), .Y(new_n1825_));
  NOR2  g01440(.A(new_n1825_), .B(new_n526_), .Y(new_n1826_));
  NOR2  g01441(.A(new_n1826_), .B(new_n530_), .Y(new_n1827_));
  NOR2  g01442(.A(new_n1827_), .B(new_n536_), .Y(new_n1828_));
  NOR2  g01443(.A(new_n1828_), .B(new_n540_), .Y(new_n1829_));
  NOR2  g01444(.A(new_n1829_), .B(new_n546_), .Y(new_n1830_));
  NOR2  g01445(.A(new_n1830_), .B(new_n550_), .Y(new_n1831_));
  NOR2  g01446(.A(new_n1831_), .B(new_n556_), .Y(new_n1832_));
  NOR2  g01447(.A(new_n1832_), .B(new_n560_), .Y(new_n1833_));
  NOR2  g01448(.A(new_n1833_), .B(new_n566_), .Y(new_n1834_));
  NOR2  g01449(.A(new_n1834_), .B(new_n570_), .Y(new_n1835_));
  NOR2  g01450(.A(new_n1835_), .B(new_n576_), .Y(new_n1836_));
  NOR2  g01451(.A(new_n1836_), .B(new_n580_), .Y(new_n1837_));
  NOR2  g01452(.A(new_n1837_), .B(new_n586_), .Y(new_n1838_));
  NOR2  g01453(.A(new_n1838_), .B(new_n590_), .Y(new_n1839_));
  NOR2  g01454(.A(new_n1839_), .B(new_n596_), .Y(new_n1840_));
  NOR2  g01455(.A(new_n1840_), .B(new_n600_), .Y(new_n1841_));
  NOR2  g01456(.A(new_n1841_), .B(new_n606_), .Y(new_n1842_));
  NOR2  g01457(.A(new_n1842_), .B(new_n610_), .Y(new_n1843_));
  NOR2  g01458(.A(new_n1843_), .B(new_n616_), .Y(new_n1844_));
  NOR2  g01459(.A(new_n1844_), .B(new_n620_), .Y(new_n1845_));
  NOR2  g01460(.A(new_n1845_), .B(new_n626_), .Y(new_n1846_));
  NOR2  g01461(.A(new_n1846_), .B(new_n630_), .Y(new_n1847_));
  NOR2  g01462(.A(new_n1847_), .B(new_n636_), .Y(new_n1848_));
  NOR2  g01463(.A(new_n1848_), .B(new_n640_), .Y(new_n1849_));
  NOR2  g01464(.A(new_n1849_), .B(new_n646_), .Y(new_n1850_));
  NOR2  g01465(.A(new_n1850_), .B(new_n650_), .Y(new_n1851_));
  NOR2  g01466(.A(new_n1851_), .B(new_n656_), .Y(new_n1852_));
  NOR2  g01467(.A(new_n1852_), .B(new_n660_), .Y(new_n1853_));
  NOR2  g01468(.A(new_n1853_), .B(new_n666_), .Y(new_n1854_));
  NOR2  g01469(.A(new_n1854_), .B(new_n670_), .Y(new_n1855_));
  NOR2  g01470(.A(new_n1855_), .B(new_n676_), .Y(new_n1856_));
  NOR2  g01471(.A(new_n1856_), .B(new_n680_), .Y(new_n1857_));
  NOR2  g01472(.A(new_n1857_), .B(new_n686_), .Y(new_n1858_));
  NOR2  g01473(.A(new_n1858_), .B(new_n690_), .Y(new_n1859_));
  NOR2  g01474(.A(new_n1859_), .B(new_n696_), .Y(new_n1860_));
  NOR2  g01475(.A(new_n1860_), .B(new_n700_), .Y(new_n1861_));
  NOR2  g01476(.A(new_n1861_), .B(new_n706_), .Y(new_n1862_));
  NOR2  g01477(.A(new_n1862_), .B(new_n710_), .Y(new_n1863_));
  NOR2  g01478(.A(new_n1863_), .B(new_n716_), .Y(new_n1864_));
  NOR2  g01479(.A(new_n1864_), .B(new_n720_), .Y(new_n1865_));
  NOR2  g01480(.A(new_n1865_), .B(new_n726_), .Y(new_n1866_));
  NOR2  g01481(.A(new_n1866_), .B(new_n730_), .Y(new_n1867_));
  NOR2  g01482(.A(new_n1867_), .B(new_n736_), .Y(new_n1868_));
  NOR2  g01483(.A(new_n1868_), .B(new_n740_), .Y(new_n1869_));
  NOR2  g01484(.A(new_n1869_), .B(new_n746_), .Y(new_n1870_));
  NOR2  g01485(.A(new_n1870_), .B(new_n750_), .Y(new_n1871_));
  NOR2  g01486(.A(new_n1871_), .B(new_n756_), .Y(new_n1872_));
  NOR2  g01487(.A(new_n1872_), .B(new_n760_), .Y(new_n1873_));
  NOR2  g01488(.A(new_n1873_), .B(new_n766_), .Y(new_n1874_));
  NOR2  g01489(.A(new_n1874_), .B(new_n770_), .Y(new_n1875_));
  NOR2  g01490(.A(new_n1875_), .B(new_n776_), .Y(new_n1876_));
  NOR2  g01491(.A(new_n1876_), .B(new_n780_), .Y(new_n1877_));
  NOR2  g01492(.A(new_n1877_), .B(new_n786_), .Y(new_n1878_));
  NOR2  g01493(.A(new_n1878_), .B(new_n790_), .Y(new_n1879_));
  NOR2  g01494(.A(new_n1879_), .B(new_n796_), .Y(new_n1880_));
  NOR2  g01495(.A(new_n1880_), .B(new_n800_), .Y(new_n1881_));
  NOR2  g01496(.A(new_n1881_), .B(new_n806_), .Y(new_n1882_));
  NOR2  g01497(.A(new_n1882_), .B(new_n1616_), .Y(new_n1883_));
  NOR2  g01498(.A(new_n1883_), .B(new_n1618_), .Y(new_n1884_));
  NAND2 g01499(.A(new_n1620_), .B(new_n814_), .Y(new_n1885_));
  NOR2  g01500(.A(new_n1885_), .B(new_n1884_), .Y(new_n1886_));
  NOR2  g01501(.A(new_n1886_), .B(new_n820_), .Y(new_n1887_));
  NAND2 g01502(.A(new_n822_), .B(\req[6] ), .Y(new_n1888_));
  NOR2  g01503(.A(new_n1888_), .B(new_n1887_), .Y(\grant[6] ));
  INV   g01504(.A(new_n832_), .Y(new_n1890_));
  NOR2  g01505(.A(new_n1206_), .B(new_n1890_), .Y(new_n1891_));
  NOR2  g01506(.A(new_n1891_), .B(new_n838_), .Y(new_n1892_));
  NOR2  g01507(.A(new_n1892_), .B(new_n842_), .Y(new_n1893_));
  NOR2  g01508(.A(new_n1893_), .B(new_n847_), .Y(new_n1894_));
  NOR2  g01509(.A(new_n1894_), .B(new_n851_), .Y(new_n1895_));
  NOR2  g01510(.A(new_n1895_), .B(new_n856_), .Y(new_n1896_));
  NOR2  g01511(.A(new_n1896_), .B(new_n860_), .Y(new_n1897_));
  NOR2  g01512(.A(new_n1897_), .B(new_n865_), .Y(new_n1898_));
  NOR2  g01513(.A(new_n1898_), .B(new_n869_), .Y(new_n1899_));
  NOR2  g01514(.A(new_n1899_), .B(new_n874_), .Y(new_n1900_));
  NOR2  g01515(.A(new_n1900_), .B(new_n878_), .Y(new_n1901_));
  NOR2  g01516(.A(new_n1901_), .B(new_n883_), .Y(new_n1902_));
  NOR2  g01517(.A(new_n1902_), .B(new_n887_), .Y(new_n1903_));
  NOR2  g01518(.A(new_n1903_), .B(new_n892_), .Y(new_n1904_));
  NOR2  g01519(.A(new_n1904_), .B(new_n896_), .Y(new_n1905_));
  NOR2  g01520(.A(new_n1905_), .B(new_n901_), .Y(new_n1906_));
  NOR2  g01521(.A(new_n1906_), .B(new_n905_), .Y(new_n1907_));
  NOR2  g01522(.A(new_n1907_), .B(new_n910_), .Y(new_n1908_));
  NOR2  g01523(.A(new_n1908_), .B(new_n914_), .Y(new_n1909_));
  NOR2  g01524(.A(new_n1909_), .B(new_n919_), .Y(new_n1910_));
  NOR2  g01525(.A(new_n1910_), .B(new_n923_), .Y(new_n1911_));
  NOR2  g01526(.A(new_n1911_), .B(new_n928_), .Y(new_n1912_));
  NOR2  g01527(.A(new_n1912_), .B(new_n932_), .Y(new_n1913_));
  NOR2  g01528(.A(new_n1913_), .B(new_n937_), .Y(new_n1914_));
  NOR2  g01529(.A(new_n1914_), .B(new_n941_), .Y(new_n1915_));
  NOR2  g01530(.A(new_n1915_), .B(new_n946_), .Y(new_n1916_));
  NOR2  g01531(.A(new_n1916_), .B(new_n950_), .Y(new_n1917_));
  NOR2  g01532(.A(new_n1917_), .B(new_n955_), .Y(new_n1918_));
  NOR2  g01533(.A(new_n1918_), .B(new_n959_), .Y(new_n1919_));
  NOR2  g01534(.A(new_n1919_), .B(new_n964_), .Y(new_n1920_));
  NOR2  g01535(.A(new_n1920_), .B(new_n968_), .Y(new_n1921_));
  NOR2  g01536(.A(new_n1921_), .B(new_n973_), .Y(new_n1922_));
  NOR2  g01537(.A(new_n1922_), .B(new_n977_), .Y(new_n1923_));
  NOR2  g01538(.A(new_n1923_), .B(new_n982_), .Y(new_n1924_));
  NOR2  g01539(.A(new_n1924_), .B(new_n986_), .Y(new_n1925_));
  NOR2  g01540(.A(new_n1925_), .B(new_n991_), .Y(new_n1926_));
  NOR2  g01541(.A(new_n1926_), .B(new_n995_), .Y(new_n1927_));
  NOR2  g01542(.A(new_n1927_), .B(new_n1000_), .Y(new_n1928_));
  NOR2  g01543(.A(new_n1928_), .B(new_n1004_), .Y(new_n1929_));
  NOR2  g01544(.A(new_n1929_), .B(new_n1009_), .Y(new_n1930_));
  NOR2  g01545(.A(new_n1930_), .B(new_n1013_), .Y(new_n1931_));
  NOR2  g01546(.A(new_n1931_), .B(new_n1018_), .Y(new_n1932_));
  NOR2  g01547(.A(new_n1932_), .B(new_n1022_), .Y(new_n1933_));
  NOR2  g01548(.A(new_n1933_), .B(new_n1027_), .Y(new_n1934_));
  NOR2  g01549(.A(new_n1934_), .B(new_n1031_), .Y(new_n1935_));
  NOR2  g01550(.A(new_n1935_), .B(new_n1036_), .Y(new_n1936_));
  NOR2  g01551(.A(new_n1936_), .B(new_n1040_), .Y(new_n1937_));
  NOR2  g01552(.A(new_n1937_), .B(new_n1045_), .Y(new_n1938_));
  NOR2  g01553(.A(new_n1938_), .B(new_n1049_), .Y(new_n1939_));
  NOR2  g01554(.A(new_n1939_), .B(new_n1054_), .Y(new_n1940_));
  NOR2  g01555(.A(new_n1940_), .B(new_n1058_), .Y(new_n1941_));
  NOR2  g01556(.A(new_n1941_), .B(new_n1063_), .Y(new_n1942_));
  NOR2  g01557(.A(new_n1942_), .B(new_n1067_), .Y(new_n1943_));
  NOR2  g01558(.A(new_n1943_), .B(new_n1072_), .Y(new_n1944_));
  NOR2  g01559(.A(new_n1944_), .B(new_n1076_), .Y(new_n1945_));
  NOR2  g01560(.A(new_n1945_), .B(new_n1081_), .Y(new_n1946_));
  NOR2  g01561(.A(new_n1946_), .B(new_n1085_), .Y(new_n1947_));
  NOR2  g01562(.A(new_n1947_), .B(new_n1090_), .Y(new_n1948_));
  NOR2  g01563(.A(new_n1948_), .B(new_n1094_), .Y(new_n1949_));
  NOR2  g01564(.A(new_n1949_), .B(new_n1099_), .Y(new_n1950_));
  NOR2  g01565(.A(new_n1950_), .B(new_n1103_), .Y(new_n1951_));
  NOR2  g01566(.A(new_n1951_), .B(new_n1108_), .Y(new_n1952_));
  NOR2  g01567(.A(new_n1952_), .B(new_n1112_), .Y(new_n1953_));
  NOR2  g01568(.A(new_n1953_), .B(new_n1117_), .Y(new_n1954_));
  NOR2  g01569(.A(new_n1954_), .B(new_n1121_), .Y(new_n1955_));
  NOR2  g01570(.A(new_n1955_), .B(new_n1126_), .Y(new_n1956_));
  NOR2  g01571(.A(new_n1956_), .B(new_n1130_), .Y(new_n1957_));
  NOR2  g01572(.A(new_n1957_), .B(new_n1135_), .Y(new_n1958_));
  NOR2  g01573(.A(new_n1958_), .B(new_n1139_), .Y(new_n1959_));
  NOR2  g01574(.A(new_n1959_), .B(new_n1144_), .Y(new_n1960_));
  NOR2  g01575(.A(new_n1960_), .B(new_n1148_), .Y(new_n1961_));
  NOR2  g01576(.A(new_n1961_), .B(new_n1153_), .Y(new_n1962_));
  NOR2  g01577(.A(new_n1962_), .B(new_n1157_), .Y(new_n1963_));
  NOR2  g01578(.A(new_n1963_), .B(new_n1162_), .Y(new_n1964_));
  NOR2  g01579(.A(new_n1964_), .B(new_n1166_), .Y(new_n1965_));
  NOR2  g01580(.A(new_n1965_), .B(new_n1171_), .Y(new_n1966_));
  NOR2  g01581(.A(new_n1966_), .B(new_n1175_), .Y(new_n1967_));
  NOR2  g01582(.A(new_n1967_), .B(new_n1180_), .Y(new_n1968_));
  NOR2  g01583(.A(new_n1968_), .B(new_n1184_), .Y(new_n1969_));
  NOR2  g01584(.A(new_n1969_), .B(new_n1189_), .Y(new_n1970_));
  NOR2  g01585(.A(new_n1970_), .B(new_n1707_), .Y(new_n1971_));
  NOR2  g01586(.A(new_n1971_), .B(new_n1709_), .Y(new_n1972_));
  NAND2 g01587(.A(new_n1711_), .B(new_n1194_), .Y(new_n1973_));
  NOR2  g01588(.A(new_n1973_), .B(new_n1972_), .Y(new_n1974_));
  NOR2  g01589(.A(new_n1974_), .B(new_n1199_), .Y(new_n1975_));
  NAND2 g01590(.A(new_n1201_), .B(\req[7] ), .Y(new_n1976_));
  NOR2  g01591(.A(new_n1976_), .B(new_n1975_), .Y(\grant[7] ));
  INV   g01592(.A(new_n1210_), .Y(new_n1978_));
  NOR2  g01593(.A(new_n1978_), .B(new_n415_), .Y(new_n1979_));
  NOR2  g01594(.A(new_n1979_), .B(new_n1215_), .Y(new_n1980_));
  NOR2  g01595(.A(new_n1980_), .B(new_n1219_), .Y(new_n1981_));
  NOR2  g01596(.A(new_n1981_), .B(new_n1223_), .Y(new_n1982_));
  NOR2  g01597(.A(new_n1982_), .B(new_n1227_), .Y(new_n1983_));
  NOR2  g01598(.A(new_n1983_), .B(new_n1231_), .Y(new_n1984_));
  NOR2  g01599(.A(new_n1984_), .B(new_n1235_), .Y(new_n1985_));
  NOR2  g01600(.A(new_n1985_), .B(new_n1239_), .Y(new_n1986_));
  NOR2  g01601(.A(new_n1986_), .B(new_n1243_), .Y(new_n1987_));
  NOR2  g01602(.A(new_n1987_), .B(new_n1247_), .Y(new_n1988_));
  NOR2  g01603(.A(new_n1988_), .B(new_n1251_), .Y(new_n1989_));
  NOR2  g01604(.A(new_n1989_), .B(new_n1255_), .Y(new_n1990_));
  NOR2  g01605(.A(new_n1990_), .B(new_n1259_), .Y(new_n1991_));
  NOR2  g01606(.A(new_n1991_), .B(new_n1263_), .Y(new_n1992_));
  NOR2  g01607(.A(new_n1992_), .B(new_n1267_), .Y(new_n1993_));
  NOR2  g01608(.A(new_n1993_), .B(new_n1271_), .Y(new_n1994_));
  NOR2  g01609(.A(new_n1994_), .B(new_n1275_), .Y(new_n1995_));
  NOR2  g01610(.A(new_n1995_), .B(new_n1279_), .Y(new_n1996_));
  NOR2  g01611(.A(new_n1996_), .B(new_n1283_), .Y(new_n1997_));
  NOR2  g01612(.A(new_n1997_), .B(new_n1287_), .Y(new_n1998_));
  NOR2  g01613(.A(new_n1998_), .B(new_n1291_), .Y(new_n1999_));
  NOR2  g01614(.A(new_n1999_), .B(new_n1295_), .Y(new_n2000_));
  NOR2  g01615(.A(new_n2000_), .B(new_n1299_), .Y(new_n2001_));
  NOR2  g01616(.A(new_n2001_), .B(new_n1303_), .Y(new_n2002_));
  NOR2  g01617(.A(new_n2002_), .B(new_n1307_), .Y(new_n2003_));
  NOR2  g01618(.A(new_n2003_), .B(new_n1311_), .Y(new_n2004_));
  NOR2  g01619(.A(new_n2004_), .B(new_n1315_), .Y(new_n2005_));
  NOR2  g01620(.A(new_n2005_), .B(new_n1319_), .Y(new_n2006_));
  NOR2  g01621(.A(new_n2006_), .B(new_n1323_), .Y(new_n2007_));
  NOR2  g01622(.A(new_n2007_), .B(new_n1327_), .Y(new_n2008_));
  NOR2  g01623(.A(new_n2008_), .B(new_n1331_), .Y(new_n2009_));
  NOR2  g01624(.A(new_n2009_), .B(new_n1335_), .Y(new_n2010_));
  NOR2  g01625(.A(new_n2010_), .B(new_n1339_), .Y(new_n2011_));
  NOR2  g01626(.A(new_n2011_), .B(new_n1343_), .Y(new_n2012_));
  NOR2  g01627(.A(new_n2012_), .B(new_n1347_), .Y(new_n2013_));
  NOR2  g01628(.A(new_n2013_), .B(new_n1351_), .Y(new_n2014_));
  NOR2  g01629(.A(new_n2014_), .B(new_n1355_), .Y(new_n2015_));
  NOR2  g01630(.A(new_n2015_), .B(new_n1359_), .Y(new_n2016_));
  NOR2  g01631(.A(new_n2016_), .B(new_n1363_), .Y(new_n2017_));
  NOR2  g01632(.A(new_n2017_), .B(new_n1367_), .Y(new_n2018_));
  NOR2  g01633(.A(new_n2018_), .B(new_n1371_), .Y(new_n2019_));
  NOR2  g01634(.A(new_n2019_), .B(new_n1375_), .Y(new_n2020_));
  NOR2  g01635(.A(new_n2020_), .B(new_n1379_), .Y(new_n2021_));
  NOR2  g01636(.A(new_n2021_), .B(new_n1383_), .Y(new_n2022_));
  NOR2  g01637(.A(new_n2022_), .B(new_n1387_), .Y(new_n2023_));
  NOR2  g01638(.A(new_n2023_), .B(new_n1391_), .Y(new_n2024_));
  NOR2  g01639(.A(new_n2024_), .B(new_n1395_), .Y(new_n2025_));
  NOR2  g01640(.A(new_n2025_), .B(new_n1399_), .Y(new_n2026_));
  NOR2  g01641(.A(new_n2026_), .B(new_n1403_), .Y(new_n2027_));
  NOR2  g01642(.A(new_n2027_), .B(new_n1407_), .Y(new_n2028_));
  NOR2  g01643(.A(new_n2028_), .B(new_n1411_), .Y(new_n2029_));
  NOR2  g01644(.A(new_n2029_), .B(new_n1415_), .Y(new_n2030_));
  NOR2  g01645(.A(new_n2030_), .B(new_n1419_), .Y(new_n2031_));
  NOR2  g01646(.A(new_n2031_), .B(new_n1423_), .Y(new_n2032_));
  NOR2  g01647(.A(new_n2032_), .B(new_n1427_), .Y(new_n2033_));
  NOR2  g01648(.A(new_n2033_), .B(new_n1431_), .Y(new_n2034_));
  NOR2  g01649(.A(new_n2034_), .B(new_n1435_), .Y(new_n2035_));
  NOR2  g01650(.A(new_n2035_), .B(new_n1439_), .Y(new_n2036_));
  NOR2  g01651(.A(new_n2036_), .B(new_n1443_), .Y(new_n2037_));
  NOR2  g01652(.A(new_n2037_), .B(new_n1447_), .Y(new_n2038_));
  NOR2  g01653(.A(new_n2038_), .B(new_n1451_), .Y(new_n2039_));
  NOR2  g01654(.A(new_n2039_), .B(new_n1455_), .Y(new_n2040_));
  NOR2  g01655(.A(new_n2040_), .B(new_n1459_), .Y(new_n2041_));
  NOR2  g01656(.A(new_n2041_), .B(new_n1463_), .Y(new_n2042_));
  NOR2  g01657(.A(new_n2042_), .B(new_n1467_), .Y(new_n2043_));
  NOR2  g01658(.A(new_n2043_), .B(new_n1471_), .Y(new_n2044_));
  NOR2  g01659(.A(new_n2044_), .B(new_n1475_), .Y(new_n2045_));
  NOR2  g01660(.A(new_n2045_), .B(new_n1479_), .Y(new_n2046_));
  NOR2  g01661(.A(new_n2046_), .B(new_n1483_), .Y(new_n2047_));
  NOR2  g01662(.A(new_n2047_), .B(new_n1487_), .Y(new_n2048_));
  NOR2  g01663(.A(new_n2048_), .B(new_n1491_), .Y(new_n2049_));
  NOR2  g01664(.A(new_n2049_), .B(new_n1495_), .Y(new_n2050_));
  NOR2  g01665(.A(new_n2050_), .B(new_n1499_), .Y(new_n2051_));
  NOR2  g01666(.A(new_n2051_), .B(new_n1503_), .Y(new_n2052_));
  NOR2  g01667(.A(new_n2052_), .B(new_n1507_), .Y(new_n2053_));
  NOR2  g01668(.A(new_n2053_), .B(new_n1511_), .Y(new_n2054_));
  NOR2  g01669(.A(new_n2054_), .B(new_n1515_), .Y(new_n2055_));
  NOR2  g01670(.A(new_n2055_), .B(new_n1519_), .Y(new_n2056_));
  NOR2  g01671(.A(new_n2056_), .B(new_n1523_), .Y(new_n2057_));
  NOR2  g01672(.A(new_n2057_), .B(new_n1527_), .Y(new_n2058_));
  NOR2  g01673(.A(new_n2058_), .B(new_n1797_), .Y(new_n2059_));
  NOR2  g01674(.A(new_n2059_), .B(new_n396_), .Y(new_n2060_));
  NOR2  g01675(.A(new_n2060_), .B(new_n400_), .Y(new_n2061_));
  NOR2  g01676(.A(new_n2061_), .B(new_n406_), .Y(new_n2062_));
  NAND2 g01677(.A(new_n408_), .B(\req[8] ), .Y(new_n2063_));
  NOR2  g01678(.A(new_n2063_), .B(new_n2062_), .Y(\grant[8] ));
  INV   g01679(.A(new_n419_), .Y(new_n2065_));
  NOR2  g01680(.A(new_n837_), .B(new_n2065_), .Y(new_n2066_));
  NOR2  g01681(.A(new_n2066_), .B(new_n426_), .Y(new_n2067_));
  NOR2  g01682(.A(new_n2067_), .B(new_n430_), .Y(new_n2068_));
  NOR2  g01683(.A(new_n2068_), .B(new_n436_), .Y(new_n2069_));
  NOR2  g01684(.A(new_n2069_), .B(new_n440_), .Y(new_n2070_));
  NOR2  g01685(.A(new_n2070_), .B(new_n446_), .Y(new_n2071_));
  NOR2  g01686(.A(new_n2071_), .B(new_n450_), .Y(new_n2072_));
  NOR2  g01687(.A(new_n2072_), .B(new_n456_), .Y(new_n2073_));
  NOR2  g01688(.A(new_n2073_), .B(new_n460_), .Y(new_n2074_));
  NOR2  g01689(.A(new_n2074_), .B(new_n466_), .Y(new_n2075_));
  NOR2  g01690(.A(new_n2075_), .B(new_n470_), .Y(new_n2076_));
  NOR2  g01691(.A(new_n2076_), .B(new_n476_), .Y(new_n2077_));
  NOR2  g01692(.A(new_n2077_), .B(new_n480_), .Y(new_n2078_));
  NOR2  g01693(.A(new_n2078_), .B(new_n486_), .Y(new_n2079_));
  NOR2  g01694(.A(new_n2079_), .B(new_n490_), .Y(new_n2080_));
  NOR2  g01695(.A(new_n2080_), .B(new_n496_), .Y(new_n2081_));
  NOR2  g01696(.A(new_n2081_), .B(new_n500_), .Y(new_n2082_));
  NOR2  g01697(.A(new_n2082_), .B(new_n506_), .Y(new_n2083_));
  NOR2  g01698(.A(new_n2083_), .B(new_n510_), .Y(new_n2084_));
  NOR2  g01699(.A(new_n2084_), .B(new_n516_), .Y(new_n2085_));
  NOR2  g01700(.A(new_n2085_), .B(new_n520_), .Y(new_n2086_));
  NOR2  g01701(.A(new_n2086_), .B(new_n526_), .Y(new_n2087_));
  NOR2  g01702(.A(new_n2087_), .B(new_n530_), .Y(new_n2088_));
  NOR2  g01703(.A(new_n2088_), .B(new_n536_), .Y(new_n2089_));
  NOR2  g01704(.A(new_n2089_), .B(new_n540_), .Y(new_n2090_));
  NOR2  g01705(.A(new_n2090_), .B(new_n546_), .Y(new_n2091_));
  NOR2  g01706(.A(new_n2091_), .B(new_n550_), .Y(new_n2092_));
  NOR2  g01707(.A(new_n2092_), .B(new_n556_), .Y(new_n2093_));
  NOR2  g01708(.A(new_n2093_), .B(new_n560_), .Y(new_n2094_));
  NOR2  g01709(.A(new_n2094_), .B(new_n566_), .Y(new_n2095_));
  NOR2  g01710(.A(new_n2095_), .B(new_n570_), .Y(new_n2096_));
  NOR2  g01711(.A(new_n2096_), .B(new_n576_), .Y(new_n2097_));
  NOR2  g01712(.A(new_n2097_), .B(new_n580_), .Y(new_n2098_));
  NOR2  g01713(.A(new_n2098_), .B(new_n586_), .Y(new_n2099_));
  NOR2  g01714(.A(new_n2099_), .B(new_n590_), .Y(new_n2100_));
  NOR2  g01715(.A(new_n2100_), .B(new_n596_), .Y(new_n2101_));
  NOR2  g01716(.A(new_n2101_), .B(new_n600_), .Y(new_n2102_));
  NOR2  g01717(.A(new_n2102_), .B(new_n606_), .Y(new_n2103_));
  NOR2  g01718(.A(new_n2103_), .B(new_n610_), .Y(new_n2104_));
  NOR2  g01719(.A(new_n2104_), .B(new_n616_), .Y(new_n2105_));
  NOR2  g01720(.A(new_n2105_), .B(new_n620_), .Y(new_n2106_));
  NOR2  g01721(.A(new_n2106_), .B(new_n626_), .Y(new_n2107_));
  NOR2  g01722(.A(new_n2107_), .B(new_n630_), .Y(new_n2108_));
  NOR2  g01723(.A(new_n2108_), .B(new_n636_), .Y(new_n2109_));
  NOR2  g01724(.A(new_n2109_), .B(new_n640_), .Y(new_n2110_));
  NOR2  g01725(.A(new_n2110_), .B(new_n646_), .Y(new_n2111_));
  NOR2  g01726(.A(new_n2111_), .B(new_n650_), .Y(new_n2112_));
  NOR2  g01727(.A(new_n2112_), .B(new_n656_), .Y(new_n2113_));
  NOR2  g01728(.A(new_n2113_), .B(new_n660_), .Y(new_n2114_));
  NOR2  g01729(.A(new_n2114_), .B(new_n666_), .Y(new_n2115_));
  NOR2  g01730(.A(new_n2115_), .B(new_n670_), .Y(new_n2116_));
  NOR2  g01731(.A(new_n2116_), .B(new_n676_), .Y(new_n2117_));
  NOR2  g01732(.A(new_n2117_), .B(new_n680_), .Y(new_n2118_));
  NOR2  g01733(.A(new_n2118_), .B(new_n686_), .Y(new_n2119_));
  NOR2  g01734(.A(new_n2119_), .B(new_n690_), .Y(new_n2120_));
  NOR2  g01735(.A(new_n2120_), .B(new_n696_), .Y(new_n2121_));
  NOR2  g01736(.A(new_n2121_), .B(new_n700_), .Y(new_n2122_));
  NOR2  g01737(.A(new_n2122_), .B(new_n706_), .Y(new_n2123_));
  NOR2  g01738(.A(new_n2123_), .B(new_n710_), .Y(new_n2124_));
  NOR2  g01739(.A(new_n2124_), .B(new_n716_), .Y(new_n2125_));
  NOR2  g01740(.A(new_n2125_), .B(new_n720_), .Y(new_n2126_));
  NOR2  g01741(.A(new_n2126_), .B(new_n726_), .Y(new_n2127_));
  NOR2  g01742(.A(new_n2127_), .B(new_n730_), .Y(new_n2128_));
  NOR2  g01743(.A(new_n2128_), .B(new_n736_), .Y(new_n2129_));
  NOR2  g01744(.A(new_n2129_), .B(new_n740_), .Y(new_n2130_));
  NOR2  g01745(.A(new_n2130_), .B(new_n746_), .Y(new_n2131_));
  NOR2  g01746(.A(new_n2131_), .B(new_n750_), .Y(new_n2132_));
  NOR2  g01747(.A(new_n2132_), .B(new_n756_), .Y(new_n2133_));
  NOR2  g01748(.A(new_n2133_), .B(new_n760_), .Y(new_n2134_));
  NOR2  g01749(.A(new_n2134_), .B(new_n766_), .Y(new_n2135_));
  NOR2  g01750(.A(new_n2135_), .B(new_n770_), .Y(new_n2136_));
  NOR2  g01751(.A(new_n2136_), .B(new_n776_), .Y(new_n2137_));
  NOR2  g01752(.A(new_n2137_), .B(new_n780_), .Y(new_n2138_));
  NOR2  g01753(.A(new_n2138_), .B(new_n786_), .Y(new_n2139_));
  NOR2  g01754(.A(new_n2139_), .B(new_n790_), .Y(new_n2140_));
  NOR2  g01755(.A(new_n2140_), .B(new_n796_), .Y(new_n2141_));
  NOR2  g01756(.A(new_n2141_), .B(new_n800_), .Y(new_n2142_));
  NOR2  g01757(.A(new_n2142_), .B(new_n806_), .Y(new_n2143_));
  NOR2  g01758(.A(new_n2143_), .B(new_n1616_), .Y(new_n2144_));
  NOR2  g01759(.A(new_n2144_), .B(new_n1618_), .Y(new_n2145_));
  NOR2  g01760(.A(new_n2145_), .B(new_n1885_), .Y(new_n2146_));
  NOR2  g01761(.A(new_n2146_), .B(new_n820_), .Y(new_n2147_));
  NOR2  g01762(.A(new_n2147_), .B(new_n824_), .Y(new_n2148_));
  NOR2  g01763(.A(new_n2148_), .B(new_n829_), .Y(new_n2149_));
  NAND2 g01764(.A(new_n831_), .B(\req[9] ), .Y(new_n2150_));
  NOR2  g01765(.A(new_n2150_), .B(new_n2149_), .Y(\grant[9] ));
  INV   g01766(.A(new_n841_), .Y(new_n2152_));
  NOR2  g01767(.A(new_n1214_), .B(new_n2152_), .Y(new_n2153_));
  NOR2  g01768(.A(new_n2153_), .B(new_n847_), .Y(new_n2154_));
  NOR2  g01769(.A(new_n2154_), .B(new_n851_), .Y(new_n2155_));
  NOR2  g01770(.A(new_n2155_), .B(new_n856_), .Y(new_n2156_));
  NOR2  g01771(.A(new_n2156_), .B(new_n860_), .Y(new_n2157_));
  NOR2  g01772(.A(new_n2157_), .B(new_n865_), .Y(new_n2158_));
  NOR2  g01773(.A(new_n2158_), .B(new_n869_), .Y(new_n2159_));
  NOR2  g01774(.A(new_n2159_), .B(new_n874_), .Y(new_n2160_));
  NOR2  g01775(.A(new_n2160_), .B(new_n878_), .Y(new_n2161_));
  NOR2  g01776(.A(new_n2161_), .B(new_n883_), .Y(new_n2162_));
  NOR2  g01777(.A(new_n2162_), .B(new_n887_), .Y(new_n2163_));
  NOR2  g01778(.A(new_n2163_), .B(new_n892_), .Y(new_n2164_));
  NOR2  g01779(.A(new_n2164_), .B(new_n896_), .Y(new_n2165_));
  NOR2  g01780(.A(new_n2165_), .B(new_n901_), .Y(new_n2166_));
  NOR2  g01781(.A(new_n2166_), .B(new_n905_), .Y(new_n2167_));
  NOR2  g01782(.A(new_n2167_), .B(new_n910_), .Y(new_n2168_));
  NOR2  g01783(.A(new_n2168_), .B(new_n914_), .Y(new_n2169_));
  NOR2  g01784(.A(new_n2169_), .B(new_n919_), .Y(new_n2170_));
  NOR2  g01785(.A(new_n2170_), .B(new_n923_), .Y(new_n2171_));
  NOR2  g01786(.A(new_n2171_), .B(new_n928_), .Y(new_n2172_));
  NOR2  g01787(.A(new_n2172_), .B(new_n932_), .Y(new_n2173_));
  NOR2  g01788(.A(new_n2173_), .B(new_n937_), .Y(new_n2174_));
  NOR2  g01789(.A(new_n2174_), .B(new_n941_), .Y(new_n2175_));
  NOR2  g01790(.A(new_n2175_), .B(new_n946_), .Y(new_n2176_));
  NOR2  g01791(.A(new_n2176_), .B(new_n950_), .Y(new_n2177_));
  NOR2  g01792(.A(new_n2177_), .B(new_n955_), .Y(new_n2178_));
  NOR2  g01793(.A(new_n2178_), .B(new_n959_), .Y(new_n2179_));
  NOR2  g01794(.A(new_n2179_), .B(new_n964_), .Y(new_n2180_));
  NOR2  g01795(.A(new_n2180_), .B(new_n968_), .Y(new_n2181_));
  NOR2  g01796(.A(new_n2181_), .B(new_n973_), .Y(new_n2182_));
  NOR2  g01797(.A(new_n2182_), .B(new_n977_), .Y(new_n2183_));
  NOR2  g01798(.A(new_n2183_), .B(new_n982_), .Y(new_n2184_));
  NOR2  g01799(.A(new_n2184_), .B(new_n986_), .Y(new_n2185_));
  NOR2  g01800(.A(new_n2185_), .B(new_n991_), .Y(new_n2186_));
  NOR2  g01801(.A(new_n2186_), .B(new_n995_), .Y(new_n2187_));
  NOR2  g01802(.A(new_n2187_), .B(new_n1000_), .Y(new_n2188_));
  NOR2  g01803(.A(new_n2188_), .B(new_n1004_), .Y(new_n2189_));
  NOR2  g01804(.A(new_n2189_), .B(new_n1009_), .Y(new_n2190_));
  NOR2  g01805(.A(new_n2190_), .B(new_n1013_), .Y(new_n2191_));
  NOR2  g01806(.A(new_n2191_), .B(new_n1018_), .Y(new_n2192_));
  NOR2  g01807(.A(new_n2192_), .B(new_n1022_), .Y(new_n2193_));
  NOR2  g01808(.A(new_n2193_), .B(new_n1027_), .Y(new_n2194_));
  NOR2  g01809(.A(new_n2194_), .B(new_n1031_), .Y(new_n2195_));
  NOR2  g01810(.A(new_n2195_), .B(new_n1036_), .Y(new_n2196_));
  NOR2  g01811(.A(new_n2196_), .B(new_n1040_), .Y(new_n2197_));
  NOR2  g01812(.A(new_n2197_), .B(new_n1045_), .Y(new_n2198_));
  NOR2  g01813(.A(new_n2198_), .B(new_n1049_), .Y(new_n2199_));
  NOR2  g01814(.A(new_n2199_), .B(new_n1054_), .Y(new_n2200_));
  NOR2  g01815(.A(new_n2200_), .B(new_n1058_), .Y(new_n2201_));
  NOR2  g01816(.A(new_n2201_), .B(new_n1063_), .Y(new_n2202_));
  NOR2  g01817(.A(new_n2202_), .B(new_n1067_), .Y(new_n2203_));
  NOR2  g01818(.A(new_n2203_), .B(new_n1072_), .Y(new_n2204_));
  NOR2  g01819(.A(new_n2204_), .B(new_n1076_), .Y(new_n2205_));
  NOR2  g01820(.A(new_n2205_), .B(new_n1081_), .Y(new_n2206_));
  NOR2  g01821(.A(new_n2206_), .B(new_n1085_), .Y(new_n2207_));
  NOR2  g01822(.A(new_n2207_), .B(new_n1090_), .Y(new_n2208_));
  NOR2  g01823(.A(new_n2208_), .B(new_n1094_), .Y(new_n2209_));
  NOR2  g01824(.A(new_n2209_), .B(new_n1099_), .Y(new_n2210_));
  NOR2  g01825(.A(new_n2210_), .B(new_n1103_), .Y(new_n2211_));
  NOR2  g01826(.A(new_n2211_), .B(new_n1108_), .Y(new_n2212_));
  NOR2  g01827(.A(new_n2212_), .B(new_n1112_), .Y(new_n2213_));
  NOR2  g01828(.A(new_n2213_), .B(new_n1117_), .Y(new_n2214_));
  NOR2  g01829(.A(new_n2214_), .B(new_n1121_), .Y(new_n2215_));
  NOR2  g01830(.A(new_n2215_), .B(new_n1126_), .Y(new_n2216_));
  NOR2  g01831(.A(new_n2216_), .B(new_n1130_), .Y(new_n2217_));
  NOR2  g01832(.A(new_n2217_), .B(new_n1135_), .Y(new_n2218_));
  NOR2  g01833(.A(new_n2218_), .B(new_n1139_), .Y(new_n2219_));
  NOR2  g01834(.A(new_n2219_), .B(new_n1144_), .Y(new_n2220_));
  NOR2  g01835(.A(new_n2220_), .B(new_n1148_), .Y(new_n2221_));
  NOR2  g01836(.A(new_n2221_), .B(new_n1153_), .Y(new_n2222_));
  NOR2  g01837(.A(new_n2222_), .B(new_n1157_), .Y(new_n2223_));
  NOR2  g01838(.A(new_n2223_), .B(new_n1162_), .Y(new_n2224_));
  NOR2  g01839(.A(new_n2224_), .B(new_n1166_), .Y(new_n2225_));
  NOR2  g01840(.A(new_n2225_), .B(new_n1171_), .Y(new_n2226_));
  NOR2  g01841(.A(new_n2226_), .B(new_n1175_), .Y(new_n2227_));
  NOR2  g01842(.A(new_n2227_), .B(new_n1180_), .Y(new_n2228_));
  NOR2  g01843(.A(new_n2228_), .B(new_n1184_), .Y(new_n2229_));
  NOR2  g01844(.A(new_n2229_), .B(new_n1189_), .Y(new_n2230_));
  NOR2  g01845(.A(new_n2230_), .B(new_n1707_), .Y(new_n2231_));
  NOR2  g01846(.A(new_n2231_), .B(new_n1709_), .Y(new_n2232_));
  NOR2  g01847(.A(new_n2232_), .B(new_n1973_), .Y(new_n2233_));
  NOR2  g01848(.A(new_n2233_), .B(new_n1199_), .Y(new_n2234_));
  NOR2  g01849(.A(new_n2234_), .B(new_n1203_), .Y(new_n2235_));
  NOR2  g01850(.A(new_n2235_), .B(new_n1207_), .Y(new_n2236_));
  NAND2 g01851(.A(new_n1209_), .B(\req[10] ), .Y(new_n2237_));
  NOR2  g01852(.A(new_n2237_), .B(new_n2236_), .Y(\grant[10] ));
  INV   g01853(.A(new_n1218_), .Y(new_n2239_));
  NOR2  g01854(.A(new_n2239_), .B(new_n425_), .Y(new_n2240_));
  NOR2  g01855(.A(new_n2240_), .B(new_n1223_), .Y(new_n2241_));
  NOR2  g01856(.A(new_n2241_), .B(new_n1227_), .Y(new_n2242_));
  NOR2  g01857(.A(new_n2242_), .B(new_n1231_), .Y(new_n2243_));
  NOR2  g01858(.A(new_n2243_), .B(new_n1235_), .Y(new_n2244_));
  NOR2  g01859(.A(new_n2244_), .B(new_n1239_), .Y(new_n2245_));
  NOR2  g01860(.A(new_n2245_), .B(new_n1243_), .Y(new_n2246_));
  NOR2  g01861(.A(new_n2246_), .B(new_n1247_), .Y(new_n2247_));
  NOR2  g01862(.A(new_n2247_), .B(new_n1251_), .Y(new_n2248_));
  NOR2  g01863(.A(new_n2248_), .B(new_n1255_), .Y(new_n2249_));
  NOR2  g01864(.A(new_n2249_), .B(new_n1259_), .Y(new_n2250_));
  NOR2  g01865(.A(new_n2250_), .B(new_n1263_), .Y(new_n2251_));
  NOR2  g01866(.A(new_n2251_), .B(new_n1267_), .Y(new_n2252_));
  NOR2  g01867(.A(new_n2252_), .B(new_n1271_), .Y(new_n2253_));
  NOR2  g01868(.A(new_n2253_), .B(new_n1275_), .Y(new_n2254_));
  NOR2  g01869(.A(new_n2254_), .B(new_n1279_), .Y(new_n2255_));
  NOR2  g01870(.A(new_n2255_), .B(new_n1283_), .Y(new_n2256_));
  NOR2  g01871(.A(new_n2256_), .B(new_n1287_), .Y(new_n2257_));
  NOR2  g01872(.A(new_n2257_), .B(new_n1291_), .Y(new_n2258_));
  NOR2  g01873(.A(new_n2258_), .B(new_n1295_), .Y(new_n2259_));
  NOR2  g01874(.A(new_n2259_), .B(new_n1299_), .Y(new_n2260_));
  NOR2  g01875(.A(new_n2260_), .B(new_n1303_), .Y(new_n2261_));
  NOR2  g01876(.A(new_n2261_), .B(new_n1307_), .Y(new_n2262_));
  NOR2  g01877(.A(new_n2262_), .B(new_n1311_), .Y(new_n2263_));
  NOR2  g01878(.A(new_n2263_), .B(new_n1315_), .Y(new_n2264_));
  NOR2  g01879(.A(new_n2264_), .B(new_n1319_), .Y(new_n2265_));
  NOR2  g01880(.A(new_n2265_), .B(new_n1323_), .Y(new_n2266_));
  NOR2  g01881(.A(new_n2266_), .B(new_n1327_), .Y(new_n2267_));
  NOR2  g01882(.A(new_n2267_), .B(new_n1331_), .Y(new_n2268_));
  NOR2  g01883(.A(new_n2268_), .B(new_n1335_), .Y(new_n2269_));
  NOR2  g01884(.A(new_n2269_), .B(new_n1339_), .Y(new_n2270_));
  NOR2  g01885(.A(new_n2270_), .B(new_n1343_), .Y(new_n2271_));
  NOR2  g01886(.A(new_n2271_), .B(new_n1347_), .Y(new_n2272_));
  NOR2  g01887(.A(new_n2272_), .B(new_n1351_), .Y(new_n2273_));
  NOR2  g01888(.A(new_n2273_), .B(new_n1355_), .Y(new_n2274_));
  NOR2  g01889(.A(new_n2274_), .B(new_n1359_), .Y(new_n2275_));
  NOR2  g01890(.A(new_n2275_), .B(new_n1363_), .Y(new_n2276_));
  NOR2  g01891(.A(new_n2276_), .B(new_n1367_), .Y(new_n2277_));
  NOR2  g01892(.A(new_n2277_), .B(new_n1371_), .Y(new_n2278_));
  NOR2  g01893(.A(new_n2278_), .B(new_n1375_), .Y(new_n2279_));
  NOR2  g01894(.A(new_n2279_), .B(new_n1379_), .Y(new_n2280_));
  NOR2  g01895(.A(new_n2280_), .B(new_n1383_), .Y(new_n2281_));
  NOR2  g01896(.A(new_n2281_), .B(new_n1387_), .Y(new_n2282_));
  NOR2  g01897(.A(new_n2282_), .B(new_n1391_), .Y(new_n2283_));
  NOR2  g01898(.A(new_n2283_), .B(new_n1395_), .Y(new_n2284_));
  NOR2  g01899(.A(new_n2284_), .B(new_n1399_), .Y(new_n2285_));
  NOR2  g01900(.A(new_n2285_), .B(new_n1403_), .Y(new_n2286_));
  NOR2  g01901(.A(new_n2286_), .B(new_n1407_), .Y(new_n2287_));
  NOR2  g01902(.A(new_n2287_), .B(new_n1411_), .Y(new_n2288_));
  NOR2  g01903(.A(new_n2288_), .B(new_n1415_), .Y(new_n2289_));
  NOR2  g01904(.A(new_n2289_), .B(new_n1419_), .Y(new_n2290_));
  NOR2  g01905(.A(new_n2290_), .B(new_n1423_), .Y(new_n2291_));
  NOR2  g01906(.A(new_n2291_), .B(new_n1427_), .Y(new_n2292_));
  NOR2  g01907(.A(new_n2292_), .B(new_n1431_), .Y(new_n2293_));
  NOR2  g01908(.A(new_n2293_), .B(new_n1435_), .Y(new_n2294_));
  NOR2  g01909(.A(new_n2294_), .B(new_n1439_), .Y(new_n2295_));
  NOR2  g01910(.A(new_n2295_), .B(new_n1443_), .Y(new_n2296_));
  NOR2  g01911(.A(new_n2296_), .B(new_n1447_), .Y(new_n2297_));
  NOR2  g01912(.A(new_n2297_), .B(new_n1451_), .Y(new_n2298_));
  NOR2  g01913(.A(new_n2298_), .B(new_n1455_), .Y(new_n2299_));
  NOR2  g01914(.A(new_n2299_), .B(new_n1459_), .Y(new_n2300_));
  NOR2  g01915(.A(new_n2300_), .B(new_n1463_), .Y(new_n2301_));
  NOR2  g01916(.A(new_n2301_), .B(new_n1467_), .Y(new_n2302_));
  NOR2  g01917(.A(new_n2302_), .B(new_n1471_), .Y(new_n2303_));
  NOR2  g01918(.A(new_n2303_), .B(new_n1475_), .Y(new_n2304_));
  NOR2  g01919(.A(new_n2304_), .B(new_n1479_), .Y(new_n2305_));
  NOR2  g01920(.A(new_n2305_), .B(new_n1483_), .Y(new_n2306_));
  NOR2  g01921(.A(new_n2306_), .B(new_n1487_), .Y(new_n2307_));
  NOR2  g01922(.A(new_n2307_), .B(new_n1491_), .Y(new_n2308_));
  NOR2  g01923(.A(new_n2308_), .B(new_n1495_), .Y(new_n2309_));
  NOR2  g01924(.A(new_n2309_), .B(new_n1499_), .Y(new_n2310_));
  NOR2  g01925(.A(new_n2310_), .B(new_n1503_), .Y(new_n2311_));
  NOR2  g01926(.A(new_n2311_), .B(new_n1507_), .Y(new_n2312_));
  NOR2  g01927(.A(new_n2312_), .B(new_n1511_), .Y(new_n2313_));
  NOR2  g01928(.A(new_n2313_), .B(new_n1515_), .Y(new_n2314_));
  NOR2  g01929(.A(new_n2314_), .B(new_n1519_), .Y(new_n2315_));
  NOR2  g01930(.A(new_n2315_), .B(new_n1523_), .Y(new_n2316_));
  NOR2  g01931(.A(new_n2316_), .B(new_n1527_), .Y(new_n2317_));
  NOR2  g01932(.A(new_n2317_), .B(new_n1797_), .Y(new_n2318_));
  NOR2  g01933(.A(new_n2318_), .B(new_n396_), .Y(new_n2319_));
  NOR2  g01934(.A(new_n2319_), .B(new_n400_), .Y(new_n2320_));
  NOR2  g01935(.A(new_n2320_), .B(new_n406_), .Y(new_n2321_));
  NOR2  g01936(.A(new_n2321_), .B(new_n410_), .Y(new_n2322_));
  NOR2  g01937(.A(new_n2322_), .B(new_n416_), .Y(new_n2323_));
  NAND2 g01938(.A(new_n418_), .B(\req[11] ), .Y(new_n2324_));
  NOR2  g01939(.A(new_n2324_), .B(new_n2323_), .Y(\grant[11] ));
  INV   g01940(.A(new_n429_), .Y(new_n2326_));
  NOR2  g01941(.A(new_n846_), .B(new_n2326_), .Y(new_n2327_));
  NOR2  g01942(.A(new_n2327_), .B(new_n436_), .Y(new_n2328_));
  NOR2  g01943(.A(new_n2328_), .B(new_n440_), .Y(new_n2329_));
  NOR2  g01944(.A(new_n2329_), .B(new_n446_), .Y(new_n2330_));
  NOR2  g01945(.A(new_n2330_), .B(new_n450_), .Y(new_n2331_));
  NOR2  g01946(.A(new_n2331_), .B(new_n456_), .Y(new_n2332_));
  NOR2  g01947(.A(new_n2332_), .B(new_n460_), .Y(new_n2333_));
  NOR2  g01948(.A(new_n2333_), .B(new_n466_), .Y(new_n2334_));
  NOR2  g01949(.A(new_n2334_), .B(new_n470_), .Y(new_n2335_));
  NOR2  g01950(.A(new_n2335_), .B(new_n476_), .Y(new_n2336_));
  NOR2  g01951(.A(new_n2336_), .B(new_n480_), .Y(new_n2337_));
  NOR2  g01952(.A(new_n2337_), .B(new_n486_), .Y(new_n2338_));
  NOR2  g01953(.A(new_n2338_), .B(new_n490_), .Y(new_n2339_));
  NOR2  g01954(.A(new_n2339_), .B(new_n496_), .Y(new_n2340_));
  NOR2  g01955(.A(new_n2340_), .B(new_n500_), .Y(new_n2341_));
  NOR2  g01956(.A(new_n2341_), .B(new_n506_), .Y(new_n2342_));
  NOR2  g01957(.A(new_n2342_), .B(new_n510_), .Y(new_n2343_));
  NOR2  g01958(.A(new_n2343_), .B(new_n516_), .Y(new_n2344_));
  NOR2  g01959(.A(new_n2344_), .B(new_n520_), .Y(new_n2345_));
  NOR2  g01960(.A(new_n2345_), .B(new_n526_), .Y(new_n2346_));
  NOR2  g01961(.A(new_n2346_), .B(new_n530_), .Y(new_n2347_));
  NOR2  g01962(.A(new_n2347_), .B(new_n536_), .Y(new_n2348_));
  NOR2  g01963(.A(new_n2348_), .B(new_n540_), .Y(new_n2349_));
  NOR2  g01964(.A(new_n2349_), .B(new_n546_), .Y(new_n2350_));
  NOR2  g01965(.A(new_n2350_), .B(new_n550_), .Y(new_n2351_));
  NOR2  g01966(.A(new_n2351_), .B(new_n556_), .Y(new_n2352_));
  NOR2  g01967(.A(new_n2352_), .B(new_n560_), .Y(new_n2353_));
  NOR2  g01968(.A(new_n2353_), .B(new_n566_), .Y(new_n2354_));
  NOR2  g01969(.A(new_n2354_), .B(new_n570_), .Y(new_n2355_));
  NOR2  g01970(.A(new_n2355_), .B(new_n576_), .Y(new_n2356_));
  NOR2  g01971(.A(new_n2356_), .B(new_n580_), .Y(new_n2357_));
  NOR2  g01972(.A(new_n2357_), .B(new_n586_), .Y(new_n2358_));
  NOR2  g01973(.A(new_n2358_), .B(new_n590_), .Y(new_n2359_));
  NOR2  g01974(.A(new_n2359_), .B(new_n596_), .Y(new_n2360_));
  NOR2  g01975(.A(new_n2360_), .B(new_n600_), .Y(new_n2361_));
  NOR2  g01976(.A(new_n2361_), .B(new_n606_), .Y(new_n2362_));
  NOR2  g01977(.A(new_n2362_), .B(new_n610_), .Y(new_n2363_));
  NOR2  g01978(.A(new_n2363_), .B(new_n616_), .Y(new_n2364_));
  NOR2  g01979(.A(new_n2364_), .B(new_n620_), .Y(new_n2365_));
  NOR2  g01980(.A(new_n2365_), .B(new_n626_), .Y(new_n2366_));
  NOR2  g01981(.A(new_n2366_), .B(new_n630_), .Y(new_n2367_));
  NOR2  g01982(.A(new_n2367_), .B(new_n636_), .Y(new_n2368_));
  NOR2  g01983(.A(new_n2368_), .B(new_n640_), .Y(new_n2369_));
  NOR2  g01984(.A(new_n2369_), .B(new_n646_), .Y(new_n2370_));
  NOR2  g01985(.A(new_n2370_), .B(new_n650_), .Y(new_n2371_));
  NOR2  g01986(.A(new_n2371_), .B(new_n656_), .Y(new_n2372_));
  NOR2  g01987(.A(new_n2372_), .B(new_n660_), .Y(new_n2373_));
  NOR2  g01988(.A(new_n2373_), .B(new_n666_), .Y(new_n2374_));
  NOR2  g01989(.A(new_n2374_), .B(new_n670_), .Y(new_n2375_));
  NOR2  g01990(.A(new_n2375_), .B(new_n676_), .Y(new_n2376_));
  NOR2  g01991(.A(new_n2376_), .B(new_n680_), .Y(new_n2377_));
  NOR2  g01992(.A(new_n2377_), .B(new_n686_), .Y(new_n2378_));
  NOR2  g01993(.A(new_n2378_), .B(new_n690_), .Y(new_n2379_));
  NOR2  g01994(.A(new_n2379_), .B(new_n696_), .Y(new_n2380_));
  NOR2  g01995(.A(new_n2380_), .B(new_n700_), .Y(new_n2381_));
  NOR2  g01996(.A(new_n2381_), .B(new_n706_), .Y(new_n2382_));
  NOR2  g01997(.A(new_n2382_), .B(new_n710_), .Y(new_n2383_));
  NOR2  g01998(.A(new_n2383_), .B(new_n716_), .Y(new_n2384_));
  NOR2  g01999(.A(new_n2384_), .B(new_n720_), .Y(new_n2385_));
  NOR2  g02000(.A(new_n2385_), .B(new_n726_), .Y(new_n2386_));
  NOR2  g02001(.A(new_n2386_), .B(new_n730_), .Y(new_n2387_));
  NOR2  g02002(.A(new_n2387_), .B(new_n736_), .Y(new_n2388_));
  NOR2  g02003(.A(new_n2388_), .B(new_n740_), .Y(new_n2389_));
  NOR2  g02004(.A(new_n2389_), .B(new_n746_), .Y(new_n2390_));
  NOR2  g02005(.A(new_n2390_), .B(new_n750_), .Y(new_n2391_));
  NOR2  g02006(.A(new_n2391_), .B(new_n756_), .Y(new_n2392_));
  NOR2  g02007(.A(new_n2392_), .B(new_n760_), .Y(new_n2393_));
  NOR2  g02008(.A(new_n2393_), .B(new_n766_), .Y(new_n2394_));
  NOR2  g02009(.A(new_n2394_), .B(new_n770_), .Y(new_n2395_));
  NOR2  g02010(.A(new_n2395_), .B(new_n776_), .Y(new_n2396_));
  NOR2  g02011(.A(new_n2396_), .B(new_n780_), .Y(new_n2397_));
  NOR2  g02012(.A(new_n2397_), .B(new_n786_), .Y(new_n2398_));
  NOR2  g02013(.A(new_n2398_), .B(new_n790_), .Y(new_n2399_));
  NOR2  g02014(.A(new_n2399_), .B(new_n796_), .Y(new_n2400_));
  NOR2  g02015(.A(new_n2400_), .B(new_n800_), .Y(new_n2401_));
  NOR2  g02016(.A(new_n2401_), .B(new_n806_), .Y(new_n2402_));
  NOR2  g02017(.A(new_n2402_), .B(new_n1616_), .Y(new_n2403_));
  NOR2  g02018(.A(new_n2403_), .B(new_n1618_), .Y(new_n2404_));
  NOR2  g02019(.A(new_n2404_), .B(new_n1885_), .Y(new_n2405_));
  NOR2  g02020(.A(new_n2405_), .B(new_n820_), .Y(new_n2406_));
  NOR2  g02021(.A(new_n2406_), .B(new_n824_), .Y(new_n2407_));
  NOR2  g02022(.A(new_n2407_), .B(new_n829_), .Y(new_n2408_));
  NOR2  g02023(.A(new_n2408_), .B(new_n833_), .Y(new_n2409_));
  NOR2  g02024(.A(new_n2409_), .B(new_n838_), .Y(new_n2410_));
  NAND2 g02025(.A(new_n840_), .B(\req[12] ), .Y(new_n2411_));
  NOR2  g02026(.A(new_n2411_), .B(new_n2410_), .Y(\grant[12] ));
  INV   g02027(.A(new_n850_), .Y(new_n2413_));
  NOR2  g02028(.A(new_n1222_), .B(new_n2413_), .Y(new_n2414_));
  NOR2  g02029(.A(new_n2414_), .B(new_n856_), .Y(new_n2415_));
  NOR2  g02030(.A(new_n2415_), .B(new_n860_), .Y(new_n2416_));
  NOR2  g02031(.A(new_n2416_), .B(new_n865_), .Y(new_n2417_));
  NOR2  g02032(.A(new_n2417_), .B(new_n869_), .Y(new_n2418_));
  NOR2  g02033(.A(new_n2418_), .B(new_n874_), .Y(new_n2419_));
  NOR2  g02034(.A(new_n2419_), .B(new_n878_), .Y(new_n2420_));
  NOR2  g02035(.A(new_n2420_), .B(new_n883_), .Y(new_n2421_));
  NOR2  g02036(.A(new_n2421_), .B(new_n887_), .Y(new_n2422_));
  NOR2  g02037(.A(new_n2422_), .B(new_n892_), .Y(new_n2423_));
  NOR2  g02038(.A(new_n2423_), .B(new_n896_), .Y(new_n2424_));
  NOR2  g02039(.A(new_n2424_), .B(new_n901_), .Y(new_n2425_));
  NOR2  g02040(.A(new_n2425_), .B(new_n905_), .Y(new_n2426_));
  NOR2  g02041(.A(new_n2426_), .B(new_n910_), .Y(new_n2427_));
  NOR2  g02042(.A(new_n2427_), .B(new_n914_), .Y(new_n2428_));
  NOR2  g02043(.A(new_n2428_), .B(new_n919_), .Y(new_n2429_));
  NOR2  g02044(.A(new_n2429_), .B(new_n923_), .Y(new_n2430_));
  NOR2  g02045(.A(new_n2430_), .B(new_n928_), .Y(new_n2431_));
  NOR2  g02046(.A(new_n2431_), .B(new_n932_), .Y(new_n2432_));
  NOR2  g02047(.A(new_n2432_), .B(new_n937_), .Y(new_n2433_));
  NOR2  g02048(.A(new_n2433_), .B(new_n941_), .Y(new_n2434_));
  NOR2  g02049(.A(new_n2434_), .B(new_n946_), .Y(new_n2435_));
  NOR2  g02050(.A(new_n2435_), .B(new_n950_), .Y(new_n2436_));
  NOR2  g02051(.A(new_n2436_), .B(new_n955_), .Y(new_n2437_));
  NOR2  g02052(.A(new_n2437_), .B(new_n959_), .Y(new_n2438_));
  NOR2  g02053(.A(new_n2438_), .B(new_n964_), .Y(new_n2439_));
  NOR2  g02054(.A(new_n2439_), .B(new_n968_), .Y(new_n2440_));
  NOR2  g02055(.A(new_n2440_), .B(new_n973_), .Y(new_n2441_));
  NOR2  g02056(.A(new_n2441_), .B(new_n977_), .Y(new_n2442_));
  NOR2  g02057(.A(new_n2442_), .B(new_n982_), .Y(new_n2443_));
  NOR2  g02058(.A(new_n2443_), .B(new_n986_), .Y(new_n2444_));
  NOR2  g02059(.A(new_n2444_), .B(new_n991_), .Y(new_n2445_));
  NOR2  g02060(.A(new_n2445_), .B(new_n995_), .Y(new_n2446_));
  NOR2  g02061(.A(new_n2446_), .B(new_n1000_), .Y(new_n2447_));
  NOR2  g02062(.A(new_n2447_), .B(new_n1004_), .Y(new_n2448_));
  NOR2  g02063(.A(new_n2448_), .B(new_n1009_), .Y(new_n2449_));
  NOR2  g02064(.A(new_n2449_), .B(new_n1013_), .Y(new_n2450_));
  NOR2  g02065(.A(new_n2450_), .B(new_n1018_), .Y(new_n2451_));
  NOR2  g02066(.A(new_n2451_), .B(new_n1022_), .Y(new_n2452_));
  NOR2  g02067(.A(new_n2452_), .B(new_n1027_), .Y(new_n2453_));
  NOR2  g02068(.A(new_n2453_), .B(new_n1031_), .Y(new_n2454_));
  NOR2  g02069(.A(new_n2454_), .B(new_n1036_), .Y(new_n2455_));
  NOR2  g02070(.A(new_n2455_), .B(new_n1040_), .Y(new_n2456_));
  NOR2  g02071(.A(new_n2456_), .B(new_n1045_), .Y(new_n2457_));
  NOR2  g02072(.A(new_n2457_), .B(new_n1049_), .Y(new_n2458_));
  NOR2  g02073(.A(new_n2458_), .B(new_n1054_), .Y(new_n2459_));
  NOR2  g02074(.A(new_n2459_), .B(new_n1058_), .Y(new_n2460_));
  NOR2  g02075(.A(new_n2460_), .B(new_n1063_), .Y(new_n2461_));
  NOR2  g02076(.A(new_n2461_), .B(new_n1067_), .Y(new_n2462_));
  NOR2  g02077(.A(new_n2462_), .B(new_n1072_), .Y(new_n2463_));
  NOR2  g02078(.A(new_n2463_), .B(new_n1076_), .Y(new_n2464_));
  NOR2  g02079(.A(new_n2464_), .B(new_n1081_), .Y(new_n2465_));
  NOR2  g02080(.A(new_n2465_), .B(new_n1085_), .Y(new_n2466_));
  NOR2  g02081(.A(new_n2466_), .B(new_n1090_), .Y(new_n2467_));
  NOR2  g02082(.A(new_n2467_), .B(new_n1094_), .Y(new_n2468_));
  NOR2  g02083(.A(new_n2468_), .B(new_n1099_), .Y(new_n2469_));
  NOR2  g02084(.A(new_n2469_), .B(new_n1103_), .Y(new_n2470_));
  NOR2  g02085(.A(new_n2470_), .B(new_n1108_), .Y(new_n2471_));
  NOR2  g02086(.A(new_n2471_), .B(new_n1112_), .Y(new_n2472_));
  NOR2  g02087(.A(new_n2472_), .B(new_n1117_), .Y(new_n2473_));
  NOR2  g02088(.A(new_n2473_), .B(new_n1121_), .Y(new_n2474_));
  NOR2  g02089(.A(new_n2474_), .B(new_n1126_), .Y(new_n2475_));
  NOR2  g02090(.A(new_n2475_), .B(new_n1130_), .Y(new_n2476_));
  NOR2  g02091(.A(new_n2476_), .B(new_n1135_), .Y(new_n2477_));
  NOR2  g02092(.A(new_n2477_), .B(new_n1139_), .Y(new_n2478_));
  NOR2  g02093(.A(new_n2478_), .B(new_n1144_), .Y(new_n2479_));
  NOR2  g02094(.A(new_n2479_), .B(new_n1148_), .Y(new_n2480_));
  NOR2  g02095(.A(new_n2480_), .B(new_n1153_), .Y(new_n2481_));
  NOR2  g02096(.A(new_n2481_), .B(new_n1157_), .Y(new_n2482_));
  NOR2  g02097(.A(new_n2482_), .B(new_n1162_), .Y(new_n2483_));
  NOR2  g02098(.A(new_n2483_), .B(new_n1166_), .Y(new_n2484_));
  NOR2  g02099(.A(new_n2484_), .B(new_n1171_), .Y(new_n2485_));
  NOR2  g02100(.A(new_n2485_), .B(new_n1175_), .Y(new_n2486_));
  NOR2  g02101(.A(new_n2486_), .B(new_n1180_), .Y(new_n2487_));
  NOR2  g02102(.A(new_n2487_), .B(new_n1184_), .Y(new_n2488_));
  NOR2  g02103(.A(new_n2488_), .B(new_n1189_), .Y(new_n2489_));
  NOR2  g02104(.A(new_n2489_), .B(new_n1707_), .Y(new_n2490_));
  NOR2  g02105(.A(new_n2490_), .B(new_n1709_), .Y(new_n2491_));
  NOR2  g02106(.A(new_n2491_), .B(new_n1973_), .Y(new_n2492_));
  NOR2  g02107(.A(new_n2492_), .B(new_n1199_), .Y(new_n2493_));
  NOR2  g02108(.A(new_n2493_), .B(new_n1203_), .Y(new_n2494_));
  NOR2  g02109(.A(new_n2494_), .B(new_n1207_), .Y(new_n2495_));
  NOR2  g02110(.A(new_n2495_), .B(new_n1211_), .Y(new_n2496_));
  NOR2  g02111(.A(new_n2496_), .B(new_n1215_), .Y(new_n2497_));
  NAND2 g02112(.A(new_n1217_), .B(\req[13] ), .Y(new_n2498_));
  NOR2  g02113(.A(new_n2498_), .B(new_n2497_), .Y(\grant[13] ));
  INV   g02114(.A(new_n1226_), .Y(new_n2500_));
  NOR2  g02115(.A(new_n2500_), .B(new_n435_), .Y(new_n2501_));
  NOR2  g02116(.A(new_n2501_), .B(new_n1231_), .Y(new_n2502_));
  NOR2  g02117(.A(new_n2502_), .B(new_n1235_), .Y(new_n2503_));
  NOR2  g02118(.A(new_n2503_), .B(new_n1239_), .Y(new_n2504_));
  NOR2  g02119(.A(new_n2504_), .B(new_n1243_), .Y(new_n2505_));
  NOR2  g02120(.A(new_n2505_), .B(new_n1247_), .Y(new_n2506_));
  NOR2  g02121(.A(new_n2506_), .B(new_n1251_), .Y(new_n2507_));
  NOR2  g02122(.A(new_n2507_), .B(new_n1255_), .Y(new_n2508_));
  NOR2  g02123(.A(new_n2508_), .B(new_n1259_), .Y(new_n2509_));
  NOR2  g02124(.A(new_n2509_), .B(new_n1263_), .Y(new_n2510_));
  NOR2  g02125(.A(new_n2510_), .B(new_n1267_), .Y(new_n2511_));
  NOR2  g02126(.A(new_n2511_), .B(new_n1271_), .Y(new_n2512_));
  NOR2  g02127(.A(new_n2512_), .B(new_n1275_), .Y(new_n2513_));
  NOR2  g02128(.A(new_n2513_), .B(new_n1279_), .Y(new_n2514_));
  NOR2  g02129(.A(new_n2514_), .B(new_n1283_), .Y(new_n2515_));
  NOR2  g02130(.A(new_n2515_), .B(new_n1287_), .Y(new_n2516_));
  NOR2  g02131(.A(new_n2516_), .B(new_n1291_), .Y(new_n2517_));
  NOR2  g02132(.A(new_n2517_), .B(new_n1295_), .Y(new_n2518_));
  NOR2  g02133(.A(new_n2518_), .B(new_n1299_), .Y(new_n2519_));
  NOR2  g02134(.A(new_n2519_), .B(new_n1303_), .Y(new_n2520_));
  NOR2  g02135(.A(new_n2520_), .B(new_n1307_), .Y(new_n2521_));
  NOR2  g02136(.A(new_n2521_), .B(new_n1311_), .Y(new_n2522_));
  NOR2  g02137(.A(new_n2522_), .B(new_n1315_), .Y(new_n2523_));
  NOR2  g02138(.A(new_n2523_), .B(new_n1319_), .Y(new_n2524_));
  NOR2  g02139(.A(new_n2524_), .B(new_n1323_), .Y(new_n2525_));
  NOR2  g02140(.A(new_n2525_), .B(new_n1327_), .Y(new_n2526_));
  NOR2  g02141(.A(new_n2526_), .B(new_n1331_), .Y(new_n2527_));
  NOR2  g02142(.A(new_n2527_), .B(new_n1335_), .Y(new_n2528_));
  NOR2  g02143(.A(new_n2528_), .B(new_n1339_), .Y(new_n2529_));
  NOR2  g02144(.A(new_n2529_), .B(new_n1343_), .Y(new_n2530_));
  NOR2  g02145(.A(new_n2530_), .B(new_n1347_), .Y(new_n2531_));
  NOR2  g02146(.A(new_n2531_), .B(new_n1351_), .Y(new_n2532_));
  NOR2  g02147(.A(new_n2532_), .B(new_n1355_), .Y(new_n2533_));
  NOR2  g02148(.A(new_n2533_), .B(new_n1359_), .Y(new_n2534_));
  NOR2  g02149(.A(new_n2534_), .B(new_n1363_), .Y(new_n2535_));
  NOR2  g02150(.A(new_n2535_), .B(new_n1367_), .Y(new_n2536_));
  NOR2  g02151(.A(new_n2536_), .B(new_n1371_), .Y(new_n2537_));
  NOR2  g02152(.A(new_n2537_), .B(new_n1375_), .Y(new_n2538_));
  NOR2  g02153(.A(new_n2538_), .B(new_n1379_), .Y(new_n2539_));
  NOR2  g02154(.A(new_n2539_), .B(new_n1383_), .Y(new_n2540_));
  NOR2  g02155(.A(new_n2540_), .B(new_n1387_), .Y(new_n2541_));
  NOR2  g02156(.A(new_n2541_), .B(new_n1391_), .Y(new_n2542_));
  NOR2  g02157(.A(new_n2542_), .B(new_n1395_), .Y(new_n2543_));
  NOR2  g02158(.A(new_n2543_), .B(new_n1399_), .Y(new_n2544_));
  NOR2  g02159(.A(new_n2544_), .B(new_n1403_), .Y(new_n2545_));
  NOR2  g02160(.A(new_n2545_), .B(new_n1407_), .Y(new_n2546_));
  NOR2  g02161(.A(new_n2546_), .B(new_n1411_), .Y(new_n2547_));
  NOR2  g02162(.A(new_n2547_), .B(new_n1415_), .Y(new_n2548_));
  NOR2  g02163(.A(new_n2548_), .B(new_n1419_), .Y(new_n2549_));
  NOR2  g02164(.A(new_n2549_), .B(new_n1423_), .Y(new_n2550_));
  NOR2  g02165(.A(new_n2550_), .B(new_n1427_), .Y(new_n2551_));
  NOR2  g02166(.A(new_n2551_), .B(new_n1431_), .Y(new_n2552_));
  NOR2  g02167(.A(new_n2552_), .B(new_n1435_), .Y(new_n2553_));
  NOR2  g02168(.A(new_n2553_), .B(new_n1439_), .Y(new_n2554_));
  NOR2  g02169(.A(new_n2554_), .B(new_n1443_), .Y(new_n2555_));
  NOR2  g02170(.A(new_n2555_), .B(new_n1447_), .Y(new_n2556_));
  NOR2  g02171(.A(new_n2556_), .B(new_n1451_), .Y(new_n2557_));
  NOR2  g02172(.A(new_n2557_), .B(new_n1455_), .Y(new_n2558_));
  NOR2  g02173(.A(new_n2558_), .B(new_n1459_), .Y(new_n2559_));
  NOR2  g02174(.A(new_n2559_), .B(new_n1463_), .Y(new_n2560_));
  NOR2  g02175(.A(new_n2560_), .B(new_n1467_), .Y(new_n2561_));
  NOR2  g02176(.A(new_n2561_), .B(new_n1471_), .Y(new_n2562_));
  NOR2  g02177(.A(new_n2562_), .B(new_n1475_), .Y(new_n2563_));
  NOR2  g02178(.A(new_n2563_), .B(new_n1479_), .Y(new_n2564_));
  NOR2  g02179(.A(new_n2564_), .B(new_n1483_), .Y(new_n2565_));
  NOR2  g02180(.A(new_n2565_), .B(new_n1487_), .Y(new_n2566_));
  NOR2  g02181(.A(new_n2566_), .B(new_n1491_), .Y(new_n2567_));
  NOR2  g02182(.A(new_n2567_), .B(new_n1495_), .Y(new_n2568_));
  NOR2  g02183(.A(new_n2568_), .B(new_n1499_), .Y(new_n2569_));
  NOR2  g02184(.A(new_n2569_), .B(new_n1503_), .Y(new_n2570_));
  NOR2  g02185(.A(new_n2570_), .B(new_n1507_), .Y(new_n2571_));
  NOR2  g02186(.A(new_n2571_), .B(new_n1511_), .Y(new_n2572_));
  NOR2  g02187(.A(new_n2572_), .B(new_n1515_), .Y(new_n2573_));
  NOR2  g02188(.A(new_n2573_), .B(new_n1519_), .Y(new_n2574_));
  NOR2  g02189(.A(new_n2574_), .B(new_n1523_), .Y(new_n2575_));
  NOR2  g02190(.A(new_n2575_), .B(new_n1527_), .Y(new_n2576_));
  NOR2  g02191(.A(new_n2576_), .B(new_n1797_), .Y(new_n2577_));
  NOR2  g02192(.A(new_n2577_), .B(new_n396_), .Y(new_n2578_));
  NOR2  g02193(.A(new_n2578_), .B(new_n400_), .Y(new_n2579_));
  NOR2  g02194(.A(new_n2579_), .B(new_n406_), .Y(new_n2580_));
  NOR2  g02195(.A(new_n2580_), .B(new_n410_), .Y(new_n2581_));
  NOR2  g02196(.A(new_n2581_), .B(new_n416_), .Y(new_n2582_));
  NOR2  g02197(.A(new_n2582_), .B(new_n420_), .Y(new_n2583_));
  NOR2  g02198(.A(new_n2583_), .B(new_n426_), .Y(new_n2584_));
  NAND2 g02199(.A(new_n428_), .B(\req[14] ), .Y(new_n2585_));
  NOR2  g02200(.A(new_n2585_), .B(new_n2584_), .Y(\grant[14] ));
  INV   g02201(.A(new_n439_), .Y(new_n2587_));
  NOR2  g02202(.A(new_n855_), .B(new_n2587_), .Y(new_n2588_));
  NOR2  g02203(.A(new_n2588_), .B(new_n446_), .Y(new_n2589_));
  NOR2  g02204(.A(new_n2589_), .B(new_n450_), .Y(new_n2590_));
  NOR2  g02205(.A(new_n2590_), .B(new_n456_), .Y(new_n2591_));
  NOR2  g02206(.A(new_n2591_), .B(new_n460_), .Y(new_n2592_));
  NOR2  g02207(.A(new_n2592_), .B(new_n466_), .Y(new_n2593_));
  NOR2  g02208(.A(new_n2593_), .B(new_n470_), .Y(new_n2594_));
  NOR2  g02209(.A(new_n2594_), .B(new_n476_), .Y(new_n2595_));
  NOR2  g02210(.A(new_n2595_), .B(new_n480_), .Y(new_n2596_));
  NOR2  g02211(.A(new_n2596_), .B(new_n486_), .Y(new_n2597_));
  NOR2  g02212(.A(new_n2597_), .B(new_n490_), .Y(new_n2598_));
  NOR2  g02213(.A(new_n2598_), .B(new_n496_), .Y(new_n2599_));
  NOR2  g02214(.A(new_n2599_), .B(new_n500_), .Y(new_n2600_));
  NOR2  g02215(.A(new_n2600_), .B(new_n506_), .Y(new_n2601_));
  NOR2  g02216(.A(new_n2601_), .B(new_n510_), .Y(new_n2602_));
  NOR2  g02217(.A(new_n2602_), .B(new_n516_), .Y(new_n2603_));
  NOR2  g02218(.A(new_n2603_), .B(new_n520_), .Y(new_n2604_));
  NOR2  g02219(.A(new_n2604_), .B(new_n526_), .Y(new_n2605_));
  NOR2  g02220(.A(new_n2605_), .B(new_n530_), .Y(new_n2606_));
  NOR2  g02221(.A(new_n2606_), .B(new_n536_), .Y(new_n2607_));
  NOR2  g02222(.A(new_n2607_), .B(new_n540_), .Y(new_n2608_));
  NOR2  g02223(.A(new_n2608_), .B(new_n546_), .Y(new_n2609_));
  NOR2  g02224(.A(new_n2609_), .B(new_n550_), .Y(new_n2610_));
  NOR2  g02225(.A(new_n2610_), .B(new_n556_), .Y(new_n2611_));
  NOR2  g02226(.A(new_n2611_), .B(new_n560_), .Y(new_n2612_));
  NOR2  g02227(.A(new_n2612_), .B(new_n566_), .Y(new_n2613_));
  NOR2  g02228(.A(new_n2613_), .B(new_n570_), .Y(new_n2614_));
  NOR2  g02229(.A(new_n2614_), .B(new_n576_), .Y(new_n2615_));
  NOR2  g02230(.A(new_n2615_), .B(new_n580_), .Y(new_n2616_));
  NOR2  g02231(.A(new_n2616_), .B(new_n586_), .Y(new_n2617_));
  NOR2  g02232(.A(new_n2617_), .B(new_n590_), .Y(new_n2618_));
  NOR2  g02233(.A(new_n2618_), .B(new_n596_), .Y(new_n2619_));
  NOR2  g02234(.A(new_n2619_), .B(new_n600_), .Y(new_n2620_));
  NOR2  g02235(.A(new_n2620_), .B(new_n606_), .Y(new_n2621_));
  NOR2  g02236(.A(new_n2621_), .B(new_n610_), .Y(new_n2622_));
  NOR2  g02237(.A(new_n2622_), .B(new_n616_), .Y(new_n2623_));
  NOR2  g02238(.A(new_n2623_), .B(new_n620_), .Y(new_n2624_));
  NOR2  g02239(.A(new_n2624_), .B(new_n626_), .Y(new_n2625_));
  NOR2  g02240(.A(new_n2625_), .B(new_n630_), .Y(new_n2626_));
  NOR2  g02241(.A(new_n2626_), .B(new_n636_), .Y(new_n2627_));
  NOR2  g02242(.A(new_n2627_), .B(new_n640_), .Y(new_n2628_));
  NOR2  g02243(.A(new_n2628_), .B(new_n646_), .Y(new_n2629_));
  NOR2  g02244(.A(new_n2629_), .B(new_n650_), .Y(new_n2630_));
  NOR2  g02245(.A(new_n2630_), .B(new_n656_), .Y(new_n2631_));
  NOR2  g02246(.A(new_n2631_), .B(new_n660_), .Y(new_n2632_));
  NOR2  g02247(.A(new_n2632_), .B(new_n666_), .Y(new_n2633_));
  NOR2  g02248(.A(new_n2633_), .B(new_n670_), .Y(new_n2634_));
  NOR2  g02249(.A(new_n2634_), .B(new_n676_), .Y(new_n2635_));
  NOR2  g02250(.A(new_n2635_), .B(new_n680_), .Y(new_n2636_));
  NOR2  g02251(.A(new_n2636_), .B(new_n686_), .Y(new_n2637_));
  NOR2  g02252(.A(new_n2637_), .B(new_n690_), .Y(new_n2638_));
  NOR2  g02253(.A(new_n2638_), .B(new_n696_), .Y(new_n2639_));
  NOR2  g02254(.A(new_n2639_), .B(new_n700_), .Y(new_n2640_));
  NOR2  g02255(.A(new_n2640_), .B(new_n706_), .Y(new_n2641_));
  NOR2  g02256(.A(new_n2641_), .B(new_n710_), .Y(new_n2642_));
  NOR2  g02257(.A(new_n2642_), .B(new_n716_), .Y(new_n2643_));
  NOR2  g02258(.A(new_n2643_), .B(new_n720_), .Y(new_n2644_));
  NOR2  g02259(.A(new_n2644_), .B(new_n726_), .Y(new_n2645_));
  NOR2  g02260(.A(new_n2645_), .B(new_n730_), .Y(new_n2646_));
  NOR2  g02261(.A(new_n2646_), .B(new_n736_), .Y(new_n2647_));
  NOR2  g02262(.A(new_n2647_), .B(new_n740_), .Y(new_n2648_));
  NOR2  g02263(.A(new_n2648_), .B(new_n746_), .Y(new_n2649_));
  NOR2  g02264(.A(new_n2649_), .B(new_n750_), .Y(new_n2650_));
  NOR2  g02265(.A(new_n2650_), .B(new_n756_), .Y(new_n2651_));
  NOR2  g02266(.A(new_n2651_), .B(new_n760_), .Y(new_n2652_));
  NOR2  g02267(.A(new_n2652_), .B(new_n766_), .Y(new_n2653_));
  NOR2  g02268(.A(new_n2653_), .B(new_n770_), .Y(new_n2654_));
  NOR2  g02269(.A(new_n2654_), .B(new_n776_), .Y(new_n2655_));
  NOR2  g02270(.A(new_n2655_), .B(new_n780_), .Y(new_n2656_));
  NOR2  g02271(.A(new_n2656_), .B(new_n786_), .Y(new_n2657_));
  NOR2  g02272(.A(new_n2657_), .B(new_n790_), .Y(new_n2658_));
  NOR2  g02273(.A(new_n2658_), .B(new_n796_), .Y(new_n2659_));
  NOR2  g02274(.A(new_n2659_), .B(new_n800_), .Y(new_n2660_));
  NOR2  g02275(.A(new_n2660_), .B(new_n806_), .Y(new_n2661_));
  NOR2  g02276(.A(new_n2661_), .B(new_n1616_), .Y(new_n2662_));
  NOR2  g02277(.A(new_n2662_), .B(new_n1618_), .Y(new_n2663_));
  NOR2  g02278(.A(new_n2663_), .B(new_n1885_), .Y(new_n2664_));
  NOR2  g02279(.A(new_n2664_), .B(new_n820_), .Y(new_n2665_));
  NOR2  g02280(.A(new_n2665_), .B(new_n824_), .Y(new_n2666_));
  NOR2  g02281(.A(new_n2666_), .B(new_n829_), .Y(new_n2667_));
  NOR2  g02282(.A(new_n2667_), .B(new_n833_), .Y(new_n2668_));
  NOR2  g02283(.A(new_n2668_), .B(new_n838_), .Y(new_n2669_));
  NOR2  g02284(.A(new_n2669_), .B(new_n842_), .Y(new_n2670_));
  NOR2  g02285(.A(new_n2670_), .B(new_n847_), .Y(new_n2671_));
  NAND2 g02286(.A(new_n849_), .B(\req[15] ), .Y(new_n2672_));
  NOR2  g02287(.A(new_n2672_), .B(new_n2671_), .Y(\grant[15] ));
  INV   g02288(.A(new_n859_), .Y(new_n2674_));
  NOR2  g02289(.A(new_n1230_), .B(new_n2674_), .Y(new_n2675_));
  NOR2  g02290(.A(new_n2675_), .B(new_n865_), .Y(new_n2676_));
  NOR2  g02291(.A(new_n2676_), .B(new_n869_), .Y(new_n2677_));
  NOR2  g02292(.A(new_n2677_), .B(new_n874_), .Y(new_n2678_));
  NOR2  g02293(.A(new_n2678_), .B(new_n878_), .Y(new_n2679_));
  NOR2  g02294(.A(new_n2679_), .B(new_n883_), .Y(new_n2680_));
  NOR2  g02295(.A(new_n2680_), .B(new_n887_), .Y(new_n2681_));
  NOR2  g02296(.A(new_n2681_), .B(new_n892_), .Y(new_n2682_));
  NOR2  g02297(.A(new_n2682_), .B(new_n896_), .Y(new_n2683_));
  NOR2  g02298(.A(new_n2683_), .B(new_n901_), .Y(new_n2684_));
  NOR2  g02299(.A(new_n2684_), .B(new_n905_), .Y(new_n2685_));
  NOR2  g02300(.A(new_n2685_), .B(new_n910_), .Y(new_n2686_));
  NOR2  g02301(.A(new_n2686_), .B(new_n914_), .Y(new_n2687_));
  NOR2  g02302(.A(new_n2687_), .B(new_n919_), .Y(new_n2688_));
  NOR2  g02303(.A(new_n2688_), .B(new_n923_), .Y(new_n2689_));
  NOR2  g02304(.A(new_n2689_), .B(new_n928_), .Y(new_n2690_));
  NOR2  g02305(.A(new_n2690_), .B(new_n932_), .Y(new_n2691_));
  NOR2  g02306(.A(new_n2691_), .B(new_n937_), .Y(new_n2692_));
  NOR2  g02307(.A(new_n2692_), .B(new_n941_), .Y(new_n2693_));
  NOR2  g02308(.A(new_n2693_), .B(new_n946_), .Y(new_n2694_));
  NOR2  g02309(.A(new_n2694_), .B(new_n950_), .Y(new_n2695_));
  NOR2  g02310(.A(new_n2695_), .B(new_n955_), .Y(new_n2696_));
  NOR2  g02311(.A(new_n2696_), .B(new_n959_), .Y(new_n2697_));
  NOR2  g02312(.A(new_n2697_), .B(new_n964_), .Y(new_n2698_));
  NOR2  g02313(.A(new_n2698_), .B(new_n968_), .Y(new_n2699_));
  NOR2  g02314(.A(new_n2699_), .B(new_n973_), .Y(new_n2700_));
  NOR2  g02315(.A(new_n2700_), .B(new_n977_), .Y(new_n2701_));
  NOR2  g02316(.A(new_n2701_), .B(new_n982_), .Y(new_n2702_));
  NOR2  g02317(.A(new_n2702_), .B(new_n986_), .Y(new_n2703_));
  NOR2  g02318(.A(new_n2703_), .B(new_n991_), .Y(new_n2704_));
  NOR2  g02319(.A(new_n2704_), .B(new_n995_), .Y(new_n2705_));
  NOR2  g02320(.A(new_n2705_), .B(new_n1000_), .Y(new_n2706_));
  NOR2  g02321(.A(new_n2706_), .B(new_n1004_), .Y(new_n2707_));
  NOR2  g02322(.A(new_n2707_), .B(new_n1009_), .Y(new_n2708_));
  NOR2  g02323(.A(new_n2708_), .B(new_n1013_), .Y(new_n2709_));
  NOR2  g02324(.A(new_n2709_), .B(new_n1018_), .Y(new_n2710_));
  NOR2  g02325(.A(new_n2710_), .B(new_n1022_), .Y(new_n2711_));
  NOR2  g02326(.A(new_n2711_), .B(new_n1027_), .Y(new_n2712_));
  NOR2  g02327(.A(new_n2712_), .B(new_n1031_), .Y(new_n2713_));
  NOR2  g02328(.A(new_n2713_), .B(new_n1036_), .Y(new_n2714_));
  NOR2  g02329(.A(new_n2714_), .B(new_n1040_), .Y(new_n2715_));
  NOR2  g02330(.A(new_n2715_), .B(new_n1045_), .Y(new_n2716_));
  NOR2  g02331(.A(new_n2716_), .B(new_n1049_), .Y(new_n2717_));
  NOR2  g02332(.A(new_n2717_), .B(new_n1054_), .Y(new_n2718_));
  NOR2  g02333(.A(new_n2718_), .B(new_n1058_), .Y(new_n2719_));
  NOR2  g02334(.A(new_n2719_), .B(new_n1063_), .Y(new_n2720_));
  NOR2  g02335(.A(new_n2720_), .B(new_n1067_), .Y(new_n2721_));
  NOR2  g02336(.A(new_n2721_), .B(new_n1072_), .Y(new_n2722_));
  NOR2  g02337(.A(new_n2722_), .B(new_n1076_), .Y(new_n2723_));
  NOR2  g02338(.A(new_n2723_), .B(new_n1081_), .Y(new_n2724_));
  NOR2  g02339(.A(new_n2724_), .B(new_n1085_), .Y(new_n2725_));
  NOR2  g02340(.A(new_n2725_), .B(new_n1090_), .Y(new_n2726_));
  NOR2  g02341(.A(new_n2726_), .B(new_n1094_), .Y(new_n2727_));
  NOR2  g02342(.A(new_n2727_), .B(new_n1099_), .Y(new_n2728_));
  NOR2  g02343(.A(new_n2728_), .B(new_n1103_), .Y(new_n2729_));
  NOR2  g02344(.A(new_n2729_), .B(new_n1108_), .Y(new_n2730_));
  NOR2  g02345(.A(new_n2730_), .B(new_n1112_), .Y(new_n2731_));
  NOR2  g02346(.A(new_n2731_), .B(new_n1117_), .Y(new_n2732_));
  NOR2  g02347(.A(new_n2732_), .B(new_n1121_), .Y(new_n2733_));
  NOR2  g02348(.A(new_n2733_), .B(new_n1126_), .Y(new_n2734_));
  NOR2  g02349(.A(new_n2734_), .B(new_n1130_), .Y(new_n2735_));
  NOR2  g02350(.A(new_n2735_), .B(new_n1135_), .Y(new_n2736_));
  NOR2  g02351(.A(new_n2736_), .B(new_n1139_), .Y(new_n2737_));
  NOR2  g02352(.A(new_n2737_), .B(new_n1144_), .Y(new_n2738_));
  NOR2  g02353(.A(new_n2738_), .B(new_n1148_), .Y(new_n2739_));
  NOR2  g02354(.A(new_n2739_), .B(new_n1153_), .Y(new_n2740_));
  NOR2  g02355(.A(new_n2740_), .B(new_n1157_), .Y(new_n2741_));
  NOR2  g02356(.A(new_n2741_), .B(new_n1162_), .Y(new_n2742_));
  NOR2  g02357(.A(new_n2742_), .B(new_n1166_), .Y(new_n2743_));
  NOR2  g02358(.A(new_n2743_), .B(new_n1171_), .Y(new_n2744_));
  NOR2  g02359(.A(new_n2744_), .B(new_n1175_), .Y(new_n2745_));
  NOR2  g02360(.A(new_n2745_), .B(new_n1180_), .Y(new_n2746_));
  NOR2  g02361(.A(new_n2746_), .B(new_n1184_), .Y(new_n2747_));
  NOR2  g02362(.A(new_n2747_), .B(new_n1189_), .Y(new_n2748_));
  NOR2  g02363(.A(new_n2748_), .B(new_n1707_), .Y(new_n2749_));
  NOR2  g02364(.A(new_n2749_), .B(new_n1709_), .Y(new_n2750_));
  NOR2  g02365(.A(new_n2750_), .B(new_n1973_), .Y(new_n2751_));
  NOR2  g02366(.A(new_n2751_), .B(new_n1199_), .Y(new_n2752_));
  NOR2  g02367(.A(new_n2752_), .B(new_n1203_), .Y(new_n2753_));
  NOR2  g02368(.A(new_n2753_), .B(new_n1207_), .Y(new_n2754_));
  NOR2  g02369(.A(new_n2754_), .B(new_n1211_), .Y(new_n2755_));
  NOR2  g02370(.A(new_n2755_), .B(new_n1215_), .Y(new_n2756_));
  NOR2  g02371(.A(new_n2756_), .B(new_n1219_), .Y(new_n2757_));
  NOR2  g02372(.A(new_n2757_), .B(new_n1223_), .Y(new_n2758_));
  NAND2 g02373(.A(new_n1225_), .B(\req[16] ), .Y(new_n2759_));
  NOR2  g02374(.A(new_n2759_), .B(new_n2758_), .Y(\grant[16] ));
  INV   g02375(.A(new_n1234_), .Y(new_n2761_));
  NOR2  g02376(.A(new_n2761_), .B(new_n445_), .Y(new_n2762_));
  NOR2  g02377(.A(new_n2762_), .B(new_n1239_), .Y(new_n2763_));
  NOR2  g02378(.A(new_n2763_), .B(new_n1243_), .Y(new_n2764_));
  NOR2  g02379(.A(new_n2764_), .B(new_n1247_), .Y(new_n2765_));
  NOR2  g02380(.A(new_n2765_), .B(new_n1251_), .Y(new_n2766_));
  NOR2  g02381(.A(new_n2766_), .B(new_n1255_), .Y(new_n2767_));
  NOR2  g02382(.A(new_n2767_), .B(new_n1259_), .Y(new_n2768_));
  NOR2  g02383(.A(new_n2768_), .B(new_n1263_), .Y(new_n2769_));
  NOR2  g02384(.A(new_n2769_), .B(new_n1267_), .Y(new_n2770_));
  NOR2  g02385(.A(new_n2770_), .B(new_n1271_), .Y(new_n2771_));
  NOR2  g02386(.A(new_n2771_), .B(new_n1275_), .Y(new_n2772_));
  NOR2  g02387(.A(new_n2772_), .B(new_n1279_), .Y(new_n2773_));
  NOR2  g02388(.A(new_n2773_), .B(new_n1283_), .Y(new_n2774_));
  NOR2  g02389(.A(new_n2774_), .B(new_n1287_), .Y(new_n2775_));
  NOR2  g02390(.A(new_n2775_), .B(new_n1291_), .Y(new_n2776_));
  NOR2  g02391(.A(new_n2776_), .B(new_n1295_), .Y(new_n2777_));
  NOR2  g02392(.A(new_n2777_), .B(new_n1299_), .Y(new_n2778_));
  NOR2  g02393(.A(new_n2778_), .B(new_n1303_), .Y(new_n2779_));
  NOR2  g02394(.A(new_n2779_), .B(new_n1307_), .Y(new_n2780_));
  NOR2  g02395(.A(new_n2780_), .B(new_n1311_), .Y(new_n2781_));
  NOR2  g02396(.A(new_n2781_), .B(new_n1315_), .Y(new_n2782_));
  NOR2  g02397(.A(new_n2782_), .B(new_n1319_), .Y(new_n2783_));
  NOR2  g02398(.A(new_n2783_), .B(new_n1323_), .Y(new_n2784_));
  NOR2  g02399(.A(new_n2784_), .B(new_n1327_), .Y(new_n2785_));
  NOR2  g02400(.A(new_n2785_), .B(new_n1331_), .Y(new_n2786_));
  NOR2  g02401(.A(new_n2786_), .B(new_n1335_), .Y(new_n2787_));
  NOR2  g02402(.A(new_n2787_), .B(new_n1339_), .Y(new_n2788_));
  NOR2  g02403(.A(new_n2788_), .B(new_n1343_), .Y(new_n2789_));
  NOR2  g02404(.A(new_n2789_), .B(new_n1347_), .Y(new_n2790_));
  NOR2  g02405(.A(new_n2790_), .B(new_n1351_), .Y(new_n2791_));
  NOR2  g02406(.A(new_n2791_), .B(new_n1355_), .Y(new_n2792_));
  NOR2  g02407(.A(new_n2792_), .B(new_n1359_), .Y(new_n2793_));
  NOR2  g02408(.A(new_n2793_), .B(new_n1363_), .Y(new_n2794_));
  NOR2  g02409(.A(new_n2794_), .B(new_n1367_), .Y(new_n2795_));
  NOR2  g02410(.A(new_n2795_), .B(new_n1371_), .Y(new_n2796_));
  NOR2  g02411(.A(new_n2796_), .B(new_n1375_), .Y(new_n2797_));
  NOR2  g02412(.A(new_n2797_), .B(new_n1379_), .Y(new_n2798_));
  NOR2  g02413(.A(new_n2798_), .B(new_n1383_), .Y(new_n2799_));
  NOR2  g02414(.A(new_n2799_), .B(new_n1387_), .Y(new_n2800_));
  NOR2  g02415(.A(new_n2800_), .B(new_n1391_), .Y(new_n2801_));
  NOR2  g02416(.A(new_n2801_), .B(new_n1395_), .Y(new_n2802_));
  NOR2  g02417(.A(new_n2802_), .B(new_n1399_), .Y(new_n2803_));
  NOR2  g02418(.A(new_n2803_), .B(new_n1403_), .Y(new_n2804_));
  NOR2  g02419(.A(new_n2804_), .B(new_n1407_), .Y(new_n2805_));
  NOR2  g02420(.A(new_n2805_), .B(new_n1411_), .Y(new_n2806_));
  NOR2  g02421(.A(new_n2806_), .B(new_n1415_), .Y(new_n2807_));
  NOR2  g02422(.A(new_n2807_), .B(new_n1419_), .Y(new_n2808_));
  NOR2  g02423(.A(new_n2808_), .B(new_n1423_), .Y(new_n2809_));
  NOR2  g02424(.A(new_n2809_), .B(new_n1427_), .Y(new_n2810_));
  NOR2  g02425(.A(new_n2810_), .B(new_n1431_), .Y(new_n2811_));
  NOR2  g02426(.A(new_n2811_), .B(new_n1435_), .Y(new_n2812_));
  NOR2  g02427(.A(new_n2812_), .B(new_n1439_), .Y(new_n2813_));
  NOR2  g02428(.A(new_n2813_), .B(new_n1443_), .Y(new_n2814_));
  NOR2  g02429(.A(new_n2814_), .B(new_n1447_), .Y(new_n2815_));
  NOR2  g02430(.A(new_n2815_), .B(new_n1451_), .Y(new_n2816_));
  NOR2  g02431(.A(new_n2816_), .B(new_n1455_), .Y(new_n2817_));
  NOR2  g02432(.A(new_n2817_), .B(new_n1459_), .Y(new_n2818_));
  NOR2  g02433(.A(new_n2818_), .B(new_n1463_), .Y(new_n2819_));
  NOR2  g02434(.A(new_n2819_), .B(new_n1467_), .Y(new_n2820_));
  NOR2  g02435(.A(new_n2820_), .B(new_n1471_), .Y(new_n2821_));
  NOR2  g02436(.A(new_n2821_), .B(new_n1475_), .Y(new_n2822_));
  NOR2  g02437(.A(new_n2822_), .B(new_n1479_), .Y(new_n2823_));
  NOR2  g02438(.A(new_n2823_), .B(new_n1483_), .Y(new_n2824_));
  NOR2  g02439(.A(new_n2824_), .B(new_n1487_), .Y(new_n2825_));
  NOR2  g02440(.A(new_n2825_), .B(new_n1491_), .Y(new_n2826_));
  NOR2  g02441(.A(new_n2826_), .B(new_n1495_), .Y(new_n2827_));
  NOR2  g02442(.A(new_n2827_), .B(new_n1499_), .Y(new_n2828_));
  NOR2  g02443(.A(new_n2828_), .B(new_n1503_), .Y(new_n2829_));
  NOR2  g02444(.A(new_n2829_), .B(new_n1507_), .Y(new_n2830_));
  NOR2  g02445(.A(new_n2830_), .B(new_n1511_), .Y(new_n2831_));
  NOR2  g02446(.A(new_n2831_), .B(new_n1515_), .Y(new_n2832_));
  NOR2  g02447(.A(new_n2832_), .B(new_n1519_), .Y(new_n2833_));
  NOR2  g02448(.A(new_n2833_), .B(new_n1523_), .Y(new_n2834_));
  NOR2  g02449(.A(new_n2834_), .B(new_n1527_), .Y(new_n2835_));
  NOR2  g02450(.A(new_n2835_), .B(new_n1797_), .Y(new_n2836_));
  NOR2  g02451(.A(new_n2836_), .B(new_n396_), .Y(new_n2837_));
  NOR2  g02452(.A(new_n2837_), .B(new_n400_), .Y(new_n2838_));
  NOR2  g02453(.A(new_n2838_), .B(new_n406_), .Y(new_n2839_));
  NOR2  g02454(.A(new_n2839_), .B(new_n410_), .Y(new_n2840_));
  NOR2  g02455(.A(new_n2840_), .B(new_n416_), .Y(new_n2841_));
  NOR2  g02456(.A(new_n2841_), .B(new_n420_), .Y(new_n2842_));
  NOR2  g02457(.A(new_n2842_), .B(new_n426_), .Y(new_n2843_));
  NOR2  g02458(.A(new_n2843_), .B(new_n430_), .Y(new_n2844_));
  NOR2  g02459(.A(new_n2844_), .B(new_n436_), .Y(new_n2845_));
  NAND2 g02460(.A(new_n438_), .B(\req[17] ), .Y(new_n2846_));
  NOR2  g02461(.A(new_n2846_), .B(new_n2845_), .Y(\grant[17] ));
  INV   g02462(.A(new_n449_), .Y(new_n2848_));
  NOR2  g02463(.A(new_n864_), .B(new_n2848_), .Y(new_n2849_));
  NOR2  g02464(.A(new_n2849_), .B(new_n456_), .Y(new_n2850_));
  NOR2  g02465(.A(new_n2850_), .B(new_n460_), .Y(new_n2851_));
  NOR2  g02466(.A(new_n2851_), .B(new_n466_), .Y(new_n2852_));
  NOR2  g02467(.A(new_n2852_), .B(new_n470_), .Y(new_n2853_));
  NOR2  g02468(.A(new_n2853_), .B(new_n476_), .Y(new_n2854_));
  NOR2  g02469(.A(new_n2854_), .B(new_n480_), .Y(new_n2855_));
  NOR2  g02470(.A(new_n2855_), .B(new_n486_), .Y(new_n2856_));
  NOR2  g02471(.A(new_n2856_), .B(new_n490_), .Y(new_n2857_));
  NOR2  g02472(.A(new_n2857_), .B(new_n496_), .Y(new_n2858_));
  NOR2  g02473(.A(new_n2858_), .B(new_n500_), .Y(new_n2859_));
  NOR2  g02474(.A(new_n2859_), .B(new_n506_), .Y(new_n2860_));
  NOR2  g02475(.A(new_n2860_), .B(new_n510_), .Y(new_n2861_));
  NOR2  g02476(.A(new_n2861_), .B(new_n516_), .Y(new_n2862_));
  NOR2  g02477(.A(new_n2862_), .B(new_n520_), .Y(new_n2863_));
  NOR2  g02478(.A(new_n2863_), .B(new_n526_), .Y(new_n2864_));
  NOR2  g02479(.A(new_n2864_), .B(new_n530_), .Y(new_n2865_));
  NOR2  g02480(.A(new_n2865_), .B(new_n536_), .Y(new_n2866_));
  NOR2  g02481(.A(new_n2866_), .B(new_n540_), .Y(new_n2867_));
  NOR2  g02482(.A(new_n2867_), .B(new_n546_), .Y(new_n2868_));
  NOR2  g02483(.A(new_n2868_), .B(new_n550_), .Y(new_n2869_));
  NOR2  g02484(.A(new_n2869_), .B(new_n556_), .Y(new_n2870_));
  NOR2  g02485(.A(new_n2870_), .B(new_n560_), .Y(new_n2871_));
  NOR2  g02486(.A(new_n2871_), .B(new_n566_), .Y(new_n2872_));
  NOR2  g02487(.A(new_n2872_), .B(new_n570_), .Y(new_n2873_));
  NOR2  g02488(.A(new_n2873_), .B(new_n576_), .Y(new_n2874_));
  NOR2  g02489(.A(new_n2874_), .B(new_n580_), .Y(new_n2875_));
  NOR2  g02490(.A(new_n2875_), .B(new_n586_), .Y(new_n2876_));
  NOR2  g02491(.A(new_n2876_), .B(new_n590_), .Y(new_n2877_));
  NOR2  g02492(.A(new_n2877_), .B(new_n596_), .Y(new_n2878_));
  NOR2  g02493(.A(new_n2878_), .B(new_n600_), .Y(new_n2879_));
  NOR2  g02494(.A(new_n2879_), .B(new_n606_), .Y(new_n2880_));
  NOR2  g02495(.A(new_n2880_), .B(new_n610_), .Y(new_n2881_));
  NOR2  g02496(.A(new_n2881_), .B(new_n616_), .Y(new_n2882_));
  NOR2  g02497(.A(new_n2882_), .B(new_n620_), .Y(new_n2883_));
  NOR2  g02498(.A(new_n2883_), .B(new_n626_), .Y(new_n2884_));
  NOR2  g02499(.A(new_n2884_), .B(new_n630_), .Y(new_n2885_));
  NOR2  g02500(.A(new_n2885_), .B(new_n636_), .Y(new_n2886_));
  NOR2  g02501(.A(new_n2886_), .B(new_n640_), .Y(new_n2887_));
  NOR2  g02502(.A(new_n2887_), .B(new_n646_), .Y(new_n2888_));
  NOR2  g02503(.A(new_n2888_), .B(new_n650_), .Y(new_n2889_));
  NOR2  g02504(.A(new_n2889_), .B(new_n656_), .Y(new_n2890_));
  NOR2  g02505(.A(new_n2890_), .B(new_n660_), .Y(new_n2891_));
  NOR2  g02506(.A(new_n2891_), .B(new_n666_), .Y(new_n2892_));
  NOR2  g02507(.A(new_n2892_), .B(new_n670_), .Y(new_n2893_));
  NOR2  g02508(.A(new_n2893_), .B(new_n676_), .Y(new_n2894_));
  NOR2  g02509(.A(new_n2894_), .B(new_n680_), .Y(new_n2895_));
  NOR2  g02510(.A(new_n2895_), .B(new_n686_), .Y(new_n2896_));
  NOR2  g02511(.A(new_n2896_), .B(new_n690_), .Y(new_n2897_));
  NOR2  g02512(.A(new_n2897_), .B(new_n696_), .Y(new_n2898_));
  NOR2  g02513(.A(new_n2898_), .B(new_n700_), .Y(new_n2899_));
  NOR2  g02514(.A(new_n2899_), .B(new_n706_), .Y(new_n2900_));
  NOR2  g02515(.A(new_n2900_), .B(new_n710_), .Y(new_n2901_));
  NOR2  g02516(.A(new_n2901_), .B(new_n716_), .Y(new_n2902_));
  NOR2  g02517(.A(new_n2902_), .B(new_n720_), .Y(new_n2903_));
  NOR2  g02518(.A(new_n2903_), .B(new_n726_), .Y(new_n2904_));
  NOR2  g02519(.A(new_n2904_), .B(new_n730_), .Y(new_n2905_));
  NOR2  g02520(.A(new_n2905_), .B(new_n736_), .Y(new_n2906_));
  NOR2  g02521(.A(new_n2906_), .B(new_n740_), .Y(new_n2907_));
  NOR2  g02522(.A(new_n2907_), .B(new_n746_), .Y(new_n2908_));
  NOR2  g02523(.A(new_n2908_), .B(new_n750_), .Y(new_n2909_));
  NOR2  g02524(.A(new_n2909_), .B(new_n756_), .Y(new_n2910_));
  NOR2  g02525(.A(new_n2910_), .B(new_n760_), .Y(new_n2911_));
  NOR2  g02526(.A(new_n2911_), .B(new_n766_), .Y(new_n2912_));
  NOR2  g02527(.A(new_n2912_), .B(new_n770_), .Y(new_n2913_));
  NOR2  g02528(.A(new_n2913_), .B(new_n776_), .Y(new_n2914_));
  NOR2  g02529(.A(new_n2914_), .B(new_n780_), .Y(new_n2915_));
  NOR2  g02530(.A(new_n2915_), .B(new_n786_), .Y(new_n2916_));
  NOR2  g02531(.A(new_n2916_), .B(new_n790_), .Y(new_n2917_));
  NOR2  g02532(.A(new_n2917_), .B(new_n796_), .Y(new_n2918_));
  NOR2  g02533(.A(new_n2918_), .B(new_n800_), .Y(new_n2919_));
  NOR2  g02534(.A(new_n2919_), .B(new_n806_), .Y(new_n2920_));
  NOR2  g02535(.A(new_n2920_), .B(new_n1616_), .Y(new_n2921_));
  NOR2  g02536(.A(new_n2921_), .B(new_n1618_), .Y(new_n2922_));
  NOR2  g02537(.A(new_n2922_), .B(new_n1885_), .Y(new_n2923_));
  NOR2  g02538(.A(new_n2923_), .B(new_n820_), .Y(new_n2924_));
  NOR2  g02539(.A(new_n2924_), .B(new_n824_), .Y(new_n2925_));
  NOR2  g02540(.A(new_n2925_), .B(new_n829_), .Y(new_n2926_));
  NOR2  g02541(.A(new_n2926_), .B(new_n833_), .Y(new_n2927_));
  NOR2  g02542(.A(new_n2927_), .B(new_n838_), .Y(new_n2928_));
  NOR2  g02543(.A(new_n2928_), .B(new_n842_), .Y(new_n2929_));
  NOR2  g02544(.A(new_n2929_), .B(new_n847_), .Y(new_n2930_));
  NOR2  g02545(.A(new_n2930_), .B(new_n851_), .Y(new_n2931_));
  NOR2  g02546(.A(new_n2931_), .B(new_n856_), .Y(new_n2932_));
  NAND2 g02547(.A(new_n858_), .B(\req[18] ), .Y(new_n2933_));
  NOR2  g02548(.A(new_n2933_), .B(new_n2932_), .Y(\grant[18] ));
  INV   g02549(.A(new_n868_), .Y(new_n2935_));
  NOR2  g02550(.A(new_n1238_), .B(new_n2935_), .Y(new_n2936_));
  NOR2  g02551(.A(new_n2936_), .B(new_n874_), .Y(new_n2937_));
  NOR2  g02552(.A(new_n2937_), .B(new_n878_), .Y(new_n2938_));
  NOR2  g02553(.A(new_n2938_), .B(new_n883_), .Y(new_n2939_));
  NOR2  g02554(.A(new_n2939_), .B(new_n887_), .Y(new_n2940_));
  NOR2  g02555(.A(new_n2940_), .B(new_n892_), .Y(new_n2941_));
  NOR2  g02556(.A(new_n2941_), .B(new_n896_), .Y(new_n2942_));
  NOR2  g02557(.A(new_n2942_), .B(new_n901_), .Y(new_n2943_));
  NOR2  g02558(.A(new_n2943_), .B(new_n905_), .Y(new_n2944_));
  NOR2  g02559(.A(new_n2944_), .B(new_n910_), .Y(new_n2945_));
  NOR2  g02560(.A(new_n2945_), .B(new_n914_), .Y(new_n2946_));
  NOR2  g02561(.A(new_n2946_), .B(new_n919_), .Y(new_n2947_));
  NOR2  g02562(.A(new_n2947_), .B(new_n923_), .Y(new_n2948_));
  NOR2  g02563(.A(new_n2948_), .B(new_n928_), .Y(new_n2949_));
  NOR2  g02564(.A(new_n2949_), .B(new_n932_), .Y(new_n2950_));
  NOR2  g02565(.A(new_n2950_), .B(new_n937_), .Y(new_n2951_));
  NOR2  g02566(.A(new_n2951_), .B(new_n941_), .Y(new_n2952_));
  NOR2  g02567(.A(new_n2952_), .B(new_n946_), .Y(new_n2953_));
  NOR2  g02568(.A(new_n2953_), .B(new_n950_), .Y(new_n2954_));
  NOR2  g02569(.A(new_n2954_), .B(new_n955_), .Y(new_n2955_));
  NOR2  g02570(.A(new_n2955_), .B(new_n959_), .Y(new_n2956_));
  NOR2  g02571(.A(new_n2956_), .B(new_n964_), .Y(new_n2957_));
  NOR2  g02572(.A(new_n2957_), .B(new_n968_), .Y(new_n2958_));
  NOR2  g02573(.A(new_n2958_), .B(new_n973_), .Y(new_n2959_));
  NOR2  g02574(.A(new_n2959_), .B(new_n977_), .Y(new_n2960_));
  NOR2  g02575(.A(new_n2960_), .B(new_n982_), .Y(new_n2961_));
  NOR2  g02576(.A(new_n2961_), .B(new_n986_), .Y(new_n2962_));
  NOR2  g02577(.A(new_n2962_), .B(new_n991_), .Y(new_n2963_));
  NOR2  g02578(.A(new_n2963_), .B(new_n995_), .Y(new_n2964_));
  NOR2  g02579(.A(new_n2964_), .B(new_n1000_), .Y(new_n2965_));
  NOR2  g02580(.A(new_n2965_), .B(new_n1004_), .Y(new_n2966_));
  NOR2  g02581(.A(new_n2966_), .B(new_n1009_), .Y(new_n2967_));
  NOR2  g02582(.A(new_n2967_), .B(new_n1013_), .Y(new_n2968_));
  NOR2  g02583(.A(new_n2968_), .B(new_n1018_), .Y(new_n2969_));
  NOR2  g02584(.A(new_n2969_), .B(new_n1022_), .Y(new_n2970_));
  NOR2  g02585(.A(new_n2970_), .B(new_n1027_), .Y(new_n2971_));
  NOR2  g02586(.A(new_n2971_), .B(new_n1031_), .Y(new_n2972_));
  NOR2  g02587(.A(new_n2972_), .B(new_n1036_), .Y(new_n2973_));
  NOR2  g02588(.A(new_n2973_), .B(new_n1040_), .Y(new_n2974_));
  NOR2  g02589(.A(new_n2974_), .B(new_n1045_), .Y(new_n2975_));
  NOR2  g02590(.A(new_n2975_), .B(new_n1049_), .Y(new_n2976_));
  NOR2  g02591(.A(new_n2976_), .B(new_n1054_), .Y(new_n2977_));
  NOR2  g02592(.A(new_n2977_), .B(new_n1058_), .Y(new_n2978_));
  NOR2  g02593(.A(new_n2978_), .B(new_n1063_), .Y(new_n2979_));
  NOR2  g02594(.A(new_n2979_), .B(new_n1067_), .Y(new_n2980_));
  NOR2  g02595(.A(new_n2980_), .B(new_n1072_), .Y(new_n2981_));
  NOR2  g02596(.A(new_n2981_), .B(new_n1076_), .Y(new_n2982_));
  NOR2  g02597(.A(new_n2982_), .B(new_n1081_), .Y(new_n2983_));
  NOR2  g02598(.A(new_n2983_), .B(new_n1085_), .Y(new_n2984_));
  NOR2  g02599(.A(new_n2984_), .B(new_n1090_), .Y(new_n2985_));
  NOR2  g02600(.A(new_n2985_), .B(new_n1094_), .Y(new_n2986_));
  NOR2  g02601(.A(new_n2986_), .B(new_n1099_), .Y(new_n2987_));
  NOR2  g02602(.A(new_n2987_), .B(new_n1103_), .Y(new_n2988_));
  NOR2  g02603(.A(new_n2988_), .B(new_n1108_), .Y(new_n2989_));
  NOR2  g02604(.A(new_n2989_), .B(new_n1112_), .Y(new_n2990_));
  NOR2  g02605(.A(new_n2990_), .B(new_n1117_), .Y(new_n2991_));
  NOR2  g02606(.A(new_n2991_), .B(new_n1121_), .Y(new_n2992_));
  NOR2  g02607(.A(new_n2992_), .B(new_n1126_), .Y(new_n2993_));
  NOR2  g02608(.A(new_n2993_), .B(new_n1130_), .Y(new_n2994_));
  NOR2  g02609(.A(new_n2994_), .B(new_n1135_), .Y(new_n2995_));
  NOR2  g02610(.A(new_n2995_), .B(new_n1139_), .Y(new_n2996_));
  NOR2  g02611(.A(new_n2996_), .B(new_n1144_), .Y(new_n2997_));
  NOR2  g02612(.A(new_n2997_), .B(new_n1148_), .Y(new_n2998_));
  NOR2  g02613(.A(new_n2998_), .B(new_n1153_), .Y(new_n2999_));
  NOR2  g02614(.A(new_n2999_), .B(new_n1157_), .Y(new_n3000_));
  NOR2  g02615(.A(new_n3000_), .B(new_n1162_), .Y(new_n3001_));
  NOR2  g02616(.A(new_n3001_), .B(new_n1166_), .Y(new_n3002_));
  NOR2  g02617(.A(new_n3002_), .B(new_n1171_), .Y(new_n3003_));
  NOR2  g02618(.A(new_n3003_), .B(new_n1175_), .Y(new_n3004_));
  NOR2  g02619(.A(new_n3004_), .B(new_n1180_), .Y(new_n3005_));
  NOR2  g02620(.A(new_n3005_), .B(new_n1184_), .Y(new_n3006_));
  NOR2  g02621(.A(new_n3006_), .B(new_n1189_), .Y(new_n3007_));
  NOR2  g02622(.A(new_n3007_), .B(new_n1707_), .Y(new_n3008_));
  NOR2  g02623(.A(new_n3008_), .B(new_n1709_), .Y(new_n3009_));
  NOR2  g02624(.A(new_n3009_), .B(new_n1973_), .Y(new_n3010_));
  NOR2  g02625(.A(new_n3010_), .B(new_n1199_), .Y(new_n3011_));
  NOR2  g02626(.A(new_n3011_), .B(new_n1203_), .Y(new_n3012_));
  NOR2  g02627(.A(new_n3012_), .B(new_n1207_), .Y(new_n3013_));
  NOR2  g02628(.A(new_n3013_), .B(new_n1211_), .Y(new_n3014_));
  NOR2  g02629(.A(new_n3014_), .B(new_n1215_), .Y(new_n3015_));
  NOR2  g02630(.A(new_n3015_), .B(new_n1219_), .Y(new_n3016_));
  NOR2  g02631(.A(new_n3016_), .B(new_n1223_), .Y(new_n3017_));
  NOR2  g02632(.A(new_n3017_), .B(new_n1227_), .Y(new_n3018_));
  NOR2  g02633(.A(new_n3018_), .B(new_n1231_), .Y(new_n3019_));
  NAND2 g02634(.A(new_n1233_), .B(\req[19] ), .Y(new_n3020_));
  NOR2  g02635(.A(new_n3020_), .B(new_n3019_), .Y(\grant[19] ));
  INV   g02636(.A(new_n1242_), .Y(new_n3022_));
  NOR2  g02637(.A(new_n3022_), .B(new_n455_), .Y(new_n3023_));
  NOR2  g02638(.A(new_n3023_), .B(new_n1247_), .Y(new_n3024_));
  NOR2  g02639(.A(new_n3024_), .B(new_n1251_), .Y(new_n3025_));
  NOR2  g02640(.A(new_n3025_), .B(new_n1255_), .Y(new_n3026_));
  NOR2  g02641(.A(new_n3026_), .B(new_n1259_), .Y(new_n3027_));
  NOR2  g02642(.A(new_n3027_), .B(new_n1263_), .Y(new_n3028_));
  NOR2  g02643(.A(new_n3028_), .B(new_n1267_), .Y(new_n3029_));
  NOR2  g02644(.A(new_n3029_), .B(new_n1271_), .Y(new_n3030_));
  NOR2  g02645(.A(new_n3030_), .B(new_n1275_), .Y(new_n3031_));
  NOR2  g02646(.A(new_n3031_), .B(new_n1279_), .Y(new_n3032_));
  NOR2  g02647(.A(new_n3032_), .B(new_n1283_), .Y(new_n3033_));
  NOR2  g02648(.A(new_n3033_), .B(new_n1287_), .Y(new_n3034_));
  NOR2  g02649(.A(new_n3034_), .B(new_n1291_), .Y(new_n3035_));
  NOR2  g02650(.A(new_n3035_), .B(new_n1295_), .Y(new_n3036_));
  NOR2  g02651(.A(new_n3036_), .B(new_n1299_), .Y(new_n3037_));
  NOR2  g02652(.A(new_n3037_), .B(new_n1303_), .Y(new_n3038_));
  NOR2  g02653(.A(new_n3038_), .B(new_n1307_), .Y(new_n3039_));
  NOR2  g02654(.A(new_n3039_), .B(new_n1311_), .Y(new_n3040_));
  NOR2  g02655(.A(new_n3040_), .B(new_n1315_), .Y(new_n3041_));
  NOR2  g02656(.A(new_n3041_), .B(new_n1319_), .Y(new_n3042_));
  NOR2  g02657(.A(new_n3042_), .B(new_n1323_), .Y(new_n3043_));
  NOR2  g02658(.A(new_n3043_), .B(new_n1327_), .Y(new_n3044_));
  NOR2  g02659(.A(new_n3044_), .B(new_n1331_), .Y(new_n3045_));
  NOR2  g02660(.A(new_n3045_), .B(new_n1335_), .Y(new_n3046_));
  NOR2  g02661(.A(new_n3046_), .B(new_n1339_), .Y(new_n3047_));
  NOR2  g02662(.A(new_n3047_), .B(new_n1343_), .Y(new_n3048_));
  NOR2  g02663(.A(new_n3048_), .B(new_n1347_), .Y(new_n3049_));
  NOR2  g02664(.A(new_n3049_), .B(new_n1351_), .Y(new_n3050_));
  NOR2  g02665(.A(new_n3050_), .B(new_n1355_), .Y(new_n3051_));
  NOR2  g02666(.A(new_n3051_), .B(new_n1359_), .Y(new_n3052_));
  NOR2  g02667(.A(new_n3052_), .B(new_n1363_), .Y(new_n3053_));
  NOR2  g02668(.A(new_n3053_), .B(new_n1367_), .Y(new_n3054_));
  NOR2  g02669(.A(new_n3054_), .B(new_n1371_), .Y(new_n3055_));
  NOR2  g02670(.A(new_n3055_), .B(new_n1375_), .Y(new_n3056_));
  NOR2  g02671(.A(new_n3056_), .B(new_n1379_), .Y(new_n3057_));
  NOR2  g02672(.A(new_n3057_), .B(new_n1383_), .Y(new_n3058_));
  NOR2  g02673(.A(new_n3058_), .B(new_n1387_), .Y(new_n3059_));
  NOR2  g02674(.A(new_n3059_), .B(new_n1391_), .Y(new_n3060_));
  NOR2  g02675(.A(new_n3060_), .B(new_n1395_), .Y(new_n3061_));
  NOR2  g02676(.A(new_n3061_), .B(new_n1399_), .Y(new_n3062_));
  NOR2  g02677(.A(new_n3062_), .B(new_n1403_), .Y(new_n3063_));
  NOR2  g02678(.A(new_n3063_), .B(new_n1407_), .Y(new_n3064_));
  NOR2  g02679(.A(new_n3064_), .B(new_n1411_), .Y(new_n3065_));
  NOR2  g02680(.A(new_n3065_), .B(new_n1415_), .Y(new_n3066_));
  NOR2  g02681(.A(new_n3066_), .B(new_n1419_), .Y(new_n3067_));
  NOR2  g02682(.A(new_n3067_), .B(new_n1423_), .Y(new_n3068_));
  NOR2  g02683(.A(new_n3068_), .B(new_n1427_), .Y(new_n3069_));
  NOR2  g02684(.A(new_n3069_), .B(new_n1431_), .Y(new_n3070_));
  NOR2  g02685(.A(new_n3070_), .B(new_n1435_), .Y(new_n3071_));
  NOR2  g02686(.A(new_n3071_), .B(new_n1439_), .Y(new_n3072_));
  NOR2  g02687(.A(new_n3072_), .B(new_n1443_), .Y(new_n3073_));
  NOR2  g02688(.A(new_n3073_), .B(new_n1447_), .Y(new_n3074_));
  NOR2  g02689(.A(new_n3074_), .B(new_n1451_), .Y(new_n3075_));
  NOR2  g02690(.A(new_n3075_), .B(new_n1455_), .Y(new_n3076_));
  NOR2  g02691(.A(new_n3076_), .B(new_n1459_), .Y(new_n3077_));
  NOR2  g02692(.A(new_n3077_), .B(new_n1463_), .Y(new_n3078_));
  NOR2  g02693(.A(new_n3078_), .B(new_n1467_), .Y(new_n3079_));
  NOR2  g02694(.A(new_n3079_), .B(new_n1471_), .Y(new_n3080_));
  NOR2  g02695(.A(new_n3080_), .B(new_n1475_), .Y(new_n3081_));
  NOR2  g02696(.A(new_n3081_), .B(new_n1479_), .Y(new_n3082_));
  NOR2  g02697(.A(new_n3082_), .B(new_n1483_), .Y(new_n3083_));
  NOR2  g02698(.A(new_n3083_), .B(new_n1487_), .Y(new_n3084_));
  NOR2  g02699(.A(new_n3084_), .B(new_n1491_), .Y(new_n3085_));
  NOR2  g02700(.A(new_n3085_), .B(new_n1495_), .Y(new_n3086_));
  NOR2  g02701(.A(new_n3086_), .B(new_n1499_), .Y(new_n3087_));
  NOR2  g02702(.A(new_n3087_), .B(new_n1503_), .Y(new_n3088_));
  NOR2  g02703(.A(new_n3088_), .B(new_n1507_), .Y(new_n3089_));
  NOR2  g02704(.A(new_n3089_), .B(new_n1511_), .Y(new_n3090_));
  NOR2  g02705(.A(new_n3090_), .B(new_n1515_), .Y(new_n3091_));
  NOR2  g02706(.A(new_n3091_), .B(new_n1519_), .Y(new_n3092_));
  NOR2  g02707(.A(new_n3092_), .B(new_n1523_), .Y(new_n3093_));
  NOR2  g02708(.A(new_n3093_), .B(new_n1527_), .Y(new_n3094_));
  NOR2  g02709(.A(new_n3094_), .B(new_n1797_), .Y(new_n3095_));
  NOR2  g02710(.A(new_n3095_), .B(new_n396_), .Y(new_n3096_));
  NOR2  g02711(.A(new_n3096_), .B(new_n400_), .Y(new_n3097_));
  NOR2  g02712(.A(new_n3097_), .B(new_n406_), .Y(new_n3098_));
  NOR2  g02713(.A(new_n3098_), .B(new_n410_), .Y(new_n3099_));
  NOR2  g02714(.A(new_n3099_), .B(new_n416_), .Y(new_n3100_));
  NOR2  g02715(.A(new_n3100_), .B(new_n420_), .Y(new_n3101_));
  NOR2  g02716(.A(new_n3101_), .B(new_n426_), .Y(new_n3102_));
  NOR2  g02717(.A(new_n3102_), .B(new_n430_), .Y(new_n3103_));
  NOR2  g02718(.A(new_n3103_), .B(new_n436_), .Y(new_n3104_));
  NOR2  g02719(.A(new_n3104_), .B(new_n440_), .Y(new_n3105_));
  NOR2  g02720(.A(new_n3105_), .B(new_n446_), .Y(new_n3106_));
  NAND2 g02721(.A(new_n448_), .B(\req[20] ), .Y(new_n3107_));
  NOR2  g02722(.A(new_n3107_), .B(new_n3106_), .Y(\grant[20] ));
  INV   g02723(.A(new_n459_), .Y(new_n3109_));
  NOR2  g02724(.A(new_n873_), .B(new_n3109_), .Y(new_n3110_));
  NOR2  g02725(.A(new_n3110_), .B(new_n466_), .Y(new_n3111_));
  NOR2  g02726(.A(new_n3111_), .B(new_n470_), .Y(new_n3112_));
  NOR2  g02727(.A(new_n3112_), .B(new_n476_), .Y(new_n3113_));
  NOR2  g02728(.A(new_n3113_), .B(new_n480_), .Y(new_n3114_));
  NOR2  g02729(.A(new_n3114_), .B(new_n486_), .Y(new_n3115_));
  NOR2  g02730(.A(new_n3115_), .B(new_n490_), .Y(new_n3116_));
  NOR2  g02731(.A(new_n3116_), .B(new_n496_), .Y(new_n3117_));
  NOR2  g02732(.A(new_n3117_), .B(new_n500_), .Y(new_n3118_));
  NOR2  g02733(.A(new_n3118_), .B(new_n506_), .Y(new_n3119_));
  NOR2  g02734(.A(new_n3119_), .B(new_n510_), .Y(new_n3120_));
  NOR2  g02735(.A(new_n3120_), .B(new_n516_), .Y(new_n3121_));
  NOR2  g02736(.A(new_n3121_), .B(new_n520_), .Y(new_n3122_));
  NOR2  g02737(.A(new_n3122_), .B(new_n526_), .Y(new_n3123_));
  NOR2  g02738(.A(new_n3123_), .B(new_n530_), .Y(new_n3124_));
  NOR2  g02739(.A(new_n3124_), .B(new_n536_), .Y(new_n3125_));
  NOR2  g02740(.A(new_n3125_), .B(new_n540_), .Y(new_n3126_));
  NOR2  g02741(.A(new_n3126_), .B(new_n546_), .Y(new_n3127_));
  NOR2  g02742(.A(new_n3127_), .B(new_n550_), .Y(new_n3128_));
  NOR2  g02743(.A(new_n3128_), .B(new_n556_), .Y(new_n3129_));
  NOR2  g02744(.A(new_n3129_), .B(new_n560_), .Y(new_n3130_));
  NOR2  g02745(.A(new_n3130_), .B(new_n566_), .Y(new_n3131_));
  NOR2  g02746(.A(new_n3131_), .B(new_n570_), .Y(new_n3132_));
  NOR2  g02747(.A(new_n3132_), .B(new_n576_), .Y(new_n3133_));
  NOR2  g02748(.A(new_n3133_), .B(new_n580_), .Y(new_n3134_));
  NOR2  g02749(.A(new_n3134_), .B(new_n586_), .Y(new_n3135_));
  NOR2  g02750(.A(new_n3135_), .B(new_n590_), .Y(new_n3136_));
  NOR2  g02751(.A(new_n3136_), .B(new_n596_), .Y(new_n3137_));
  NOR2  g02752(.A(new_n3137_), .B(new_n600_), .Y(new_n3138_));
  NOR2  g02753(.A(new_n3138_), .B(new_n606_), .Y(new_n3139_));
  NOR2  g02754(.A(new_n3139_), .B(new_n610_), .Y(new_n3140_));
  NOR2  g02755(.A(new_n3140_), .B(new_n616_), .Y(new_n3141_));
  NOR2  g02756(.A(new_n3141_), .B(new_n620_), .Y(new_n3142_));
  NOR2  g02757(.A(new_n3142_), .B(new_n626_), .Y(new_n3143_));
  NOR2  g02758(.A(new_n3143_), .B(new_n630_), .Y(new_n3144_));
  NOR2  g02759(.A(new_n3144_), .B(new_n636_), .Y(new_n3145_));
  NOR2  g02760(.A(new_n3145_), .B(new_n640_), .Y(new_n3146_));
  NOR2  g02761(.A(new_n3146_), .B(new_n646_), .Y(new_n3147_));
  NOR2  g02762(.A(new_n3147_), .B(new_n650_), .Y(new_n3148_));
  NOR2  g02763(.A(new_n3148_), .B(new_n656_), .Y(new_n3149_));
  NOR2  g02764(.A(new_n3149_), .B(new_n660_), .Y(new_n3150_));
  NOR2  g02765(.A(new_n3150_), .B(new_n666_), .Y(new_n3151_));
  NOR2  g02766(.A(new_n3151_), .B(new_n670_), .Y(new_n3152_));
  NOR2  g02767(.A(new_n3152_), .B(new_n676_), .Y(new_n3153_));
  NOR2  g02768(.A(new_n3153_), .B(new_n680_), .Y(new_n3154_));
  NOR2  g02769(.A(new_n3154_), .B(new_n686_), .Y(new_n3155_));
  NOR2  g02770(.A(new_n3155_), .B(new_n690_), .Y(new_n3156_));
  NOR2  g02771(.A(new_n3156_), .B(new_n696_), .Y(new_n3157_));
  NOR2  g02772(.A(new_n3157_), .B(new_n700_), .Y(new_n3158_));
  NOR2  g02773(.A(new_n3158_), .B(new_n706_), .Y(new_n3159_));
  NOR2  g02774(.A(new_n3159_), .B(new_n710_), .Y(new_n3160_));
  NOR2  g02775(.A(new_n3160_), .B(new_n716_), .Y(new_n3161_));
  NOR2  g02776(.A(new_n3161_), .B(new_n720_), .Y(new_n3162_));
  NOR2  g02777(.A(new_n3162_), .B(new_n726_), .Y(new_n3163_));
  NOR2  g02778(.A(new_n3163_), .B(new_n730_), .Y(new_n3164_));
  NOR2  g02779(.A(new_n3164_), .B(new_n736_), .Y(new_n3165_));
  NOR2  g02780(.A(new_n3165_), .B(new_n740_), .Y(new_n3166_));
  NOR2  g02781(.A(new_n3166_), .B(new_n746_), .Y(new_n3167_));
  NOR2  g02782(.A(new_n3167_), .B(new_n750_), .Y(new_n3168_));
  NOR2  g02783(.A(new_n3168_), .B(new_n756_), .Y(new_n3169_));
  NOR2  g02784(.A(new_n3169_), .B(new_n760_), .Y(new_n3170_));
  NOR2  g02785(.A(new_n3170_), .B(new_n766_), .Y(new_n3171_));
  NOR2  g02786(.A(new_n3171_), .B(new_n770_), .Y(new_n3172_));
  NOR2  g02787(.A(new_n3172_), .B(new_n776_), .Y(new_n3173_));
  NOR2  g02788(.A(new_n3173_), .B(new_n780_), .Y(new_n3174_));
  NOR2  g02789(.A(new_n3174_), .B(new_n786_), .Y(new_n3175_));
  NOR2  g02790(.A(new_n3175_), .B(new_n790_), .Y(new_n3176_));
  NOR2  g02791(.A(new_n3176_), .B(new_n796_), .Y(new_n3177_));
  NOR2  g02792(.A(new_n3177_), .B(new_n800_), .Y(new_n3178_));
  NOR2  g02793(.A(new_n3178_), .B(new_n806_), .Y(new_n3179_));
  NOR2  g02794(.A(new_n3179_), .B(new_n1616_), .Y(new_n3180_));
  NOR2  g02795(.A(new_n3180_), .B(new_n1618_), .Y(new_n3181_));
  NOR2  g02796(.A(new_n3181_), .B(new_n1885_), .Y(new_n3182_));
  NOR2  g02797(.A(new_n3182_), .B(new_n820_), .Y(new_n3183_));
  NOR2  g02798(.A(new_n3183_), .B(new_n824_), .Y(new_n3184_));
  NOR2  g02799(.A(new_n3184_), .B(new_n829_), .Y(new_n3185_));
  NOR2  g02800(.A(new_n3185_), .B(new_n833_), .Y(new_n3186_));
  NOR2  g02801(.A(new_n3186_), .B(new_n838_), .Y(new_n3187_));
  NOR2  g02802(.A(new_n3187_), .B(new_n842_), .Y(new_n3188_));
  NOR2  g02803(.A(new_n3188_), .B(new_n847_), .Y(new_n3189_));
  NOR2  g02804(.A(new_n3189_), .B(new_n851_), .Y(new_n3190_));
  NOR2  g02805(.A(new_n3190_), .B(new_n856_), .Y(new_n3191_));
  NOR2  g02806(.A(new_n3191_), .B(new_n860_), .Y(new_n3192_));
  NOR2  g02807(.A(new_n3192_), .B(new_n865_), .Y(new_n3193_));
  NAND2 g02808(.A(new_n867_), .B(\req[21] ), .Y(new_n3194_));
  NOR2  g02809(.A(new_n3194_), .B(new_n3193_), .Y(\grant[21] ));
  INV   g02810(.A(new_n877_), .Y(new_n3196_));
  NOR2  g02811(.A(new_n1246_), .B(new_n3196_), .Y(new_n3197_));
  NOR2  g02812(.A(new_n3197_), .B(new_n883_), .Y(new_n3198_));
  NOR2  g02813(.A(new_n3198_), .B(new_n887_), .Y(new_n3199_));
  NOR2  g02814(.A(new_n3199_), .B(new_n892_), .Y(new_n3200_));
  NOR2  g02815(.A(new_n3200_), .B(new_n896_), .Y(new_n3201_));
  NOR2  g02816(.A(new_n3201_), .B(new_n901_), .Y(new_n3202_));
  NOR2  g02817(.A(new_n3202_), .B(new_n905_), .Y(new_n3203_));
  NOR2  g02818(.A(new_n3203_), .B(new_n910_), .Y(new_n3204_));
  NOR2  g02819(.A(new_n3204_), .B(new_n914_), .Y(new_n3205_));
  NOR2  g02820(.A(new_n3205_), .B(new_n919_), .Y(new_n3206_));
  NOR2  g02821(.A(new_n3206_), .B(new_n923_), .Y(new_n3207_));
  NOR2  g02822(.A(new_n3207_), .B(new_n928_), .Y(new_n3208_));
  NOR2  g02823(.A(new_n3208_), .B(new_n932_), .Y(new_n3209_));
  NOR2  g02824(.A(new_n3209_), .B(new_n937_), .Y(new_n3210_));
  NOR2  g02825(.A(new_n3210_), .B(new_n941_), .Y(new_n3211_));
  NOR2  g02826(.A(new_n3211_), .B(new_n946_), .Y(new_n3212_));
  NOR2  g02827(.A(new_n3212_), .B(new_n950_), .Y(new_n3213_));
  NOR2  g02828(.A(new_n3213_), .B(new_n955_), .Y(new_n3214_));
  NOR2  g02829(.A(new_n3214_), .B(new_n959_), .Y(new_n3215_));
  NOR2  g02830(.A(new_n3215_), .B(new_n964_), .Y(new_n3216_));
  NOR2  g02831(.A(new_n3216_), .B(new_n968_), .Y(new_n3217_));
  NOR2  g02832(.A(new_n3217_), .B(new_n973_), .Y(new_n3218_));
  NOR2  g02833(.A(new_n3218_), .B(new_n977_), .Y(new_n3219_));
  NOR2  g02834(.A(new_n3219_), .B(new_n982_), .Y(new_n3220_));
  NOR2  g02835(.A(new_n3220_), .B(new_n986_), .Y(new_n3221_));
  NOR2  g02836(.A(new_n3221_), .B(new_n991_), .Y(new_n3222_));
  NOR2  g02837(.A(new_n3222_), .B(new_n995_), .Y(new_n3223_));
  NOR2  g02838(.A(new_n3223_), .B(new_n1000_), .Y(new_n3224_));
  NOR2  g02839(.A(new_n3224_), .B(new_n1004_), .Y(new_n3225_));
  NOR2  g02840(.A(new_n3225_), .B(new_n1009_), .Y(new_n3226_));
  NOR2  g02841(.A(new_n3226_), .B(new_n1013_), .Y(new_n3227_));
  NOR2  g02842(.A(new_n3227_), .B(new_n1018_), .Y(new_n3228_));
  NOR2  g02843(.A(new_n3228_), .B(new_n1022_), .Y(new_n3229_));
  NOR2  g02844(.A(new_n3229_), .B(new_n1027_), .Y(new_n3230_));
  NOR2  g02845(.A(new_n3230_), .B(new_n1031_), .Y(new_n3231_));
  NOR2  g02846(.A(new_n3231_), .B(new_n1036_), .Y(new_n3232_));
  NOR2  g02847(.A(new_n3232_), .B(new_n1040_), .Y(new_n3233_));
  NOR2  g02848(.A(new_n3233_), .B(new_n1045_), .Y(new_n3234_));
  NOR2  g02849(.A(new_n3234_), .B(new_n1049_), .Y(new_n3235_));
  NOR2  g02850(.A(new_n3235_), .B(new_n1054_), .Y(new_n3236_));
  NOR2  g02851(.A(new_n3236_), .B(new_n1058_), .Y(new_n3237_));
  NOR2  g02852(.A(new_n3237_), .B(new_n1063_), .Y(new_n3238_));
  NOR2  g02853(.A(new_n3238_), .B(new_n1067_), .Y(new_n3239_));
  NOR2  g02854(.A(new_n3239_), .B(new_n1072_), .Y(new_n3240_));
  NOR2  g02855(.A(new_n3240_), .B(new_n1076_), .Y(new_n3241_));
  NOR2  g02856(.A(new_n3241_), .B(new_n1081_), .Y(new_n3242_));
  NOR2  g02857(.A(new_n3242_), .B(new_n1085_), .Y(new_n3243_));
  NOR2  g02858(.A(new_n3243_), .B(new_n1090_), .Y(new_n3244_));
  NOR2  g02859(.A(new_n3244_), .B(new_n1094_), .Y(new_n3245_));
  NOR2  g02860(.A(new_n3245_), .B(new_n1099_), .Y(new_n3246_));
  NOR2  g02861(.A(new_n3246_), .B(new_n1103_), .Y(new_n3247_));
  NOR2  g02862(.A(new_n3247_), .B(new_n1108_), .Y(new_n3248_));
  NOR2  g02863(.A(new_n3248_), .B(new_n1112_), .Y(new_n3249_));
  NOR2  g02864(.A(new_n3249_), .B(new_n1117_), .Y(new_n3250_));
  NOR2  g02865(.A(new_n3250_), .B(new_n1121_), .Y(new_n3251_));
  NOR2  g02866(.A(new_n3251_), .B(new_n1126_), .Y(new_n3252_));
  NOR2  g02867(.A(new_n3252_), .B(new_n1130_), .Y(new_n3253_));
  NOR2  g02868(.A(new_n3253_), .B(new_n1135_), .Y(new_n3254_));
  NOR2  g02869(.A(new_n3254_), .B(new_n1139_), .Y(new_n3255_));
  NOR2  g02870(.A(new_n3255_), .B(new_n1144_), .Y(new_n3256_));
  NOR2  g02871(.A(new_n3256_), .B(new_n1148_), .Y(new_n3257_));
  NOR2  g02872(.A(new_n3257_), .B(new_n1153_), .Y(new_n3258_));
  NOR2  g02873(.A(new_n3258_), .B(new_n1157_), .Y(new_n3259_));
  NOR2  g02874(.A(new_n3259_), .B(new_n1162_), .Y(new_n3260_));
  NOR2  g02875(.A(new_n3260_), .B(new_n1166_), .Y(new_n3261_));
  NOR2  g02876(.A(new_n3261_), .B(new_n1171_), .Y(new_n3262_));
  NOR2  g02877(.A(new_n3262_), .B(new_n1175_), .Y(new_n3263_));
  NOR2  g02878(.A(new_n3263_), .B(new_n1180_), .Y(new_n3264_));
  NOR2  g02879(.A(new_n3264_), .B(new_n1184_), .Y(new_n3265_));
  NOR2  g02880(.A(new_n3265_), .B(new_n1189_), .Y(new_n3266_));
  NOR2  g02881(.A(new_n3266_), .B(new_n1707_), .Y(new_n3267_));
  NOR2  g02882(.A(new_n3267_), .B(new_n1709_), .Y(new_n3268_));
  NOR2  g02883(.A(new_n3268_), .B(new_n1973_), .Y(new_n3269_));
  NOR2  g02884(.A(new_n3269_), .B(new_n1199_), .Y(new_n3270_));
  NOR2  g02885(.A(new_n3270_), .B(new_n1203_), .Y(new_n3271_));
  NOR2  g02886(.A(new_n3271_), .B(new_n1207_), .Y(new_n3272_));
  NOR2  g02887(.A(new_n3272_), .B(new_n1211_), .Y(new_n3273_));
  NOR2  g02888(.A(new_n3273_), .B(new_n1215_), .Y(new_n3274_));
  NOR2  g02889(.A(new_n3274_), .B(new_n1219_), .Y(new_n3275_));
  NOR2  g02890(.A(new_n3275_), .B(new_n1223_), .Y(new_n3276_));
  NOR2  g02891(.A(new_n3276_), .B(new_n1227_), .Y(new_n3277_));
  NOR2  g02892(.A(new_n3277_), .B(new_n1231_), .Y(new_n3278_));
  NOR2  g02893(.A(new_n3278_), .B(new_n1235_), .Y(new_n3279_));
  NOR2  g02894(.A(new_n3279_), .B(new_n1239_), .Y(new_n3280_));
  NAND2 g02895(.A(new_n1241_), .B(\req[22] ), .Y(new_n3281_));
  NOR2  g02896(.A(new_n3281_), .B(new_n3280_), .Y(\grant[22] ));
  INV   g02897(.A(new_n1250_), .Y(new_n3283_));
  NOR2  g02898(.A(new_n3283_), .B(new_n465_), .Y(new_n3284_));
  NOR2  g02899(.A(new_n3284_), .B(new_n1255_), .Y(new_n3285_));
  NOR2  g02900(.A(new_n3285_), .B(new_n1259_), .Y(new_n3286_));
  NOR2  g02901(.A(new_n3286_), .B(new_n1263_), .Y(new_n3287_));
  NOR2  g02902(.A(new_n3287_), .B(new_n1267_), .Y(new_n3288_));
  NOR2  g02903(.A(new_n3288_), .B(new_n1271_), .Y(new_n3289_));
  NOR2  g02904(.A(new_n3289_), .B(new_n1275_), .Y(new_n3290_));
  NOR2  g02905(.A(new_n3290_), .B(new_n1279_), .Y(new_n3291_));
  NOR2  g02906(.A(new_n3291_), .B(new_n1283_), .Y(new_n3292_));
  NOR2  g02907(.A(new_n3292_), .B(new_n1287_), .Y(new_n3293_));
  NOR2  g02908(.A(new_n3293_), .B(new_n1291_), .Y(new_n3294_));
  NOR2  g02909(.A(new_n3294_), .B(new_n1295_), .Y(new_n3295_));
  NOR2  g02910(.A(new_n3295_), .B(new_n1299_), .Y(new_n3296_));
  NOR2  g02911(.A(new_n3296_), .B(new_n1303_), .Y(new_n3297_));
  NOR2  g02912(.A(new_n3297_), .B(new_n1307_), .Y(new_n3298_));
  NOR2  g02913(.A(new_n3298_), .B(new_n1311_), .Y(new_n3299_));
  NOR2  g02914(.A(new_n3299_), .B(new_n1315_), .Y(new_n3300_));
  NOR2  g02915(.A(new_n3300_), .B(new_n1319_), .Y(new_n3301_));
  NOR2  g02916(.A(new_n3301_), .B(new_n1323_), .Y(new_n3302_));
  NOR2  g02917(.A(new_n3302_), .B(new_n1327_), .Y(new_n3303_));
  NOR2  g02918(.A(new_n3303_), .B(new_n1331_), .Y(new_n3304_));
  NOR2  g02919(.A(new_n3304_), .B(new_n1335_), .Y(new_n3305_));
  NOR2  g02920(.A(new_n3305_), .B(new_n1339_), .Y(new_n3306_));
  NOR2  g02921(.A(new_n3306_), .B(new_n1343_), .Y(new_n3307_));
  NOR2  g02922(.A(new_n3307_), .B(new_n1347_), .Y(new_n3308_));
  NOR2  g02923(.A(new_n3308_), .B(new_n1351_), .Y(new_n3309_));
  NOR2  g02924(.A(new_n3309_), .B(new_n1355_), .Y(new_n3310_));
  NOR2  g02925(.A(new_n3310_), .B(new_n1359_), .Y(new_n3311_));
  NOR2  g02926(.A(new_n3311_), .B(new_n1363_), .Y(new_n3312_));
  NOR2  g02927(.A(new_n3312_), .B(new_n1367_), .Y(new_n3313_));
  NOR2  g02928(.A(new_n3313_), .B(new_n1371_), .Y(new_n3314_));
  NOR2  g02929(.A(new_n3314_), .B(new_n1375_), .Y(new_n3315_));
  NOR2  g02930(.A(new_n3315_), .B(new_n1379_), .Y(new_n3316_));
  NOR2  g02931(.A(new_n3316_), .B(new_n1383_), .Y(new_n3317_));
  NOR2  g02932(.A(new_n3317_), .B(new_n1387_), .Y(new_n3318_));
  NOR2  g02933(.A(new_n3318_), .B(new_n1391_), .Y(new_n3319_));
  NOR2  g02934(.A(new_n3319_), .B(new_n1395_), .Y(new_n3320_));
  NOR2  g02935(.A(new_n3320_), .B(new_n1399_), .Y(new_n3321_));
  NOR2  g02936(.A(new_n3321_), .B(new_n1403_), .Y(new_n3322_));
  NOR2  g02937(.A(new_n3322_), .B(new_n1407_), .Y(new_n3323_));
  NOR2  g02938(.A(new_n3323_), .B(new_n1411_), .Y(new_n3324_));
  NOR2  g02939(.A(new_n3324_), .B(new_n1415_), .Y(new_n3325_));
  NOR2  g02940(.A(new_n3325_), .B(new_n1419_), .Y(new_n3326_));
  NOR2  g02941(.A(new_n3326_), .B(new_n1423_), .Y(new_n3327_));
  NOR2  g02942(.A(new_n3327_), .B(new_n1427_), .Y(new_n3328_));
  NOR2  g02943(.A(new_n3328_), .B(new_n1431_), .Y(new_n3329_));
  NOR2  g02944(.A(new_n3329_), .B(new_n1435_), .Y(new_n3330_));
  NOR2  g02945(.A(new_n3330_), .B(new_n1439_), .Y(new_n3331_));
  NOR2  g02946(.A(new_n3331_), .B(new_n1443_), .Y(new_n3332_));
  NOR2  g02947(.A(new_n3332_), .B(new_n1447_), .Y(new_n3333_));
  NOR2  g02948(.A(new_n3333_), .B(new_n1451_), .Y(new_n3334_));
  NOR2  g02949(.A(new_n3334_), .B(new_n1455_), .Y(new_n3335_));
  NOR2  g02950(.A(new_n3335_), .B(new_n1459_), .Y(new_n3336_));
  NOR2  g02951(.A(new_n3336_), .B(new_n1463_), .Y(new_n3337_));
  NOR2  g02952(.A(new_n3337_), .B(new_n1467_), .Y(new_n3338_));
  NOR2  g02953(.A(new_n3338_), .B(new_n1471_), .Y(new_n3339_));
  NOR2  g02954(.A(new_n3339_), .B(new_n1475_), .Y(new_n3340_));
  NOR2  g02955(.A(new_n3340_), .B(new_n1479_), .Y(new_n3341_));
  NOR2  g02956(.A(new_n3341_), .B(new_n1483_), .Y(new_n3342_));
  NOR2  g02957(.A(new_n3342_), .B(new_n1487_), .Y(new_n3343_));
  NOR2  g02958(.A(new_n3343_), .B(new_n1491_), .Y(new_n3344_));
  NOR2  g02959(.A(new_n3344_), .B(new_n1495_), .Y(new_n3345_));
  NOR2  g02960(.A(new_n3345_), .B(new_n1499_), .Y(new_n3346_));
  NOR2  g02961(.A(new_n3346_), .B(new_n1503_), .Y(new_n3347_));
  NOR2  g02962(.A(new_n3347_), .B(new_n1507_), .Y(new_n3348_));
  NOR2  g02963(.A(new_n3348_), .B(new_n1511_), .Y(new_n3349_));
  NOR2  g02964(.A(new_n3349_), .B(new_n1515_), .Y(new_n3350_));
  NOR2  g02965(.A(new_n3350_), .B(new_n1519_), .Y(new_n3351_));
  NOR2  g02966(.A(new_n3351_), .B(new_n1523_), .Y(new_n3352_));
  NOR2  g02967(.A(new_n3352_), .B(new_n1527_), .Y(new_n3353_));
  NOR2  g02968(.A(new_n3353_), .B(new_n1797_), .Y(new_n3354_));
  NOR2  g02969(.A(new_n3354_), .B(new_n396_), .Y(new_n3355_));
  NOR2  g02970(.A(new_n3355_), .B(new_n400_), .Y(new_n3356_));
  NOR2  g02971(.A(new_n3356_), .B(new_n406_), .Y(new_n3357_));
  NOR2  g02972(.A(new_n3357_), .B(new_n410_), .Y(new_n3358_));
  NOR2  g02973(.A(new_n3358_), .B(new_n416_), .Y(new_n3359_));
  NOR2  g02974(.A(new_n3359_), .B(new_n420_), .Y(new_n3360_));
  NOR2  g02975(.A(new_n3360_), .B(new_n426_), .Y(new_n3361_));
  NOR2  g02976(.A(new_n3361_), .B(new_n430_), .Y(new_n3362_));
  NOR2  g02977(.A(new_n3362_), .B(new_n436_), .Y(new_n3363_));
  NOR2  g02978(.A(new_n3363_), .B(new_n440_), .Y(new_n3364_));
  NOR2  g02979(.A(new_n3364_), .B(new_n446_), .Y(new_n3365_));
  NOR2  g02980(.A(new_n3365_), .B(new_n450_), .Y(new_n3366_));
  NOR2  g02981(.A(new_n3366_), .B(new_n456_), .Y(new_n3367_));
  NAND2 g02982(.A(new_n458_), .B(\req[23] ), .Y(new_n3368_));
  NOR2  g02983(.A(new_n3368_), .B(new_n3367_), .Y(\grant[23] ));
  INV   g02984(.A(new_n469_), .Y(new_n3370_));
  NOR2  g02985(.A(new_n882_), .B(new_n3370_), .Y(new_n3371_));
  NOR2  g02986(.A(new_n3371_), .B(new_n476_), .Y(new_n3372_));
  NOR2  g02987(.A(new_n3372_), .B(new_n480_), .Y(new_n3373_));
  NOR2  g02988(.A(new_n3373_), .B(new_n486_), .Y(new_n3374_));
  NOR2  g02989(.A(new_n3374_), .B(new_n490_), .Y(new_n3375_));
  NOR2  g02990(.A(new_n3375_), .B(new_n496_), .Y(new_n3376_));
  NOR2  g02991(.A(new_n3376_), .B(new_n500_), .Y(new_n3377_));
  NOR2  g02992(.A(new_n3377_), .B(new_n506_), .Y(new_n3378_));
  NOR2  g02993(.A(new_n3378_), .B(new_n510_), .Y(new_n3379_));
  NOR2  g02994(.A(new_n3379_), .B(new_n516_), .Y(new_n3380_));
  NOR2  g02995(.A(new_n3380_), .B(new_n520_), .Y(new_n3381_));
  NOR2  g02996(.A(new_n3381_), .B(new_n526_), .Y(new_n3382_));
  NOR2  g02997(.A(new_n3382_), .B(new_n530_), .Y(new_n3383_));
  NOR2  g02998(.A(new_n3383_), .B(new_n536_), .Y(new_n3384_));
  NOR2  g02999(.A(new_n3384_), .B(new_n540_), .Y(new_n3385_));
  NOR2  g03000(.A(new_n3385_), .B(new_n546_), .Y(new_n3386_));
  NOR2  g03001(.A(new_n3386_), .B(new_n550_), .Y(new_n3387_));
  NOR2  g03002(.A(new_n3387_), .B(new_n556_), .Y(new_n3388_));
  NOR2  g03003(.A(new_n3388_), .B(new_n560_), .Y(new_n3389_));
  NOR2  g03004(.A(new_n3389_), .B(new_n566_), .Y(new_n3390_));
  NOR2  g03005(.A(new_n3390_), .B(new_n570_), .Y(new_n3391_));
  NOR2  g03006(.A(new_n3391_), .B(new_n576_), .Y(new_n3392_));
  NOR2  g03007(.A(new_n3392_), .B(new_n580_), .Y(new_n3393_));
  NOR2  g03008(.A(new_n3393_), .B(new_n586_), .Y(new_n3394_));
  NOR2  g03009(.A(new_n3394_), .B(new_n590_), .Y(new_n3395_));
  NOR2  g03010(.A(new_n3395_), .B(new_n596_), .Y(new_n3396_));
  NOR2  g03011(.A(new_n3396_), .B(new_n600_), .Y(new_n3397_));
  NOR2  g03012(.A(new_n3397_), .B(new_n606_), .Y(new_n3398_));
  NOR2  g03013(.A(new_n3398_), .B(new_n610_), .Y(new_n3399_));
  NOR2  g03014(.A(new_n3399_), .B(new_n616_), .Y(new_n3400_));
  NOR2  g03015(.A(new_n3400_), .B(new_n620_), .Y(new_n3401_));
  NOR2  g03016(.A(new_n3401_), .B(new_n626_), .Y(new_n3402_));
  NOR2  g03017(.A(new_n3402_), .B(new_n630_), .Y(new_n3403_));
  NOR2  g03018(.A(new_n3403_), .B(new_n636_), .Y(new_n3404_));
  NOR2  g03019(.A(new_n3404_), .B(new_n640_), .Y(new_n3405_));
  NOR2  g03020(.A(new_n3405_), .B(new_n646_), .Y(new_n3406_));
  NOR2  g03021(.A(new_n3406_), .B(new_n650_), .Y(new_n3407_));
  NOR2  g03022(.A(new_n3407_), .B(new_n656_), .Y(new_n3408_));
  NOR2  g03023(.A(new_n3408_), .B(new_n660_), .Y(new_n3409_));
  NOR2  g03024(.A(new_n3409_), .B(new_n666_), .Y(new_n3410_));
  NOR2  g03025(.A(new_n3410_), .B(new_n670_), .Y(new_n3411_));
  NOR2  g03026(.A(new_n3411_), .B(new_n676_), .Y(new_n3412_));
  NOR2  g03027(.A(new_n3412_), .B(new_n680_), .Y(new_n3413_));
  NOR2  g03028(.A(new_n3413_), .B(new_n686_), .Y(new_n3414_));
  NOR2  g03029(.A(new_n3414_), .B(new_n690_), .Y(new_n3415_));
  NOR2  g03030(.A(new_n3415_), .B(new_n696_), .Y(new_n3416_));
  NOR2  g03031(.A(new_n3416_), .B(new_n700_), .Y(new_n3417_));
  NOR2  g03032(.A(new_n3417_), .B(new_n706_), .Y(new_n3418_));
  NOR2  g03033(.A(new_n3418_), .B(new_n710_), .Y(new_n3419_));
  NOR2  g03034(.A(new_n3419_), .B(new_n716_), .Y(new_n3420_));
  NOR2  g03035(.A(new_n3420_), .B(new_n720_), .Y(new_n3421_));
  NOR2  g03036(.A(new_n3421_), .B(new_n726_), .Y(new_n3422_));
  NOR2  g03037(.A(new_n3422_), .B(new_n730_), .Y(new_n3423_));
  NOR2  g03038(.A(new_n3423_), .B(new_n736_), .Y(new_n3424_));
  NOR2  g03039(.A(new_n3424_), .B(new_n740_), .Y(new_n3425_));
  NOR2  g03040(.A(new_n3425_), .B(new_n746_), .Y(new_n3426_));
  NOR2  g03041(.A(new_n3426_), .B(new_n750_), .Y(new_n3427_));
  NOR2  g03042(.A(new_n3427_), .B(new_n756_), .Y(new_n3428_));
  NOR2  g03043(.A(new_n3428_), .B(new_n760_), .Y(new_n3429_));
  NOR2  g03044(.A(new_n3429_), .B(new_n766_), .Y(new_n3430_));
  NOR2  g03045(.A(new_n3430_), .B(new_n770_), .Y(new_n3431_));
  NOR2  g03046(.A(new_n3431_), .B(new_n776_), .Y(new_n3432_));
  NOR2  g03047(.A(new_n3432_), .B(new_n780_), .Y(new_n3433_));
  NOR2  g03048(.A(new_n3433_), .B(new_n786_), .Y(new_n3434_));
  NOR2  g03049(.A(new_n3434_), .B(new_n790_), .Y(new_n3435_));
  NOR2  g03050(.A(new_n3435_), .B(new_n796_), .Y(new_n3436_));
  NOR2  g03051(.A(new_n3436_), .B(new_n800_), .Y(new_n3437_));
  NOR2  g03052(.A(new_n3437_), .B(new_n806_), .Y(new_n3438_));
  NOR2  g03053(.A(new_n3438_), .B(new_n1616_), .Y(new_n3439_));
  NOR2  g03054(.A(new_n3439_), .B(new_n1618_), .Y(new_n3440_));
  NOR2  g03055(.A(new_n3440_), .B(new_n1885_), .Y(new_n3441_));
  NOR2  g03056(.A(new_n3441_), .B(new_n820_), .Y(new_n3442_));
  NOR2  g03057(.A(new_n3442_), .B(new_n824_), .Y(new_n3443_));
  NOR2  g03058(.A(new_n3443_), .B(new_n829_), .Y(new_n3444_));
  NOR2  g03059(.A(new_n3444_), .B(new_n833_), .Y(new_n3445_));
  NOR2  g03060(.A(new_n3445_), .B(new_n838_), .Y(new_n3446_));
  NOR2  g03061(.A(new_n3446_), .B(new_n842_), .Y(new_n3447_));
  NOR2  g03062(.A(new_n3447_), .B(new_n847_), .Y(new_n3448_));
  NOR2  g03063(.A(new_n3448_), .B(new_n851_), .Y(new_n3449_));
  NOR2  g03064(.A(new_n3449_), .B(new_n856_), .Y(new_n3450_));
  NOR2  g03065(.A(new_n3450_), .B(new_n860_), .Y(new_n3451_));
  NOR2  g03066(.A(new_n3451_), .B(new_n865_), .Y(new_n3452_));
  NOR2  g03067(.A(new_n3452_), .B(new_n869_), .Y(new_n3453_));
  NOR2  g03068(.A(new_n3453_), .B(new_n874_), .Y(new_n3454_));
  NAND2 g03069(.A(new_n876_), .B(\req[24] ), .Y(new_n3455_));
  NOR2  g03070(.A(new_n3455_), .B(new_n3454_), .Y(\grant[24] ));
  INV   g03071(.A(new_n886_), .Y(new_n3457_));
  NOR2  g03072(.A(new_n1254_), .B(new_n3457_), .Y(new_n3458_));
  NOR2  g03073(.A(new_n3458_), .B(new_n892_), .Y(new_n3459_));
  NOR2  g03074(.A(new_n3459_), .B(new_n896_), .Y(new_n3460_));
  NOR2  g03075(.A(new_n3460_), .B(new_n901_), .Y(new_n3461_));
  NOR2  g03076(.A(new_n3461_), .B(new_n905_), .Y(new_n3462_));
  NOR2  g03077(.A(new_n3462_), .B(new_n910_), .Y(new_n3463_));
  NOR2  g03078(.A(new_n3463_), .B(new_n914_), .Y(new_n3464_));
  NOR2  g03079(.A(new_n3464_), .B(new_n919_), .Y(new_n3465_));
  NOR2  g03080(.A(new_n3465_), .B(new_n923_), .Y(new_n3466_));
  NOR2  g03081(.A(new_n3466_), .B(new_n928_), .Y(new_n3467_));
  NOR2  g03082(.A(new_n3467_), .B(new_n932_), .Y(new_n3468_));
  NOR2  g03083(.A(new_n3468_), .B(new_n937_), .Y(new_n3469_));
  NOR2  g03084(.A(new_n3469_), .B(new_n941_), .Y(new_n3470_));
  NOR2  g03085(.A(new_n3470_), .B(new_n946_), .Y(new_n3471_));
  NOR2  g03086(.A(new_n3471_), .B(new_n950_), .Y(new_n3472_));
  NOR2  g03087(.A(new_n3472_), .B(new_n955_), .Y(new_n3473_));
  NOR2  g03088(.A(new_n3473_), .B(new_n959_), .Y(new_n3474_));
  NOR2  g03089(.A(new_n3474_), .B(new_n964_), .Y(new_n3475_));
  NOR2  g03090(.A(new_n3475_), .B(new_n968_), .Y(new_n3476_));
  NOR2  g03091(.A(new_n3476_), .B(new_n973_), .Y(new_n3477_));
  NOR2  g03092(.A(new_n3477_), .B(new_n977_), .Y(new_n3478_));
  NOR2  g03093(.A(new_n3478_), .B(new_n982_), .Y(new_n3479_));
  NOR2  g03094(.A(new_n3479_), .B(new_n986_), .Y(new_n3480_));
  NOR2  g03095(.A(new_n3480_), .B(new_n991_), .Y(new_n3481_));
  NOR2  g03096(.A(new_n3481_), .B(new_n995_), .Y(new_n3482_));
  NOR2  g03097(.A(new_n3482_), .B(new_n1000_), .Y(new_n3483_));
  NOR2  g03098(.A(new_n3483_), .B(new_n1004_), .Y(new_n3484_));
  NOR2  g03099(.A(new_n3484_), .B(new_n1009_), .Y(new_n3485_));
  NOR2  g03100(.A(new_n3485_), .B(new_n1013_), .Y(new_n3486_));
  NOR2  g03101(.A(new_n3486_), .B(new_n1018_), .Y(new_n3487_));
  NOR2  g03102(.A(new_n3487_), .B(new_n1022_), .Y(new_n3488_));
  NOR2  g03103(.A(new_n3488_), .B(new_n1027_), .Y(new_n3489_));
  NOR2  g03104(.A(new_n3489_), .B(new_n1031_), .Y(new_n3490_));
  NOR2  g03105(.A(new_n3490_), .B(new_n1036_), .Y(new_n3491_));
  NOR2  g03106(.A(new_n3491_), .B(new_n1040_), .Y(new_n3492_));
  NOR2  g03107(.A(new_n3492_), .B(new_n1045_), .Y(new_n3493_));
  NOR2  g03108(.A(new_n3493_), .B(new_n1049_), .Y(new_n3494_));
  NOR2  g03109(.A(new_n3494_), .B(new_n1054_), .Y(new_n3495_));
  NOR2  g03110(.A(new_n3495_), .B(new_n1058_), .Y(new_n3496_));
  NOR2  g03111(.A(new_n3496_), .B(new_n1063_), .Y(new_n3497_));
  NOR2  g03112(.A(new_n3497_), .B(new_n1067_), .Y(new_n3498_));
  NOR2  g03113(.A(new_n3498_), .B(new_n1072_), .Y(new_n3499_));
  NOR2  g03114(.A(new_n3499_), .B(new_n1076_), .Y(new_n3500_));
  NOR2  g03115(.A(new_n3500_), .B(new_n1081_), .Y(new_n3501_));
  NOR2  g03116(.A(new_n3501_), .B(new_n1085_), .Y(new_n3502_));
  NOR2  g03117(.A(new_n3502_), .B(new_n1090_), .Y(new_n3503_));
  NOR2  g03118(.A(new_n3503_), .B(new_n1094_), .Y(new_n3504_));
  NOR2  g03119(.A(new_n3504_), .B(new_n1099_), .Y(new_n3505_));
  NOR2  g03120(.A(new_n3505_), .B(new_n1103_), .Y(new_n3506_));
  NOR2  g03121(.A(new_n3506_), .B(new_n1108_), .Y(new_n3507_));
  NOR2  g03122(.A(new_n3507_), .B(new_n1112_), .Y(new_n3508_));
  NOR2  g03123(.A(new_n3508_), .B(new_n1117_), .Y(new_n3509_));
  NOR2  g03124(.A(new_n3509_), .B(new_n1121_), .Y(new_n3510_));
  NOR2  g03125(.A(new_n3510_), .B(new_n1126_), .Y(new_n3511_));
  NOR2  g03126(.A(new_n3511_), .B(new_n1130_), .Y(new_n3512_));
  NOR2  g03127(.A(new_n3512_), .B(new_n1135_), .Y(new_n3513_));
  NOR2  g03128(.A(new_n3513_), .B(new_n1139_), .Y(new_n3514_));
  NOR2  g03129(.A(new_n3514_), .B(new_n1144_), .Y(new_n3515_));
  NOR2  g03130(.A(new_n3515_), .B(new_n1148_), .Y(new_n3516_));
  NOR2  g03131(.A(new_n3516_), .B(new_n1153_), .Y(new_n3517_));
  NOR2  g03132(.A(new_n3517_), .B(new_n1157_), .Y(new_n3518_));
  NOR2  g03133(.A(new_n3518_), .B(new_n1162_), .Y(new_n3519_));
  NOR2  g03134(.A(new_n3519_), .B(new_n1166_), .Y(new_n3520_));
  NOR2  g03135(.A(new_n3520_), .B(new_n1171_), .Y(new_n3521_));
  NOR2  g03136(.A(new_n3521_), .B(new_n1175_), .Y(new_n3522_));
  NOR2  g03137(.A(new_n3522_), .B(new_n1180_), .Y(new_n3523_));
  NOR2  g03138(.A(new_n3523_), .B(new_n1184_), .Y(new_n3524_));
  NOR2  g03139(.A(new_n3524_), .B(new_n1189_), .Y(new_n3525_));
  NOR2  g03140(.A(new_n3525_), .B(new_n1707_), .Y(new_n3526_));
  NOR2  g03141(.A(new_n3526_), .B(new_n1709_), .Y(new_n3527_));
  NOR2  g03142(.A(new_n3527_), .B(new_n1973_), .Y(new_n3528_));
  NOR2  g03143(.A(new_n3528_), .B(new_n1199_), .Y(new_n3529_));
  NOR2  g03144(.A(new_n3529_), .B(new_n1203_), .Y(new_n3530_));
  NOR2  g03145(.A(new_n3530_), .B(new_n1207_), .Y(new_n3531_));
  NOR2  g03146(.A(new_n3531_), .B(new_n1211_), .Y(new_n3532_));
  NOR2  g03147(.A(new_n3532_), .B(new_n1215_), .Y(new_n3533_));
  NOR2  g03148(.A(new_n3533_), .B(new_n1219_), .Y(new_n3534_));
  NOR2  g03149(.A(new_n3534_), .B(new_n1223_), .Y(new_n3535_));
  NOR2  g03150(.A(new_n3535_), .B(new_n1227_), .Y(new_n3536_));
  NOR2  g03151(.A(new_n3536_), .B(new_n1231_), .Y(new_n3537_));
  NOR2  g03152(.A(new_n3537_), .B(new_n1235_), .Y(new_n3538_));
  NOR2  g03153(.A(new_n3538_), .B(new_n1239_), .Y(new_n3539_));
  NOR2  g03154(.A(new_n3539_), .B(new_n1243_), .Y(new_n3540_));
  NOR2  g03155(.A(new_n3540_), .B(new_n1247_), .Y(new_n3541_));
  NAND2 g03156(.A(new_n1249_), .B(\req[25] ), .Y(new_n3542_));
  NOR2  g03157(.A(new_n3542_), .B(new_n3541_), .Y(\grant[25] ));
  INV   g03158(.A(new_n1258_), .Y(new_n3544_));
  NOR2  g03159(.A(new_n3544_), .B(new_n475_), .Y(new_n3545_));
  NOR2  g03160(.A(new_n3545_), .B(new_n1263_), .Y(new_n3546_));
  NOR2  g03161(.A(new_n3546_), .B(new_n1267_), .Y(new_n3547_));
  NOR2  g03162(.A(new_n3547_), .B(new_n1271_), .Y(new_n3548_));
  NOR2  g03163(.A(new_n3548_), .B(new_n1275_), .Y(new_n3549_));
  NOR2  g03164(.A(new_n3549_), .B(new_n1279_), .Y(new_n3550_));
  NOR2  g03165(.A(new_n3550_), .B(new_n1283_), .Y(new_n3551_));
  NOR2  g03166(.A(new_n3551_), .B(new_n1287_), .Y(new_n3552_));
  NOR2  g03167(.A(new_n3552_), .B(new_n1291_), .Y(new_n3553_));
  NOR2  g03168(.A(new_n3553_), .B(new_n1295_), .Y(new_n3554_));
  NOR2  g03169(.A(new_n3554_), .B(new_n1299_), .Y(new_n3555_));
  NOR2  g03170(.A(new_n3555_), .B(new_n1303_), .Y(new_n3556_));
  NOR2  g03171(.A(new_n3556_), .B(new_n1307_), .Y(new_n3557_));
  NOR2  g03172(.A(new_n3557_), .B(new_n1311_), .Y(new_n3558_));
  NOR2  g03173(.A(new_n3558_), .B(new_n1315_), .Y(new_n3559_));
  NOR2  g03174(.A(new_n3559_), .B(new_n1319_), .Y(new_n3560_));
  NOR2  g03175(.A(new_n3560_), .B(new_n1323_), .Y(new_n3561_));
  NOR2  g03176(.A(new_n3561_), .B(new_n1327_), .Y(new_n3562_));
  NOR2  g03177(.A(new_n3562_), .B(new_n1331_), .Y(new_n3563_));
  NOR2  g03178(.A(new_n3563_), .B(new_n1335_), .Y(new_n3564_));
  NOR2  g03179(.A(new_n3564_), .B(new_n1339_), .Y(new_n3565_));
  NOR2  g03180(.A(new_n3565_), .B(new_n1343_), .Y(new_n3566_));
  NOR2  g03181(.A(new_n3566_), .B(new_n1347_), .Y(new_n3567_));
  NOR2  g03182(.A(new_n3567_), .B(new_n1351_), .Y(new_n3568_));
  NOR2  g03183(.A(new_n3568_), .B(new_n1355_), .Y(new_n3569_));
  NOR2  g03184(.A(new_n3569_), .B(new_n1359_), .Y(new_n3570_));
  NOR2  g03185(.A(new_n3570_), .B(new_n1363_), .Y(new_n3571_));
  NOR2  g03186(.A(new_n3571_), .B(new_n1367_), .Y(new_n3572_));
  NOR2  g03187(.A(new_n3572_), .B(new_n1371_), .Y(new_n3573_));
  NOR2  g03188(.A(new_n3573_), .B(new_n1375_), .Y(new_n3574_));
  NOR2  g03189(.A(new_n3574_), .B(new_n1379_), .Y(new_n3575_));
  NOR2  g03190(.A(new_n3575_), .B(new_n1383_), .Y(new_n3576_));
  NOR2  g03191(.A(new_n3576_), .B(new_n1387_), .Y(new_n3577_));
  NOR2  g03192(.A(new_n3577_), .B(new_n1391_), .Y(new_n3578_));
  NOR2  g03193(.A(new_n3578_), .B(new_n1395_), .Y(new_n3579_));
  NOR2  g03194(.A(new_n3579_), .B(new_n1399_), .Y(new_n3580_));
  NOR2  g03195(.A(new_n3580_), .B(new_n1403_), .Y(new_n3581_));
  NOR2  g03196(.A(new_n3581_), .B(new_n1407_), .Y(new_n3582_));
  NOR2  g03197(.A(new_n3582_), .B(new_n1411_), .Y(new_n3583_));
  NOR2  g03198(.A(new_n3583_), .B(new_n1415_), .Y(new_n3584_));
  NOR2  g03199(.A(new_n3584_), .B(new_n1419_), .Y(new_n3585_));
  NOR2  g03200(.A(new_n3585_), .B(new_n1423_), .Y(new_n3586_));
  NOR2  g03201(.A(new_n3586_), .B(new_n1427_), .Y(new_n3587_));
  NOR2  g03202(.A(new_n3587_), .B(new_n1431_), .Y(new_n3588_));
  NOR2  g03203(.A(new_n3588_), .B(new_n1435_), .Y(new_n3589_));
  NOR2  g03204(.A(new_n3589_), .B(new_n1439_), .Y(new_n3590_));
  NOR2  g03205(.A(new_n3590_), .B(new_n1443_), .Y(new_n3591_));
  NOR2  g03206(.A(new_n3591_), .B(new_n1447_), .Y(new_n3592_));
  NOR2  g03207(.A(new_n3592_), .B(new_n1451_), .Y(new_n3593_));
  NOR2  g03208(.A(new_n3593_), .B(new_n1455_), .Y(new_n3594_));
  NOR2  g03209(.A(new_n3594_), .B(new_n1459_), .Y(new_n3595_));
  NOR2  g03210(.A(new_n3595_), .B(new_n1463_), .Y(new_n3596_));
  NOR2  g03211(.A(new_n3596_), .B(new_n1467_), .Y(new_n3597_));
  NOR2  g03212(.A(new_n3597_), .B(new_n1471_), .Y(new_n3598_));
  NOR2  g03213(.A(new_n3598_), .B(new_n1475_), .Y(new_n3599_));
  NOR2  g03214(.A(new_n3599_), .B(new_n1479_), .Y(new_n3600_));
  NOR2  g03215(.A(new_n3600_), .B(new_n1483_), .Y(new_n3601_));
  NOR2  g03216(.A(new_n3601_), .B(new_n1487_), .Y(new_n3602_));
  NOR2  g03217(.A(new_n3602_), .B(new_n1491_), .Y(new_n3603_));
  NOR2  g03218(.A(new_n3603_), .B(new_n1495_), .Y(new_n3604_));
  NOR2  g03219(.A(new_n3604_), .B(new_n1499_), .Y(new_n3605_));
  NOR2  g03220(.A(new_n3605_), .B(new_n1503_), .Y(new_n3606_));
  NOR2  g03221(.A(new_n3606_), .B(new_n1507_), .Y(new_n3607_));
  NOR2  g03222(.A(new_n3607_), .B(new_n1511_), .Y(new_n3608_));
  NOR2  g03223(.A(new_n3608_), .B(new_n1515_), .Y(new_n3609_));
  NOR2  g03224(.A(new_n3609_), .B(new_n1519_), .Y(new_n3610_));
  NOR2  g03225(.A(new_n3610_), .B(new_n1523_), .Y(new_n3611_));
  NOR2  g03226(.A(new_n3611_), .B(new_n1527_), .Y(new_n3612_));
  NOR2  g03227(.A(new_n3612_), .B(new_n1797_), .Y(new_n3613_));
  NOR2  g03228(.A(new_n3613_), .B(new_n396_), .Y(new_n3614_));
  NOR2  g03229(.A(new_n3614_), .B(new_n400_), .Y(new_n3615_));
  NOR2  g03230(.A(new_n3615_), .B(new_n406_), .Y(new_n3616_));
  NOR2  g03231(.A(new_n3616_), .B(new_n410_), .Y(new_n3617_));
  NOR2  g03232(.A(new_n3617_), .B(new_n416_), .Y(new_n3618_));
  NOR2  g03233(.A(new_n3618_), .B(new_n420_), .Y(new_n3619_));
  NOR2  g03234(.A(new_n3619_), .B(new_n426_), .Y(new_n3620_));
  NOR2  g03235(.A(new_n3620_), .B(new_n430_), .Y(new_n3621_));
  NOR2  g03236(.A(new_n3621_), .B(new_n436_), .Y(new_n3622_));
  NOR2  g03237(.A(new_n3622_), .B(new_n440_), .Y(new_n3623_));
  NOR2  g03238(.A(new_n3623_), .B(new_n446_), .Y(new_n3624_));
  NOR2  g03239(.A(new_n3624_), .B(new_n450_), .Y(new_n3625_));
  NOR2  g03240(.A(new_n3625_), .B(new_n456_), .Y(new_n3626_));
  NOR2  g03241(.A(new_n3626_), .B(new_n460_), .Y(new_n3627_));
  NOR2  g03242(.A(new_n3627_), .B(new_n466_), .Y(new_n3628_));
  NAND2 g03243(.A(new_n468_), .B(\req[26] ), .Y(new_n3629_));
  NOR2  g03244(.A(new_n3629_), .B(new_n3628_), .Y(\grant[26] ));
  INV   g03245(.A(new_n479_), .Y(new_n3631_));
  NOR2  g03246(.A(new_n891_), .B(new_n3631_), .Y(new_n3632_));
  NOR2  g03247(.A(new_n3632_), .B(new_n486_), .Y(new_n3633_));
  NOR2  g03248(.A(new_n3633_), .B(new_n490_), .Y(new_n3634_));
  NOR2  g03249(.A(new_n3634_), .B(new_n496_), .Y(new_n3635_));
  NOR2  g03250(.A(new_n3635_), .B(new_n500_), .Y(new_n3636_));
  NOR2  g03251(.A(new_n3636_), .B(new_n506_), .Y(new_n3637_));
  NOR2  g03252(.A(new_n3637_), .B(new_n510_), .Y(new_n3638_));
  NOR2  g03253(.A(new_n3638_), .B(new_n516_), .Y(new_n3639_));
  NOR2  g03254(.A(new_n3639_), .B(new_n520_), .Y(new_n3640_));
  NOR2  g03255(.A(new_n3640_), .B(new_n526_), .Y(new_n3641_));
  NOR2  g03256(.A(new_n3641_), .B(new_n530_), .Y(new_n3642_));
  NOR2  g03257(.A(new_n3642_), .B(new_n536_), .Y(new_n3643_));
  NOR2  g03258(.A(new_n3643_), .B(new_n540_), .Y(new_n3644_));
  NOR2  g03259(.A(new_n3644_), .B(new_n546_), .Y(new_n3645_));
  NOR2  g03260(.A(new_n3645_), .B(new_n550_), .Y(new_n3646_));
  NOR2  g03261(.A(new_n3646_), .B(new_n556_), .Y(new_n3647_));
  NOR2  g03262(.A(new_n3647_), .B(new_n560_), .Y(new_n3648_));
  NOR2  g03263(.A(new_n3648_), .B(new_n566_), .Y(new_n3649_));
  NOR2  g03264(.A(new_n3649_), .B(new_n570_), .Y(new_n3650_));
  NOR2  g03265(.A(new_n3650_), .B(new_n576_), .Y(new_n3651_));
  NOR2  g03266(.A(new_n3651_), .B(new_n580_), .Y(new_n3652_));
  NOR2  g03267(.A(new_n3652_), .B(new_n586_), .Y(new_n3653_));
  NOR2  g03268(.A(new_n3653_), .B(new_n590_), .Y(new_n3654_));
  NOR2  g03269(.A(new_n3654_), .B(new_n596_), .Y(new_n3655_));
  NOR2  g03270(.A(new_n3655_), .B(new_n600_), .Y(new_n3656_));
  NOR2  g03271(.A(new_n3656_), .B(new_n606_), .Y(new_n3657_));
  NOR2  g03272(.A(new_n3657_), .B(new_n610_), .Y(new_n3658_));
  NOR2  g03273(.A(new_n3658_), .B(new_n616_), .Y(new_n3659_));
  NOR2  g03274(.A(new_n3659_), .B(new_n620_), .Y(new_n3660_));
  NOR2  g03275(.A(new_n3660_), .B(new_n626_), .Y(new_n3661_));
  NOR2  g03276(.A(new_n3661_), .B(new_n630_), .Y(new_n3662_));
  NOR2  g03277(.A(new_n3662_), .B(new_n636_), .Y(new_n3663_));
  NOR2  g03278(.A(new_n3663_), .B(new_n640_), .Y(new_n3664_));
  NOR2  g03279(.A(new_n3664_), .B(new_n646_), .Y(new_n3665_));
  NOR2  g03280(.A(new_n3665_), .B(new_n650_), .Y(new_n3666_));
  NOR2  g03281(.A(new_n3666_), .B(new_n656_), .Y(new_n3667_));
  NOR2  g03282(.A(new_n3667_), .B(new_n660_), .Y(new_n3668_));
  NOR2  g03283(.A(new_n3668_), .B(new_n666_), .Y(new_n3669_));
  NOR2  g03284(.A(new_n3669_), .B(new_n670_), .Y(new_n3670_));
  NOR2  g03285(.A(new_n3670_), .B(new_n676_), .Y(new_n3671_));
  NOR2  g03286(.A(new_n3671_), .B(new_n680_), .Y(new_n3672_));
  NOR2  g03287(.A(new_n3672_), .B(new_n686_), .Y(new_n3673_));
  NOR2  g03288(.A(new_n3673_), .B(new_n690_), .Y(new_n3674_));
  NOR2  g03289(.A(new_n3674_), .B(new_n696_), .Y(new_n3675_));
  NOR2  g03290(.A(new_n3675_), .B(new_n700_), .Y(new_n3676_));
  NOR2  g03291(.A(new_n3676_), .B(new_n706_), .Y(new_n3677_));
  NOR2  g03292(.A(new_n3677_), .B(new_n710_), .Y(new_n3678_));
  NOR2  g03293(.A(new_n3678_), .B(new_n716_), .Y(new_n3679_));
  NOR2  g03294(.A(new_n3679_), .B(new_n720_), .Y(new_n3680_));
  NOR2  g03295(.A(new_n3680_), .B(new_n726_), .Y(new_n3681_));
  NOR2  g03296(.A(new_n3681_), .B(new_n730_), .Y(new_n3682_));
  NOR2  g03297(.A(new_n3682_), .B(new_n736_), .Y(new_n3683_));
  NOR2  g03298(.A(new_n3683_), .B(new_n740_), .Y(new_n3684_));
  NOR2  g03299(.A(new_n3684_), .B(new_n746_), .Y(new_n3685_));
  NOR2  g03300(.A(new_n3685_), .B(new_n750_), .Y(new_n3686_));
  NOR2  g03301(.A(new_n3686_), .B(new_n756_), .Y(new_n3687_));
  NOR2  g03302(.A(new_n3687_), .B(new_n760_), .Y(new_n3688_));
  NOR2  g03303(.A(new_n3688_), .B(new_n766_), .Y(new_n3689_));
  NOR2  g03304(.A(new_n3689_), .B(new_n770_), .Y(new_n3690_));
  NOR2  g03305(.A(new_n3690_), .B(new_n776_), .Y(new_n3691_));
  NOR2  g03306(.A(new_n3691_), .B(new_n780_), .Y(new_n3692_));
  NOR2  g03307(.A(new_n3692_), .B(new_n786_), .Y(new_n3693_));
  NOR2  g03308(.A(new_n3693_), .B(new_n790_), .Y(new_n3694_));
  NOR2  g03309(.A(new_n3694_), .B(new_n796_), .Y(new_n3695_));
  NOR2  g03310(.A(new_n3695_), .B(new_n800_), .Y(new_n3696_));
  NOR2  g03311(.A(new_n3696_), .B(new_n806_), .Y(new_n3697_));
  NOR2  g03312(.A(new_n3697_), .B(new_n1616_), .Y(new_n3698_));
  NOR2  g03313(.A(new_n3698_), .B(new_n1618_), .Y(new_n3699_));
  NOR2  g03314(.A(new_n3699_), .B(new_n1885_), .Y(new_n3700_));
  NOR2  g03315(.A(new_n3700_), .B(new_n820_), .Y(new_n3701_));
  NOR2  g03316(.A(new_n3701_), .B(new_n824_), .Y(new_n3702_));
  NOR2  g03317(.A(new_n3702_), .B(new_n829_), .Y(new_n3703_));
  NOR2  g03318(.A(new_n3703_), .B(new_n833_), .Y(new_n3704_));
  NOR2  g03319(.A(new_n3704_), .B(new_n838_), .Y(new_n3705_));
  NOR2  g03320(.A(new_n3705_), .B(new_n842_), .Y(new_n3706_));
  NOR2  g03321(.A(new_n3706_), .B(new_n847_), .Y(new_n3707_));
  NOR2  g03322(.A(new_n3707_), .B(new_n851_), .Y(new_n3708_));
  NOR2  g03323(.A(new_n3708_), .B(new_n856_), .Y(new_n3709_));
  NOR2  g03324(.A(new_n3709_), .B(new_n860_), .Y(new_n3710_));
  NOR2  g03325(.A(new_n3710_), .B(new_n865_), .Y(new_n3711_));
  NOR2  g03326(.A(new_n3711_), .B(new_n869_), .Y(new_n3712_));
  NOR2  g03327(.A(new_n3712_), .B(new_n874_), .Y(new_n3713_));
  NOR2  g03328(.A(new_n3713_), .B(new_n878_), .Y(new_n3714_));
  NOR2  g03329(.A(new_n3714_), .B(new_n883_), .Y(new_n3715_));
  NAND2 g03330(.A(new_n885_), .B(\req[27] ), .Y(new_n3716_));
  NOR2  g03331(.A(new_n3716_), .B(new_n3715_), .Y(\grant[27] ));
  INV   g03332(.A(new_n895_), .Y(new_n3718_));
  NOR2  g03333(.A(new_n1262_), .B(new_n3718_), .Y(new_n3719_));
  NOR2  g03334(.A(new_n3719_), .B(new_n901_), .Y(new_n3720_));
  NOR2  g03335(.A(new_n3720_), .B(new_n905_), .Y(new_n3721_));
  NOR2  g03336(.A(new_n3721_), .B(new_n910_), .Y(new_n3722_));
  NOR2  g03337(.A(new_n3722_), .B(new_n914_), .Y(new_n3723_));
  NOR2  g03338(.A(new_n3723_), .B(new_n919_), .Y(new_n3724_));
  NOR2  g03339(.A(new_n3724_), .B(new_n923_), .Y(new_n3725_));
  NOR2  g03340(.A(new_n3725_), .B(new_n928_), .Y(new_n3726_));
  NOR2  g03341(.A(new_n3726_), .B(new_n932_), .Y(new_n3727_));
  NOR2  g03342(.A(new_n3727_), .B(new_n937_), .Y(new_n3728_));
  NOR2  g03343(.A(new_n3728_), .B(new_n941_), .Y(new_n3729_));
  NOR2  g03344(.A(new_n3729_), .B(new_n946_), .Y(new_n3730_));
  NOR2  g03345(.A(new_n3730_), .B(new_n950_), .Y(new_n3731_));
  NOR2  g03346(.A(new_n3731_), .B(new_n955_), .Y(new_n3732_));
  NOR2  g03347(.A(new_n3732_), .B(new_n959_), .Y(new_n3733_));
  NOR2  g03348(.A(new_n3733_), .B(new_n964_), .Y(new_n3734_));
  NOR2  g03349(.A(new_n3734_), .B(new_n968_), .Y(new_n3735_));
  NOR2  g03350(.A(new_n3735_), .B(new_n973_), .Y(new_n3736_));
  NOR2  g03351(.A(new_n3736_), .B(new_n977_), .Y(new_n3737_));
  NOR2  g03352(.A(new_n3737_), .B(new_n982_), .Y(new_n3738_));
  NOR2  g03353(.A(new_n3738_), .B(new_n986_), .Y(new_n3739_));
  NOR2  g03354(.A(new_n3739_), .B(new_n991_), .Y(new_n3740_));
  NOR2  g03355(.A(new_n3740_), .B(new_n995_), .Y(new_n3741_));
  NOR2  g03356(.A(new_n3741_), .B(new_n1000_), .Y(new_n3742_));
  NOR2  g03357(.A(new_n3742_), .B(new_n1004_), .Y(new_n3743_));
  NOR2  g03358(.A(new_n3743_), .B(new_n1009_), .Y(new_n3744_));
  NOR2  g03359(.A(new_n3744_), .B(new_n1013_), .Y(new_n3745_));
  NOR2  g03360(.A(new_n3745_), .B(new_n1018_), .Y(new_n3746_));
  NOR2  g03361(.A(new_n3746_), .B(new_n1022_), .Y(new_n3747_));
  NOR2  g03362(.A(new_n3747_), .B(new_n1027_), .Y(new_n3748_));
  NOR2  g03363(.A(new_n3748_), .B(new_n1031_), .Y(new_n3749_));
  NOR2  g03364(.A(new_n3749_), .B(new_n1036_), .Y(new_n3750_));
  NOR2  g03365(.A(new_n3750_), .B(new_n1040_), .Y(new_n3751_));
  NOR2  g03366(.A(new_n3751_), .B(new_n1045_), .Y(new_n3752_));
  NOR2  g03367(.A(new_n3752_), .B(new_n1049_), .Y(new_n3753_));
  NOR2  g03368(.A(new_n3753_), .B(new_n1054_), .Y(new_n3754_));
  NOR2  g03369(.A(new_n3754_), .B(new_n1058_), .Y(new_n3755_));
  NOR2  g03370(.A(new_n3755_), .B(new_n1063_), .Y(new_n3756_));
  NOR2  g03371(.A(new_n3756_), .B(new_n1067_), .Y(new_n3757_));
  NOR2  g03372(.A(new_n3757_), .B(new_n1072_), .Y(new_n3758_));
  NOR2  g03373(.A(new_n3758_), .B(new_n1076_), .Y(new_n3759_));
  NOR2  g03374(.A(new_n3759_), .B(new_n1081_), .Y(new_n3760_));
  NOR2  g03375(.A(new_n3760_), .B(new_n1085_), .Y(new_n3761_));
  NOR2  g03376(.A(new_n3761_), .B(new_n1090_), .Y(new_n3762_));
  NOR2  g03377(.A(new_n3762_), .B(new_n1094_), .Y(new_n3763_));
  NOR2  g03378(.A(new_n3763_), .B(new_n1099_), .Y(new_n3764_));
  NOR2  g03379(.A(new_n3764_), .B(new_n1103_), .Y(new_n3765_));
  NOR2  g03380(.A(new_n3765_), .B(new_n1108_), .Y(new_n3766_));
  NOR2  g03381(.A(new_n3766_), .B(new_n1112_), .Y(new_n3767_));
  NOR2  g03382(.A(new_n3767_), .B(new_n1117_), .Y(new_n3768_));
  NOR2  g03383(.A(new_n3768_), .B(new_n1121_), .Y(new_n3769_));
  NOR2  g03384(.A(new_n3769_), .B(new_n1126_), .Y(new_n3770_));
  NOR2  g03385(.A(new_n3770_), .B(new_n1130_), .Y(new_n3771_));
  NOR2  g03386(.A(new_n3771_), .B(new_n1135_), .Y(new_n3772_));
  NOR2  g03387(.A(new_n3772_), .B(new_n1139_), .Y(new_n3773_));
  NOR2  g03388(.A(new_n3773_), .B(new_n1144_), .Y(new_n3774_));
  NOR2  g03389(.A(new_n3774_), .B(new_n1148_), .Y(new_n3775_));
  NOR2  g03390(.A(new_n3775_), .B(new_n1153_), .Y(new_n3776_));
  NOR2  g03391(.A(new_n3776_), .B(new_n1157_), .Y(new_n3777_));
  NOR2  g03392(.A(new_n3777_), .B(new_n1162_), .Y(new_n3778_));
  NOR2  g03393(.A(new_n3778_), .B(new_n1166_), .Y(new_n3779_));
  NOR2  g03394(.A(new_n3779_), .B(new_n1171_), .Y(new_n3780_));
  NOR2  g03395(.A(new_n3780_), .B(new_n1175_), .Y(new_n3781_));
  NOR2  g03396(.A(new_n3781_), .B(new_n1180_), .Y(new_n3782_));
  NOR2  g03397(.A(new_n3782_), .B(new_n1184_), .Y(new_n3783_));
  NOR2  g03398(.A(new_n3783_), .B(new_n1189_), .Y(new_n3784_));
  NOR2  g03399(.A(new_n3784_), .B(new_n1707_), .Y(new_n3785_));
  NOR2  g03400(.A(new_n3785_), .B(new_n1709_), .Y(new_n3786_));
  NOR2  g03401(.A(new_n3786_), .B(new_n1973_), .Y(new_n3787_));
  NOR2  g03402(.A(new_n3787_), .B(new_n1199_), .Y(new_n3788_));
  NOR2  g03403(.A(new_n3788_), .B(new_n1203_), .Y(new_n3789_));
  NOR2  g03404(.A(new_n3789_), .B(new_n1207_), .Y(new_n3790_));
  NOR2  g03405(.A(new_n3790_), .B(new_n1211_), .Y(new_n3791_));
  NOR2  g03406(.A(new_n3791_), .B(new_n1215_), .Y(new_n3792_));
  NOR2  g03407(.A(new_n3792_), .B(new_n1219_), .Y(new_n3793_));
  NOR2  g03408(.A(new_n3793_), .B(new_n1223_), .Y(new_n3794_));
  NOR2  g03409(.A(new_n3794_), .B(new_n1227_), .Y(new_n3795_));
  NOR2  g03410(.A(new_n3795_), .B(new_n1231_), .Y(new_n3796_));
  NOR2  g03411(.A(new_n3796_), .B(new_n1235_), .Y(new_n3797_));
  NOR2  g03412(.A(new_n3797_), .B(new_n1239_), .Y(new_n3798_));
  NOR2  g03413(.A(new_n3798_), .B(new_n1243_), .Y(new_n3799_));
  NOR2  g03414(.A(new_n3799_), .B(new_n1247_), .Y(new_n3800_));
  NOR2  g03415(.A(new_n3800_), .B(new_n1251_), .Y(new_n3801_));
  NOR2  g03416(.A(new_n3801_), .B(new_n1255_), .Y(new_n3802_));
  NAND2 g03417(.A(new_n1257_), .B(\req[28] ), .Y(new_n3803_));
  NOR2  g03418(.A(new_n3803_), .B(new_n3802_), .Y(\grant[28] ));
  INV   g03419(.A(new_n1266_), .Y(new_n3805_));
  NOR2  g03420(.A(new_n3805_), .B(new_n485_), .Y(new_n3806_));
  NOR2  g03421(.A(new_n3806_), .B(new_n1271_), .Y(new_n3807_));
  NOR2  g03422(.A(new_n3807_), .B(new_n1275_), .Y(new_n3808_));
  NOR2  g03423(.A(new_n3808_), .B(new_n1279_), .Y(new_n3809_));
  NOR2  g03424(.A(new_n3809_), .B(new_n1283_), .Y(new_n3810_));
  NOR2  g03425(.A(new_n3810_), .B(new_n1287_), .Y(new_n3811_));
  NOR2  g03426(.A(new_n3811_), .B(new_n1291_), .Y(new_n3812_));
  NOR2  g03427(.A(new_n3812_), .B(new_n1295_), .Y(new_n3813_));
  NOR2  g03428(.A(new_n3813_), .B(new_n1299_), .Y(new_n3814_));
  NOR2  g03429(.A(new_n3814_), .B(new_n1303_), .Y(new_n3815_));
  NOR2  g03430(.A(new_n3815_), .B(new_n1307_), .Y(new_n3816_));
  NOR2  g03431(.A(new_n3816_), .B(new_n1311_), .Y(new_n3817_));
  NOR2  g03432(.A(new_n3817_), .B(new_n1315_), .Y(new_n3818_));
  NOR2  g03433(.A(new_n3818_), .B(new_n1319_), .Y(new_n3819_));
  NOR2  g03434(.A(new_n3819_), .B(new_n1323_), .Y(new_n3820_));
  NOR2  g03435(.A(new_n3820_), .B(new_n1327_), .Y(new_n3821_));
  NOR2  g03436(.A(new_n3821_), .B(new_n1331_), .Y(new_n3822_));
  NOR2  g03437(.A(new_n3822_), .B(new_n1335_), .Y(new_n3823_));
  NOR2  g03438(.A(new_n3823_), .B(new_n1339_), .Y(new_n3824_));
  NOR2  g03439(.A(new_n3824_), .B(new_n1343_), .Y(new_n3825_));
  NOR2  g03440(.A(new_n3825_), .B(new_n1347_), .Y(new_n3826_));
  NOR2  g03441(.A(new_n3826_), .B(new_n1351_), .Y(new_n3827_));
  NOR2  g03442(.A(new_n3827_), .B(new_n1355_), .Y(new_n3828_));
  NOR2  g03443(.A(new_n3828_), .B(new_n1359_), .Y(new_n3829_));
  NOR2  g03444(.A(new_n3829_), .B(new_n1363_), .Y(new_n3830_));
  NOR2  g03445(.A(new_n3830_), .B(new_n1367_), .Y(new_n3831_));
  NOR2  g03446(.A(new_n3831_), .B(new_n1371_), .Y(new_n3832_));
  NOR2  g03447(.A(new_n3832_), .B(new_n1375_), .Y(new_n3833_));
  NOR2  g03448(.A(new_n3833_), .B(new_n1379_), .Y(new_n3834_));
  NOR2  g03449(.A(new_n3834_), .B(new_n1383_), .Y(new_n3835_));
  NOR2  g03450(.A(new_n3835_), .B(new_n1387_), .Y(new_n3836_));
  NOR2  g03451(.A(new_n3836_), .B(new_n1391_), .Y(new_n3837_));
  NOR2  g03452(.A(new_n3837_), .B(new_n1395_), .Y(new_n3838_));
  NOR2  g03453(.A(new_n3838_), .B(new_n1399_), .Y(new_n3839_));
  NOR2  g03454(.A(new_n3839_), .B(new_n1403_), .Y(new_n3840_));
  NOR2  g03455(.A(new_n3840_), .B(new_n1407_), .Y(new_n3841_));
  NOR2  g03456(.A(new_n3841_), .B(new_n1411_), .Y(new_n3842_));
  NOR2  g03457(.A(new_n3842_), .B(new_n1415_), .Y(new_n3843_));
  NOR2  g03458(.A(new_n3843_), .B(new_n1419_), .Y(new_n3844_));
  NOR2  g03459(.A(new_n3844_), .B(new_n1423_), .Y(new_n3845_));
  NOR2  g03460(.A(new_n3845_), .B(new_n1427_), .Y(new_n3846_));
  NOR2  g03461(.A(new_n3846_), .B(new_n1431_), .Y(new_n3847_));
  NOR2  g03462(.A(new_n3847_), .B(new_n1435_), .Y(new_n3848_));
  NOR2  g03463(.A(new_n3848_), .B(new_n1439_), .Y(new_n3849_));
  NOR2  g03464(.A(new_n3849_), .B(new_n1443_), .Y(new_n3850_));
  NOR2  g03465(.A(new_n3850_), .B(new_n1447_), .Y(new_n3851_));
  NOR2  g03466(.A(new_n3851_), .B(new_n1451_), .Y(new_n3852_));
  NOR2  g03467(.A(new_n3852_), .B(new_n1455_), .Y(new_n3853_));
  NOR2  g03468(.A(new_n3853_), .B(new_n1459_), .Y(new_n3854_));
  NOR2  g03469(.A(new_n3854_), .B(new_n1463_), .Y(new_n3855_));
  NOR2  g03470(.A(new_n3855_), .B(new_n1467_), .Y(new_n3856_));
  NOR2  g03471(.A(new_n3856_), .B(new_n1471_), .Y(new_n3857_));
  NOR2  g03472(.A(new_n3857_), .B(new_n1475_), .Y(new_n3858_));
  NOR2  g03473(.A(new_n3858_), .B(new_n1479_), .Y(new_n3859_));
  NOR2  g03474(.A(new_n3859_), .B(new_n1483_), .Y(new_n3860_));
  NOR2  g03475(.A(new_n3860_), .B(new_n1487_), .Y(new_n3861_));
  NOR2  g03476(.A(new_n3861_), .B(new_n1491_), .Y(new_n3862_));
  NOR2  g03477(.A(new_n3862_), .B(new_n1495_), .Y(new_n3863_));
  NOR2  g03478(.A(new_n3863_), .B(new_n1499_), .Y(new_n3864_));
  NOR2  g03479(.A(new_n3864_), .B(new_n1503_), .Y(new_n3865_));
  NOR2  g03480(.A(new_n3865_), .B(new_n1507_), .Y(new_n3866_));
  NOR2  g03481(.A(new_n3866_), .B(new_n1511_), .Y(new_n3867_));
  NOR2  g03482(.A(new_n3867_), .B(new_n1515_), .Y(new_n3868_));
  NOR2  g03483(.A(new_n3868_), .B(new_n1519_), .Y(new_n3869_));
  NOR2  g03484(.A(new_n3869_), .B(new_n1523_), .Y(new_n3870_));
  NOR2  g03485(.A(new_n3870_), .B(new_n1527_), .Y(new_n3871_));
  NOR2  g03486(.A(new_n3871_), .B(new_n1797_), .Y(new_n3872_));
  NOR2  g03487(.A(new_n3872_), .B(new_n396_), .Y(new_n3873_));
  NOR2  g03488(.A(new_n3873_), .B(new_n400_), .Y(new_n3874_));
  NOR2  g03489(.A(new_n3874_), .B(new_n406_), .Y(new_n3875_));
  NOR2  g03490(.A(new_n3875_), .B(new_n410_), .Y(new_n3876_));
  NOR2  g03491(.A(new_n3876_), .B(new_n416_), .Y(new_n3877_));
  NOR2  g03492(.A(new_n3877_), .B(new_n420_), .Y(new_n3878_));
  NOR2  g03493(.A(new_n3878_), .B(new_n426_), .Y(new_n3879_));
  NOR2  g03494(.A(new_n3879_), .B(new_n430_), .Y(new_n3880_));
  NOR2  g03495(.A(new_n3880_), .B(new_n436_), .Y(new_n3881_));
  NOR2  g03496(.A(new_n3881_), .B(new_n440_), .Y(new_n3882_));
  NOR2  g03497(.A(new_n3882_), .B(new_n446_), .Y(new_n3883_));
  NOR2  g03498(.A(new_n3883_), .B(new_n450_), .Y(new_n3884_));
  NOR2  g03499(.A(new_n3884_), .B(new_n456_), .Y(new_n3885_));
  NOR2  g03500(.A(new_n3885_), .B(new_n460_), .Y(new_n3886_));
  NOR2  g03501(.A(new_n3886_), .B(new_n466_), .Y(new_n3887_));
  NOR2  g03502(.A(new_n3887_), .B(new_n470_), .Y(new_n3888_));
  NOR2  g03503(.A(new_n3888_), .B(new_n476_), .Y(new_n3889_));
  NAND2 g03504(.A(new_n478_), .B(\req[29] ), .Y(new_n3890_));
  NOR2  g03505(.A(new_n3890_), .B(new_n3889_), .Y(\grant[29] ));
  INV   g03506(.A(new_n489_), .Y(new_n3892_));
  NOR2  g03507(.A(new_n900_), .B(new_n3892_), .Y(new_n3893_));
  NOR2  g03508(.A(new_n3893_), .B(new_n496_), .Y(new_n3894_));
  NOR2  g03509(.A(new_n3894_), .B(new_n500_), .Y(new_n3895_));
  NOR2  g03510(.A(new_n3895_), .B(new_n506_), .Y(new_n3896_));
  NOR2  g03511(.A(new_n3896_), .B(new_n510_), .Y(new_n3897_));
  NOR2  g03512(.A(new_n3897_), .B(new_n516_), .Y(new_n3898_));
  NOR2  g03513(.A(new_n3898_), .B(new_n520_), .Y(new_n3899_));
  NOR2  g03514(.A(new_n3899_), .B(new_n526_), .Y(new_n3900_));
  NOR2  g03515(.A(new_n3900_), .B(new_n530_), .Y(new_n3901_));
  NOR2  g03516(.A(new_n3901_), .B(new_n536_), .Y(new_n3902_));
  NOR2  g03517(.A(new_n3902_), .B(new_n540_), .Y(new_n3903_));
  NOR2  g03518(.A(new_n3903_), .B(new_n546_), .Y(new_n3904_));
  NOR2  g03519(.A(new_n3904_), .B(new_n550_), .Y(new_n3905_));
  NOR2  g03520(.A(new_n3905_), .B(new_n556_), .Y(new_n3906_));
  NOR2  g03521(.A(new_n3906_), .B(new_n560_), .Y(new_n3907_));
  NOR2  g03522(.A(new_n3907_), .B(new_n566_), .Y(new_n3908_));
  NOR2  g03523(.A(new_n3908_), .B(new_n570_), .Y(new_n3909_));
  NOR2  g03524(.A(new_n3909_), .B(new_n576_), .Y(new_n3910_));
  NOR2  g03525(.A(new_n3910_), .B(new_n580_), .Y(new_n3911_));
  NOR2  g03526(.A(new_n3911_), .B(new_n586_), .Y(new_n3912_));
  NOR2  g03527(.A(new_n3912_), .B(new_n590_), .Y(new_n3913_));
  NOR2  g03528(.A(new_n3913_), .B(new_n596_), .Y(new_n3914_));
  NOR2  g03529(.A(new_n3914_), .B(new_n600_), .Y(new_n3915_));
  NOR2  g03530(.A(new_n3915_), .B(new_n606_), .Y(new_n3916_));
  NOR2  g03531(.A(new_n3916_), .B(new_n610_), .Y(new_n3917_));
  NOR2  g03532(.A(new_n3917_), .B(new_n616_), .Y(new_n3918_));
  NOR2  g03533(.A(new_n3918_), .B(new_n620_), .Y(new_n3919_));
  NOR2  g03534(.A(new_n3919_), .B(new_n626_), .Y(new_n3920_));
  NOR2  g03535(.A(new_n3920_), .B(new_n630_), .Y(new_n3921_));
  NOR2  g03536(.A(new_n3921_), .B(new_n636_), .Y(new_n3922_));
  NOR2  g03537(.A(new_n3922_), .B(new_n640_), .Y(new_n3923_));
  NOR2  g03538(.A(new_n3923_), .B(new_n646_), .Y(new_n3924_));
  NOR2  g03539(.A(new_n3924_), .B(new_n650_), .Y(new_n3925_));
  NOR2  g03540(.A(new_n3925_), .B(new_n656_), .Y(new_n3926_));
  NOR2  g03541(.A(new_n3926_), .B(new_n660_), .Y(new_n3927_));
  NOR2  g03542(.A(new_n3927_), .B(new_n666_), .Y(new_n3928_));
  NOR2  g03543(.A(new_n3928_), .B(new_n670_), .Y(new_n3929_));
  NOR2  g03544(.A(new_n3929_), .B(new_n676_), .Y(new_n3930_));
  NOR2  g03545(.A(new_n3930_), .B(new_n680_), .Y(new_n3931_));
  NOR2  g03546(.A(new_n3931_), .B(new_n686_), .Y(new_n3932_));
  NOR2  g03547(.A(new_n3932_), .B(new_n690_), .Y(new_n3933_));
  NOR2  g03548(.A(new_n3933_), .B(new_n696_), .Y(new_n3934_));
  NOR2  g03549(.A(new_n3934_), .B(new_n700_), .Y(new_n3935_));
  NOR2  g03550(.A(new_n3935_), .B(new_n706_), .Y(new_n3936_));
  NOR2  g03551(.A(new_n3936_), .B(new_n710_), .Y(new_n3937_));
  NOR2  g03552(.A(new_n3937_), .B(new_n716_), .Y(new_n3938_));
  NOR2  g03553(.A(new_n3938_), .B(new_n720_), .Y(new_n3939_));
  NOR2  g03554(.A(new_n3939_), .B(new_n726_), .Y(new_n3940_));
  NOR2  g03555(.A(new_n3940_), .B(new_n730_), .Y(new_n3941_));
  NOR2  g03556(.A(new_n3941_), .B(new_n736_), .Y(new_n3942_));
  NOR2  g03557(.A(new_n3942_), .B(new_n740_), .Y(new_n3943_));
  NOR2  g03558(.A(new_n3943_), .B(new_n746_), .Y(new_n3944_));
  NOR2  g03559(.A(new_n3944_), .B(new_n750_), .Y(new_n3945_));
  NOR2  g03560(.A(new_n3945_), .B(new_n756_), .Y(new_n3946_));
  NOR2  g03561(.A(new_n3946_), .B(new_n760_), .Y(new_n3947_));
  NOR2  g03562(.A(new_n3947_), .B(new_n766_), .Y(new_n3948_));
  NOR2  g03563(.A(new_n3948_), .B(new_n770_), .Y(new_n3949_));
  NOR2  g03564(.A(new_n3949_), .B(new_n776_), .Y(new_n3950_));
  NOR2  g03565(.A(new_n3950_), .B(new_n780_), .Y(new_n3951_));
  NOR2  g03566(.A(new_n3951_), .B(new_n786_), .Y(new_n3952_));
  NOR2  g03567(.A(new_n3952_), .B(new_n790_), .Y(new_n3953_));
  NOR2  g03568(.A(new_n3953_), .B(new_n796_), .Y(new_n3954_));
  NOR2  g03569(.A(new_n3954_), .B(new_n800_), .Y(new_n3955_));
  NOR2  g03570(.A(new_n3955_), .B(new_n806_), .Y(new_n3956_));
  NOR2  g03571(.A(new_n3956_), .B(new_n1616_), .Y(new_n3957_));
  NOR2  g03572(.A(new_n3957_), .B(new_n1618_), .Y(new_n3958_));
  NOR2  g03573(.A(new_n3958_), .B(new_n1885_), .Y(new_n3959_));
  NOR2  g03574(.A(new_n3959_), .B(new_n820_), .Y(new_n3960_));
  NOR2  g03575(.A(new_n3960_), .B(new_n824_), .Y(new_n3961_));
  NOR2  g03576(.A(new_n3961_), .B(new_n829_), .Y(new_n3962_));
  NOR2  g03577(.A(new_n3962_), .B(new_n833_), .Y(new_n3963_));
  NOR2  g03578(.A(new_n3963_), .B(new_n838_), .Y(new_n3964_));
  NOR2  g03579(.A(new_n3964_), .B(new_n842_), .Y(new_n3965_));
  NOR2  g03580(.A(new_n3965_), .B(new_n847_), .Y(new_n3966_));
  NOR2  g03581(.A(new_n3966_), .B(new_n851_), .Y(new_n3967_));
  NOR2  g03582(.A(new_n3967_), .B(new_n856_), .Y(new_n3968_));
  NOR2  g03583(.A(new_n3968_), .B(new_n860_), .Y(new_n3969_));
  NOR2  g03584(.A(new_n3969_), .B(new_n865_), .Y(new_n3970_));
  NOR2  g03585(.A(new_n3970_), .B(new_n869_), .Y(new_n3971_));
  NOR2  g03586(.A(new_n3971_), .B(new_n874_), .Y(new_n3972_));
  NOR2  g03587(.A(new_n3972_), .B(new_n878_), .Y(new_n3973_));
  NOR2  g03588(.A(new_n3973_), .B(new_n883_), .Y(new_n3974_));
  NOR2  g03589(.A(new_n3974_), .B(new_n887_), .Y(new_n3975_));
  NOR2  g03590(.A(new_n3975_), .B(new_n892_), .Y(new_n3976_));
  NAND2 g03591(.A(new_n894_), .B(\req[30] ), .Y(new_n3977_));
  NOR2  g03592(.A(new_n3977_), .B(new_n3976_), .Y(\grant[30] ));
  INV   g03593(.A(new_n904_), .Y(new_n3979_));
  NOR2  g03594(.A(new_n1270_), .B(new_n3979_), .Y(new_n3980_));
  NOR2  g03595(.A(new_n3980_), .B(new_n910_), .Y(new_n3981_));
  NOR2  g03596(.A(new_n3981_), .B(new_n914_), .Y(new_n3982_));
  NOR2  g03597(.A(new_n3982_), .B(new_n919_), .Y(new_n3983_));
  NOR2  g03598(.A(new_n3983_), .B(new_n923_), .Y(new_n3984_));
  NOR2  g03599(.A(new_n3984_), .B(new_n928_), .Y(new_n3985_));
  NOR2  g03600(.A(new_n3985_), .B(new_n932_), .Y(new_n3986_));
  NOR2  g03601(.A(new_n3986_), .B(new_n937_), .Y(new_n3987_));
  NOR2  g03602(.A(new_n3987_), .B(new_n941_), .Y(new_n3988_));
  NOR2  g03603(.A(new_n3988_), .B(new_n946_), .Y(new_n3989_));
  NOR2  g03604(.A(new_n3989_), .B(new_n950_), .Y(new_n3990_));
  NOR2  g03605(.A(new_n3990_), .B(new_n955_), .Y(new_n3991_));
  NOR2  g03606(.A(new_n3991_), .B(new_n959_), .Y(new_n3992_));
  NOR2  g03607(.A(new_n3992_), .B(new_n964_), .Y(new_n3993_));
  NOR2  g03608(.A(new_n3993_), .B(new_n968_), .Y(new_n3994_));
  NOR2  g03609(.A(new_n3994_), .B(new_n973_), .Y(new_n3995_));
  NOR2  g03610(.A(new_n3995_), .B(new_n977_), .Y(new_n3996_));
  NOR2  g03611(.A(new_n3996_), .B(new_n982_), .Y(new_n3997_));
  NOR2  g03612(.A(new_n3997_), .B(new_n986_), .Y(new_n3998_));
  NOR2  g03613(.A(new_n3998_), .B(new_n991_), .Y(new_n3999_));
  NOR2  g03614(.A(new_n3999_), .B(new_n995_), .Y(new_n4000_));
  NOR2  g03615(.A(new_n4000_), .B(new_n1000_), .Y(new_n4001_));
  NOR2  g03616(.A(new_n4001_), .B(new_n1004_), .Y(new_n4002_));
  NOR2  g03617(.A(new_n4002_), .B(new_n1009_), .Y(new_n4003_));
  NOR2  g03618(.A(new_n4003_), .B(new_n1013_), .Y(new_n4004_));
  NOR2  g03619(.A(new_n4004_), .B(new_n1018_), .Y(new_n4005_));
  NOR2  g03620(.A(new_n4005_), .B(new_n1022_), .Y(new_n4006_));
  NOR2  g03621(.A(new_n4006_), .B(new_n1027_), .Y(new_n4007_));
  NOR2  g03622(.A(new_n4007_), .B(new_n1031_), .Y(new_n4008_));
  NOR2  g03623(.A(new_n4008_), .B(new_n1036_), .Y(new_n4009_));
  NOR2  g03624(.A(new_n4009_), .B(new_n1040_), .Y(new_n4010_));
  NOR2  g03625(.A(new_n4010_), .B(new_n1045_), .Y(new_n4011_));
  NOR2  g03626(.A(new_n4011_), .B(new_n1049_), .Y(new_n4012_));
  NOR2  g03627(.A(new_n4012_), .B(new_n1054_), .Y(new_n4013_));
  NOR2  g03628(.A(new_n4013_), .B(new_n1058_), .Y(new_n4014_));
  NOR2  g03629(.A(new_n4014_), .B(new_n1063_), .Y(new_n4015_));
  NOR2  g03630(.A(new_n4015_), .B(new_n1067_), .Y(new_n4016_));
  NOR2  g03631(.A(new_n4016_), .B(new_n1072_), .Y(new_n4017_));
  NOR2  g03632(.A(new_n4017_), .B(new_n1076_), .Y(new_n4018_));
  NOR2  g03633(.A(new_n4018_), .B(new_n1081_), .Y(new_n4019_));
  NOR2  g03634(.A(new_n4019_), .B(new_n1085_), .Y(new_n4020_));
  NOR2  g03635(.A(new_n4020_), .B(new_n1090_), .Y(new_n4021_));
  NOR2  g03636(.A(new_n4021_), .B(new_n1094_), .Y(new_n4022_));
  NOR2  g03637(.A(new_n4022_), .B(new_n1099_), .Y(new_n4023_));
  NOR2  g03638(.A(new_n4023_), .B(new_n1103_), .Y(new_n4024_));
  NOR2  g03639(.A(new_n4024_), .B(new_n1108_), .Y(new_n4025_));
  NOR2  g03640(.A(new_n4025_), .B(new_n1112_), .Y(new_n4026_));
  NOR2  g03641(.A(new_n4026_), .B(new_n1117_), .Y(new_n4027_));
  NOR2  g03642(.A(new_n4027_), .B(new_n1121_), .Y(new_n4028_));
  NOR2  g03643(.A(new_n4028_), .B(new_n1126_), .Y(new_n4029_));
  NOR2  g03644(.A(new_n4029_), .B(new_n1130_), .Y(new_n4030_));
  NOR2  g03645(.A(new_n4030_), .B(new_n1135_), .Y(new_n4031_));
  NOR2  g03646(.A(new_n4031_), .B(new_n1139_), .Y(new_n4032_));
  NOR2  g03647(.A(new_n4032_), .B(new_n1144_), .Y(new_n4033_));
  NOR2  g03648(.A(new_n4033_), .B(new_n1148_), .Y(new_n4034_));
  NOR2  g03649(.A(new_n4034_), .B(new_n1153_), .Y(new_n4035_));
  NOR2  g03650(.A(new_n4035_), .B(new_n1157_), .Y(new_n4036_));
  NOR2  g03651(.A(new_n4036_), .B(new_n1162_), .Y(new_n4037_));
  NOR2  g03652(.A(new_n4037_), .B(new_n1166_), .Y(new_n4038_));
  NOR2  g03653(.A(new_n4038_), .B(new_n1171_), .Y(new_n4039_));
  NOR2  g03654(.A(new_n4039_), .B(new_n1175_), .Y(new_n4040_));
  NOR2  g03655(.A(new_n4040_), .B(new_n1180_), .Y(new_n4041_));
  NOR2  g03656(.A(new_n4041_), .B(new_n1184_), .Y(new_n4042_));
  NOR2  g03657(.A(new_n4042_), .B(new_n1189_), .Y(new_n4043_));
  NOR2  g03658(.A(new_n4043_), .B(new_n1707_), .Y(new_n4044_));
  NOR2  g03659(.A(new_n4044_), .B(new_n1709_), .Y(new_n4045_));
  NOR2  g03660(.A(new_n4045_), .B(new_n1973_), .Y(new_n4046_));
  NOR2  g03661(.A(new_n4046_), .B(new_n1199_), .Y(new_n4047_));
  NOR2  g03662(.A(new_n4047_), .B(new_n1203_), .Y(new_n4048_));
  NOR2  g03663(.A(new_n4048_), .B(new_n1207_), .Y(new_n4049_));
  NOR2  g03664(.A(new_n4049_), .B(new_n1211_), .Y(new_n4050_));
  NOR2  g03665(.A(new_n4050_), .B(new_n1215_), .Y(new_n4051_));
  NOR2  g03666(.A(new_n4051_), .B(new_n1219_), .Y(new_n4052_));
  NOR2  g03667(.A(new_n4052_), .B(new_n1223_), .Y(new_n4053_));
  NOR2  g03668(.A(new_n4053_), .B(new_n1227_), .Y(new_n4054_));
  NOR2  g03669(.A(new_n4054_), .B(new_n1231_), .Y(new_n4055_));
  NOR2  g03670(.A(new_n4055_), .B(new_n1235_), .Y(new_n4056_));
  NOR2  g03671(.A(new_n4056_), .B(new_n1239_), .Y(new_n4057_));
  NOR2  g03672(.A(new_n4057_), .B(new_n1243_), .Y(new_n4058_));
  NOR2  g03673(.A(new_n4058_), .B(new_n1247_), .Y(new_n4059_));
  NOR2  g03674(.A(new_n4059_), .B(new_n1251_), .Y(new_n4060_));
  NOR2  g03675(.A(new_n4060_), .B(new_n1255_), .Y(new_n4061_));
  NOR2  g03676(.A(new_n4061_), .B(new_n1259_), .Y(new_n4062_));
  NOR2  g03677(.A(new_n4062_), .B(new_n1263_), .Y(new_n4063_));
  NAND2 g03678(.A(new_n1265_), .B(\req[31] ), .Y(new_n4064_));
  NOR2  g03679(.A(new_n4064_), .B(new_n4063_), .Y(\grant[31] ));
  INV   g03680(.A(new_n1274_), .Y(new_n4066_));
  NOR2  g03681(.A(new_n4066_), .B(new_n495_), .Y(new_n4067_));
  NOR2  g03682(.A(new_n4067_), .B(new_n1279_), .Y(new_n4068_));
  NOR2  g03683(.A(new_n4068_), .B(new_n1283_), .Y(new_n4069_));
  NOR2  g03684(.A(new_n4069_), .B(new_n1287_), .Y(new_n4070_));
  NOR2  g03685(.A(new_n4070_), .B(new_n1291_), .Y(new_n4071_));
  NOR2  g03686(.A(new_n4071_), .B(new_n1295_), .Y(new_n4072_));
  NOR2  g03687(.A(new_n4072_), .B(new_n1299_), .Y(new_n4073_));
  NOR2  g03688(.A(new_n4073_), .B(new_n1303_), .Y(new_n4074_));
  NOR2  g03689(.A(new_n4074_), .B(new_n1307_), .Y(new_n4075_));
  NOR2  g03690(.A(new_n4075_), .B(new_n1311_), .Y(new_n4076_));
  NOR2  g03691(.A(new_n4076_), .B(new_n1315_), .Y(new_n4077_));
  NOR2  g03692(.A(new_n4077_), .B(new_n1319_), .Y(new_n4078_));
  NOR2  g03693(.A(new_n4078_), .B(new_n1323_), .Y(new_n4079_));
  NOR2  g03694(.A(new_n4079_), .B(new_n1327_), .Y(new_n4080_));
  NOR2  g03695(.A(new_n4080_), .B(new_n1331_), .Y(new_n4081_));
  NOR2  g03696(.A(new_n4081_), .B(new_n1335_), .Y(new_n4082_));
  NOR2  g03697(.A(new_n4082_), .B(new_n1339_), .Y(new_n4083_));
  NOR2  g03698(.A(new_n4083_), .B(new_n1343_), .Y(new_n4084_));
  NOR2  g03699(.A(new_n4084_), .B(new_n1347_), .Y(new_n4085_));
  NOR2  g03700(.A(new_n4085_), .B(new_n1351_), .Y(new_n4086_));
  NOR2  g03701(.A(new_n4086_), .B(new_n1355_), .Y(new_n4087_));
  NOR2  g03702(.A(new_n4087_), .B(new_n1359_), .Y(new_n4088_));
  NOR2  g03703(.A(new_n4088_), .B(new_n1363_), .Y(new_n4089_));
  NOR2  g03704(.A(new_n4089_), .B(new_n1367_), .Y(new_n4090_));
  NOR2  g03705(.A(new_n4090_), .B(new_n1371_), .Y(new_n4091_));
  NOR2  g03706(.A(new_n4091_), .B(new_n1375_), .Y(new_n4092_));
  NOR2  g03707(.A(new_n4092_), .B(new_n1379_), .Y(new_n4093_));
  NOR2  g03708(.A(new_n4093_), .B(new_n1383_), .Y(new_n4094_));
  NOR2  g03709(.A(new_n4094_), .B(new_n1387_), .Y(new_n4095_));
  NOR2  g03710(.A(new_n4095_), .B(new_n1391_), .Y(new_n4096_));
  NOR2  g03711(.A(new_n4096_), .B(new_n1395_), .Y(new_n4097_));
  NOR2  g03712(.A(new_n4097_), .B(new_n1399_), .Y(new_n4098_));
  NOR2  g03713(.A(new_n4098_), .B(new_n1403_), .Y(new_n4099_));
  NOR2  g03714(.A(new_n4099_), .B(new_n1407_), .Y(new_n4100_));
  NOR2  g03715(.A(new_n4100_), .B(new_n1411_), .Y(new_n4101_));
  NOR2  g03716(.A(new_n4101_), .B(new_n1415_), .Y(new_n4102_));
  NOR2  g03717(.A(new_n4102_), .B(new_n1419_), .Y(new_n4103_));
  NOR2  g03718(.A(new_n4103_), .B(new_n1423_), .Y(new_n4104_));
  NOR2  g03719(.A(new_n4104_), .B(new_n1427_), .Y(new_n4105_));
  NOR2  g03720(.A(new_n4105_), .B(new_n1431_), .Y(new_n4106_));
  NOR2  g03721(.A(new_n4106_), .B(new_n1435_), .Y(new_n4107_));
  NOR2  g03722(.A(new_n4107_), .B(new_n1439_), .Y(new_n4108_));
  NOR2  g03723(.A(new_n4108_), .B(new_n1443_), .Y(new_n4109_));
  NOR2  g03724(.A(new_n4109_), .B(new_n1447_), .Y(new_n4110_));
  NOR2  g03725(.A(new_n4110_), .B(new_n1451_), .Y(new_n4111_));
  NOR2  g03726(.A(new_n4111_), .B(new_n1455_), .Y(new_n4112_));
  NOR2  g03727(.A(new_n4112_), .B(new_n1459_), .Y(new_n4113_));
  NOR2  g03728(.A(new_n4113_), .B(new_n1463_), .Y(new_n4114_));
  NOR2  g03729(.A(new_n4114_), .B(new_n1467_), .Y(new_n4115_));
  NOR2  g03730(.A(new_n4115_), .B(new_n1471_), .Y(new_n4116_));
  NOR2  g03731(.A(new_n4116_), .B(new_n1475_), .Y(new_n4117_));
  NOR2  g03732(.A(new_n4117_), .B(new_n1479_), .Y(new_n4118_));
  NOR2  g03733(.A(new_n4118_), .B(new_n1483_), .Y(new_n4119_));
  NOR2  g03734(.A(new_n4119_), .B(new_n1487_), .Y(new_n4120_));
  NOR2  g03735(.A(new_n4120_), .B(new_n1491_), .Y(new_n4121_));
  NOR2  g03736(.A(new_n4121_), .B(new_n1495_), .Y(new_n4122_));
  NOR2  g03737(.A(new_n4122_), .B(new_n1499_), .Y(new_n4123_));
  NOR2  g03738(.A(new_n4123_), .B(new_n1503_), .Y(new_n4124_));
  NOR2  g03739(.A(new_n4124_), .B(new_n1507_), .Y(new_n4125_));
  NOR2  g03740(.A(new_n4125_), .B(new_n1511_), .Y(new_n4126_));
  NOR2  g03741(.A(new_n4126_), .B(new_n1515_), .Y(new_n4127_));
  NOR2  g03742(.A(new_n4127_), .B(new_n1519_), .Y(new_n4128_));
  NOR2  g03743(.A(new_n4128_), .B(new_n1523_), .Y(new_n4129_));
  NOR2  g03744(.A(new_n4129_), .B(new_n1527_), .Y(new_n4130_));
  NOR2  g03745(.A(new_n4130_), .B(new_n1797_), .Y(new_n4131_));
  NOR2  g03746(.A(new_n4131_), .B(new_n396_), .Y(new_n4132_));
  NOR2  g03747(.A(new_n4132_), .B(new_n400_), .Y(new_n4133_));
  NOR2  g03748(.A(new_n4133_), .B(new_n406_), .Y(new_n4134_));
  NOR2  g03749(.A(new_n4134_), .B(new_n410_), .Y(new_n4135_));
  NOR2  g03750(.A(new_n4135_), .B(new_n416_), .Y(new_n4136_));
  NOR2  g03751(.A(new_n4136_), .B(new_n420_), .Y(new_n4137_));
  NOR2  g03752(.A(new_n4137_), .B(new_n426_), .Y(new_n4138_));
  NOR2  g03753(.A(new_n4138_), .B(new_n430_), .Y(new_n4139_));
  NOR2  g03754(.A(new_n4139_), .B(new_n436_), .Y(new_n4140_));
  NOR2  g03755(.A(new_n4140_), .B(new_n440_), .Y(new_n4141_));
  NOR2  g03756(.A(new_n4141_), .B(new_n446_), .Y(new_n4142_));
  NOR2  g03757(.A(new_n4142_), .B(new_n450_), .Y(new_n4143_));
  NOR2  g03758(.A(new_n4143_), .B(new_n456_), .Y(new_n4144_));
  NOR2  g03759(.A(new_n4144_), .B(new_n460_), .Y(new_n4145_));
  NOR2  g03760(.A(new_n4145_), .B(new_n466_), .Y(new_n4146_));
  NOR2  g03761(.A(new_n4146_), .B(new_n470_), .Y(new_n4147_));
  NOR2  g03762(.A(new_n4147_), .B(new_n476_), .Y(new_n4148_));
  NOR2  g03763(.A(new_n4148_), .B(new_n480_), .Y(new_n4149_));
  NOR2  g03764(.A(new_n4149_), .B(new_n486_), .Y(new_n4150_));
  NAND2 g03765(.A(new_n488_), .B(\req[32] ), .Y(new_n4151_));
  NOR2  g03766(.A(new_n4151_), .B(new_n4150_), .Y(\grant[32] ));
  INV   g03767(.A(new_n499_), .Y(new_n4153_));
  NOR2  g03768(.A(new_n909_), .B(new_n4153_), .Y(new_n4154_));
  NOR2  g03769(.A(new_n4154_), .B(new_n506_), .Y(new_n4155_));
  NOR2  g03770(.A(new_n4155_), .B(new_n510_), .Y(new_n4156_));
  NOR2  g03771(.A(new_n4156_), .B(new_n516_), .Y(new_n4157_));
  NOR2  g03772(.A(new_n4157_), .B(new_n520_), .Y(new_n4158_));
  NOR2  g03773(.A(new_n4158_), .B(new_n526_), .Y(new_n4159_));
  NOR2  g03774(.A(new_n4159_), .B(new_n530_), .Y(new_n4160_));
  NOR2  g03775(.A(new_n4160_), .B(new_n536_), .Y(new_n4161_));
  NOR2  g03776(.A(new_n4161_), .B(new_n540_), .Y(new_n4162_));
  NOR2  g03777(.A(new_n4162_), .B(new_n546_), .Y(new_n4163_));
  NOR2  g03778(.A(new_n4163_), .B(new_n550_), .Y(new_n4164_));
  NOR2  g03779(.A(new_n4164_), .B(new_n556_), .Y(new_n4165_));
  NOR2  g03780(.A(new_n4165_), .B(new_n560_), .Y(new_n4166_));
  NOR2  g03781(.A(new_n4166_), .B(new_n566_), .Y(new_n4167_));
  NOR2  g03782(.A(new_n4167_), .B(new_n570_), .Y(new_n4168_));
  NOR2  g03783(.A(new_n4168_), .B(new_n576_), .Y(new_n4169_));
  NOR2  g03784(.A(new_n4169_), .B(new_n580_), .Y(new_n4170_));
  NOR2  g03785(.A(new_n4170_), .B(new_n586_), .Y(new_n4171_));
  NOR2  g03786(.A(new_n4171_), .B(new_n590_), .Y(new_n4172_));
  NOR2  g03787(.A(new_n4172_), .B(new_n596_), .Y(new_n4173_));
  NOR2  g03788(.A(new_n4173_), .B(new_n600_), .Y(new_n4174_));
  NOR2  g03789(.A(new_n4174_), .B(new_n606_), .Y(new_n4175_));
  NOR2  g03790(.A(new_n4175_), .B(new_n610_), .Y(new_n4176_));
  NOR2  g03791(.A(new_n4176_), .B(new_n616_), .Y(new_n4177_));
  NOR2  g03792(.A(new_n4177_), .B(new_n620_), .Y(new_n4178_));
  NOR2  g03793(.A(new_n4178_), .B(new_n626_), .Y(new_n4179_));
  NOR2  g03794(.A(new_n4179_), .B(new_n630_), .Y(new_n4180_));
  NOR2  g03795(.A(new_n4180_), .B(new_n636_), .Y(new_n4181_));
  NOR2  g03796(.A(new_n4181_), .B(new_n640_), .Y(new_n4182_));
  NOR2  g03797(.A(new_n4182_), .B(new_n646_), .Y(new_n4183_));
  NOR2  g03798(.A(new_n4183_), .B(new_n650_), .Y(new_n4184_));
  NOR2  g03799(.A(new_n4184_), .B(new_n656_), .Y(new_n4185_));
  NOR2  g03800(.A(new_n4185_), .B(new_n660_), .Y(new_n4186_));
  NOR2  g03801(.A(new_n4186_), .B(new_n666_), .Y(new_n4187_));
  NOR2  g03802(.A(new_n4187_), .B(new_n670_), .Y(new_n4188_));
  NOR2  g03803(.A(new_n4188_), .B(new_n676_), .Y(new_n4189_));
  NOR2  g03804(.A(new_n4189_), .B(new_n680_), .Y(new_n4190_));
  NOR2  g03805(.A(new_n4190_), .B(new_n686_), .Y(new_n4191_));
  NOR2  g03806(.A(new_n4191_), .B(new_n690_), .Y(new_n4192_));
  NOR2  g03807(.A(new_n4192_), .B(new_n696_), .Y(new_n4193_));
  NOR2  g03808(.A(new_n4193_), .B(new_n700_), .Y(new_n4194_));
  NOR2  g03809(.A(new_n4194_), .B(new_n706_), .Y(new_n4195_));
  NOR2  g03810(.A(new_n4195_), .B(new_n710_), .Y(new_n4196_));
  NOR2  g03811(.A(new_n4196_), .B(new_n716_), .Y(new_n4197_));
  NOR2  g03812(.A(new_n4197_), .B(new_n720_), .Y(new_n4198_));
  NOR2  g03813(.A(new_n4198_), .B(new_n726_), .Y(new_n4199_));
  NOR2  g03814(.A(new_n4199_), .B(new_n730_), .Y(new_n4200_));
  NOR2  g03815(.A(new_n4200_), .B(new_n736_), .Y(new_n4201_));
  NOR2  g03816(.A(new_n4201_), .B(new_n740_), .Y(new_n4202_));
  NOR2  g03817(.A(new_n4202_), .B(new_n746_), .Y(new_n4203_));
  NOR2  g03818(.A(new_n4203_), .B(new_n750_), .Y(new_n4204_));
  NOR2  g03819(.A(new_n4204_), .B(new_n756_), .Y(new_n4205_));
  NOR2  g03820(.A(new_n4205_), .B(new_n760_), .Y(new_n4206_));
  NOR2  g03821(.A(new_n4206_), .B(new_n766_), .Y(new_n4207_));
  NOR2  g03822(.A(new_n4207_), .B(new_n770_), .Y(new_n4208_));
  NOR2  g03823(.A(new_n4208_), .B(new_n776_), .Y(new_n4209_));
  NOR2  g03824(.A(new_n4209_), .B(new_n780_), .Y(new_n4210_));
  NOR2  g03825(.A(new_n4210_), .B(new_n786_), .Y(new_n4211_));
  NOR2  g03826(.A(new_n4211_), .B(new_n790_), .Y(new_n4212_));
  NOR2  g03827(.A(new_n4212_), .B(new_n796_), .Y(new_n4213_));
  NOR2  g03828(.A(new_n4213_), .B(new_n800_), .Y(new_n4214_));
  NOR2  g03829(.A(new_n4214_), .B(new_n806_), .Y(new_n4215_));
  NOR2  g03830(.A(new_n4215_), .B(new_n1616_), .Y(new_n4216_));
  NOR2  g03831(.A(new_n4216_), .B(new_n1618_), .Y(new_n4217_));
  NOR2  g03832(.A(new_n4217_), .B(new_n1885_), .Y(new_n4218_));
  NOR2  g03833(.A(new_n4218_), .B(new_n820_), .Y(new_n4219_));
  NOR2  g03834(.A(new_n4219_), .B(new_n824_), .Y(new_n4220_));
  NOR2  g03835(.A(new_n4220_), .B(new_n829_), .Y(new_n4221_));
  NOR2  g03836(.A(new_n4221_), .B(new_n833_), .Y(new_n4222_));
  NOR2  g03837(.A(new_n4222_), .B(new_n838_), .Y(new_n4223_));
  NOR2  g03838(.A(new_n4223_), .B(new_n842_), .Y(new_n4224_));
  NOR2  g03839(.A(new_n4224_), .B(new_n847_), .Y(new_n4225_));
  NOR2  g03840(.A(new_n4225_), .B(new_n851_), .Y(new_n4226_));
  NOR2  g03841(.A(new_n4226_), .B(new_n856_), .Y(new_n4227_));
  NOR2  g03842(.A(new_n4227_), .B(new_n860_), .Y(new_n4228_));
  NOR2  g03843(.A(new_n4228_), .B(new_n865_), .Y(new_n4229_));
  NOR2  g03844(.A(new_n4229_), .B(new_n869_), .Y(new_n4230_));
  NOR2  g03845(.A(new_n4230_), .B(new_n874_), .Y(new_n4231_));
  NOR2  g03846(.A(new_n4231_), .B(new_n878_), .Y(new_n4232_));
  NOR2  g03847(.A(new_n4232_), .B(new_n883_), .Y(new_n4233_));
  NOR2  g03848(.A(new_n4233_), .B(new_n887_), .Y(new_n4234_));
  NOR2  g03849(.A(new_n4234_), .B(new_n892_), .Y(new_n4235_));
  NOR2  g03850(.A(new_n4235_), .B(new_n896_), .Y(new_n4236_));
  NOR2  g03851(.A(new_n4236_), .B(new_n901_), .Y(new_n4237_));
  NAND2 g03852(.A(new_n903_), .B(\req[33] ), .Y(new_n4238_));
  NOR2  g03853(.A(new_n4238_), .B(new_n4237_), .Y(\grant[33] ));
  INV   g03854(.A(new_n913_), .Y(new_n4240_));
  NOR2  g03855(.A(new_n1278_), .B(new_n4240_), .Y(new_n4241_));
  NOR2  g03856(.A(new_n4241_), .B(new_n919_), .Y(new_n4242_));
  NOR2  g03857(.A(new_n4242_), .B(new_n923_), .Y(new_n4243_));
  NOR2  g03858(.A(new_n4243_), .B(new_n928_), .Y(new_n4244_));
  NOR2  g03859(.A(new_n4244_), .B(new_n932_), .Y(new_n4245_));
  NOR2  g03860(.A(new_n4245_), .B(new_n937_), .Y(new_n4246_));
  NOR2  g03861(.A(new_n4246_), .B(new_n941_), .Y(new_n4247_));
  NOR2  g03862(.A(new_n4247_), .B(new_n946_), .Y(new_n4248_));
  NOR2  g03863(.A(new_n4248_), .B(new_n950_), .Y(new_n4249_));
  NOR2  g03864(.A(new_n4249_), .B(new_n955_), .Y(new_n4250_));
  NOR2  g03865(.A(new_n4250_), .B(new_n959_), .Y(new_n4251_));
  NOR2  g03866(.A(new_n4251_), .B(new_n964_), .Y(new_n4252_));
  NOR2  g03867(.A(new_n4252_), .B(new_n968_), .Y(new_n4253_));
  NOR2  g03868(.A(new_n4253_), .B(new_n973_), .Y(new_n4254_));
  NOR2  g03869(.A(new_n4254_), .B(new_n977_), .Y(new_n4255_));
  NOR2  g03870(.A(new_n4255_), .B(new_n982_), .Y(new_n4256_));
  NOR2  g03871(.A(new_n4256_), .B(new_n986_), .Y(new_n4257_));
  NOR2  g03872(.A(new_n4257_), .B(new_n991_), .Y(new_n4258_));
  NOR2  g03873(.A(new_n4258_), .B(new_n995_), .Y(new_n4259_));
  NOR2  g03874(.A(new_n4259_), .B(new_n1000_), .Y(new_n4260_));
  NOR2  g03875(.A(new_n4260_), .B(new_n1004_), .Y(new_n4261_));
  NOR2  g03876(.A(new_n4261_), .B(new_n1009_), .Y(new_n4262_));
  NOR2  g03877(.A(new_n4262_), .B(new_n1013_), .Y(new_n4263_));
  NOR2  g03878(.A(new_n4263_), .B(new_n1018_), .Y(new_n4264_));
  NOR2  g03879(.A(new_n4264_), .B(new_n1022_), .Y(new_n4265_));
  NOR2  g03880(.A(new_n4265_), .B(new_n1027_), .Y(new_n4266_));
  NOR2  g03881(.A(new_n4266_), .B(new_n1031_), .Y(new_n4267_));
  NOR2  g03882(.A(new_n4267_), .B(new_n1036_), .Y(new_n4268_));
  NOR2  g03883(.A(new_n4268_), .B(new_n1040_), .Y(new_n4269_));
  NOR2  g03884(.A(new_n4269_), .B(new_n1045_), .Y(new_n4270_));
  NOR2  g03885(.A(new_n4270_), .B(new_n1049_), .Y(new_n4271_));
  NOR2  g03886(.A(new_n4271_), .B(new_n1054_), .Y(new_n4272_));
  NOR2  g03887(.A(new_n4272_), .B(new_n1058_), .Y(new_n4273_));
  NOR2  g03888(.A(new_n4273_), .B(new_n1063_), .Y(new_n4274_));
  NOR2  g03889(.A(new_n4274_), .B(new_n1067_), .Y(new_n4275_));
  NOR2  g03890(.A(new_n4275_), .B(new_n1072_), .Y(new_n4276_));
  NOR2  g03891(.A(new_n4276_), .B(new_n1076_), .Y(new_n4277_));
  NOR2  g03892(.A(new_n4277_), .B(new_n1081_), .Y(new_n4278_));
  NOR2  g03893(.A(new_n4278_), .B(new_n1085_), .Y(new_n4279_));
  NOR2  g03894(.A(new_n4279_), .B(new_n1090_), .Y(new_n4280_));
  NOR2  g03895(.A(new_n4280_), .B(new_n1094_), .Y(new_n4281_));
  NOR2  g03896(.A(new_n4281_), .B(new_n1099_), .Y(new_n4282_));
  NOR2  g03897(.A(new_n4282_), .B(new_n1103_), .Y(new_n4283_));
  NOR2  g03898(.A(new_n4283_), .B(new_n1108_), .Y(new_n4284_));
  NOR2  g03899(.A(new_n4284_), .B(new_n1112_), .Y(new_n4285_));
  NOR2  g03900(.A(new_n4285_), .B(new_n1117_), .Y(new_n4286_));
  NOR2  g03901(.A(new_n4286_), .B(new_n1121_), .Y(new_n4287_));
  NOR2  g03902(.A(new_n4287_), .B(new_n1126_), .Y(new_n4288_));
  NOR2  g03903(.A(new_n4288_), .B(new_n1130_), .Y(new_n4289_));
  NOR2  g03904(.A(new_n4289_), .B(new_n1135_), .Y(new_n4290_));
  NOR2  g03905(.A(new_n4290_), .B(new_n1139_), .Y(new_n4291_));
  NOR2  g03906(.A(new_n4291_), .B(new_n1144_), .Y(new_n4292_));
  NOR2  g03907(.A(new_n4292_), .B(new_n1148_), .Y(new_n4293_));
  NOR2  g03908(.A(new_n4293_), .B(new_n1153_), .Y(new_n4294_));
  NOR2  g03909(.A(new_n4294_), .B(new_n1157_), .Y(new_n4295_));
  NOR2  g03910(.A(new_n4295_), .B(new_n1162_), .Y(new_n4296_));
  NOR2  g03911(.A(new_n4296_), .B(new_n1166_), .Y(new_n4297_));
  NOR2  g03912(.A(new_n4297_), .B(new_n1171_), .Y(new_n4298_));
  NOR2  g03913(.A(new_n4298_), .B(new_n1175_), .Y(new_n4299_));
  NOR2  g03914(.A(new_n4299_), .B(new_n1180_), .Y(new_n4300_));
  NOR2  g03915(.A(new_n4300_), .B(new_n1184_), .Y(new_n4301_));
  NOR2  g03916(.A(new_n4301_), .B(new_n1189_), .Y(new_n4302_));
  NOR2  g03917(.A(new_n4302_), .B(new_n1707_), .Y(new_n4303_));
  NOR2  g03918(.A(new_n4303_), .B(new_n1709_), .Y(new_n4304_));
  NOR2  g03919(.A(new_n4304_), .B(new_n1973_), .Y(new_n4305_));
  NOR2  g03920(.A(new_n4305_), .B(new_n1199_), .Y(new_n4306_));
  NOR2  g03921(.A(new_n4306_), .B(new_n1203_), .Y(new_n4307_));
  NOR2  g03922(.A(new_n4307_), .B(new_n1207_), .Y(new_n4308_));
  NOR2  g03923(.A(new_n4308_), .B(new_n1211_), .Y(new_n4309_));
  NOR2  g03924(.A(new_n4309_), .B(new_n1215_), .Y(new_n4310_));
  NOR2  g03925(.A(new_n4310_), .B(new_n1219_), .Y(new_n4311_));
  NOR2  g03926(.A(new_n4311_), .B(new_n1223_), .Y(new_n4312_));
  NOR2  g03927(.A(new_n4312_), .B(new_n1227_), .Y(new_n4313_));
  NOR2  g03928(.A(new_n4313_), .B(new_n1231_), .Y(new_n4314_));
  NOR2  g03929(.A(new_n4314_), .B(new_n1235_), .Y(new_n4315_));
  NOR2  g03930(.A(new_n4315_), .B(new_n1239_), .Y(new_n4316_));
  NOR2  g03931(.A(new_n4316_), .B(new_n1243_), .Y(new_n4317_));
  NOR2  g03932(.A(new_n4317_), .B(new_n1247_), .Y(new_n4318_));
  NOR2  g03933(.A(new_n4318_), .B(new_n1251_), .Y(new_n4319_));
  NOR2  g03934(.A(new_n4319_), .B(new_n1255_), .Y(new_n4320_));
  NOR2  g03935(.A(new_n4320_), .B(new_n1259_), .Y(new_n4321_));
  NOR2  g03936(.A(new_n4321_), .B(new_n1263_), .Y(new_n4322_));
  NOR2  g03937(.A(new_n4322_), .B(new_n1267_), .Y(new_n4323_));
  NOR2  g03938(.A(new_n4323_), .B(new_n1271_), .Y(new_n4324_));
  NAND2 g03939(.A(new_n1273_), .B(\req[34] ), .Y(new_n4325_));
  NOR2  g03940(.A(new_n4325_), .B(new_n4324_), .Y(\grant[34] ));
  INV   g03941(.A(new_n1282_), .Y(new_n4327_));
  NOR2  g03942(.A(new_n4327_), .B(new_n505_), .Y(new_n4328_));
  NOR2  g03943(.A(new_n4328_), .B(new_n1287_), .Y(new_n4329_));
  NOR2  g03944(.A(new_n4329_), .B(new_n1291_), .Y(new_n4330_));
  NOR2  g03945(.A(new_n4330_), .B(new_n1295_), .Y(new_n4331_));
  NOR2  g03946(.A(new_n4331_), .B(new_n1299_), .Y(new_n4332_));
  NOR2  g03947(.A(new_n4332_), .B(new_n1303_), .Y(new_n4333_));
  NOR2  g03948(.A(new_n4333_), .B(new_n1307_), .Y(new_n4334_));
  NOR2  g03949(.A(new_n4334_), .B(new_n1311_), .Y(new_n4335_));
  NOR2  g03950(.A(new_n4335_), .B(new_n1315_), .Y(new_n4336_));
  NOR2  g03951(.A(new_n4336_), .B(new_n1319_), .Y(new_n4337_));
  NOR2  g03952(.A(new_n4337_), .B(new_n1323_), .Y(new_n4338_));
  NOR2  g03953(.A(new_n4338_), .B(new_n1327_), .Y(new_n4339_));
  NOR2  g03954(.A(new_n4339_), .B(new_n1331_), .Y(new_n4340_));
  NOR2  g03955(.A(new_n4340_), .B(new_n1335_), .Y(new_n4341_));
  NOR2  g03956(.A(new_n4341_), .B(new_n1339_), .Y(new_n4342_));
  NOR2  g03957(.A(new_n4342_), .B(new_n1343_), .Y(new_n4343_));
  NOR2  g03958(.A(new_n4343_), .B(new_n1347_), .Y(new_n4344_));
  NOR2  g03959(.A(new_n4344_), .B(new_n1351_), .Y(new_n4345_));
  NOR2  g03960(.A(new_n4345_), .B(new_n1355_), .Y(new_n4346_));
  NOR2  g03961(.A(new_n4346_), .B(new_n1359_), .Y(new_n4347_));
  NOR2  g03962(.A(new_n4347_), .B(new_n1363_), .Y(new_n4348_));
  NOR2  g03963(.A(new_n4348_), .B(new_n1367_), .Y(new_n4349_));
  NOR2  g03964(.A(new_n4349_), .B(new_n1371_), .Y(new_n4350_));
  NOR2  g03965(.A(new_n4350_), .B(new_n1375_), .Y(new_n4351_));
  NOR2  g03966(.A(new_n4351_), .B(new_n1379_), .Y(new_n4352_));
  NOR2  g03967(.A(new_n4352_), .B(new_n1383_), .Y(new_n4353_));
  NOR2  g03968(.A(new_n4353_), .B(new_n1387_), .Y(new_n4354_));
  NOR2  g03969(.A(new_n4354_), .B(new_n1391_), .Y(new_n4355_));
  NOR2  g03970(.A(new_n4355_), .B(new_n1395_), .Y(new_n4356_));
  NOR2  g03971(.A(new_n4356_), .B(new_n1399_), .Y(new_n4357_));
  NOR2  g03972(.A(new_n4357_), .B(new_n1403_), .Y(new_n4358_));
  NOR2  g03973(.A(new_n4358_), .B(new_n1407_), .Y(new_n4359_));
  NOR2  g03974(.A(new_n4359_), .B(new_n1411_), .Y(new_n4360_));
  NOR2  g03975(.A(new_n4360_), .B(new_n1415_), .Y(new_n4361_));
  NOR2  g03976(.A(new_n4361_), .B(new_n1419_), .Y(new_n4362_));
  NOR2  g03977(.A(new_n4362_), .B(new_n1423_), .Y(new_n4363_));
  NOR2  g03978(.A(new_n4363_), .B(new_n1427_), .Y(new_n4364_));
  NOR2  g03979(.A(new_n4364_), .B(new_n1431_), .Y(new_n4365_));
  NOR2  g03980(.A(new_n4365_), .B(new_n1435_), .Y(new_n4366_));
  NOR2  g03981(.A(new_n4366_), .B(new_n1439_), .Y(new_n4367_));
  NOR2  g03982(.A(new_n4367_), .B(new_n1443_), .Y(new_n4368_));
  NOR2  g03983(.A(new_n4368_), .B(new_n1447_), .Y(new_n4369_));
  NOR2  g03984(.A(new_n4369_), .B(new_n1451_), .Y(new_n4370_));
  NOR2  g03985(.A(new_n4370_), .B(new_n1455_), .Y(new_n4371_));
  NOR2  g03986(.A(new_n4371_), .B(new_n1459_), .Y(new_n4372_));
  NOR2  g03987(.A(new_n4372_), .B(new_n1463_), .Y(new_n4373_));
  NOR2  g03988(.A(new_n4373_), .B(new_n1467_), .Y(new_n4374_));
  NOR2  g03989(.A(new_n4374_), .B(new_n1471_), .Y(new_n4375_));
  NOR2  g03990(.A(new_n4375_), .B(new_n1475_), .Y(new_n4376_));
  NOR2  g03991(.A(new_n4376_), .B(new_n1479_), .Y(new_n4377_));
  NOR2  g03992(.A(new_n4377_), .B(new_n1483_), .Y(new_n4378_));
  NOR2  g03993(.A(new_n4378_), .B(new_n1487_), .Y(new_n4379_));
  NOR2  g03994(.A(new_n4379_), .B(new_n1491_), .Y(new_n4380_));
  NOR2  g03995(.A(new_n4380_), .B(new_n1495_), .Y(new_n4381_));
  NOR2  g03996(.A(new_n4381_), .B(new_n1499_), .Y(new_n4382_));
  NOR2  g03997(.A(new_n4382_), .B(new_n1503_), .Y(new_n4383_));
  NOR2  g03998(.A(new_n4383_), .B(new_n1507_), .Y(new_n4384_));
  NOR2  g03999(.A(new_n4384_), .B(new_n1511_), .Y(new_n4385_));
  NOR2  g04000(.A(new_n4385_), .B(new_n1515_), .Y(new_n4386_));
  NOR2  g04001(.A(new_n4386_), .B(new_n1519_), .Y(new_n4387_));
  NOR2  g04002(.A(new_n4387_), .B(new_n1523_), .Y(new_n4388_));
  NOR2  g04003(.A(new_n4388_), .B(new_n1527_), .Y(new_n4389_));
  NOR2  g04004(.A(new_n4389_), .B(new_n1797_), .Y(new_n4390_));
  NOR2  g04005(.A(new_n4390_), .B(new_n396_), .Y(new_n4391_));
  NOR2  g04006(.A(new_n4391_), .B(new_n400_), .Y(new_n4392_));
  NOR2  g04007(.A(new_n4392_), .B(new_n406_), .Y(new_n4393_));
  NOR2  g04008(.A(new_n4393_), .B(new_n410_), .Y(new_n4394_));
  NOR2  g04009(.A(new_n4394_), .B(new_n416_), .Y(new_n4395_));
  NOR2  g04010(.A(new_n4395_), .B(new_n420_), .Y(new_n4396_));
  NOR2  g04011(.A(new_n4396_), .B(new_n426_), .Y(new_n4397_));
  NOR2  g04012(.A(new_n4397_), .B(new_n430_), .Y(new_n4398_));
  NOR2  g04013(.A(new_n4398_), .B(new_n436_), .Y(new_n4399_));
  NOR2  g04014(.A(new_n4399_), .B(new_n440_), .Y(new_n4400_));
  NOR2  g04015(.A(new_n4400_), .B(new_n446_), .Y(new_n4401_));
  NOR2  g04016(.A(new_n4401_), .B(new_n450_), .Y(new_n4402_));
  NOR2  g04017(.A(new_n4402_), .B(new_n456_), .Y(new_n4403_));
  NOR2  g04018(.A(new_n4403_), .B(new_n460_), .Y(new_n4404_));
  NOR2  g04019(.A(new_n4404_), .B(new_n466_), .Y(new_n4405_));
  NOR2  g04020(.A(new_n4405_), .B(new_n470_), .Y(new_n4406_));
  NOR2  g04021(.A(new_n4406_), .B(new_n476_), .Y(new_n4407_));
  NOR2  g04022(.A(new_n4407_), .B(new_n480_), .Y(new_n4408_));
  NOR2  g04023(.A(new_n4408_), .B(new_n486_), .Y(new_n4409_));
  NOR2  g04024(.A(new_n4409_), .B(new_n490_), .Y(new_n4410_));
  NOR2  g04025(.A(new_n4410_), .B(new_n496_), .Y(new_n4411_));
  NAND2 g04026(.A(new_n498_), .B(\req[35] ), .Y(new_n4412_));
  NOR2  g04027(.A(new_n4412_), .B(new_n4411_), .Y(\grant[35] ));
  INV   g04028(.A(new_n509_), .Y(new_n4414_));
  NOR2  g04029(.A(new_n918_), .B(new_n4414_), .Y(new_n4415_));
  NOR2  g04030(.A(new_n4415_), .B(new_n516_), .Y(new_n4416_));
  NOR2  g04031(.A(new_n4416_), .B(new_n520_), .Y(new_n4417_));
  NOR2  g04032(.A(new_n4417_), .B(new_n526_), .Y(new_n4418_));
  NOR2  g04033(.A(new_n4418_), .B(new_n530_), .Y(new_n4419_));
  NOR2  g04034(.A(new_n4419_), .B(new_n536_), .Y(new_n4420_));
  NOR2  g04035(.A(new_n4420_), .B(new_n540_), .Y(new_n4421_));
  NOR2  g04036(.A(new_n4421_), .B(new_n546_), .Y(new_n4422_));
  NOR2  g04037(.A(new_n4422_), .B(new_n550_), .Y(new_n4423_));
  NOR2  g04038(.A(new_n4423_), .B(new_n556_), .Y(new_n4424_));
  NOR2  g04039(.A(new_n4424_), .B(new_n560_), .Y(new_n4425_));
  NOR2  g04040(.A(new_n4425_), .B(new_n566_), .Y(new_n4426_));
  NOR2  g04041(.A(new_n4426_), .B(new_n570_), .Y(new_n4427_));
  NOR2  g04042(.A(new_n4427_), .B(new_n576_), .Y(new_n4428_));
  NOR2  g04043(.A(new_n4428_), .B(new_n580_), .Y(new_n4429_));
  NOR2  g04044(.A(new_n4429_), .B(new_n586_), .Y(new_n4430_));
  NOR2  g04045(.A(new_n4430_), .B(new_n590_), .Y(new_n4431_));
  NOR2  g04046(.A(new_n4431_), .B(new_n596_), .Y(new_n4432_));
  NOR2  g04047(.A(new_n4432_), .B(new_n600_), .Y(new_n4433_));
  NOR2  g04048(.A(new_n4433_), .B(new_n606_), .Y(new_n4434_));
  NOR2  g04049(.A(new_n4434_), .B(new_n610_), .Y(new_n4435_));
  NOR2  g04050(.A(new_n4435_), .B(new_n616_), .Y(new_n4436_));
  NOR2  g04051(.A(new_n4436_), .B(new_n620_), .Y(new_n4437_));
  NOR2  g04052(.A(new_n4437_), .B(new_n626_), .Y(new_n4438_));
  NOR2  g04053(.A(new_n4438_), .B(new_n630_), .Y(new_n4439_));
  NOR2  g04054(.A(new_n4439_), .B(new_n636_), .Y(new_n4440_));
  NOR2  g04055(.A(new_n4440_), .B(new_n640_), .Y(new_n4441_));
  NOR2  g04056(.A(new_n4441_), .B(new_n646_), .Y(new_n4442_));
  NOR2  g04057(.A(new_n4442_), .B(new_n650_), .Y(new_n4443_));
  NOR2  g04058(.A(new_n4443_), .B(new_n656_), .Y(new_n4444_));
  NOR2  g04059(.A(new_n4444_), .B(new_n660_), .Y(new_n4445_));
  NOR2  g04060(.A(new_n4445_), .B(new_n666_), .Y(new_n4446_));
  NOR2  g04061(.A(new_n4446_), .B(new_n670_), .Y(new_n4447_));
  NOR2  g04062(.A(new_n4447_), .B(new_n676_), .Y(new_n4448_));
  NOR2  g04063(.A(new_n4448_), .B(new_n680_), .Y(new_n4449_));
  NOR2  g04064(.A(new_n4449_), .B(new_n686_), .Y(new_n4450_));
  NOR2  g04065(.A(new_n4450_), .B(new_n690_), .Y(new_n4451_));
  NOR2  g04066(.A(new_n4451_), .B(new_n696_), .Y(new_n4452_));
  NOR2  g04067(.A(new_n4452_), .B(new_n700_), .Y(new_n4453_));
  NOR2  g04068(.A(new_n4453_), .B(new_n706_), .Y(new_n4454_));
  NOR2  g04069(.A(new_n4454_), .B(new_n710_), .Y(new_n4455_));
  NOR2  g04070(.A(new_n4455_), .B(new_n716_), .Y(new_n4456_));
  NOR2  g04071(.A(new_n4456_), .B(new_n720_), .Y(new_n4457_));
  NOR2  g04072(.A(new_n4457_), .B(new_n726_), .Y(new_n4458_));
  NOR2  g04073(.A(new_n4458_), .B(new_n730_), .Y(new_n4459_));
  NOR2  g04074(.A(new_n4459_), .B(new_n736_), .Y(new_n4460_));
  NOR2  g04075(.A(new_n4460_), .B(new_n740_), .Y(new_n4461_));
  NOR2  g04076(.A(new_n4461_), .B(new_n746_), .Y(new_n4462_));
  NOR2  g04077(.A(new_n4462_), .B(new_n750_), .Y(new_n4463_));
  NOR2  g04078(.A(new_n4463_), .B(new_n756_), .Y(new_n4464_));
  NOR2  g04079(.A(new_n4464_), .B(new_n760_), .Y(new_n4465_));
  NOR2  g04080(.A(new_n4465_), .B(new_n766_), .Y(new_n4466_));
  NOR2  g04081(.A(new_n4466_), .B(new_n770_), .Y(new_n4467_));
  NOR2  g04082(.A(new_n4467_), .B(new_n776_), .Y(new_n4468_));
  NOR2  g04083(.A(new_n4468_), .B(new_n780_), .Y(new_n4469_));
  NOR2  g04084(.A(new_n4469_), .B(new_n786_), .Y(new_n4470_));
  NOR2  g04085(.A(new_n4470_), .B(new_n790_), .Y(new_n4471_));
  NOR2  g04086(.A(new_n4471_), .B(new_n796_), .Y(new_n4472_));
  NOR2  g04087(.A(new_n4472_), .B(new_n800_), .Y(new_n4473_));
  NOR2  g04088(.A(new_n4473_), .B(new_n806_), .Y(new_n4474_));
  NOR2  g04089(.A(new_n4474_), .B(new_n1616_), .Y(new_n4475_));
  NOR2  g04090(.A(new_n4475_), .B(new_n1618_), .Y(new_n4476_));
  NOR2  g04091(.A(new_n4476_), .B(new_n1885_), .Y(new_n4477_));
  NOR2  g04092(.A(new_n4477_), .B(new_n820_), .Y(new_n4478_));
  NOR2  g04093(.A(new_n4478_), .B(new_n824_), .Y(new_n4479_));
  NOR2  g04094(.A(new_n4479_), .B(new_n829_), .Y(new_n4480_));
  NOR2  g04095(.A(new_n4480_), .B(new_n833_), .Y(new_n4481_));
  NOR2  g04096(.A(new_n4481_), .B(new_n838_), .Y(new_n4482_));
  NOR2  g04097(.A(new_n4482_), .B(new_n842_), .Y(new_n4483_));
  NOR2  g04098(.A(new_n4483_), .B(new_n847_), .Y(new_n4484_));
  NOR2  g04099(.A(new_n4484_), .B(new_n851_), .Y(new_n4485_));
  NOR2  g04100(.A(new_n4485_), .B(new_n856_), .Y(new_n4486_));
  NOR2  g04101(.A(new_n4486_), .B(new_n860_), .Y(new_n4487_));
  NOR2  g04102(.A(new_n4487_), .B(new_n865_), .Y(new_n4488_));
  NOR2  g04103(.A(new_n4488_), .B(new_n869_), .Y(new_n4489_));
  NOR2  g04104(.A(new_n4489_), .B(new_n874_), .Y(new_n4490_));
  NOR2  g04105(.A(new_n4490_), .B(new_n878_), .Y(new_n4491_));
  NOR2  g04106(.A(new_n4491_), .B(new_n883_), .Y(new_n4492_));
  NOR2  g04107(.A(new_n4492_), .B(new_n887_), .Y(new_n4493_));
  NOR2  g04108(.A(new_n4493_), .B(new_n892_), .Y(new_n4494_));
  NOR2  g04109(.A(new_n4494_), .B(new_n896_), .Y(new_n4495_));
  NOR2  g04110(.A(new_n4495_), .B(new_n901_), .Y(new_n4496_));
  NOR2  g04111(.A(new_n4496_), .B(new_n905_), .Y(new_n4497_));
  NOR2  g04112(.A(new_n4497_), .B(new_n910_), .Y(new_n4498_));
  NAND2 g04113(.A(new_n912_), .B(\req[36] ), .Y(new_n4499_));
  NOR2  g04114(.A(new_n4499_), .B(new_n4498_), .Y(\grant[36] ));
  INV   g04115(.A(new_n922_), .Y(new_n4501_));
  NOR2  g04116(.A(new_n1286_), .B(new_n4501_), .Y(new_n4502_));
  NOR2  g04117(.A(new_n4502_), .B(new_n928_), .Y(new_n4503_));
  NOR2  g04118(.A(new_n4503_), .B(new_n932_), .Y(new_n4504_));
  NOR2  g04119(.A(new_n4504_), .B(new_n937_), .Y(new_n4505_));
  NOR2  g04120(.A(new_n4505_), .B(new_n941_), .Y(new_n4506_));
  NOR2  g04121(.A(new_n4506_), .B(new_n946_), .Y(new_n4507_));
  NOR2  g04122(.A(new_n4507_), .B(new_n950_), .Y(new_n4508_));
  NOR2  g04123(.A(new_n4508_), .B(new_n955_), .Y(new_n4509_));
  NOR2  g04124(.A(new_n4509_), .B(new_n959_), .Y(new_n4510_));
  NOR2  g04125(.A(new_n4510_), .B(new_n964_), .Y(new_n4511_));
  NOR2  g04126(.A(new_n4511_), .B(new_n968_), .Y(new_n4512_));
  NOR2  g04127(.A(new_n4512_), .B(new_n973_), .Y(new_n4513_));
  NOR2  g04128(.A(new_n4513_), .B(new_n977_), .Y(new_n4514_));
  NOR2  g04129(.A(new_n4514_), .B(new_n982_), .Y(new_n4515_));
  NOR2  g04130(.A(new_n4515_), .B(new_n986_), .Y(new_n4516_));
  NOR2  g04131(.A(new_n4516_), .B(new_n991_), .Y(new_n4517_));
  NOR2  g04132(.A(new_n4517_), .B(new_n995_), .Y(new_n4518_));
  NOR2  g04133(.A(new_n4518_), .B(new_n1000_), .Y(new_n4519_));
  NOR2  g04134(.A(new_n4519_), .B(new_n1004_), .Y(new_n4520_));
  NOR2  g04135(.A(new_n4520_), .B(new_n1009_), .Y(new_n4521_));
  NOR2  g04136(.A(new_n4521_), .B(new_n1013_), .Y(new_n4522_));
  NOR2  g04137(.A(new_n4522_), .B(new_n1018_), .Y(new_n4523_));
  NOR2  g04138(.A(new_n4523_), .B(new_n1022_), .Y(new_n4524_));
  NOR2  g04139(.A(new_n4524_), .B(new_n1027_), .Y(new_n4525_));
  NOR2  g04140(.A(new_n4525_), .B(new_n1031_), .Y(new_n4526_));
  NOR2  g04141(.A(new_n4526_), .B(new_n1036_), .Y(new_n4527_));
  NOR2  g04142(.A(new_n4527_), .B(new_n1040_), .Y(new_n4528_));
  NOR2  g04143(.A(new_n4528_), .B(new_n1045_), .Y(new_n4529_));
  NOR2  g04144(.A(new_n4529_), .B(new_n1049_), .Y(new_n4530_));
  NOR2  g04145(.A(new_n4530_), .B(new_n1054_), .Y(new_n4531_));
  NOR2  g04146(.A(new_n4531_), .B(new_n1058_), .Y(new_n4532_));
  NOR2  g04147(.A(new_n4532_), .B(new_n1063_), .Y(new_n4533_));
  NOR2  g04148(.A(new_n4533_), .B(new_n1067_), .Y(new_n4534_));
  NOR2  g04149(.A(new_n4534_), .B(new_n1072_), .Y(new_n4535_));
  NOR2  g04150(.A(new_n4535_), .B(new_n1076_), .Y(new_n4536_));
  NOR2  g04151(.A(new_n4536_), .B(new_n1081_), .Y(new_n4537_));
  NOR2  g04152(.A(new_n4537_), .B(new_n1085_), .Y(new_n4538_));
  NOR2  g04153(.A(new_n4538_), .B(new_n1090_), .Y(new_n4539_));
  NOR2  g04154(.A(new_n4539_), .B(new_n1094_), .Y(new_n4540_));
  NOR2  g04155(.A(new_n4540_), .B(new_n1099_), .Y(new_n4541_));
  NOR2  g04156(.A(new_n4541_), .B(new_n1103_), .Y(new_n4542_));
  NOR2  g04157(.A(new_n4542_), .B(new_n1108_), .Y(new_n4543_));
  NOR2  g04158(.A(new_n4543_), .B(new_n1112_), .Y(new_n4544_));
  NOR2  g04159(.A(new_n4544_), .B(new_n1117_), .Y(new_n4545_));
  NOR2  g04160(.A(new_n4545_), .B(new_n1121_), .Y(new_n4546_));
  NOR2  g04161(.A(new_n4546_), .B(new_n1126_), .Y(new_n4547_));
  NOR2  g04162(.A(new_n4547_), .B(new_n1130_), .Y(new_n4548_));
  NOR2  g04163(.A(new_n4548_), .B(new_n1135_), .Y(new_n4549_));
  NOR2  g04164(.A(new_n4549_), .B(new_n1139_), .Y(new_n4550_));
  NOR2  g04165(.A(new_n4550_), .B(new_n1144_), .Y(new_n4551_));
  NOR2  g04166(.A(new_n4551_), .B(new_n1148_), .Y(new_n4552_));
  NOR2  g04167(.A(new_n4552_), .B(new_n1153_), .Y(new_n4553_));
  NOR2  g04168(.A(new_n4553_), .B(new_n1157_), .Y(new_n4554_));
  NOR2  g04169(.A(new_n4554_), .B(new_n1162_), .Y(new_n4555_));
  NOR2  g04170(.A(new_n4555_), .B(new_n1166_), .Y(new_n4556_));
  NOR2  g04171(.A(new_n4556_), .B(new_n1171_), .Y(new_n4557_));
  NOR2  g04172(.A(new_n4557_), .B(new_n1175_), .Y(new_n4558_));
  NOR2  g04173(.A(new_n4558_), .B(new_n1180_), .Y(new_n4559_));
  NOR2  g04174(.A(new_n4559_), .B(new_n1184_), .Y(new_n4560_));
  NOR2  g04175(.A(new_n4560_), .B(new_n1189_), .Y(new_n4561_));
  NOR2  g04176(.A(new_n4561_), .B(new_n1707_), .Y(new_n4562_));
  NOR2  g04177(.A(new_n4562_), .B(new_n1709_), .Y(new_n4563_));
  NOR2  g04178(.A(new_n4563_), .B(new_n1973_), .Y(new_n4564_));
  NOR2  g04179(.A(new_n4564_), .B(new_n1199_), .Y(new_n4565_));
  NOR2  g04180(.A(new_n4565_), .B(new_n1203_), .Y(new_n4566_));
  NOR2  g04181(.A(new_n4566_), .B(new_n1207_), .Y(new_n4567_));
  NOR2  g04182(.A(new_n4567_), .B(new_n1211_), .Y(new_n4568_));
  NOR2  g04183(.A(new_n4568_), .B(new_n1215_), .Y(new_n4569_));
  NOR2  g04184(.A(new_n4569_), .B(new_n1219_), .Y(new_n4570_));
  NOR2  g04185(.A(new_n4570_), .B(new_n1223_), .Y(new_n4571_));
  NOR2  g04186(.A(new_n4571_), .B(new_n1227_), .Y(new_n4572_));
  NOR2  g04187(.A(new_n4572_), .B(new_n1231_), .Y(new_n4573_));
  NOR2  g04188(.A(new_n4573_), .B(new_n1235_), .Y(new_n4574_));
  NOR2  g04189(.A(new_n4574_), .B(new_n1239_), .Y(new_n4575_));
  NOR2  g04190(.A(new_n4575_), .B(new_n1243_), .Y(new_n4576_));
  NOR2  g04191(.A(new_n4576_), .B(new_n1247_), .Y(new_n4577_));
  NOR2  g04192(.A(new_n4577_), .B(new_n1251_), .Y(new_n4578_));
  NOR2  g04193(.A(new_n4578_), .B(new_n1255_), .Y(new_n4579_));
  NOR2  g04194(.A(new_n4579_), .B(new_n1259_), .Y(new_n4580_));
  NOR2  g04195(.A(new_n4580_), .B(new_n1263_), .Y(new_n4581_));
  NOR2  g04196(.A(new_n4581_), .B(new_n1267_), .Y(new_n4582_));
  NOR2  g04197(.A(new_n4582_), .B(new_n1271_), .Y(new_n4583_));
  NOR2  g04198(.A(new_n4583_), .B(new_n1275_), .Y(new_n4584_));
  NOR2  g04199(.A(new_n4584_), .B(new_n1279_), .Y(new_n4585_));
  NAND2 g04200(.A(new_n1281_), .B(\req[37] ), .Y(new_n4586_));
  NOR2  g04201(.A(new_n4586_), .B(new_n4585_), .Y(\grant[37] ));
  INV   g04202(.A(new_n1290_), .Y(new_n4588_));
  NOR2  g04203(.A(new_n4588_), .B(new_n515_), .Y(new_n4589_));
  NOR2  g04204(.A(new_n4589_), .B(new_n1295_), .Y(new_n4590_));
  NOR2  g04205(.A(new_n4590_), .B(new_n1299_), .Y(new_n4591_));
  NOR2  g04206(.A(new_n4591_), .B(new_n1303_), .Y(new_n4592_));
  NOR2  g04207(.A(new_n4592_), .B(new_n1307_), .Y(new_n4593_));
  NOR2  g04208(.A(new_n4593_), .B(new_n1311_), .Y(new_n4594_));
  NOR2  g04209(.A(new_n4594_), .B(new_n1315_), .Y(new_n4595_));
  NOR2  g04210(.A(new_n4595_), .B(new_n1319_), .Y(new_n4596_));
  NOR2  g04211(.A(new_n4596_), .B(new_n1323_), .Y(new_n4597_));
  NOR2  g04212(.A(new_n4597_), .B(new_n1327_), .Y(new_n4598_));
  NOR2  g04213(.A(new_n4598_), .B(new_n1331_), .Y(new_n4599_));
  NOR2  g04214(.A(new_n4599_), .B(new_n1335_), .Y(new_n4600_));
  NOR2  g04215(.A(new_n4600_), .B(new_n1339_), .Y(new_n4601_));
  NOR2  g04216(.A(new_n4601_), .B(new_n1343_), .Y(new_n4602_));
  NOR2  g04217(.A(new_n4602_), .B(new_n1347_), .Y(new_n4603_));
  NOR2  g04218(.A(new_n4603_), .B(new_n1351_), .Y(new_n4604_));
  NOR2  g04219(.A(new_n4604_), .B(new_n1355_), .Y(new_n4605_));
  NOR2  g04220(.A(new_n4605_), .B(new_n1359_), .Y(new_n4606_));
  NOR2  g04221(.A(new_n4606_), .B(new_n1363_), .Y(new_n4607_));
  NOR2  g04222(.A(new_n4607_), .B(new_n1367_), .Y(new_n4608_));
  NOR2  g04223(.A(new_n4608_), .B(new_n1371_), .Y(new_n4609_));
  NOR2  g04224(.A(new_n4609_), .B(new_n1375_), .Y(new_n4610_));
  NOR2  g04225(.A(new_n4610_), .B(new_n1379_), .Y(new_n4611_));
  NOR2  g04226(.A(new_n4611_), .B(new_n1383_), .Y(new_n4612_));
  NOR2  g04227(.A(new_n4612_), .B(new_n1387_), .Y(new_n4613_));
  NOR2  g04228(.A(new_n4613_), .B(new_n1391_), .Y(new_n4614_));
  NOR2  g04229(.A(new_n4614_), .B(new_n1395_), .Y(new_n4615_));
  NOR2  g04230(.A(new_n4615_), .B(new_n1399_), .Y(new_n4616_));
  NOR2  g04231(.A(new_n4616_), .B(new_n1403_), .Y(new_n4617_));
  NOR2  g04232(.A(new_n4617_), .B(new_n1407_), .Y(new_n4618_));
  NOR2  g04233(.A(new_n4618_), .B(new_n1411_), .Y(new_n4619_));
  NOR2  g04234(.A(new_n4619_), .B(new_n1415_), .Y(new_n4620_));
  NOR2  g04235(.A(new_n4620_), .B(new_n1419_), .Y(new_n4621_));
  NOR2  g04236(.A(new_n4621_), .B(new_n1423_), .Y(new_n4622_));
  NOR2  g04237(.A(new_n4622_), .B(new_n1427_), .Y(new_n4623_));
  NOR2  g04238(.A(new_n4623_), .B(new_n1431_), .Y(new_n4624_));
  NOR2  g04239(.A(new_n4624_), .B(new_n1435_), .Y(new_n4625_));
  NOR2  g04240(.A(new_n4625_), .B(new_n1439_), .Y(new_n4626_));
  NOR2  g04241(.A(new_n4626_), .B(new_n1443_), .Y(new_n4627_));
  NOR2  g04242(.A(new_n4627_), .B(new_n1447_), .Y(new_n4628_));
  NOR2  g04243(.A(new_n4628_), .B(new_n1451_), .Y(new_n4629_));
  NOR2  g04244(.A(new_n4629_), .B(new_n1455_), .Y(new_n4630_));
  NOR2  g04245(.A(new_n4630_), .B(new_n1459_), .Y(new_n4631_));
  NOR2  g04246(.A(new_n4631_), .B(new_n1463_), .Y(new_n4632_));
  NOR2  g04247(.A(new_n4632_), .B(new_n1467_), .Y(new_n4633_));
  NOR2  g04248(.A(new_n4633_), .B(new_n1471_), .Y(new_n4634_));
  NOR2  g04249(.A(new_n4634_), .B(new_n1475_), .Y(new_n4635_));
  NOR2  g04250(.A(new_n4635_), .B(new_n1479_), .Y(new_n4636_));
  NOR2  g04251(.A(new_n4636_), .B(new_n1483_), .Y(new_n4637_));
  NOR2  g04252(.A(new_n4637_), .B(new_n1487_), .Y(new_n4638_));
  NOR2  g04253(.A(new_n4638_), .B(new_n1491_), .Y(new_n4639_));
  NOR2  g04254(.A(new_n4639_), .B(new_n1495_), .Y(new_n4640_));
  NOR2  g04255(.A(new_n4640_), .B(new_n1499_), .Y(new_n4641_));
  NOR2  g04256(.A(new_n4641_), .B(new_n1503_), .Y(new_n4642_));
  NOR2  g04257(.A(new_n4642_), .B(new_n1507_), .Y(new_n4643_));
  NOR2  g04258(.A(new_n4643_), .B(new_n1511_), .Y(new_n4644_));
  NOR2  g04259(.A(new_n4644_), .B(new_n1515_), .Y(new_n4645_));
  NOR2  g04260(.A(new_n4645_), .B(new_n1519_), .Y(new_n4646_));
  NOR2  g04261(.A(new_n4646_), .B(new_n1523_), .Y(new_n4647_));
  NOR2  g04262(.A(new_n4647_), .B(new_n1527_), .Y(new_n4648_));
  NOR2  g04263(.A(new_n4648_), .B(new_n1797_), .Y(new_n4649_));
  NOR2  g04264(.A(new_n4649_), .B(new_n396_), .Y(new_n4650_));
  NOR2  g04265(.A(new_n4650_), .B(new_n400_), .Y(new_n4651_));
  NOR2  g04266(.A(new_n4651_), .B(new_n406_), .Y(new_n4652_));
  NOR2  g04267(.A(new_n4652_), .B(new_n410_), .Y(new_n4653_));
  NOR2  g04268(.A(new_n4653_), .B(new_n416_), .Y(new_n4654_));
  NOR2  g04269(.A(new_n4654_), .B(new_n420_), .Y(new_n4655_));
  NOR2  g04270(.A(new_n4655_), .B(new_n426_), .Y(new_n4656_));
  NOR2  g04271(.A(new_n4656_), .B(new_n430_), .Y(new_n4657_));
  NOR2  g04272(.A(new_n4657_), .B(new_n436_), .Y(new_n4658_));
  NOR2  g04273(.A(new_n4658_), .B(new_n440_), .Y(new_n4659_));
  NOR2  g04274(.A(new_n4659_), .B(new_n446_), .Y(new_n4660_));
  NOR2  g04275(.A(new_n4660_), .B(new_n450_), .Y(new_n4661_));
  NOR2  g04276(.A(new_n4661_), .B(new_n456_), .Y(new_n4662_));
  NOR2  g04277(.A(new_n4662_), .B(new_n460_), .Y(new_n4663_));
  NOR2  g04278(.A(new_n4663_), .B(new_n466_), .Y(new_n4664_));
  NOR2  g04279(.A(new_n4664_), .B(new_n470_), .Y(new_n4665_));
  NOR2  g04280(.A(new_n4665_), .B(new_n476_), .Y(new_n4666_));
  NOR2  g04281(.A(new_n4666_), .B(new_n480_), .Y(new_n4667_));
  NOR2  g04282(.A(new_n4667_), .B(new_n486_), .Y(new_n4668_));
  NOR2  g04283(.A(new_n4668_), .B(new_n490_), .Y(new_n4669_));
  NOR2  g04284(.A(new_n4669_), .B(new_n496_), .Y(new_n4670_));
  NOR2  g04285(.A(new_n4670_), .B(new_n500_), .Y(new_n4671_));
  NOR2  g04286(.A(new_n4671_), .B(new_n506_), .Y(new_n4672_));
  NAND2 g04287(.A(new_n508_), .B(\req[38] ), .Y(new_n4673_));
  NOR2  g04288(.A(new_n4673_), .B(new_n4672_), .Y(\grant[38] ));
  INV   g04289(.A(new_n519_), .Y(new_n4675_));
  NOR2  g04290(.A(new_n927_), .B(new_n4675_), .Y(new_n4676_));
  NOR2  g04291(.A(new_n4676_), .B(new_n526_), .Y(new_n4677_));
  NOR2  g04292(.A(new_n4677_), .B(new_n530_), .Y(new_n4678_));
  NOR2  g04293(.A(new_n4678_), .B(new_n536_), .Y(new_n4679_));
  NOR2  g04294(.A(new_n4679_), .B(new_n540_), .Y(new_n4680_));
  NOR2  g04295(.A(new_n4680_), .B(new_n546_), .Y(new_n4681_));
  NOR2  g04296(.A(new_n4681_), .B(new_n550_), .Y(new_n4682_));
  NOR2  g04297(.A(new_n4682_), .B(new_n556_), .Y(new_n4683_));
  NOR2  g04298(.A(new_n4683_), .B(new_n560_), .Y(new_n4684_));
  NOR2  g04299(.A(new_n4684_), .B(new_n566_), .Y(new_n4685_));
  NOR2  g04300(.A(new_n4685_), .B(new_n570_), .Y(new_n4686_));
  NOR2  g04301(.A(new_n4686_), .B(new_n576_), .Y(new_n4687_));
  NOR2  g04302(.A(new_n4687_), .B(new_n580_), .Y(new_n4688_));
  NOR2  g04303(.A(new_n4688_), .B(new_n586_), .Y(new_n4689_));
  NOR2  g04304(.A(new_n4689_), .B(new_n590_), .Y(new_n4690_));
  NOR2  g04305(.A(new_n4690_), .B(new_n596_), .Y(new_n4691_));
  NOR2  g04306(.A(new_n4691_), .B(new_n600_), .Y(new_n4692_));
  NOR2  g04307(.A(new_n4692_), .B(new_n606_), .Y(new_n4693_));
  NOR2  g04308(.A(new_n4693_), .B(new_n610_), .Y(new_n4694_));
  NOR2  g04309(.A(new_n4694_), .B(new_n616_), .Y(new_n4695_));
  NOR2  g04310(.A(new_n4695_), .B(new_n620_), .Y(new_n4696_));
  NOR2  g04311(.A(new_n4696_), .B(new_n626_), .Y(new_n4697_));
  NOR2  g04312(.A(new_n4697_), .B(new_n630_), .Y(new_n4698_));
  NOR2  g04313(.A(new_n4698_), .B(new_n636_), .Y(new_n4699_));
  NOR2  g04314(.A(new_n4699_), .B(new_n640_), .Y(new_n4700_));
  NOR2  g04315(.A(new_n4700_), .B(new_n646_), .Y(new_n4701_));
  NOR2  g04316(.A(new_n4701_), .B(new_n650_), .Y(new_n4702_));
  NOR2  g04317(.A(new_n4702_), .B(new_n656_), .Y(new_n4703_));
  NOR2  g04318(.A(new_n4703_), .B(new_n660_), .Y(new_n4704_));
  NOR2  g04319(.A(new_n4704_), .B(new_n666_), .Y(new_n4705_));
  NOR2  g04320(.A(new_n4705_), .B(new_n670_), .Y(new_n4706_));
  NOR2  g04321(.A(new_n4706_), .B(new_n676_), .Y(new_n4707_));
  NOR2  g04322(.A(new_n4707_), .B(new_n680_), .Y(new_n4708_));
  NOR2  g04323(.A(new_n4708_), .B(new_n686_), .Y(new_n4709_));
  NOR2  g04324(.A(new_n4709_), .B(new_n690_), .Y(new_n4710_));
  NOR2  g04325(.A(new_n4710_), .B(new_n696_), .Y(new_n4711_));
  NOR2  g04326(.A(new_n4711_), .B(new_n700_), .Y(new_n4712_));
  NOR2  g04327(.A(new_n4712_), .B(new_n706_), .Y(new_n4713_));
  NOR2  g04328(.A(new_n4713_), .B(new_n710_), .Y(new_n4714_));
  NOR2  g04329(.A(new_n4714_), .B(new_n716_), .Y(new_n4715_));
  NOR2  g04330(.A(new_n4715_), .B(new_n720_), .Y(new_n4716_));
  NOR2  g04331(.A(new_n4716_), .B(new_n726_), .Y(new_n4717_));
  NOR2  g04332(.A(new_n4717_), .B(new_n730_), .Y(new_n4718_));
  NOR2  g04333(.A(new_n4718_), .B(new_n736_), .Y(new_n4719_));
  NOR2  g04334(.A(new_n4719_), .B(new_n740_), .Y(new_n4720_));
  NOR2  g04335(.A(new_n4720_), .B(new_n746_), .Y(new_n4721_));
  NOR2  g04336(.A(new_n4721_), .B(new_n750_), .Y(new_n4722_));
  NOR2  g04337(.A(new_n4722_), .B(new_n756_), .Y(new_n4723_));
  NOR2  g04338(.A(new_n4723_), .B(new_n760_), .Y(new_n4724_));
  NOR2  g04339(.A(new_n4724_), .B(new_n766_), .Y(new_n4725_));
  NOR2  g04340(.A(new_n4725_), .B(new_n770_), .Y(new_n4726_));
  NOR2  g04341(.A(new_n4726_), .B(new_n776_), .Y(new_n4727_));
  NOR2  g04342(.A(new_n4727_), .B(new_n780_), .Y(new_n4728_));
  NOR2  g04343(.A(new_n4728_), .B(new_n786_), .Y(new_n4729_));
  NOR2  g04344(.A(new_n4729_), .B(new_n790_), .Y(new_n4730_));
  NOR2  g04345(.A(new_n4730_), .B(new_n796_), .Y(new_n4731_));
  NOR2  g04346(.A(new_n4731_), .B(new_n800_), .Y(new_n4732_));
  NOR2  g04347(.A(new_n4732_), .B(new_n806_), .Y(new_n4733_));
  NOR2  g04348(.A(new_n4733_), .B(new_n1616_), .Y(new_n4734_));
  NOR2  g04349(.A(new_n4734_), .B(new_n1618_), .Y(new_n4735_));
  NOR2  g04350(.A(new_n4735_), .B(new_n1885_), .Y(new_n4736_));
  NOR2  g04351(.A(new_n4736_), .B(new_n820_), .Y(new_n4737_));
  NOR2  g04352(.A(new_n4737_), .B(new_n824_), .Y(new_n4738_));
  NOR2  g04353(.A(new_n4738_), .B(new_n829_), .Y(new_n4739_));
  NOR2  g04354(.A(new_n4739_), .B(new_n833_), .Y(new_n4740_));
  NOR2  g04355(.A(new_n4740_), .B(new_n838_), .Y(new_n4741_));
  NOR2  g04356(.A(new_n4741_), .B(new_n842_), .Y(new_n4742_));
  NOR2  g04357(.A(new_n4742_), .B(new_n847_), .Y(new_n4743_));
  NOR2  g04358(.A(new_n4743_), .B(new_n851_), .Y(new_n4744_));
  NOR2  g04359(.A(new_n4744_), .B(new_n856_), .Y(new_n4745_));
  NOR2  g04360(.A(new_n4745_), .B(new_n860_), .Y(new_n4746_));
  NOR2  g04361(.A(new_n4746_), .B(new_n865_), .Y(new_n4747_));
  NOR2  g04362(.A(new_n4747_), .B(new_n869_), .Y(new_n4748_));
  NOR2  g04363(.A(new_n4748_), .B(new_n874_), .Y(new_n4749_));
  NOR2  g04364(.A(new_n4749_), .B(new_n878_), .Y(new_n4750_));
  NOR2  g04365(.A(new_n4750_), .B(new_n883_), .Y(new_n4751_));
  NOR2  g04366(.A(new_n4751_), .B(new_n887_), .Y(new_n4752_));
  NOR2  g04367(.A(new_n4752_), .B(new_n892_), .Y(new_n4753_));
  NOR2  g04368(.A(new_n4753_), .B(new_n896_), .Y(new_n4754_));
  NOR2  g04369(.A(new_n4754_), .B(new_n901_), .Y(new_n4755_));
  NOR2  g04370(.A(new_n4755_), .B(new_n905_), .Y(new_n4756_));
  NOR2  g04371(.A(new_n4756_), .B(new_n910_), .Y(new_n4757_));
  NOR2  g04372(.A(new_n4757_), .B(new_n914_), .Y(new_n4758_));
  NOR2  g04373(.A(new_n4758_), .B(new_n919_), .Y(new_n4759_));
  NAND2 g04374(.A(new_n921_), .B(\req[39] ), .Y(new_n4760_));
  NOR2  g04375(.A(new_n4760_), .B(new_n4759_), .Y(\grant[39] ));
  INV   g04376(.A(new_n931_), .Y(new_n4762_));
  NOR2  g04377(.A(new_n1294_), .B(new_n4762_), .Y(new_n4763_));
  NOR2  g04378(.A(new_n4763_), .B(new_n937_), .Y(new_n4764_));
  NOR2  g04379(.A(new_n4764_), .B(new_n941_), .Y(new_n4765_));
  NOR2  g04380(.A(new_n4765_), .B(new_n946_), .Y(new_n4766_));
  NOR2  g04381(.A(new_n4766_), .B(new_n950_), .Y(new_n4767_));
  NOR2  g04382(.A(new_n4767_), .B(new_n955_), .Y(new_n4768_));
  NOR2  g04383(.A(new_n4768_), .B(new_n959_), .Y(new_n4769_));
  NOR2  g04384(.A(new_n4769_), .B(new_n964_), .Y(new_n4770_));
  NOR2  g04385(.A(new_n4770_), .B(new_n968_), .Y(new_n4771_));
  NOR2  g04386(.A(new_n4771_), .B(new_n973_), .Y(new_n4772_));
  NOR2  g04387(.A(new_n4772_), .B(new_n977_), .Y(new_n4773_));
  NOR2  g04388(.A(new_n4773_), .B(new_n982_), .Y(new_n4774_));
  NOR2  g04389(.A(new_n4774_), .B(new_n986_), .Y(new_n4775_));
  NOR2  g04390(.A(new_n4775_), .B(new_n991_), .Y(new_n4776_));
  NOR2  g04391(.A(new_n4776_), .B(new_n995_), .Y(new_n4777_));
  NOR2  g04392(.A(new_n4777_), .B(new_n1000_), .Y(new_n4778_));
  NOR2  g04393(.A(new_n4778_), .B(new_n1004_), .Y(new_n4779_));
  NOR2  g04394(.A(new_n4779_), .B(new_n1009_), .Y(new_n4780_));
  NOR2  g04395(.A(new_n4780_), .B(new_n1013_), .Y(new_n4781_));
  NOR2  g04396(.A(new_n4781_), .B(new_n1018_), .Y(new_n4782_));
  NOR2  g04397(.A(new_n4782_), .B(new_n1022_), .Y(new_n4783_));
  NOR2  g04398(.A(new_n4783_), .B(new_n1027_), .Y(new_n4784_));
  NOR2  g04399(.A(new_n4784_), .B(new_n1031_), .Y(new_n4785_));
  NOR2  g04400(.A(new_n4785_), .B(new_n1036_), .Y(new_n4786_));
  NOR2  g04401(.A(new_n4786_), .B(new_n1040_), .Y(new_n4787_));
  NOR2  g04402(.A(new_n4787_), .B(new_n1045_), .Y(new_n4788_));
  NOR2  g04403(.A(new_n4788_), .B(new_n1049_), .Y(new_n4789_));
  NOR2  g04404(.A(new_n4789_), .B(new_n1054_), .Y(new_n4790_));
  NOR2  g04405(.A(new_n4790_), .B(new_n1058_), .Y(new_n4791_));
  NOR2  g04406(.A(new_n4791_), .B(new_n1063_), .Y(new_n4792_));
  NOR2  g04407(.A(new_n4792_), .B(new_n1067_), .Y(new_n4793_));
  NOR2  g04408(.A(new_n4793_), .B(new_n1072_), .Y(new_n4794_));
  NOR2  g04409(.A(new_n4794_), .B(new_n1076_), .Y(new_n4795_));
  NOR2  g04410(.A(new_n4795_), .B(new_n1081_), .Y(new_n4796_));
  NOR2  g04411(.A(new_n4796_), .B(new_n1085_), .Y(new_n4797_));
  NOR2  g04412(.A(new_n4797_), .B(new_n1090_), .Y(new_n4798_));
  NOR2  g04413(.A(new_n4798_), .B(new_n1094_), .Y(new_n4799_));
  NOR2  g04414(.A(new_n4799_), .B(new_n1099_), .Y(new_n4800_));
  NOR2  g04415(.A(new_n4800_), .B(new_n1103_), .Y(new_n4801_));
  NOR2  g04416(.A(new_n4801_), .B(new_n1108_), .Y(new_n4802_));
  NOR2  g04417(.A(new_n4802_), .B(new_n1112_), .Y(new_n4803_));
  NOR2  g04418(.A(new_n4803_), .B(new_n1117_), .Y(new_n4804_));
  NOR2  g04419(.A(new_n4804_), .B(new_n1121_), .Y(new_n4805_));
  NOR2  g04420(.A(new_n4805_), .B(new_n1126_), .Y(new_n4806_));
  NOR2  g04421(.A(new_n4806_), .B(new_n1130_), .Y(new_n4807_));
  NOR2  g04422(.A(new_n4807_), .B(new_n1135_), .Y(new_n4808_));
  NOR2  g04423(.A(new_n4808_), .B(new_n1139_), .Y(new_n4809_));
  NOR2  g04424(.A(new_n4809_), .B(new_n1144_), .Y(new_n4810_));
  NOR2  g04425(.A(new_n4810_), .B(new_n1148_), .Y(new_n4811_));
  NOR2  g04426(.A(new_n4811_), .B(new_n1153_), .Y(new_n4812_));
  NOR2  g04427(.A(new_n4812_), .B(new_n1157_), .Y(new_n4813_));
  NOR2  g04428(.A(new_n4813_), .B(new_n1162_), .Y(new_n4814_));
  NOR2  g04429(.A(new_n4814_), .B(new_n1166_), .Y(new_n4815_));
  NOR2  g04430(.A(new_n4815_), .B(new_n1171_), .Y(new_n4816_));
  NOR2  g04431(.A(new_n4816_), .B(new_n1175_), .Y(new_n4817_));
  NOR2  g04432(.A(new_n4817_), .B(new_n1180_), .Y(new_n4818_));
  NOR2  g04433(.A(new_n4818_), .B(new_n1184_), .Y(new_n4819_));
  NOR2  g04434(.A(new_n4819_), .B(new_n1189_), .Y(new_n4820_));
  NOR2  g04435(.A(new_n4820_), .B(new_n1707_), .Y(new_n4821_));
  NOR2  g04436(.A(new_n4821_), .B(new_n1709_), .Y(new_n4822_));
  NOR2  g04437(.A(new_n4822_), .B(new_n1973_), .Y(new_n4823_));
  NOR2  g04438(.A(new_n4823_), .B(new_n1199_), .Y(new_n4824_));
  NOR2  g04439(.A(new_n4824_), .B(new_n1203_), .Y(new_n4825_));
  NOR2  g04440(.A(new_n4825_), .B(new_n1207_), .Y(new_n4826_));
  NOR2  g04441(.A(new_n4826_), .B(new_n1211_), .Y(new_n4827_));
  NOR2  g04442(.A(new_n4827_), .B(new_n1215_), .Y(new_n4828_));
  NOR2  g04443(.A(new_n4828_), .B(new_n1219_), .Y(new_n4829_));
  NOR2  g04444(.A(new_n4829_), .B(new_n1223_), .Y(new_n4830_));
  NOR2  g04445(.A(new_n4830_), .B(new_n1227_), .Y(new_n4831_));
  NOR2  g04446(.A(new_n4831_), .B(new_n1231_), .Y(new_n4832_));
  NOR2  g04447(.A(new_n4832_), .B(new_n1235_), .Y(new_n4833_));
  NOR2  g04448(.A(new_n4833_), .B(new_n1239_), .Y(new_n4834_));
  NOR2  g04449(.A(new_n4834_), .B(new_n1243_), .Y(new_n4835_));
  NOR2  g04450(.A(new_n4835_), .B(new_n1247_), .Y(new_n4836_));
  NOR2  g04451(.A(new_n4836_), .B(new_n1251_), .Y(new_n4837_));
  NOR2  g04452(.A(new_n4837_), .B(new_n1255_), .Y(new_n4838_));
  NOR2  g04453(.A(new_n4838_), .B(new_n1259_), .Y(new_n4839_));
  NOR2  g04454(.A(new_n4839_), .B(new_n1263_), .Y(new_n4840_));
  NOR2  g04455(.A(new_n4840_), .B(new_n1267_), .Y(new_n4841_));
  NOR2  g04456(.A(new_n4841_), .B(new_n1271_), .Y(new_n4842_));
  NOR2  g04457(.A(new_n4842_), .B(new_n1275_), .Y(new_n4843_));
  NOR2  g04458(.A(new_n4843_), .B(new_n1279_), .Y(new_n4844_));
  NOR2  g04459(.A(new_n4844_), .B(new_n1283_), .Y(new_n4845_));
  NOR2  g04460(.A(new_n4845_), .B(new_n1287_), .Y(new_n4846_));
  NAND2 g04461(.A(new_n1289_), .B(\req[40] ), .Y(new_n4847_));
  NOR2  g04462(.A(new_n4847_), .B(new_n4846_), .Y(\grant[40] ));
  INV   g04463(.A(new_n1298_), .Y(new_n4849_));
  NOR2  g04464(.A(new_n4849_), .B(new_n525_), .Y(new_n4850_));
  NOR2  g04465(.A(new_n4850_), .B(new_n1303_), .Y(new_n4851_));
  NOR2  g04466(.A(new_n4851_), .B(new_n1307_), .Y(new_n4852_));
  NOR2  g04467(.A(new_n4852_), .B(new_n1311_), .Y(new_n4853_));
  NOR2  g04468(.A(new_n4853_), .B(new_n1315_), .Y(new_n4854_));
  NOR2  g04469(.A(new_n4854_), .B(new_n1319_), .Y(new_n4855_));
  NOR2  g04470(.A(new_n4855_), .B(new_n1323_), .Y(new_n4856_));
  NOR2  g04471(.A(new_n4856_), .B(new_n1327_), .Y(new_n4857_));
  NOR2  g04472(.A(new_n4857_), .B(new_n1331_), .Y(new_n4858_));
  NOR2  g04473(.A(new_n4858_), .B(new_n1335_), .Y(new_n4859_));
  NOR2  g04474(.A(new_n4859_), .B(new_n1339_), .Y(new_n4860_));
  NOR2  g04475(.A(new_n4860_), .B(new_n1343_), .Y(new_n4861_));
  NOR2  g04476(.A(new_n4861_), .B(new_n1347_), .Y(new_n4862_));
  NOR2  g04477(.A(new_n4862_), .B(new_n1351_), .Y(new_n4863_));
  NOR2  g04478(.A(new_n4863_), .B(new_n1355_), .Y(new_n4864_));
  NOR2  g04479(.A(new_n4864_), .B(new_n1359_), .Y(new_n4865_));
  NOR2  g04480(.A(new_n4865_), .B(new_n1363_), .Y(new_n4866_));
  NOR2  g04481(.A(new_n4866_), .B(new_n1367_), .Y(new_n4867_));
  NOR2  g04482(.A(new_n4867_), .B(new_n1371_), .Y(new_n4868_));
  NOR2  g04483(.A(new_n4868_), .B(new_n1375_), .Y(new_n4869_));
  NOR2  g04484(.A(new_n4869_), .B(new_n1379_), .Y(new_n4870_));
  NOR2  g04485(.A(new_n4870_), .B(new_n1383_), .Y(new_n4871_));
  NOR2  g04486(.A(new_n4871_), .B(new_n1387_), .Y(new_n4872_));
  NOR2  g04487(.A(new_n4872_), .B(new_n1391_), .Y(new_n4873_));
  NOR2  g04488(.A(new_n4873_), .B(new_n1395_), .Y(new_n4874_));
  NOR2  g04489(.A(new_n4874_), .B(new_n1399_), .Y(new_n4875_));
  NOR2  g04490(.A(new_n4875_), .B(new_n1403_), .Y(new_n4876_));
  NOR2  g04491(.A(new_n4876_), .B(new_n1407_), .Y(new_n4877_));
  NOR2  g04492(.A(new_n4877_), .B(new_n1411_), .Y(new_n4878_));
  NOR2  g04493(.A(new_n4878_), .B(new_n1415_), .Y(new_n4879_));
  NOR2  g04494(.A(new_n4879_), .B(new_n1419_), .Y(new_n4880_));
  NOR2  g04495(.A(new_n4880_), .B(new_n1423_), .Y(new_n4881_));
  NOR2  g04496(.A(new_n4881_), .B(new_n1427_), .Y(new_n4882_));
  NOR2  g04497(.A(new_n4882_), .B(new_n1431_), .Y(new_n4883_));
  NOR2  g04498(.A(new_n4883_), .B(new_n1435_), .Y(new_n4884_));
  NOR2  g04499(.A(new_n4884_), .B(new_n1439_), .Y(new_n4885_));
  NOR2  g04500(.A(new_n4885_), .B(new_n1443_), .Y(new_n4886_));
  NOR2  g04501(.A(new_n4886_), .B(new_n1447_), .Y(new_n4887_));
  NOR2  g04502(.A(new_n4887_), .B(new_n1451_), .Y(new_n4888_));
  NOR2  g04503(.A(new_n4888_), .B(new_n1455_), .Y(new_n4889_));
  NOR2  g04504(.A(new_n4889_), .B(new_n1459_), .Y(new_n4890_));
  NOR2  g04505(.A(new_n4890_), .B(new_n1463_), .Y(new_n4891_));
  NOR2  g04506(.A(new_n4891_), .B(new_n1467_), .Y(new_n4892_));
  NOR2  g04507(.A(new_n4892_), .B(new_n1471_), .Y(new_n4893_));
  NOR2  g04508(.A(new_n4893_), .B(new_n1475_), .Y(new_n4894_));
  NOR2  g04509(.A(new_n4894_), .B(new_n1479_), .Y(new_n4895_));
  NOR2  g04510(.A(new_n4895_), .B(new_n1483_), .Y(new_n4896_));
  NOR2  g04511(.A(new_n4896_), .B(new_n1487_), .Y(new_n4897_));
  NOR2  g04512(.A(new_n4897_), .B(new_n1491_), .Y(new_n4898_));
  NOR2  g04513(.A(new_n4898_), .B(new_n1495_), .Y(new_n4899_));
  NOR2  g04514(.A(new_n4899_), .B(new_n1499_), .Y(new_n4900_));
  NOR2  g04515(.A(new_n4900_), .B(new_n1503_), .Y(new_n4901_));
  NOR2  g04516(.A(new_n4901_), .B(new_n1507_), .Y(new_n4902_));
  NOR2  g04517(.A(new_n4902_), .B(new_n1511_), .Y(new_n4903_));
  NOR2  g04518(.A(new_n4903_), .B(new_n1515_), .Y(new_n4904_));
  NOR2  g04519(.A(new_n4904_), .B(new_n1519_), .Y(new_n4905_));
  NOR2  g04520(.A(new_n4905_), .B(new_n1523_), .Y(new_n4906_));
  NOR2  g04521(.A(new_n4906_), .B(new_n1527_), .Y(new_n4907_));
  NOR2  g04522(.A(new_n4907_), .B(new_n1797_), .Y(new_n4908_));
  NOR2  g04523(.A(new_n4908_), .B(new_n396_), .Y(new_n4909_));
  NOR2  g04524(.A(new_n4909_), .B(new_n400_), .Y(new_n4910_));
  NOR2  g04525(.A(new_n4910_), .B(new_n406_), .Y(new_n4911_));
  NOR2  g04526(.A(new_n4911_), .B(new_n410_), .Y(new_n4912_));
  NOR2  g04527(.A(new_n4912_), .B(new_n416_), .Y(new_n4913_));
  NOR2  g04528(.A(new_n4913_), .B(new_n420_), .Y(new_n4914_));
  NOR2  g04529(.A(new_n4914_), .B(new_n426_), .Y(new_n4915_));
  NOR2  g04530(.A(new_n4915_), .B(new_n430_), .Y(new_n4916_));
  NOR2  g04531(.A(new_n4916_), .B(new_n436_), .Y(new_n4917_));
  NOR2  g04532(.A(new_n4917_), .B(new_n440_), .Y(new_n4918_));
  NOR2  g04533(.A(new_n4918_), .B(new_n446_), .Y(new_n4919_));
  NOR2  g04534(.A(new_n4919_), .B(new_n450_), .Y(new_n4920_));
  NOR2  g04535(.A(new_n4920_), .B(new_n456_), .Y(new_n4921_));
  NOR2  g04536(.A(new_n4921_), .B(new_n460_), .Y(new_n4922_));
  NOR2  g04537(.A(new_n4922_), .B(new_n466_), .Y(new_n4923_));
  NOR2  g04538(.A(new_n4923_), .B(new_n470_), .Y(new_n4924_));
  NOR2  g04539(.A(new_n4924_), .B(new_n476_), .Y(new_n4925_));
  NOR2  g04540(.A(new_n4925_), .B(new_n480_), .Y(new_n4926_));
  NOR2  g04541(.A(new_n4926_), .B(new_n486_), .Y(new_n4927_));
  NOR2  g04542(.A(new_n4927_), .B(new_n490_), .Y(new_n4928_));
  NOR2  g04543(.A(new_n4928_), .B(new_n496_), .Y(new_n4929_));
  NOR2  g04544(.A(new_n4929_), .B(new_n500_), .Y(new_n4930_));
  NOR2  g04545(.A(new_n4930_), .B(new_n506_), .Y(new_n4931_));
  NOR2  g04546(.A(new_n4931_), .B(new_n510_), .Y(new_n4932_));
  NOR2  g04547(.A(new_n4932_), .B(new_n516_), .Y(new_n4933_));
  NAND2 g04548(.A(new_n518_), .B(\req[41] ), .Y(new_n4934_));
  NOR2  g04549(.A(new_n4934_), .B(new_n4933_), .Y(\grant[41] ));
  INV   g04550(.A(new_n529_), .Y(new_n4936_));
  NOR2  g04551(.A(new_n936_), .B(new_n4936_), .Y(new_n4937_));
  NOR2  g04552(.A(new_n4937_), .B(new_n536_), .Y(new_n4938_));
  NOR2  g04553(.A(new_n4938_), .B(new_n540_), .Y(new_n4939_));
  NOR2  g04554(.A(new_n4939_), .B(new_n546_), .Y(new_n4940_));
  NOR2  g04555(.A(new_n4940_), .B(new_n550_), .Y(new_n4941_));
  NOR2  g04556(.A(new_n4941_), .B(new_n556_), .Y(new_n4942_));
  NOR2  g04557(.A(new_n4942_), .B(new_n560_), .Y(new_n4943_));
  NOR2  g04558(.A(new_n4943_), .B(new_n566_), .Y(new_n4944_));
  NOR2  g04559(.A(new_n4944_), .B(new_n570_), .Y(new_n4945_));
  NOR2  g04560(.A(new_n4945_), .B(new_n576_), .Y(new_n4946_));
  NOR2  g04561(.A(new_n4946_), .B(new_n580_), .Y(new_n4947_));
  NOR2  g04562(.A(new_n4947_), .B(new_n586_), .Y(new_n4948_));
  NOR2  g04563(.A(new_n4948_), .B(new_n590_), .Y(new_n4949_));
  NOR2  g04564(.A(new_n4949_), .B(new_n596_), .Y(new_n4950_));
  NOR2  g04565(.A(new_n4950_), .B(new_n600_), .Y(new_n4951_));
  NOR2  g04566(.A(new_n4951_), .B(new_n606_), .Y(new_n4952_));
  NOR2  g04567(.A(new_n4952_), .B(new_n610_), .Y(new_n4953_));
  NOR2  g04568(.A(new_n4953_), .B(new_n616_), .Y(new_n4954_));
  NOR2  g04569(.A(new_n4954_), .B(new_n620_), .Y(new_n4955_));
  NOR2  g04570(.A(new_n4955_), .B(new_n626_), .Y(new_n4956_));
  NOR2  g04571(.A(new_n4956_), .B(new_n630_), .Y(new_n4957_));
  NOR2  g04572(.A(new_n4957_), .B(new_n636_), .Y(new_n4958_));
  NOR2  g04573(.A(new_n4958_), .B(new_n640_), .Y(new_n4959_));
  NOR2  g04574(.A(new_n4959_), .B(new_n646_), .Y(new_n4960_));
  NOR2  g04575(.A(new_n4960_), .B(new_n650_), .Y(new_n4961_));
  NOR2  g04576(.A(new_n4961_), .B(new_n656_), .Y(new_n4962_));
  NOR2  g04577(.A(new_n4962_), .B(new_n660_), .Y(new_n4963_));
  NOR2  g04578(.A(new_n4963_), .B(new_n666_), .Y(new_n4964_));
  NOR2  g04579(.A(new_n4964_), .B(new_n670_), .Y(new_n4965_));
  NOR2  g04580(.A(new_n4965_), .B(new_n676_), .Y(new_n4966_));
  NOR2  g04581(.A(new_n4966_), .B(new_n680_), .Y(new_n4967_));
  NOR2  g04582(.A(new_n4967_), .B(new_n686_), .Y(new_n4968_));
  NOR2  g04583(.A(new_n4968_), .B(new_n690_), .Y(new_n4969_));
  NOR2  g04584(.A(new_n4969_), .B(new_n696_), .Y(new_n4970_));
  NOR2  g04585(.A(new_n4970_), .B(new_n700_), .Y(new_n4971_));
  NOR2  g04586(.A(new_n4971_), .B(new_n706_), .Y(new_n4972_));
  NOR2  g04587(.A(new_n4972_), .B(new_n710_), .Y(new_n4973_));
  NOR2  g04588(.A(new_n4973_), .B(new_n716_), .Y(new_n4974_));
  NOR2  g04589(.A(new_n4974_), .B(new_n720_), .Y(new_n4975_));
  NOR2  g04590(.A(new_n4975_), .B(new_n726_), .Y(new_n4976_));
  NOR2  g04591(.A(new_n4976_), .B(new_n730_), .Y(new_n4977_));
  NOR2  g04592(.A(new_n4977_), .B(new_n736_), .Y(new_n4978_));
  NOR2  g04593(.A(new_n4978_), .B(new_n740_), .Y(new_n4979_));
  NOR2  g04594(.A(new_n4979_), .B(new_n746_), .Y(new_n4980_));
  NOR2  g04595(.A(new_n4980_), .B(new_n750_), .Y(new_n4981_));
  NOR2  g04596(.A(new_n4981_), .B(new_n756_), .Y(new_n4982_));
  NOR2  g04597(.A(new_n4982_), .B(new_n760_), .Y(new_n4983_));
  NOR2  g04598(.A(new_n4983_), .B(new_n766_), .Y(new_n4984_));
  NOR2  g04599(.A(new_n4984_), .B(new_n770_), .Y(new_n4985_));
  NOR2  g04600(.A(new_n4985_), .B(new_n776_), .Y(new_n4986_));
  NOR2  g04601(.A(new_n4986_), .B(new_n780_), .Y(new_n4987_));
  NOR2  g04602(.A(new_n4987_), .B(new_n786_), .Y(new_n4988_));
  NOR2  g04603(.A(new_n4988_), .B(new_n790_), .Y(new_n4989_));
  NOR2  g04604(.A(new_n4989_), .B(new_n796_), .Y(new_n4990_));
  NOR2  g04605(.A(new_n4990_), .B(new_n800_), .Y(new_n4991_));
  NOR2  g04606(.A(new_n4991_), .B(new_n806_), .Y(new_n4992_));
  NOR2  g04607(.A(new_n4992_), .B(new_n1616_), .Y(new_n4993_));
  NOR2  g04608(.A(new_n4993_), .B(new_n1618_), .Y(new_n4994_));
  NOR2  g04609(.A(new_n4994_), .B(new_n1885_), .Y(new_n4995_));
  NOR2  g04610(.A(new_n4995_), .B(new_n820_), .Y(new_n4996_));
  NOR2  g04611(.A(new_n4996_), .B(new_n824_), .Y(new_n4997_));
  NOR2  g04612(.A(new_n4997_), .B(new_n829_), .Y(new_n4998_));
  NOR2  g04613(.A(new_n4998_), .B(new_n833_), .Y(new_n4999_));
  NOR2  g04614(.A(new_n4999_), .B(new_n838_), .Y(new_n5000_));
  NOR2  g04615(.A(new_n5000_), .B(new_n842_), .Y(new_n5001_));
  NOR2  g04616(.A(new_n5001_), .B(new_n847_), .Y(new_n5002_));
  NOR2  g04617(.A(new_n5002_), .B(new_n851_), .Y(new_n5003_));
  NOR2  g04618(.A(new_n5003_), .B(new_n856_), .Y(new_n5004_));
  NOR2  g04619(.A(new_n5004_), .B(new_n860_), .Y(new_n5005_));
  NOR2  g04620(.A(new_n5005_), .B(new_n865_), .Y(new_n5006_));
  NOR2  g04621(.A(new_n5006_), .B(new_n869_), .Y(new_n5007_));
  NOR2  g04622(.A(new_n5007_), .B(new_n874_), .Y(new_n5008_));
  NOR2  g04623(.A(new_n5008_), .B(new_n878_), .Y(new_n5009_));
  NOR2  g04624(.A(new_n5009_), .B(new_n883_), .Y(new_n5010_));
  NOR2  g04625(.A(new_n5010_), .B(new_n887_), .Y(new_n5011_));
  NOR2  g04626(.A(new_n5011_), .B(new_n892_), .Y(new_n5012_));
  NOR2  g04627(.A(new_n5012_), .B(new_n896_), .Y(new_n5013_));
  NOR2  g04628(.A(new_n5013_), .B(new_n901_), .Y(new_n5014_));
  NOR2  g04629(.A(new_n5014_), .B(new_n905_), .Y(new_n5015_));
  NOR2  g04630(.A(new_n5015_), .B(new_n910_), .Y(new_n5016_));
  NOR2  g04631(.A(new_n5016_), .B(new_n914_), .Y(new_n5017_));
  NOR2  g04632(.A(new_n5017_), .B(new_n919_), .Y(new_n5018_));
  NOR2  g04633(.A(new_n5018_), .B(new_n923_), .Y(new_n5019_));
  NOR2  g04634(.A(new_n5019_), .B(new_n928_), .Y(new_n5020_));
  NAND2 g04635(.A(new_n930_), .B(\req[42] ), .Y(new_n5021_));
  NOR2  g04636(.A(new_n5021_), .B(new_n5020_), .Y(\grant[42] ));
  INV   g04637(.A(new_n940_), .Y(new_n5023_));
  NOR2  g04638(.A(new_n1302_), .B(new_n5023_), .Y(new_n5024_));
  NOR2  g04639(.A(new_n5024_), .B(new_n946_), .Y(new_n5025_));
  NOR2  g04640(.A(new_n5025_), .B(new_n950_), .Y(new_n5026_));
  NOR2  g04641(.A(new_n5026_), .B(new_n955_), .Y(new_n5027_));
  NOR2  g04642(.A(new_n5027_), .B(new_n959_), .Y(new_n5028_));
  NOR2  g04643(.A(new_n5028_), .B(new_n964_), .Y(new_n5029_));
  NOR2  g04644(.A(new_n5029_), .B(new_n968_), .Y(new_n5030_));
  NOR2  g04645(.A(new_n5030_), .B(new_n973_), .Y(new_n5031_));
  NOR2  g04646(.A(new_n5031_), .B(new_n977_), .Y(new_n5032_));
  NOR2  g04647(.A(new_n5032_), .B(new_n982_), .Y(new_n5033_));
  NOR2  g04648(.A(new_n5033_), .B(new_n986_), .Y(new_n5034_));
  NOR2  g04649(.A(new_n5034_), .B(new_n991_), .Y(new_n5035_));
  NOR2  g04650(.A(new_n5035_), .B(new_n995_), .Y(new_n5036_));
  NOR2  g04651(.A(new_n5036_), .B(new_n1000_), .Y(new_n5037_));
  NOR2  g04652(.A(new_n5037_), .B(new_n1004_), .Y(new_n5038_));
  NOR2  g04653(.A(new_n5038_), .B(new_n1009_), .Y(new_n5039_));
  NOR2  g04654(.A(new_n5039_), .B(new_n1013_), .Y(new_n5040_));
  NOR2  g04655(.A(new_n5040_), .B(new_n1018_), .Y(new_n5041_));
  NOR2  g04656(.A(new_n5041_), .B(new_n1022_), .Y(new_n5042_));
  NOR2  g04657(.A(new_n5042_), .B(new_n1027_), .Y(new_n5043_));
  NOR2  g04658(.A(new_n5043_), .B(new_n1031_), .Y(new_n5044_));
  NOR2  g04659(.A(new_n5044_), .B(new_n1036_), .Y(new_n5045_));
  NOR2  g04660(.A(new_n5045_), .B(new_n1040_), .Y(new_n5046_));
  NOR2  g04661(.A(new_n5046_), .B(new_n1045_), .Y(new_n5047_));
  NOR2  g04662(.A(new_n5047_), .B(new_n1049_), .Y(new_n5048_));
  NOR2  g04663(.A(new_n5048_), .B(new_n1054_), .Y(new_n5049_));
  NOR2  g04664(.A(new_n5049_), .B(new_n1058_), .Y(new_n5050_));
  NOR2  g04665(.A(new_n5050_), .B(new_n1063_), .Y(new_n5051_));
  NOR2  g04666(.A(new_n5051_), .B(new_n1067_), .Y(new_n5052_));
  NOR2  g04667(.A(new_n5052_), .B(new_n1072_), .Y(new_n5053_));
  NOR2  g04668(.A(new_n5053_), .B(new_n1076_), .Y(new_n5054_));
  NOR2  g04669(.A(new_n5054_), .B(new_n1081_), .Y(new_n5055_));
  NOR2  g04670(.A(new_n5055_), .B(new_n1085_), .Y(new_n5056_));
  NOR2  g04671(.A(new_n5056_), .B(new_n1090_), .Y(new_n5057_));
  NOR2  g04672(.A(new_n5057_), .B(new_n1094_), .Y(new_n5058_));
  NOR2  g04673(.A(new_n5058_), .B(new_n1099_), .Y(new_n5059_));
  NOR2  g04674(.A(new_n5059_), .B(new_n1103_), .Y(new_n5060_));
  NOR2  g04675(.A(new_n5060_), .B(new_n1108_), .Y(new_n5061_));
  NOR2  g04676(.A(new_n5061_), .B(new_n1112_), .Y(new_n5062_));
  NOR2  g04677(.A(new_n5062_), .B(new_n1117_), .Y(new_n5063_));
  NOR2  g04678(.A(new_n5063_), .B(new_n1121_), .Y(new_n5064_));
  NOR2  g04679(.A(new_n5064_), .B(new_n1126_), .Y(new_n5065_));
  NOR2  g04680(.A(new_n5065_), .B(new_n1130_), .Y(new_n5066_));
  NOR2  g04681(.A(new_n5066_), .B(new_n1135_), .Y(new_n5067_));
  NOR2  g04682(.A(new_n5067_), .B(new_n1139_), .Y(new_n5068_));
  NOR2  g04683(.A(new_n5068_), .B(new_n1144_), .Y(new_n5069_));
  NOR2  g04684(.A(new_n5069_), .B(new_n1148_), .Y(new_n5070_));
  NOR2  g04685(.A(new_n5070_), .B(new_n1153_), .Y(new_n5071_));
  NOR2  g04686(.A(new_n5071_), .B(new_n1157_), .Y(new_n5072_));
  NOR2  g04687(.A(new_n5072_), .B(new_n1162_), .Y(new_n5073_));
  NOR2  g04688(.A(new_n5073_), .B(new_n1166_), .Y(new_n5074_));
  NOR2  g04689(.A(new_n5074_), .B(new_n1171_), .Y(new_n5075_));
  NOR2  g04690(.A(new_n5075_), .B(new_n1175_), .Y(new_n5076_));
  NOR2  g04691(.A(new_n5076_), .B(new_n1180_), .Y(new_n5077_));
  NOR2  g04692(.A(new_n5077_), .B(new_n1184_), .Y(new_n5078_));
  NOR2  g04693(.A(new_n5078_), .B(new_n1189_), .Y(new_n5079_));
  NOR2  g04694(.A(new_n5079_), .B(new_n1707_), .Y(new_n5080_));
  NOR2  g04695(.A(new_n5080_), .B(new_n1709_), .Y(new_n5081_));
  NOR2  g04696(.A(new_n5081_), .B(new_n1973_), .Y(new_n5082_));
  NOR2  g04697(.A(new_n5082_), .B(new_n1199_), .Y(new_n5083_));
  NOR2  g04698(.A(new_n5083_), .B(new_n1203_), .Y(new_n5084_));
  NOR2  g04699(.A(new_n5084_), .B(new_n1207_), .Y(new_n5085_));
  NOR2  g04700(.A(new_n5085_), .B(new_n1211_), .Y(new_n5086_));
  NOR2  g04701(.A(new_n5086_), .B(new_n1215_), .Y(new_n5087_));
  NOR2  g04702(.A(new_n5087_), .B(new_n1219_), .Y(new_n5088_));
  NOR2  g04703(.A(new_n5088_), .B(new_n1223_), .Y(new_n5089_));
  NOR2  g04704(.A(new_n5089_), .B(new_n1227_), .Y(new_n5090_));
  NOR2  g04705(.A(new_n5090_), .B(new_n1231_), .Y(new_n5091_));
  NOR2  g04706(.A(new_n5091_), .B(new_n1235_), .Y(new_n5092_));
  NOR2  g04707(.A(new_n5092_), .B(new_n1239_), .Y(new_n5093_));
  NOR2  g04708(.A(new_n5093_), .B(new_n1243_), .Y(new_n5094_));
  NOR2  g04709(.A(new_n5094_), .B(new_n1247_), .Y(new_n5095_));
  NOR2  g04710(.A(new_n5095_), .B(new_n1251_), .Y(new_n5096_));
  NOR2  g04711(.A(new_n5096_), .B(new_n1255_), .Y(new_n5097_));
  NOR2  g04712(.A(new_n5097_), .B(new_n1259_), .Y(new_n5098_));
  NOR2  g04713(.A(new_n5098_), .B(new_n1263_), .Y(new_n5099_));
  NOR2  g04714(.A(new_n5099_), .B(new_n1267_), .Y(new_n5100_));
  NOR2  g04715(.A(new_n5100_), .B(new_n1271_), .Y(new_n5101_));
  NOR2  g04716(.A(new_n5101_), .B(new_n1275_), .Y(new_n5102_));
  NOR2  g04717(.A(new_n5102_), .B(new_n1279_), .Y(new_n5103_));
  NOR2  g04718(.A(new_n5103_), .B(new_n1283_), .Y(new_n5104_));
  NOR2  g04719(.A(new_n5104_), .B(new_n1287_), .Y(new_n5105_));
  NOR2  g04720(.A(new_n5105_), .B(new_n1291_), .Y(new_n5106_));
  NOR2  g04721(.A(new_n5106_), .B(new_n1295_), .Y(new_n5107_));
  NAND2 g04722(.A(new_n1297_), .B(\req[43] ), .Y(new_n5108_));
  NOR2  g04723(.A(new_n5108_), .B(new_n5107_), .Y(\grant[43] ));
  INV   g04724(.A(new_n1306_), .Y(new_n5110_));
  NOR2  g04725(.A(new_n5110_), .B(new_n535_), .Y(new_n5111_));
  NOR2  g04726(.A(new_n5111_), .B(new_n1311_), .Y(new_n5112_));
  NOR2  g04727(.A(new_n5112_), .B(new_n1315_), .Y(new_n5113_));
  NOR2  g04728(.A(new_n5113_), .B(new_n1319_), .Y(new_n5114_));
  NOR2  g04729(.A(new_n5114_), .B(new_n1323_), .Y(new_n5115_));
  NOR2  g04730(.A(new_n5115_), .B(new_n1327_), .Y(new_n5116_));
  NOR2  g04731(.A(new_n5116_), .B(new_n1331_), .Y(new_n5117_));
  NOR2  g04732(.A(new_n5117_), .B(new_n1335_), .Y(new_n5118_));
  NOR2  g04733(.A(new_n5118_), .B(new_n1339_), .Y(new_n5119_));
  NOR2  g04734(.A(new_n5119_), .B(new_n1343_), .Y(new_n5120_));
  NOR2  g04735(.A(new_n5120_), .B(new_n1347_), .Y(new_n5121_));
  NOR2  g04736(.A(new_n5121_), .B(new_n1351_), .Y(new_n5122_));
  NOR2  g04737(.A(new_n5122_), .B(new_n1355_), .Y(new_n5123_));
  NOR2  g04738(.A(new_n5123_), .B(new_n1359_), .Y(new_n5124_));
  NOR2  g04739(.A(new_n5124_), .B(new_n1363_), .Y(new_n5125_));
  NOR2  g04740(.A(new_n5125_), .B(new_n1367_), .Y(new_n5126_));
  NOR2  g04741(.A(new_n5126_), .B(new_n1371_), .Y(new_n5127_));
  NOR2  g04742(.A(new_n5127_), .B(new_n1375_), .Y(new_n5128_));
  NOR2  g04743(.A(new_n5128_), .B(new_n1379_), .Y(new_n5129_));
  NOR2  g04744(.A(new_n5129_), .B(new_n1383_), .Y(new_n5130_));
  NOR2  g04745(.A(new_n5130_), .B(new_n1387_), .Y(new_n5131_));
  NOR2  g04746(.A(new_n5131_), .B(new_n1391_), .Y(new_n5132_));
  NOR2  g04747(.A(new_n5132_), .B(new_n1395_), .Y(new_n5133_));
  NOR2  g04748(.A(new_n5133_), .B(new_n1399_), .Y(new_n5134_));
  NOR2  g04749(.A(new_n5134_), .B(new_n1403_), .Y(new_n5135_));
  NOR2  g04750(.A(new_n5135_), .B(new_n1407_), .Y(new_n5136_));
  NOR2  g04751(.A(new_n5136_), .B(new_n1411_), .Y(new_n5137_));
  NOR2  g04752(.A(new_n5137_), .B(new_n1415_), .Y(new_n5138_));
  NOR2  g04753(.A(new_n5138_), .B(new_n1419_), .Y(new_n5139_));
  NOR2  g04754(.A(new_n5139_), .B(new_n1423_), .Y(new_n5140_));
  NOR2  g04755(.A(new_n5140_), .B(new_n1427_), .Y(new_n5141_));
  NOR2  g04756(.A(new_n5141_), .B(new_n1431_), .Y(new_n5142_));
  NOR2  g04757(.A(new_n5142_), .B(new_n1435_), .Y(new_n5143_));
  NOR2  g04758(.A(new_n5143_), .B(new_n1439_), .Y(new_n5144_));
  NOR2  g04759(.A(new_n5144_), .B(new_n1443_), .Y(new_n5145_));
  NOR2  g04760(.A(new_n5145_), .B(new_n1447_), .Y(new_n5146_));
  NOR2  g04761(.A(new_n5146_), .B(new_n1451_), .Y(new_n5147_));
  NOR2  g04762(.A(new_n5147_), .B(new_n1455_), .Y(new_n5148_));
  NOR2  g04763(.A(new_n5148_), .B(new_n1459_), .Y(new_n5149_));
  NOR2  g04764(.A(new_n5149_), .B(new_n1463_), .Y(new_n5150_));
  NOR2  g04765(.A(new_n5150_), .B(new_n1467_), .Y(new_n5151_));
  NOR2  g04766(.A(new_n5151_), .B(new_n1471_), .Y(new_n5152_));
  NOR2  g04767(.A(new_n5152_), .B(new_n1475_), .Y(new_n5153_));
  NOR2  g04768(.A(new_n5153_), .B(new_n1479_), .Y(new_n5154_));
  NOR2  g04769(.A(new_n5154_), .B(new_n1483_), .Y(new_n5155_));
  NOR2  g04770(.A(new_n5155_), .B(new_n1487_), .Y(new_n5156_));
  NOR2  g04771(.A(new_n5156_), .B(new_n1491_), .Y(new_n5157_));
  NOR2  g04772(.A(new_n5157_), .B(new_n1495_), .Y(new_n5158_));
  NOR2  g04773(.A(new_n5158_), .B(new_n1499_), .Y(new_n5159_));
  NOR2  g04774(.A(new_n5159_), .B(new_n1503_), .Y(new_n5160_));
  NOR2  g04775(.A(new_n5160_), .B(new_n1507_), .Y(new_n5161_));
  NOR2  g04776(.A(new_n5161_), .B(new_n1511_), .Y(new_n5162_));
  NOR2  g04777(.A(new_n5162_), .B(new_n1515_), .Y(new_n5163_));
  NOR2  g04778(.A(new_n5163_), .B(new_n1519_), .Y(new_n5164_));
  NOR2  g04779(.A(new_n5164_), .B(new_n1523_), .Y(new_n5165_));
  NOR2  g04780(.A(new_n5165_), .B(new_n1527_), .Y(new_n5166_));
  NOR2  g04781(.A(new_n5166_), .B(new_n1797_), .Y(new_n5167_));
  NOR2  g04782(.A(new_n5167_), .B(new_n396_), .Y(new_n5168_));
  NOR2  g04783(.A(new_n5168_), .B(new_n400_), .Y(new_n5169_));
  NOR2  g04784(.A(new_n5169_), .B(new_n406_), .Y(new_n5170_));
  NOR2  g04785(.A(new_n5170_), .B(new_n410_), .Y(new_n5171_));
  NOR2  g04786(.A(new_n5171_), .B(new_n416_), .Y(new_n5172_));
  NOR2  g04787(.A(new_n5172_), .B(new_n420_), .Y(new_n5173_));
  NOR2  g04788(.A(new_n5173_), .B(new_n426_), .Y(new_n5174_));
  NOR2  g04789(.A(new_n5174_), .B(new_n430_), .Y(new_n5175_));
  NOR2  g04790(.A(new_n5175_), .B(new_n436_), .Y(new_n5176_));
  NOR2  g04791(.A(new_n5176_), .B(new_n440_), .Y(new_n5177_));
  NOR2  g04792(.A(new_n5177_), .B(new_n446_), .Y(new_n5178_));
  NOR2  g04793(.A(new_n5178_), .B(new_n450_), .Y(new_n5179_));
  NOR2  g04794(.A(new_n5179_), .B(new_n456_), .Y(new_n5180_));
  NOR2  g04795(.A(new_n5180_), .B(new_n460_), .Y(new_n5181_));
  NOR2  g04796(.A(new_n5181_), .B(new_n466_), .Y(new_n5182_));
  NOR2  g04797(.A(new_n5182_), .B(new_n470_), .Y(new_n5183_));
  NOR2  g04798(.A(new_n5183_), .B(new_n476_), .Y(new_n5184_));
  NOR2  g04799(.A(new_n5184_), .B(new_n480_), .Y(new_n5185_));
  NOR2  g04800(.A(new_n5185_), .B(new_n486_), .Y(new_n5186_));
  NOR2  g04801(.A(new_n5186_), .B(new_n490_), .Y(new_n5187_));
  NOR2  g04802(.A(new_n5187_), .B(new_n496_), .Y(new_n5188_));
  NOR2  g04803(.A(new_n5188_), .B(new_n500_), .Y(new_n5189_));
  NOR2  g04804(.A(new_n5189_), .B(new_n506_), .Y(new_n5190_));
  NOR2  g04805(.A(new_n5190_), .B(new_n510_), .Y(new_n5191_));
  NOR2  g04806(.A(new_n5191_), .B(new_n516_), .Y(new_n5192_));
  NOR2  g04807(.A(new_n5192_), .B(new_n520_), .Y(new_n5193_));
  NOR2  g04808(.A(new_n5193_), .B(new_n526_), .Y(new_n5194_));
  NAND2 g04809(.A(new_n528_), .B(\req[44] ), .Y(new_n5195_));
  NOR2  g04810(.A(new_n5195_), .B(new_n5194_), .Y(\grant[44] ));
  INV   g04811(.A(new_n539_), .Y(new_n5197_));
  NOR2  g04812(.A(new_n945_), .B(new_n5197_), .Y(new_n5198_));
  NOR2  g04813(.A(new_n5198_), .B(new_n546_), .Y(new_n5199_));
  NOR2  g04814(.A(new_n5199_), .B(new_n550_), .Y(new_n5200_));
  NOR2  g04815(.A(new_n5200_), .B(new_n556_), .Y(new_n5201_));
  NOR2  g04816(.A(new_n5201_), .B(new_n560_), .Y(new_n5202_));
  NOR2  g04817(.A(new_n5202_), .B(new_n566_), .Y(new_n5203_));
  NOR2  g04818(.A(new_n5203_), .B(new_n570_), .Y(new_n5204_));
  NOR2  g04819(.A(new_n5204_), .B(new_n576_), .Y(new_n5205_));
  NOR2  g04820(.A(new_n5205_), .B(new_n580_), .Y(new_n5206_));
  NOR2  g04821(.A(new_n5206_), .B(new_n586_), .Y(new_n5207_));
  NOR2  g04822(.A(new_n5207_), .B(new_n590_), .Y(new_n5208_));
  NOR2  g04823(.A(new_n5208_), .B(new_n596_), .Y(new_n5209_));
  NOR2  g04824(.A(new_n5209_), .B(new_n600_), .Y(new_n5210_));
  NOR2  g04825(.A(new_n5210_), .B(new_n606_), .Y(new_n5211_));
  NOR2  g04826(.A(new_n5211_), .B(new_n610_), .Y(new_n5212_));
  NOR2  g04827(.A(new_n5212_), .B(new_n616_), .Y(new_n5213_));
  NOR2  g04828(.A(new_n5213_), .B(new_n620_), .Y(new_n5214_));
  NOR2  g04829(.A(new_n5214_), .B(new_n626_), .Y(new_n5215_));
  NOR2  g04830(.A(new_n5215_), .B(new_n630_), .Y(new_n5216_));
  NOR2  g04831(.A(new_n5216_), .B(new_n636_), .Y(new_n5217_));
  NOR2  g04832(.A(new_n5217_), .B(new_n640_), .Y(new_n5218_));
  NOR2  g04833(.A(new_n5218_), .B(new_n646_), .Y(new_n5219_));
  NOR2  g04834(.A(new_n5219_), .B(new_n650_), .Y(new_n5220_));
  NOR2  g04835(.A(new_n5220_), .B(new_n656_), .Y(new_n5221_));
  NOR2  g04836(.A(new_n5221_), .B(new_n660_), .Y(new_n5222_));
  NOR2  g04837(.A(new_n5222_), .B(new_n666_), .Y(new_n5223_));
  NOR2  g04838(.A(new_n5223_), .B(new_n670_), .Y(new_n5224_));
  NOR2  g04839(.A(new_n5224_), .B(new_n676_), .Y(new_n5225_));
  NOR2  g04840(.A(new_n5225_), .B(new_n680_), .Y(new_n5226_));
  NOR2  g04841(.A(new_n5226_), .B(new_n686_), .Y(new_n5227_));
  NOR2  g04842(.A(new_n5227_), .B(new_n690_), .Y(new_n5228_));
  NOR2  g04843(.A(new_n5228_), .B(new_n696_), .Y(new_n5229_));
  NOR2  g04844(.A(new_n5229_), .B(new_n700_), .Y(new_n5230_));
  NOR2  g04845(.A(new_n5230_), .B(new_n706_), .Y(new_n5231_));
  NOR2  g04846(.A(new_n5231_), .B(new_n710_), .Y(new_n5232_));
  NOR2  g04847(.A(new_n5232_), .B(new_n716_), .Y(new_n5233_));
  NOR2  g04848(.A(new_n5233_), .B(new_n720_), .Y(new_n5234_));
  NOR2  g04849(.A(new_n5234_), .B(new_n726_), .Y(new_n5235_));
  NOR2  g04850(.A(new_n5235_), .B(new_n730_), .Y(new_n5236_));
  NOR2  g04851(.A(new_n5236_), .B(new_n736_), .Y(new_n5237_));
  NOR2  g04852(.A(new_n5237_), .B(new_n740_), .Y(new_n5238_));
  NOR2  g04853(.A(new_n5238_), .B(new_n746_), .Y(new_n5239_));
  NOR2  g04854(.A(new_n5239_), .B(new_n750_), .Y(new_n5240_));
  NOR2  g04855(.A(new_n5240_), .B(new_n756_), .Y(new_n5241_));
  NOR2  g04856(.A(new_n5241_), .B(new_n760_), .Y(new_n5242_));
  NOR2  g04857(.A(new_n5242_), .B(new_n766_), .Y(new_n5243_));
  NOR2  g04858(.A(new_n5243_), .B(new_n770_), .Y(new_n5244_));
  NOR2  g04859(.A(new_n5244_), .B(new_n776_), .Y(new_n5245_));
  NOR2  g04860(.A(new_n5245_), .B(new_n780_), .Y(new_n5246_));
  NOR2  g04861(.A(new_n5246_), .B(new_n786_), .Y(new_n5247_));
  NOR2  g04862(.A(new_n5247_), .B(new_n790_), .Y(new_n5248_));
  NOR2  g04863(.A(new_n5248_), .B(new_n796_), .Y(new_n5249_));
  NOR2  g04864(.A(new_n5249_), .B(new_n800_), .Y(new_n5250_));
  NOR2  g04865(.A(new_n5250_), .B(new_n806_), .Y(new_n5251_));
  NOR2  g04866(.A(new_n5251_), .B(new_n1616_), .Y(new_n5252_));
  NOR2  g04867(.A(new_n5252_), .B(new_n1618_), .Y(new_n5253_));
  NOR2  g04868(.A(new_n5253_), .B(new_n1885_), .Y(new_n5254_));
  NOR2  g04869(.A(new_n5254_), .B(new_n820_), .Y(new_n5255_));
  NOR2  g04870(.A(new_n5255_), .B(new_n824_), .Y(new_n5256_));
  NOR2  g04871(.A(new_n5256_), .B(new_n829_), .Y(new_n5257_));
  NOR2  g04872(.A(new_n5257_), .B(new_n833_), .Y(new_n5258_));
  NOR2  g04873(.A(new_n5258_), .B(new_n838_), .Y(new_n5259_));
  NOR2  g04874(.A(new_n5259_), .B(new_n842_), .Y(new_n5260_));
  NOR2  g04875(.A(new_n5260_), .B(new_n847_), .Y(new_n5261_));
  NOR2  g04876(.A(new_n5261_), .B(new_n851_), .Y(new_n5262_));
  NOR2  g04877(.A(new_n5262_), .B(new_n856_), .Y(new_n5263_));
  NOR2  g04878(.A(new_n5263_), .B(new_n860_), .Y(new_n5264_));
  NOR2  g04879(.A(new_n5264_), .B(new_n865_), .Y(new_n5265_));
  NOR2  g04880(.A(new_n5265_), .B(new_n869_), .Y(new_n5266_));
  NOR2  g04881(.A(new_n5266_), .B(new_n874_), .Y(new_n5267_));
  NOR2  g04882(.A(new_n5267_), .B(new_n878_), .Y(new_n5268_));
  NOR2  g04883(.A(new_n5268_), .B(new_n883_), .Y(new_n5269_));
  NOR2  g04884(.A(new_n5269_), .B(new_n887_), .Y(new_n5270_));
  NOR2  g04885(.A(new_n5270_), .B(new_n892_), .Y(new_n5271_));
  NOR2  g04886(.A(new_n5271_), .B(new_n896_), .Y(new_n5272_));
  NOR2  g04887(.A(new_n5272_), .B(new_n901_), .Y(new_n5273_));
  NOR2  g04888(.A(new_n5273_), .B(new_n905_), .Y(new_n5274_));
  NOR2  g04889(.A(new_n5274_), .B(new_n910_), .Y(new_n5275_));
  NOR2  g04890(.A(new_n5275_), .B(new_n914_), .Y(new_n5276_));
  NOR2  g04891(.A(new_n5276_), .B(new_n919_), .Y(new_n5277_));
  NOR2  g04892(.A(new_n5277_), .B(new_n923_), .Y(new_n5278_));
  NOR2  g04893(.A(new_n5278_), .B(new_n928_), .Y(new_n5279_));
  NOR2  g04894(.A(new_n5279_), .B(new_n932_), .Y(new_n5280_));
  NOR2  g04895(.A(new_n5280_), .B(new_n937_), .Y(new_n5281_));
  NAND2 g04896(.A(new_n939_), .B(\req[45] ), .Y(new_n5282_));
  NOR2  g04897(.A(new_n5282_), .B(new_n5281_), .Y(\grant[45] ));
  INV   g04898(.A(new_n949_), .Y(new_n5284_));
  NOR2  g04899(.A(new_n1310_), .B(new_n5284_), .Y(new_n5285_));
  NOR2  g04900(.A(new_n5285_), .B(new_n955_), .Y(new_n5286_));
  NOR2  g04901(.A(new_n5286_), .B(new_n959_), .Y(new_n5287_));
  NOR2  g04902(.A(new_n5287_), .B(new_n964_), .Y(new_n5288_));
  NOR2  g04903(.A(new_n5288_), .B(new_n968_), .Y(new_n5289_));
  NOR2  g04904(.A(new_n5289_), .B(new_n973_), .Y(new_n5290_));
  NOR2  g04905(.A(new_n5290_), .B(new_n977_), .Y(new_n5291_));
  NOR2  g04906(.A(new_n5291_), .B(new_n982_), .Y(new_n5292_));
  NOR2  g04907(.A(new_n5292_), .B(new_n986_), .Y(new_n5293_));
  NOR2  g04908(.A(new_n5293_), .B(new_n991_), .Y(new_n5294_));
  NOR2  g04909(.A(new_n5294_), .B(new_n995_), .Y(new_n5295_));
  NOR2  g04910(.A(new_n5295_), .B(new_n1000_), .Y(new_n5296_));
  NOR2  g04911(.A(new_n5296_), .B(new_n1004_), .Y(new_n5297_));
  NOR2  g04912(.A(new_n5297_), .B(new_n1009_), .Y(new_n5298_));
  NOR2  g04913(.A(new_n5298_), .B(new_n1013_), .Y(new_n5299_));
  NOR2  g04914(.A(new_n5299_), .B(new_n1018_), .Y(new_n5300_));
  NOR2  g04915(.A(new_n5300_), .B(new_n1022_), .Y(new_n5301_));
  NOR2  g04916(.A(new_n5301_), .B(new_n1027_), .Y(new_n5302_));
  NOR2  g04917(.A(new_n5302_), .B(new_n1031_), .Y(new_n5303_));
  NOR2  g04918(.A(new_n5303_), .B(new_n1036_), .Y(new_n5304_));
  NOR2  g04919(.A(new_n5304_), .B(new_n1040_), .Y(new_n5305_));
  NOR2  g04920(.A(new_n5305_), .B(new_n1045_), .Y(new_n5306_));
  NOR2  g04921(.A(new_n5306_), .B(new_n1049_), .Y(new_n5307_));
  NOR2  g04922(.A(new_n5307_), .B(new_n1054_), .Y(new_n5308_));
  NOR2  g04923(.A(new_n5308_), .B(new_n1058_), .Y(new_n5309_));
  NOR2  g04924(.A(new_n5309_), .B(new_n1063_), .Y(new_n5310_));
  NOR2  g04925(.A(new_n5310_), .B(new_n1067_), .Y(new_n5311_));
  NOR2  g04926(.A(new_n5311_), .B(new_n1072_), .Y(new_n5312_));
  NOR2  g04927(.A(new_n5312_), .B(new_n1076_), .Y(new_n5313_));
  NOR2  g04928(.A(new_n5313_), .B(new_n1081_), .Y(new_n5314_));
  NOR2  g04929(.A(new_n5314_), .B(new_n1085_), .Y(new_n5315_));
  NOR2  g04930(.A(new_n5315_), .B(new_n1090_), .Y(new_n5316_));
  NOR2  g04931(.A(new_n5316_), .B(new_n1094_), .Y(new_n5317_));
  NOR2  g04932(.A(new_n5317_), .B(new_n1099_), .Y(new_n5318_));
  NOR2  g04933(.A(new_n5318_), .B(new_n1103_), .Y(new_n5319_));
  NOR2  g04934(.A(new_n5319_), .B(new_n1108_), .Y(new_n5320_));
  NOR2  g04935(.A(new_n5320_), .B(new_n1112_), .Y(new_n5321_));
  NOR2  g04936(.A(new_n5321_), .B(new_n1117_), .Y(new_n5322_));
  NOR2  g04937(.A(new_n5322_), .B(new_n1121_), .Y(new_n5323_));
  NOR2  g04938(.A(new_n5323_), .B(new_n1126_), .Y(new_n5324_));
  NOR2  g04939(.A(new_n5324_), .B(new_n1130_), .Y(new_n5325_));
  NOR2  g04940(.A(new_n5325_), .B(new_n1135_), .Y(new_n5326_));
  NOR2  g04941(.A(new_n5326_), .B(new_n1139_), .Y(new_n5327_));
  NOR2  g04942(.A(new_n5327_), .B(new_n1144_), .Y(new_n5328_));
  NOR2  g04943(.A(new_n5328_), .B(new_n1148_), .Y(new_n5329_));
  NOR2  g04944(.A(new_n5329_), .B(new_n1153_), .Y(new_n5330_));
  NOR2  g04945(.A(new_n5330_), .B(new_n1157_), .Y(new_n5331_));
  NOR2  g04946(.A(new_n5331_), .B(new_n1162_), .Y(new_n5332_));
  NOR2  g04947(.A(new_n5332_), .B(new_n1166_), .Y(new_n5333_));
  NOR2  g04948(.A(new_n5333_), .B(new_n1171_), .Y(new_n5334_));
  NOR2  g04949(.A(new_n5334_), .B(new_n1175_), .Y(new_n5335_));
  NOR2  g04950(.A(new_n5335_), .B(new_n1180_), .Y(new_n5336_));
  NOR2  g04951(.A(new_n5336_), .B(new_n1184_), .Y(new_n5337_));
  NOR2  g04952(.A(new_n5337_), .B(new_n1189_), .Y(new_n5338_));
  NOR2  g04953(.A(new_n5338_), .B(new_n1707_), .Y(new_n5339_));
  NOR2  g04954(.A(new_n5339_), .B(new_n1709_), .Y(new_n5340_));
  NOR2  g04955(.A(new_n5340_), .B(new_n1973_), .Y(new_n5341_));
  NOR2  g04956(.A(new_n5341_), .B(new_n1199_), .Y(new_n5342_));
  NOR2  g04957(.A(new_n5342_), .B(new_n1203_), .Y(new_n5343_));
  NOR2  g04958(.A(new_n5343_), .B(new_n1207_), .Y(new_n5344_));
  NOR2  g04959(.A(new_n5344_), .B(new_n1211_), .Y(new_n5345_));
  NOR2  g04960(.A(new_n5345_), .B(new_n1215_), .Y(new_n5346_));
  NOR2  g04961(.A(new_n5346_), .B(new_n1219_), .Y(new_n5347_));
  NOR2  g04962(.A(new_n5347_), .B(new_n1223_), .Y(new_n5348_));
  NOR2  g04963(.A(new_n5348_), .B(new_n1227_), .Y(new_n5349_));
  NOR2  g04964(.A(new_n5349_), .B(new_n1231_), .Y(new_n5350_));
  NOR2  g04965(.A(new_n5350_), .B(new_n1235_), .Y(new_n5351_));
  NOR2  g04966(.A(new_n5351_), .B(new_n1239_), .Y(new_n5352_));
  NOR2  g04967(.A(new_n5352_), .B(new_n1243_), .Y(new_n5353_));
  NOR2  g04968(.A(new_n5353_), .B(new_n1247_), .Y(new_n5354_));
  NOR2  g04969(.A(new_n5354_), .B(new_n1251_), .Y(new_n5355_));
  NOR2  g04970(.A(new_n5355_), .B(new_n1255_), .Y(new_n5356_));
  NOR2  g04971(.A(new_n5356_), .B(new_n1259_), .Y(new_n5357_));
  NOR2  g04972(.A(new_n5357_), .B(new_n1263_), .Y(new_n5358_));
  NOR2  g04973(.A(new_n5358_), .B(new_n1267_), .Y(new_n5359_));
  NOR2  g04974(.A(new_n5359_), .B(new_n1271_), .Y(new_n5360_));
  NOR2  g04975(.A(new_n5360_), .B(new_n1275_), .Y(new_n5361_));
  NOR2  g04976(.A(new_n5361_), .B(new_n1279_), .Y(new_n5362_));
  NOR2  g04977(.A(new_n5362_), .B(new_n1283_), .Y(new_n5363_));
  NOR2  g04978(.A(new_n5363_), .B(new_n1287_), .Y(new_n5364_));
  NOR2  g04979(.A(new_n5364_), .B(new_n1291_), .Y(new_n5365_));
  NOR2  g04980(.A(new_n5365_), .B(new_n1295_), .Y(new_n5366_));
  NOR2  g04981(.A(new_n5366_), .B(new_n1299_), .Y(new_n5367_));
  NOR2  g04982(.A(new_n5367_), .B(new_n1303_), .Y(new_n5368_));
  NAND2 g04983(.A(new_n1305_), .B(\req[46] ), .Y(new_n5369_));
  NOR2  g04984(.A(new_n5369_), .B(new_n5368_), .Y(\grant[46] ));
  INV   g04985(.A(new_n1314_), .Y(new_n5371_));
  NOR2  g04986(.A(new_n5371_), .B(new_n545_), .Y(new_n5372_));
  NOR2  g04987(.A(new_n5372_), .B(new_n1319_), .Y(new_n5373_));
  NOR2  g04988(.A(new_n5373_), .B(new_n1323_), .Y(new_n5374_));
  NOR2  g04989(.A(new_n5374_), .B(new_n1327_), .Y(new_n5375_));
  NOR2  g04990(.A(new_n5375_), .B(new_n1331_), .Y(new_n5376_));
  NOR2  g04991(.A(new_n5376_), .B(new_n1335_), .Y(new_n5377_));
  NOR2  g04992(.A(new_n5377_), .B(new_n1339_), .Y(new_n5378_));
  NOR2  g04993(.A(new_n5378_), .B(new_n1343_), .Y(new_n5379_));
  NOR2  g04994(.A(new_n5379_), .B(new_n1347_), .Y(new_n5380_));
  NOR2  g04995(.A(new_n5380_), .B(new_n1351_), .Y(new_n5381_));
  NOR2  g04996(.A(new_n5381_), .B(new_n1355_), .Y(new_n5382_));
  NOR2  g04997(.A(new_n5382_), .B(new_n1359_), .Y(new_n5383_));
  NOR2  g04998(.A(new_n5383_), .B(new_n1363_), .Y(new_n5384_));
  NOR2  g04999(.A(new_n5384_), .B(new_n1367_), .Y(new_n5385_));
  NOR2  g05000(.A(new_n5385_), .B(new_n1371_), .Y(new_n5386_));
  NOR2  g05001(.A(new_n5386_), .B(new_n1375_), .Y(new_n5387_));
  NOR2  g05002(.A(new_n5387_), .B(new_n1379_), .Y(new_n5388_));
  NOR2  g05003(.A(new_n5388_), .B(new_n1383_), .Y(new_n5389_));
  NOR2  g05004(.A(new_n5389_), .B(new_n1387_), .Y(new_n5390_));
  NOR2  g05005(.A(new_n5390_), .B(new_n1391_), .Y(new_n5391_));
  NOR2  g05006(.A(new_n5391_), .B(new_n1395_), .Y(new_n5392_));
  NOR2  g05007(.A(new_n5392_), .B(new_n1399_), .Y(new_n5393_));
  NOR2  g05008(.A(new_n5393_), .B(new_n1403_), .Y(new_n5394_));
  NOR2  g05009(.A(new_n5394_), .B(new_n1407_), .Y(new_n5395_));
  NOR2  g05010(.A(new_n5395_), .B(new_n1411_), .Y(new_n5396_));
  NOR2  g05011(.A(new_n5396_), .B(new_n1415_), .Y(new_n5397_));
  NOR2  g05012(.A(new_n5397_), .B(new_n1419_), .Y(new_n5398_));
  NOR2  g05013(.A(new_n5398_), .B(new_n1423_), .Y(new_n5399_));
  NOR2  g05014(.A(new_n5399_), .B(new_n1427_), .Y(new_n5400_));
  NOR2  g05015(.A(new_n5400_), .B(new_n1431_), .Y(new_n5401_));
  NOR2  g05016(.A(new_n5401_), .B(new_n1435_), .Y(new_n5402_));
  NOR2  g05017(.A(new_n5402_), .B(new_n1439_), .Y(new_n5403_));
  NOR2  g05018(.A(new_n5403_), .B(new_n1443_), .Y(new_n5404_));
  NOR2  g05019(.A(new_n5404_), .B(new_n1447_), .Y(new_n5405_));
  NOR2  g05020(.A(new_n5405_), .B(new_n1451_), .Y(new_n5406_));
  NOR2  g05021(.A(new_n5406_), .B(new_n1455_), .Y(new_n5407_));
  NOR2  g05022(.A(new_n5407_), .B(new_n1459_), .Y(new_n5408_));
  NOR2  g05023(.A(new_n5408_), .B(new_n1463_), .Y(new_n5409_));
  NOR2  g05024(.A(new_n5409_), .B(new_n1467_), .Y(new_n5410_));
  NOR2  g05025(.A(new_n5410_), .B(new_n1471_), .Y(new_n5411_));
  NOR2  g05026(.A(new_n5411_), .B(new_n1475_), .Y(new_n5412_));
  NOR2  g05027(.A(new_n5412_), .B(new_n1479_), .Y(new_n5413_));
  NOR2  g05028(.A(new_n5413_), .B(new_n1483_), .Y(new_n5414_));
  NOR2  g05029(.A(new_n5414_), .B(new_n1487_), .Y(new_n5415_));
  NOR2  g05030(.A(new_n5415_), .B(new_n1491_), .Y(new_n5416_));
  NOR2  g05031(.A(new_n5416_), .B(new_n1495_), .Y(new_n5417_));
  NOR2  g05032(.A(new_n5417_), .B(new_n1499_), .Y(new_n5418_));
  NOR2  g05033(.A(new_n5418_), .B(new_n1503_), .Y(new_n5419_));
  NOR2  g05034(.A(new_n5419_), .B(new_n1507_), .Y(new_n5420_));
  NOR2  g05035(.A(new_n5420_), .B(new_n1511_), .Y(new_n5421_));
  NOR2  g05036(.A(new_n5421_), .B(new_n1515_), .Y(new_n5422_));
  NOR2  g05037(.A(new_n5422_), .B(new_n1519_), .Y(new_n5423_));
  NOR2  g05038(.A(new_n5423_), .B(new_n1523_), .Y(new_n5424_));
  NOR2  g05039(.A(new_n5424_), .B(new_n1527_), .Y(new_n5425_));
  NOR2  g05040(.A(new_n5425_), .B(new_n1797_), .Y(new_n5426_));
  NOR2  g05041(.A(new_n5426_), .B(new_n396_), .Y(new_n5427_));
  NOR2  g05042(.A(new_n5427_), .B(new_n400_), .Y(new_n5428_));
  NOR2  g05043(.A(new_n5428_), .B(new_n406_), .Y(new_n5429_));
  NOR2  g05044(.A(new_n5429_), .B(new_n410_), .Y(new_n5430_));
  NOR2  g05045(.A(new_n5430_), .B(new_n416_), .Y(new_n5431_));
  NOR2  g05046(.A(new_n5431_), .B(new_n420_), .Y(new_n5432_));
  NOR2  g05047(.A(new_n5432_), .B(new_n426_), .Y(new_n5433_));
  NOR2  g05048(.A(new_n5433_), .B(new_n430_), .Y(new_n5434_));
  NOR2  g05049(.A(new_n5434_), .B(new_n436_), .Y(new_n5435_));
  NOR2  g05050(.A(new_n5435_), .B(new_n440_), .Y(new_n5436_));
  NOR2  g05051(.A(new_n5436_), .B(new_n446_), .Y(new_n5437_));
  NOR2  g05052(.A(new_n5437_), .B(new_n450_), .Y(new_n5438_));
  NOR2  g05053(.A(new_n5438_), .B(new_n456_), .Y(new_n5439_));
  NOR2  g05054(.A(new_n5439_), .B(new_n460_), .Y(new_n5440_));
  NOR2  g05055(.A(new_n5440_), .B(new_n466_), .Y(new_n5441_));
  NOR2  g05056(.A(new_n5441_), .B(new_n470_), .Y(new_n5442_));
  NOR2  g05057(.A(new_n5442_), .B(new_n476_), .Y(new_n5443_));
  NOR2  g05058(.A(new_n5443_), .B(new_n480_), .Y(new_n5444_));
  NOR2  g05059(.A(new_n5444_), .B(new_n486_), .Y(new_n5445_));
  NOR2  g05060(.A(new_n5445_), .B(new_n490_), .Y(new_n5446_));
  NOR2  g05061(.A(new_n5446_), .B(new_n496_), .Y(new_n5447_));
  NOR2  g05062(.A(new_n5447_), .B(new_n500_), .Y(new_n5448_));
  NOR2  g05063(.A(new_n5448_), .B(new_n506_), .Y(new_n5449_));
  NOR2  g05064(.A(new_n5449_), .B(new_n510_), .Y(new_n5450_));
  NOR2  g05065(.A(new_n5450_), .B(new_n516_), .Y(new_n5451_));
  NOR2  g05066(.A(new_n5451_), .B(new_n520_), .Y(new_n5452_));
  NOR2  g05067(.A(new_n5452_), .B(new_n526_), .Y(new_n5453_));
  NOR2  g05068(.A(new_n5453_), .B(new_n530_), .Y(new_n5454_));
  NOR2  g05069(.A(new_n5454_), .B(new_n536_), .Y(new_n5455_));
  NAND2 g05070(.A(new_n538_), .B(\req[47] ), .Y(new_n5456_));
  NOR2  g05071(.A(new_n5456_), .B(new_n5455_), .Y(\grant[47] ));
  INV   g05072(.A(new_n549_), .Y(new_n5458_));
  NOR2  g05073(.A(new_n954_), .B(new_n5458_), .Y(new_n5459_));
  NOR2  g05074(.A(new_n5459_), .B(new_n556_), .Y(new_n5460_));
  NOR2  g05075(.A(new_n5460_), .B(new_n560_), .Y(new_n5461_));
  NOR2  g05076(.A(new_n5461_), .B(new_n566_), .Y(new_n5462_));
  NOR2  g05077(.A(new_n5462_), .B(new_n570_), .Y(new_n5463_));
  NOR2  g05078(.A(new_n5463_), .B(new_n576_), .Y(new_n5464_));
  NOR2  g05079(.A(new_n5464_), .B(new_n580_), .Y(new_n5465_));
  NOR2  g05080(.A(new_n5465_), .B(new_n586_), .Y(new_n5466_));
  NOR2  g05081(.A(new_n5466_), .B(new_n590_), .Y(new_n5467_));
  NOR2  g05082(.A(new_n5467_), .B(new_n596_), .Y(new_n5468_));
  NOR2  g05083(.A(new_n5468_), .B(new_n600_), .Y(new_n5469_));
  NOR2  g05084(.A(new_n5469_), .B(new_n606_), .Y(new_n5470_));
  NOR2  g05085(.A(new_n5470_), .B(new_n610_), .Y(new_n5471_));
  NOR2  g05086(.A(new_n5471_), .B(new_n616_), .Y(new_n5472_));
  NOR2  g05087(.A(new_n5472_), .B(new_n620_), .Y(new_n5473_));
  NOR2  g05088(.A(new_n5473_), .B(new_n626_), .Y(new_n5474_));
  NOR2  g05089(.A(new_n5474_), .B(new_n630_), .Y(new_n5475_));
  NOR2  g05090(.A(new_n5475_), .B(new_n636_), .Y(new_n5476_));
  NOR2  g05091(.A(new_n5476_), .B(new_n640_), .Y(new_n5477_));
  NOR2  g05092(.A(new_n5477_), .B(new_n646_), .Y(new_n5478_));
  NOR2  g05093(.A(new_n5478_), .B(new_n650_), .Y(new_n5479_));
  NOR2  g05094(.A(new_n5479_), .B(new_n656_), .Y(new_n5480_));
  NOR2  g05095(.A(new_n5480_), .B(new_n660_), .Y(new_n5481_));
  NOR2  g05096(.A(new_n5481_), .B(new_n666_), .Y(new_n5482_));
  NOR2  g05097(.A(new_n5482_), .B(new_n670_), .Y(new_n5483_));
  NOR2  g05098(.A(new_n5483_), .B(new_n676_), .Y(new_n5484_));
  NOR2  g05099(.A(new_n5484_), .B(new_n680_), .Y(new_n5485_));
  NOR2  g05100(.A(new_n5485_), .B(new_n686_), .Y(new_n5486_));
  NOR2  g05101(.A(new_n5486_), .B(new_n690_), .Y(new_n5487_));
  NOR2  g05102(.A(new_n5487_), .B(new_n696_), .Y(new_n5488_));
  NOR2  g05103(.A(new_n5488_), .B(new_n700_), .Y(new_n5489_));
  NOR2  g05104(.A(new_n5489_), .B(new_n706_), .Y(new_n5490_));
  NOR2  g05105(.A(new_n5490_), .B(new_n710_), .Y(new_n5491_));
  NOR2  g05106(.A(new_n5491_), .B(new_n716_), .Y(new_n5492_));
  NOR2  g05107(.A(new_n5492_), .B(new_n720_), .Y(new_n5493_));
  NOR2  g05108(.A(new_n5493_), .B(new_n726_), .Y(new_n5494_));
  NOR2  g05109(.A(new_n5494_), .B(new_n730_), .Y(new_n5495_));
  NOR2  g05110(.A(new_n5495_), .B(new_n736_), .Y(new_n5496_));
  NOR2  g05111(.A(new_n5496_), .B(new_n740_), .Y(new_n5497_));
  NOR2  g05112(.A(new_n5497_), .B(new_n746_), .Y(new_n5498_));
  NOR2  g05113(.A(new_n5498_), .B(new_n750_), .Y(new_n5499_));
  NOR2  g05114(.A(new_n5499_), .B(new_n756_), .Y(new_n5500_));
  NOR2  g05115(.A(new_n5500_), .B(new_n760_), .Y(new_n5501_));
  NOR2  g05116(.A(new_n5501_), .B(new_n766_), .Y(new_n5502_));
  NOR2  g05117(.A(new_n5502_), .B(new_n770_), .Y(new_n5503_));
  NOR2  g05118(.A(new_n5503_), .B(new_n776_), .Y(new_n5504_));
  NOR2  g05119(.A(new_n5504_), .B(new_n780_), .Y(new_n5505_));
  NOR2  g05120(.A(new_n5505_), .B(new_n786_), .Y(new_n5506_));
  NOR2  g05121(.A(new_n5506_), .B(new_n790_), .Y(new_n5507_));
  NOR2  g05122(.A(new_n5507_), .B(new_n796_), .Y(new_n5508_));
  NOR2  g05123(.A(new_n5508_), .B(new_n800_), .Y(new_n5509_));
  NOR2  g05124(.A(new_n5509_), .B(new_n806_), .Y(new_n5510_));
  NOR2  g05125(.A(new_n5510_), .B(new_n1616_), .Y(new_n5511_));
  NOR2  g05126(.A(new_n5511_), .B(new_n1618_), .Y(new_n5512_));
  NOR2  g05127(.A(new_n5512_), .B(new_n1885_), .Y(new_n5513_));
  NOR2  g05128(.A(new_n5513_), .B(new_n820_), .Y(new_n5514_));
  NOR2  g05129(.A(new_n5514_), .B(new_n824_), .Y(new_n5515_));
  NOR2  g05130(.A(new_n5515_), .B(new_n829_), .Y(new_n5516_));
  NOR2  g05131(.A(new_n5516_), .B(new_n833_), .Y(new_n5517_));
  NOR2  g05132(.A(new_n5517_), .B(new_n838_), .Y(new_n5518_));
  NOR2  g05133(.A(new_n5518_), .B(new_n842_), .Y(new_n5519_));
  NOR2  g05134(.A(new_n5519_), .B(new_n847_), .Y(new_n5520_));
  NOR2  g05135(.A(new_n5520_), .B(new_n851_), .Y(new_n5521_));
  NOR2  g05136(.A(new_n5521_), .B(new_n856_), .Y(new_n5522_));
  NOR2  g05137(.A(new_n5522_), .B(new_n860_), .Y(new_n5523_));
  NOR2  g05138(.A(new_n5523_), .B(new_n865_), .Y(new_n5524_));
  NOR2  g05139(.A(new_n5524_), .B(new_n869_), .Y(new_n5525_));
  NOR2  g05140(.A(new_n5525_), .B(new_n874_), .Y(new_n5526_));
  NOR2  g05141(.A(new_n5526_), .B(new_n878_), .Y(new_n5527_));
  NOR2  g05142(.A(new_n5527_), .B(new_n883_), .Y(new_n5528_));
  NOR2  g05143(.A(new_n5528_), .B(new_n887_), .Y(new_n5529_));
  NOR2  g05144(.A(new_n5529_), .B(new_n892_), .Y(new_n5530_));
  NOR2  g05145(.A(new_n5530_), .B(new_n896_), .Y(new_n5531_));
  NOR2  g05146(.A(new_n5531_), .B(new_n901_), .Y(new_n5532_));
  NOR2  g05147(.A(new_n5532_), .B(new_n905_), .Y(new_n5533_));
  NOR2  g05148(.A(new_n5533_), .B(new_n910_), .Y(new_n5534_));
  NOR2  g05149(.A(new_n5534_), .B(new_n914_), .Y(new_n5535_));
  NOR2  g05150(.A(new_n5535_), .B(new_n919_), .Y(new_n5536_));
  NOR2  g05151(.A(new_n5536_), .B(new_n923_), .Y(new_n5537_));
  NOR2  g05152(.A(new_n5537_), .B(new_n928_), .Y(new_n5538_));
  NOR2  g05153(.A(new_n5538_), .B(new_n932_), .Y(new_n5539_));
  NOR2  g05154(.A(new_n5539_), .B(new_n937_), .Y(new_n5540_));
  NOR2  g05155(.A(new_n5540_), .B(new_n941_), .Y(new_n5541_));
  NOR2  g05156(.A(new_n5541_), .B(new_n946_), .Y(new_n5542_));
  NAND2 g05157(.A(new_n948_), .B(\req[48] ), .Y(new_n5543_));
  NOR2  g05158(.A(new_n5543_), .B(new_n5542_), .Y(\grant[48] ));
  INV   g05159(.A(new_n958_), .Y(new_n5545_));
  NOR2  g05160(.A(new_n1318_), .B(new_n5545_), .Y(new_n5546_));
  NOR2  g05161(.A(new_n5546_), .B(new_n964_), .Y(new_n5547_));
  NOR2  g05162(.A(new_n5547_), .B(new_n968_), .Y(new_n5548_));
  NOR2  g05163(.A(new_n5548_), .B(new_n973_), .Y(new_n5549_));
  NOR2  g05164(.A(new_n5549_), .B(new_n977_), .Y(new_n5550_));
  NOR2  g05165(.A(new_n5550_), .B(new_n982_), .Y(new_n5551_));
  NOR2  g05166(.A(new_n5551_), .B(new_n986_), .Y(new_n5552_));
  NOR2  g05167(.A(new_n5552_), .B(new_n991_), .Y(new_n5553_));
  NOR2  g05168(.A(new_n5553_), .B(new_n995_), .Y(new_n5554_));
  NOR2  g05169(.A(new_n5554_), .B(new_n1000_), .Y(new_n5555_));
  NOR2  g05170(.A(new_n5555_), .B(new_n1004_), .Y(new_n5556_));
  NOR2  g05171(.A(new_n5556_), .B(new_n1009_), .Y(new_n5557_));
  NOR2  g05172(.A(new_n5557_), .B(new_n1013_), .Y(new_n5558_));
  NOR2  g05173(.A(new_n5558_), .B(new_n1018_), .Y(new_n5559_));
  NOR2  g05174(.A(new_n5559_), .B(new_n1022_), .Y(new_n5560_));
  NOR2  g05175(.A(new_n5560_), .B(new_n1027_), .Y(new_n5561_));
  NOR2  g05176(.A(new_n5561_), .B(new_n1031_), .Y(new_n5562_));
  NOR2  g05177(.A(new_n5562_), .B(new_n1036_), .Y(new_n5563_));
  NOR2  g05178(.A(new_n5563_), .B(new_n1040_), .Y(new_n5564_));
  NOR2  g05179(.A(new_n5564_), .B(new_n1045_), .Y(new_n5565_));
  NOR2  g05180(.A(new_n5565_), .B(new_n1049_), .Y(new_n5566_));
  NOR2  g05181(.A(new_n5566_), .B(new_n1054_), .Y(new_n5567_));
  NOR2  g05182(.A(new_n5567_), .B(new_n1058_), .Y(new_n5568_));
  NOR2  g05183(.A(new_n5568_), .B(new_n1063_), .Y(new_n5569_));
  NOR2  g05184(.A(new_n5569_), .B(new_n1067_), .Y(new_n5570_));
  NOR2  g05185(.A(new_n5570_), .B(new_n1072_), .Y(new_n5571_));
  NOR2  g05186(.A(new_n5571_), .B(new_n1076_), .Y(new_n5572_));
  NOR2  g05187(.A(new_n5572_), .B(new_n1081_), .Y(new_n5573_));
  NOR2  g05188(.A(new_n5573_), .B(new_n1085_), .Y(new_n5574_));
  NOR2  g05189(.A(new_n5574_), .B(new_n1090_), .Y(new_n5575_));
  NOR2  g05190(.A(new_n5575_), .B(new_n1094_), .Y(new_n5576_));
  NOR2  g05191(.A(new_n5576_), .B(new_n1099_), .Y(new_n5577_));
  NOR2  g05192(.A(new_n5577_), .B(new_n1103_), .Y(new_n5578_));
  NOR2  g05193(.A(new_n5578_), .B(new_n1108_), .Y(new_n5579_));
  NOR2  g05194(.A(new_n5579_), .B(new_n1112_), .Y(new_n5580_));
  NOR2  g05195(.A(new_n5580_), .B(new_n1117_), .Y(new_n5581_));
  NOR2  g05196(.A(new_n5581_), .B(new_n1121_), .Y(new_n5582_));
  NOR2  g05197(.A(new_n5582_), .B(new_n1126_), .Y(new_n5583_));
  NOR2  g05198(.A(new_n5583_), .B(new_n1130_), .Y(new_n5584_));
  NOR2  g05199(.A(new_n5584_), .B(new_n1135_), .Y(new_n5585_));
  NOR2  g05200(.A(new_n5585_), .B(new_n1139_), .Y(new_n5586_));
  NOR2  g05201(.A(new_n5586_), .B(new_n1144_), .Y(new_n5587_));
  NOR2  g05202(.A(new_n5587_), .B(new_n1148_), .Y(new_n5588_));
  NOR2  g05203(.A(new_n5588_), .B(new_n1153_), .Y(new_n5589_));
  NOR2  g05204(.A(new_n5589_), .B(new_n1157_), .Y(new_n5590_));
  NOR2  g05205(.A(new_n5590_), .B(new_n1162_), .Y(new_n5591_));
  NOR2  g05206(.A(new_n5591_), .B(new_n1166_), .Y(new_n5592_));
  NOR2  g05207(.A(new_n5592_), .B(new_n1171_), .Y(new_n5593_));
  NOR2  g05208(.A(new_n5593_), .B(new_n1175_), .Y(new_n5594_));
  NOR2  g05209(.A(new_n5594_), .B(new_n1180_), .Y(new_n5595_));
  NOR2  g05210(.A(new_n5595_), .B(new_n1184_), .Y(new_n5596_));
  NOR2  g05211(.A(new_n5596_), .B(new_n1189_), .Y(new_n5597_));
  NOR2  g05212(.A(new_n5597_), .B(new_n1707_), .Y(new_n5598_));
  NOR2  g05213(.A(new_n5598_), .B(new_n1709_), .Y(new_n5599_));
  NOR2  g05214(.A(new_n5599_), .B(new_n1973_), .Y(new_n5600_));
  NOR2  g05215(.A(new_n5600_), .B(new_n1199_), .Y(new_n5601_));
  NOR2  g05216(.A(new_n5601_), .B(new_n1203_), .Y(new_n5602_));
  NOR2  g05217(.A(new_n5602_), .B(new_n1207_), .Y(new_n5603_));
  NOR2  g05218(.A(new_n5603_), .B(new_n1211_), .Y(new_n5604_));
  NOR2  g05219(.A(new_n5604_), .B(new_n1215_), .Y(new_n5605_));
  NOR2  g05220(.A(new_n5605_), .B(new_n1219_), .Y(new_n5606_));
  NOR2  g05221(.A(new_n5606_), .B(new_n1223_), .Y(new_n5607_));
  NOR2  g05222(.A(new_n5607_), .B(new_n1227_), .Y(new_n5608_));
  NOR2  g05223(.A(new_n5608_), .B(new_n1231_), .Y(new_n5609_));
  NOR2  g05224(.A(new_n5609_), .B(new_n1235_), .Y(new_n5610_));
  NOR2  g05225(.A(new_n5610_), .B(new_n1239_), .Y(new_n5611_));
  NOR2  g05226(.A(new_n5611_), .B(new_n1243_), .Y(new_n5612_));
  NOR2  g05227(.A(new_n5612_), .B(new_n1247_), .Y(new_n5613_));
  NOR2  g05228(.A(new_n5613_), .B(new_n1251_), .Y(new_n5614_));
  NOR2  g05229(.A(new_n5614_), .B(new_n1255_), .Y(new_n5615_));
  NOR2  g05230(.A(new_n5615_), .B(new_n1259_), .Y(new_n5616_));
  NOR2  g05231(.A(new_n5616_), .B(new_n1263_), .Y(new_n5617_));
  NOR2  g05232(.A(new_n5617_), .B(new_n1267_), .Y(new_n5618_));
  NOR2  g05233(.A(new_n5618_), .B(new_n1271_), .Y(new_n5619_));
  NOR2  g05234(.A(new_n5619_), .B(new_n1275_), .Y(new_n5620_));
  NOR2  g05235(.A(new_n5620_), .B(new_n1279_), .Y(new_n5621_));
  NOR2  g05236(.A(new_n5621_), .B(new_n1283_), .Y(new_n5622_));
  NOR2  g05237(.A(new_n5622_), .B(new_n1287_), .Y(new_n5623_));
  NOR2  g05238(.A(new_n5623_), .B(new_n1291_), .Y(new_n5624_));
  NOR2  g05239(.A(new_n5624_), .B(new_n1295_), .Y(new_n5625_));
  NOR2  g05240(.A(new_n5625_), .B(new_n1299_), .Y(new_n5626_));
  NOR2  g05241(.A(new_n5626_), .B(new_n1303_), .Y(new_n5627_));
  NOR2  g05242(.A(new_n5627_), .B(new_n1307_), .Y(new_n5628_));
  NOR2  g05243(.A(new_n5628_), .B(new_n1311_), .Y(new_n5629_));
  NAND2 g05244(.A(new_n1313_), .B(\req[49] ), .Y(new_n5630_));
  NOR2  g05245(.A(new_n5630_), .B(new_n5629_), .Y(\grant[49] ));
  INV   g05246(.A(new_n1322_), .Y(new_n5632_));
  NOR2  g05247(.A(new_n5632_), .B(new_n555_), .Y(new_n5633_));
  NOR2  g05248(.A(new_n5633_), .B(new_n1327_), .Y(new_n5634_));
  NOR2  g05249(.A(new_n5634_), .B(new_n1331_), .Y(new_n5635_));
  NOR2  g05250(.A(new_n5635_), .B(new_n1335_), .Y(new_n5636_));
  NOR2  g05251(.A(new_n5636_), .B(new_n1339_), .Y(new_n5637_));
  NOR2  g05252(.A(new_n5637_), .B(new_n1343_), .Y(new_n5638_));
  NOR2  g05253(.A(new_n5638_), .B(new_n1347_), .Y(new_n5639_));
  NOR2  g05254(.A(new_n5639_), .B(new_n1351_), .Y(new_n5640_));
  NOR2  g05255(.A(new_n5640_), .B(new_n1355_), .Y(new_n5641_));
  NOR2  g05256(.A(new_n5641_), .B(new_n1359_), .Y(new_n5642_));
  NOR2  g05257(.A(new_n5642_), .B(new_n1363_), .Y(new_n5643_));
  NOR2  g05258(.A(new_n5643_), .B(new_n1367_), .Y(new_n5644_));
  NOR2  g05259(.A(new_n5644_), .B(new_n1371_), .Y(new_n5645_));
  NOR2  g05260(.A(new_n5645_), .B(new_n1375_), .Y(new_n5646_));
  NOR2  g05261(.A(new_n5646_), .B(new_n1379_), .Y(new_n5647_));
  NOR2  g05262(.A(new_n5647_), .B(new_n1383_), .Y(new_n5648_));
  NOR2  g05263(.A(new_n5648_), .B(new_n1387_), .Y(new_n5649_));
  NOR2  g05264(.A(new_n5649_), .B(new_n1391_), .Y(new_n5650_));
  NOR2  g05265(.A(new_n5650_), .B(new_n1395_), .Y(new_n5651_));
  NOR2  g05266(.A(new_n5651_), .B(new_n1399_), .Y(new_n5652_));
  NOR2  g05267(.A(new_n5652_), .B(new_n1403_), .Y(new_n5653_));
  NOR2  g05268(.A(new_n5653_), .B(new_n1407_), .Y(new_n5654_));
  NOR2  g05269(.A(new_n5654_), .B(new_n1411_), .Y(new_n5655_));
  NOR2  g05270(.A(new_n5655_), .B(new_n1415_), .Y(new_n5656_));
  NOR2  g05271(.A(new_n5656_), .B(new_n1419_), .Y(new_n5657_));
  NOR2  g05272(.A(new_n5657_), .B(new_n1423_), .Y(new_n5658_));
  NOR2  g05273(.A(new_n5658_), .B(new_n1427_), .Y(new_n5659_));
  NOR2  g05274(.A(new_n5659_), .B(new_n1431_), .Y(new_n5660_));
  NOR2  g05275(.A(new_n5660_), .B(new_n1435_), .Y(new_n5661_));
  NOR2  g05276(.A(new_n5661_), .B(new_n1439_), .Y(new_n5662_));
  NOR2  g05277(.A(new_n5662_), .B(new_n1443_), .Y(new_n5663_));
  NOR2  g05278(.A(new_n5663_), .B(new_n1447_), .Y(new_n5664_));
  NOR2  g05279(.A(new_n5664_), .B(new_n1451_), .Y(new_n5665_));
  NOR2  g05280(.A(new_n5665_), .B(new_n1455_), .Y(new_n5666_));
  NOR2  g05281(.A(new_n5666_), .B(new_n1459_), .Y(new_n5667_));
  NOR2  g05282(.A(new_n5667_), .B(new_n1463_), .Y(new_n5668_));
  NOR2  g05283(.A(new_n5668_), .B(new_n1467_), .Y(new_n5669_));
  NOR2  g05284(.A(new_n5669_), .B(new_n1471_), .Y(new_n5670_));
  NOR2  g05285(.A(new_n5670_), .B(new_n1475_), .Y(new_n5671_));
  NOR2  g05286(.A(new_n5671_), .B(new_n1479_), .Y(new_n5672_));
  NOR2  g05287(.A(new_n5672_), .B(new_n1483_), .Y(new_n5673_));
  NOR2  g05288(.A(new_n5673_), .B(new_n1487_), .Y(new_n5674_));
  NOR2  g05289(.A(new_n5674_), .B(new_n1491_), .Y(new_n5675_));
  NOR2  g05290(.A(new_n5675_), .B(new_n1495_), .Y(new_n5676_));
  NOR2  g05291(.A(new_n5676_), .B(new_n1499_), .Y(new_n5677_));
  NOR2  g05292(.A(new_n5677_), .B(new_n1503_), .Y(new_n5678_));
  NOR2  g05293(.A(new_n5678_), .B(new_n1507_), .Y(new_n5679_));
  NOR2  g05294(.A(new_n5679_), .B(new_n1511_), .Y(new_n5680_));
  NOR2  g05295(.A(new_n5680_), .B(new_n1515_), .Y(new_n5681_));
  NOR2  g05296(.A(new_n5681_), .B(new_n1519_), .Y(new_n5682_));
  NOR2  g05297(.A(new_n5682_), .B(new_n1523_), .Y(new_n5683_));
  NOR2  g05298(.A(new_n5683_), .B(new_n1527_), .Y(new_n5684_));
  NOR2  g05299(.A(new_n5684_), .B(new_n1797_), .Y(new_n5685_));
  NOR2  g05300(.A(new_n5685_), .B(new_n396_), .Y(new_n5686_));
  NOR2  g05301(.A(new_n5686_), .B(new_n400_), .Y(new_n5687_));
  NOR2  g05302(.A(new_n5687_), .B(new_n406_), .Y(new_n5688_));
  NOR2  g05303(.A(new_n5688_), .B(new_n410_), .Y(new_n5689_));
  NOR2  g05304(.A(new_n5689_), .B(new_n416_), .Y(new_n5690_));
  NOR2  g05305(.A(new_n5690_), .B(new_n420_), .Y(new_n5691_));
  NOR2  g05306(.A(new_n5691_), .B(new_n426_), .Y(new_n5692_));
  NOR2  g05307(.A(new_n5692_), .B(new_n430_), .Y(new_n5693_));
  NOR2  g05308(.A(new_n5693_), .B(new_n436_), .Y(new_n5694_));
  NOR2  g05309(.A(new_n5694_), .B(new_n440_), .Y(new_n5695_));
  NOR2  g05310(.A(new_n5695_), .B(new_n446_), .Y(new_n5696_));
  NOR2  g05311(.A(new_n5696_), .B(new_n450_), .Y(new_n5697_));
  NOR2  g05312(.A(new_n5697_), .B(new_n456_), .Y(new_n5698_));
  NOR2  g05313(.A(new_n5698_), .B(new_n460_), .Y(new_n5699_));
  NOR2  g05314(.A(new_n5699_), .B(new_n466_), .Y(new_n5700_));
  NOR2  g05315(.A(new_n5700_), .B(new_n470_), .Y(new_n5701_));
  NOR2  g05316(.A(new_n5701_), .B(new_n476_), .Y(new_n5702_));
  NOR2  g05317(.A(new_n5702_), .B(new_n480_), .Y(new_n5703_));
  NOR2  g05318(.A(new_n5703_), .B(new_n486_), .Y(new_n5704_));
  NOR2  g05319(.A(new_n5704_), .B(new_n490_), .Y(new_n5705_));
  NOR2  g05320(.A(new_n5705_), .B(new_n496_), .Y(new_n5706_));
  NOR2  g05321(.A(new_n5706_), .B(new_n500_), .Y(new_n5707_));
  NOR2  g05322(.A(new_n5707_), .B(new_n506_), .Y(new_n5708_));
  NOR2  g05323(.A(new_n5708_), .B(new_n510_), .Y(new_n5709_));
  NOR2  g05324(.A(new_n5709_), .B(new_n516_), .Y(new_n5710_));
  NOR2  g05325(.A(new_n5710_), .B(new_n520_), .Y(new_n5711_));
  NOR2  g05326(.A(new_n5711_), .B(new_n526_), .Y(new_n5712_));
  NOR2  g05327(.A(new_n5712_), .B(new_n530_), .Y(new_n5713_));
  NOR2  g05328(.A(new_n5713_), .B(new_n536_), .Y(new_n5714_));
  NOR2  g05329(.A(new_n5714_), .B(new_n540_), .Y(new_n5715_));
  NOR2  g05330(.A(new_n5715_), .B(new_n546_), .Y(new_n5716_));
  NAND2 g05331(.A(new_n548_), .B(\req[50] ), .Y(new_n5717_));
  NOR2  g05332(.A(new_n5717_), .B(new_n5716_), .Y(\grant[50] ));
  INV   g05333(.A(new_n559_), .Y(new_n5719_));
  NOR2  g05334(.A(new_n963_), .B(new_n5719_), .Y(new_n5720_));
  NOR2  g05335(.A(new_n5720_), .B(new_n566_), .Y(new_n5721_));
  NOR2  g05336(.A(new_n5721_), .B(new_n570_), .Y(new_n5722_));
  NOR2  g05337(.A(new_n5722_), .B(new_n576_), .Y(new_n5723_));
  NOR2  g05338(.A(new_n5723_), .B(new_n580_), .Y(new_n5724_));
  NOR2  g05339(.A(new_n5724_), .B(new_n586_), .Y(new_n5725_));
  NOR2  g05340(.A(new_n5725_), .B(new_n590_), .Y(new_n5726_));
  NOR2  g05341(.A(new_n5726_), .B(new_n596_), .Y(new_n5727_));
  NOR2  g05342(.A(new_n5727_), .B(new_n600_), .Y(new_n5728_));
  NOR2  g05343(.A(new_n5728_), .B(new_n606_), .Y(new_n5729_));
  NOR2  g05344(.A(new_n5729_), .B(new_n610_), .Y(new_n5730_));
  NOR2  g05345(.A(new_n5730_), .B(new_n616_), .Y(new_n5731_));
  NOR2  g05346(.A(new_n5731_), .B(new_n620_), .Y(new_n5732_));
  NOR2  g05347(.A(new_n5732_), .B(new_n626_), .Y(new_n5733_));
  NOR2  g05348(.A(new_n5733_), .B(new_n630_), .Y(new_n5734_));
  NOR2  g05349(.A(new_n5734_), .B(new_n636_), .Y(new_n5735_));
  NOR2  g05350(.A(new_n5735_), .B(new_n640_), .Y(new_n5736_));
  NOR2  g05351(.A(new_n5736_), .B(new_n646_), .Y(new_n5737_));
  NOR2  g05352(.A(new_n5737_), .B(new_n650_), .Y(new_n5738_));
  NOR2  g05353(.A(new_n5738_), .B(new_n656_), .Y(new_n5739_));
  NOR2  g05354(.A(new_n5739_), .B(new_n660_), .Y(new_n5740_));
  NOR2  g05355(.A(new_n5740_), .B(new_n666_), .Y(new_n5741_));
  NOR2  g05356(.A(new_n5741_), .B(new_n670_), .Y(new_n5742_));
  NOR2  g05357(.A(new_n5742_), .B(new_n676_), .Y(new_n5743_));
  NOR2  g05358(.A(new_n5743_), .B(new_n680_), .Y(new_n5744_));
  NOR2  g05359(.A(new_n5744_), .B(new_n686_), .Y(new_n5745_));
  NOR2  g05360(.A(new_n5745_), .B(new_n690_), .Y(new_n5746_));
  NOR2  g05361(.A(new_n5746_), .B(new_n696_), .Y(new_n5747_));
  NOR2  g05362(.A(new_n5747_), .B(new_n700_), .Y(new_n5748_));
  NOR2  g05363(.A(new_n5748_), .B(new_n706_), .Y(new_n5749_));
  NOR2  g05364(.A(new_n5749_), .B(new_n710_), .Y(new_n5750_));
  NOR2  g05365(.A(new_n5750_), .B(new_n716_), .Y(new_n5751_));
  NOR2  g05366(.A(new_n5751_), .B(new_n720_), .Y(new_n5752_));
  NOR2  g05367(.A(new_n5752_), .B(new_n726_), .Y(new_n5753_));
  NOR2  g05368(.A(new_n5753_), .B(new_n730_), .Y(new_n5754_));
  NOR2  g05369(.A(new_n5754_), .B(new_n736_), .Y(new_n5755_));
  NOR2  g05370(.A(new_n5755_), .B(new_n740_), .Y(new_n5756_));
  NOR2  g05371(.A(new_n5756_), .B(new_n746_), .Y(new_n5757_));
  NOR2  g05372(.A(new_n5757_), .B(new_n750_), .Y(new_n5758_));
  NOR2  g05373(.A(new_n5758_), .B(new_n756_), .Y(new_n5759_));
  NOR2  g05374(.A(new_n5759_), .B(new_n760_), .Y(new_n5760_));
  NOR2  g05375(.A(new_n5760_), .B(new_n766_), .Y(new_n5761_));
  NOR2  g05376(.A(new_n5761_), .B(new_n770_), .Y(new_n5762_));
  NOR2  g05377(.A(new_n5762_), .B(new_n776_), .Y(new_n5763_));
  NOR2  g05378(.A(new_n5763_), .B(new_n780_), .Y(new_n5764_));
  NOR2  g05379(.A(new_n5764_), .B(new_n786_), .Y(new_n5765_));
  NOR2  g05380(.A(new_n5765_), .B(new_n790_), .Y(new_n5766_));
  NOR2  g05381(.A(new_n5766_), .B(new_n796_), .Y(new_n5767_));
  NOR2  g05382(.A(new_n5767_), .B(new_n800_), .Y(new_n5768_));
  NOR2  g05383(.A(new_n5768_), .B(new_n806_), .Y(new_n5769_));
  NOR2  g05384(.A(new_n5769_), .B(new_n1616_), .Y(new_n5770_));
  NOR2  g05385(.A(new_n5770_), .B(new_n1618_), .Y(new_n5771_));
  NOR2  g05386(.A(new_n5771_), .B(new_n1885_), .Y(new_n5772_));
  NOR2  g05387(.A(new_n5772_), .B(new_n820_), .Y(new_n5773_));
  NOR2  g05388(.A(new_n5773_), .B(new_n824_), .Y(new_n5774_));
  NOR2  g05389(.A(new_n5774_), .B(new_n829_), .Y(new_n5775_));
  NOR2  g05390(.A(new_n5775_), .B(new_n833_), .Y(new_n5776_));
  NOR2  g05391(.A(new_n5776_), .B(new_n838_), .Y(new_n5777_));
  NOR2  g05392(.A(new_n5777_), .B(new_n842_), .Y(new_n5778_));
  NOR2  g05393(.A(new_n5778_), .B(new_n847_), .Y(new_n5779_));
  NOR2  g05394(.A(new_n5779_), .B(new_n851_), .Y(new_n5780_));
  NOR2  g05395(.A(new_n5780_), .B(new_n856_), .Y(new_n5781_));
  NOR2  g05396(.A(new_n5781_), .B(new_n860_), .Y(new_n5782_));
  NOR2  g05397(.A(new_n5782_), .B(new_n865_), .Y(new_n5783_));
  NOR2  g05398(.A(new_n5783_), .B(new_n869_), .Y(new_n5784_));
  NOR2  g05399(.A(new_n5784_), .B(new_n874_), .Y(new_n5785_));
  NOR2  g05400(.A(new_n5785_), .B(new_n878_), .Y(new_n5786_));
  NOR2  g05401(.A(new_n5786_), .B(new_n883_), .Y(new_n5787_));
  NOR2  g05402(.A(new_n5787_), .B(new_n887_), .Y(new_n5788_));
  NOR2  g05403(.A(new_n5788_), .B(new_n892_), .Y(new_n5789_));
  NOR2  g05404(.A(new_n5789_), .B(new_n896_), .Y(new_n5790_));
  NOR2  g05405(.A(new_n5790_), .B(new_n901_), .Y(new_n5791_));
  NOR2  g05406(.A(new_n5791_), .B(new_n905_), .Y(new_n5792_));
  NOR2  g05407(.A(new_n5792_), .B(new_n910_), .Y(new_n5793_));
  NOR2  g05408(.A(new_n5793_), .B(new_n914_), .Y(new_n5794_));
  NOR2  g05409(.A(new_n5794_), .B(new_n919_), .Y(new_n5795_));
  NOR2  g05410(.A(new_n5795_), .B(new_n923_), .Y(new_n5796_));
  NOR2  g05411(.A(new_n5796_), .B(new_n928_), .Y(new_n5797_));
  NOR2  g05412(.A(new_n5797_), .B(new_n932_), .Y(new_n5798_));
  NOR2  g05413(.A(new_n5798_), .B(new_n937_), .Y(new_n5799_));
  NOR2  g05414(.A(new_n5799_), .B(new_n941_), .Y(new_n5800_));
  NOR2  g05415(.A(new_n5800_), .B(new_n946_), .Y(new_n5801_));
  NOR2  g05416(.A(new_n5801_), .B(new_n950_), .Y(new_n5802_));
  NOR2  g05417(.A(new_n5802_), .B(new_n955_), .Y(new_n5803_));
  NAND2 g05418(.A(new_n957_), .B(\req[51] ), .Y(new_n5804_));
  NOR2  g05419(.A(new_n5804_), .B(new_n5803_), .Y(\grant[51] ));
  INV   g05420(.A(new_n967_), .Y(new_n5806_));
  NOR2  g05421(.A(new_n1326_), .B(new_n5806_), .Y(new_n5807_));
  NOR2  g05422(.A(new_n5807_), .B(new_n973_), .Y(new_n5808_));
  NOR2  g05423(.A(new_n5808_), .B(new_n977_), .Y(new_n5809_));
  NOR2  g05424(.A(new_n5809_), .B(new_n982_), .Y(new_n5810_));
  NOR2  g05425(.A(new_n5810_), .B(new_n986_), .Y(new_n5811_));
  NOR2  g05426(.A(new_n5811_), .B(new_n991_), .Y(new_n5812_));
  NOR2  g05427(.A(new_n5812_), .B(new_n995_), .Y(new_n5813_));
  NOR2  g05428(.A(new_n5813_), .B(new_n1000_), .Y(new_n5814_));
  NOR2  g05429(.A(new_n5814_), .B(new_n1004_), .Y(new_n5815_));
  NOR2  g05430(.A(new_n5815_), .B(new_n1009_), .Y(new_n5816_));
  NOR2  g05431(.A(new_n5816_), .B(new_n1013_), .Y(new_n5817_));
  NOR2  g05432(.A(new_n5817_), .B(new_n1018_), .Y(new_n5818_));
  NOR2  g05433(.A(new_n5818_), .B(new_n1022_), .Y(new_n5819_));
  NOR2  g05434(.A(new_n5819_), .B(new_n1027_), .Y(new_n5820_));
  NOR2  g05435(.A(new_n5820_), .B(new_n1031_), .Y(new_n5821_));
  NOR2  g05436(.A(new_n5821_), .B(new_n1036_), .Y(new_n5822_));
  NOR2  g05437(.A(new_n5822_), .B(new_n1040_), .Y(new_n5823_));
  NOR2  g05438(.A(new_n5823_), .B(new_n1045_), .Y(new_n5824_));
  NOR2  g05439(.A(new_n5824_), .B(new_n1049_), .Y(new_n5825_));
  NOR2  g05440(.A(new_n5825_), .B(new_n1054_), .Y(new_n5826_));
  NOR2  g05441(.A(new_n5826_), .B(new_n1058_), .Y(new_n5827_));
  NOR2  g05442(.A(new_n5827_), .B(new_n1063_), .Y(new_n5828_));
  NOR2  g05443(.A(new_n5828_), .B(new_n1067_), .Y(new_n5829_));
  NOR2  g05444(.A(new_n5829_), .B(new_n1072_), .Y(new_n5830_));
  NOR2  g05445(.A(new_n5830_), .B(new_n1076_), .Y(new_n5831_));
  NOR2  g05446(.A(new_n5831_), .B(new_n1081_), .Y(new_n5832_));
  NOR2  g05447(.A(new_n5832_), .B(new_n1085_), .Y(new_n5833_));
  NOR2  g05448(.A(new_n5833_), .B(new_n1090_), .Y(new_n5834_));
  NOR2  g05449(.A(new_n5834_), .B(new_n1094_), .Y(new_n5835_));
  NOR2  g05450(.A(new_n5835_), .B(new_n1099_), .Y(new_n5836_));
  NOR2  g05451(.A(new_n5836_), .B(new_n1103_), .Y(new_n5837_));
  NOR2  g05452(.A(new_n5837_), .B(new_n1108_), .Y(new_n5838_));
  NOR2  g05453(.A(new_n5838_), .B(new_n1112_), .Y(new_n5839_));
  NOR2  g05454(.A(new_n5839_), .B(new_n1117_), .Y(new_n5840_));
  NOR2  g05455(.A(new_n5840_), .B(new_n1121_), .Y(new_n5841_));
  NOR2  g05456(.A(new_n5841_), .B(new_n1126_), .Y(new_n5842_));
  NOR2  g05457(.A(new_n5842_), .B(new_n1130_), .Y(new_n5843_));
  NOR2  g05458(.A(new_n5843_), .B(new_n1135_), .Y(new_n5844_));
  NOR2  g05459(.A(new_n5844_), .B(new_n1139_), .Y(new_n5845_));
  NOR2  g05460(.A(new_n5845_), .B(new_n1144_), .Y(new_n5846_));
  NOR2  g05461(.A(new_n5846_), .B(new_n1148_), .Y(new_n5847_));
  NOR2  g05462(.A(new_n5847_), .B(new_n1153_), .Y(new_n5848_));
  NOR2  g05463(.A(new_n5848_), .B(new_n1157_), .Y(new_n5849_));
  NOR2  g05464(.A(new_n5849_), .B(new_n1162_), .Y(new_n5850_));
  NOR2  g05465(.A(new_n5850_), .B(new_n1166_), .Y(new_n5851_));
  NOR2  g05466(.A(new_n5851_), .B(new_n1171_), .Y(new_n5852_));
  NOR2  g05467(.A(new_n5852_), .B(new_n1175_), .Y(new_n5853_));
  NOR2  g05468(.A(new_n5853_), .B(new_n1180_), .Y(new_n5854_));
  NOR2  g05469(.A(new_n5854_), .B(new_n1184_), .Y(new_n5855_));
  NOR2  g05470(.A(new_n5855_), .B(new_n1189_), .Y(new_n5856_));
  NOR2  g05471(.A(new_n5856_), .B(new_n1707_), .Y(new_n5857_));
  NOR2  g05472(.A(new_n5857_), .B(new_n1709_), .Y(new_n5858_));
  NOR2  g05473(.A(new_n5858_), .B(new_n1973_), .Y(new_n5859_));
  NOR2  g05474(.A(new_n5859_), .B(new_n1199_), .Y(new_n5860_));
  NOR2  g05475(.A(new_n5860_), .B(new_n1203_), .Y(new_n5861_));
  NOR2  g05476(.A(new_n5861_), .B(new_n1207_), .Y(new_n5862_));
  NOR2  g05477(.A(new_n5862_), .B(new_n1211_), .Y(new_n5863_));
  NOR2  g05478(.A(new_n5863_), .B(new_n1215_), .Y(new_n5864_));
  NOR2  g05479(.A(new_n5864_), .B(new_n1219_), .Y(new_n5865_));
  NOR2  g05480(.A(new_n5865_), .B(new_n1223_), .Y(new_n5866_));
  NOR2  g05481(.A(new_n5866_), .B(new_n1227_), .Y(new_n5867_));
  NOR2  g05482(.A(new_n5867_), .B(new_n1231_), .Y(new_n5868_));
  NOR2  g05483(.A(new_n5868_), .B(new_n1235_), .Y(new_n5869_));
  NOR2  g05484(.A(new_n5869_), .B(new_n1239_), .Y(new_n5870_));
  NOR2  g05485(.A(new_n5870_), .B(new_n1243_), .Y(new_n5871_));
  NOR2  g05486(.A(new_n5871_), .B(new_n1247_), .Y(new_n5872_));
  NOR2  g05487(.A(new_n5872_), .B(new_n1251_), .Y(new_n5873_));
  NOR2  g05488(.A(new_n5873_), .B(new_n1255_), .Y(new_n5874_));
  NOR2  g05489(.A(new_n5874_), .B(new_n1259_), .Y(new_n5875_));
  NOR2  g05490(.A(new_n5875_), .B(new_n1263_), .Y(new_n5876_));
  NOR2  g05491(.A(new_n5876_), .B(new_n1267_), .Y(new_n5877_));
  NOR2  g05492(.A(new_n5877_), .B(new_n1271_), .Y(new_n5878_));
  NOR2  g05493(.A(new_n5878_), .B(new_n1275_), .Y(new_n5879_));
  NOR2  g05494(.A(new_n5879_), .B(new_n1279_), .Y(new_n5880_));
  NOR2  g05495(.A(new_n5880_), .B(new_n1283_), .Y(new_n5881_));
  NOR2  g05496(.A(new_n5881_), .B(new_n1287_), .Y(new_n5882_));
  NOR2  g05497(.A(new_n5882_), .B(new_n1291_), .Y(new_n5883_));
  NOR2  g05498(.A(new_n5883_), .B(new_n1295_), .Y(new_n5884_));
  NOR2  g05499(.A(new_n5884_), .B(new_n1299_), .Y(new_n5885_));
  NOR2  g05500(.A(new_n5885_), .B(new_n1303_), .Y(new_n5886_));
  NOR2  g05501(.A(new_n5886_), .B(new_n1307_), .Y(new_n5887_));
  NOR2  g05502(.A(new_n5887_), .B(new_n1311_), .Y(new_n5888_));
  NOR2  g05503(.A(new_n5888_), .B(new_n1315_), .Y(new_n5889_));
  NOR2  g05504(.A(new_n5889_), .B(new_n1319_), .Y(new_n5890_));
  NAND2 g05505(.A(new_n1321_), .B(\req[52] ), .Y(new_n5891_));
  NOR2  g05506(.A(new_n5891_), .B(new_n5890_), .Y(\grant[52] ));
  INV   g05507(.A(new_n1330_), .Y(new_n5893_));
  NOR2  g05508(.A(new_n5893_), .B(new_n565_), .Y(new_n5894_));
  NOR2  g05509(.A(new_n5894_), .B(new_n1335_), .Y(new_n5895_));
  NOR2  g05510(.A(new_n5895_), .B(new_n1339_), .Y(new_n5896_));
  NOR2  g05511(.A(new_n5896_), .B(new_n1343_), .Y(new_n5897_));
  NOR2  g05512(.A(new_n5897_), .B(new_n1347_), .Y(new_n5898_));
  NOR2  g05513(.A(new_n5898_), .B(new_n1351_), .Y(new_n5899_));
  NOR2  g05514(.A(new_n5899_), .B(new_n1355_), .Y(new_n5900_));
  NOR2  g05515(.A(new_n5900_), .B(new_n1359_), .Y(new_n5901_));
  NOR2  g05516(.A(new_n5901_), .B(new_n1363_), .Y(new_n5902_));
  NOR2  g05517(.A(new_n5902_), .B(new_n1367_), .Y(new_n5903_));
  NOR2  g05518(.A(new_n5903_), .B(new_n1371_), .Y(new_n5904_));
  NOR2  g05519(.A(new_n5904_), .B(new_n1375_), .Y(new_n5905_));
  NOR2  g05520(.A(new_n5905_), .B(new_n1379_), .Y(new_n5906_));
  NOR2  g05521(.A(new_n5906_), .B(new_n1383_), .Y(new_n5907_));
  NOR2  g05522(.A(new_n5907_), .B(new_n1387_), .Y(new_n5908_));
  NOR2  g05523(.A(new_n5908_), .B(new_n1391_), .Y(new_n5909_));
  NOR2  g05524(.A(new_n5909_), .B(new_n1395_), .Y(new_n5910_));
  NOR2  g05525(.A(new_n5910_), .B(new_n1399_), .Y(new_n5911_));
  NOR2  g05526(.A(new_n5911_), .B(new_n1403_), .Y(new_n5912_));
  NOR2  g05527(.A(new_n5912_), .B(new_n1407_), .Y(new_n5913_));
  NOR2  g05528(.A(new_n5913_), .B(new_n1411_), .Y(new_n5914_));
  NOR2  g05529(.A(new_n5914_), .B(new_n1415_), .Y(new_n5915_));
  NOR2  g05530(.A(new_n5915_), .B(new_n1419_), .Y(new_n5916_));
  NOR2  g05531(.A(new_n5916_), .B(new_n1423_), .Y(new_n5917_));
  NOR2  g05532(.A(new_n5917_), .B(new_n1427_), .Y(new_n5918_));
  NOR2  g05533(.A(new_n5918_), .B(new_n1431_), .Y(new_n5919_));
  NOR2  g05534(.A(new_n5919_), .B(new_n1435_), .Y(new_n5920_));
  NOR2  g05535(.A(new_n5920_), .B(new_n1439_), .Y(new_n5921_));
  NOR2  g05536(.A(new_n5921_), .B(new_n1443_), .Y(new_n5922_));
  NOR2  g05537(.A(new_n5922_), .B(new_n1447_), .Y(new_n5923_));
  NOR2  g05538(.A(new_n5923_), .B(new_n1451_), .Y(new_n5924_));
  NOR2  g05539(.A(new_n5924_), .B(new_n1455_), .Y(new_n5925_));
  NOR2  g05540(.A(new_n5925_), .B(new_n1459_), .Y(new_n5926_));
  NOR2  g05541(.A(new_n5926_), .B(new_n1463_), .Y(new_n5927_));
  NOR2  g05542(.A(new_n5927_), .B(new_n1467_), .Y(new_n5928_));
  NOR2  g05543(.A(new_n5928_), .B(new_n1471_), .Y(new_n5929_));
  NOR2  g05544(.A(new_n5929_), .B(new_n1475_), .Y(new_n5930_));
  NOR2  g05545(.A(new_n5930_), .B(new_n1479_), .Y(new_n5931_));
  NOR2  g05546(.A(new_n5931_), .B(new_n1483_), .Y(new_n5932_));
  NOR2  g05547(.A(new_n5932_), .B(new_n1487_), .Y(new_n5933_));
  NOR2  g05548(.A(new_n5933_), .B(new_n1491_), .Y(new_n5934_));
  NOR2  g05549(.A(new_n5934_), .B(new_n1495_), .Y(new_n5935_));
  NOR2  g05550(.A(new_n5935_), .B(new_n1499_), .Y(new_n5936_));
  NOR2  g05551(.A(new_n5936_), .B(new_n1503_), .Y(new_n5937_));
  NOR2  g05552(.A(new_n5937_), .B(new_n1507_), .Y(new_n5938_));
  NOR2  g05553(.A(new_n5938_), .B(new_n1511_), .Y(new_n5939_));
  NOR2  g05554(.A(new_n5939_), .B(new_n1515_), .Y(new_n5940_));
  NOR2  g05555(.A(new_n5940_), .B(new_n1519_), .Y(new_n5941_));
  NOR2  g05556(.A(new_n5941_), .B(new_n1523_), .Y(new_n5942_));
  NOR2  g05557(.A(new_n5942_), .B(new_n1527_), .Y(new_n5943_));
  NOR2  g05558(.A(new_n5943_), .B(new_n1797_), .Y(new_n5944_));
  NOR2  g05559(.A(new_n5944_), .B(new_n396_), .Y(new_n5945_));
  NOR2  g05560(.A(new_n5945_), .B(new_n400_), .Y(new_n5946_));
  NOR2  g05561(.A(new_n5946_), .B(new_n406_), .Y(new_n5947_));
  NOR2  g05562(.A(new_n5947_), .B(new_n410_), .Y(new_n5948_));
  NOR2  g05563(.A(new_n5948_), .B(new_n416_), .Y(new_n5949_));
  NOR2  g05564(.A(new_n5949_), .B(new_n420_), .Y(new_n5950_));
  NOR2  g05565(.A(new_n5950_), .B(new_n426_), .Y(new_n5951_));
  NOR2  g05566(.A(new_n5951_), .B(new_n430_), .Y(new_n5952_));
  NOR2  g05567(.A(new_n5952_), .B(new_n436_), .Y(new_n5953_));
  NOR2  g05568(.A(new_n5953_), .B(new_n440_), .Y(new_n5954_));
  NOR2  g05569(.A(new_n5954_), .B(new_n446_), .Y(new_n5955_));
  NOR2  g05570(.A(new_n5955_), .B(new_n450_), .Y(new_n5956_));
  NOR2  g05571(.A(new_n5956_), .B(new_n456_), .Y(new_n5957_));
  NOR2  g05572(.A(new_n5957_), .B(new_n460_), .Y(new_n5958_));
  NOR2  g05573(.A(new_n5958_), .B(new_n466_), .Y(new_n5959_));
  NOR2  g05574(.A(new_n5959_), .B(new_n470_), .Y(new_n5960_));
  NOR2  g05575(.A(new_n5960_), .B(new_n476_), .Y(new_n5961_));
  NOR2  g05576(.A(new_n5961_), .B(new_n480_), .Y(new_n5962_));
  NOR2  g05577(.A(new_n5962_), .B(new_n486_), .Y(new_n5963_));
  NOR2  g05578(.A(new_n5963_), .B(new_n490_), .Y(new_n5964_));
  NOR2  g05579(.A(new_n5964_), .B(new_n496_), .Y(new_n5965_));
  NOR2  g05580(.A(new_n5965_), .B(new_n500_), .Y(new_n5966_));
  NOR2  g05581(.A(new_n5966_), .B(new_n506_), .Y(new_n5967_));
  NOR2  g05582(.A(new_n5967_), .B(new_n510_), .Y(new_n5968_));
  NOR2  g05583(.A(new_n5968_), .B(new_n516_), .Y(new_n5969_));
  NOR2  g05584(.A(new_n5969_), .B(new_n520_), .Y(new_n5970_));
  NOR2  g05585(.A(new_n5970_), .B(new_n526_), .Y(new_n5971_));
  NOR2  g05586(.A(new_n5971_), .B(new_n530_), .Y(new_n5972_));
  NOR2  g05587(.A(new_n5972_), .B(new_n536_), .Y(new_n5973_));
  NOR2  g05588(.A(new_n5973_), .B(new_n540_), .Y(new_n5974_));
  NOR2  g05589(.A(new_n5974_), .B(new_n546_), .Y(new_n5975_));
  NOR2  g05590(.A(new_n5975_), .B(new_n550_), .Y(new_n5976_));
  NOR2  g05591(.A(new_n5976_), .B(new_n556_), .Y(new_n5977_));
  NAND2 g05592(.A(new_n558_), .B(\req[53] ), .Y(new_n5978_));
  NOR2  g05593(.A(new_n5978_), .B(new_n5977_), .Y(\grant[53] ));
  INV   g05594(.A(new_n569_), .Y(new_n5980_));
  NOR2  g05595(.A(new_n972_), .B(new_n5980_), .Y(new_n5981_));
  NOR2  g05596(.A(new_n5981_), .B(new_n576_), .Y(new_n5982_));
  NOR2  g05597(.A(new_n5982_), .B(new_n580_), .Y(new_n5983_));
  NOR2  g05598(.A(new_n5983_), .B(new_n586_), .Y(new_n5984_));
  NOR2  g05599(.A(new_n5984_), .B(new_n590_), .Y(new_n5985_));
  NOR2  g05600(.A(new_n5985_), .B(new_n596_), .Y(new_n5986_));
  NOR2  g05601(.A(new_n5986_), .B(new_n600_), .Y(new_n5987_));
  NOR2  g05602(.A(new_n5987_), .B(new_n606_), .Y(new_n5988_));
  NOR2  g05603(.A(new_n5988_), .B(new_n610_), .Y(new_n5989_));
  NOR2  g05604(.A(new_n5989_), .B(new_n616_), .Y(new_n5990_));
  NOR2  g05605(.A(new_n5990_), .B(new_n620_), .Y(new_n5991_));
  NOR2  g05606(.A(new_n5991_), .B(new_n626_), .Y(new_n5992_));
  NOR2  g05607(.A(new_n5992_), .B(new_n630_), .Y(new_n5993_));
  NOR2  g05608(.A(new_n5993_), .B(new_n636_), .Y(new_n5994_));
  NOR2  g05609(.A(new_n5994_), .B(new_n640_), .Y(new_n5995_));
  NOR2  g05610(.A(new_n5995_), .B(new_n646_), .Y(new_n5996_));
  NOR2  g05611(.A(new_n5996_), .B(new_n650_), .Y(new_n5997_));
  NOR2  g05612(.A(new_n5997_), .B(new_n656_), .Y(new_n5998_));
  NOR2  g05613(.A(new_n5998_), .B(new_n660_), .Y(new_n5999_));
  NOR2  g05614(.A(new_n5999_), .B(new_n666_), .Y(new_n6000_));
  NOR2  g05615(.A(new_n6000_), .B(new_n670_), .Y(new_n6001_));
  NOR2  g05616(.A(new_n6001_), .B(new_n676_), .Y(new_n6002_));
  NOR2  g05617(.A(new_n6002_), .B(new_n680_), .Y(new_n6003_));
  NOR2  g05618(.A(new_n6003_), .B(new_n686_), .Y(new_n6004_));
  NOR2  g05619(.A(new_n6004_), .B(new_n690_), .Y(new_n6005_));
  NOR2  g05620(.A(new_n6005_), .B(new_n696_), .Y(new_n6006_));
  NOR2  g05621(.A(new_n6006_), .B(new_n700_), .Y(new_n6007_));
  NOR2  g05622(.A(new_n6007_), .B(new_n706_), .Y(new_n6008_));
  NOR2  g05623(.A(new_n6008_), .B(new_n710_), .Y(new_n6009_));
  NOR2  g05624(.A(new_n6009_), .B(new_n716_), .Y(new_n6010_));
  NOR2  g05625(.A(new_n6010_), .B(new_n720_), .Y(new_n6011_));
  NOR2  g05626(.A(new_n6011_), .B(new_n726_), .Y(new_n6012_));
  NOR2  g05627(.A(new_n6012_), .B(new_n730_), .Y(new_n6013_));
  NOR2  g05628(.A(new_n6013_), .B(new_n736_), .Y(new_n6014_));
  NOR2  g05629(.A(new_n6014_), .B(new_n740_), .Y(new_n6015_));
  NOR2  g05630(.A(new_n6015_), .B(new_n746_), .Y(new_n6016_));
  NOR2  g05631(.A(new_n6016_), .B(new_n750_), .Y(new_n6017_));
  NOR2  g05632(.A(new_n6017_), .B(new_n756_), .Y(new_n6018_));
  NOR2  g05633(.A(new_n6018_), .B(new_n760_), .Y(new_n6019_));
  NOR2  g05634(.A(new_n6019_), .B(new_n766_), .Y(new_n6020_));
  NOR2  g05635(.A(new_n6020_), .B(new_n770_), .Y(new_n6021_));
  NOR2  g05636(.A(new_n6021_), .B(new_n776_), .Y(new_n6022_));
  NOR2  g05637(.A(new_n6022_), .B(new_n780_), .Y(new_n6023_));
  NOR2  g05638(.A(new_n6023_), .B(new_n786_), .Y(new_n6024_));
  NOR2  g05639(.A(new_n6024_), .B(new_n790_), .Y(new_n6025_));
  NOR2  g05640(.A(new_n6025_), .B(new_n796_), .Y(new_n6026_));
  NOR2  g05641(.A(new_n6026_), .B(new_n800_), .Y(new_n6027_));
  NOR2  g05642(.A(new_n6027_), .B(new_n806_), .Y(new_n6028_));
  NOR2  g05643(.A(new_n6028_), .B(new_n1616_), .Y(new_n6029_));
  NOR2  g05644(.A(new_n6029_), .B(new_n1618_), .Y(new_n6030_));
  NOR2  g05645(.A(new_n6030_), .B(new_n1885_), .Y(new_n6031_));
  NOR2  g05646(.A(new_n6031_), .B(new_n820_), .Y(new_n6032_));
  NOR2  g05647(.A(new_n6032_), .B(new_n824_), .Y(new_n6033_));
  NOR2  g05648(.A(new_n6033_), .B(new_n829_), .Y(new_n6034_));
  NOR2  g05649(.A(new_n6034_), .B(new_n833_), .Y(new_n6035_));
  NOR2  g05650(.A(new_n6035_), .B(new_n838_), .Y(new_n6036_));
  NOR2  g05651(.A(new_n6036_), .B(new_n842_), .Y(new_n6037_));
  NOR2  g05652(.A(new_n6037_), .B(new_n847_), .Y(new_n6038_));
  NOR2  g05653(.A(new_n6038_), .B(new_n851_), .Y(new_n6039_));
  NOR2  g05654(.A(new_n6039_), .B(new_n856_), .Y(new_n6040_));
  NOR2  g05655(.A(new_n6040_), .B(new_n860_), .Y(new_n6041_));
  NOR2  g05656(.A(new_n6041_), .B(new_n865_), .Y(new_n6042_));
  NOR2  g05657(.A(new_n6042_), .B(new_n869_), .Y(new_n6043_));
  NOR2  g05658(.A(new_n6043_), .B(new_n874_), .Y(new_n6044_));
  NOR2  g05659(.A(new_n6044_), .B(new_n878_), .Y(new_n6045_));
  NOR2  g05660(.A(new_n6045_), .B(new_n883_), .Y(new_n6046_));
  NOR2  g05661(.A(new_n6046_), .B(new_n887_), .Y(new_n6047_));
  NOR2  g05662(.A(new_n6047_), .B(new_n892_), .Y(new_n6048_));
  NOR2  g05663(.A(new_n6048_), .B(new_n896_), .Y(new_n6049_));
  NOR2  g05664(.A(new_n6049_), .B(new_n901_), .Y(new_n6050_));
  NOR2  g05665(.A(new_n6050_), .B(new_n905_), .Y(new_n6051_));
  NOR2  g05666(.A(new_n6051_), .B(new_n910_), .Y(new_n6052_));
  NOR2  g05667(.A(new_n6052_), .B(new_n914_), .Y(new_n6053_));
  NOR2  g05668(.A(new_n6053_), .B(new_n919_), .Y(new_n6054_));
  NOR2  g05669(.A(new_n6054_), .B(new_n923_), .Y(new_n6055_));
  NOR2  g05670(.A(new_n6055_), .B(new_n928_), .Y(new_n6056_));
  NOR2  g05671(.A(new_n6056_), .B(new_n932_), .Y(new_n6057_));
  NOR2  g05672(.A(new_n6057_), .B(new_n937_), .Y(new_n6058_));
  NOR2  g05673(.A(new_n6058_), .B(new_n941_), .Y(new_n6059_));
  NOR2  g05674(.A(new_n6059_), .B(new_n946_), .Y(new_n6060_));
  NOR2  g05675(.A(new_n6060_), .B(new_n950_), .Y(new_n6061_));
  NOR2  g05676(.A(new_n6061_), .B(new_n955_), .Y(new_n6062_));
  NOR2  g05677(.A(new_n6062_), .B(new_n959_), .Y(new_n6063_));
  NOR2  g05678(.A(new_n6063_), .B(new_n964_), .Y(new_n6064_));
  NAND2 g05679(.A(new_n966_), .B(\req[54] ), .Y(new_n6065_));
  NOR2  g05680(.A(new_n6065_), .B(new_n6064_), .Y(\grant[54] ));
  INV   g05681(.A(new_n976_), .Y(new_n6067_));
  NOR2  g05682(.A(new_n1334_), .B(new_n6067_), .Y(new_n6068_));
  NOR2  g05683(.A(new_n6068_), .B(new_n982_), .Y(new_n6069_));
  NOR2  g05684(.A(new_n6069_), .B(new_n986_), .Y(new_n6070_));
  NOR2  g05685(.A(new_n6070_), .B(new_n991_), .Y(new_n6071_));
  NOR2  g05686(.A(new_n6071_), .B(new_n995_), .Y(new_n6072_));
  NOR2  g05687(.A(new_n6072_), .B(new_n1000_), .Y(new_n6073_));
  NOR2  g05688(.A(new_n6073_), .B(new_n1004_), .Y(new_n6074_));
  NOR2  g05689(.A(new_n6074_), .B(new_n1009_), .Y(new_n6075_));
  NOR2  g05690(.A(new_n6075_), .B(new_n1013_), .Y(new_n6076_));
  NOR2  g05691(.A(new_n6076_), .B(new_n1018_), .Y(new_n6077_));
  NOR2  g05692(.A(new_n6077_), .B(new_n1022_), .Y(new_n6078_));
  NOR2  g05693(.A(new_n6078_), .B(new_n1027_), .Y(new_n6079_));
  NOR2  g05694(.A(new_n6079_), .B(new_n1031_), .Y(new_n6080_));
  NOR2  g05695(.A(new_n6080_), .B(new_n1036_), .Y(new_n6081_));
  NOR2  g05696(.A(new_n6081_), .B(new_n1040_), .Y(new_n6082_));
  NOR2  g05697(.A(new_n6082_), .B(new_n1045_), .Y(new_n6083_));
  NOR2  g05698(.A(new_n6083_), .B(new_n1049_), .Y(new_n6084_));
  NOR2  g05699(.A(new_n6084_), .B(new_n1054_), .Y(new_n6085_));
  NOR2  g05700(.A(new_n6085_), .B(new_n1058_), .Y(new_n6086_));
  NOR2  g05701(.A(new_n6086_), .B(new_n1063_), .Y(new_n6087_));
  NOR2  g05702(.A(new_n6087_), .B(new_n1067_), .Y(new_n6088_));
  NOR2  g05703(.A(new_n6088_), .B(new_n1072_), .Y(new_n6089_));
  NOR2  g05704(.A(new_n6089_), .B(new_n1076_), .Y(new_n6090_));
  NOR2  g05705(.A(new_n6090_), .B(new_n1081_), .Y(new_n6091_));
  NOR2  g05706(.A(new_n6091_), .B(new_n1085_), .Y(new_n6092_));
  NOR2  g05707(.A(new_n6092_), .B(new_n1090_), .Y(new_n6093_));
  NOR2  g05708(.A(new_n6093_), .B(new_n1094_), .Y(new_n6094_));
  NOR2  g05709(.A(new_n6094_), .B(new_n1099_), .Y(new_n6095_));
  NOR2  g05710(.A(new_n6095_), .B(new_n1103_), .Y(new_n6096_));
  NOR2  g05711(.A(new_n6096_), .B(new_n1108_), .Y(new_n6097_));
  NOR2  g05712(.A(new_n6097_), .B(new_n1112_), .Y(new_n6098_));
  NOR2  g05713(.A(new_n6098_), .B(new_n1117_), .Y(new_n6099_));
  NOR2  g05714(.A(new_n6099_), .B(new_n1121_), .Y(new_n6100_));
  NOR2  g05715(.A(new_n6100_), .B(new_n1126_), .Y(new_n6101_));
  NOR2  g05716(.A(new_n6101_), .B(new_n1130_), .Y(new_n6102_));
  NOR2  g05717(.A(new_n6102_), .B(new_n1135_), .Y(new_n6103_));
  NOR2  g05718(.A(new_n6103_), .B(new_n1139_), .Y(new_n6104_));
  NOR2  g05719(.A(new_n6104_), .B(new_n1144_), .Y(new_n6105_));
  NOR2  g05720(.A(new_n6105_), .B(new_n1148_), .Y(new_n6106_));
  NOR2  g05721(.A(new_n6106_), .B(new_n1153_), .Y(new_n6107_));
  NOR2  g05722(.A(new_n6107_), .B(new_n1157_), .Y(new_n6108_));
  NOR2  g05723(.A(new_n6108_), .B(new_n1162_), .Y(new_n6109_));
  NOR2  g05724(.A(new_n6109_), .B(new_n1166_), .Y(new_n6110_));
  NOR2  g05725(.A(new_n6110_), .B(new_n1171_), .Y(new_n6111_));
  NOR2  g05726(.A(new_n6111_), .B(new_n1175_), .Y(new_n6112_));
  NOR2  g05727(.A(new_n6112_), .B(new_n1180_), .Y(new_n6113_));
  NOR2  g05728(.A(new_n6113_), .B(new_n1184_), .Y(new_n6114_));
  NOR2  g05729(.A(new_n6114_), .B(new_n1189_), .Y(new_n6115_));
  NOR2  g05730(.A(new_n6115_), .B(new_n1707_), .Y(new_n6116_));
  NOR2  g05731(.A(new_n6116_), .B(new_n1709_), .Y(new_n6117_));
  NOR2  g05732(.A(new_n6117_), .B(new_n1973_), .Y(new_n6118_));
  NOR2  g05733(.A(new_n6118_), .B(new_n1199_), .Y(new_n6119_));
  NOR2  g05734(.A(new_n6119_), .B(new_n1203_), .Y(new_n6120_));
  NOR2  g05735(.A(new_n6120_), .B(new_n1207_), .Y(new_n6121_));
  NOR2  g05736(.A(new_n6121_), .B(new_n1211_), .Y(new_n6122_));
  NOR2  g05737(.A(new_n6122_), .B(new_n1215_), .Y(new_n6123_));
  NOR2  g05738(.A(new_n6123_), .B(new_n1219_), .Y(new_n6124_));
  NOR2  g05739(.A(new_n6124_), .B(new_n1223_), .Y(new_n6125_));
  NOR2  g05740(.A(new_n6125_), .B(new_n1227_), .Y(new_n6126_));
  NOR2  g05741(.A(new_n6126_), .B(new_n1231_), .Y(new_n6127_));
  NOR2  g05742(.A(new_n6127_), .B(new_n1235_), .Y(new_n6128_));
  NOR2  g05743(.A(new_n6128_), .B(new_n1239_), .Y(new_n6129_));
  NOR2  g05744(.A(new_n6129_), .B(new_n1243_), .Y(new_n6130_));
  NOR2  g05745(.A(new_n6130_), .B(new_n1247_), .Y(new_n6131_));
  NOR2  g05746(.A(new_n6131_), .B(new_n1251_), .Y(new_n6132_));
  NOR2  g05747(.A(new_n6132_), .B(new_n1255_), .Y(new_n6133_));
  NOR2  g05748(.A(new_n6133_), .B(new_n1259_), .Y(new_n6134_));
  NOR2  g05749(.A(new_n6134_), .B(new_n1263_), .Y(new_n6135_));
  NOR2  g05750(.A(new_n6135_), .B(new_n1267_), .Y(new_n6136_));
  NOR2  g05751(.A(new_n6136_), .B(new_n1271_), .Y(new_n6137_));
  NOR2  g05752(.A(new_n6137_), .B(new_n1275_), .Y(new_n6138_));
  NOR2  g05753(.A(new_n6138_), .B(new_n1279_), .Y(new_n6139_));
  NOR2  g05754(.A(new_n6139_), .B(new_n1283_), .Y(new_n6140_));
  NOR2  g05755(.A(new_n6140_), .B(new_n1287_), .Y(new_n6141_));
  NOR2  g05756(.A(new_n6141_), .B(new_n1291_), .Y(new_n6142_));
  NOR2  g05757(.A(new_n6142_), .B(new_n1295_), .Y(new_n6143_));
  NOR2  g05758(.A(new_n6143_), .B(new_n1299_), .Y(new_n6144_));
  NOR2  g05759(.A(new_n6144_), .B(new_n1303_), .Y(new_n6145_));
  NOR2  g05760(.A(new_n6145_), .B(new_n1307_), .Y(new_n6146_));
  NOR2  g05761(.A(new_n6146_), .B(new_n1311_), .Y(new_n6147_));
  NOR2  g05762(.A(new_n6147_), .B(new_n1315_), .Y(new_n6148_));
  NOR2  g05763(.A(new_n6148_), .B(new_n1319_), .Y(new_n6149_));
  NOR2  g05764(.A(new_n6149_), .B(new_n1323_), .Y(new_n6150_));
  NOR2  g05765(.A(new_n6150_), .B(new_n1327_), .Y(new_n6151_));
  NAND2 g05766(.A(new_n1329_), .B(\req[55] ), .Y(new_n6152_));
  NOR2  g05767(.A(new_n6152_), .B(new_n6151_), .Y(\grant[55] ));
  INV   g05768(.A(new_n1338_), .Y(new_n6154_));
  NOR2  g05769(.A(new_n6154_), .B(new_n575_), .Y(new_n6155_));
  NOR2  g05770(.A(new_n6155_), .B(new_n1343_), .Y(new_n6156_));
  NOR2  g05771(.A(new_n6156_), .B(new_n1347_), .Y(new_n6157_));
  NOR2  g05772(.A(new_n6157_), .B(new_n1351_), .Y(new_n6158_));
  NOR2  g05773(.A(new_n6158_), .B(new_n1355_), .Y(new_n6159_));
  NOR2  g05774(.A(new_n6159_), .B(new_n1359_), .Y(new_n6160_));
  NOR2  g05775(.A(new_n6160_), .B(new_n1363_), .Y(new_n6161_));
  NOR2  g05776(.A(new_n6161_), .B(new_n1367_), .Y(new_n6162_));
  NOR2  g05777(.A(new_n6162_), .B(new_n1371_), .Y(new_n6163_));
  NOR2  g05778(.A(new_n6163_), .B(new_n1375_), .Y(new_n6164_));
  NOR2  g05779(.A(new_n6164_), .B(new_n1379_), .Y(new_n6165_));
  NOR2  g05780(.A(new_n6165_), .B(new_n1383_), .Y(new_n6166_));
  NOR2  g05781(.A(new_n6166_), .B(new_n1387_), .Y(new_n6167_));
  NOR2  g05782(.A(new_n6167_), .B(new_n1391_), .Y(new_n6168_));
  NOR2  g05783(.A(new_n6168_), .B(new_n1395_), .Y(new_n6169_));
  NOR2  g05784(.A(new_n6169_), .B(new_n1399_), .Y(new_n6170_));
  NOR2  g05785(.A(new_n6170_), .B(new_n1403_), .Y(new_n6171_));
  NOR2  g05786(.A(new_n6171_), .B(new_n1407_), .Y(new_n6172_));
  NOR2  g05787(.A(new_n6172_), .B(new_n1411_), .Y(new_n6173_));
  NOR2  g05788(.A(new_n6173_), .B(new_n1415_), .Y(new_n6174_));
  NOR2  g05789(.A(new_n6174_), .B(new_n1419_), .Y(new_n6175_));
  NOR2  g05790(.A(new_n6175_), .B(new_n1423_), .Y(new_n6176_));
  NOR2  g05791(.A(new_n6176_), .B(new_n1427_), .Y(new_n6177_));
  NOR2  g05792(.A(new_n6177_), .B(new_n1431_), .Y(new_n6178_));
  NOR2  g05793(.A(new_n6178_), .B(new_n1435_), .Y(new_n6179_));
  NOR2  g05794(.A(new_n6179_), .B(new_n1439_), .Y(new_n6180_));
  NOR2  g05795(.A(new_n6180_), .B(new_n1443_), .Y(new_n6181_));
  NOR2  g05796(.A(new_n6181_), .B(new_n1447_), .Y(new_n6182_));
  NOR2  g05797(.A(new_n6182_), .B(new_n1451_), .Y(new_n6183_));
  NOR2  g05798(.A(new_n6183_), .B(new_n1455_), .Y(new_n6184_));
  NOR2  g05799(.A(new_n6184_), .B(new_n1459_), .Y(new_n6185_));
  NOR2  g05800(.A(new_n6185_), .B(new_n1463_), .Y(new_n6186_));
  NOR2  g05801(.A(new_n6186_), .B(new_n1467_), .Y(new_n6187_));
  NOR2  g05802(.A(new_n6187_), .B(new_n1471_), .Y(new_n6188_));
  NOR2  g05803(.A(new_n6188_), .B(new_n1475_), .Y(new_n6189_));
  NOR2  g05804(.A(new_n6189_), .B(new_n1479_), .Y(new_n6190_));
  NOR2  g05805(.A(new_n6190_), .B(new_n1483_), .Y(new_n6191_));
  NOR2  g05806(.A(new_n6191_), .B(new_n1487_), .Y(new_n6192_));
  NOR2  g05807(.A(new_n6192_), .B(new_n1491_), .Y(new_n6193_));
  NOR2  g05808(.A(new_n6193_), .B(new_n1495_), .Y(new_n6194_));
  NOR2  g05809(.A(new_n6194_), .B(new_n1499_), .Y(new_n6195_));
  NOR2  g05810(.A(new_n6195_), .B(new_n1503_), .Y(new_n6196_));
  NOR2  g05811(.A(new_n6196_), .B(new_n1507_), .Y(new_n6197_));
  NOR2  g05812(.A(new_n6197_), .B(new_n1511_), .Y(new_n6198_));
  NOR2  g05813(.A(new_n6198_), .B(new_n1515_), .Y(new_n6199_));
  NOR2  g05814(.A(new_n6199_), .B(new_n1519_), .Y(new_n6200_));
  NOR2  g05815(.A(new_n6200_), .B(new_n1523_), .Y(new_n6201_));
  NOR2  g05816(.A(new_n6201_), .B(new_n1527_), .Y(new_n6202_));
  NOR2  g05817(.A(new_n6202_), .B(new_n1797_), .Y(new_n6203_));
  NOR2  g05818(.A(new_n6203_), .B(new_n396_), .Y(new_n6204_));
  NOR2  g05819(.A(new_n6204_), .B(new_n400_), .Y(new_n6205_));
  NOR2  g05820(.A(new_n6205_), .B(new_n406_), .Y(new_n6206_));
  NOR2  g05821(.A(new_n6206_), .B(new_n410_), .Y(new_n6207_));
  NOR2  g05822(.A(new_n6207_), .B(new_n416_), .Y(new_n6208_));
  NOR2  g05823(.A(new_n6208_), .B(new_n420_), .Y(new_n6209_));
  NOR2  g05824(.A(new_n6209_), .B(new_n426_), .Y(new_n6210_));
  NOR2  g05825(.A(new_n6210_), .B(new_n430_), .Y(new_n6211_));
  NOR2  g05826(.A(new_n6211_), .B(new_n436_), .Y(new_n6212_));
  NOR2  g05827(.A(new_n6212_), .B(new_n440_), .Y(new_n6213_));
  NOR2  g05828(.A(new_n6213_), .B(new_n446_), .Y(new_n6214_));
  NOR2  g05829(.A(new_n6214_), .B(new_n450_), .Y(new_n6215_));
  NOR2  g05830(.A(new_n6215_), .B(new_n456_), .Y(new_n6216_));
  NOR2  g05831(.A(new_n6216_), .B(new_n460_), .Y(new_n6217_));
  NOR2  g05832(.A(new_n6217_), .B(new_n466_), .Y(new_n6218_));
  NOR2  g05833(.A(new_n6218_), .B(new_n470_), .Y(new_n6219_));
  NOR2  g05834(.A(new_n6219_), .B(new_n476_), .Y(new_n6220_));
  NOR2  g05835(.A(new_n6220_), .B(new_n480_), .Y(new_n6221_));
  NOR2  g05836(.A(new_n6221_), .B(new_n486_), .Y(new_n6222_));
  NOR2  g05837(.A(new_n6222_), .B(new_n490_), .Y(new_n6223_));
  NOR2  g05838(.A(new_n6223_), .B(new_n496_), .Y(new_n6224_));
  NOR2  g05839(.A(new_n6224_), .B(new_n500_), .Y(new_n6225_));
  NOR2  g05840(.A(new_n6225_), .B(new_n506_), .Y(new_n6226_));
  NOR2  g05841(.A(new_n6226_), .B(new_n510_), .Y(new_n6227_));
  NOR2  g05842(.A(new_n6227_), .B(new_n516_), .Y(new_n6228_));
  NOR2  g05843(.A(new_n6228_), .B(new_n520_), .Y(new_n6229_));
  NOR2  g05844(.A(new_n6229_), .B(new_n526_), .Y(new_n6230_));
  NOR2  g05845(.A(new_n6230_), .B(new_n530_), .Y(new_n6231_));
  NOR2  g05846(.A(new_n6231_), .B(new_n536_), .Y(new_n6232_));
  NOR2  g05847(.A(new_n6232_), .B(new_n540_), .Y(new_n6233_));
  NOR2  g05848(.A(new_n6233_), .B(new_n546_), .Y(new_n6234_));
  NOR2  g05849(.A(new_n6234_), .B(new_n550_), .Y(new_n6235_));
  NOR2  g05850(.A(new_n6235_), .B(new_n556_), .Y(new_n6236_));
  NOR2  g05851(.A(new_n6236_), .B(new_n560_), .Y(new_n6237_));
  NOR2  g05852(.A(new_n6237_), .B(new_n566_), .Y(new_n6238_));
  NAND2 g05853(.A(new_n568_), .B(\req[56] ), .Y(new_n6239_));
  NOR2  g05854(.A(new_n6239_), .B(new_n6238_), .Y(\grant[56] ));
  INV   g05855(.A(new_n579_), .Y(new_n6241_));
  NOR2  g05856(.A(new_n981_), .B(new_n6241_), .Y(new_n6242_));
  NOR2  g05857(.A(new_n6242_), .B(new_n586_), .Y(new_n6243_));
  NOR2  g05858(.A(new_n6243_), .B(new_n590_), .Y(new_n6244_));
  NOR2  g05859(.A(new_n6244_), .B(new_n596_), .Y(new_n6245_));
  NOR2  g05860(.A(new_n6245_), .B(new_n600_), .Y(new_n6246_));
  NOR2  g05861(.A(new_n6246_), .B(new_n606_), .Y(new_n6247_));
  NOR2  g05862(.A(new_n6247_), .B(new_n610_), .Y(new_n6248_));
  NOR2  g05863(.A(new_n6248_), .B(new_n616_), .Y(new_n6249_));
  NOR2  g05864(.A(new_n6249_), .B(new_n620_), .Y(new_n6250_));
  NOR2  g05865(.A(new_n6250_), .B(new_n626_), .Y(new_n6251_));
  NOR2  g05866(.A(new_n6251_), .B(new_n630_), .Y(new_n6252_));
  NOR2  g05867(.A(new_n6252_), .B(new_n636_), .Y(new_n6253_));
  NOR2  g05868(.A(new_n6253_), .B(new_n640_), .Y(new_n6254_));
  NOR2  g05869(.A(new_n6254_), .B(new_n646_), .Y(new_n6255_));
  NOR2  g05870(.A(new_n6255_), .B(new_n650_), .Y(new_n6256_));
  NOR2  g05871(.A(new_n6256_), .B(new_n656_), .Y(new_n6257_));
  NOR2  g05872(.A(new_n6257_), .B(new_n660_), .Y(new_n6258_));
  NOR2  g05873(.A(new_n6258_), .B(new_n666_), .Y(new_n6259_));
  NOR2  g05874(.A(new_n6259_), .B(new_n670_), .Y(new_n6260_));
  NOR2  g05875(.A(new_n6260_), .B(new_n676_), .Y(new_n6261_));
  NOR2  g05876(.A(new_n6261_), .B(new_n680_), .Y(new_n6262_));
  NOR2  g05877(.A(new_n6262_), .B(new_n686_), .Y(new_n6263_));
  NOR2  g05878(.A(new_n6263_), .B(new_n690_), .Y(new_n6264_));
  NOR2  g05879(.A(new_n6264_), .B(new_n696_), .Y(new_n6265_));
  NOR2  g05880(.A(new_n6265_), .B(new_n700_), .Y(new_n6266_));
  NOR2  g05881(.A(new_n6266_), .B(new_n706_), .Y(new_n6267_));
  NOR2  g05882(.A(new_n6267_), .B(new_n710_), .Y(new_n6268_));
  NOR2  g05883(.A(new_n6268_), .B(new_n716_), .Y(new_n6269_));
  NOR2  g05884(.A(new_n6269_), .B(new_n720_), .Y(new_n6270_));
  NOR2  g05885(.A(new_n6270_), .B(new_n726_), .Y(new_n6271_));
  NOR2  g05886(.A(new_n6271_), .B(new_n730_), .Y(new_n6272_));
  NOR2  g05887(.A(new_n6272_), .B(new_n736_), .Y(new_n6273_));
  NOR2  g05888(.A(new_n6273_), .B(new_n740_), .Y(new_n6274_));
  NOR2  g05889(.A(new_n6274_), .B(new_n746_), .Y(new_n6275_));
  NOR2  g05890(.A(new_n6275_), .B(new_n750_), .Y(new_n6276_));
  NOR2  g05891(.A(new_n6276_), .B(new_n756_), .Y(new_n6277_));
  NOR2  g05892(.A(new_n6277_), .B(new_n760_), .Y(new_n6278_));
  NOR2  g05893(.A(new_n6278_), .B(new_n766_), .Y(new_n6279_));
  NOR2  g05894(.A(new_n6279_), .B(new_n770_), .Y(new_n6280_));
  NOR2  g05895(.A(new_n6280_), .B(new_n776_), .Y(new_n6281_));
  NOR2  g05896(.A(new_n6281_), .B(new_n780_), .Y(new_n6282_));
  NOR2  g05897(.A(new_n6282_), .B(new_n786_), .Y(new_n6283_));
  NOR2  g05898(.A(new_n6283_), .B(new_n790_), .Y(new_n6284_));
  NOR2  g05899(.A(new_n6284_), .B(new_n796_), .Y(new_n6285_));
  NOR2  g05900(.A(new_n6285_), .B(new_n800_), .Y(new_n6286_));
  NOR2  g05901(.A(new_n6286_), .B(new_n806_), .Y(new_n6287_));
  NOR2  g05902(.A(new_n6287_), .B(new_n1616_), .Y(new_n6288_));
  NOR2  g05903(.A(new_n6288_), .B(new_n1618_), .Y(new_n6289_));
  NOR2  g05904(.A(new_n6289_), .B(new_n1885_), .Y(new_n6290_));
  NOR2  g05905(.A(new_n6290_), .B(new_n820_), .Y(new_n6291_));
  NOR2  g05906(.A(new_n6291_), .B(new_n824_), .Y(new_n6292_));
  NOR2  g05907(.A(new_n6292_), .B(new_n829_), .Y(new_n6293_));
  NOR2  g05908(.A(new_n6293_), .B(new_n833_), .Y(new_n6294_));
  NOR2  g05909(.A(new_n6294_), .B(new_n838_), .Y(new_n6295_));
  NOR2  g05910(.A(new_n6295_), .B(new_n842_), .Y(new_n6296_));
  NOR2  g05911(.A(new_n6296_), .B(new_n847_), .Y(new_n6297_));
  NOR2  g05912(.A(new_n6297_), .B(new_n851_), .Y(new_n6298_));
  NOR2  g05913(.A(new_n6298_), .B(new_n856_), .Y(new_n6299_));
  NOR2  g05914(.A(new_n6299_), .B(new_n860_), .Y(new_n6300_));
  NOR2  g05915(.A(new_n6300_), .B(new_n865_), .Y(new_n6301_));
  NOR2  g05916(.A(new_n6301_), .B(new_n869_), .Y(new_n6302_));
  NOR2  g05917(.A(new_n6302_), .B(new_n874_), .Y(new_n6303_));
  NOR2  g05918(.A(new_n6303_), .B(new_n878_), .Y(new_n6304_));
  NOR2  g05919(.A(new_n6304_), .B(new_n883_), .Y(new_n6305_));
  NOR2  g05920(.A(new_n6305_), .B(new_n887_), .Y(new_n6306_));
  NOR2  g05921(.A(new_n6306_), .B(new_n892_), .Y(new_n6307_));
  NOR2  g05922(.A(new_n6307_), .B(new_n896_), .Y(new_n6308_));
  NOR2  g05923(.A(new_n6308_), .B(new_n901_), .Y(new_n6309_));
  NOR2  g05924(.A(new_n6309_), .B(new_n905_), .Y(new_n6310_));
  NOR2  g05925(.A(new_n6310_), .B(new_n910_), .Y(new_n6311_));
  NOR2  g05926(.A(new_n6311_), .B(new_n914_), .Y(new_n6312_));
  NOR2  g05927(.A(new_n6312_), .B(new_n919_), .Y(new_n6313_));
  NOR2  g05928(.A(new_n6313_), .B(new_n923_), .Y(new_n6314_));
  NOR2  g05929(.A(new_n6314_), .B(new_n928_), .Y(new_n6315_));
  NOR2  g05930(.A(new_n6315_), .B(new_n932_), .Y(new_n6316_));
  NOR2  g05931(.A(new_n6316_), .B(new_n937_), .Y(new_n6317_));
  NOR2  g05932(.A(new_n6317_), .B(new_n941_), .Y(new_n6318_));
  NOR2  g05933(.A(new_n6318_), .B(new_n946_), .Y(new_n6319_));
  NOR2  g05934(.A(new_n6319_), .B(new_n950_), .Y(new_n6320_));
  NOR2  g05935(.A(new_n6320_), .B(new_n955_), .Y(new_n6321_));
  NOR2  g05936(.A(new_n6321_), .B(new_n959_), .Y(new_n6322_));
  NOR2  g05937(.A(new_n6322_), .B(new_n964_), .Y(new_n6323_));
  NOR2  g05938(.A(new_n6323_), .B(new_n968_), .Y(new_n6324_));
  NOR2  g05939(.A(new_n6324_), .B(new_n973_), .Y(new_n6325_));
  NAND2 g05940(.A(new_n975_), .B(\req[57] ), .Y(new_n6326_));
  NOR2  g05941(.A(new_n6326_), .B(new_n6325_), .Y(\grant[57] ));
  INV   g05942(.A(new_n985_), .Y(new_n6328_));
  NOR2  g05943(.A(new_n1342_), .B(new_n6328_), .Y(new_n6329_));
  NOR2  g05944(.A(new_n6329_), .B(new_n991_), .Y(new_n6330_));
  NOR2  g05945(.A(new_n6330_), .B(new_n995_), .Y(new_n6331_));
  NOR2  g05946(.A(new_n6331_), .B(new_n1000_), .Y(new_n6332_));
  NOR2  g05947(.A(new_n6332_), .B(new_n1004_), .Y(new_n6333_));
  NOR2  g05948(.A(new_n6333_), .B(new_n1009_), .Y(new_n6334_));
  NOR2  g05949(.A(new_n6334_), .B(new_n1013_), .Y(new_n6335_));
  NOR2  g05950(.A(new_n6335_), .B(new_n1018_), .Y(new_n6336_));
  NOR2  g05951(.A(new_n6336_), .B(new_n1022_), .Y(new_n6337_));
  NOR2  g05952(.A(new_n6337_), .B(new_n1027_), .Y(new_n6338_));
  NOR2  g05953(.A(new_n6338_), .B(new_n1031_), .Y(new_n6339_));
  NOR2  g05954(.A(new_n6339_), .B(new_n1036_), .Y(new_n6340_));
  NOR2  g05955(.A(new_n6340_), .B(new_n1040_), .Y(new_n6341_));
  NOR2  g05956(.A(new_n6341_), .B(new_n1045_), .Y(new_n6342_));
  NOR2  g05957(.A(new_n6342_), .B(new_n1049_), .Y(new_n6343_));
  NOR2  g05958(.A(new_n6343_), .B(new_n1054_), .Y(new_n6344_));
  NOR2  g05959(.A(new_n6344_), .B(new_n1058_), .Y(new_n6345_));
  NOR2  g05960(.A(new_n6345_), .B(new_n1063_), .Y(new_n6346_));
  NOR2  g05961(.A(new_n6346_), .B(new_n1067_), .Y(new_n6347_));
  NOR2  g05962(.A(new_n6347_), .B(new_n1072_), .Y(new_n6348_));
  NOR2  g05963(.A(new_n6348_), .B(new_n1076_), .Y(new_n6349_));
  NOR2  g05964(.A(new_n6349_), .B(new_n1081_), .Y(new_n6350_));
  NOR2  g05965(.A(new_n6350_), .B(new_n1085_), .Y(new_n6351_));
  NOR2  g05966(.A(new_n6351_), .B(new_n1090_), .Y(new_n6352_));
  NOR2  g05967(.A(new_n6352_), .B(new_n1094_), .Y(new_n6353_));
  NOR2  g05968(.A(new_n6353_), .B(new_n1099_), .Y(new_n6354_));
  NOR2  g05969(.A(new_n6354_), .B(new_n1103_), .Y(new_n6355_));
  NOR2  g05970(.A(new_n6355_), .B(new_n1108_), .Y(new_n6356_));
  NOR2  g05971(.A(new_n6356_), .B(new_n1112_), .Y(new_n6357_));
  NOR2  g05972(.A(new_n6357_), .B(new_n1117_), .Y(new_n6358_));
  NOR2  g05973(.A(new_n6358_), .B(new_n1121_), .Y(new_n6359_));
  NOR2  g05974(.A(new_n6359_), .B(new_n1126_), .Y(new_n6360_));
  NOR2  g05975(.A(new_n6360_), .B(new_n1130_), .Y(new_n6361_));
  NOR2  g05976(.A(new_n6361_), .B(new_n1135_), .Y(new_n6362_));
  NOR2  g05977(.A(new_n6362_), .B(new_n1139_), .Y(new_n6363_));
  NOR2  g05978(.A(new_n6363_), .B(new_n1144_), .Y(new_n6364_));
  NOR2  g05979(.A(new_n6364_), .B(new_n1148_), .Y(new_n6365_));
  NOR2  g05980(.A(new_n6365_), .B(new_n1153_), .Y(new_n6366_));
  NOR2  g05981(.A(new_n6366_), .B(new_n1157_), .Y(new_n6367_));
  NOR2  g05982(.A(new_n6367_), .B(new_n1162_), .Y(new_n6368_));
  NOR2  g05983(.A(new_n6368_), .B(new_n1166_), .Y(new_n6369_));
  NOR2  g05984(.A(new_n6369_), .B(new_n1171_), .Y(new_n6370_));
  NOR2  g05985(.A(new_n6370_), .B(new_n1175_), .Y(new_n6371_));
  NOR2  g05986(.A(new_n6371_), .B(new_n1180_), .Y(new_n6372_));
  NOR2  g05987(.A(new_n6372_), .B(new_n1184_), .Y(new_n6373_));
  NOR2  g05988(.A(new_n6373_), .B(new_n1189_), .Y(new_n6374_));
  NOR2  g05989(.A(new_n6374_), .B(new_n1707_), .Y(new_n6375_));
  NOR2  g05990(.A(new_n6375_), .B(new_n1709_), .Y(new_n6376_));
  NOR2  g05991(.A(new_n6376_), .B(new_n1973_), .Y(new_n6377_));
  NOR2  g05992(.A(new_n6377_), .B(new_n1199_), .Y(new_n6378_));
  NOR2  g05993(.A(new_n6378_), .B(new_n1203_), .Y(new_n6379_));
  NOR2  g05994(.A(new_n6379_), .B(new_n1207_), .Y(new_n6380_));
  NOR2  g05995(.A(new_n6380_), .B(new_n1211_), .Y(new_n6381_));
  NOR2  g05996(.A(new_n6381_), .B(new_n1215_), .Y(new_n6382_));
  NOR2  g05997(.A(new_n6382_), .B(new_n1219_), .Y(new_n6383_));
  NOR2  g05998(.A(new_n6383_), .B(new_n1223_), .Y(new_n6384_));
  NOR2  g05999(.A(new_n6384_), .B(new_n1227_), .Y(new_n6385_));
  NOR2  g06000(.A(new_n6385_), .B(new_n1231_), .Y(new_n6386_));
  NOR2  g06001(.A(new_n6386_), .B(new_n1235_), .Y(new_n6387_));
  NOR2  g06002(.A(new_n6387_), .B(new_n1239_), .Y(new_n6388_));
  NOR2  g06003(.A(new_n6388_), .B(new_n1243_), .Y(new_n6389_));
  NOR2  g06004(.A(new_n6389_), .B(new_n1247_), .Y(new_n6390_));
  NOR2  g06005(.A(new_n6390_), .B(new_n1251_), .Y(new_n6391_));
  NOR2  g06006(.A(new_n6391_), .B(new_n1255_), .Y(new_n6392_));
  NOR2  g06007(.A(new_n6392_), .B(new_n1259_), .Y(new_n6393_));
  NOR2  g06008(.A(new_n6393_), .B(new_n1263_), .Y(new_n6394_));
  NOR2  g06009(.A(new_n6394_), .B(new_n1267_), .Y(new_n6395_));
  NOR2  g06010(.A(new_n6395_), .B(new_n1271_), .Y(new_n6396_));
  NOR2  g06011(.A(new_n6396_), .B(new_n1275_), .Y(new_n6397_));
  NOR2  g06012(.A(new_n6397_), .B(new_n1279_), .Y(new_n6398_));
  NOR2  g06013(.A(new_n6398_), .B(new_n1283_), .Y(new_n6399_));
  NOR2  g06014(.A(new_n6399_), .B(new_n1287_), .Y(new_n6400_));
  NOR2  g06015(.A(new_n6400_), .B(new_n1291_), .Y(new_n6401_));
  NOR2  g06016(.A(new_n6401_), .B(new_n1295_), .Y(new_n6402_));
  NOR2  g06017(.A(new_n6402_), .B(new_n1299_), .Y(new_n6403_));
  NOR2  g06018(.A(new_n6403_), .B(new_n1303_), .Y(new_n6404_));
  NOR2  g06019(.A(new_n6404_), .B(new_n1307_), .Y(new_n6405_));
  NOR2  g06020(.A(new_n6405_), .B(new_n1311_), .Y(new_n6406_));
  NOR2  g06021(.A(new_n6406_), .B(new_n1315_), .Y(new_n6407_));
  NOR2  g06022(.A(new_n6407_), .B(new_n1319_), .Y(new_n6408_));
  NOR2  g06023(.A(new_n6408_), .B(new_n1323_), .Y(new_n6409_));
  NOR2  g06024(.A(new_n6409_), .B(new_n1327_), .Y(new_n6410_));
  NOR2  g06025(.A(new_n6410_), .B(new_n1331_), .Y(new_n6411_));
  NOR2  g06026(.A(new_n6411_), .B(new_n1335_), .Y(new_n6412_));
  NAND2 g06027(.A(new_n1337_), .B(\req[58] ), .Y(new_n6413_));
  NOR2  g06028(.A(new_n6413_), .B(new_n6412_), .Y(\grant[58] ));
  INV   g06029(.A(new_n1346_), .Y(new_n6415_));
  NOR2  g06030(.A(new_n6415_), .B(new_n585_), .Y(new_n6416_));
  NOR2  g06031(.A(new_n6416_), .B(new_n1351_), .Y(new_n6417_));
  NOR2  g06032(.A(new_n6417_), .B(new_n1355_), .Y(new_n6418_));
  NOR2  g06033(.A(new_n6418_), .B(new_n1359_), .Y(new_n6419_));
  NOR2  g06034(.A(new_n6419_), .B(new_n1363_), .Y(new_n6420_));
  NOR2  g06035(.A(new_n6420_), .B(new_n1367_), .Y(new_n6421_));
  NOR2  g06036(.A(new_n6421_), .B(new_n1371_), .Y(new_n6422_));
  NOR2  g06037(.A(new_n6422_), .B(new_n1375_), .Y(new_n6423_));
  NOR2  g06038(.A(new_n6423_), .B(new_n1379_), .Y(new_n6424_));
  NOR2  g06039(.A(new_n6424_), .B(new_n1383_), .Y(new_n6425_));
  NOR2  g06040(.A(new_n6425_), .B(new_n1387_), .Y(new_n6426_));
  NOR2  g06041(.A(new_n6426_), .B(new_n1391_), .Y(new_n6427_));
  NOR2  g06042(.A(new_n6427_), .B(new_n1395_), .Y(new_n6428_));
  NOR2  g06043(.A(new_n6428_), .B(new_n1399_), .Y(new_n6429_));
  NOR2  g06044(.A(new_n6429_), .B(new_n1403_), .Y(new_n6430_));
  NOR2  g06045(.A(new_n6430_), .B(new_n1407_), .Y(new_n6431_));
  NOR2  g06046(.A(new_n6431_), .B(new_n1411_), .Y(new_n6432_));
  NOR2  g06047(.A(new_n6432_), .B(new_n1415_), .Y(new_n6433_));
  NOR2  g06048(.A(new_n6433_), .B(new_n1419_), .Y(new_n6434_));
  NOR2  g06049(.A(new_n6434_), .B(new_n1423_), .Y(new_n6435_));
  NOR2  g06050(.A(new_n6435_), .B(new_n1427_), .Y(new_n6436_));
  NOR2  g06051(.A(new_n6436_), .B(new_n1431_), .Y(new_n6437_));
  NOR2  g06052(.A(new_n6437_), .B(new_n1435_), .Y(new_n6438_));
  NOR2  g06053(.A(new_n6438_), .B(new_n1439_), .Y(new_n6439_));
  NOR2  g06054(.A(new_n6439_), .B(new_n1443_), .Y(new_n6440_));
  NOR2  g06055(.A(new_n6440_), .B(new_n1447_), .Y(new_n6441_));
  NOR2  g06056(.A(new_n6441_), .B(new_n1451_), .Y(new_n6442_));
  NOR2  g06057(.A(new_n6442_), .B(new_n1455_), .Y(new_n6443_));
  NOR2  g06058(.A(new_n6443_), .B(new_n1459_), .Y(new_n6444_));
  NOR2  g06059(.A(new_n6444_), .B(new_n1463_), .Y(new_n6445_));
  NOR2  g06060(.A(new_n6445_), .B(new_n1467_), .Y(new_n6446_));
  NOR2  g06061(.A(new_n6446_), .B(new_n1471_), .Y(new_n6447_));
  NOR2  g06062(.A(new_n6447_), .B(new_n1475_), .Y(new_n6448_));
  NOR2  g06063(.A(new_n6448_), .B(new_n1479_), .Y(new_n6449_));
  NOR2  g06064(.A(new_n6449_), .B(new_n1483_), .Y(new_n6450_));
  NOR2  g06065(.A(new_n6450_), .B(new_n1487_), .Y(new_n6451_));
  NOR2  g06066(.A(new_n6451_), .B(new_n1491_), .Y(new_n6452_));
  NOR2  g06067(.A(new_n6452_), .B(new_n1495_), .Y(new_n6453_));
  NOR2  g06068(.A(new_n6453_), .B(new_n1499_), .Y(new_n6454_));
  NOR2  g06069(.A(new_n6454_), .B(new_n1503_), .Y(new_n6455_));
  NOR2  g06070(.A(new_n6455_), .B(new_n1507_), .Y(new_n6456_));
  NOR2  g06071(.A(new_n6456_), .B(new_n1511_), .Y(new_n6457_));
  NOR2  g06072(.A(new_n6457_), .B(new_n1515_), .Y(new_n6458_));
  NOR2  g06073(.A(new_n6458_), .B(new_n1519_), .Y(new_n6459_));
  NOR2  g06074(.A(new_n6459_), .B(new_n1523_), .Y(new_n6460_));
  NOR2  g06075(.A(new_n6460_), .B(new_n1527_), .Y(new_n6461_));
  NOR2  g06076(.A(new_n6461_), .B(new_n1797_), .Y(new_n6462_));
  NOR2  g06077(.A(new_n6462_), .B(new_n396_), .Y(new_n6463_));
  NOR2  g06078(.A(new_n6463_), .B(new_n400_), .Y(new_n6464_));
  NOR2  g06079(.A(new_n6464_), .B(new_n406_), .Y(new_n6465_));
  NOR2  g06080(.A(new_n6465_), .B(new_n410_), .Y(new_n6466_));
  NOR2  g06081(.A(new_n6466_), .B(new_n416_), .Y(new_n6467_));
  NOR2  g06082(.A(new_n6467_), .B(new_n420_), .Y(new_n6468_));
  NOR2  g06083(.A(new_n6468_), .B(new_n426_), .Y(new_n6469_));
  NOR2  g06084(.A(new_n6469_), .B(new_n430_), .Y(new_n6470_));
  NOR2  g06085(.A(new_n6470_), .B(new_n436_), .Y(new_n6471_));
  NOR2  g06086(.A(new_n6471_), .B(new_n440_), .Y(new_n6472_));
  NOR2  g06087(.A(new_n6472_), .B(new_n446_), .Y(new_n6473_));
  NOR2  g06088(.A(new_n6473_), .B(new_n450_), .Y(new_n6474_));
  NOR2  g06089(.A(new_n6474_), .B(new_n456_), .Y(new_n6475_));
  NOR2  g06090(.A(new_n6475_), .B(new_n460_), .Y(new_n6476_));
  NOR2  g06091(.A(new_n6476_), .B(new_n466_), .Y(new_n6477_));
  NOR2  g06092(.A(new_n6477_), .B(new_n470_), .Y(new_n6478_));
  NOR2  g06093(.A(new_n6478_), .B(new_n476_), .Y(new_n6479_));
  NOR2  g06094(.A(new_n6479_), .B(new_n480_), .Y(new_n6480_));
  NOR2  g06095(.A(new_n6480_), .B(new_n486_), .Y(new_n6481_));
  NOR2  g06096(.A(new_n6481_), .B(new_n490_), .Y(new_n6482_));
  NOR2  g06097(.A(new_n6482_), .B(new_n496_), .Y(new_n6483_));
  NOR2  g06098(.A(new_n6483_), .B(new_n500_), .Y(new_n6484_));
  NOR2  g06099(.A(new_n6484_), .B(new_n506_), .Y(new_n6485_));
  NOR2  g06100(.A(new_n6485_), .B(new_n510_), .Y(new_n6486_));
  NOR2  g06101(.A(new_n6486_), .B(new_n516_), .Y(new_n6487_));
  NOR2  g06102(.A(new_n6487_), .B(new_n520_), .Y(new_n6488_));
  NOR2  g06103(.A(new_n6488_), .B(new_n526_), .Y(new_n6489_));
  NOR2  g06104(.A(new_n6489_), .B(new_n530_), .Y(new_n6490_));
  NOR2  g06105(.A(new_n6490_), .B(new_n536_), .Y(new_n6491_));
  NOR2  g06106(.A(new_n6491_), .B(new_n540_), .Y(new_n6492_));
  NOR2  g06107(.A(new_n6492_), .B(new_n546_), .Y(new_n6493_));
  NOR2  g06108(.A(new_n6493_), .B(new_n550_), .Y(new_n6494_));
  NOR2  g06109(.A(new_n6494_), .B(new_n556_), .Y(new_n6495_));
  NOR2  g06110(.A(new_n6495_), .B(new_n560_), .Y(new_n6496_));
  NOR2  g06111(.A(new_n6496_), .B(new_n566_), .Y(new_n6497_));
  NOR2  g06112(.A(new_n6497_), .B(new_n570_), .Y(new_n6498_));
  NOR2  g06113(.A(new_n6498_), .B(new_n576_), .Y(new_n6499_));
  NAND2 g06114(.A(new_n578_), .B(\req[59] ), .Y(new_n6500_));
  NOR2  g06115(.A(new_n6500_), .B(new_n6499_), .Y(\grant[59] ));
  INV   g06116(.A(new_n589_), .Y(new_n6502_));
  NOR2  g06117(.A(new_n990_), .B(new_n6502_), .Y(new_n6503_));
  NOR2  g06118(.A(new_n6503_), .B(new_n596_), .Y(new_n6504_));
  NOR2  g06119(.A(new_n6504_), .B(new_n600_), .Y(new_n6505_));
  NOR2  g06120(.A(new_n6505_), .B(new_n606_), .Y(new_n6506_));
  NOR2  g06121(.A(new_n6506_), .B(new_n610_), .Y(new_n6507_));
  NOR2  g06122(.A(new_n6507_), .B(new_n616_), .Y(new_n6508_));
  NOR2  g06123(.A(new_n6508_), .B(new_n620_), .Y(new_n6509_));
  NOR2  g06124(.A(new_n6509_), .B(new_n626_), .Y(new_n6510_));
  NOR2  g06125(.A(new_n6510_), .B(new_n630_), .Y(new_n6511_));
  NOR2  g06126(.A(new_n6511_), .B(new_n636_), .Y(new_n6512_));
  NOR2  g06127(.A(new_n6512_), .B(new_n640_), .Y(new_n6513_));
  NOR2  g06128(.A(new_n6513_), .B(new_n646_), .Y(new_n6514_));
  NOR2  g06129(.A(new_n6514_), .B(new_n650_), .Y(new_n6515_));
  NOR2  g06130(.A(new_n6515_), .B(new_n656_), .Y(new_n6516_));
  NOR2  g06131(.A(new_n6516_), .B(new_n660_), .Y(new_n6517_));
  NOR2  g06132(.A(new_n6517_), .B(new_n666_), .Y(new_n6518_));
  NOR2  g06133(.A(new_n6518_), .B(new_n670_), .Y(new_n6519_));
  NOR2  g06134(.A(new_n6519_), .B(new_n676_), .Y(new_n6520_));
  NOR2  g06135(.A(new_n6520_), .B(new_n680_), .Y(new_n6521_));
  NOR2  g06136(.A(new_n6521_), .B(new_n686_), .Y(new_n6522_));
  NOR2  g06137(.A(new_n6522_), .B(new_n690_), .Y(new_n6523_));
  NOR2  g06138(.A(new_n6523_), .B(new_n696_), .Y(new_n6524_));
  NOR2  g06139(.A(new_n6524_), .B(new_n700_), .Y(new_n6525_));
  NOR2  g06140(.A(new_n6525_), .B(new_n706_), .Y(new_n6526_));
  NOR2  g06141(.A(new_n6526_), .B(new_n710_), .Y(new_n6527_));
  NOR2  g06142(.A(new_n6527_), .B(new_n716_), .Y(new_n6528_));
  NOR2  g06143(.A(new_n6528_), .B(new_n720_), .Y(new_n6529_));
  NOR2  g06144(.A(new_n6529_), .B(new_n726_), .Y(new_n6530_));
  NOR2  g06145(.A(new_n6530_), .B(new_n730_), .Y(new_n6531_));
  NOR2  g06146(.A(new_n6531_), .B(new_n736_), .Y(new_n6532_));
  NOR2  g06147(.A(new_n6532_), .B(new_n740_), .Y(new_n6533_));
  NOR2  g06148(.A(new_n6533_), .B(new_n746_), .Y(new_n6534_));
  NOR2  g06149(.A(new_n6534_), .B(new_n750_), .Y(new_n6535_));
  NOR2  g06150(.A(new_n6535_), .B(new_n756_), .Y(new_n6536_));
  NOR2  g06151(.A(new_n6536_), .B(new_n760_), .Y(new_n6537_));
  NOR2  g06152(.A(new_n6537_), .B(new_n766_), .Y(new_n6538_));
  NOR2  g06153(.A(new_n6538_), .B(new_n770_), .Y(new_n6539_));
  NOR2  g06154(.A(new_n6539_), .B(new_n776_), .Y(new_n6540_));
  NOR2  g06155(.A(new_n6540_), .B(new_n780_), .Y(new_n6541_));
  NOR2  g06156(.A(new_n6541_), .B(new_n786_), .Y(new_n6542_));
  NOR2  g06157(.A(new_n6542_), .B(new_n790_), .Y(new_n6543_));
  NOR2  g06158(.A(new_n6543_), .B(new_n796_), .Y(new_n6544_));
  NOR2  g06159(.A(new_n6544_), .B(new_n800_), .Y(new_n6545_));
  NOR2  g06160(.A(new_n6545_), .B(new_n806_), .Y(new_n6546_));
  NOR2  g06161(.A(new_n6546_), .B(new_n1616_), .Y(new_n6547_));
  NOR2  g06162(.A(new_n6547_), .B(new_n1618_), .Y(new_n6548_));
  NOR2  g06163(.A(new_n6548_), .B(new_n1885_), .Y(new_n6549_));
  NOR2  g06164(.A(new_n6549_), .B(new_n820_), .Y(new_n6550_));
  NOR2  g06165(.A(new_n6550_), .B(new_n824_), .Y(new_n6551_));
  NOR2  g06166(.A(new_n6551_), .B(new_n829_), .Y(new_n6552_));
  NOR2  g06167(.A(new_n6552_), .B(new_n833_), .Y(new_n6553_));
  NOR2  g06168(.A(new_n6553_), .B(new_n838_), .Y(new_n6554_));
  NOR2  g06169(.A(new_n6554_), .B(new_n842_), .Y(new_n6555_));
  NOR2  g06170(.A(new_n6555_), .B(new_n847_), .Y(new_n6556_));
  NOR2  g06171(.A(new_n6556_), .B(new_n851_), .Y(new_n6557_));
  NOR2  g06172(.A(new_n6557_), .B(new_n856_), .Y(new_n6558_));
  NOR2  g06173(.A(new_n6558_), .B(new_n860_), .Y(new_n6559_));
  NOR2  g06174(.A(new_n6559_), .B(new_n865_), .Y(new_n6560_));
  NOR2  g06175(.A(new_n6560_), .B(new_n869_), .Y(new_n6561_));
  NOR2  g06176(.A(new_n6561_), .B(new_n874_), .Y(new_n6562_));
  NOR2  g06177(.A(new_n6562_), .B(new_n878_), .Y(new_n6563_));
  NOR2  g06178(.A(new_n6563_), .B(new_n883_), .Y(new_n6564_));
  NOR2  g06179(.A(new_n6564_), .B(new_n887_), .Y(new_n6565_));
  NOR2  g06180(.A(new_n6565_), .B(new_n892_), .Y(new_n6566_));
  NOR2  g06181(.A(new_n6566_), .B(new_n896_), .Y(new_n6567_));
  NOR2  g06182(.A(new_n6567_), .B(new_n901_), .Y(new_n6568_));
  NOR2  g06183(.A(new_n6568_), .B(new_n905_), .Y(new_n6569_));
  NOR2  g06184(.A(new_n6569_), .B(new_n910_), .Y(new_n6570_));
  NOR2  g06185(.A(new_n6570_), .B(new_n914_), .Y(new_n6571_));
  NOR2  g06186(.A(new_n6571_), .B(new_n919_), .Y(new_n6572_));
  NOR2  g06187(.A(new_n6572_), .B(new_n923_), .Y(new_n6573_));
  NOR2  g06188(.A(new_n6573_), .B(new_n928_), .Y(new_n6574_));
  NOR2  g06189(.A(new_n6574_), .B(new_n932_), .Y(new_n6575_));
  NOR2  g06190(.A(new_n6575_), .B(new_n937_), .Y(new_n6576_));
  NOR2  g06191(.A(new_n6576_), .B(new_n941_), .Y(new_n6577_));
  NOR2  g06192(.A(new_n6577_), .B(new_n946_), .Y(new_n6578_));
  NOR2  g06193(.A(new_n6578_), .B(new_n950_), .Y(new_n6579_));
  NOR2  g06194(.A(new_n6579_), .B(new_n955_), .Y(new_n6580_));
  NOR2  g06195(.A(new_n6580_), .B(new_n959_), .Y(new_n6581_));
  NOR2  g06196(.A(new_n6581_), .B(new_n964_), .Y(new_n6582_));
  NOR2  g06197(.A(new_n6582_), .B(new_n968_), .Y(new_n6583_));
  NOR2  g06198(.A(new_n6583_), .B(new_n973_), .Y(new_n6584_));
  NOR2  g06199(.A(new_n6584_), .B(new_n977_), .Y(new_n6585_));
  NOR2  g06200(.A(new_n6585_), .B(new_n982_), .Y(new_n6586_));
  NAND2 g06201(.A(new_n984_), .B(\req[60] ), .Y(new_n6587_));
  NOR2  g06202(.A(new_n6587_), .B(new_n6586_), .Y(\grant[60] ));
  INV   g06203(.A(new_n994_), .Y(new_n6589_));
  NOR2  g06204(.A(new_n1350_), .B(new_n6589_), .Y(new_n6590_));
  NOR2  g06205(.A(new_n6590_), .B(new_n1000_), .Y(new_n6591_));
  NOR2  g06206(.A(new_n6591_), .B(new_n1004_), .Y(new_n6592_));
  NOR2  g06207(.A(new_n6592_), .B(new_n1009_), .Y(new_n6593_));
  NOR2  g06208(.A(new_n6593_), .B(new_n1013_), .Y(new_n6594_));
  NOR2  g06209(.A(new_n6594_), .B(new_n1018_), .Y(new_n6595_));
  NOR2  g06210(.A(new_n6595_), .B(new_n1022_), .Y(new_n6596_));
  NOR2  g06211(.A(new_n6596_), .B(new_n1027_), .Y(new_n6597_));
  NOR2  g06212(.A(new_n6597_), .B(new_n1031_), .Y(new_n6598_));
  NOR2  g06213(.A(new_n6598_), .B(new_n1036_), .Y(new_n6599_));
  NOR2  g06214(.A(new_n6599_), .B(new_n1040_), .Y(new_n6600_));
  NOR2  g06215(.A(new_n6600_), .B(new_n1045_), .Y(new_n6601_));
  NOR2  g06216(.A(new_n6601_), .B(new_n1049_), .Y(new_n6602_));
  NOR2  g06217(.A(new_n6602_), .B(new_n1054_), .Y(new_n6603_));
  NOR2  g06218(.A(new_n6603_), .B(new_n1058_), .Y(new_n6604_));
  NOR2  g06219(.A(new_n6604_), .B(new_n1063_), .Y(new_n6605_));
  NOR2  g06220(.A(new_n6605_), .B(new_n1067_), .Y(new_n6606_));
  NOR2  g06221(.A(new_n6606_), .B(new_n1072_), .Y(new_n6607_));
  NOR2  g06222(.A(new_n6607_), .B(new_n1076_), .Y(new_n6608_));
  NOR2  g06223(.A(new_n6608_), .B(new_n1081_), .Y(new_n6609_));
  NOR2  g06224(.A(new_n6609_), .B(new_n1085_), .Y(new_n6610_));
  NOR2  g06225(.A(new_n6610_), .B(new_n1090_), .Y(new_n6611_));
  NOR2  g06226(.A(new_n6611_), .B(new_n1094_), .Y(new_n6612_));
  NOR2  g06227(.A(new_n6612_), .B(new_n1099_), .Y(new_n6613_));
  NOR2  g06228(.A(new_n6613_), .B(new_n1103_), .Y(new_n6614_));
  NOR2  g06229(.A(new_n6614_), .B(new_n1108_), .Y(new_n6615_));
  NOR2  g06230(.A(new_n6615_), .B(new_n1112_), .Y(new_n6616_));
  NOR2  g06231(.A(new_n6616_), .B(new_n1117_), .Y(new_n6617_));
  NOR2  g06232(.A(new_n6617_), .B(new_n1121_), .Y(new_n6618_));
  NOR2  g06233(.A(new_n6618_), .B(new_n1126_), .Y(new_n6619_));
  NOR2  g06234(.A(new_n6619_), .B(new_n1130_), .Y(new_n6620_));
  NOR2  g06235(.A(new_n6620_), .B(new_n1135_), .Y(new_n6621_));
  NOR2  g06236(.A(new_n6621_), .B(new_n1139_), .Y(new_n6622_));
  NOR2  g06237(.A(new_n6622_), .B(new_n1144_), .Y(new_n6623_));
  NOR2  g06238(.A(new_n6623_), .B(new_n1148_), .Y(new_n6624_));
  NOR2  g06239(.A(new_n6624_), .B(new_n1153_), .Y(new_n6625_));
  NOR2  g06240(.A(new_n6625_), .B(new_n1157_), .Y(new_n6626_));
  NOR2  g06241(.A(new_n6626_), .B(new_n1162_), .Y(new_n6627_));
  NOR2  g06242(.A(new_n6627_), .B(new_n1166_), .Y(new_n6628_));
  NOR2  g06243(.A(new_n6628_), .B(new_n1171_), .Y(new_n6629_));
  NOR2  g06244(.A(new_n6629_), .B(new_n1175_), .Y(new_n6630_));
  NOR2  g06245(.A(new_n6630_), .B(new_n1180_), .Y(new_n6631_));
  NOR2  g06246(.A(new_n6631_), .B(new_n1184_), .Y(new_n6632_));
  NOR2  g06247(.A(new_n6632_), .B(new_n1189_), .Y(new_n6633_));
  NOR2  g06248(.A(new_n6633_), .B(new_n1707_), .Y(new_n6634_));
  NOR2  g06249(.A(new_n6634_), .B(new_n1709_), .Y(new_n6635_));
  NOR2  g06250(.A(new_n6635_), .B(new_n1973_), .Y(new_n6636_));
  NOR2  g06251(.A(new_n6636_), .B(new_n1199_), .Y(new_n6637_));
  NOR2  g06252(.A(new_n6637_), .B(new_n1203_), .Y(new_n6638_));
  NOR2  g06253(.A(new_n6638_), .B(new_n1207_), .Y(new_n6639_));
  NOR2  g06254(.A(new_n6639_), .B(new_n1211_), .Y(new_n6640_));
  NOR2  g06255(.A(new_n6640_), .B(new_n1215_), .Y(new_n6641_));
  NOR2  g06256(.A(new_n6641_), .B(new_n1219_), .Y(new_n6642_));
  NOR2  g06257(.A(new_n6642_), .B(new_n1223_), .Y(new_n6643_));
  NOR2  g06258(.A(new_n6643_), .B(new_n1227_), .Y(new_n6644_));
  NOR2  g06259(.A(new_n6644_), .B(new_n1231_), .Y(new_n6645_));
  NOR2  g06260(.A(new_n6645_), .B(new_n1235_), .Y(new_n6646_));
  NOR2  g06261(.A(new_n6646_), .B(new_n1239_), .Y(new_n6647_));
  NOR2  g06262(.A(new_n6647_), .B(new_n1243_), .Y(new_n6648_));
  NOR2  g06263(.A(new_n6648_), .B(new_n1247_), .Y(new_n6649_));
  NOR2  g06264(.A(new_n6649_), .B(new_n1251_), .Y(new_n6650_));
  NOR2  g06265(.A(new_n6650_), .B(new_n1255_), .Y(new_n6651_));
  NOR2  g06266(.A(new_n6651_), .B(new_n1259_), .Y(new_n6652_));
  NOR2  g06267(.A(new_n6652_), .B(new_n1263_), .Y(new_n6653_));
  NOR2  g06268(.A(new_n6653_), .B(new_n1267_), .Y(new_n6654_));
  NOR2  g06269(.A(new_n6654_), .B(new_n1271_), .Y(new_n6655_));
  NOR2  g06270(.A(new_n6655_), .B(new_n1275_), .Y(new_n6656_));
  NOR2  g06271(.A(new_n6656_), .B(new_n1279_), .Y(new_n6657_));
  NOR2  g06272(.A(new_n6657_), .B(new_n1283_), .Y(new_n6658_));
  NOR2  g06273(.A(new_n6658_), .B(new_n1287_), .Y(new_n6659_));
  NOR2  g06274(.A(new_n6659_), .B(new_n1291_), .Y(new_n6660_));
  NOR2  g06275(.A(new_n6660_), .B(new_n1295_), .Y(new_n6661_));
  NOR2  g06276(.A(new_n6661_), .B(new_n1299_), .Y(new_n6662_));
  NOR2  g06277(.A(new_n6662_), .B(new_n1303_), .Y(new_n6663_));
  NOR2  g06278(.A(new_n6663_), .B(new_n1307_), .Y(new_n6664_));
  NOR2  g06279(.A(new_n6664_), .B(new_n1311_), .Y(new_n6665_));
  NOR2  g06280(.A(new_n6665_), .B(new_n1315_), .Y(new_n6666_));
  NOR2  g06281(.A(new_n6666_), .B(new_n1319_), .Y(new_n6667_));
  NOR2  g06282(.A(new_n6667_), .B(new_n1323_), .Y(new_n6668_));
  NOR2  g06283(.A(new_n6668_), .B(new_n1327_), .Y(new_n6669_));
  NOR2  g06284(.A(new_n6669_), .B(new_n1331_), .Y(new_n6670_));
  NOR2  g06285(.A(new_n6670_), .B(new_n1335_), .Y(new_n6671_));
  NOR2  g06286(.A(new_n6671_), .B(new_n1339_), .Y(new_n6672_));
  NOR2  g06287(.A(new_n6672_), .B(new_n1343_), .Y(new_n6673_));
  NAND2 g06288(.A(new_n1345_), .B(\req[61] ), .Y(new_n6674_));
  NOR2  g06289(.A(new_n6674_), .B(new_n6673_), .Y(\grant[61] ));
  INV   g06290(.A(new_n1354_), .Y(new_n6676_));
  NOR2  g06291(.A(new_n6676_), .B(new_n595_), .Y(new_n6677_));
  NOR2  g06292(.A(new_n6677_), .B(new_n1359_), .Y(new_n6678_));
  NOR2  g06293(.A(new_n6678_), .B(new_n1363_), .Y(new_n6679_));
  NOR2  g06294(.A(new_n6679_), .B(new_n1367_), .Y(new_n6680_));
  NOR2  g06295(.A(new_n6680_), .B(new_n1371_), .Y(new_n6681_));
  NOR2  g06296(.A(new_n6681_), .B(new_n1375_), .Y(new_n6682_));
  NOR2  g06297(.A(new_n6682_), .B(new_n1379_), .Y(new_n6683_));
  NOR2  g06298(.A(new_n6683_), .B(new_n1383_), .Y(new_n6684_));
  NOR2  g06299(.A(new_n6684_), .B(new_n1387_), .Y(new_n6685_));
  NOR2  g06300(.A(new_n6685_), .B(new_n1391_), .Y(new_n6686_));
  NOR2  g06301(.A(new_n6686_), .B(new_n1395_), .Y(new_n6687_));
  NOR2  g06302(.A(new_n6687_), .B(new_n1399_), .Y(new_n6688_));
  NOR2  g06303(.A(new_n6688_), .B(new_n1403_), .Y(new_n6689_));
  NOR2  g06304(.A(new_n6689_), .B(new_n1407_), .Y(new_n6690_));
  NOR2  g06305(.A(new_n6690_), .B(new_n1411_), .Y(new_n6691_));
  NOR2  g06306(.A(new_n6691_), .B(new_n1415_), .Y(new_n6692_));
  NOR2  g06307(.A(new_n6692_), .B(new_n1419_), .Y(new_n6693_));
  NOR2  g06308(.A(new_n6693_), .B(new_n1423_), .Y(new_n6694_));
  NOR2  g06309(.A(new_n6694_), .B(new_n1427_), .Y(new_n6695_));
  NOR2  g06310(.A(new_n6695_), .B(new_n1431_), .Y(new_n6696_));
  NOR2  g06311(.A(new_n6696_), .B(new_n1435_), .Y(new_n6697_));
  NOR2  g06312(.A(new_n6697_), .B(new_n1439_), .Y(new_n6698_));
  NOR2  g06313(.A(new_n6698_), .B(new_n1443_), .Y(new_n6699_));
  NOR2  g06314(.A(new_n6699_), .B(new_n1447_), .Y(new_n6700_));
  NOR2  g06315(.A(new_n6700_), .B(new_n1451_), .Y(new_n6701_));
  NOR2  g06316(.A(new_n6701_), .B(new_n1455_), .Y(new_n6702_));
  NOR2  g06317(.A(new_n6702_), .B(new_n1459_), .Y(new_n6703_));
  NOR2  g06318(.A(new_n6703_), .B(new_n1463_), .Y(new_n6704_));
  NOR2  g06319(.A(new_n6704_), .B(new_n1467_), .Y(new_n6705_));
  NOR2  g06320(.A(new_n6705_), .B(new_n1471_), .Y(new_n6706_));
  NOR2  g06321(.A(new_n6706_), .B(new_n1475_), .Y(new_n6707_));
  NOR2  g06322(.A(new_n6707_), .B(new_n1479_), .Y(new_n6708_));
  NOR2  g06323(.A(new_n6708_), .B(new_n1483_), .Y(new_n6709_));
  NOR2  g06324(.A(new_n6709_), .B(new_n1487_), .Y(new_n6710_));
  NOR2  g06325(.A(new_n6710_), .B(new_n1491_), .Y(new_n6711_));
  NOR2  g06326(.A(new_n6711_), .B(new_n1495_), .Y(new_n6712_));
  NOR2  g06327(.A(new_n6712_), .B(new_n1499_), .Y(new_n6713_));
  NOR2  g06328(.A(new_n6713_), .B(new_n1503_), .Y(new_n6714_));
  NOR2  g06329(.A(new_n6714_), .B(new_n1507_), .Y(new_n6715_));
  NOR2  g06330(.A(new_n6715_), .B(new_n1511_), .Y(new_n6716_));
  NOR2  g06331(.A(new_n6716_), .B(new_n1515_), .Y(new_n6717_));
  NOR2  g06332(.A(new_n6717_), .B(new_n1519_), .Y(new_n6718_));
  NOR2  g06333(.A(new_n6718_), .B(new_n1523_), .Y(new_n6719_));
  NOR2  g06334(.A(new_n6719_), .B(new_n1527_), .Y(new_n6720_));
  NOR2  g06335(.A(new_n6720_), .B(new_n1797_), .Y(new_n6721_));
  NOR2  g06336(.A(new_n6721_), .B(new_n396_), .Y(new_n6722_));
  NOR2  g06337(.A(new_n6722_), .B(new_n400_), .Y(new_n6723_));
  NOR2  g06338(.A(new_n6723_), .B(new_n406_), .Y(new_n6724_));
  NOR2  g06339(.A(new_n6724_), .B(new_n410_), .Y(new_n6725_));
  NOR2  g06340(.A(new_n6725_), .B(new_n416_), .Y(new_n6726_));
  NOR2  g06341(.A(new_n6726_), .B(new_n420_), .Y(new_n6727_));
  NOR2  g06342(.A(new_n6727_), .B(new_n426_), .Y(new_n6728_));
  NOR2  g06343(.A(new_n6728_), .B(new_n430_), .Y(new_n6729_));
  NOR2  g06344(.A(new_n6729_), .B(new_n436_), .Y(new_n6730_));
  NOR2  g06345(.A(new_n6730_), .B(new_n440_), .Y(new_n6731_));
  NOR2  g06346(.A(new_n6731_), .B(new_n446_), .Y(new_n6732_));
  NOR2  g06347(.A(new_n6732_), .B(new_n450_), .Y(new_n6733_));
  NOR2  g06348(.A(new_n6733_), .B(new_n456_), .Y(new_n6734_));
  NOR2  g06349(.A(new_n6734_), .B(new_n460_), .Y(new_n6735_));
  NOR2  g06350(.A(new_n6735_), .B(new_n466_), .Y(new_n6736_));
  NOR2  g06351(.A(new_n6736_), .B(new_n470_), .Y(new_n6737_));
  NOR2  g06352(.A(new_n6737_), .B(new_n476_), .Y(new_n6738_));
  NOR2  g06353(.A(new_n6738_), .B(new_n480_), .Y(new_n6739_));
  NOR2  g06354(.A(new_n6739_), .B(new_n486_), .Y(new_n6740_));
  NOR2  g06355(.A(new_n6740_), .B(new_n490_), .Y(new_n6741_));
  NOR2  g06356(.A(new_n6741_), .B(new_n496_), .Y(new_n6742_));
  NOR2  g06357(.A(new_n6742_), .B(new_n500_), .Y(new_n6743_));
  NOR2  g06358(.A(new_n6743_), .B(new_n506_), .Y(new_n6744_));
  NOR2  g06359(.A(new_n6744_), .B(new_n510_), .Y(new_n6745_));
  NOR2  g06360(.A(new_n6745_), .B(new_n516_), .Y(new_n6746_));
  NOR2  g06361(.A(new_n6746_), .B(new_n520_), .Y(new_n6747_));
  NOR2  g06362(.A(new_n6747_), .B(new_n526_), .Y(new_n6748_));
  NOR2  g06363(.A(new_n6748_), .B(new_n530_), .Y(new_n6749_));
  NOR2  g06364(.A(new_n6749_), .B(new_n536_), .Y(new_n6750_));
  NOR2  g06365(.A(new_n6750_), .B(new_n540_), .Y(new_n6751_));
  NOR2  g06366(.A(new_n6751_), .B(new_n546_), .Y(new_n6752_));
  NOR2  g06367(.A(new_n6752_), .B(new_n550_), .Y(new_n6753_));
  NOR2  g06368(.A(new_n6753_), .B(new_n556_), .Y(new_n6754_));
  NOR2  g06369(.A(new_n6754_), .B(new_n560_), .Y(new_n6755_));
  NOR2  g06370(.A(new_n6755_), .B(new_n566_), .Y(new_n6756_));
  NOR2  g06371(.A(new_n6756_), .B(new_n570_), .Y(new_n6757_));
  NOR2  g06372(.A(new_n6757_), .B(new_n576_), .Y(new_n6758_));
  NOR2  g06373(.A(new_n6758_), .B(new_n580_), .Y(new_n6759_));
  NOR2  g06374(.A(new_n6759_), .B(new_n586_), .Y(new_n6760_));
  NAND2 g06375(.A(new_n588_), .B(\req[62] ), .Y(new_n6761_));
  NOR2  g06376(.A(new_n6761_), .B(new_n6760_), .Y(\grant[62] ));
  INV   g06377(.A(new_n599_), .Y(new_n6763_));
  NOR2  g06378(.A(new_n999_), .B(new_n6763_), .Y(new_n6764_));
  NOR2  g06379(.A(new_n6764_), .B(new_n606_), .Y(new_n6765_));
  NOR2  g06380(.A(new_n6765_), .B(new_n610_), .Y(new_n6766_));
  NOR2  g06381(.A(new_n6766_), .B(new_n616_), .Y(new_n6767_));
  NOR2  g06382(.A(new_n6767_), .B(new_n620_), .Y(new_n6768_));
  NOR2  g06383(.A(new_n6768_), .B(new_n626_), .Y(new_n6769_));
  NOR2  g06384(.A(new_n6769_), .B(new_n630_), .Y(new_n6770_));
  NOR2  g06385(.A(new_n6770_), .B(new_n636_), .Y(new_n6771_));
  NOR2  g06386(.A(new_n6771_), .B(new_n640_), .Y(new_n6772_));
  NOR2  g06387(.A(new_n6772_), .B(new_n646_), .Y(new_n6773_));
  NOR2  g06388(.A(new_n6773_), .B(new_n650_), .Y(new_n6774_));
  NOR2  g06389(.A(new_n6774_), .B(new_n656_), .Y(new_n6775_));
  NOR2  g06390(.A(new_n6775_), .B(new_n660_), .Y(new_n6776_));
  NOR2  g06391(.A(new_n6776_), .B(new_n666_), .Y(new_n6777_));
  NOR2  g06392(.A(new_n6777_), .B(new_n670_), .Y(new_n6778_));
  NOR2  g06393(.A(new_n6778_), .B(new_n676_), .Y(new_n6779_));
  NOR2  g06394(.A(new_n6779_), .B(new_n680_), .Y(new_n6780_));
  NOR2  g06395(.A(new_n6780_), .B(new_n686_), .Y(new_n6781_));
  NOR2  g06396(.A(new_n6781_), .B(new_n690_), .Y(new_n6782_));
  NOR2  g06397(.A(new_n6782_), .B(new_n696_), .Y(new_n6783_));
  NOR2  g06398(.A(new_n6783_), .B(new_n700_), .Y(new_n6784_));
  NOR2  g06399(.A(new_n6784_), .B(new_n706_), .Y(new_n6785_));
  NOR2  g06400(.A(new_n6785_), .B(new_n710_), .Y(new_n6786_));
  NOR2  g06401(.A(new_n6786_), .B(new_n716_), .Y(new_n6787_));
  NOR2  g06402(.A(new_n6787_), .B(new_n720_), .Y(new_n6788_));
  NOR2  g06403(.A(new_n6788_), .B(new_n726_), .Y(new_n6789_));
  NOR2  g06404(.A(new_n6789_), .B(new_n730_), .Y(new_n6790_));
  NOR2  g06405(.A(new_n6790_), .B(new_n736_), .Y(new_n6791_));
  NOR2  g06406(.A(new_n6791_), .B(new_n740_), .Y(new_n6792_));
  NOR2  g06407(.A(new_n6792_), .B(new_n746_), .Y(new_n6793_));
  NOR2  g06408(.A(new_n6793_), .B(new_n750_), .Y(new_n6794_));
  NOR2  g06409(.A(new_n6794_), .B(new_n756_), .Y(new_n6795_));
  NOR2  g06410(.A(new_n6795_), .B(new_n760_), .Y(new_n6796_));
  NOR2  g06411(.A(new_n6796_), .B(new_n766_), .Y(new_n6797_));
  NOR2  g06412(.A(new_n6797_), .B(new_n770_), .Y(new_n6798_));
  NOR2  g06413(.A(new_n6798_), .B(new_n776_), .Y(new_n6799_));
  NOR2  g06414(.A(new_n6799_), .B(new_n780_), .Y(new_n6800_));
  NOR2  g06415(.A(new_n6800_), .B(new_n786_), .Y(new_n6801_));
  NOR2  g06416(.A(new_n6801_), .B(new_n790_), .Y(new_n6802_));
  NOR2  g06417(.A(new_n6802_), .B(new_n796_), .Y(new_n6803_));
  NOR2  g06418(.A(new_n6803_), .B(new_n800_), .Y(new_n6804_));
  NOR2  g06419(.A(new_n6804_), .B(new_n806_), .Y(new_n6805_));
  NOR2  g06420(.A(new_n6805_), .B(new_n1616_), .Y(new_n6806_));
  NOR2  g06421(.A(new_n6806_), .B(new_n1618_), .Y(new_n6807_));
  NOR2  g06422(.A(new_n6807_), .B(new_n1885_), .Y(new_n6808_));
  NOR2  g06423(.A(new_n6808_), .B(new_n820_), .Y(new_n6809_));
  NOR2  g06424(.A(new_n6809_), .B(new_n824_), .Y(new_n6810_));
  NOR2  g06425(.A(new_n6810_), .B(new_n829_), .Y(new_n6811_));
  NOR2  g06426(.A(new_n6811_), .B(new_n833_), .Y(new_n6812_));
  NOR2  g06427(.A(new_n6812_), .B(new_n838_), .Y(new_n6813_));
  NOR2  g06428(.A(new_n6813_), .B(new_n842_), .Y(new_n6814_));
  NOR2  g06429(.A(new_n6814_), .B(new_n847_), .Y(new_n6815_));
  NOR2  g06430(.A(new_n6815_), .B(new_n851_), .Y(new_n6816_));
  NOR2  g06431(.A(new_n6816_), .B(new_n856_), .Y(new_n6817_));
  NOR2  g06432(.A(new_n6817_), .B(new_n860_), .Y(new_n6818_));
  NOR2  g06433(.A(new_n6818_), .B(new_n865_), .Y(new_n6819_));
  NOR2  g06434(.A(new_n6819_), .B(new_n869_), .Y(new_n6820_));
  NOR2  g06435(.A(new_n6820_), .B(new_n874_), .Y(new_n6821_));
  NOR2  g06436(.A(new_n6821_), .B(new_n878_), .Y(new_n6822_));
  NOR2  g06437(.A(new_n6822_), .B(new_n883_), .Y(new_n6823_));
  NOR2  g06438(.A(new_n6823_), .B(new_n887_), .Y(new_n6824_));
  NOR2  g06439(.A(new_n6824_), .B(new_n892_), .Y(new_n6825_));
  NOR2  g06440(.A(new_n6825_), .B(new_n896_), .Y(new_n6826_));
  NOR2  g06441(.A(new_n6826_), .B(new_n901_), .Y(new_n6827_));
  NOR2  g06442(.A(new_n6827_), .B(new_n905_), .Y(new_n6828_));
  NOR2  g06443(.A(new_n6828_), .B(new_n910_), .Y(new_n6829_));
  NOR2  g06444(.A(new_n6829_), .B(new_n914_), .Y(new_n6830_));
  NOR2  g06445(.A(new_n6830_), .B(new_n919_), .Y(new_n6831_));
  NOR2  g06446(.A(new_n6831_), .B(new_n923_), .Y(new_n6832_));
  NOR2  g06447(.A(new_n6832_), .B(new_n928_), .Y(new_n6833_));
  NOR2  g06448(.A(new_n6833_), .B(new_n932_), .Y(new_n6834_));
  NOR2  g06449(.A(new_n6834_), .B(new_n937_), .Y(new_n6835_));
  NOR2  g06450(.A(new_n6835_), .B(new_n941_), .Y(new_n6836_));
  NOR2  g06451(.A(new_n6836_), .B(new_n946_), .Y(new_n6837_));
  NOR2  g06452(.A(new_n6837_), .B(new_n950_), .Y(new_n6838_));
  NOR2  g06453(.A(new_n6838_), .B(new_n955_), .Y(new_n6839_));
  NOR2  g06454(.A(new_n6839_), .B(new_n959_), .Y(new_n6840_));
  NOR2  g06455(.A(new_n6840_), .B(new_n964_), .Y(new_n6841_));
  NOR2  g06456(.A(new_n6841_), .B(new_n968_), .Y(new_n6842_));
  NOR2  g06457(.A(new_n6842_), .B(new_n973_), .Y(new_n6843_));
  NOR2  g06458(.A(new_n6843_), .B(new_n977_), .Y(new_n6844_));
  NOR2  g06459(.A(new_n6844_), .B(new_n982_), .Y(new_n6845_));
  NOR2  g06460(.A(new_n6845_), .B(new_n986_), .Y(new_n6846_));
  NOR2  g06461(.A(new_n6846_), .B(new_n991_), .Y(new_n6847_));
  NAND2 g06462(.A(new_n993_), .B(\req[63] ), .Y(new_n6848_));
  NOR2  g06463(.A(new_n6848_), .B(new_n6847_), .Y(\grant[63] ));
  INV   g06464(.A(new_n1003_), .Y(new_n6850_));
  NOR2  g06465(.A(new_n1358_), .B(new_n6850_), .Y(new_n6851_));
  NOR2  g06466(.A(new_n6851_), .B(new_n1009_), .Y(new_n6852_));
  NOR2  g06467(.A(new_n6852_), .B(new_n1013_), .Y(new_n6853_));
  NOR2  g06468(.A(new_n6853_), .B(new_n1018_), .Y(new_n6854_));
  NOR2  g06469(.A(new_n6854_), .B(new_n1022_), .Y(new_n6855_));
  NOR2  g06470(.A(new_n6855_), .B(new_n1027_), .Y(new_n6856_));
  NOR2  g06471(.A(new_n6856_), .B(new_n1031_), .Y(new_n6857_));
  NOR2  g06472(.A(new_n6857_), .B(new_n1036_), .Y(new_n6858_));
  NOR2  g06473(.A(new_n6858_), .B(new_n1040_), .Y(new_n6859_));
  NOR2  g06474(.A(new_n6859_), .B(new_n1045_), .Y(new_n6860_));
  NOR2  g06475(.A(new_n6860_), .B(new_n1049_), .Y(new_n6861_));
  NOR2  g06476(.A(new_n6861_), .B(new_n1054_), .Y(new_n6862_));
  NOR2  g06477(.A(new_n6862_), .B(new_n1058_), .Y(new_n6863_));
  NOR2  g06478(.A(new_n6863_), .B(new_n1063_), .Y(new_n6864_));
  NOR2  g06479(.A(new_n6864_), .B(new_n1067_), .Y(new_n6865_));
  NOR2  g06480(.A(new_n6865_), .B(new_n1072_), .Y(new_n6866_));
  NOR2  g06481(.A(new_n6866_), .B(new_n1076_), .Y(new_n6867_));
  NOR2  g06482(.A(new_n6867_), .B(new_n1081_), .Y(new_n6868_));
  NOR2  g06483(.A(new_n6868_), .B(new_n1085_), .Y(new_n6869_));
  NOR2  g06484(.A(new_n6869_), .B(new_n1090_), .Y(new_n6870_));
  NOR2  g06485(.A(new_n6870_), .B(new_n1094_), .Y(new_n6871_));
  NOR2  g06486(.A(new_n6871_), .B(new_n1099_), .Y(new_n6872_));
  NOR2  g06487(.A(new_n6872_), .B(new_n1103_), .Y(new_n6873_));
  NOR2  g06488(.A(new_n6873_), .B(new_n1108_), .Y(new_n6874_));
  NOR2  g06489(.A(new_n6874_), .B(new_n1112_), .Y(new_n6875_));
  NOR2  g06490(.A(new_n6875_), .B(new_n1117_), .Y(new_n6876_));
  NOR2  g06491(.A(new_n6876_), .B(new_n1121_), .Y(new_n6877_));
  NOR2  g06492(.A(new_n6877_), .B(new_n1126_), .Y(new_n6878_));
  NOR2  g06493(.A(new_n6878_), .B(new_n1130_), .Y(new_n6879_));
  NOR2  g06494(.A(new_n6879_), .B(new_n1135_), .Y(new_n6880_));
  NOR2  g06495(.A(new_n6880_), .B(new_n1139_), .Y(new_n6881_));
  NOR2  g06496(.A(new_n6881_), .B(new_n1144_), .Y(new_n6882_));
  NOR2  g06497(.A(new_n6882_), .B(new_n1148_), .Y(new_n6883_));
  NOR2  g06498(.A(new_n6883_), .B(new_n1153_), .Y(new_n6884_));
  NOR2  g06499(.A(new_n6884_), .B(new_n1157_), .Y(new_n6885_));
  NOR2  g06500(.A(new_n6885_), .B(new_n1162_), .Y(new_n6886_));
  NOR2  g06501(.A(new_n6886_), .B(new_n1166_), .Y(new_n6887_));
  NOR2  g06502(.A(new_n6887_), .B(new_n1171_), .Y(new_n6888_));
  NOR2  g06503(.A(new_n6888_), .B(new_n1175_), .Y(new_n6889_));
  NOR2  g06504(.A(new_n6889_), .B(new_n1180_), .Y(new_n6890_));
  NOR2  g06505(.A(new_n6890_), .B(new_n1184_), .Y(new_n6891_));
  NOR2  g06506(.A(new_n6891_), .B(new_n1189_), .Y(new_n6892_));
  NOR2  g06507(.A(new_n6892_), .B(new_n1707_), .Y(new_n6893_));
  NOR2  g06508(.A(new_n6893_), .B(new_n1709_), .Y(new_n6894_));
  NOR2  g06509(.A(new_n6894_), .B(new_n1973_), .Y(new_n6895_));
  NOR2  g06510(.A(new_n6895_), .B(new_n1199_), .Y(new_n6896_));
  NOR2  g06511(.A(new_n6896_), .B(new_n1203_), .Y(new_n6897_));
  NOR2  g06512(.A(new_n6897_), .B(new_n1207_), .Y(new_n6898_));
  NOR2  g06513(.A(new_n6898_), .B(new_n1211_), .Y(new_n6899_));
  NOR2  g06514(.A(new_n6899_), .B(new_n1215_), .Y(new_n6900_));
  NOR2  g06515(.A(new_n6900_), .B(new_n1219_), .Y(new_n6901_));
  NOR2  g06516(.A(new_n6901_), .B(new_n1223_), .Y(new_n6902_));
  NOR2  g06517(.A(new_n6902_), .B(new_n1227_), .Y(new_n6903_));
  NOR2  g06518(.A(new_n6903_), .B(new_n1231_), .Y(new_n6904_));
  NOR2  g06519(.A(new_n6904_), .B(new_n1235_), .Y(new_n6905_));
  NOR2  g06520(.A(new_n6905_), .B(new_n1239_), .Y(new_n6906_));
  NOR2  g06521(.A(new_n6906_), .B(new_n1243_), .Y(new_n6907_));
  NOR2  g06522(.A(new_n6907_), .B(new_n1247_), .Y(new_n6908_));
  NOR2  g06523(.A(new_n6908_), .B(new_n1251_), .Y(new_n6909_));
  NOR2  g06524(.A(new_n6909_), .B(new_n1255_), .Y(new_n6910_));
  NOR2  g06525(.A(new_n6910_), .B(new_n1259_), .Y(new_n6911_));
  NOR2  g06526(.A(new_n6911_), .B(new_n1263_), .Y(new_n6912_));
  NOR2  g06527(.A(new_n6912_), .B(new_n1267_), .Y(new_n6913_));
  NOR2  g06528(.A(new_n6913_), .B(new_n1271_), .Y(new_n6914_));
  NOR2  g06529(.A(new_n6914_), .B(new_n1275_), .Y(new_n6915_));
  NOR2  g06530(.A(new_n6915_), .B(new_n1279_), .Y(new_n6916_));
  NOR2  g06531(.A(new_n6916_), .B(new_n1283_), .Y(new_n6917_));
  NOR2  g06532(.A(new_n6917_), .B(new_n1287_), .Y(new_n6918_));
  NOR2  g06533(.A(new_n6918_), .B(new_n1291_), .Y(new_n6919_));
  NOR2  g06534(.A(new_n6919_), .B(new_n1295_), .Y(new_n6920_));
  NOR2  g06535(.A(new_n6920_), .B(new_n1299_), .Y(new_n6921_));
  NOR2  g06536(.A(new_n6921_), .B(new_n1303_), .Y(new_n6922_));
  NOR2  g06537(.A(new_n6922_), .B(new_n1307_), .Y(new_n6923_));
  NOR2  g06538(.A(new_n6923_), .B(new_n1311_), .Y(new_n6924_));
  NOR2  g06539(.A(new_n6924_), .B(new_n1315_), .Y(new_n6925_));
  NOR2  g06540(.A(new_n6925_), .B(new_n1319_), .Y(new_n6926_));
  NOR2  g06541(.A(new_n6926_), .B(new_n1323_), .Y(new_n6927_));
  NOR2  g06542(.A(new_n6927_), .B(new_n1327_), .Y(new_n6928_));
  NOR2  g06543(.A(new_n6928_), .B(new_n1331_), .Y(new_n6929_));
  NOR2  g06544(.A(new_n6929_), .B(new_n1335_), .Y(new_n6930_));
  NOR2  g06545(.A(new_n6930_), .B(new_n1339_), .Y(new_n6931_));
  NOR2  g06546(.A(new_n6931_), .B(new_n1343_), .Y(new_n6932_));
  NOR2  g06547(.A(new_n6932_), .B(new_n1347_), .Y(new_n6933_));
  NOR2  g06548(.A(new_n6933_), .B(new_n1351_), .Y(new_n6934_));
  NAND2 g06549(.A(new_n1353_), .B(\req[64] ), .Y(new_n6935_));
  NOR2  g06550(.A(new_n6935_), .B(new_n6934_), .Y(\grant[64] ));
  INV   g06551(.A(new_n1362_), .Y(new_n6937_));
  NOR2  g06552(.A(new_n6937_), .B(new_n605_), .Y(new_n6938_));
  NOR2  g06553(.A(new_n6938_), .B(new_n1367_), .Y(new_n6939_));
  NOR2  g06554(.A(new_n6939_), .B(new_n1371_), .Y(new_n6940_));
  NOR2  g06555(.A(new_n6940_), .B(new_n1375_), .Y(new_n6941_));
  NOR2  g06556(.A(new_n6941_), .B(new_n1379_), .Y(new_n6942_));
  NOR2  g06557(.A(new_n6942_), .B(new_n1383_), .Y(new_n6943_));
  NOR2  g06558(.A(new_n6943_), .B(new_n1387_), .Y(new_n6944_));
  NOR2  g06559(.A(new_n6944_), .B(new_n1391_), .Y(new_n6945_));
  NOR2  g06560(.A(new_n6945_), .B(new_n1395_), .Y(new_n6946_));
  NOR2  g06561(.A(new_n6946_), .B(new_n1399_), .Y(new_n6947_));
  NOR2  g06562(.A(new_n6947_), .B(new_n1403_), .Y(new_n6948_));
  NOR2  g06563(.A(new_n6948_), .B(new_n1407_), .Y(new_n6949_));
  NOR2  g06564(.A(new_n6949_), .B(new_n1411_), .Y(new_n6950_));
  NOR2  g06565(.A(new_n6950_), .B(new_n1415_), .Y(new_n6951_));
  NOR2  g06566(.A(new_n6951_), .B(new_n1419_), .Y(new_n6952_));
  NOR2  g06567(.A(new_n6952_), .B(new_n1423_), .Y(new_n6953_));
  NOR2  g06568(.A(new_n6953_), .B(new_n1427_), .Y(new_n6954_));
  NOR2  g06569(.A(new_n6954_), .B(new_n1431_), .Y(new_n6955_));
  NOR2  g06570(.A(new_n6955_), .B(new_n1435_), .Y(new_n6956_));
  NOR2  g06571(.A(new_n6956_), .B(new_n1439_), .Y(new_n6957_));
  NOR2  g06572(.A(new_n6957_), .B(new_n1443_), .Y(new_n6958_));
  NOR2  g06573(.A(new_n6958_), .B(new_n1447_), .Y(new_n6959_));
  NOR2  g06574(.A(new_n6959_), .B(new_n1451_), .Y(new_n6960_));
  NOR2  g06575(.A(new_n6960_), .B(new_n1455_), .Y(new_n6961_));
  NOR2  g06576(.A(new_n6961_), .B(new_n1459_), .Y(new_n6962_));
  NOR2  g06577(.A(new_n6962_), .B(new_n1463_), .Y(new_n6963_));
  NOR2  g06578(.A(new_n6963_), .B(new_n1467_), .Y(new_n6964_));
  NOR2  g06579(.A(new_n6964_), .B(new_n1471_), .Y(new_n6965_));
  NOR2  g06580(.A(new_n6965_), .B(new_n1475_), .Y(new_n6966_));
  NOR2  g06581(.A(new_n6966_), .B(new_n1479_), .Y(new_n6967_));
  NOR2  g06582(.A(new_n6967_), .B(new_n1483_), .Y(new_n6968_));
  NOR2  g06583(.A(new_n6968_), .B(new_n1487_), .Y(new_n6969_));
  NOR2  g06584(.A(new_n6969_), .B(new_n1491_), .Y(new_n6970_));
  NOR2  g06585(.A(new_n6970_), .B(new_n1495_), .Y(new_n6971_));
  NOR2  g06586(.A(new_n6971_), .B(new_n1499_), .Y(new_n6972_));
  NOR2  g06587(.A(new_n6972_), .B(new_n1503_), .Y(new_n6973_));
  NOR2  g06588(.A(new_n6973_), .B(new_n1507_), .Y(new_n6974_));
  NOR2  g06589(.A(new_n6974_), .B(new_n1511_), .Y(new_n6975_));
  NOR2  g06590(.A(new_n6975_), .B(new_n1515_), .Y(new_n6976_));
  NOR2  g06591(.A(new_n6976_), .B(new_n1519_), .Y(new_n6977_));
  NOR2  g06592(.A(new_n6977_), .B(new_n1523_), .Y(new_n6978_));
  NOR2  g06593(.A(new_n6978_), .B(new_n1527_), .Y(new_n6979_));
  NOR2  g06594(.A(new_n6979_), .B(new_n1797_), .Y(new_n6980_));
  NOR2  g06595(.A(new_n6980_), .B(new_n396_), .Y(new_n6981_));
  NOR2  g06596(.A(new_n6981_), .B(new_n400_), .Y(new_n6982_));
  NOR2  g06597(.A(new_n6982_), .B(new_n406_), .Y(new_n6983_));
  NOR2  g06598(.A(new_n6983_), .B(new_n410_), .Y(new_n6984_));
  NOR2  g06599(.A(new_n6984_), .B(new_n416_), .Y(new_n6985_));
  NOR2  g06600(.A(new_n6985_), .B(new_n420_), .Y(new_n6986_));
  NOR2  g06601(.A(new_n6986_), .B(new_n426_), .Y(new_n6987_));
  NOR2  g06602(.A(new_n6987_), .B(new_n430_), .Y(new_n6988_));
  NOR2  g06603(.A(new_n6988_), .B(new_n436_), .Y(new_n6989_));
  NOR2  g06604(.A(new_n6989_), .B(new_n440_), .Y(new_n6990_));
  NOR2  g06605(.A(new_n6990_), .B(new_n446_), .Y(new_n6991_));
  NOR2  g06606(.A(new_n6991_), .B(new_n450_), .Y(new_n6992_));
  NOR2  g06607(.A(new_n6992_), .B(new_n456_), .Y(new_n6993_));
  NOR2  g06608(.A(new_n6993_), .B(new_n460_), .Y(new_n6994_));
  NOR2  g06609(.A(new_n6994_), .B(new_n466_), .Y(new_n6995_));
  NOR2  g06610(.A(new_n6995_), .B(new_n470_), .Y(new_n6996_));
  NOR2  g06611(.A(new_n6996_), .B(new_n476_), .Y(new_n6997_));
  NOR2  g06612(.A(new_n6997_), .B(new_n480_), .Y(new_n6998_));
  NOR2  g06613(.A(new_n6998_), .B(new_n486_), .Y(new_n6999_));
  NOR2  g06614(.A(new_n6999_), .B(new_n490_), .Y(new_n7000_));
  NOR2  g06615(.A(new_n7000_), .B(new_n496_), .Y(new_n7001_));
  NOR2  g06616(.A(new_n7001_), .B(new_n500_), .Y(new_n7002_));
  NOR2  g06617(.A(new_n7002_), .B(new_n506_), .Y(new_n7003_));
  NOR2  g06618(.A(new_n7003_), .B(new_n510_), .Y(new_n7004_));
  NOR2  g06619(.A(new_n7004_), .B(new_n516_), .Y(new_n7005_));
  NOR2  g06620(.A(new_n7005_), .B(new_n520_), .Y(new_n7006_));
  NOR2  g06621(.A(new_n7006_), .B(new_n526_), .Y(new_n7007_));
  NOR2  g06622(.A(new_n7007_), .B(new_n530_), .Y(new_n7008_));
  NOR2  g06623(.A(new_n7008_), .B(new_n536_), .Y(new_n7009_));
  NOR2  g06624(.A(new_n7009_), .B(new_n540_), .Y(new_n7010_));
  NOR2  g06625(.A(new_n7010_), .B(new_n546_), .Y(new_n7011_));
  NOR2  g06626(.A(new_n7011_), .B(new_n550_), .Y(new_n7012_));
  NOR2  g06627(.A(new_n7012_), .B(new_n556_), .Y(new_n7013_));
  NOR2  g06628(.A(new_n7013_), .B(new_n560_), .Y(new_n7014_));
  NOR2  g06629(.A(new_n7014_), .B(new_n566_), .Y(new_n7015_));
  NOR2  g06630(.A(new_n7015_), .B(new_n570_), .Y(new_n7016_));
  NOR2  g06631(.A(new_n7016_), .B(new_n576_), .Y(new_n7017_));
  NOR2  g06632(.A(new_n7017_), .B(new_n580_), .Y(new_n7018_));
  NOR2  g06633(.A(new_n7018_), .B(new_n586_), .Y(new_n7019_));
  NOR2  g06634(.A(new_n7019_), .B(new_n590_), .Y(new_n7020_));
  NOR2  g06635(.A(new_n7020_), .B(new_n596_), .Y(new_n7021_));
  NAND2 g06636(.A(new_n598_), .B(\req[65] ), .Y(new_n7022_));
  NOR2  g06637(.A(new_n7022_), .B(new_n7021_), .Y(\grant[65] ));
  INV   g06638(.A(new_n609_), .Y(new_n7024_));
  NOR2  g06639(.A(new_n1008_), .B(new_n7024_), .Y(new_n7025_));
  NOR2  g06640(.A(new_n7025_), .B(new_n616_), .Y(new_n7026_));
  NOR2  g06641(.A(new_n7026_), .B(new_n620_), .Y(new_n7027_));
  NOR2  g06642(.A(new_n7027_), .B(new_n626_), .Y(new_n7028_));
  NOR2  g06643(.A(new_n7028_), .B(new_n630_), .Y(new_n7029_));
  NOR2  g06644(.A(new_n7029_), .B(new_n636_), .Y(new_n7030_));
  NOR2  g06645(.A(new_n7030_), .B(new_n640_), .Y(new_n7031_));
  NOR2  g06646(.A(new_n7031_), .B(new_n646_), .Y(new_n7032_));
  NOR2  g06647(.A(new_n7032_), .B(new_n650_), .Y(new_n7033_));
  NOR2  g06648(.A(new_n7033_), .B(new_n656_), .Y(new_n7034_));
  NOR2  g06649(.A(new_n7034_), .B(new_n660_), .Y(new_n7035_));
  NOR2  g06650(.A(new_n7035_), .B(new_n666_), .Y(new_n7036_));
  NOR2  g06651(.A(new_n7036_), .B(new_n670_), .Y(new_n7037_));
  NOR2  g06652(.A(new_n7037_), .B(new_n676_), .Y(new_n7038_));
  NOR2  g06653(.A(new_n7038_), .B(new_n680_), .Y(new_n7039_));
  NOR2  g06654(.A(new_n7039_), .B(new_n686_), .Y(new_n7040_));
  NOR2  g06655(.A(new_n7040_), .B(new_n690_), .Y(new_n7041_));
  NOR2  g06656(.A(new_n7041_), .B(new_n696_), .Y(new_n7042_));
  NOR2  g06657(.A(new_n7042_), .B(new_n700_), .Y(new_n7043_));
  NOR2  g06658(.A(new_n7043_), .B(new_n706_), .Y(new_n7044_));
  NOR2  g06659(.A(new_n7044_), .B(new_n710_), .Y(new_n7045_));
  NOR2  g06660(.A(new_n7045_), .B(new_n716_), .Y(new_n7046_));
  NOR2  g06661(.A(new_n7046_), .B(new_n720_), .Y(new_n7047_));
  NOR2  g06662(.A(new_n7047_), .B(new_n726_), .Y(new_n7048_));
  NOR2  g06663(.A(new_n7048_), .B(new_n730_), .Y(new_n7049_));
  NOR2  g06664(.A(new_n7049_), .B(new_n736_), .Y(new_n7050_));
  NOR2  g06665(.A(new_n7050_), .B(new_n740_), .Y(new_n7051_));
  NOR2  g06666(.A(new_n7051_), .B(new_n746_), .Y(new_n7052_));
  NOR2  g06667(.A(new_n7052_), .B(new_n750_), .Y(new_n7053_));
  NOR2  g06668(.A(new_n7053_), .B(new_n756_), .Y(new_n7054_));
  NOR2  g06669(.A(new_n7054_), .B(new_n760_), .Y(new_n7055_));
  NOR2  g06670(.A(new_n7055_), .B(new_n766_), .Y(new_n7056_));
  NOR2  g06671(.A(new_n7056_), .B(new_n770_), .Y(new_n7057_));
  NOR2  g06672(.A(new_n7057_), .B(new_n776_), .Y(new_n7058_));
  NOR2  g06673(.A(new_n7058_), .B(new_n780_), .Y(new_n7059_));
  NOR2  g06674(.A(new_n7059_), .B(new_n786_), .Y(new_n7060_));
  NOR2  g06675(.A(new_n7060_), .B(new_n790_), .Y(new_n7061_));
  NOR2  g06676(.A(new_n7061_), .B(new_n796_), .Y(new_n7062_));
  NOR2  g06677(.A(new_n7062_), .B(new_n800_), .Y(new_n7063_));
  NOR2  g06678(.A(new_n7063_), .B(new_n806_), .Y(new_n7064_));
  NOR2  g06679(.A(new_n7064_), .B(new_n1616_), .Y(new_n7065_));
  NOR2  g06680(.A(new_n7065_), .B(new_n1618_), .Y(new_n7066_));
  NOR2  g06681(.A(new_n7066_), .B(new_n1885_), .Y(new_n7067_));
  NOR2  g06682(.A(new_n7067_), .B(new_n820_), .Y(new_n7068_));
  NOR2  g06683(.A(new_n7068_), .B(new_n824_), .Y(new_n7069_));
  NOR2  g06684(.A(new_n7069_), .B(new_n829_), .Y(new_n7070_));
  NOR2  g06685(.A(new_n7070_), .B(new_n833_), .Y(new_n7071_));
  NOR2  g06686(.A(new_n7071_), .B(new_n838_), .Y(new_n7072_));
  NOR2  g06687(.A(new_n7072_), .B(new_n842_), .Y(new_n7073_));
  NOR2  g06688(.A(new_n7073_), .B(new_n847_), .Y(new_n7074_));
  NOR2  g06689(.A(new_n7074_), .B(new_n851_), .Y(new_n7075_));
  NOR2  g06690(.A(new_n7075_), .B(new_n856_), .Y(new_n7076_));
  NOR2  g06691(.A(new_n7076_), .B(new_n860_), .Y(new_n7077_));
  NOR2  g06692(.A(new_n7077_), .B(new_n865_), .Y(new_n7078_));
  NOR2  g06693(.A(new_n7078_), .B(new_n869_), .Y(new_n7079_));
  NOR2  g06694(.A(new_n7079_), .B(new_n874_), .Y(new_n7080_));
  NOR2  g06695(.A(new_n7080_), .B(new_n878_), .Y(new_n7081_));
  NOR2  g06696(.A(new_n7081_), .B(new_n883_), .Y(new_n7082_));
  NOR2  g06697(.A(new_n7082_), .B(new_n887_), .Y(new_n7083_));
  NOR2  g06698(.A(new_n7083_), .B(new_n892_), .Y(new_n7084_));
  NOR2  g06699(.A(new_n7084_), .B(new_n896_), .Y(new_n7085_));
  NOR2  g06700(.A(new_n7085_), .B(new_n901_), .Y(new_n7086_));
  NOR2  g06701(.A(new_n7086_), .B(new_n905_), .Y(new_n7087_));
  NOR2  g06702(.A(new_n7087_), .B(new_n910_), .Y(new_n7088_));
  NOR2  g06703(.A(new_n7088_), .B(new_n914_), .Y(new_n7089_));
  NOR2  g06704(.A(new_n7089_), .B(new_n919_), .Y(new_n7090_));
  NOR2  g06705(.A(new_n7090_), .B(new_n923_), .Y(new_n7091_));
  NOR2  g06706(.A(new_n7091_), .B(new_n928_), .Y(new_n7092_));
  NOR2  g06707(.A(new_n7092_), .B(new_n932_), .Y(new_n7093_));
  NOR2  g06708(.A(new_n7093_), .B(new_n937_), .Y(new_n7094_));
  NOR2  g06709(.A(new_n7094_), .B(new_n941_), .Y(new_n7095_));
  NOR2  g06710(.A(new_n7095_), .B(new_n946_), .Y(new_n7096_));
  NOR2  g06711(.A(new_n7096_), .B(new_n950_), .Y(new_n7097_));
  NOR2  g06712(.A(new_n7097_), .B(new_n955_), .Y(new_n7098_));
  NOR2  g06713(.A(new_n7098_), .B(new_n959_), .Y(new_n7099_));
  NOR2  g06714(.A(new_n7099_), .B(new_n964_), .Y(new_n7100_));
  NOR2  g06715(.A(new_n7100_), .B(new_n968_), .Y(new_n7101_));
  NOR2  g06716(.A(new_n7101_), .B(new_n973_), .Y(new_n7102_));
  NOR2  g06717(.A(new_n7102_), .B(new_n977_), .Y(new_n7103_));
  NOR2  g06718(.A(new_n7103_), .B(new_n982_), .Y(new_n7104_));
  NOR2  g06719(.A(new_n7104_), .B(new_n986_), .Y(new_n7105_));
  NOR2  g06720(.A(new_n7105_), .B(new_n991_), .Y(new_n7106_));
  NOR2  g06721(.A(new_n7106_), .B(new_n995_), .Y(new_n7107_));
  NOR2  g06722(.A(new_n7107_), .B(new_n1000_), .Y(new_n7108_));
  NAND2 g06723(.A(new_n1002_), .B(\req[66] ), .Y(new_n7109_));
  NOR2  g06724(.A(new_n7109_), .B(new_n7108_), .Y(\grant[66] ));
  INV   g06725(.A(new_n1012_), .Y(new_n7111_));
  NOR2  g06726(.A(new_n1366_), .B(new_n7111_), .Y(new_n7112_));
  NOR2  g06727(.A(new_n7112_), .B(new_n1018_), .Y(new_n7113_));
  NOR2  g06728(.A(new_n7113_), .B(new_n1022_), .Y(new_n7114_));
  NOR2  g06729(.A(new_n7114_), .B(new_n1027_), .Y(new_n7115_));
  NOR2  g06730(.A(new_n7115_), .B(new_n1031_), .Y(new_n7116_));
  NOR2  g06731(.A(new_n7116_), .B(new_n1036_), .Y(new_n7117_));
  NOR2  g06732(.A(new_n7117_), .B(new_n1040_), .Y(new_n7118_));
  NOR2  g06733(.A(new_n7118_), .B(new_n1045_), .Y(new_n7119_));
  NOR2  g06734(.A(new_n7119_), .B(new_n1049_), .Y(new_n7120_));
  NOR2  g06735(.A(new_n7120_), .B(new_n1054_), .Y(new_n7121_));
  NOR2  g06736(.A(new_n7121_), .B(new_n1058_), .Y(new_n7122_));
  NOR2  g06737(.A(new_n7122_), .B(new_n1063_), .Y(new_n7123_));
  NOR2  g06738(.A(new_n7123_), .B(new_n1067_), .Y(new_n7124_));
  NOR2  g06739(.A(new_n7124_), .B(new_n1072_), .Y(new_n7125_));
  NOR2  g06740(.A(new_n7125_), .B(new_n1076_), .Y(new_n7126_));
  NOR2  g06741(.A(new_n7126_), .B(new_n1081_), .Y(new_n7127_));
  NOR2  g06742(.A(new_n7127_), .B(new_n1085_), .Y(new_n7128_));
  NOR2  g06743(.A(new_n7128_), .B(new_n1090_), .Y(new_n7129_));
  NOR2  g06744(.A(new_n7129_), .B(new_n1094_), .Y(new_n7130_));
  NOR2  g06745(.A(new_n7130_), .B(new_n1099_), .Y(new_n7131_));
  NOR2  g06746(.A(new_n7131_), .B(new_n1103_), .Y(new_n7132_));
  NOR2  g06747(.A(new_n7132_), .B(new_n1108_), .Y(new_n7133_));
  NOR2  g06748(.A(new_n7133_), .B(new_n1112_), .Y(new_n7134_));
  NOR2  g06749(.A(new_n7134_), .B(new_n1117_), .Y(new_n7135_));
  NOR2  g06750(.A(new_n7135_), .B(new_n1121_), .Y(new_n7136_));
  NOR2  g06751(.A(new_n7136_), .B(new_n1126_), .Y(new_n7137_));
  NOR2  g06752(.A(new_n7137_), .B(new_n1130_), .Y(new_n7138_));
  NOR2  g06753(.A(new_n7138_), .B(new_n1135_), .Y(new_n7139_));
  NOR2  g06754(.A(new_n7139_), .B(new_n1139_), .Y(new_n7140_));
  NOR2  g06755(.A(new_n7140_), .B(new_n1144_), .Y(new_n7141_));
  NOR2  g06756(.A(new_n7141_), .B(new_n1148_), .Y(new_n7142_));
  NOR2  g06757(.A(new_n7142_), .B(new_n1153_), .Y(new_n7143_));
  NOR2  g06758(.A(new_n7143_), .B(new_n1157_), .Y(new_n7144_));
  NOR2  g06759(.A(new_n7144_), .B(new_n1162_), .Y(new_n7145_));
  NOR2  g06760(.A(new_n7145_), .B(new_n1166_), .Y(new_n7146_));
  NOR2  g06761(.A(new_n7146_), .B(new_n1171_), .Y(new_n7147_));
  NOR2  g06762(.A(new_n7147_), .B(new_n1175_), .Y(new_n7148_));
  NOR2  g06763(.A(new_n7148_), .B(new_n1180_), .Y(new_n7149_));
  NOR2  g06764(.A(new_n7149_), .B(new_n1184_), .Y(new_n7150_));
  NOR2  g06765(.A(new_n7150_), .B(new_n1189_), .Y(new_n7151_));
  NOR2  g06766(.A(new_n7151_), .B(new_n1707_), .Y(new_n7152_));
  NOR2  g06767(.A(new_n7152_), .B(new_n1709_), .Y(new_n7153_));
  NOR2  g06768(.A(new_n7153_), .B(new_n1973_), .Y(new_n7154_));
  NOR2  g06769(.A(new_n7154_), .B(new_n1199_), .Y(new_n7155_));
  NOR2  g06770(.A(new_n7155_), .B(new_n1203_), .Y(new_n7156_));
  NOR2  g06771(.A(new_n7156_), .B(new_n1207_), .Y(new_n7157_));
  NOR2  g06772(.A(new_n7157_), .B(new_n1211_), .Y(new_n7158_));
  NOR2  g06773(.A(new_n7158_), .B(new_n1215_), .Y(new_n7159_));
  NOR2  g06774(.A(new_n7159_), .B(new_n1219_), .Y(new_n7160_));
  NOR2  g06775(.A(new_n7160_), .B(new_n1223_), .Y(new_n7161_));
  NOR2  g06776(.A(new_n7161_), .B(new_n1227_), .Y(new_n7162_));
  NOR2  g06777(.A(new_n7162_), .B(new_n1231_), .Y(new_n7163_));
  NOR2  g06778(.A(new_n7163_), .B(new_n1235_), .Y(new_n7164_));
  NOR2  g06779(.A(new_n7164_), .B(new_n1239_), .Y(new_n7165_));
  NOR2  g06780(.A(new_n7165_), .B(new_n1243_), .Y(new_n7166_));
  NOR2  g06781(.A(new_n7166_), .B(new_n1247_), .Y(new_n7167_));
  NOR2  g06782(.A(new_n7167_), .B(new_n1251_), .Y(new_n7168_));
  NOR2  g06783(.A(new_n7168_), .B(new_n1255_), .Y(new_n7169_));
  NOR2  g06784(.A(new_n7169_), .B(new_n1259_), .Y(new_n7170_));
  NOR2  g06785(.A(new_n7170_), .B(new_n1263_), .Y(new_n7171_));
  NOR2  g06786(.A(new_n7171_), .B(new_n1267_), .Y(new_n7172_));
  NOR2  g06787(.A(new_n7172_), .B(new_n1271_), .Y(new_n7173_));
  NOR2  g06788(.A(new_n7173_), .B(new_n1275_), .Y(new_n7174_));
  NOR2  g06789(.A(new_n7174_), .B(new_n1279_), .Y(new_n7175_));
  NOR2  g06790(.A(new_n7175_), .B(new_n1283_), .Y(new_n7176_));
  NOR2  g06791(.A(new_n7176_), .B(new_n1287_), .Y(new_n7177_));
  NOR2  g06792(.A(new_n7177_), .B(new_n1291_), .Y(new_n7178_));
  NOR2  g06793(.A(new_n7178_), .B(new_n1295_), .Y(new_n7179_));
  NOR2  g06794(.A(new_n7179_), .B(new_n1299_), .Y(new_n7180_));
  NOR2  g06795(.A(new_n7180_), .B(new_n1303_), .Y(new_n7181_));
  NOR2  g06796(.A(new_n7181_), .B(new_n1307_), .Y(new_n7182_));
  NOR2  g06797(.A(new_n7182_), .B(new_n1311_), .Y(new_n7183_));
  NOR2  g06798(.A(new_n7183_), .B(new_n1315_), .Y(new_n7184_));
  NOR2  g06799(.A(new_n7184_), .B(new_n1319_), .Y(new_n7185_));
  NOR2  g06800(.A(new_n7185_), .B(new_n1323_), .Y(new_n7186_));
  NOR2  g06801(.A(new_n7186_), .B(new_n1327_), .Y(new_n7187_));
  NOR2  g06802(.A(new_n7187_), .B(new_n1331_), .Y(new_n7188_));
  NOR2  g06803(.A(new_n7188_), .B(new_n1335_), .Y(new_n7189_));
  NOR2  g06804(.A(new_n7189_), .B(new_n1339_), .Y(new_n7190_));
  NOR2  g06805(.A(new_n7190_), .B(new_n1343_), .Y(new_n7191_));
  NOR2  g06806(.A(new_n7191_), .B(new_n1347_), .Y(new_n7192_));
  NOR2  g06807(.A(new_n7192_), .B(new_n1351_), .Y(new_n7193_));
  NOR2  g06808(.A(new_n7193_), .B(new_n1355_), .Y(new_n7194_));
  NOR2  g06809(.A(new_n7194_), .B(new_n1359_), .Y(new_n7195_));
  NAND2 g06810(.A(new_n1361_), .B(\req[67] ), .Y(new_n7196_));
  NOR2  g06811(.A(new_n7196_), .B(new_n7195_), .Y(\grant[67] ));
  INV   g06812(.A(new_n1370_), .Y(new_n7198_));
  NOR2  g06813(.A(new_n7198_), .B(new_n615_), .Y(new_n7199_));
  NOR2  g06814(.A(new_n7199_), .B(new_n1375_), .Y(new_n7200_));
  NOR2  g06815(.A(new_n7200_), .B(new_n1379_), .Y(new_n7201_));
  NOR2  g06816(.A(new_n7201_), .B(new_n1383_), .Y(new_n7202_));
  NOR2  g06817(.A(new_n7202_), .B(new_n1387_), .Y(new_n7203_));
  NOR2  g06818(.A(new_n7203_), .B(new_n1391_), .Y(new_n7204_));
  NOR2  g06819(.A(new_n7204_), .B(new_n1395_), .Y(new_n7205_));
  NOR2  g06820(.A(new_n7205_), .B(new_n1399_), .Y(new_n7206_));
  NOR2  g06821(.A(new_n7206_), .B(new_n1403_), .Y(new_n7207_));
  NOR2  g06822(.A(new_n7207_), .B(new_n1407_), .Y(new_n7208_));
  NOR2  g06823(.A(new_n7208_), .B(new_n1411_), .Y(new_n7209_));
  NOR2  g06824(.A(new_n7209_), .B(new_n1415_), .Y(new_n7210_));
  NOR2  g06825(.A(new_n7210_), .B(new_n1419_), .Y(new_n7211_));
  NOR2  g06826(.A(new_n7211_), .B(new_n1423_), .Y(new_n7212_));
  NOR2  g06827(.A(new_n7212_), .B(new_n1427_), .Y(new_n7213_));
  NOR2  g06828(.A(new_n7213_), .B(new_n1431_), .Y(new_n7214_));
  NOR2  g06829(.A(new_n7214_), .B(new_n1435_), .Y(new_n7215_));
  NOR2  g06830(.A(new_n7215_), .B(new_n1439_), .Y(new_n7216_));
  NOR2  g06831(.A(new_n7216_), .B(new_n1443_), .Y(new_n7217_));
  NOR2  g06832(.A(new_n7217_), .B(new_n1447_), .Y(new_n7218_));
  NOR2  g06833(.A(new_n7218_), .B(new_n1451_), .Y(new_n7219_));
  NOR2  g06834(.A(new_n7219_), .B(new_n1455_), .Y(new_n7220_));
  NOR2  g06835(.A(new_n7220_), .B(new_n1459_), .Y(new_n7221_));
  NOR2  g06836(.A(new_n7221_), .B(new_n1463_), .Y(new_n7222_));
  NOR2  g06837(.A(new_n7222_), .B(new_n1467_), .Y(new_n7223_));
  NOR2  g06838(.A(new_n7223_), .B(new_n1471_), .Y(new_n7224_));
  NOR2  g06839(.A(new_n7224_), .B(new_n1475_), .Y(new_n7225_));
  NOR2  g06840(.A(new_n7225_), .B(new_n1479_), .Y(new_n7226_));
  NOR2  g06841(.A(new_n7226_), .B(new_n1483_), .Y(new_n7227_));
  NOR2  g06842(.A(new_n7227_), .B(new_n1487_), .Y(new_n7228_));
  NOR2  g06843(.A(new_n7228_), .B(new_n1491_), .Y(new_n7229_));
  NOR2  g06844(.A(new_n7229_), .B(new_n1495_), .Y(new_n7230_));
  NOR2  g06845(.A(new_n7230_), .B(new_n1499_), .Y(new_n7231_));
  NOR2  g06846(.A(new_n7231_), .B(new_n1503_), .Y(new_n7232_));
  NOR2  g06847(.A(new_n7232_), .B(new_n1507_), .Y(new_n7233_));
  NOR2  g06848(.A(new_n7233_), .B(new_n1511_), .Y(new_n7234_));
  NOR2  g06849(.A(new_n7234_), .B(new_n1515_), .Y(new_n7235_));
  NOR2  g06850(.A(new_n7235_), .B(new_n1519_), .Y(new_n7236_));
  NOR2  g06851(.A(new_n7236_), .B(new_n1523_), .Y(new_n7237_));
  NOR2  g06852(.A(new_n7237_), .B(new_n1527_), .Y(new_n7238_));
  NOR2  g06853(.A(new_n7238_), .B(new_n1797_), .Y(new_n7239_));
  NOR2  g06854(.A(new_n7239_), .B(new_n396_), .Y(new_n7240_));
  NOR2  g06855(.A(new_n7240_), .B(new_n400_), .Y(new_n7241_));
  NOR2  g06856(.A(new_n7241_), .B(new_n406_), .Y(new_n7242_));
  NOR2  g06857(.A(new_n7242_), .B(new_n410_), .Y(new_n7243_));
  NOR2  g06858(.A(new_n7243_), .B(new_n416_), .Y(new_n7244_));
  NOR2  g06859(.A(new_n7244_), .B(new_n420_), .Y(new_n7245_));
  NOR2  g06860(.A(new_n7245_), .B(new_n426_), .Y(new_n7246_));
  NOR2  g06861(.A(new_n7246_), .B(new_n430_), .Y(new_n7247_));
  NOR2  g06862(.A(new_n7247_), .B(new_n436_), .Y(new_n7248_));
  NOR2  g06863(.A(new_n7248_), .B(new_n440_), .Y(new_n7249_));
  NOR2  g06864(.A(new_n7249_), .B(new_n446_), .Y(new_n7250_));
  NOR2  g06865(.A(new_n7250_), .B(new_n450_), .Y(new_n7251_));
  NOR2  g06866(.A(new_n7251_), .B(new_n456_), .Y(new_n7252_));
  NOR2  g06867(.A(new_n7252_), .B(new_n460_), .Y(new_n7253_));
  NOR2  g06868(.A(new_n7253_), .B(new_n466_), .Y(new_n7254_));
  NOR2  g06869(.A(new_n7254_), .B(new_n470_), .Y(new_n7255_));
  NOR2  g06870(.A(new_n7255_), .B(new_n476_), .Y(new_n7256_));
  NOR2  g06871(.A(new_n7256_), .B(new_n480_), .Y(new_n7257_));
  NOR2  g06872(.A(new_n7257_), .B(new_n486_), .Y(new_n7258_));
  NOR2  g06873(.A(new_n7258_), .B(new_n490_), .Y(new_n7259_));
  NOR2  g06874(.A(new_n7259_), .B(new_n496_), .Y(new_n7260_));
  NOR2  g06875(.A(new_n7260_), .B(new_n500_), .Y(new_n7261_));
  NOR2  g06876(.A(new_n7261_), .B(new_n506_), .Y(new_n7262_));
  NOR2  g06877(.A(new_n7262_), .B(new_n510_), .Y(new_n7263_));
  NOR2  g06878(.A(new_n7263_), .B(new_n516_), .Y(new_n7264_));
  NOR2  g06879(.A(new_n7264_), .B(new_n520_), .Y(new_n7265_));
  NOR2  g06880(.A(new_n7265_), .B(new_n526_), .Y(new_n7266_));
  NOR2  g06881(.A(new_n7266_), .B(new_n530_), .Y(new_n7267_));
  NOR2  g06882(.A(new_n7267_), .B(new_n536_), .Y(new_n7268_));
  NOR2  g06883(.A(new_n7268_), .B(new_n540_), .Y(new_n7269_));
  NOR2  g06884(.A(new_n7269_), .B(new_n546_), .Y(new_n7270_));
  NOR2  g06885(.A(new_n7270_), .B(new_n550_), .Y(new_n7271_));
  NOR2  g06886(.A(new_n7271_), .B(new_n556_), .Y(new_n7272_));
  NOR2  g06887(.A(new_n7272_), .B(new_n560_), .Y(new_n7273_));
  NOR2  g06888(.A(new_n7273_), .B(new_n566_), .Y(new_n7274_));
  NOR2  g06889(.A(new_n7274_), .B(new_n570_), .Y(new_n7275_));
  NOR2  g06890(.A(new_n7275_), .B(new_n576_), .Y(new_n7276_));
  NOR2  g06891(.A(new_n7276_), .B(new_n580_), .Y(new_n7277_));
  NOR2  g06892(.A(new_n7277_), .B(new_n586_), .Y(new_n7278_));
  NOR2  g06893(.A(new_n7278_), .B(new_n590_), .Y(new_n7279_));
  NOR2  g06894(.A(new_n7279_), .B(new_n596_), .Y(new_n7280_));
  NOR2  g06895(.A(new_n7280_), .B(new_n600_), .Y(new_n7281_));
  NOR2  g06896(.A(new_n7281_), .B(new_n606_), .Y(new_n7282_));
  NAND2 g06897(.A(new_n608_), .B(\req[68] ), .Y(new_n7283_));
  NOR2  g06898(.A(new_n7283_), .B(new_n7282_), .Y(\grant[68] ));
  INV   g06899(.A(new_n619_), .Y(new_n7285_));
  NOR2  g06900(.A(new_n1017_), .B(new_n7285_), .Y(new_n7286_));
  NOR2  g06901(.A(new_n7286_), .B(new_n626_), .Y(new_n7287_));
  NOR2  g06902(.A(new_n7287_), .B(new_n630_), .Y(new_n7288_));
  NOR2  g06903(.A(new_n7288_), .B(new_n636_), .Y(new_n7289_));
  NOR2  g06904(.A(new_n7289_), .B(new_n640_), .Y(new_n7290_));
  NOR2  g06905(.A(new_n7290_), .B(new_n646_), .Y(new_n7291_));
  NOR2  g06906(.A(new_n7291_), .B(new_n650_), .Y(new_n7292_));
  NOR2  g06907(.A(new_n7292_), .B(new_n656_), .Y(new_n7293_));
  NOR2  g06908(.A(new_n7293_), .B(new_n660_), .Y(new_n7294_));
  NOR2  g06909(.A(new_n7294_), .B(new_n666_), .Y(new_n7295_));
  NOR2  g06910(.A(new_n7295_), .B(new_n670_), .Y(new_n7296_));
  NOR2  g06911(.A(new_n7296_), .B(new_n676_), .Y(new_n7297_));
  NOR2  g06912(.A(new_n7297_), .B(new_n680_), .Y(new_n7298_));
  NOR2  g06913(.A(new_n7298_), .B(new_n686_), .Y(new_n7299_));
  NOR2  g06914(.A(new_n7299_), .B(new_n690_), .Y(new_n7300_));
  NOR2  g06915(.A(new_n7300_), .B(new_n696_), .Y(new_n7301_));
  NOR2  g06916(.A(new_n7301_), .B(new_n700_), .Y(new_n7302_));
  NOR2  g06917(.A(new_n7302_), .B(new_n706_), .Y(new_n7303_));
  NOR2  g06918(.A(new_n7303_), .B(new_n710_), .Y(new_n7304_));
  NOR2  g06919(.A(new_n7304_), .B(new_n716_), .Y(new_n7305_));
  NOR2  g06920(.A(new_n7305_), .B(new_n720_), .Y(new_n7306_));
  NOR2  g06921(.A(new_n7306_), .B(new_n726_), .Y(new_n7307_));
  NOR2  g06922(.A(new_n7307_), .B(new_n730_), .Y(new_n7308_));
  NOR2  g06923(.A(new_n7308_), .B(new_n736_), .Y(new_n7309_));
  NOR2  g06924(.A(new_n7309_), .B(new_n740_), .Y(new_n7310_));
  NOR2  g06925(.A(new_n7310_), .B(new_n746_), .Y(new_n7311_));
  NOR2  g06926(.A(new_n7311_), .B(new_n750_), .Y(new_n7312_));
  NOR2  g06927(.A(new_n7312_), .B(new_n756_), .Y(new_n7313_));
  NOR2  g06928(.A(new_n7313_), .B(new_n760_), .Y(new_n7314_));
  NOR2  g06929(.A(new_n7314_), .B(new_n766_), .Y(new_n7315_));
  NOR2  g06930(.A(new_n7315_), .B(new_n770_), .Y(new_n7316_));
  NOR2  g06931(.A(new_n7316_), .B(new_n776_), .Y(new_n7317_));
  NOR2  g06932(.A(new_n7317_), .B(new_n780_), .Y(new_n7318_));
  NOR2  g06933(.A(new_n7318_), .B(new_n786_), .Y(new_n7319_));
  NOR2  g06934(.A(new_n7319_), .B(new_n790_), .Y(new_n7320_));
  NOR2  g06935(.A(new_n7320_), .B(new_n796_), .Y(new_n7321_));
  NOR2  g06936(.A(new_n7321_), .B(new_n800_), .Y(new_n7322_));
  NOR2  g06937(.A(new_n7322_), .B(new_n806_), .Y(new_n7323_));
  NOR2  g06938(.A(new_n7323_), .B(new_n1616_), .Y(new_n7324_));
  NOR2  g06939(.A(new_n7324_), .B(new_n1618_), .Y(new_n7325_));
  NOR2  g06940(.A(new_n7325_), .B(new_n1885_), .Y(new_n7326_));
  NOR2  g06941(.A(new_n7326_), .B(new_n820_), .Y(new_n7327_));
  NOR2  g06942(.A(new_n7327_), .B(new_n824_), .Y(new_n7328_));
  NOR2  g06943(.A(new_n7328_), .B(new_n829_), .Y(new_n7329_));
  NOR2  g06944(.A(new_n7329_), .B(new_n833_), .Y(new_n7330_));
  NOR2  g06945(.A(new_n7330_), .B(new_n838_), .Y(new_n7331_));
  NOR2  g06946(.A(new_n7331_), .B(new_n842_), .Y(new_n7332_));
  NOR2  g06947(.A(new_n7332_), .B(new_n847_), .Y(new_n7333_));
  NOR2  g06948(.A(new_n7333_), .B(new_n851_), .Y(new_n7334_));
  NOR2  g06949(.A(new_n7334_), .B(new_n856_), .Y(new_n7335_));
  NOR2  g06950(.A(new_n7335_), .B(new_n860_), .Y(new_n7336_));
  NOR2  g06951(.A(new_n7336_), .B(new_n865_), .Y(new_n7337_));
  NOR2  g06952(.A(new_n7337_), .B(new_n869_), .Y(new_n7338_));
  NOR2  g06953(.A(new_n7338_), .B(new_n874_), .Y(new_n7339_));
  NOR2  g06954(.A(new_n7339_), .B(new_n878_), .Y(new_n7340_));
  NOR2  g06955(.A(new_n7340_), .B(new_n883_), .Y(new_n7341_));
  NOR2  g06956(.A(new_n7341_), .B(new_n887_), .Y(new_n7342_));
  NOR2  g06957(.A(new_n7342_), .B(new_n892_), .Y(new_n7343_));
  NOR2  g06958(.A(new_n7343_), .B(new_n896_), .Y(new_n7344_));
  NOR2  g06959(.A(new_n7344_), .B(new_n901_), .Y(new_n7345_));
  NOR2  g06960(.A(new_n7345_), .B(new_n905_), .Y(new_n7346_));
  NOR2  g06961(.A(new_n7346_), .B(new_n910_), .Y(new_n7347_));
  NOR2  g06962(.A(new_n7347_), .B(new_n914_), .Y(new_n7348_));
  NOR2  g06963(.A(new_n7348_), .B(new_n919_), .Y(new_n7349_));
  NOR2  g06964(.A(new_n7349_), .B(new_n923_), .Y(new_n7350_));
  NOR2  g06965(.A(new_n7350_), .B(new_n928_), .Y(new_n7351_));
  NOR2  g06966(.A(new_n7351_), .B(new_n932_), .Y(new_n7352_));
  NOR2  g06967(.A(new_n7352_), .B(new_n937_), .Y(new_n7353_));
  NOR2  g06968(.A(new_n7353_), .B(new_n941_), .Y(new_n7354_));
  NOR2  g06969(.A(new_n7354_), .B(new_n946_), .Y(new_n7355_));
  NOR2  g06970(.A(new_n7355_), .B(new_n950_), .Y(new_n7356_));
  NOR2  g06971(.A(new_n7356_), .B(new_n955_), .Y(new_n7357_));
  NOR2  g06972(.A(new_n7357_), .B(new_n959_), .Y(new_n7358_));
  NOR2  g06973(.A(new_n7358_), .B(new_n964_), .Y(new_n7359_));
  NOR2  g06974(.A(new_n7359_), .B(new_n968_), .Y(new_n7360_));
  NOR2  g06975(.A(new_n7360_), .B(new_n973_), .Y(new_n7361_));
  NOR2  g06976(.A(new_n7361_), .B(new_n977_), .Y(new_n7362_));
  NOR2  g06977(.A(new_n7362_), .B(new_n982_), .Y(new_n7363_));
  NOR2  g06978(.A(new_n7363_), .B(new_n986_), .Y(new_n7364_));
  NOR2  g06979(.A(new_n7364_), .B(new_n991_), .Y(new_n7365_));
  NOR2  g06980(.A(new_n7365_), .B(new_n995_), .Y(new_n7366_));
  NOR2  g06981(.A(new_n7366_), .B(new_n1000_), .Y(new_n7367_));
  NOR2  g06982(.A(new_n7367_), .B(new_n1004_), .Y(new_n7368_));
  NOR2  g06983(.A(new_n7368_), .B(new_n1009_), .Y(new_n7369_));
  NAND2 g06984(.A(new_n1011_), .B(\req[69] ), .Y(new_n7370_));
  NOR2  g06985(.A(new_n7370_), .B(new_n7369_), .Y(\grant[69] ));
  INV   g06986(.A(new_n1021_), .Y(new_n7372_));
  NOR2  g06987(.A(new_n1374_), .B(new_n7372_), .Y(new_n7373_));
  NOR2  g06988(.A(new_n7373_), .B(new_n1027_), .Y(new_n7374_));
  NOR2  g06989(.A(new_n7374_), .B(new_n1031_), .Y(new_n7375_));
  NOR2  g06990(.A(new_n7375_), .B(new_n1036_), .Y(new_n7376_));
  NOR2  g06991(.A(new_n7376_), .B(new_n1040_), .Y(new_n7377_));
  NOR2  g06992(.A(new_n7377_), .B(new_n1045_), .Y(new_n7378_));
  NOR2  g06993(.A(new_n7378_), .B(new_n1049_), .Y(new_n7379_));
  NOR2  g06994(.A(new_n7379_), .B(new_n1054_), .Y(new_n7380_));
  NOR2  g06995(.A(new_n7380_), .B(new_n1058_), .Y(new_n7381_));
  NOR2  g06996(.A(new_n7381_), .B(new_n1063_), .Y(new_n7382_));
  NOR2  g06997(.A(new_n7382_), .B(new_n1067_), .Y(new_n7383_));
  NOR2  g06998(.A(new_n7383_), .B(new_n1072_), .Y(new_n7384_));
  NOR2  g06999(.A(new_n7384_), .B(new_n1076_), .Y(new_n7385_));
  NOR2  g07000(.A(new_n7385_), .B(new_n1081_), .Y(new_n7386_));
  NOR2  g07001(.A(new_n7386_), .B(new_n1085_), .Y(new_n7387_));
  NOR2  g07002(.A(new_n7387_), .B(new_n1090_), .Y(new_n7388_));
  NOR2  g07003(.A(new_n7388_), .B(new_n1094_), .Y(new_n7389_));
  NOR2  g07004(.A(new_n7389_), .B(new_n1099_), .Y(new_n7390_));
  NOR2  g07005(.A(new_n7390_), .B(new_n1103_), .Y(new_n7391_));
  NOR2  g07006(.A(new_n7391_), .B(new_n1108_), .Y(new_n7392_));
  NOR2  g07007(.A(new_n7392_), .B(new_n1112_), .Y(new_n7393_));
  NOR2  g07008(.A(new_n7393_), .B(new_n1117_), .Y(new_n7394_));
  NOR2  g07009(.A(new_n7394_), .B(new_n1121_), .Y(new_n7395_));
  NOR2  g07010(.A(new_n7395_), .B(new_n1126_), .Y(new_n7396_));
  NOR2  g07011(.A(new_n7396_), .B(new_n1130_), .Y(new_n7397_));
  NOR2  g07012(.A(new_n7397_), .B(new_n1135_), .Y(new_n7398_));
  NOR2  g07013(.A(new_n7398_), .B(new_n1139_), .Y(new_n7399_));
  NOR2  g07014(.A(new_n7399_), .B(new_n1144_), .Y(new_n7400_));
  NOR2  g07015(.A(new_n7400_), .B(new_n1148_), .Y(new_n7401_));
  NOR2  g07016(.A(new_n7401_), .B(new_n1153_), .Y(new_n7402_));
  NOR2  g07017(.A(new_n7402_), .B(new_n1157_), .Y(new_n7403_));
  NOR2  g07018(.A(new_n7403_), .B(new_n1162_), .Y(new_n7404_));
  NOR2  g07019(.A(new_n7404_), .B(new_n1166_), .Y(new_n7405_));
  NOR2  g07020(.A(new_n7405_), .B(new_n1171_), .Y(new_n7406_));
  NOR2  g07021(.A(new_n7406_), .B(new_n1175_), .Y(new_n7407_));
  NOR2  g07022(.A(new_n7407_), .B(new_n1180_), .Y(new_n7408_));
  NOR2  g07023(.A(new_n7408_), .B(new_n1184_), .Y(new_n7409_));
  NOR2  g07024(.A(new_n7409_), .B(new_n1189_), .Y(new_n7410_));
  NOR2  g07025(.A(new_n7410_), .B(new_n1707_), .Y(new_n7411_));
  NOR2  g07026(.A(new_n7411_), .B(new_n1709_), .Y(new_n7412_));
  NOR2  g07027(.A(new_n7412_), .B(new_n1973_), .Y(new_n7413_));
  NOR2  g07028(.A(new_n7413_), .B(new_n1199_), .Y(new_n7414_));
  NOR2  g07029(.A(new_n7414_), .B(new_n1203_), .Y(new_n7415_));
  NOR2  g07030(.A(new_n7415_), .B(new_n1207_), .Y(new_n7416_));
  NOR2  g07031(.A(new_n7416_), .B(new_n1211_), .Y(new_n7417_));
  NOR2  g07032(.A(new_n7417_), .B(new_n1215_), .Y(new_n7418_));
  NOR2  g07033(.A(new_n7418_), .B(new_n1219_), .Y(new_n7419_));
  NOR2  g07034(.A(new_n7419_), .B(new_n1223_), .Y(new_n7420_));
  NOR2  g07035(.A(new_n7420_), .B(new_n1227_), .Y(new_n7421_));
  NOR2  g07036(.A(new_n7421_), .B(new_n1231_), .Y(new_n7422_));
  NOR2  g07037(.A(new_n7422_), .B(new_n1235_), .Y(new_n7423_));
  NOR2  g07038(.A(new_n7423_), .B(new_n1239_), .Y(new_n7424_));
  NOR2  g07039(.A(new_n7424_), .B(new_n1243_), .Y(new_n7425_));
  NOR2  g07040(.A(new_n7425_), .B(new_n1247_), .Y(new_n7426_));
  NOR2  g07041(.A(new_n7426_), .B(new_n1251_), .Y(new_n7427_));
  NOR2  g07042(.A(new_n7427_), .B(new_n1255_), .Y(new_n7428_));
  NOR2  g07043(.A(new_n7428_), .B(new_n1259_), .Y(new_n7429_));
  NOR2  g07044(.A(new_n7429_), .B(new_n1263_), .Y(new_n7430_));
  NOR2  g07045(.A(new_n7430_), .B(new_n1267_), .Y(new_n7431_));
  NOR2  g07046(.A(new_n7431_), .B(new_n1271_), .Y(new_n7432_));
  NOR2  g07047(.A(new_n7432_), .B(new_n1275_), .Y(new_n7433_));
  NOR2  g07048(.A(new_n7433_), .B(new_n1279_), .Y(new_n7434_));
  NOR2  g07049(.A(new_n7434_), .B(new_n1283_), .Y(new_n7435_));
  NOR2  g07050(.A(new_n7435_), .B(new_n1287_), .Y(new_n7436_));
  NOR2  g07051(.A(new_n7436_), .B(new_n1291_), .Y(new_n7437_));
  NOR2  g07052(.A(new_n7437_), .B(new_n1295_), .Y(new_n7438_));
  NOR2  g07053(.A(new_n7438_), .B(new_n1299_), .Y(new_n7439_));
  NOR2  g07054(.A(new_n7439_), .B(new_n1303_), .Y(new_n7440_));
  NOR2  g07055(.A(new_n7440_), .B(new_n1307_), .Y(new_n7441_));
  NOR2  g07056(.A(new_n7441_), .B(new_n1311_), .Y(new_n7442_));
  NOR2  g07057(.A(new_n7442_), .B(new_n1315_), .Y(new_n7443_));
  NOR2  g07058(.A(new_n7443_), .B(new_n1319_), .Y(new_n7444_));
  NOR2  g07059(.A(new_n7444_), .B(new_n1323_), .Y(new_n7445_));
  NOR2  g07060(.A(new_n7445_), .B(new_n1327_), .Y(new_n7446_));
  NOR2  g07061(.A(new_n7446_), .B(new_n1331_), .Y(new_n7447_));
  NOR2  g07062(.A(new_n7447_), .B(new_n1335_), .Y(new_n7448_));
  NOR2  g07063(.A(new_n7448_), .B(new_n1339_), .Y(new_n7449_));
  NOR2  g07064(.A(new_n7449_), .B(new_n1343_), .Y(new_n7450_));
  NOR2  g07065(.A(new_n7450_), .B(new_n1347_), .Y(new_n7451_));
  NOR2  g07066(.A(new_n7451_), .B(new_n1351_), .Y(new_n7452_));
  NOR2  g07067(.A(new_n7452_), .B(new_n1355_), .Y(new_n7453_));
  NOR2  g07068(.A(new_n7453_), .B(new_n1359_), .Y(new_n7454_));
  NOR2  g07069(.A(new_n7454_), .B(new_n1363_), .Y(new_n7455_));
  NOR2  g07070(.A(new_n7455_), .B(new_n1367_), .Y(new_n7456_));
  NAND2 g07071(.A(new_n1369_), .B(\req[70] ), .Y(new_n7457_));
  NOR2  g07072(.A(new_n7457_), .B(new_n7456_), .Y(\grant[70] ));
  INV   g07073(.A(new_n1378_), .Y(new_n7459_));
  NOR2  g07074(.A(new_n7459_), .B(new_n625_), .Y(new_n7460_));
  NOR2  g07075(.A(new_n7460_), .B(new_n1383_), .Y(new_n7461_));
  NOR2  g07076(.A(new_n7461_), .B(new_n1387_), .Y(new_n7462_));
  NOR2  g07077(.A(new_n7462_), .B(new_n1391_), .Y(new_n7463_));
  NOR2  g07078(.A(new_n7463_), .B(new_n1395_), .Y(new_n7464_));
  NOR2  g07079(.A(new_n7464_), .B(new_n1399_), .Y(new_n7465_));
  NOR2  g07080(.A(new_n7465_), .B(new_n1403_), .Y(new_n7466_));
  NOR2  g07081(.A(new_n7466_), .B(new_n1407_), .Y(new_n7467_));
  NOR2  g07082(.A(new_n7467_), .B(new_n1411_), .Y(new_n7468_));
  NOR2  g07083(.A(new_n7468_), .B(new_n1415_), .Y(new_n7469_));
  NOR2  g07084(.A(new_n7469_), .B(new_n1419_), .Y(new_n7470_));
  NOR2  g07085(.A(new_n7470_), .B(new_n1423_), .Y(new_n7471_));
  NOR2  g07086(.A(new_n7471_), .B(new_n1427_), .Y(new_n7472_));
  NOR2  g07087(.A(new_n7472_), .B(new_n1431_), .Y(new_n7473_));
  NOR2  g07088(.A(new_n7473_), .B(new_n1435_), .Y(new_n7474_));
  NOR2  g07089(.A(new_n7474_), .B(new_n1439_), .Y(new_n7475_));
  NOR2  g07090(.A(new_n7475_), .B(new_n1443_), .Y(new_n7476_));
  NOR2  g07091(.A(new_n7476_), .B(new_n1447_), .Y(new_n7477_));
  NOR2  g07092(.A(new_n7477_), .B(new_n1451_), .Y(new_n7478_));
  NOR2  g07093(.A(new_n7478_), .B(new_n1455_), .Y(new_n7479_));
  NOR2  g07094(.A(new_n7479_), .B(new_n1459_), .Y(new_n7480_));
  NOR2  g07095(.A(new_n7480_), .B(new_n1463_), .Y(new_n7481_));
  NOR2  g07096(.A(new_n7481_), .B(new_n1467_), .Y(new_n7482_));
  NOR2  g07097(.A(new_n7482_), .B(new_n1471_), .Y(new_n7483_));
  NOR2  g07098(.A(new_n7483_), .B(new_n1475_), .Y(new_n7484_));
  NOR2  g07099(.A(new_n7484_), .B(new_n1479_), .Y(new_n7485_));
  NOR2  g07100(.A(new_n7485_), .B(new_n1483_), .Y(new_n7486_));
  NOR2  g07101(.A(new_n7486_), .B(new_n1487_), .Y(new_n7487_));
  NOR2  g07102(.A(new_n7487_), .B(new_n1491_), .Y(new_n7488_));
  NOR2  g07103(.A(new_n7488_), .B(new_n1495_), .Y(new_n7489_));
  NOR2  g07104(.A(new_n7489_), .B(new_n1499_), .Y(new_n7490_));
  NOR2  g07105(.A(new_n7490_), .B(new_n1503_), .Y(new_n7491_));
  NOR2  g07106(.A(new_n7491_), .B(new_n1507_), .Y(new_n7492_));
  NOR2  g07107(.A(new_n7492_), .B(new_n1511_), .Y(new_n7493_));
  NOR2  g07108(.A(new_n7493_), .B(new_n1515_), .Y(new_n7494_));
  NOR2  g07109(.A(new_n7494_), .B(new_n1519_), .Y(new_n7495_));
  NOR2  g07110(.A(new_n7495_), .B(new_n1523_), .Y(new_n7496_));
  NOR2  g07111(.A(new_n7496_), .B(new_n1527_), .Y(new_n7497_));
  NOR2  g07112(.A(new_n7497_), .B(new_n1797_), .Y(new_n7498_));
  NOR2  g07113(.A(new_n7498_), .B(new_n396_), .Y(new_n7499_));
  NOR2  g07114(.A(new_n7499_), .B(new_n400_), .Y(new_n7500_));
  NOR2  g07115(.A(new_n7500_), .B(new_n406_), .Y(new_n7501_));
  NOR2  g07116(.A(new_n7501_), .B(new_n410_), .Y(new_n7502_));
  NOR2  g07117(.A(new_n7502_), .B(new_n416_), .Y(new_n7503_));
  NOR2  g07118(.A(new_n7503_), .B(new_n420_), .Y(new_n7504_));
  NOR2  g07119(.A(new_n7504_), .B(new_n426_), .Y(new_n7505_));
  NOR2  g07120(.A(new_n7505_), .B(new_n430_), .Y(new_n7506_));
  NOR2  g07121(.A(new_n7506_), .B(new_n436_), .Y(new_n7507_));
  NOR2  g07122(.A(new_n7507_), .B(new_n440_), .Y(new_n7508_));
  NOR2  g07123(.A(new_n7508_), .B(new_n446_), .Y(new_n7509_));
  NOR2  g07124(.A(new_n7509_), .B(new_n450_), .Y(new_n7510_));
  NOR2  g07125(.A(new_n7510_), .B(new_n456_), .Y(new_n7511_));
  NOR2  g07126(.A(new_n7511_), .B(new_n460_), .Y(new_n7512_));
  NOR2  g07127(.A(new_n7512_), .B(new_n466_), .Y(new_n7513_));
  NOR2  g07128(.A(new_n7513_), .B(new_n470_), .Y(new_n7514_));
  NOR2  g07129(.A(new_n7514_), .B(new_n476_), .Y(new_n7515_));
  NOR2  g07130(.A(new_n7515_), .B(new_n480_), .Y(new_n7516_));
  NOR2  g07131(.A(new_n7516_), .B(new_n486_), .Y(new_n7517_));
  NOR2  g07132(.A(new_n7517_), .B(new_n490_), .Y(new_n7518_));
  NOR2  g07133(.A(new_n7518_), .B(new_n496_), .Y(new_n7519_));
  NOR2  g07134(.A(new_n7519_), .B(new_n500_), .Y(new_n7520_));
  NOR2  g07135(.A(new_n7520_), .B(new_n506_), .Y(new_n7521_));
  NOR2  g07136(.A(new_n7521_), .B(new_n510_), .Y(new_n7522_));
  NOR2  g07137(.A(new_n7522_), .B(new_n516_), .Y(new_n7523_));
  NOR2  g07138(.A(new_n7523_), .B(new_n520_), .Y(new_n7524_));
  NOR2  g07139(.A(new_n7524_), .B(new_n526_), .Y(new_n7525_));
  NOR2  g07140(.A(new_n7525_), .B(new_n530_), .Y(new_n7526_));
  NOR2  g07141(.A(new_n7526_), .B(new_n536_), .Y(new_n7527_));
  NOR2  g07142(.A(new_n7527_), .B(new_n540_), .Y(new_n7528_));
  NOR2  g07143(.A(new_n7528_), .B(new_n546_), .Y(new_n7529_));
  NOR2  g07144(.A(new_n7529_), .B(new_n550_), .Y(new_n7530_));
  NOR2  g07145(.A(new_n7530_), .B(new_n556_), .Y(new_n7531_));
  NOR2  g07146(.A(new_n7531_), .B(new_n560_), .Y(new_n7532_));
  NOR2  g07147(.A(new_n7532_), .B(new_n566_), .Y(new_n7533_));
  NOR2  g07148(.A(new_n7533_), .B(new_n570_), .Y(new_n7534_));
  NOR2  g07149(.A(new_n7534_), .B(new_n576_), .Y(new_n7535_));
  NOR2  g07150(.A(new_n7535_), .B(new_n580_), .Y(new_n7536_));
  NOR2  g07151(.A(new_n7536_), .B(new_n586_), .Y(new_n7537_));
  NOR2  g07152(.A(new_n7537_), .B(new_n590_), .Y(new_n7538_));
  NOR2  g07153(.A(new_n7538_), .B(new_n596_), .Y(new_n7539_));
  NOR2  g07154(.A(new_n7539_), .B(new_n600_), .Y(new_n7540_));
  NOR2  g07155(.A(new_n7540_), .B(new_n606_), .Y(new_n7541_));
  NOR2  g07156(.A(new_n7541_), .B(new_n610_), .Y(new_n7542_));
  NOR2  g07157(.A(new_n7542_), .B(new_n616_), .Y(new_n7543_));
  NAND2 g07158(.A(new_n618_), .B(\req[71] ), .Y(new_n7544_));
  NOR2  g07159(.A(new_n7544_), .B(new_n7543_), .Y(\grant[71] ));
  INV   g07160(.A(new_n629_), .Y(new_n7546_));
  NOR2  g07161(.A(new_n1026_), .B(new_n7546_), .Y(new_n7547_));
  NOR2  g07162(.A(new_n7547_), .B(new_n636_), .Y(new_n7548_));
  NOR2  g07163(.A(new_n7548_), .B(new_n640_), .Y(new_n7549_));
  NOR2  g07164(.A(new_n7549_), .B(new_n646_), .Y(new_n7550_));
  NOR2  g07165(.A(new_n7550_), .B(new_n650_), .Y(new_n7551_));
  NOR2  g07166(.A(new_n7551_), .B(new_n656_), .Y(new_n7552_));
  NOR2  g07167(.A(new_n7552_), .B(new_n660_), .Y(new_n7553_));
  NOR2  g07168(.A(new_n7553_), .B(new_n666_), .Y(new_n7554_));
  NOR2  g07169(.A(new_n7554_), .B(new_n670_), .Y(new_n7555_));
  NOR2  g07170(.A(new_n7555_), .B(new_n676_), .Y(new_n7556_));
  NOR2  g07171(.A(new_n7556_), .B(new_n680_), .Y(new_n7557_));
  NOR2  g07172(.A(new_n7557_), .B(new_n686_), .Y(new_n7558_));
  NOR2  g07173(.A(new_n7558_), .B(new_n690_), .Y(new_n7559_));
  NOR2  g07174(.A(new_n7559_), .B(new_n696_), .Y(new_n7560_));
  NOR2  g07175(.A(new_n7560_), .B(new_n700_), .Y(new_n7561_));
  NOR2  g07176(.A(new_n7561_), .B(new_n706_), .Y(new_n7562_));
  NOR2  g07177(.A(new_n7562_), .B(new_n710_), .Y(new_n7563_));
  NOR2  g07178(.A(new_n7563_), .B(new_n716_), .Y(new_n7564_));
  NOR2  g07179(.A(new_n7564_), .B(new_n720_), .Y(new_n7565_));
  NOR2  g07180(.A(new_n7565_), .B(new_n726_), .Y(new_n7566_));
  NOR2  g07181(.A(new_n7566_), .B(new_n730_), .Y(new_n7567_));
  NOR2  g07182(.A(new_n7567_), .B(new_n736_), .Y(new_n7568_));
  NOR2  g07183(.A(new_n7568_), .B(new_n740_), .Y(new_n7569_));
  NOR2  g07184(.A(new_n7569_), .B(new_n746_), .Y(new_n7570_));
  NOR2  g07185(.A(new_n7570_), .B(new_n750_), .Y(new_n7571_));
  NOR2  g07186(.A(new_n7571_), .B(new_n756_), .Y(new_n7572_));
  NOR2  g07187(.A(new_n7572_), .B(new_n760_), .Y(new_n7573_));
  NOR2  g07188(.A(new_n7573_), .B(new_n766_), .Y(new_n7574_));
  NOR2  g07189(.A(new_n7574_), .B(new_n770_), .Y(new_n7575_));
  NOR2  g07190(.A(new_n7575_), .B(new_n776_), .Y(new_n7576_));
  NOR2  g07191(.A(new_n7576_), .B(new_n780_), .Y(new_n7577_));
  NOR2  g07192(.A(new_n7577_), .B(new_n786_), .Y(new_n7578_));
  NOR2  g07193(.A(new_n7578_), .B(new_n790_), .Y(new_n7579_));
  NOR2  g07194(.A(new_n7579_), .B(new_n796_), .Y(new_n7580_));
  NOR2  g07195(.A(new_n7580_), .B(new_n800_), .Y(new_n7581_));
  NOR2  g07196(.A(new_n7581_), .B(new_n806_), .Y(new_n7582_));
  NOR2  g07197(.A(new_n7582_), .B(new_n1616_), .Y(new_n7583_));
  NOR2  g07198(.A(new_n7583_), .B(new_n1618_), .Y(new_n7584_));
  NOR2  g07199(.A(new_n7584_), .B(new_n1885_), .Y(new_n7585_));
  NOR2  g07200(.A(new_n7585_), .B(new_n820_), .Y(new_n7586_));
  NOR2  g07201(.A(new_n7586_), .B(new_n824_), .Y(new_n7587_));
  NOR2  g07202(.A(new_n7587_), .B(new_n829_), .Y(new_n7588_));
  NOR2  g07203(.A(new_n7588_), .B(new_n833_), .Y(new_n7589_));
  NOR2  g07204(.A(new_n7589_), .B(new_n838_), .Y(new_n7590_));
  NOR2  g07205(.A(new_n7590_), .B(new_n842_), .Y(new_n7591_));
  NOR2  g07206(.A(new_n7591_), .B(new_n847_), .Y(new_n7592_));
  NOR2  g07207(.A(new_n7592_), .B(new_n851_), .Y(new_n7593_));
  NOR2  g07208(.A(new_n7593_), .B(new_n856_), .Y(new_n7594_));
  NOR2  g07209(.A(new_n7594_), .B(new_n860_), .Y(new_n7595_));
  NOR2  g07210(.A(new_n7595_), .B(new_n865_), .Y(new_n7596_));
  NOR2  g07211(.A(new_n7596_), .B(new_n869_), .Y(new_n7597_));
  NOR2  g07212(.A(new_n7597_), .B(new_n874_), .Y(new_n7598_));
  NOR2  g07213(.A(new_n7598_), .B(new_n878_), .Y(new_n7599_));
  NOR2  g07214(.A(new_n7599_), .B(new_n883_), .Y(new_n7600_));
  NOR2  g07215(.A(new_n7600_), .B(new_n887_), .Y(new_n7601_));
  NOR2  g07216(.A(new_n7601_), .B(new_n892_), .Y(new_n7602_));
  NOR2  g07217(.A(new_n7602_), .B(new_n896_), .Y(new_n7603_));
  NOR2  g07218(.A(new_n7603_), .B(new_n901_), .Y(new_n7604_));
  NOR2  g07219(.A(new_n7604_), .B(new_n905_), .Y(new_n7605_));
  NOR2  g07220(.A(new_n7605_), .B(new_n910_), .Y(new_n7606_));
  NOR2  g07221(.A(new_n7606_), .B(new_n914_), .Y(new_n7607_));
  NOR2  g07222(.A(new_n7607_), .B(new_n919_), .Y(new_n7608_));
  NOR2  g07223(.A(new_n7608_), .B(new_n923_), .Y(new_n7609_));
  NOR2  g07224(.A(new_n7609_), .B(new_n928_), .Y(new_n7610_));
  NOR2  g07225(.A(new_n7610_), .B(new_n932_), .Y(new_n7611_));
  NOR2  g07226(.A(new_n7611_), .B(new_n937_), .Y(new_n7612_));
  NOR2  g07227(.A(new_n7612_), .B(new_n941_), .Y(new_n7613_));
  NOR2  g07228(.A(new_n7613_), .B(new_n946_), .Y(new_n7614_));
  NOR2  g07229(.A(new_n7614_), .B(new_n950_), .Y(new_n7615_));
  NOR2  g07230(.A(new_n7615_), .B(new_n955_), .Y(new_n7616_));
  NOR2  g07231(.A(new_n7616_), .B(new_n959_), .Y(new_n7617_));
  NOR2  g07232(.A(new_n7617_), .B(new_n964_), .Y(new_n7618_));
  NOR2  g07233(.A(new_n7618_), .B(new_n968_), .Y(new_n7619_));
  NOR2  g07234(.A(new_n7619_), .B(new_n973_), .Y(new_n7620_));
  NOR2  g07235(.A(new_n7620_), .B(new_n977_), .Y(new_n7621_));
  NOR2  g07236(.A(new_n7621_), .B(new_n982_), .Y(new_n7622_));
  NOR2  g07237(.A(new_n7622_), .B(new_n986_), .Y(new_n7623_));
  NOR2  g07238(.A(new_n7623_), .B(new_n991_), .Y(new_n7624_));
  NOR2  g07239(.A(new_n7624_), .B(new_n995_), .Y(new_n7625_));
  NOR2  g07240(.A(new_n7625_), .B(new_n1000_), .Y(new_n7626_));
  NOR2  g07241(.A(new_n7626_), .B(new_n1004_), .Y(new_n7627_));
  NOR2  g07242(.A(new_n7627_), .B(new_n1009_), .Y(new_n7628_));
  NOR2  g07243(.A(new_n7628_), .B(new_n1013_), .Y(new_n7629_));
  NOR2  g07244(.A(new_n7629_), .B(new_n1018_), .Y(new_n7630_));
  NAND2 g07245(.A(new_n1020_), .B(\req[72] ), .Y(new_n7631_));
  NOR2  g07246(.A(new_n7631_), .B(new_n7630_), .Y(\grant[72] ));
  INV   g07247(.A(new_n1030_), .Y(new_n7633_));
  NOR2  g07248(.A(new_n1382_), .B(new_n7633_), .Y(new_n7634_));
  NOR2  g07249(.A(new_n7634_), .B(new_n1036_), .Y(new_n7635_));
  NOR2  g07250(.A(new_n7635_), .B(new_n1040_), .Y(new_n7636_));
  NOR2  g07251(.A(new_n7636_), .B(new_n1045_), .Y(new_n7637_));
  NOR2  g07252(.A(new_n7637_), .B(new_n1049_), .Y(new_n7638_));
  NOR2  g07253(.A(new_n7638_), .B(new_n1054_), .Y(new_n7639_));
  NOR2  g07254(.A(new_n7639_), .B(new_n1058_), .Y(new_n7640_));
  NOR2  g07255(.A(new_n7640_), .B(new_n1063_), .Y(new_n7641_));
  NOR2  g07256(.A(new_n7641_), .B(new_n1067_), .Y(new_n7642_));
  NOR2  g07257(.A(new_n7642_), .B(new_n1072_), .Y(new_n7643_));
  NOR2  g07258(.A(new_n7643_), .B(new_n1076_), .Y(new_n7644_));
  NOR2  g07259(.A(new_n7644_), .B(new_n1081_), .Y(new_n7645_));
  NOR2  g07260(.A(new_n7645_), .B(new_n1085_), .Y(new_n7646_));
  NOR2  g07261(.A(new_n7646_), .B(new_n1090_), .Y(new_n7647_));
  NOR2  g07262(.A(new_n7647_), .B(new_n1094_), .Y(new_n7648_));
  NOR2  g07263(.A(new_n7648_), .B(new_n1099_), .Y(new_n7649_));
  NOR2  g07264(.A(new_n7649_), .B(new_n1103_), .Y(new_n7650_));
  NOR2  g07265(.A(new_n7650_), .B(new_n1108_), .Y(new_n7651_));
  NOR2  g07266(.A(new_n7651_), .B(new_n1112_), .Y(new_n7652_));
  NOR2  g07267(.A(new_n7652_), .B(new_n1117_), .Y(new_n7653_));
  NOR2  g07268(.A(new_n7653_), .B(new_n1121_), .Y(new_n7654_));
  NOR2  g07269(.A(new_n7654_), .B(new_n1126_), .Y(new_n7655_));
  NOR2  g07270(.A(new_n7655_), .B(new_n1130_), .Y(new_n7656_));
  NOR2  g07271(.A(new_n7656_), .B(new_n1135_), .Y(new_n7657_));
  NOR2  g07272(.A(new_n7657_), .B(new_n1139_), .Y(new_n7658_));
  NOR2  g07273(.A(new_n7658_), .B(new_n1144_), .Y(new_n7659_));
  NOR2  g07274(.A(new_n7659_), .B(new_n1148_), .Y(new_n7660_));
  NOR2  g07275(.A(new_n7660_), .B(new_n1153_), .Y(new_n7661_));
  NOR2  g07276(.A(new_n7661_), .B(new_n1157_), .Y(new_n7662_));
  NOR2  g07277(.A(new_n7662_), .B(new_n1162_), .Y(new_n7663_));
  NOR2  g07278(.A(new_n7663_), .B(new_n1166_), .Y(new_n7664_));
  NOR2  g07279(.A(new_n7664_), .B(new_n1171_), .Y(new_n7665_));
  NOR2  g07280(.A(new_n7665_), .B(new_n1175_), .Y(new_n7666_));
  NOR2  g07281(.A(new_n7666_), .B(new_n1180_), .Y(new_n7667_));
  NOR2  g07282(.A(new_n7667_), .B(new_n1184_), .Y(new_n7668_));
  NOR2  g07283(.A(new_n7668_), .B(new_n1189_), .Y(new_n7669_));
  NOR2  g07284(.A(new_n7669_), .B(new_n1707_), .Y(new_n7670_));
  NOR2  g07285(.A(new_n7670_), .B(new_n1709_), .Y(new_n7671_));
  NOR2  g07286(.A(new_n7671_), .B(new_n1973_), .Y(new_n7672_));
  NOR2  g07287(.A(new_n7672_), .B(new_n1199_), .Y(new_n7673_));
  NOR2  g07288(.A(new_n7673_), .B(new_n1203_), .Y(new_n7674_));
  NOR2  g07289(.A(new_n7674_), .B(new_n1207_), .Y(new_n7675_));
  NOR2  g07290(.A(new_n7675_), .B(new_n1211_), .Y(new_n7676_));
  NOR2  g07291(.A(new_n7676_), .B(new_n1215_), .Y(new_n7677_));
  NOR2  g07292(.A(new_n7677_), .B(new_n1219_), .Y(new_n7678_));
  NOR2  g07293(.A(new_n7678_), .B(new_n1223_), .Y(new_n7679_));
  NOR2  g07294(.A(new_n7679_), .B(new_n1227_), .Y(new_n7680_));
  NOR2  g07295(.A(new_n7680_), .B(new_n1231_), .Y(new_n7681_));
  NOR2  g07296(.A(new_n7681_), .B(new_n1235_), .Y(new_n7682_));
  NOR2  g07297(.A(new_n7682_), .B(new_n1239_), .Y(new_n7683_));
  NOR2  g07298(.A(new_n7683_), .B(new_n1243_), .Y(new_n7684_));
  NOR2  g07299(.A(new_n7684_), .B(new_n1247_), .Y(new_n7685_));
  NOR2  g07300(.A(new_n7685_), .B(new_n1251_), .Y(new_n7686_));
  NOR2  g07301(.A(new_n7686_), .B(new_n1255_), .Y(new_n7687_));
  NOR2  g07302(.A(new_n7687_), .B(new_n1259_), .Y(new_n7688_));
  NOR2  g07303(.A(new_n7688_), .B(new_n1263_), .Y(new_n7689_));
  NOR2  g07304(.A(new_n7689_), .B(new_n1267_), .Y(new_n7690_));
  NOR2  g07305(.A(new_n7690_), .B(new_n1271_), .Y(new_n7691_));
  NOR2  g07306(.A(new_n7691_), .B(new_n1275_), .Y(new_n7692_));
  NOR2  g07307(.A(new_n7692_), .B(new_n1279_), .Y(new_n7693_));
  NOR2  g07308(.A(new_n7693_), .B(new_n1283_), .Y(new_n7694_));
  NOR2  g07309(.A(new_n7694_), .B(new_n1287_), .Y(new_n7695_));
  NOR2  g07310(.A(new_n7695_), .B(new_n1291_), .Y(new_n7696_));
  NOR2  g07311(.A(new_n7696_), .B(new_n1295_), .Y(new_n7697_));
  NOR2  g07312(.A(new_n7697_), .B(new_n1299_), .Y(new_n7698_));
  NOR2  g07313(.A(new_n7698_), .B(new_n1303_), .Y(new_n7699_));
  NOR2  g07314(.A(new_n7699_), .B(new_n1307_), .Y(new_n7700_));
  NOR2  g07315(.A(new_n7700_), .B(new_n1311_), .Y(new_n7701_));
  NOR2  g07316(.A(new_n7701_), .B(new_n1315_), .Y(new_n7702_));
  NOR2  g07317(.A(new_n7702_), .B(new_n1319_), .Y(new_n7703_));
  NOR2  g07318(.A(new_n7703_), .B(new_n1323_), .Y(new_n7704_));
  NOR2  g07319(.A(new_n7704_), .B(new_n1327_), .Y(new_n7705_));
  NOR2  g07320(.A(new_n7705_), .B(new_n1331_), .Y(new_n7706_));
  NOR2  g07321(.A(new_n7706_), .B(new_n1335_), .Y(new_n7707_));
  NOR2  g07322(.A(new_n7707_), .B(new_n1339_), .Y(new_n7708_));
  NOR2  g07323(.A(new_n7708_), .B(new_n1343_), .Y(new_n7709_));
  NOR2  g07324(.A(new_n7709_), .B(new_n1347_), .Y(new_n7710_));
  NOR2  g07325(.A(new_n7710_), .B(new_n1351_), .Y(new_n7711_));
  NOR2  g07326(.A(new_n7711_), .B(new_n1355_), .Y(new_n7712_));
  NOR2  g07327(.A(new_n7712_), .B(new_n1359_), .Y(new_n7713_));
  NOR2  g07328(.A(new_n7713_), .B(new_n1363_), .Y(new_n7714_));
  NOR2  g07329(.A(new_n7714_), .B(new_n1367_), .Y(new_n7715_));
  NOR2  g07330(.A(new_n7715_), .B(new_n1371_), .Y(new_n7716_));
  NOR2  g07331(.A(new_n7716_), .B(new_n1375_), .Y(new_n7717_));
  NAND2 g07332(.A(new_n1377_), .B(\req[73] ), .Y(new_n7718_));
  NOR2  g07333(.A(new_n7718_), .B(new_n7717_), .Y(\grant[73] ));
  INV   g07334(.A(new_n1386_), .Y(new_n7720_));
  NOR2  g07335(.A(new_n7720_), .B(new_n635_), .Y(new_n7721_));
  NOR2  g07336(.A(new_n7721_), .B(new_n1391_), .Y(new_n7722_));
  NOR2  g07337(.A(new_n7722_), .B(new_n1395_), .Y(new_n7723_));
  NOR2  g07338(.A(new_n7723_), .B(new_n1399_), .Y(new_n7724_));
  NOR2  g07339(.A(new_n7724_), .B(new_n1403_), .Y(new_n7725_));
  NOR2  g07340(.A(new_n7725_), .B(new_n1407_), .Y(new_n7726_));
  NOR2  g07341(.A(new_n7726_), .B(new_n1411_), .Y(new_n7727_));
  NOR2  g07342(.A(new_n7727_), .B(new_n1415_), .Y(new_n7728_));
  NOR2  g07343(.A(new_n7728_), .B(new_n1419_), .Y(new_n7729_));
  NOR2  g07344(.A(new_n7729_), .B(new_n1423_), .Y(new_n7730_));
  NOR2  g07345(.A(new_n7730_), .B(new_n1427_), .Y(new_n7731_));
  NOR2  g07346(.A(new_n7731_), .B(new_n1431_), .Y(new_n7732_));
  NOR2  g07347(.A(new_n7732_), .B(new_n1435_), .Y(new_n7733_));
  NOR2  g07348(.A(new_n7733_), .B(new_n1439_), .Y(new_n7734_));
  NOR2  g07349(.A(new_n7734_), .B(new_n1443_), .Y(new_n7735_));
  NOR2  g07350(.A(new_n7735_), .B(new_n1447_), .Y(new_n7736_));
  NOR2  g07351(.A(new_n7736_), .B(new_n1451_), .Y(new_n7737_));
  NOR2  g07352(.A(new_n7737_), .B(new_n1455_), .Y(new_n7738_));
  NOR2  g07353(.A(new_n7738_), .B(new_n1459_), .Y(new_n7739_));
  NOR2  g07354(.A(new_n7739_), .B(new_n1463_), .Y(new_n7740_));
  NOR2  g07355(.A(new_n7740_), .B(new_n1467_), .Y(new_n7741_));
  NOR2  g07356(.A(new_n7741_), .B(new_n1471_), .Y(new_n7742_));
  NOR2  g07357(.A(new_n7742_), .B(new_n1475_), .Y(new_n7743_));
  NOR2  g07358(.A(new_n7743_), .B(new_n1479_), .Y(new_n7744_));
  NOR2  g07359(.A(new_n7744_), .B(new_n1483_), .Y(new_n7745_));
  NOR2  g07360(.A(new_n7745_), .B(new_n1487_), .Y(new_n7746_));
  NOR2  g07361(.A(new_n7746_), .B(new_n1491_), .Y(new_n7747_));
  NOR2  g07362(.A(new_n7747_), .B(new_n1495_), .Y(new_n7748_));
  NOR2  g07363(.A(new_n7748_), .B(new_n1499_), .Y(new_n7749_));
  NOR2  g07364(.A(new_n7749_), .B(new_n1503_), .Y(new_n7750_));
  NOR2  g07365(.A(new_n7750_), .B(new_n1507_), .Y(new_n7751_));
  NOR2  g07366(.A(new_n7751_), .B(new_n1511_), .Y(new_n7752_));
  NOR2  g07367(.A(new_n7752_), .B(new_n1515_), .Y(new_n7753_));
  NOR2  g07368(.A(new_n7753_), .B(new_n1519_), .Y(new_n7754_));
  NOR2  g07369(.A(new_n7754_), .B(new_n1523_), .Y(new_n7755_));
  NOR2  g07370(.A(new_n7755_), .B(new_n1527_), .Y(new_n7756_));
  NOR2  g07371(.A(new_n7756_), .B(new_n1797_), .Y(new_n7757_));
  NOR2  g07372(.A(new_n7757_), .B(new_n396_), .Y(new_n7758_));
  NOR2  g07373(.A(new_n7758_), .B(new_n400_), .Y(new_n7759_));
  NOR2  g07374(.A(new_n7759_), .B(new_n406_), .Y(new_n7760_));
  NOR2  g07375(.A(new_n7760_), .B(new_n410_), .Y(new_n7761_));
  NOR2  g07376(.A(new_n7761_), .B(new_n416_), .Y(new_n7762_));
  NOR2  g07377(.A(new_n7762_), .B(new_n420_), .Y(new_n7763_));
  NOR2  g07378(.A(new_n7763_), .B(new_n426_), .Y(new_n7764_));
  NOR2  g07379(.A(new_n7764_), .B(new_n430_), .Y(new_n7765_));
  NOR2  g07380(.A(new_n7765_), .B(new_n436_), .Y(new_n7766_));
  NOR2  g07381(.A(new_n7766_), .B(new_n440_), .Y(new_n7767_));
  NOR2  g07382(.A(new_n7767_), .B(new_n446_), .Y(new_n7768_));
  NOR2  g07383(.A(new_n7768_), .B(new_n450_), .Y(new_n7769_));
  NOR2  g07384(.A(new_n7769_), .B(new_n456_), .Y(new_n7770_));
  NOR2  g07385(.A(new_n7770_), .B(new_n460_), .Y(new_n7771_));
  NOR2  g07386(.A(new_n7771_), .B(new_n466_), .Y(new_n7772_));
  NOR2  g07387(.A(new_n7772_), .B(new_n470_), .Y(new_n7773_));
  NOR2  g07388(.A(new_n7773_), .B(new_n476_), .Y(new_n7774_));
  NOR2  g07389(.A(new_n7774_), .B(new_n480_), .Y(new_n7775_));
  NOR2  g07390(.A(new_n7775_), .B(new_n486_), .Y(new_n7776_));
  NOR2  g07391(.A(new_n7776_), .B(new_n490_), .Y(new_n7777_));
  NOR2  g07392(.A(new_n7777_), .B(new_n496_), .Y(new_n7778_));
  NOR2  g07393(.A(new_n7778_), .B(new_n500_), .Y(new_n7779_));
  NOR2  g07394(.A(new_n7779_), .B(new_n506_), .Y(new_n7780_));
  NOR2  g07395(.A(new_n7780_), .B(new_n510_), .Y(new_n7781_));
  NOR2  g07396(.A(new_n7781_), .B(new_n516_), .Y(new_n7782_));
  NOR2  g07397(.A(new_n7782_), .B(new_n520_), .Y(new_n7783_));
  NOR2  g07398(.A(new_n7783_), .B(new_n526_), .Y(new_n7784_));
  NOR2  g07399(.A(new_n7784_), .B(new_n530_), .Y(new_n7785_));
  NOR2  g07400(.A(new_n7785_), .B(new_n536_), .Y(new_n7786_));
  NOR2  g07401(.A(new_n7786_), .B(new_n540_), .Y(new_n7787_));
  NOR2  g07402(.A(new_n7787_), .B(new_n546_), .Y(new_n7788_));
  NOR2  g07403(.A(new_n7788_), .B(new_n550_), .Y(new_n7789_));
  NOR2  g07404(.A(new_n7789_), .B(new_n556_), .Y(new_n7790_));
  NOR2  g07405(.A(new_n7790_), .B(new_n560_), .Y(new_n7791_));
  NOR2  g07406(.A(new_n7791_), .B(new_n566_), .Y(new_n7792_));
  NOR2  g07407(.A(new_n7792_), .B(new_n570_), .Y(new_n7793_));
  NOR2  g07408(.A(new_n7793_), .B(new_n576_), .Y(new_n7794_));
  NOR2  g07409(.A(new_n7794_), .B(new_n580_), .Y(new_n7795_));
  NOR2  g07410(.A(new_n7795_), .B(new_n586_), .Y(new_n7796_));
  NOR2  g07411(.A(new_n7796_), .B(new_n590_), .Y(new_n7797_));
  NOR2  g07412(.A(new_n7797_), .B(new_n596_), .Y(new_n7798_));
  NOR2  g07413(.A(new_n7798_), .B(new_n600_), .Y(new_n7799_));
  NOR2  g07414(.A(new_n7799_), .B(new_n606_), .Y(new_n7800_));
  NOR2  g07415(.A(new_n7800_), .B(new_n610_), .Y(new_n7801_));
  NOR2  g07416(.A(new_n7801_), .B(new_n616_), .Y(new_n7802_));
  NOR2  g07417(.A(new_n7802_), .B(new_n620_), .Y(new_n7803_));
  NOR2  g07418(.A(new_n7803_), .B(new_n626_), .Y(new_n7804_));
  NAND2 g07419(.A(new_n628_), .B(\req[74] ), .Y(new_n7805_));
  NOR2  g07420(.A(new_n7805_), .B(new_n7804_), .Y(\grant[74] ));
  INV   g07421(.A(new_n639_), .Y(new_n7807_));
  NOR2  g07422(.A(new_n1035_), .B(new_n7807_), .Y(new_n7808_));
  NOR2  g07423(.A(new_n7808_), .B(new_n646_), .Y(new_n7809_));
  NOR2  g07424(.A(new_n7809_), .B(new_n650_), .Y(new_n7810_));
  NOR2  g07425(.A(new_n7810_), .B(new_n656_), .Y(new_n7811_));
  NOR2  g07426(.A(new_n7811_), .B(new_n660_), .Y(new_n7812_));
  NOR2  g07427(.A(new_n7812_), .B(new_n666_), .Y(new_n7813_));
  NOR2  g07428(.A(new_n7813_), .B(new_n670_), .Y(new_n7814_));
  NOR2  g07429(.A(new_n7814_), .B(new_n676_), .Y(new_n7815_));
  NOR2  g07430(.A(new_n7815_), .B(new_n680_), .Y(new_n7816_));
  NOR2  g07431(.A(new_n7816_), .B(new_n686_), .Y(new_n7817_));
  NOR2  g07432(.A(new_n7817_), .B(new_n690_), .Y(new_n7818_));
  NOR2  g07433(.A(new_n7818_), .B(new_n696_), .Y(new_n7819_));
  NOR2  g07434(.A(new_n7819_), .B(new_n700_), .Y(new_n7820_));
  NOR2  g07435(.A(new_n7820_), .B(new_n706_), .Y(new_n7821_));
  NOR2  g07436(.A(new_n7821_), .B(new_n710_), .Y(new_n7822_));
  NOR2  g07437(.A(new_n7822_), .B(new_n716_), .Y(new_n7823_));
  NOR2  g07438(.A(new_n7823_), .B(new_n720_), .Y(new_n7824_));
  NOR2  g07439(.A(new_n7824_), .B(new_n726_), .Y(new_n7825_));
  NOR2  g07440(.A(new_n7825_), .B(new_n730_), .Y(new_n7826_));
  NOR2  g07441(.A(new_n7826_), .B(new_n736_), .Y(new_n7827_));
  NOR2  g07442(.A(new_n7827_), .B(new_n740_), .Y(new_n7828_));
  NOR2  g07443(.A(new_n7828_), .B(new_n746_), .Y(new_n7829_));
  NOR2  g07444(.A(new_n7829_), .B(new_n750_), .Y(new_n7830_));
  NOR2  g07445(.A(new_n7830_), .B(new_n756_), .Y(new_n7831_));
  NOR2  g07446(.A(new_n7831_), .B(new_n760_), .Y(new_n7832_));
  NOR2  g07447(.A(new_n7832_), .B(new_n766_), .Y(new_n7833_));
  NOR2  g07448(.A(new_n7833_), .B(new_n770_), .Y(new_n7834_));
  NOR2  g07449(.A(new_n7834_), .B(new_n776_), .Y(new_n7835_));
  NOR2  g07450(.A(new_n7835_), .B(new_n780_), .Y(new_n7836_));
  NOR2  g07451(.A(new_n7836_), .B(new_n786_), .Y(new_n7837_));
  NOR2  g07452(.A(new_n7837_), .B(new_n790_), .Y(new_n7838_));
  NOR2  g07453(.A(new_n7838_), .B(new_n796_), .Y(new_n7839_));
  NOR2  g07454(.A(new_n7839_), .B(new_n800_), .Y(new_n7840_));
  NOR2  g07455(.A(new_n7840_), .B(new_n806_), .Y(new_n7841_));
  NOR2  g07456(.A(new_n7841_), .B(new_n1616_), .Y(new_n7842_));
  NOR2  g07457(.A(new_n7842_), .B(new_n1618_), .Y(new_n7843_));
  NOR2  g07458(.A(new_n7843_), .B(new_n1885_), .Y(new_n7844_));
  NOR2  g07459(.A(new_n7844_), .B(new_n820_), .Y(new_n7845_));
  NOR2  g07460(.A(new_n7845_), .B(new_n824_), .Y(new_n7846_));
  NOR2  g07461(.A(new_n7846_), .B(new_n829_), .Y(new_n7847_));
  NOR2  g07462(.A(new_n7847_), .B(new_n833_), .Y(new_n7848_));
  NOR2  g07463(.A(new_n7848_), .B(new_n838_), .Y(new_n7849_));
  NOR2  g07464(.A(new_n7849_), .B(new_n842_), .Y(new_n7850_));
  NOR2  g07465(.A(new_n7850_), .B(new_n847_), .Y(new_n7851_));
  NOR2  g07466(.A(new_n7851_), .B(new_n851_), .Y(new_n7852_));
  NOR2  g07467(.A(new_n7852_), .B(new_n856_), .Y(new_n7853_));
  NOR2  g07468(.A(new_n7853_), .B(new_n860_), .Y(new_n7854_));
  NOR2  g07469(.A(new_n7854_), .B(new_n865_), .Y(new_n7855_));
  NOR2  g07470(.A(new_n7855_), .B(new_n869_), .Y(new_n7856_));
  NOR2  g07471(.A(new_n7856_), .B(new_n874_), .Y(new_n7857_));
  NOR2  g07472(.A(new_n7857_), .B(new_n878_), .Y(new_n7858_));
  NOR2  g07473(.A(new_n7858_), .B(new_n883_), .Y(new_n7859_));
  NOR2  g07474(.A(new_n7859_), .B(new_n887_), .Y(new_n7860_));
  NOR2  g07475(.A(new_n7860_), .B(new_n892_), .Y(new_n7861_));
  NOR2  g07476(.A(new_n7861_), .B(new_n896_), .Y(new_n7862_));
  NOR2  g07477(.A(new_n7862_), .B(new_n901_), .Y(new_n7863_));
  NOR2  g07478(.A(new_n7863_), .B(new_n905_), .Y(new_n7864_));
  NOR2  g07479(.A(new_n7864_), .B(new_n910_), .Y(new_n7865_));
  NOR2  g07480(.A(new_n7865_), .B(new_n914_), .Y(new_n7866_));
  NOR2  g07481(.A(new_n7866_), .B(new_n919_), .Y(new_n7867_));
  NOR2  g07482(.A(new_n7867_), .B(new_n923_), .Y(new_n7868_));
  NOR2  g07483(.A(new_n7868_), .B(new_n928_), .Y(new_n7869_));
  NOR2  g07484(.A(new_n7869_), .B(new_n932_), .Y(new_n7870_));
  NOR2  g07485(.A(new_n7870_), .B(new_n937_), .Y(new_n7871_));
  NOR2  g07486(.A(new_n7871_), .B(new_n941_), .Y(new_n7872_));
  NOR2  g07487(.A(new_n7872_), .B(new_n946_), .Y(new_n7873_));
  NOR2  g07488(.A(new_n7873_), .B(new_n950_), .Y(new_n7874_));
  NOR2  g07489(.A(new_n7874_), .B(new_n955_), .Y(new_n7875_));
  NOR2  g07490(.A(new_n7875_), .B(new_n959_), .Y(new_n7876_));
  NOR2  g07491(.A(new_n7876_), .B(new_n964_), .Y(new_n7877_));
  NOR2  g07492(.A(new_n7877_), .B(new_n968_), .Y(new_n7878_));
  NOR2  g07493(.A(new_n7878_), .B(new_n973_), .Y(new_n7879_));
  NOR2  g07494(.A(new_n7879_), .B(new_n977_), .Y(new_n7880_));
  NOR2  g07495(.A(new_n7880_), .B(new_n982_), .Y(new_n7881_));
  NOR2  g07496(.A(new_n7881_), .B(new_n986_), .Y(new_n7882_));
  NOR2  g07497(.A(new_n7882_), .B(new_n991_), .Y(new_n7883_));
  NOR2  g07498(.A(new_n7883_), .B(new_n995_), .Y(new_n7884_));
  NOR2  g07499(.A(new_n7884_), .B(new_n1000_), .Y(new_n7885_));
  NOR2  g07500(.A(new_n7885_), .B(new_n1004_), .Y(new_n7886_));
  NOR2  g07501(.A(new_n7886_), .B(new_n1009_), .Y(new_n7887_));
  NOR2  g07502(.A(new_n7887_), .B(new_n1013_), .Y(new_n7888_));
  NOR2  g07503(.A(new_n7888_), .B(new_n1018_), .Y(new_n7889_));
  NOR2  g07504(.A(new_n7889_), .B(new_n1022_), .Y(new_n7890_));
  NOR2  g07505(.A(new_n7890_), .B(new_n1027_), .Y(new_n7891_));
  NAND2 g07506(.A(new_n1029_), .B(\req[75] ), .Y(new_n7892_));
  NOR2  g07507(.A(new_n7892_), .B(new_n7891_), .Y(\grant[75] ));
  INV   g07508(.A(new_n1039_), .Y(new_n7894_));
  NOR2  g07509(.A(new_n1390_), .B(new_n7894_), .Y(new_n7895_));
  NOR2  g07510(.A(new_n7895_), .B(new_n1045_), .Y(new_n7896_));
  NOR2  g07511(.A(new_n7896_), .B(new_n1049_), .Y(new_n7897_));
  NOR2  g07512(.A(new_n7897_), .B(new_n1054_), .Y(new_n7898_));
  NOR2  g07513(.A(new_n7898_), .B(new_n1058_), .Y(new_n7899_));
  NOR2  g07514(.A(new_n7899_), .B(new_n1063_), .Y(new_n7900_));
  NOR2  g07515(.A(new_n7900_), .B(new_n1067_), .Y(new_n7901_));
  NOR2  g07516(.A(new_n7901_), .B(new_n1072_), .Y(new_n7902_));
  NOR2  g07517(.A(new_n7902_), .B(new_n1076_), .Y(new_n7903_));
  NOR2  g07518(.A(new_n7903_), .B(new_n1081_), .Y(new_n7904_));
  NOR2  g07519(.A(new_n7904_), .B(new_n1085_), .Y(new_n7905_));
  NOR2  g07520(.A(new_n7905_), .B(new_n1090_), .Y(new_n7906_));
  NOR2  g07521(.A(new_n7906_), .B(new_n1094_), .Y(new_n7907_));
  NOR2  g07522(.A(new_n7907_), .B(new_n1099_), .Y(new_n7908_));
  NOR2  g07523(.A(new_n7908_), .B(new_n1103_), .Y(new_n7909_));
  NOR2  g07524(.A(new_n7909_), .B(new_n1108_), .Y(new_n7910_));
  NOR2  g07525(.A(new_n7910_), .B(new_n1112_), .Y(new_n7911_));
  NOR2  g07526(.A(new_n7911_), .B(new_n1117_), .Y(new_n7912_));
  NOR2  g07527(.A(new_n7912_), .B(new_n1121_), .Y(new_n7913_));
  NOR2  g07528(.A(new_n7913_), .B(new_n1126_), .Y(new_n7914_));
  NOR2  g07529(.A(new_n7914_), .B(new_n1130_), .Y(new_n7915_));
  NOR2  g07530(.A(new_n7915_), .B(new_n1135_), .Y(new_n7916_));
  NOR2  g07531(.A(new_n7916_), .B(new_n1139_), .Y(new_n7917_));
  NOR2  g07532(.A(new_n7917_), .B(new_n1144_), .Y(new_n7918_));
  NOR2  g07533(.A(new_n7918_), .B(new_n1148_), .Y(new_n7919_));
  NOR2  g07534(.A(new_n7919_), .B(new_n1153_), .Y(new_n7920_));
  NOR2  g07535(.A(new_n7920_), .B(new_n1157_), .Y(new_n7921_));
  NOR2  g07536(.A(new_n7921_), .B(new_n1162_), .Y(new_n7922_));
  NOR2  g07537(.A(new_n7922_), .B(new_n1166_), .Y(new_n7923_));
  NOR2  g07538(.A(new_n7923_), .B(new_n1171_), .Y(new_n7924_));
  NOR2  g07539(.A(new_n7924_), .B(new_n1175_), .Y(new_n7925_));
  NOR2  g07540(.A(new_n7925_), .B(new_n1180_), .Y(new_n7926_));
  NOR2  g07541(.A(new_n7926_), .B(new_n1184_), .Y(new_n7927_));
  NOR2  g07542(.A(new_n7927_), .B(new_n1189_), .Y(new_n7928_));
  NOR2  g07543(.A(new_n7928_), .B(new_n1707_), .Y(new_n7929_));
  NOR2  g07544(.A(new_n7929_), .B(new_n1709_), .Y(new_n7930_));
  NOR2  g07545(.A(new_n7930_), .B(new_n1973_), .Y(new_n7931_));
  NOR2  g07546(.A(new_n7931_), .B(new_n1199_), .Y(new_n7932_));
  NOR2  g07547(.A(new_n7932_), .B(new_n1203_), .Y(new_n7933_));
  NOR2  g07548(.A(new_n7933_), .B(new_n1207_), .Y(new_n7934_));
  NOR2  g07549(.A(new_n7934_), .B(new_n1211_), .Y(new_n7935_));
  NOR2  g07550(.A(new_n7935_), .B(new_n1215_), .Y(new_n7936_));
  NOR2  g07551(.A(new_n7936_), .B(new_n1219_), .Y(new_n7937_));
  NOR2  g07552(.A(new_n7937_), .B(new_n1223_), .Y(new_n7938_));
  NOR2  g07553(.A(new_n7938_), .B(new_n1227_), .Y(new_n7939_));
  NOR2  g07554(.A(new_n7939_), .B(new_n1231_), .Y(new_n7940_));
  NOR2  g07555(.A(new_n7940_), .B(new_n1235_), .Y(new_n7941_));
  NOR2  g07556(.A(new_n7941_), .B(new_n1239_), .Y(new_n7942_));
  NOR2  g07557(.A(new_n7942_), .B(new_n1243_), .Y(new_n7943_));
  NOR2  g07558(.A(new_n7943_), .B(new_n1247_), .Y(new_n7944_));
  NOR2  g07559(.A(new_n7944_), .B(new_n1251_), .Y(new_n7945_));
  NOR2  g07560(.A(new_n7945_), .B(new_n1255_), .Y(new_n7946_));
  NOR2  g07561(.A(new_n7946_), .B(new_n1259_), .Y(new_n7947_));
  NOR2  g07562(.A(new_n7947_), .B(new_n1263_), .Y(new_n7948_));
  NOR2  g07563(.A(new_n7948_), .B(new_n1267_), .Y(new_n7949_));
  NOR2  g07564(.A(new_n7949_), .B(new_n1271_), .Y(new_n7950_));
  NOR2  g07565(.A(new_n7950_), .B(new_n1275_), .Y(new_n7951_));
  NOR2  g07566(.A(new_n7951_), .B(new_n1279_), .Y(new_n7952_));
  NOR2  g07567(.A(new_n7952_), .B(new_n1283_), .Y(new_n7953_));
  NOR2  g07568(.A(new_n7953_), .B(new_n1287_), .Y(new_n7954_));
  NOR2  g07569(.A(new_n7954_), .B(new_n1291_), .Y(new_n7955_));
  NOR2  g07570(.A(new_n7955_), .B(new_n1295_), .Y(new_n7956_));
  NOR2  g07571(.A(new_n7956_), .B(new_n1299_), .Y(new_n7957_));
  NOR2  g07572(.A(new_n7957_), .B(new_n1303_), .Y(new_n7958_));
  NOR2  g07573(.A(new_n7958_), .B(new_n1307_), .Y(new_n7959_));
  NOR2  g07574(.A(new_n7959_), .B(new_n1311_), .Y(new_n7960_));
  NOR2  g07575(.A(new_n7960_), .B(new_n1315_), .Y(new_n7961_));
  NOR2  g07576(.A(new_n7961_), .B(new_n1319_), .Y(new_n7962_));
  NOR2  g07577(.A(new_n7962_), .B(new_n1323_), .Y(new_n7963_));
  NOR2  g07578(.A(new_n7963_), .B(new_n1327_), .Y(new_n7964_));
  NOR2  g07579(.A(new_n7964_), .B(new_n1331_), .Y(new_n7965_));
  NOR2  g07580(.A(new_n7965_), .B(new_n1335_), .Y(new_n7966_));
  NOR2  g07581(.A(new_n7966_), .B(new_n1339_), .Y(new_n7967_));
  NOR2  g07582(.A(new_n7967_), .B(new_n1343_), .Y(new_n7968_));
  NOR2  g07583(.A(new_n7968_), .B(new_n1347_), .Y(new_n7969_));
  NOR2  g07584(.A(new_n7969_), .B(new_n1351_), .Y(new_n7970_));
  NOR2  g07585(.A(new_n7970_), .B(new_n1355_), .Y(new_n7971_));
  NOR2  g07586(.A(new_n7971_), .B(new_n1359_), .Y(new_n7972_));
  NOR2  g07587(.A(new_n7972_), .B(new_n1363_), .Y(new_n7973_));
  NOR2  g07588(.A(new_n7973_), .B(new_n1367_), .Y(new_n7974_));
  NOR2  g07589(.A(new_n7974_), .B(new_n1371_), .Y(new_n7975_));
  NOR2  g07590(.A(new_n7975_), .B(new_n1375_), .Y(new_n7976_));
  NOR2  g07591(.A(new_n7976_), .B(new_n1379_), .Y(new_n7977_));
  NOR2  g07592(.A(new_n7977_), .B(new_n1383_), .Y(new_n7978_));
  NAND2 g07593(.A(new_n1385_), .B(\req[76] ), .Y(new_n7979_));
  NOR2  g07594(.A(new_n7979_), .B(new_n7978_), .Y(\grant[76] ));
  INV   g07595(.A(new_n1394_), .Y(new_n7981_));
  NOR2  g07596(.A(new_n7981_), .B(new_n645_), .Y(new_n7982_));
  NOR2  g07597(.A(new_n7982_), .B(new_n1399_), .Y(new_n7983_));
  NOR2  g07598(.A(new_n7983_), .B(new_n1403_), .Y(new_n7984_));
  NOR2  g07599(.A(new_n7984_), .B(new_n1407_), .Y(new_n7985_));
  NOR2  g07600(.A(new_n7985_), .B(new_n1411_), .Y(new_n7986_));
  NOR2  g07601(.A(new_n7986_), .B(new_n1415_), .Y(new_n7987_));
  NOR2  g07602(.A(new_n7987_), .B(new_n1419_), .Y(new_n7988_));
  NOR2  g07603(.A(new_n7988_), .B(new_n1423_), .Y(new_n7989_));
  NOR2  g07604(.A(new_n7989_), .B(new_n1427_), .Y(new_n7990_));
  NOR2  g07605(.A(new_n7990_), .B(new_n1431_), .Y(new_n7991_));
  NOR2  g07606(.A(new_n7991_), .B(new_n1435_), .Y(new_n7992_));
  NOR2  g07607(.A(new_n7992_), .B(new_n1439_), .Y(new_n7993_));
  NOR2  g07608(.A(new_n7993_), .B(new_n1443_), .Y(new_n7994_));
  NOR2  g07609(.A(new_n7994_), .B(new_n1447_), .Y(new_n7995_));
  NOR2  g07610(.A(new_n7995_), .B(new_n1451_), .Y(new_n7996_));
  NOR2  g07611(.A(new_n7996_), .B(new_n1455_), .Y(new_n7997_));
  NOR2  g07612(.A(new_n7997_), .B(new_n1459_), .Y(new_n7998_));
  NOR2  g07613(.A(new_n7998_), .B(new_n1463_), .Y(new_n7999_));
  NOR2  g07614(.A(new_n7999_), .B(new_n1467_), .Y(new_n8000_));
  NOR2  g07615(.A(new_n8000_), .B(new_n1471_), .Y(new_n8001_));
  NOR2  g07616(.A(new_n8001_), .B(new_n1475_), .Y(new_n8002_));
  NOR2  g07617(.A(new_n8002_), .B(new_n1479_), .Y(new_n8003_));
  NOR2  g07618(.A(new_n8003_), .B(new_n1483_), .Y(new_n8004_));
  NOR2  g07619(.A(new_n8004_), .B(new_n1487_), .Y(new_n8005_));
  NOR2  g07620(.A(new_n8005_), .B(new_n1491_), .Y(new_n8006_));
  NOR2  g07621(.A(new_n8006_), .B(new_n1495_), .Y(new_n8007_));
  NOR2  g07622(.A(new_n8007_), .B(new_n1499_), .Y(new_n8008_));
  NOR2  g07623(.A(new_n8008_), .B(new_n1503_), .Y(new_n8009_));
  NOR2  g07624(.A(new_n8009_), .B(new_n1507_), .Y(new_n8010_));
  NOR2  g07625(.A(new_n8010_), .B(new_n1511_), .Y(new_n8011_));
  NOR2  g07626(.A(new_n8011_), .B(new_n1515_), .Y(new_n8012_));
  NOR2  g07627(.A(new_n8012_), .B(new_n1519_), .Y(new_n8013_));
  NOR2  g07628(.A(new_n8013_), .B(new_n1523_), .Y(new_n8014_));
  NOR2  g07629(.A(new_n8014_), .B(new_n1527_), .Y(new_n8015_));
  NOR2  g07630(.A(new_n8015_), .B(new_n1797_), .Y(new_n8016_));
  NOR2  g07631(.A(new_n8016_), .B(new_n396_), .Y(new_n8017_));
  NOR2  g07632(.A(new_n8017_), .B(new_n400_), .Y(new_n8018_));
  NOR2  g07633(.A(new_n8018_), .B(new_n406_), .Y(new_n8019_));
  NOR2  g07634(.A(new_n8019_), .B(new_n410_), .Y(new_n8020_));
  NOR2  g07635(.A(new_n8020_), .B(new_n416_), .Y(new_n8021_));
  NOR2  g07636(.A(new_n8021_), .B(new_n420_), .Y(new_n8022_));
  NOR2  g07637(.A(new_n8022_), .B(new_n426_), .Y(new_n8023_));
  NOR2  g07638(.A(new_n8023_), .B(new_n430_), .Y(new_n8024_));
  NOR2  g07639(.A(new_n8024_), .B(new_n436_), .Y(new_n8025_));
  NOR2  g07640(.A(new_n8025_), .B(new_n440_), .Y(new_n8026_));
  NOR2  g07641(.A(new_n8026_), .B(new_n446_), .Y(new_n8027_));
  NOR2  g07642(.A(new_n8027_), .B(new_n450_), .Y(new_n8028_));
  NOR2  g07643(.A(new_n8028_), .B(new_n456_), .Y(new_n8029_));
  NOR2  g07644(.A(new_n8029_), .B(new_n460_), .Y(new_n8030_));
  NOR2  g07645(.A(new_n8030_), .B(new_n466_), .Y(new_n8031_));
  NOR2  g07646(.A(new_n8031_), .B(new_n470_), .Y(new_n8032_));
  NOR2  g07647(.A(new_n8032_), .B(new_n476_), .Y(new_n8033_));
  NOR2  g07648(.A(new_n8033_), .B(new_n480_), .Y(new_n8034_));
  NOR2  g07649(.A(new_n8034_), .B(new_n486_), .Y(new_n8035_));
  NOR2  g07650(.A(new_n8035_), .B(new_n490_), .Y(new_n8036_));
  NOR2  g07651(.A(new_n8036_), .B(new_n496_), .Y(new_n8037_));
  NOR2  g07652(.A(new_n8037_), .B(new_n500_), .Y(new_n8038_));
  NOR2  g07653(.A(new_n8038_), .B(new_n506_), .Y(new_n8039_));
  NOR2  g07654(.A(new_n8039_), .B(new_n510_), .Y(new_n8040_));
  NOR2  g07655(.A(new_n8040_), .B(new_n516_), .Y(new_n8041_));
  NOR2  g07656(.A(new_n8041_), .B(new_n520_), .Y(new_n8042_));
  NOR2  g07657(.A(new_n8042_), .B(new_n526_), .Y(new_n8043_));
  NOR2  g07658(.A(new_n8043_), .B(new_n530_), .Y(new_n8044_));
  NOR2  g07659(.A(new_n8044_), .B(new_n536_), .Y(new_n8045_));
  NOR2  g07660(.A(new_n8045_), .B(new_n540_), .Y(new_n8046_));
  NOR2  g07661(.A(new_n8046_), .B(new_n546_), .Y(new_n8047_));
  NOR2  g07662(.A(new_n8047_), .B(new_n550_), .Y(new_n8048_));
  NOR2  g07663(.A(new_n8048_), .B(new_n556_), .Y(new_n8049_));
  NOR2  g07664(.A(new_n8049_), .B(new_n560_), .Y(new_n8050_));
  NOR2  g07665(.A(new_n8050_), .B(new_n566_), .Y(new_n8051_));
  NOR2  g07666(.A(new_n8051_), .B(new_n570_), .Y(new_n8052_));
  NOR2  g07667(.A(new_n8052_), .B(new_n576_), .Y(new_n8053_));
  NOR2  g07668(.A(new_n8053_), .B(new_n580_), .Y(new_n8054_));
  NOR2  g07669(.A(new_n8054_), .B(new_n586_), .Y(new_n8055_));
  NOR2  g07670(.A(new_n8055_), .B(new_n590_), .Y(new_n8056_));
  NOR2  g07671(.A(new_n8056_), .B(new_n596_), .Y(new_n8057_));
  NOR2  g07672(.A(new_n8057_), .B(new_n600_), .Y(new_n8058_));
  NOR2  g07673(.A(new_n8058_), .B(new_n606_), .Y(new_n8059_));
  NOR2  g07674(.A(new_n8059_), .B(new_n610_), .Y(new_n8060_));
  NOR2  g07675(.A(new_n8060_), .B(new_n616_), .Y(new_n8061_));
  NOR2  g07676(.A(new_n8061_), .B(new_n620_), .Y(new_n8062_));
  NOR2  g07677(.A(new_n8062_), .B(new_n626_), .Y(new_n8063_));
  NOR2  g07678(.A(new_n8063_), .B(new_n630_), .Y(new_n8064_));
  NOR2  g07679(.A(new_n8064_), .B(new_n636_), .Y(new_n8065_));
  NAND2 g07680(.A(new_n638_), .B(\req[77] ), .Y(new_n8066_));
  NOR2  g07681(.A(new_n8066_), .B(new_n8065_), .Y(\grant[77] ));
  INV   g07682(.A(new_n649_), .Y(new_n8068_));
  NOR2  g07683(.A(new_n1044_), .B(new_n8068_), .Y(new_n8069_));
  NOR2  g07684(.A(new_n8069_), .B(new_n656_), .Y(new_n8070_));
  NOR2  g07685(.A(new_n8070_), .B(new_n660_), .Y(new_n8071_));
  NOR2  g07686(.A(new_n8071_), .B(new_n666_), .Y(new_n8072_));
  NOR2  g07687(.A(new_n8072_), .B(new_n670_), .Y(new_n8073_));
  NOR2  g07688(.A(new_n8073_), .B(new_n676_), .Y(new_n8074_));
  NOR2  g07689(.A(new_n8074_), .B(new_n680_), .Y(new_n8075_));
  NOR2  g07690(.A(new_n8075_), .B(new_n686_), .Y(new_n8076_));
  NOR2  g07691(.A(new_n8076_), .B(new_n690_), .Y(new_n8077_));
  NOR2  g07692(.A(new_n8077_), .B(new_n696_), .Y(new_n8078_));
  NOR2  g07693(.A(new_n8078_), .B(new_n700_), .Y(new_n8079_));
  NOR2  g07694(.A(new_n8079_), .B(new_n706_), .Y(new_n8080_));
  NOR2  g07695(.A(new_n8080_), .B(new_n710_), .Y(new_n8081_));
  NOR2  g07696(.A(new_n8081_), .B(new_n716_), .Y(new_n8082_));
  NOR2  g07697(.A(new_n8082_), .B(new_n720_), .Y(new_n8083_));
  NOR2  g07698(.A(new_n8083_), .B(new_n726_), .Y(new_n8084_));
  NOR2  g07699(.A(new_n8084_), .B(new_n730_), .Y(new_n8085_));
  NOR2  g07700(.A(new_n8085_), .B(new_n736_), .Y(new_n8086_));
  NOR2  g07701(.A(new_n8086_), .B(new_n740_), .Y(new_n8087_));
  NOR2  g07702(.A(new_n8087_), .B(new_n746_), .Y(new_n8088_));
  NOR2  g07703(.A(new_n8088_), .B(new_n750_), .Y(new_n8089_));
  NOR2  g07704(.A(new_n8089_), .B(new_n756_), .Y(new_n8090_));
  NOR2  g07705(.A(new_n8090_), .B(new_n760_), .Y(new_n8091_));
  NOR2  g07706(.A(new_n8091_), .B(new_n766_), .Y(new_n8092_));
  NOR2  g07707(.A(new_n8092_), .B(new_n770_), .Y(new_n8093_));
  NOR2  g07708(.A(new_n8093_), .B(new_n776_), .Y(new_n8094_));
  NOR2  g07709(.A(new_n8094_), .B(new_n780_), .Y(new_n8095_));
  NOR2  g07710(.A(new_n8095_), .B(new_n786_), .Y(new_n8096_));
  NOR2  g07711(.A(new_n8096_), .B(new_n790_), .Y(new_n8097_));
  NOR2  g07712(.A(new_n8097_), .B(new_n796_), .Y(new_n8098_));
  NOR2  g07713(.A(new_n8098_), .B(new_n800_), .Y(new_n8099_));
  NOR2  g07714(.A(new_n8099_), .B(new_n806_), .Y(new_n8100_));
  NOR2  g07715(.A(new_n8100_), .B(new_n1616_), .Y(new_n8101_));
  NOR2  g07716(.A(new_n8101_), .B(new_n1618_), .Y(new_n8102_));
  NOR2  g07717(.A(new_n8102_), .B(new_n1885_), .Y(new_n8103_));
  NOR2  g07718(.A(new_n8103_), .B(new_n820_), .Y(new_n8104_));
  NOR2  g07719(.A(new_n8104_), .B(new_n824_), .Y(new_n8105_));
  NOR2  g07720(.A(new_n8105_), .B(new_n829_), .Y(new_n8106_));
  NOR2  g07721(.A(new_n8106_), .B(new_n833_), .Y(new_n8107_));
  NOR2  g07722(.A(new_n8107_), .B(new_n838_), .Y(new_n8108_));
  NOR2  g07723(.A(new_n8108_), .B(new_n842_), .Y(new_n8109_));
  NOR2  g07724(.A(new_n8109_), .B(new_n847_), .Y(new_n8110_));
  NOR2  g07725(.A(new_n8110_), .B(new_n851_), .Y(new_n8111_));
  NOR2  g07726(.A(new_n8111_), .B(new_n856_), .Y(new_n8112_));
  NOR2  g07727(.A(new_n8112_), .B(new_n860_), .Y(new_n8113_));
  NOR2  g07728(.A(new_n8113_), .B(new_n865_), .Y(new_n8114_));
  NOR2  g07729(.A(new_n8114_), .B(new_n869_), .Y(new_n8115_));
  NOR2  g07730(.A(new_n8115_), .B(new_n874_), .Y(new_n8116_));
  NOR2  g07731(.A(new_n8116_), .B(new_n878_), .Y(new_n8117_));
  NOR2  g07732(.A(new_n8117_), .B(new_n883_), .Y(new_n8118_));
  NOR2  g07733(.A(new_n8118_), .B(new_n887_), .Y(new_n8119_));
  NOR2  g07734(.A(new_n8119_), .B(new_n892_), .Y(new_n8120_));
  NOR2  g07735(.A(new_n8120_), .B(new_n896_), .Y(new_n8121_));
  NOR2  g07736(.A(new_n8121_), .B(new_n901_), .Y(new_n8122_));
  NOR2  g07737(.A(new_n8122_), .B(new_n905_), .Y(new_n8123_));
  NOR2  g07738(.A(new_n8123_), .B(new_n910_), .Y(new_n8124_));
  NOR2  g07739(.A(new_n8124_), .B(new_n914_), .Y(new_n8125_));
  NOR2  g07740(.A(new_n8125_), .B(new_n919_), .Y(new_n8126_));
  NOR2  g07741(.A(new_n8126_), .B(new_n923_), .Y(new_n8127_));
  NOR2  g07742(.A(new_n8127_), .B(new_n928_), .Y(new_n8128_));
  NOR2  g07743(.A(new_n8128_), .B(new_n932_), .Y(new_n8129_));
  NOR2  g07744(.A(new_n8129_), .B(new_n937_), .Y(new_n8130_));
  NOR2  g07745(.A(new_n8130_), .B(new_n941_), .Y(new_n8131_));
  NOR2  g07746(.A(new_n8131_), .B(new_n946_), .Y(new_n8132_));
  NOR2  g07747(.A(new_n8132_), .B(new_n950_), .Y(new_n8133_));
  NOR2  g07748(.A(new_n8133_), .B(new_n955_), .Y(new_n8134_));
  NOR2  g07749(.A(new_n8134_), .B(new_n959_), .Y(new_n8135_));
  NOR2  g07750(.A(new_n8135_), .B(new_n964_), .Y(new_n8136_));
  NOR2  g07751(.A(new_n8136_), .B(new_n968_), .Y(new_n8137_));
  NOR2  g07752(.A(new_n8137_), .B(new_n973_), .Y(new_n8138_));
  NOR2  g07753(.A(new_n8138_), .B(new_n977_), .Y(new_n8139_));
  NOR2  g07754(.A(new_n8139_), .B(new_n982_), .Y(new_n8140_));
  NOR2  g07755(.A(new_n8140_), .B(new_n986_), .Y(new_n8141_));
  NOR2  g07756(.A(new_n8141_), .B(new_n991_), .Y(new_n8142_));
  NOR2  g07757(.A(new_n8142_), .B(new_n995_), .Y(new_n8143_));
  NOR2  g07758(.A(new_n8143_), .B(new_n1000_), .Y(new_n8144_));
  NOR2  g07759(.A(new_n8144_), .B(new_n1004_), .Y(new_n8145_));
  NOR2  g07760(.A(new_n8145_), .B(new_n1009_), .Y(new_n8146_));
  NOR2  g07761(.A(new_n8146_), .B(new_n1013_), .Y(new_n8147_));
  NOR2  g07762(.A(new_n8147_), .B(new_n1018_), .Y(new_n8148_));
  NOR2  g07763(.A(new_n8148_), .B(new_n1022_), .Y(new_n8149_));
  NOR2  g07764(.A(new_n8149_), .B(new_n1027_), .Y(new_n8150_));
  NOR2  g07765(.A(new_n8150_), .B(new_n1031_), .Y(new_n8151_));
  NOR2  g07766(.A(new_n8151_), .B(new_n1036_), .Y(new_n8152_));
  NAND2 g07767(.A(new_n1038_), .B(\req[78] ), .Y(new_n8153_));
  NOR2  g07768(.A(new_n8153_), .B(new_n8152_), .Y(\grant[78] ));
  INV   g07769(.A(new_n1048_), .Y(new_n8155_));
  NOR2  g07770(.A(new_n1398_), .B(new_n8155_), .Y(new_n8156_));
  NOR2  g07771(.A(new_n8156_), .B(new_n1054_), .Y(new_n8157_));
  NOR2  g07772(.A(new_n8157_), .B(new_n1058_), .Y(new_n8158_));
  NOR2  g07773(.A(new_n8158_), .B(new_n1063_), .Y(new_n8159_));
  NOR2  g07774(.A(new_n8159_), .B(new_n1067_), .Y(new_n8160_));
  NOR2  g07775(.A(new_n8160_), .B(new_n1072_), .Y(new_n8161_));
  NOR2  g07776(.A(new_n8161_), .B(new_n1076_), .Y(new_n8162_));
  NOR2  g07777(.A(new_n8162_), .B(new_n1081_), .Y(new_n8163_));
  NOR2  g07778(.A(new_n8163_), .B(new_n1085_), .Y(new_n8164_));
  NOR2  g07779(.A(new_n8164_), .B(new_n1090_), .Y(new_n8165_));
  NOR2  g07780(.A(new_n8165_), .B(new_n1094_), .Y(new_n8166_));
  NOR2  g07781(.A(new_n8166_), .B(new_n1099_), .Y(new_n8167_));
  NOR2  g07782(.A(new_n8167_), .B(new_n1103_), .Y(new_n8168_));
  NOR2  g07783(.A(new_n8168_), .B(new_n1108_), .Y(new_n8169_));
  NOR2  g07784(.A(new_n8169_), .B(new_n1112_), .Y(new_n8170_));
  NOR2  g07785(.A(new_n8170_), .B(new_n1117_), .Y(new_n8171_));
  NOR2  g07786(.A(new_n8171_), .B(new_n1121_), .Y(new_n8172_));
  NOR2  g07787(.A(new_n8172_), .B(new_n1126_), .Y(new_n8173_));
  NOR2  g07788(.A(new_n8173_), .B(new_n1130_), .Y(new_n8174_));
  NOR2  g07789(.A(new_n8174_), .B(new_n1135_), .Y(new_n8175_));
  NOR2  g07790(.A(new_n8175_), .B(new_n1139_), .Y(new_n8176_));
  NOR2  g07791(.A(new_n8176_), .B(new_n1144_), .Y(new_n8177_));
  NOR2  g07792(.A(new_n8177_), .B(new_n1148_), .Y(new_n8178_));
  NOR2  g07793(.A(new_n8178_), .B(new_n1153_), .Y(new_n8179_));
  NOR2  g07794(.A(new_n8179_), .B(new_n1157_), .Y(new_n8180_));
  NOR2  g07795(.A(new_n8180_), .B(new_n1162_), .Y(new_n8181_));
  NOR2  g07796(.A(new_n8181_), .B(new_n1166_), .Y(new_n8182_));
  NOR2  g07797(.A(new_n8182_), .B(new_n1171_), .Y(new_n8183_));
  NOR2  g07798(.A(new_n8183_), .B(new_n1175_), .Y(new_n8184_));
  NOR2  g07799(.A(new_n8184_), .B(new_n1180_), .Y(new_n8185_));
  NOR2  g07800(.A(new_n8185_), .B(new_n1184_), .Y(new_n8186_));
  NOR2  g07801(.A(new_n8186_), .B(new_n1189_), .Y(new_n8187_));
  NOR2  g07802(.A(new_n8187_), .B(new_n1707_), .Y(new_n8188_));
  NOR2  g07803(.A(new_n8188_), .B(new_n1709_), .Y(new_n8189_));
  NOR2  g07804(.A(new_n8189_), .B(new_n1973_), .Y(new_n8190_));
  NOR2  g07805(.A(new_n8190_), .B(new_n1199_), .Y(new_n8191_));
  NOR2  g07806(.A(new_n8191_), .B(new_n1203_), .Y(new_n8192_));
  NOR2  g07807(.A(new_n8192_), .B(new_n1207_), .Y(new_n8193_));
  NOR2  g07808(.A(new_n8193_), .B(new_n1211_), .Y(new_n8194_));
  NOR2  g07809(.A(new_n8194_), .B(new_n1215_), .Y(new_n8195_));
  NOR2  g07810(.A(new_n8195_), .B(new_n1219_), .Y(new_n8196_));
  NOR2  g07811(.A(new_n8196_), .B(new_n1223_), .Y(new_n8197_));
  NOR2  g07812(.A(new_n8197_), .B(new_n1227_), .Y(new_n8198_));
  NOR2  g07813(.A(new_n8198_), .B(new_n1231_), .Y(new_n8199_));
  NOR2  g07814(.A(new_n8199_), .B(new_n1235_), .Y(new_n8200_));
  NOR2  g07815(.A(new_n8200_), .B(new_n1239_), .Y(new_n8201_));
  NOR2  g07816(.A(new_n8201_), .B(new_n1243_), .Y(new_n8202_));
  NOR2  g07817(.A(new_n8202_), .B(new_n1247_), .Y(new_n8203_));
  NOR2  g07818(.A(new_n8203_), .B(new_n1251_), .Y(new_n8204_));
  NOR2  g07819(.A(new_n8204_), .B(new_n1255_), .Y(new_n8205_));
  NOR2  g07820(.A(new_n8205_), .B(new_n1259_), .Y(new_n8206_));
  NOR2  g07821(.A(new_n8206_), .B(new_n1263_), .Y(new_n8207_));
  NOR2  g07822(.A(new_n8207_), .B(new_n1267_), .Y(new_n8208_));
  NOR2  g07823(.A(new_n8208_), .B(new_n1271_), .Y(new_n8209_));
  NOR2  g07824(.A(new_n8209_), .B(new_n1275_), .Y(new_n8210_));
  NOR2  g07825(.A(new_n8210_), .B(new_n1279_), .Y(new_n8211_));
  NOR2  g07826(.A(new_n8211_), .B(new_n1283_), .Y(new_n8212_));
  NOR2  g07827(.A(new_n8212_), .B(new_n1287_), .Y(new_n8213_));
  NOR2  g07828(.A(new_n8213_), .B(new_n1291_), .Y(new_n8214_));
  NOR2  g07829(.A(new_n8214_), .B(new_n1295_), .Y(new_n8215_));
  NOR2  g07830(.A(new_n8215_), .B(new_n1299_), .Y(new_n8216_));
  NOR2  g07831(.A(new_n8216_), .B(new_n1303_), .Y(new_n8217_));
  NOR2  g07832(.A(new_n8217_), .B(new_n1307_), .Y(new_n8218_));
  NOR2  g07833(.A(new_n8218_), .B(new_n1311_), .Y(new_n8219_));
  NOR2  g07834(.A(new_n8219_), .B(new_n1315_), .Y(new_n8220_));
  NOR2  g07835(.A(new_n8220_), .B(new_n1319_), .Y(new_n8221_));
  NOR2  g07836(.A(new_n8221_), .B(new_n1323_), .Y(new_n8222_));
  NOR2  g07837(.A(new_n8222_), .B(new_n1327_), .Y(new_n8223_));
  NOR2  g07838(.A(new_n8223_), .B(new_n1331_), .Y(new_n8224_));
  NOR2  g07839(.A(new_n8224_), .B(new_n1335_), .Y(new_n8225_));
  NOR2  g07840(.A(new_n8225_), .B(new_n1339_), .Y(new_n8226_));
  NOR2  g07841(.A(new_n8226_), .B(new_n1343_), .Y(new_n8227_));
  NOR2  g07842(.A(new_n8227_), .B(new_n1347_), .Y(new_n8228_));
  NOR2  g07843(.A(new_n8228_), .B(new_n1351_), .Y(new_n8229_));
  NOR2  g07844(.A(new_n8229_), .B(new_n1355_), .Y(new_n8230_));
  NOR2  g07845(.A(new_n8230_), .B(new_n1359_), .Y(new_n8231_));
  NOR2  g07846(.A(new_n8231_), .B(new_n1363_), .Y(new_n8232_));
  NOR2  g07847(.A(new_n8232_), .B(new_n1367_), .Y(new_n8233_));
  NOR2  g07848(.A(new_n8233_), .B(new_n1371_), .Y(new_n8234_));
  NOR2  g07849(.A(new_n8234_), .B(new_n1375_), .Y(new_n8235_));
  NOR2  g07850(.A(new_n8235_), .B(new_n1379_), .Y(new_n8236_));
  NOR2  g07851(.A(new_n8236_), .B(new_n1383_), .Y(new_n8237_));
  NOR2  g07852(.A(new_n8237_), .B(new_n1387_), .Y(new_n8238_));
  NOR2  g07853(.A(new_n8238_), .B(new_n1391_), .Y(new_n8239_));
  NAND2 g07854(.A(new_n1393_), .B(\req[79] ), .Y(new_n8240_));
  NOR2  g07855(.A(new_n8240_), .B(new_n8239_), .Y(\grant[79] ));
  INV   g07856(.A(new_n1402_), .Y(new_n8242_));
  NOR2  g07857(.A(new_n8242_), .B(new_n655_), .Y(new_n8243_));
  NOR2  g07858(.A(new_n8243_), .B(new_n1407_), .Y(new_n8244_));
  NOR2  g07859(.A(new_n8244_), .B(new_n1411_), .Y(new_n8245_));
  NOR2  g07860(.A(new_n8245_), .B(new_n1415_), .Y(new_n8246_));
  NOR2  g07861(.A(new_n8246_), .B(new_n1419_), .Y(new_n8247_));
  NOR2  g07862(.A(new_n8247_), .B(new_n1423_), .Y(new_n8248_));
  NOR2  g07863(.A(new_n8248_), .B(new_n1427_), .Y(new_n8249_));
  NOR2  g07864(.A(new_n8249_), .B(new_n1431_), .Y(new_n8250_));
  NOR2  g07865(.A(new_n8250_), .B(new_n1435_), .Y(new_n8251_));
  NOR2  g07866(.A(new_n8251_), .B(new_n1439_), .Y(new_n8252_));
  NOR2  g07867(.A(new_n8252_), .B(new_n1443_), .Y(new_n8253_));
  NOR2  g07868(.A(new_n8253_), .B(new_n1447_), .Y(new_n8254_));
  NOR2  g07869(.A(new_n8254_), .B(new_n1451_), .Y(new_n8255_));
  NOR2  g07870(.A(new_n8255_), .B(new_n1455_), .Y(new_n8256_));
  NOR2  g07871(.A(new_n8256_), .B(new_n1459_), .Y(new_n8257_));
  NOR2  g07872(.A(new_n8257_), .B(new_n1463_), .Y(new_n8258_));
  NOR2  g07873(.A(new_n8258_), .B(new_n1467_), .Y(new_n8259_));
  NOR2  g07874(.A(new_n8259_), .B(new_n1471_), .Y(new_n8260_));
  NOR2  g07875(.A(new_n8260_), .B(new_n1475_), .Y(new_n8261_));
  NOR2  g07876(.A(new_n8261_), .B(new_n1479_), .Y(new_n8262_));
  NOR2  g07877(.A(new_n8262_), .B(new_n1483_), .Y(new_n8263_));
  NOR2  g07878(.A(new_n8263_), .B(new_n1487_), .Y(new_n8264_));
  NOR2  g07879(.A(new_n8264_), .B(new_n1491_), .Y(new_n8265_));
  NOR2  g07880(.A(new_n8265_), .B(new_n1495_), .Y(new_n8266_));
  NOR2  g07881(.A(new_n8266_), .B(new_n1499_), .Y(new_n8267_));
  NOR2  g07882(.A(new_n8267_), .B(new_n1503_), .Y(new_n8268_));
  NOR2  g07883(.A(new_n8268_), .B(new_n1507_), .Y(new_n8269_));
  NOR2  g07884(.A(new_n8269_), .B(new_n1511_), .Y(new_n8270_));
  NOR2  g07885(.A(new_n8270_), .B(new_n1515_), .Y(new_n8271_));
  NOR2  g07886(.A(new_n8271_), .B(new_n1519_), .Y(new_n8272_));
  NOR2  g07887(.A(new_n8272_), .B(new_n1523_), .Y(new_n8273_));
  NOR2  g07888(.A(new_n8273_), .B(new_n1527_), .Y(new_n8274_));
  NOR2  g07889(.A(new_n8274_), .B(new_n1797_), .Y(new_n8275_));
  NOR2  g07890(.A(new_n8275_), .B(new_n396_), .Y(new_n8276_));
  NOR2  g07891(.A(new_n8276_), .B(new_n400_), .Y(new_n8277_));
  NOR2  g07892(.A(new_n8277_), .B(new_n406_), .Y(new_n8278_));
  NOR2  g07893(.A(new_n8278_), .B(new_n410_), .Y(new_n8279_));
  NOR2  g07894(.A(new_n8279_), .B(new_n416_), .Y(new_n8280_));
  NOR2  g07895(.A(new_n8280_), .B(new_n420_), .Y(new_n8281_));
  NOR2  g07896(.A(new_n8281_), .B(new_n426_), .Y(new_n8282_));
  NOR2  g07897(.A(new_n8282_), .B(new_n430_), .Y(new_n8283_));
  NOR2  g07898(.A(new_n8283_), .B(new_n436_), .Y(new_n8284_));
  NOR2  g07899(.A(new_n8284_), .B(new_n440_), .Y(new_n8285_));
  NOR2  g07900(.A(new_n8285_), .B(new_n446_), .Y(new_n8286_));
  NOR2  g07901(.A(new_n8286_), .B(new_n450_), .Y(new_n8287_));
  NOR2  g07902(.A(new_n8287_), .B(new_n456_), .Y(new_n8288_));
  NOR2  g07903(.A(new_n8288_), .B(new_n460_), .Y(new_n8289_));
  NOR2  g07904(.A(new_n8289_), .B(new_n466_), .Y(new_n8290_));
  NOR2  g07905(.A(new_n8290_), .B(new_n470_), .Y(new_n8291_));
  NOR2  g07906(.A(new_n8291_), .B(new_n476_), .Y(new_n8292_));
  NOR2  g07907(.A(new_n8292_), .B(new_n480_), .Y(new_n8293_));
  NOR2  g07908(.A(new_n8293_), .B(new_n486_), .Y(new_n8294_));
  NOR2  g07909(.A(new_n8294_), .B(new_n490_), .Y(new_n8295_));
  NOR2  g07910(.A(new_n8295_), .B(new_n496_), .Y(new_n8296_));
  NOR2  g07911(.A(new_n8296_), .B(new_n500_), .Y(new_n8297_));
  NOR2  g07912(.A(new_n8297_), .B(new_n506_), .Y(new_n8298_));
  NOR2  g07913(.A(new_n8298_), .B(new_n510_), .Y(new_n8299_));
  NOR2  g07914(.A(new_n8299_), .B(new_n516_), .Y(new_n8300_));
  NOR2  g07915(.A(new_n8300_), .B(new_n520_), .Y(new_n8301_));
  NOR2  g07916(.A(new_n8301_), .B(new_n526_), .Y(new_n8302_));
  NOR2  g07917(.A(new_n8302_), .B(new_n530_), .Y(new_n8303_));
  NOR2  g07918(.A(new_n8303_), .B(new_n536_), .Y(new_n8304_));
  NOR2  g07919(.A(new_n8304_), .B(new_n540_), .Y(new_n8305_));
  NOR2  g07920(.A(new_n8305_), .B(new_n546_), .Y(new_n8306_));
  NOR2  g07921(.A(new_n8306_), .B(new_n550_), .Y(new_n8307_));
  NOR2  g07922(.A(new_n8307_), .B(new_n556_), .Y(new_n8308_));
  NOR2  g07923(.A(new_n8308_), .B(new_n560_), .Y(new_n8309_));
  NOR2  g07924(.A(new_n8309_), .B(new_n566_), .Y(new_n8310_));
  NOR2  g07925(.A(new_n8310_), .B(new_n570_), .Y(new_n8311_));
  NOR2  g07926(.A(new_n8311_), .B(new_n576_), .Y(new_n8312_));
  NOR2  g07927(.A(new_n8312_), .B(new_n580_), .Y(new_n8313_));
  NOR2  g07928(.A(new_n8313_), .B(new_n586_), .Y(new_n8314_));
  NOR2  g07929(.A(new_n8314_), .B(new_n590_), .Y(new_n8315_));
  NOR2  g07930(.A(new_n8315_), .B(new_n596_), .Y(new_n8316_));
  NOR2  g07931(.A(new_n8316_), .B(new_n600_), .Y(new_n8317_));
  NOR2  g07932(.A(new_n8317_), .B(new_n606_), .Y(new_n8318_));
  NOR2  g07933(.A(new_n8318_), .B(new_n610_), .Y(new_n8319_));
  NOR2  g07934(.A(new_n8319_), .B(new_n616_), .Y(new_n8320_));
  NOR2  g07935(.A(new_n8320_), .B(new_n620_), .Y(new_n8321_));
  NOR2  g07936(.A(new_n8321_), .B(new_n626_), .Y(new_n8322_));
  NOR2  g07937(.A(new_n8322_), .B(new_n630_), .Y(new_n8323_));
  NOR2  g07938(.A(new_n8323_), .B(new_n636_), .Y(new_n8324_));
  NOR2  g07939(.A(new_n8324_), .B(new_n640_), .Y(new_n8325_));
  NOR2  g07940(.A(new_n8325_), .B(new_n646_), .Y(new_n8326_));
  NAND2 g07941(.A(new_n648_), .B(\req[80] ), .Y(new_n8327_));
  NOR2  g07942(.A(new_n8327_), .B(new_n8326_), .Y(\grant[80] ));
  INV   g07943(.A(new_n659_), .Y(new_n8329_));
  NOR2  g07944(.A(new_n1053_), .B(new_n8329_), .Y(new_n8330_));
  NOR2  g07945(.A(new_n8330_), .B(new_n666_), .Y(new_n8331_));
  NOR2  g07946(.A(new_n8331_), .B(new_n670_), .Y(new_n8332_));
  NOR2  g07947(.A(new_n8332_), .B(new_n676_), .Y(new_n8333_));
  NOR2  g07948(.A(new_n8333_), .B(new_n680_), .Y(new_n8334_));
  NOR2  g07949(.A(new_n8334_), .B(new_n686_), .Y(new_n8335_));
  NOR2  g07950(.A(new_n8335_), .B(new_n690_), .Y(new_n8336_));
  NOR2  g07951(.A(new_n8336_), .B(new_n696_), .Y(new_n8337_));
  NOR2  g07952(.A(new_n8337_), .B(new_n700_), .Y(new_n8338_));
  NOR2  g07953(.A(new_n8338_), .B(new_n706_), .Y(new_n8339_));
  NOR2  g07954(.A(new_n8339_), .B(new_n710_), .Y(new_n8340_));
  NOR2  g07955(.A(new_n8340_), .B(new_n716_), .Y(new_n8341_));
  NOR2  g07956(.A(new_n8341_), .B(new_n720_), .Y(new_n8342_));
  NOR2  g07957(.A(new_n8342_), .B(new_n726_), .Y(new_n8343_));
  NOR2  g07958(.A(new_n8343_), .B(new_n730_), .Y(new_n8344_));
  NOR2  g07959(.A(new_n8344_), .B(new_n736_), .Y(new_n8345_));
  NOR2  g07960(.A(new_n8345_), .B(new_n740_), .Y(new_n8346_));
  NOR2  g07961(.A(new_n8346_), .B(new_n746_), .Y(new_n8347_));
  NOR2  g07962(.A(new_n8347_), .B(new_n750_), .Y(new_n8348_));
  NOR2  g07963(.A(new_n8348_), .B(new_n756_), .Y(new_n8349_));
  NOR2  g07964(.A(new_n8349_), .B(new_n760_), .Y(new_n8350_));
  NOR2  g07965(.A(new_n8350_), .B(new_n766_), .Y(new_n8351_));
  NOR2  g07966(.A(new_n8351_), .B(new_n770_), .Y(new_n8352_));
  NOR2  g07967(.A(new_n8352_), .B(new_n776_), .Y(new_n8353_));
  NOR2  g07968(.A(new_n8353_), .B(new_n780_), .Y(new_n8354_));
  NOR2  g07969(.A(new_n8354_), .B(new_n786_), .Y(new_n8355_));
  NOR2  g07970(.A(new_n8355_), .B(new_n790_), .Y(new_n8356_));
  NOR2  g07971(.A(new_n8356_), .B(new_n796_), .Y(new_n8357_));
  NOR2  g07972(.A(new_n8357_), .B(new_n800_), .Y(new_n8358_));
  NOR2  g07973(.A(new_n8358_), .B(new_n806_), .Y(new_n8359_));
  NOR2  g07974(.A(new_n8359_), .B(new_n1616_), .Y(new_n8360_));
  NOR2  g07975(.A(new_n8360_), .B(new_n1618_), .Y(new_n8361_));
  NOR2  g07976(.A(new_n8361_), .B(new_n1885_), .Y(new_n8362_));
  NOR2  g07977(.A(new_n8362_), .B(new_n820_), .Y(new_n8363_));
  NOR2  g07978(.A(new_n8363_), .B(new_n824_), .Y(new_n8364_));
  NOR2  g07979(.A(new_n8364_), .B(new_n829_), .Y(new_n8365_));
  NOR2  g07980(.A(new_n8365_), .B(new_n833_), .Y(new_n8366_));
  NOR2  g07981(.A(new_n8366_), .B(new_n838_), .Y(new_n8367_));
  NOR2  g07982(.A(new_n8367_), .B(new_n842_), .Y(new_n8368_));
  NOR2  g07983(.A(new_n8368_), .B(new_n847_), .Y(new_n8369_));
  NOR2  g07984(.A(new_n8369_), .B(new_n851_), .Y(new_n8370_));
  NOR2  g07985(.A(new_n8370_), .B(new_n856_), .Y(new_n8371_));
  NOR2  g07986(.A(new_n8371_), .B(new_n860_), .Y(new_n8372_));
  NOR2  g07987(.A(new_n8372_), .B(new_n865_), .Y(new_n8373_));
  NOR2  g07988(.A(new_n8373_), .B(new_n869_), .Y(new_n8374_));
  NOR2  g07989(.A(new_n8374_), .B(new_n874_), .Y(new_n8375_));
  NOR2  g07990(.A(new_n8375_), .B(new_n878_), .Y(new_n8376_));
  NOR2  g07991(.A(new_n8376_), .B(new_n883_), .Y(new_n8377_));
  NOR2  g07992(.A(new_n8377_), .B(new_n887_), .Y(new_n8378_));
  NOR2  g07993(.A(new_n8378_), .B(new_n892_), .Y(new_n8379_));
  NOR2  g07994(.A(new_n8379_), .B(new_n896_), .Y(new_n8380_));
  NOR2  g07995(.A(new_n8380_), .B(new_n901_), .Y(new_n8381_));
  NOR2  g07996(.A(new_n8381_), .B(new_n905_), .Y(new_n8382_));
  NOR2  g07997(.A(new_n8382_), .B(new_n910_), .Y(new_n8383_));
  NOR2  g07998(.A(new_n8383_), .B(new_n914_), .Y(new_n8384_));
  NOR2  g07999(.A(new_n8384_), .B(new_n919_), .Y(new_n8385_));
  NOR2  g08000(.A(new_n8385_), .B(new_n923_), .Y(new_n8386_));
  NOR2  g08001(.A(new_n8386_), .B(new_n928_), .Y(new_n8387_));
  NOR2  g08002(.A(new_n8387_), .B(new_n932_), .Y(new_n8388_));
  NOR2  g08003(.A(new_n8388_), .B(new_n937_), .Y(new_n8389_));
  NOR2  g08004(.A(new_n8389_), .B(new_n941_), .Y(new_n8390_));
  NOR2  g08005(.A(new_n8390_), .B(new_n946_), .Y(new_n8391_));
  NOR2  g08006(.A(new_n8391_), .B(new_n950_), .Y(new_n8392_));
  NOR2  g08007(.A(new_n8392_), .B(new_n955_), .Y(new_n8393_));
  NOR2  g08008(.A(new_n8393_), .B(new_n959_), .Y(new_n8394_));
  NOR2  g08009(.A(new_n8394_), .B(new_n964_), .Y(new_n8395_));
  NOR2  g08010(.A(new_n8395_), .B(new_n968_), .Y(new_n8396_));
  NOR2  g08011(.A(new_n8396_), .B(new_n973_), .Y(new_n8397_));
  NOR2  g08012(.A(new_n8397_), .B(new_n977_), .Y(new_n8398_));
  NOR2  g08013(.A(new_n8398_), .B(new_n982_), .Y(new_n8399_));
  NOR2  g08014(.A(new_n8399_), .B(new_n986_), .Y(new_n8400_));
  NOR2  g08015(.A(new_n8400_), .B(new_n991_), .Y(new_n8401_));
  NOR2  g08016(.A(new_n8401_), .B(new_n995_), .Y(new_n8402_));
  NOR2  g08017(.A(new_n8402_), .B(new_n1000_), .Y(new_n8403_));
  NOR2  g08018(.A(new_n8403_), .B(new_n1004_), .Y(new_n8404_));
  NOR2  g08019(.A(new_n8404_), .B(new_n1009_), .Y(new_n8405_));
  NOR2  g08020(.A(new_n8405_), .B(new_n1013_), .Y(new_n8406_));
  NOR2  g08021(.A(new_n8406_), .B(new_n1018_), .Y(new_n8407_));
  NOR2  g08022(.A(new_n8407_), .B(new_n1022_), .Y(new_n8408_));
  NOR2  g08023(.A(new_n8408_), .B(new_n1027_), .Y(new_n8409_));
  NOR2  g08024(.A(new_n8409_), .B(new_n1031_), .Y(new_n8410_));
  NOR2  g08025(.A(new_n8410_), .B(new_n1036_), .Y(new_n8411_));
  NOR2  g08026(.A(new_n8411_), .B(new_n1040_), .Y(new_n8412_));
  NOR2  g08027(.A(new_n8412_), .B(new_n1045_), .Y(new_n8413_));
  NAND2 g08028(.A(new_n1047_), .B(\req[81] ), .Y(new_n8414_));
  NOR2  g08029(.A(new_n8414_), .B(new_n8413_), .Y(\grant[81] ));
  INV   g08030(.A(new_n1057_), .Y(new_n8416_));
  NOR2  g08031(.A(new_n1406_), .B(new_n8416_), .Y(new_n8417_));
  NOR2  g08032(.A(new_n8417_), .B(new_n1063_), .Y(new_n8418_));
  NOR2  g08033(.A(new_n8418_), .B(new_n1067_), .Y(new_n8419_));
  NOR2  g08034(.A(new_n8419_), .B(new_n1072_), .Y(new_n8420_));
  NOR2  g08035(.A(new_n8420_), .B(new_n1076_), .Y(new_n8421_));
  NOR2  g08036(.A(new_n8421_), .B(new_n1081_), .Y(new_n8422_));
  NOR2  g08037(.A(new_n8422_), .B(new_n1085_), .Y(new_n8423_));
  NOR2  g08038(.A(new_n8423_), .B(new_n1090_), .Y(new_n8424_));
  NOR2  g08039(.A(new_n8424_), .B(new_n1094_), .Y(new_n8425_));
  NOR2  g08040(.A(new_n8425_), .B(new_n1099_), .Y(new_n8426_));
  NOR2  g08041(.A(new_n8426_), .B(new_n1103_), .Y(new_n8427_));
  NOR2  g08042(.A(new_n8427_), .B(new_n1108_), .Y(new_n8428_));
  NOR2  g08043(.A(new_n8428_), .B(new_n1112_), .Y(new_n8429_));
  NOR2  g08044(.A(new_n8429_), .B(new_n1117_), .Y(new_n8430_));
  NOR2  g08045(.A(new_n8430_), .B(new_n1121_), .Y(new_n8431_));
  NOR2  g08046(.A(new_n8431_), .B(new_n1126_), .Y(new_n8432_));
  NOR2  g08047(.A(new_n8432_), .B(new_n1130_), .Y(new_n8433_));
  NOR2  g08048(.A(new_n8433_), .B(new_n1135_), .Y(new_n8434_));
  NOR2  g08049(.A(new_n8434_), .B(new_n1139_), .Y(new_n8435_));
  NOR2  g08050(.A(new_n8435_), .B(new_n1144_), .Y(new_n8436_));
  NOR2  g08051(.A(new_n8436_), .B(new_n1148_), .Y(new_n8437_));
  NOR2  g08052(.A(new_n8437_), .B(new_n1153_), .Y(new_n8438_));
  NOR2  g08053(.A(new_n8438_), .B(new_n1157_), .Y(new_n8439_));
  NOR2  g08054(.A(new_n8439_), .B(new_n1162_), .Y(new_n8440_));
  NOR2  g08055(.A(new_n8440_), .B(new_n1166_), .Y(new_n8441_));
  NOR2  g08056(.A(new_n8441_), .B(new_n1171_), .Y(new_n8442_));
  NOR2  g08057(.A(new_n8442_), .B(new_n1175_), .Y(new_n8443_));
  NOR2  g08058(.A(new_n8443_), .B(new_n1180_), .Y(new_n8444_));
  NOR2  g08059(.A(new_n8444_), .B(new_n1184_), .Y(new_n8445_));
  NOR2  g08060(.A(new_n8445_), .B(new_n1189_), .Y(new_n8446_));
  NOR2  g08061(.A(new_n8446_), .B(new_n1707_), .Y(new_n8447_));
  NOR2  g08062(.A(new_n8447_), .B(new_n1709_), .Y(new_n8448_));
  NOR2  g08063(.A(new_n8448_), .B(new_n1973_), .Y(new_n8449_));
  NOR2  g08064(.A(new_n8449_), .B(new_n1199_), .Y(new_n8450_));
  NOR2  g08065(.A(new_n8450_), .B(new_n1203_), .Y(new_n8451_));
  NOR2  g08066(.A(new_n8451_), .B(new_n1207_), .Y(new_n8452_));
  NOR2  g08067(.A(new_n8452_), .B(new_n1211_), .Y(new_n8453_));
  NOR2  g08068(.A(new_n8453_), .B(new_n1215_), .Y(new_n8454_));
  NOR2  g08069(.A(new_n8454_), .B(new_n1219_), .Y(new_n8455_));
  NOR2  g08070(.A(new_n8455_), .B(new_n1223_), .Y(new_n8456_));
  NOR2  g08071(.A(new_n8456_), .B(new_n1227_), .Y(new_n8457_));
  NOR2  g08072(.A(new_n8457_), .B(new_n1231_), .Y(new_n8458_));
  NOR2  g08073(.A(new_n8458_), .B(new_n1235_), .Y(new_n8459_));
  NOR2  g08074(.A(new_n8459_), .B(new_n1239_), .Y(new_n8460_));
  NOR2  g08075(.A(new_n8460_), .B(new_n1243_), .Y(new_n8461_));
  NOR2  g08076(.A(new_n8461_), .B(new_n1247_), .Y(new_n8462_));
  NOR2  g08077(.A(new_n8462_), .B(new_n1251_), .Y(new_n8463_));
  NOR2  g08078(.A(new_n8463_), .B(new_n1255_), .Y(new_n8464_));
  NOR2  g08079(.A(new_n8464_), .B(new_n1259_), .Y(new_n8465_));
  NOR2  g08080(.A(new_n8465_), .B(new_n1263_), .Y(new_n8466_));
  NOR2  g08081(.A(new_n8466_), .B(new_n1267_), .Y(new_n8467_));
  NOR2  g08082(.A(new_n8467_), .B(new_n1271_), .Y(new_n8468_));
  NOR2  g08083(.A(new_n8468_), .B(new_n1275_), .Y(new_n8469_));
  NOR2  g08084(.A(new_n8469_), .B(new_n1279_), .Y(new_n8470_));
  NOR2  g08085(.A(new_n8470_), .B(new_n1283_), .Y(new_n8471_));
  NOR2  g08086(.A(new_n8471_), .B(new_n1287_), .Y(new_n8472_));
  NOR2  g08087(.A(new_n8472_), .B(new_n1291_), .Y(new_n8473_));
  NOR2  g08088(.A(new_n8473_), .B(new_n1295_), .Y(new_n8474_));
  NOR2  g08089(.A(new_n8474_), .B(new_n1299_), .Y(new_n8475_));
  NOR2  g08090(.A(new_n8475_), .B(new_n1303_), .Y(new_n8476_));
  NOR2  g08091(.A(new_n8476_), .B(new_n1307_), .Y(new_n8477_));
  NOR2  g08092(.A(new_n8477_), .B(new_n1311_), .Y(new_n8478_));
  NOR2  g08093(.A(new_n8478_), .B(new_n1315_), .Y(new_n8479_));
  NOR2  g08094(.A(new_n8479_), .B(new_n1319_), .Y(new_n8480_));
  NOR2  g08095(.A(new_n8480_), .B(new_n1323_), .Y(new_n8481_));
  NOR2  g08096(.A(new_n8481_), .B(new_n1327_), .Y(new_n8482_));
  NOR2  g08097(.A(new_n8482_), .B(new_n1331_), .Y(new_n8483_));
  NOR2  g08098(.A(new_n8483_), .B(new_n1335_), .Y(new_n8484_));
  NOR2  g08099(.A(new_n8484_), .B(new_n1339_), .Y(new_n8485_));
  NOR2  g08100(.A(new_n8485_), .B(new_n1343_), .Y(new_n8486_));
  NOR2  g08101(.A(new_n8486_), .B(new_n1347_), .Y(new_n8487_));
  NOR2  g08102(.A(new_n8487_), .B(new_n1351_), .Y(new_n8488_));
  NOR2  g08103(.A(new_n8488_), .B(new_n1355_), .Y(new_n8489_));
  NOR2  g08104(.A(new_n8489_), .B(new_n1359_), .Y(new_n8490_));
  NOR2  g08105(.A(new_n8490_), .B(new_n1363_), .Y(new_n8491_));
  NOR2  g08106(.A(new_n8491_), .B(new_n1367_), .Y(new_n8492_));
  NOR2  g08107(.A(new_n8492_), .B(new_n1371_), .Y(new_n8493_));
  NOR2  g08108(.A(new_n8493_), .B(new_n1375_), .Y(new_n8494_));
  NOR2  g08109(.A(new_n8494_), .B(new_n1379_), .Y(new_n8495_));
  NOR2  g08110(.A(new_n8495_), .B(new_n1383_), .Y(new_n8496_));
  NOR2  g08111(.A(new_n8496_), .B(new_n1387_), .Y(new_n8497_));
  NOR2  g08112(.A(new_n8497_), .B(new_n1391_), .Y(new_n8498_));
  NOR2  g08113(.A(new_n8498_), .B(new_n1395_), .Y(new_n8499_));
  NOR2  g08114(.A(new_n8499_), .B(new_n1399_), .Y(new_n8500_));
  NAND2 g08115(.A(new_n1401_), .B(\req[82] ), .Y(new_n8501_));
  NOR2  g08116(.A(new_n8501_), .B(new_n8500_), .Y(\grant[82] ));
  INV   g08117(.A(new_n1410_), .Y(new_n8503_));
  NOR2  g08118(.A(new_n8503_), .B(new_n665_), .Y(new_n8504_));
  NOR2  g08119(.A(new_n8504_), .B(new_n1415_), .Y(new_n8505_));
  NOR2  g08120(.A(new_n8505_), .B(new_n1419_), .Y(new_n8506_));
  NOR2  g08121(.A(new_n8506_), .B(new_n1423_), .Y(new_n8507_));
  NOR2  g08122(.A(new_n8507_), .B(new_n1427_), .Y(new_n8508_));
  NOR2  g08123(.A(new_n8508_), .B(new_n1431_), .Y(new_n8509_));
  NOR2  g08124(.A(new_n8509_), .B(new_n1435_), .Y(new_n8510_));
  NOR2  g08125(.A(new_n8510_), .B(new_n1439_), .Y(new_n8511_));
  NOR2  g08126(.A(new_n8511_), .B(new_n1443_), .Y(new_n8512_));
  NOR2  g08127(.A(new_n8512_), .B(new_n1447_), .Y(new_n8513_));
  NOR2  g08128(.A(new_n8513_), .B(new_n1451_), .Y(new_n8514_));
  NOR2  g08129(.A(new_n8514_), .B(new_n1455_), .Y(new_n8515_));
  NOR2  g08130(.A(new_n8515_), .B(new_n1459_), .Y(new_n8516_));
  NOR2  g08131(.A(new_n8516_), .B(new_n1463_), .Y(new_n8517_));
  NOR2  g08132(.A(new_n8517_), .B(new_n1467_), .Y(new_n8518_));
  NOR2  g08133(.A(new_n8518_), .B(new_n1471_), .Y(new_n8519_));
  NOR2  g08134(.A(new_n8519_), .B(new_n1475_), .Y(new_n8520_));
  NOR2  g08135(.A(new_n8520_), .B(new_n1479_), .Y(new_n8521_));
  NOR2  g08136(.A(new_n8521_), .B(new_n1483_), .Y(new_n8522_));
  NOR2  g08137(.A(new_n8522_), .B(new_n1487_), .Y(new_n8523_));
  NOR2  g08138(.A(new_n8523_), .B(new_n1491_), .Y(new_n8524_));
  NOR2  g08139(.A(new_n8524_), .B(new_n1495_), .Y(new_n8525_));
  NOR2  g08140(.A(new_n8525_), .B(new_n1499_), .Y(new_n8526_));
  NOR2  g08141(.A(new_n8526_), .B(new_n1503_), .Y(new_n8527_));
  NOR2  g08142(.A(new_n8527_), .B(new_n1507_), .Y(new_n8528_));
  NOR2  g08143(.A(new_n8528_), .B(new_n1511_), .Y(new_n8529_));
  NOR2  g08144(.A(new_n8529_), .B(new_n1515_), .Y(new_n8530_));
  NOR2  g08145(.A(new_n8530_), .B(new_n1519_), .Y(new_n8531_));
  NOR2  g08146(.A(new_n8531_), .B(new_n1523_), .Y(new_n8532_));
  NOR2  g08147(.A(new_n8532_), .B(new_n1527_), .Y(new_n8533_));
  NOR2  g08148(.A(new_n8533_), .B(new_n1797_), .Y(new_n8534_));
  NOR2  g08149(.A(new_n8534_), .B(new_n396_), .Y(new_n8535_));
  NOR2  g08150(.A(new_n8535_), .B(new_n400_), .Y(new_n8536_));
  NOR2  g08151(.A(new_n8536_), .B(new_n406_), .Y(new_n8537_));
  NOR2  g08152(.A(new_n8537_), .B(new_n410_), .Y(new_n8538_));
  NOR2  g08153(.A(new_n8538_), .B(new_n416_), .Y(new_n8539_));
  NOR2  g08154(.A(new_n8539_), .B(new_n420_), .Y(new_n8540_));
  NOR2  g08155(.A(new_n8540_), .B(new_n426_), .Y(new_n8541_));
  NOR2  g08156(.A(new_n8541_), .B(new_n430_), .Y(new_n8542_));
  NOR2  g08157(.A(new_n8542_), .B(new_n436_), .Y(new_n8543_));
  NOR2  g08158(.A(new_n8543_), .B(new_n440_), .Y(new_n8544_));
  NOR2  g08159(.A(new_n8544_), .B(new_n446_), .Y(new_n8545_));
  NOR2  g08160(.A(new_n8545_), .B(new_n450_), .Y(new_n8546_));
  NOR2  g08161(.A(new_n8546_), .B(new_n456_), .Y(new_n8547_));
  NOR2  g08162(.A(new_n8547_), .B(new_n460_), .Y(new_n8548_));
  NOR2  g08163(.A(new_n8548_), .B(new_n466_), .Y(new_n8549_));
  NOR2  g08164(.A(new_n8549_), .B(new_n470_), .Y(new_n8550_));
  NOR2  g08165(.A(new_n8550_), .B(new_n476_), .Y(new_n8551_));
  NOR2  g08166(.A(new_n8551_), .B(new_n480_), .Y(new_n8552_));
  NOR2  g08167(.A(new_n8552_), .B(new_n486_), .Y(new_n8553_));
  NOR2  g08168(.A(new_n8553_), .B(new_n490_), .Y(new_n8554_));
  NOR2  g08169(.A(new_n8554_), .B(new_n496_), .Y(new_n8555_));
  NOR2  g08170(.A(new_n8555_), .B(new_n500_), .Y(new_n8556_));
  NOR2  g08171(.A(new_n8556_), .B(new_n506_), .Y(new_n8557_));
  NOR2  g08172(.A(new_n8557_), .B(new_n510_), .Y(new_n8558_));
  NOR2  g08173(.A(new_n8558_), .B(new_n516_), .Y(new_n8559_));
  NOR2  g08174(.A(new_n8559_), .B(new_n520_), .Y(new_n8560_));
  NOR2  g08175(.A(new_n8560_), .B(new_n526_), .Y(new_n8561_));
  NOR2  g08176(.A(new_n8561_), .B(new_n530_), .Y(new_n8562_));
  NOR2  g08177(.A(new_n8562_), .B(new_n536_), .Y(new_n8563_));
  NOR2  g08178(.A(new_n8563_), .B(new_n540_), .Y(new_n8564_));
  NOR2  g08179(.A(new_n8564_), .B(new_n546_), .Y(new_n8565_));
  NOR2  g08180(.A(new_n8565_), .B(new_n550_), .Y(new_n8566_));
  NOR2  g08181(.A(new_n8566_), .B(new_n556_), .Y(new_n8567_));
  NOR2  g08182(.A(new_n8567_), .B(new_n560_), .Y(new_n8568_));
  NOR2  g08183(.A(new_n8568_), .B(new_n566_), .Y(new_n8569_));
  NOR2  g08184(.A(new_n8569_), .B(new_n570_), .Y(new_n8570_));
  NOR2  g08185(.A(new_n8570_), .B(new_n576_), .Y(new_n8571_));
  NOR2  g08186(.A(new_n8571_), .B(new_n580_), .Y(new_n8572_));
  NOR2  g08187(.A(new_n8572_), .B(new_n586_), .Y(new_n8573_));
  NOR2  g08188(.A(new_n8573_), .B(new_n590_), .Y(new_n8574_));
  NOR2  g08189(.A(new_n8574_), .B(new_n596_), .Y(new_n8575_));
  NOR2  g08190(.A(new_n8575_), .B(new_n600_), .Y(new_n8576_));
  NOR2  g08191(.A(new_n8576_), .B(new_n606_), .Y(new_n8577_));
  NOR2  g08192(.A(new_n8577_), .B(new_n610_), .Y(new_n8578_));
  NOR2  g08193(.A(new_n8578_), .B(new_n616_), .Y(new_n8579_));
  NOR2  g08194(.A(new_n8579_), .B(new_n620_), .Y(new_n8580_));
  NOR2  g08195(.A(new_n8580_), .B(new_n626_), .Y(new_n8581_));
  NOR2  g08196(.A(new_n8581_), .B(new_n630_), .Y(new_n8582_));
  NOR2  g08197(.A(new_n8582_), .B(new_n636_), .Y(new_n8583_));
  NOR2  g08198(.A(new_n8583_), .B(new_n640_), .Y(new_n8584_));
  NOR2  g08199(.A(new_n8584_), .B(new_n646_), .Y(new_n8585_));
  NOR2  g08200(.A(new_n8585_), .B(new_n650_), .Y(new_n8586_));
  NOR2  g08201(.A(new_n8586_), .B(new_n656_), .Y(new_n8587_));
  NAND2 g08202(.A(new_n658_), .B(\req[83] ), .Y(new_n8588_));
  NOR2  g08203(.A(new_n8588_), .B(new_n8587_), .Y(\grant[83] ));
  INV   g08204(.A(new_n669_), .Y(new_n8590_));
  NOR2  g08205(.A(new_n1062_), .B(new_n8590_), .Y(new_n8591_));
  NOR2  g08206(.A(new_n8591_), .B(new_n676_), .Y(new_n8592_));
  NOR2  g08207(.A(new_n8592_), .B(new_n680_), .Y(new_n8593_));
  NOR2  g08208(.A(new_n8593_), .B(new_n686_), .Y(new_n8594_));
  NOR2  g08209(.A(new_n8594_), .B(new_n690_), .Y(new_n8595_));
  NOR2  g08210(.A(new_n8595_), .B(new_n696_), .Y(new_n8596_));
  NOR2  g08211(.A(new_n8596_), .B(new_n700_), .Y(new_n8597_));
  NOR2  g08212(.A(new_n8597_), .B(new_n706_), .Y(new_n8598_));
  NOR2  g08213(.A(new_n8598_), .B(new_n710_), .Y(new_n8599_));
  NOR2  g08214(.A(new_n8599_), .B(new_n716_), .Y(new_n8600_));
  NOR2  g08215(.A(new_n8600_), .B(new_n720_), .Y(new_n8601_));
  NOR2  g08216(.A(new_n8601_), .B(new_n726_), .Y(new_n8602_));
  NOR2  g08217(.A(new_n8602_), .B(new_n730_), .Y(new_n8603_));
  NOR2  g08218(.A(new_n8603_), .B(new_n736_), .Y(new_n8604_));
  NOR2  g08219(.A(new_n8604_), .B(new_n740_), .Y(new_n8605_));
  NOR2  g08220(.A(new_n8605_), .B(new_n746_), .Y(new_n8606_));
  NOR2  g08221(.A(new_n8606_), .B(new_n750_), .Y(new_n8607_));
  NOR2  g08222(.A(new_n8607_), .B(new_n756_), .Y(new_n8608_));
  NOR2  g08223(.A(new_n8608_), .B(new_n760_), .Y(new_n8609_));
  NOR2  g08224(.A(new_n8609_), .B(new_n766_), .Y(new_n8610_));
  NOR2  g08225(.A(new_n8610_), .B(new_n770_), .Y(new_n8611_));
  NOR2  g08226(.A(new_n8611_), .B(new_n776_), .Y(new_n8612_));
  NOR2  g08227(.A(new_n8612_), .B(new_n780_), .Y(new_n8613_));
  NOR2  g08228(.A(new_n8613_), .B(new_n786_), .Y(new_n8614_));
  NOR2  g08229(.A(new_n8614_), .B(new_n790_), .Y(new_n8615_));
  NOR2  g08230(.A(new_n8615_), .B(new_n796_), .Y(new_n8616_));
  NOR2  g08231(.A(new_n8616_), .B(new_n800_), .Y(new_n8617_));
  NOR2  g08232(.A(new_n8617_), .B(new_n806_), .Y(new_n8618_));
  NOR2  g08233(.A(new_n8618_), .B(new_n1616_), .Y(new_n8619_));
  NOR2  g08234(.A(new_n8619_), .B(new_n1618_), .Y(new_n8620_));
  NOR2  g08235(.A(new_n8620_), .B(new_n1885_), .Y(new_n8621_));
  NOR2  g08236(.A(new_n8621_), .B(new_n820_), .Y(new_n8622_));
  NOR2  g08237(.A(new_n8622_), .B(new_n824_), .Y(new_n8623_));
  NOR2  g08238(.A(new_n8623_), .B(new_n829_), .Y(new_n8624_));
  NOR2  g08239(.A(new_n8624_), .B(new_n833_), .Y(new_n8625_));
  NOR2  g08240(.A(new_n8625_), .B(new_n838_), .Y(new_n8626_));
  NOR2  g08241(.A(new_n8626_), .B(new_n842_), .Y(new_n8627_));
  NOR2  g08242(.A(new_n8627_), .B(new_n847_), .Y(new_n8628_));
  NOR2  g08243(.A(new_n8628_), .B(new_n851_), .Y(new_n8629_));
  NOR2  g08244(.A(new_n8629_), .B(new_n856_), .Y(new_n8630_));
  NOR2  g08245(.A(new_n8630_), .B(new_n860_), .Y(new_n8631_));
  NOR2  g08246(.A(new_n8631_), .B(new_n865_), .Y(new_n8632_));
  NOR2  g08247(.A(new_n8632_), .B(new_n869_), .Y(new_n8633_));
  NOR2  g08248(.A(new_n8633_), .B(new_n874_), .Y(new_n8634_));
  NOR2  g08249(.A(new_n8634_), .B(new_n878_), .Y(new_n8635_));
  NOR2  g08250(.A(new_n8635_), .B(new_n883_), .Y(new_n8636_));
  NOR2  g08251(.A(new_n8636_), .B(new_n887_), .Y(new_n8637_));
  NOR2  g08252(.A(new_n8637_), .B(new_n892_), .Y(new_n8638_));
  NOR2  g08253(.A(new_n8638_), .B(new_n896_), .Y(new_n8639_));
  NOR2  g08254(.A(new_n8639_), .B(new_n901_), .Y(new_n8640_));
  NOR2  g08255(.A(new_n8640_), .B(new_n905_), .Y(new_n8641_));
  NOR2  g08256(.A(new_n8641_), .B(new_n910_), .Y(new_n8642_));
  NOR2  g08257(.A(new_n8642_), .B(new_n914_), .Y(new_n8643_));
  NOR2  g08258(.A(new_n8643_), .B(new_n919_), .Y(new_n8644_));
  NOR2  g08259(.A(new_n8644_), .B(new_n923_), .Y(new_n8645_));
  NOR2  g08260(.A(new_n8645_), .B(new_n928_), .Y(new_n8646_));
  NOR2  g08261(.A(new_n8646_), .B(new_n932_), .Y(new_n8647_));
  NOR2  g08262(.A(new_n8647_), .B(new_n937_), .Y(new_n8648_));
  NOR2  g08263(.A(new_n8648_), .B(new_n941_), .Y(new_n8649_));
  NOR2  g08264(.A(new_n8649_), .B(new_n946_), .Y(new_n8650_));
  NOR2  g08265(.A(new_n8650_), .B(new_n950_), .Y(new_n8651_));
  NOR2  g08266(.A(new_n8651_), .B(new_n955_), .Y(new_n8652_));
  NOR2  g08267(.A(new_n8652_), .B(new_n959_), .Y(new_n8653_));
  NOR2  g08268(.A(new_n8653_), .B(new_n964_), .Y(new_n8654_));
  NOR2  g08269(.A(new_n8654_), .B(new_n968_), .Y(new_n8655_));
  NOR2  g08270(.A(new_n8655_), .B(new_n973_), .Y(new_n8656_));
  NOR2  g08271(.A(new_n8656_), .B(new_n977_), .Y(new_n8657_));
  NOR2  g08272(.A(new_n8657_), .B(new_n982_), .Y(new_n8658_));
  NOR2  g08273(.A(new_n8658_), .B(new_n986_), .Y(new_n8659_));
  NOR2  g08274(.A(new_n8659_), .B(new_n991_), .Y(new_n8660_));
  NOR2  g08275(.A(new_n8660_), .B(new_n995_), .Y(new_n8661_));
  NOR2  g08276(.A(new_n8661_), .B(new_n1000_), .Y(new_n8662_));
  NOR2  g08277(.A(new_n8662_), .B(new_n1004_), .Y(new_n8663_));
  NOR2  g08278(.A(new_n8663_), .B(new_n1009_), .Y(new_n8664_));
  NOR2  g08279(.A(new_n8664_), .B(new_n1013_), .Y(new_n8665_));
  NOR2  g08280(.A(new_n8665_), .B(new_n1018_), .Y(new_n8666_));
  NOR2  g08281(.A(new_n8666_), .B(new_n1022_), .Y(new_n8667_));
  NOR2  g08282(.A(new_n8667_), .B(new_n1027_), .Y(new_n8668_));
  NOR2  g08283(.A(new_n8668_), .B(new_n1031_), .Y(new_n8669_));
  NOR2  g08284(.A(new_n8669_), .B(new_n1036_), .Y(new_n8670_));
  NOR2  g08285(.A(new_n8670_), .B(new_n1040_), .Y(new_n8671_));
  NOR2  g08286(.A(new_n8671_), .B(new_n1045_), .Y(new_n8672_));
  NOR2  g08287(.A(new_n8672_), .B(new_n1049_), .Y(new_n8673_));
  NOR2  g08288(.A(new_n8673_), .B(new_n1054_), .Y(new_n8674_));
  NAND2 g08289(.A(new_n1056_), .B(\req[84] ), .Y(new_n8675_));
  NOR2  g08290(.A(new_n8675_), .B(new_n8674_), .Y(\grant[84] ));
  INV   g08291(.A(new_n1066_), .Y(new_n8677_));
  NOR2  g08292(.A(new_n1414_), .B(new_n8677_), .Y(new_n8678_));
  NOR2  g08293(.A(new_n8678_), .B(new_n1072_), .Y(new_n8679_));
  NOR2  g08294(.A(new_n8679_), .B(new_n1076_), .Y(new_n8680_));
  NOR2  g08295(.A(new_n8680_), .B(new_n1081_), .Y(new_n8681_));
  NOR2  g08296(.A(new_n8681_), .B(new_n1085_), .Y(new_n8682_));
  NOR2  g08297(.A(new_n8682_), .B(new_n1090_), .Y(new_n8683_));
  NOR2  g08298(.A(new_n8683_), .B(new_n1094_), .Y(new_n8684_));
  NOR2  g08299(.A(new_n8684_), .B(new_n1099_), .Y(new_n8685_));
  NOR2  g08300(.A(new_n8685_), .B(new_n1103_), .Y(new_n8686_));
  NOR2  g08301(.A(new_n8686_), .B(new_n1108_), .Y(new_n8687_));
  NOR2  g08302(.A(new_n8687_), .B(new_n1112_), .Y(new_n8688_));
  NOR2  g08303(.A(new_n8688_), .B(new_n1117_), .Y(new_n8689_));
  NOR2  g08304(.A(new_n8689_), .B(new_n1121_), .Y(new_n8690_));
  NOR2  g08305(.A(new_n8690_), .B(new_n1126_), .Y(new_n8691_));
  NOR2  g08306(.A(new_n8691_), .B(new_n1130_), .Y(new_n8692_));
  NOR2  g08307(.A(new_n8692_), .B(new_n1135_), .Y(new_n8693_));
  NOR2  g08308(.A(new_n8693_), .B(new_n1139_), .Y(new_n8694_));
  NOR2  g08309(.A(new_n8694_), .B(new_n1144_), .Y(new_n8695_));
  NOR2  g08310(.A(new_n8695_), .B(new_n1148_), .Y(new_n8696_));
  NOR2  g08311(.A(new_n8696_), .B(new_n1153_), .Y(new_n8697_));
  NOR2  g08312(.A(new_n8697_), .B(new_n1157_), .Y(new_n8698_));
  NOR2  g08313(.A(new_n8698_), .B(new_n1162_), .Y(new_n8699_));
  NOR2  g08314(.A(new_n8699_), .B(new_n1166_), .Y(new_n8700_));
  NOR2  g08315(.A(new_n8700_), .B(new_n1171_), .Y(new_n8701_));
  NOR2  g08316(.A(new_n8701_), .B(new_n1175_), .Y(new_n8702_));
  NOR2  g08317(.A(new_n8702_), .B(new_n1180_), .Y(new_n8703_));
  NOR2  g08318(.A(new_n8703_), .B(new_n1184_), .Y(new_n8704_));
  NOR2  g08319(.A(new_n8704_), .B(new_n1189_), .Y(new_n8705_));
  NOR2  g08320(.A(new_n8705_), .B(new_n1707_), .Y(new_n8706_));
  NOR2  g08321(.A(new_n8706_), .B(new_n1709_), .Y(new_n8707_));
  NOR2  g08322(.A(new_n8707_), .B(new_n1973_), .Y(new_n8708_));
  NOR2  g08323(.A(new_n8708_), .B(new_n1199_), .Y(new_n8709_));
  NOR2  g08324(.A(new_n8709_), .B(new_n1203_), .Y(new_n8710_));
  NOR2  g08325(.A(new_n8710_), .B(new_n1207_), .Y(new_n8711_));
  NOR2  g08326(.A(new_n8711_), .B(new_n1211_), .Y(new_n8712_));
  NOR2  g08327(.A(new_n8712_), .B(new_n1215_), .Y(new_n8713_));
  NOR2  g08328(.A(new_n8713_), .B(new_n1219_), .Y(new_n8714_));
  NOR2  g08329(.A(new_n8714_), .B(new_n1223_), .Y(new_n8715_));
  NOR2  g08330(.A(new_n8715_), .B(new_n1227_), .Y(new_n8716_));
  NOR2  g08331(.A(new_n8716_), .B(new_n1231_), .Y(new_n8717_));
  NOR2  g08332(.A(new_n8717_), .B(new_n1235_), .Y(new_n8718_));
  NOR2  g08333(.A(new_n8718_), .B(new_n1239_), .Y(new_n8719_));
  NOR2  g08334(.A(new_n8719_), .B(new_n1243_), .Y(new_n8720_));
  NOR2  g08335(.A(new_n8720_), .B(new_n1247_), .Y(new_n8721_));
  NOR2  g08336(.A(new_n8721_), .B(new_n1251_), .Y(new_n8722_));
  NOR2  g08337(.A(new_n8722_), .B(new_n1255_), .Y(new_n8723_));
  NOR2  g08338(.A(new_n8723_), .B(new_n1259_), .Y(new_n8724_));
  NOR2  g08339(.A(new_n8724_), .B(new_n1263_), .Y(new_n8725_));
  NOR2  g08340(.A(new_n8725_), .B(new_n1267_), .Y(new_n8726_));
  NOR2  g08341(.A(new_n8726_), .B(new_n1271_), .Y(new_n8727_));
  NOR2  g08342(.A(new_n8727_), .B(new_n1275_), .Y(new_n8728_));
  NOR2  g08343(.A(new_n8728_), .B(new_n1279_), .Y(new_n8729_));
  NOR2  g08344(.A(new_n8729_), .B(new_n1283_), .Y(new_n8730_));
  NOR2  g08345(.A(new_n8730_), .B(new_n1287_), .Y(new_n8731_));
  NOR2  g08346(.A(new_n8731_), .B(new_n1291_), .Y(new_n8732_));
  NOR2  g08347(.A(new_n8732_), .B(new_n1295_), .Y(new_n8733_));
  NOR2  g08348(.A(new_n8733_), .B(new_n1299_), .Y(new_n8734_));
  NOR2  g08349(.A(new_n8734_), .B(new_n1303_), .Y(new_n8735_));
  NOR2  g08350(.A(new_n8735_), .B(new_n1307_), .Y(new_n8736_));
  NOR2  g08351(.A(new_n8736_), .B(new_n1311_), .Y(new_n8737_));
  NOR2  g08352(.A(new_n8737_), .B(new_n1315_), .Y(new_n8738_));
  NOR2  g08353(.A(new_n8738_), .B(new_n1319_), .Y(new_n8739_));
  NOR2  g08354(.A(new_n8739_), .B(new_n1323_), .Y(new_n8740_));
  NOR2  g08355(.A(new_n8740_), .B(new_n1327_), .Y(new_n8741_));
  NOR2  g08356(.A(new_n8741_), .B(new_n1331_), .Y(new_n8742_));
  NOR2  g08357(.A(new_n8742_), .B(new_n1335_), .Y(new_n8743_));
  NOR2  g08358(.A(new_n8743_), .B(new_n1339_), .Y(new_n8744_));
  NOR2  g08359(.A(new_n8744_), .B(new_n1343_), .Y(new_n8745_));
  NOR2  g08360(.A(new_n8745_), .B(new_n1347_), .Y(new_n8746_));
  NOR2  g08361(.A(new_n8746_), .B(new_n1351_), .Y(new_n8747_));
  NOR2  g08362(.A(new_n8747_), .B(new_n1355_), .Y(new_n8748_));
  NOR2  g08363(.A(new_n8748_), .B(new_n1359_), .Y(new_n8749_));
  NOR2  g08364(.A(new_n8749_), .B(new_n1363_), .Y(new_n8750_));
  NOR2  g08365(.A(new_n8750_), .B(new_n1367_), .Y(new_n8751_));
  NOR2  g08366(.A(new_n8751_), .B(new_n1371_), .Y(new_n8752_));
  NOR2  g08367(.A(new_n8752_), .B(new_n1375_), .Y(new_n8753_));
  NOR2  g08368(.A(new_n8753_), .B(new_n1379_), .Y(new_n8754_));
  NOR2  g08369(.A(new_n8754_), .B(new_n1383_), .Y(new_n8755_));
  NOR2  g08370(.A(new_n8755_), .B(new_n1387_), .Y(new_n8756_));
  NOR2  g08371(.A(new_n8756_), .B(new_n1391_), .Y(new_n8757_));
  NOR2  g08372(.A(new_n8757_), .B(new_n1395_), .Y(new_n8758_));
  NOR2  g08373(.A(new_n8758_), .B(new_n1399_), .Y(new_n8759_));
  NOR2  g08374(.A(new_n8759_), .B(new_n1403_), .Y(new_n8760_));
  NOR2  g08375(.A(new_n8760_), .B(new_n1407_), .Y(new_n8761_));
  NAND2 g08376(.A(new_n1409_), .B(\req[85] ), .Y(new_n8762_));
  NOR2  g08377(.A(new_n8762_), .B(new_n8761_), .Y(\grant[85] ));
  INV   g08378(.A(new_n1418_), .Y(new_n8764_));
  NOR2  g08379(.A(new_n8764_), .B(new_n675_), .Y(new_n8765_));
  NOR2  g08380(.A(new_n8765_), .B(new_n1423_), .Y(new_n8766_));
  NOR2  g08381(.A(new_n8766_), .B(new_n1427_), .Y(new_n8767_));
  NOR2  g08382(.A(new_n8767_), .B(new_n1431_), .Y(new_n8768_));
  NOR2  g08383(.A(new_n8768_), .B(new_n1435_), .Y(new_n8769_));
  NOR2  g08384(.A(new_n8769_), .B(new_n1439_), .Y(new_n8770_));
  NOR2  g08385(.A(new_n8770_), .B(new_n1443_), .Y(new_n8771_));
  NOR2  g08386(.A(new_n8771_), .B(new_n1447_), .Y(new_n8772_));
  NOR2  g08387(.A(new_n8772_), .B(new_n1451_), .Y(new_n8773_));
  NOR2  g08388(.A(new_n8773_), .B(new_n1455_), .Y(new_n8774_));
  NOR2  g08389(.A(new_n8774_), .B(new_n1459_), .Y(new_n8775_));
  NOR2  g08390(.A(new_n8775_), .B(new_n1463_), .Y(new_n8776_));
  NOR2  g08391(.A(new_n8776_), .B(new_n1467_), .Y(new_n8777_));
  NOR2  g08392(.A(new_n8777_), .B(new_n1471_), .Y(new_n8778_));
  NOR2  g08393(.A(new_n8778_), .B(new_n1475_), .Y(new_n8779_));
  NOR2  g08394(.A(new_n8779_), .B(new_n1479_), .Y(new_n8780_));
  NOR2  g08395(.A(new_n8780_), .B(new_n1483_), .Y(new_n8781_));
  NOR2  g08396(.A(new_n8781_), .B(new_n1487_), .Y(new_n8782_));
  NOR2  g08397(.A(new_n8782_), .B(new_n1491_), .Y(new_n8783_));
  NOR2  g08398(.A(new_n8783_), .B(new_n1495_), .Y(new_n8784_));
  NOR2  g08399(.A(new_n8784_), .B(new_n1499_), .Y(new_n8785_));
  NOR2  g08400(.A(new_n8785_), .B(new_n1503_), .Y(new_n8786_));
  NOR2  g08401(.A(new_n8786_), .B(new_n1507_), .Y(new_n8787_));
  NOR2  g08402(.A(new_n8787_), .B(new_n1511_), .Y(new_n8788_));
  NOR2  g08403(.A(new_n8788_), .B(new_n1515_), .Y(new_n8789_));
  NOR2  g08404(.A(new_n8789_), .B(new_n1519_), .Y(new_n8790_));
  NOR2  g08405(.A(new_n8790_), .B(new_n1523_), .Y(new_n8791_));
  NOR2  g08406(.A(new_n8791_), .B(new_n1527_), .Y(new_n8792_));
  NOR2  g08407(.A(new_n8792_), .B(new_n1797_), .Y(new_n8793_));
  NOR2  g08408(.A(new_n8793_), .B(new_n396_), .Y(new_n8794_));
  NOR2  g08409(.A(new_n8794_), .B(new_n400_), .Y(new_n8795_));
  NOR2  g08410(.A(new_n8795_), .B(new_n406_), .Y(new_n8796_));
  NOR2  g08411(.A(new_n8796_), .B(new_n410_), .Y(new_n8797_));
  NOR2  g08412(.A(new_n8797_), .B(new_n416_), .Y(new_n8798_));
  NOR2  g08413(.A(new_n8798_), .B(new_n420_), .Y(new_n8799_));
  NOR2  g08414(.A(new_n8799_), .B(new_n426_), .Y(new_n8800_));
  NOR2  g08415(.A(new_n8800_), .B(new_n430_), .Y(new_n8801_));
  NOR2  g08416(.A(new_n8801_), .B(new_n436_), .Y(new_n8802_));
  NOR2  g08417(.A(new_n8802_), .B(new_n440_), .Y(new_n8803_));
  NOR2  g08418(.A(new_n8803_), .B(new_n446_), .Y(new_n8804_));
  NOR2  g08419(.A(new_n8804_), .B(new_n450_), .Y(new_n8805_));
  NOR2  g08420(.A(new_n8805_), .B(new_n456_), .Y(new_n8806_));
  NOR2  g08421(.A(new_n8806_), .B(new_n460_), .Y(new_n8807_));
  NOR2  g08422(.A(new_n8807_), .B(new_n466_), .Y(new_n8808_));
  NOR2  g08423(.A(new_n8808_), .B(new_n470_), .Y(new_n8809_));
  NOR2  g08424(.A(new_n8809_), .B(new_n476_), .Y(new_n8810_));
  NOR2  g08425(.A(new_n8810_), .B(new_n480_), .Y(new_n8811_));
  NOR2  g08426(.A(new_n8811_), .B(new_n486_), .Y(new_n8812_));
  NOR2  g08427(.A(new_n8812_), .B(new_n490_), .Y(new_n8813_));
  NOR2  g08428(.A(new_n8813_), .B(new_n496_), .Y(new_n8814_));
  NOR2  g08429(.A(new_n8814_), .B(new_n500_), .Y(new_n8815_));
  NOR2  g08430(.A(new_n8815_), .B(new_n506_), .Y(new_n8816_));
  NOR2  g08431(.A(new_n8816_), .B(new_n510_), .Y(new_n8817_));
  NOR2  g08432(.A(new_n8817_), .B(new_n516_), .Y(new_n8818_));
  NOR2  g08433(.A(new_n8818_), .B(new_n520_), .Y(new_n8819_));
  NOR2  g08434(.A(new_n8819_), .B(new_n526_), .Y(new_n8820_));
  NOR2  g08435(.A(new_n8820_), .B(new_n530_), .Y(new_n8821_));
  NOR2  g08436(.A(new_n8821_), .B(new_n536_), .Y(new_n8822_));
  NOR2  g08437(.A(new_n8822_), .B(new_n540_), .Y(new_n8823_));
  NOR2  g08438(.A(new_n8823_), .B(new_n546_), .Y(new_n8824_));
  NOR2  g08439(.A(new_n8824_), .B(new_n550_), .Y(new_n8825_));
  NOR2  g08440(.A(new_n8825_), .B(new_n556_), .Y(new_n8826_));
  NOR2  g08441(.A(new_n8826_), .B(new_n560_), .Y(new_n8827_));
  NOR2  g08442(.A(new_n8827_), .B(new_n566_), .Y(new_n8828_));
  NOR2  g08443(.A(new_n8828_), .B(new_n570_), .Y(new_n8829_));
  NOR2  g08444(.A(new_n8829_), .B(new_n576_), .Y(new_n8830_));
  NOR2  g08445(.A(new_n8830_), .B(new_n580_), .Y(new_n8831_));
  NOR2  g08446(.A(new_n8831_), .B(new_n586_), .Y(new_n8832_));
  NOR2  g08447(.A(new_n8832_), .B(new_n590_), .Y(new_n8833_));
  NOR2  g08448(.A(new_n8833_), .B(new_n596_), .Y(new_n8834_));
  NOR2  g08449(.A(new_n8834_), .B(new_n600_), .Y(new_n8835_));
  NOR2  g08450(.A(new_n8835_), .B(new_n606_), .Y(new_n8836_));
  NOR2  g08451(.A(new_n8836_), .B(new_n610_), .Y(new_n8837_));
  NOR2  g08452(.A(new_n8837_), .B(new_n616_), .Y(new_n8838_));
  NOR2  g08453(.A(new_n8838_), .B(new_n620_), .Y(new_n8839_));
  NOR2  g08454(.A(new_n8839_), .B(new_n626_), .Y(new_n8840_));
  NOR2  g08455(.A(new_n8840_), .B(new_n630_), .Y(new_n8841_));
  NOR2  g08456(.A(new_n8841_), .B(new_n636_), .Y(new_n8842_));
  NOR2  g08457(.A(new_n8842_), .B(new_n640_), .Y(new_n8843_));
  NOR2  g08458(.A(new_n8843_), .B(new_n646_), .Y(new_n8844_));
  NOR2  g08459(.A(new_n8844_), .B(new_n650_), .Y(new_n8845_));
  NOR2  g08460(.A(new_n8845_), .B(new_n656_), .Y(new_n8846_));
  NOR2  g08461(.A(new_n8846_), .B(new_n660_), .Y(new_n8847_));
  NOR2  g08462(.A(new_n8847_), .B(new_n666_), .Y(new_n8848_));
  NAND2 g08463(.A(new_n668_), .B(\req[86] ), .Y(new_n8849_));
  NOR2  g08464(.A(new_n8849_), .B(new_n8848_), .Y(\grant[86] ));
  INV   g08465(.A(new_n679_), .Y(new_n8851_));
  NOR2  g08466(.A(new_n1071_), .B(new_n8851_), .Y(new_n8852_));
  NOR2  g08467(.A(new_n8852_), .B(new_n686_), .Y(new_n8853_));
  NOR2  g08468(.A(new_n8853_), .B(new_n690_), .Y(new_n8854_));
  NOR2  g08469(.A(new_n8854_), .B(new_n696_), .Y(new_n8855_));
  NOR2  g08470(.A(new_n8855_), .B(new_n700_), .Y(new_n8856_));
  NOR2  g08471(.A(new_n8856_), .B(new_n706_), .Y(new_n8857_));
  NOR2  g08472(.A(new_n8857_), .B(new_n710_), .Y(new_n8858_));
  NOR2  g08473(.A(new_n8858_), .B(new_n716_), .Y(new_n8859_));
  NOR2  g08474(.A(new_n8859_), .B(new_n720_), .Y(new_n8860_));
  NOR2  g08475(.A(new_n8860_), .B(new_n726_), .Y(new_n8861_));
  NOR2  g08476(.A(new_n8861_), .B(new_n730_), .Y(new_n8862_));
  NOR2  g08477(.A(new_n8862_), .B(new_n736_), .Y(new_n8863_));
  NOR2  g08478(.A(new_n8863_), .B(new_n740_), .Y(new_n8864_));
  NOR2  g08479(.A(new_n8864_), .B(new_n746_), .Y(new_n8865_));
  NOR2  g08480(.A(new_n8865_), .B(new_n750_), .Y(new_n8866_));
  NOR2  g08481(.A(new_n8866_), .B(new_n756_), .Y(new_n8867_));
  NOR2  g08482(.A(new_n8867_), .B(new_n760_), .Y(new_n8868_));
  NOR2  g08483(.A(new_n8868_), .B(new_n766_), .Y(new_n8869_));
  NOR2  g08484(.A(new_n8869_), .B(new_n770_), .Y(new_n8870_));
  NOR2  g08485(.A(new_n8870_), .B(new_n776_), .Y(new_n8871_));
  NOR2  g08486(.A(new_n8871_), .B(new_n780_), .Y(new_n8872_));
  NOR2  g08487(.A(new_n8872_), .B(new_n786_), .Y(new_n8873_));
  NOR2  g08488(.A(new_n8873_), .B(new_n790_), .Y(new_n8874_));
  NOR2  g08489(.A(new_n8874_), .B(new_n796_), .Y(new_n8875_));
  NOR2  g08490(.A(new_n8875_), .B(new_n800_), .Y(new_n8876_));
  NOR2  g08491(.A(new_n8876_), .B(new_n806_), .Y(new_n8877_));
  NOR2  g08492(.A(new_n8877_), .B(new_n1616_), .Y(new_n8878_));
  NOR2  g08493(.A(new_n8878_), .B(new_n1618_), .Y(new_n8879_));
  NOR2  g08494(.A(new_n8879_), .B(new_n1885_), .Y(new_n8880_));
  NOR2  g08495(.A(new_n8880_), .B(new_n820_), .Y(new_n8881_));
  NOR2  g08496(.A(new_n8881_), .B(new_n824_), .Y(new_n8882_));
  NOR2  g08497(.A(new_n8882_), .B(new_n829_), .Y(new_n8883_));
  NOR2  g08498(.A(new_n8883_), .B(new_n833_), .Y(new_n8884_));
  NOR2  g08499(.A(new_n8884_), .B(new_n838_), .Y(new_n8885_));
  NOR2  g08500(.A(new_n8885_), .B(new_n842_), .Y(new_n8886_));
  NOR2  g08501(.A(new_n8886_), .B(new_n847_), .Y(new_n8887_));
  NOR2  g08502(.A(new_n8887_), .B(new_n851_), .Y(new_n8888_));
  NOR2  g08503(.A(new_n8888_), .B(new_n856_), .Y(new_n8889_));
  NOR2  g08504(.A(new_n8889_), .B(new_n860_), .Y(new_n8890_));
  NOR2  g08505(.A(new_n8890_), .B(new_n865_), .Y(new_n8891_));
  NOR2  g08506(.A(new_n8891_), .B(new_n869_), .Y(new_n8892_));
  NOR2  g08507(.A(new_n8892_), .B(new_n874_), .Y(new_n8893_));
  NOR2  g08508(.A(new_n8893_), .B(new_n878_), .Y(new_n8894_));
  NOR2  g08509(.A(new_n8894_), .B(new_n883_), .Y(new_n8895_));
  NOR2  g08510(.A(new_n8895_), .B(new_n887_), .Y(new_n8896_));
  NOR2  g08511(.A(new_n8896_), .B(new_n892_), .Y(new_n8897_));
  NOR2  g08512(.A(new_n8897_), .B(new_n896_), .Y(new_n8898_));
  NOR2  g08513(.A(new_n8898_), .B(new_n901_), .Y(new_n8899_));
  NOR2  g08514(.A(new_n8899_), .B(new_n905_), .Y(new_n8900_));
  NOR2  g08515(.A(new_n8900_), .B(new_n910_), .Y(new_n8901_));
  NOR2  g08516(.A(new_n8901_), .B(new_n914_), .Y(new_n8902_));
  NOR2  g08517(.A(new_n8902_), .B(new_n919_), .Y(new_n8903_));
  NOR2  g08518(.A(new_n8903_), .B(new_n923_), .Y(new_n8904_));
  NOR2  g08519(.A(new_n8904_), .B(new_n928_), .Y(new_n8905_));
  NOR2  g08520(.A(new_n8905_), .B(new_n932_), .Y(new_n8906_));
  NOR2  g08521(.A(new_n8906_), .B(new_n937_), .Y(new_n8907_));
  NOR2  g08522(.A(new_n8907_), .B(new_n941_), .Y(new_n8908_));
  NOR2  g08523(.A(new_n8908_), .B(new_n946_), .Y(new_n8909_));
  NOR2  g08524(.A(new_n8909_), .B(new_n950_), .Y(new_n8910_));
  NOR2  g08525(.A(new_n8910_), .B(new_n955_), .Y(new_n8911_));
  NOR2  g08526(.A(new_n8911_), .B(new_n959_), .Y(new_n8912_));
  NOR2  g08527(.A(new_n8912_), .B(new_n964_), .Y(new_n8913_));
  NOR2  g08528(.A(new_n8913_), .B(new_n968_), .Y(new_n8914_));
  NOR2  g08529(.A(new_n8914_), .B(new_n973_), .Y(new_n8915_));
  NOR2  g08530(.A(new_n8915_), .B(new_n977_), .Y(new_n8916_));
  NOR2  g08531(.A(new_n8916_), .B(new_n982_), .Y(new_n8917_));
  NOR2  g08532(.A(new_n8917_), .B(new_n986_), .Y(new_n8918_));
  NOR2  g08533(.A(new_n8918_), .B(new_n991_), .Y(new_n8919_));
  NOR2  g08534(.A(new_n8919_), .B(new_n995_), .Y(new_n8920_));
  NOR2  g08535(.A(new_n8920_), .B(new_n1000_), .Y(new_n8921_));
  NOR2  g08536(.A(new_n8921_), .B(new_n1004_), .Y(new_n8922_));
  NOR2  g08537(.A(new_n8922_), .B(new_n1009_), .Y(new_n8923_));
  NOR2  g08538(.A(new_n8923_), .B(new_n1013_), .Y(new_n8924_));
  NOR2  g08539(.A(new_n8924_), .B(new_n1018_), .Y(new_n8925_));
  NOR2  g08540(.A(new_n8925_), .B(new_n1022_), .Y(new_n8926_));
  NOR2  g08541(.A(new_n8926_), .B(new_n1027_), .Y(new_n8927_));
  NOR2  g08542(.A(new_n8927_), .B(new_n1031_), .Y(new_n8928_));
  NOR2  g08543(.A(new_n8928_), .B(new_n1036_), .Y(new_n8929_));
  NOR2  g08544(.A(new_n8929_), .B(new_n1040_), .Y(new_n8930_));
  NOR2  g08545(.A(new_n8930_), .B(new_n1045_), .Y(new_n8931_));
  NOR2  g08546(.A(new_n8931_), .B(new_n1049_), .Y(new_n8932_));
  NOR2  g08547(.A(new_n8932_), .B(new_n1054_), .Y(new_n8933_));
  NOR2  g08548(.A(new_n8933_), .B(new_n1058_), .Y(new_n8934_));
  NOR2  g08549(.A(new_n8934_), .B(new_n1063_), .Y(new_n8935_));
  NAND2 g08550(.A(new_n1065_), .B(\req[87] ), .Y(new_n8936_));
  NOR2  g08551(.A(new_n8936_), .B(new_n8935_), .Y(\grant[87] ));
  INV   g08552(.A(new_n1075_), .Y(new_n8938_));
  NOR2  g08553(.A(new_n1422_), .B(new_n8938_), .Y(new_n8939_));
  NOR2  g08554(.A(new_n8939_), .B(new_n1081_), .Y(new_n8940_));
  NOR2  g08555(.A(new_n8940_), .B(new_n1085_), .Y(new_n8941_));
  NOR2  g08556(.A(new_n8941_), .B(new_n1090_), .Y(new_n8942_));
  NOR2  g08557(.A(new_n8942_), .B(new_n1094_), .Y(new_n8943_));
  NOR2  g08558(.A(new_n8943_), .B(new_n1099_), .Y(new_n8944_));
  NOR2  g08559(.A(new_n8944_), .B(new_n1103_), .Y(new_n8945_));
  NOR2  g08560(.A(new_n8945_), .B(new_n1108_), .Y(new_n8946_));
  NOR2  g08561(.A(new_n8946_), .B(new_n1112_), .Y(new_n8947_));
  NOR2  g08562(.A(new_n8947_), .B(new_n1117_), .Y(new_n8948_));
  NOR2  g08563(.A(new_n8948_), .B(new_n1121_), .Y(new_n8949_));
  NOR2  g08564(.A(new_n8949_), .B(new_n1126_), .Y(new_n8950_));
  NOR2  g08565(.A(new_n8950_), .B(new_n1130_), .Y(new_n8951_));
  NOR2  g08566(.A(new_n8951_), .B(new_n1135_), .Y(new_n8952_));
  NOR2  g08567(.A(new_n8952_), .B(new_n1139_), .Y(new_n8953_));
  NOR2  g08568(.A(new_n8953_), .B(new_n1144_), .Y(new_n8954_));
  NOR2  g08569(.A(new_n8954_), .B(new_n1148_), .Y(new_n8955_));
  NOR2  g08570(.A(new_n8955_), .B(new_n1153_), .Y(new_n8956_));
  NOR2  g08571(.A(new_n8956_), .B(new_n1157_), .Y(new_n8957_));
  NOR2  g08572(.A(new_n8957_), .B(new_n1162_), .Y(new_n8958_));
  NOR2  g08573(.A(new_n8958_), .B(new_n1166_), .Y(new_n8959_));
  NOR2  g08574(.A(new_n8959_), .B(new_n1171_), .Y(new_n8960_));
  NOR2  g08575(.A(new_n8960_), .B(new_n1175_), .Y(new_n8961_));
  NOR2  g08576(.A(new_n8961_), .B(new_n1180_), .Y(new_n8962_));
  NOR2  g08577(.A(new_n8962_), .B(new_n1184_), .Y(new_n8963_));
  NOR2  g08578(.A(new_n8963_), .B(new_n1189_), .Y(new_n8964_));
  NOR2  g08579(.A(new_n8964_), .B(new_n1707_), .Y(new_n8965_));
  NOR2  g08580(.A(new_n8965_), .B(new_n1709_), .Y(new_n8966_));
  NOR2  g08581(.A(new_n8966_), .B(new_n1973_), .Y(new_n8967_));
  NOR2  g08582(.A(new_n8967_), .B(new_n1199_), .Y(new_n8968_));
  NOR2  g08583(.A(new_n8968_), .B(new_n1203_), .Y(new_n8969_));
  NOR2  g08584(.A(new_n8969_), .B(new_n1207_), .Y(new_n8970_));
  NOR2  g08585(.A(new_n8970_), .B(new_n1211_), .Y(new_n8971_));
  NOR2  g08586(.A(new_n8971_), .B(new_n1215_), .Y(new_n8972_));
  NOR2  g08587(.A(new_n8972_), .B(new_n1219_), .Y(new_n8973_));
  NOR2  g08588(.A(new_n8973_), .B(new_n1223_), .Y(new_n8974_));
  NOR2  g08589(.A(new_n8974_), .B(new_n1227_), .Y(new_n8975_));
  NOR2  g08590(.A(new_n8975_), .B(new_n1231_), .Y(new_n8976_));
  NOR2  g08591(.A(new_n8976_), .B(new_n1235_), .Y(new_n8977_));
  NOR2  g08592(.A(new_n8977_), .B(new_n1239_), .Y(new_n8978_));
  NOR2  g08593(.A(new_n8978_), .B(new_n1243_), .Y(new_n8979_));
  NOR2  g08594(.A(new_n8979_), .B(new_n1247_), .Y(new_n8980_));
  NOR2  g08595(.A(new_n8980_), .B(new_n1251_), .Y(new_n8981_));
  NOR2  g08596(.A(new_n8981_), .B(new_n1255_), .Y(new_n8982_));
  NOR2  g08597(.A(new_n8982_), .B(new_n1259_), .Y(new_n8983_));
  NOR2  g08598(.A(new_n8983_), .B(new_n1263_), .Y(new_n8984_));
  NOR2  g08599(.A(new_n8984_), .B(new_n1267_), .Y(new_n8985_));
  NOR2  g08600(.A(new_n8985_), .B(new_n1271_), .Y(new_n8986_));
  NOR2  g08601(.A(new_n8986_), .B(new_n1275_), .Y(new_n8987_));
  NOR2  g08602(.A(new_n8987_), .B(new_n1279_), .Y(new_n8988_));
  NOR2  g08603(.A(new_n8988_), .B(new_n1283_), .Y(new_n8989_));
  NOR2  g08604(.A(new_n8989_), .B(new_n1287_), .Y(new_n8990_));
  NOR2  g08605(.A(new_n8990_), .B(new_n1291_), .Y(new_n8991_));
  NOR2  g08606(.A(new_n8991_), .B(new_n1295_), .Y(new_n8992_));
  NOR2  g08607(.A(new_n8992_), .B(new_n1299_), .Y(new_n8993_));
  NOR2  g08608(.A(new_n8993_), .B(new_n1303_), .Y(new_n8994_));
  NOR2  g08609(.A(new_n8994_), .B(new_n1307_), .Y(new_n8995_));
  NOR2  g08610(.A(new_n8995_), .B(new_n1311_), .Y(new_n8996_));
  NOR2  g08611(.A(new_n8996_), .B(new_n1315_), .Y(new_n8997_));
  NOR2  g08612(.A(new_n8997_), .B(new_n1319_), .Y(new_n8998_));
  NOR2  g08613(.A(new_n8998_), .B(new_n1323_), .Y(new_n8999_));
  NOR2  g08614(.A(new_n8999_), .B(new_n1327_), .Y(new_n9000_));
  NOR2  g08615(.A(new_n9000_), .B(new_n1331_), .Y(new_n9001_));
  NOR2  g08616(.A(new_n9001_), .B(new_n1335_), .Y(new_n9002_));
  NOR2  g08617(.A(new_n9002_), .B(new_n1339_), .Y(new_n9003_));
  NOR2  g08618(.A(new_n9003_), .B(new_n1343_), .Y(new_n9004_));
  NOR2  g08619(.A(new_n9004_), .B(new_n1347_), .Y(new_n9005_));
  NOR2  g08620(.A(new_n9005_), .B(new_n1351_), .Y(new_n9006_));
  NOR2  g08621(.A(new_n9006_), .B(new_n1355_), .Y(new_n9007_));
  NOR2  g08622(.A(new_n9007_), .B(new_n1359_), .Y(new_n9008_));
  NOR2  g08623(.A(new_n9008_), .B(new_n1363_), .Y(new_n9009_));
  NOR2  g08624(.A(new_n9009_), .B(new_n1367_), .Y(new_n9010_));
  NOR2  g08625(.A(new_n9010_), .B(new_n1371_), .Y(new_n9011_));
  NOR2  g08626(.A(new_n9011_), .B(new_n1375_), .Y(new_n9012_));
  NOR2  g08627(.A(new_n9012_), .B(new_n1379_), .Y(new_n9013_));
  NOR2  g08628(.A(new_n9013_), .B(new_n1383_), .Y(new_n9014_));
  NOR2  g08629(.A(new_n9014_), .B(new_n1387_), .Y(new_n9015_));
  NOR2  g08630(.A(new_n9015_), .B(new_n1391_), .Y(new_n9016_));
  NOR2  g08631(.A(new_n9016_), .B(new_n1395_), .Y(new_n9017_));
  NOR2  g08632(.A(new_n9017_), .B(new_n1399_), .Y(new_n9018_));
  NOR2  g08633(.A(new_n9018_), .B(new_n1403_), .Y(new_n9019_));
  NOR2  g08634(.A(new_n9019_), .B(new_n1407_), .Y(new_n9020_));
  NOR2  g08635(.A(new_n9020_), .B(new_n1411_), .Y(new_n9021_));
  NOR2  g08636(.A(new_n9021_), .B(new_n1415_), .Y(new_n9022_));
  NAND2 g08637(.A(new_n1417_), .B(\req[88] ), .Y(new_n9023_));
  NOR2  g08638(.A(new_n9023_), .B(new_n9022_), .Y(\grant[88] ));
  INV   g08639(.A(new_n1426_), .Y(new_n9025_));
  NOR2  g08640(.A(new_n9025_), .B(new_n685_), .Y(new_n9026_));
  NOR2  g08641(.A(new_n9026_), .B(new_n1431_), .Y(new_n9027_));
  NOR2  g08642(.A(new_n9027_), .B(new_n1435_), .Y(new_n9028_));
  NOR2  g08643(.A(new_n9028_), .B(new_n1439_), .Y(new_n9029_));
  NOR2  g08644(.A(new_n9029_), .B(new_n1443_), .Y(new_n9030_));
  NOR2  g08645(.A(new_n9030_), .B(new_n1447_), .Y(new_n9031_));
  NOR2  g08646(.A(new_n9031_), .B(new_n1451_), .Y(new_n9032_));
  NOR2  g08647(.A(new_n9032_), .B(new_n1455_), .Y(new_n9033_));
  NOR2  g08648(.A(new_n9033_), .B(new_n1459_), .Y(new_n9034_));
  NOR2  g08649(.A(new_n9034_), .B(new_n1463_), .Y(new_n9035_));
  NOR2  g08650(.A(new_n9035_), .B(new_n1467_), .Y(new_n9036_));
  NOR2  g08651(.A(new_n9036_), .B(new_n1471_), .Y(new_n9037_));
  NOR2  g08652(.A(new_n9037_), .B(new_n1475_), .Y(new_n9038_));
  NOR2  g08653(.A(new_n9038_), .B(new_n1479_), .Y(new_n9039_));
  NOR2  g08654(.A(new_n9039_), .B(new_n1483_), .Y(new_n9040_));
  NOR2  g08655(.A(new_n9040_), .B(new_n1487_), .Y(new_n9041_));
  NOR2  g08656(.A(new_n9041_), .B(new_n1491_), .Y(new_n9042_));
  NOR2  g08657(.A(new_n9042_), .B(new_n1495_), .Y(new_n9043_));
  NOR2  g08658(.A(new_n9043_), .B(new_n1499_), .Y(new_n9044_));
  NOR2  g08659(.A(new_n9044_), .B(new_n1503_), .Y(new_n9045_));
  NOR2  g08660(.A(new_n9045_), .B(new_n1507_), .Y(new_n9046_));
  NOR2  g08661(.A(new_n9046_), .B(new_n1511_), .Y(new_n9047_));
  NOR2  g08662(.A(new_n9047_), .B(new_n1515_), .Y(new_n9048_));
  NOR2  g08663(.A(new_n9048_), .B(new_n1519_), .Y(new_n9049_));
  NOR2  g08664(.A(new_n9049_), .B(new_n1523_), .Y(new_n9050_));
  NOR2  g08665(.A(new_n9050_), .B(new_n1527_), .Y(new_n9051_));
  NOR2  g08666(.A(new_n9051_), .B(new_n1797_), .Y(new_n9052_));
  NOR2  g08667(.A(new_n9052_), .B(new_n396_), .Y(new_n9053_));
  NOR2  g08668(.A(new_n9053_), .B(new_n400_), .Y(new_n9054_));
  NOR2  g08669(.A(new_n9054_), .B(new_n406_), .Y(new_n9055_));
  NOR2  g08670(.A(new_n9055_), .B(new_n410_), .Y(new_n9056_));
  NOR2  g08671(.A(new_n9056_), .B(new_n416_), .Y(new_n9057_));
  NOR2  g08672(.A(new_n9057_), .B(new_n420_), .Y(new_n9058_));
  NOR2  g08673(.A(new_n9058_), .B(new_n426_), .Y(new_n9059_));
  NOR2  g08674(.A(new_n9059_), .B(new_n430_), .Y(new_n9060_));
  NOR2  g08675(.A(new_n9060_), .B(new_n436_), .Y(new_n9061_));
  NOR2  g08676(.A(new_n9061_), .B(new_n440_), .Y(new_n9062_));
  NOR2  g08677(.A(new_n9062_), .B(new_n446_), .Y(new_n9063_));
  NOR2  g08678(.A(new_n9063_), .B(new_n450_), .Y(new_n9064_));
  NOR2  g08679(.A(new_n9064_), .B(new_n456_), .Y(new_n9065_));
  NOR2  g08680(.A(new_n9065_), .B(new_n460_), .Y(new_n9066_));
  NOR2  g08681(.A(new_n9066_), .B(new_n466_), .Y(new_n9067_));
  NOR2  g08682(.A(new_n9067_), .B(new_n470_), .Y(new_n9068_));
  NOR2  g08683(.A(new_n9068_), .B(new_n476_), .Y(new_n9069_));
  NOR2  g08684(.A(new_n9069_), .B(new_n480_), .Y(new_n9070_));
  NOR2  g08685(.A(new_n9070_), .B(new_n486_), .Y(new_n9071_));
  NOR2  g08686(.A(new_n9071_), .B(new_n490_), .Y(new_n9072_));
  NOR2  g08687(.A(new_n9072_), .B(new_n496_), .Y(new_n9073_));
  NOR2  g08688(.A(new_n9073_), .B(new_n500_), .Y(new_n9074_));
  NOR2  g08689(.A(new_n9074_), .B(new_n506_), .Y(new_n9075_));
  NOR2  g08690(.A(new_n9075_), .B(new_n510_), .Y(new_n9076_));
  NOR2  g08691(.A(new_n9076_), .B(new_n516_), .Y(new_n9077_));
  NOR2  g08692(.A(new_n9077_), .B(new_n520_), .Y(new_n9078_));
  NOR2  g08693(.A(new_n9078_), .B(new_n526_), .Y(new_n9079_));
  NOR2  g08694(.A(new_n9079_), .B(new_n530_), .Y(new_n9080_));
  NOR2  g08695(.A(new_n9080_), .B(new_n536_), .Y(new_n9081_));
  NOR2  g08696(.A(new_n9081_), .B(new_n540_), .Y(new_n9082_));
  NOR2  g08697(.A(new_n9082_), .B(new_n546_), .Y(new_n9083_));
  NOR2  g08698(.A(new_n9083_), .B(new_n550_), .Y(new_n9084_));
  NOR2  g08699(.A(new_n9084_), .B(new_n556_), .Y(new_n9085_));
  NOR2  g08700(.A(new_n9085_), .B(new_n560_), .Y(new_n9086_));
  NOR2  g08701(.A(new_n9086_), .B(new_n566_), .Y(new_n9087_));
  NOR2  g08702(.A(new_n9087_), .B(new_n570_), .Y(new_n9088_));
  NOR2  g08703(.A(new_n9088_), .B(new_n576_), .Y(new_n9089_));
  NOR2  g08704(.A(new_n9089_), .B(new_n580_), .Y(new_n9090_));
  NOR2  g08705(.A(new_n9090_), .B(new_n586_), .Y(new_n9091_));
  NOR2  g08706(.A(new_n9091_), .B(new_n590_), .Y(new_n9092_));
  NOR2  g08707(.A(new_n9092_), .B(new_n596_), .Y(new_n9093_));
  NOR2  g08708(.A(new_n9093_), .B(new_n600_), .Y(new_n9094_));
  NOR2  g08709(.A(new_n9094_), .B(new_n606_), .Y(new_n9095_));
  NOR2  g08710(.A(new_n9095_), .B(new_n610_), .Y(new_n9096_));
  NOR2  g08711(.A(new_n9096_), .B(new_n616_), .Y(new_n9097_));
  NOR2  g08712(.A(new_n9097_), .B(new_n620_), .Y(new_n9098_));
  NOR2  g08713(.A(new_n9098_), .B(new_n626_), .Y(new_n9099_));
  NOR2  g08714(.A(new_n9099_), .B(new_n630_), .Y(new_n9100_));
  NOR2  g08715(.A(new_n9100_), .B(new_n636_), .Y(new_n9101_));
  NOR2  g08716(.A(new_n9101_), .B(new_n640_), .Y(new_n9102_));
  NOR2  g08717(.A(new_n9102_), .B(new_n646_), .Y(new_n9103_));
  NOR2  g08718(.A(new_n9103_), .B(new_n650_), .Y(new_n9104_));
  NOR2  g08719(.A(new_n9104_), .B(new_n656_), .Y(new_n9105_));
  NOR2  g08720(.A(new_n9105_), .B(new_n660_), .Y(new_n9106_));
  NOR2  g08721(.A(new_n9106_), .B(new_n666_), .Y(new_n9107_));
  NOR2  g08722(.A(new_n9107_), .B(new_n670_), .Y(new_n9108_));
  NOR2  g08723(.A(new_n9108_), .B(new_n676_), .Y(new_n9109_));
  NAND2 g08724(.A(new_n678_), .B(\req[89] ), .Y(new_n9110_));
  NOR2  g08725(.A(new_n9110_), .B(new_n9109_), .Y(\grant[89] ));
  INV   g08726(.A(new_n689_), .Y(new_n9112_));
  NOR2  g08727(.A(new_n1080_), .B(new_n9112_), .Y(new_n9113_));
  NOR2  g08728(.A(new_n9113_), .B(new_n696_), .Y(new_n9114_));
  NOR2  g08729(.A(new_n9114_), .B(new_n700_), .Y(new_n9115_));
  NOR2  g08730(.A(new_n9115_), .B(new_n706_), .Y(new_n9116_));
  NOR2  g08731(.A(new_n9116_), .B(new_n710_), .Y(new_n9117_));
  NOR2  g08732(.A(new_n9117_), .B(new_n716_), .Y(new_n9118_));
  NOR2  g08733(.A(new_n9118_), .B(new_n720_), .Y(new_n9119_));
  NOR2  g08734(.A(new_n9119_), .B(new_n726_), .Y(new_n9120_));
  NOR2  g08735(.A(new_n9120_), .B(new_n730_), .Y(new_n9121_));
  NOR2  g08736(.A(new_n9121_), .B(new_n736_), .Y(new_n9122_));
  NOR2  g08737(.A(new_n9122_), .B(new_n740_), .Y(new_n9123_));
  NOR2  g08738(.A(new_n9123_), .B(new_n746_), .Y(new_n9124_));
  NOR2  g08739(.A(new_n9124_), .B(new_n750_), .Y(new_n9125_));
  NOR2  g08740(.A(new_n9125_), .B(new_n756_), .Y(new_n9126_));
  NOR2  g08741(.A(new_n9126_), .B(new_n760_), .Y(new_n9127_));
  NOR2  g08742(.A(new_n9127_), .B(new_n766_), .Y(new_n9128_));
  NOR2  g08743(.A(new_n9128_), .B(new_n770_), .Y(new_n9129_));
  NOR2  g08744(.A(new_n9129_), .B(new_n776_), .Y(new_n9130_));
  NOR2  g08745(.A(new_n9130_), .B(new_n780_), .Y(new_n9131_));
  NOR2  g08746(.A(new_n9131_), .B(new_n786_), .Y(new_n9132_));
  NOR2  g08747(.A(new_n9132_), .B(new_n790_), .Y(new_n9133_));
  NOR2  g08748(.A(new_n9133_), .B(new_n796_), .Y(new_n9134_));
  NOR2  g08749(.A(new_n9134_), .B(new_n800_), .Y(new_n9135_));
  NOR2  g08750(.A(new_n9135_), .B(new_n806_), .Y(new_n9136_));
  NOR2  g08751(.A(new_n9136_), .B(new_n1616_), .Y(new_n9137_));
  NOR2  g08752(.A(new_n9137_), .B(new_n1618_), .Y(new_n9138_));
  NOR2  g08753(.A(new_n9138_), .B(new_n1885_), .Y(new_n9139_));
  NOR2  g08754(.A(new_n9139_), .B(new_n820_), .Y(new_n9140_));
  NOR2  g08755(.A(new_n9140_), .B(new_n824_), .Y(new_n9141_));
  NOR2  g08756(.A(new_n9141_), .B(new_n829_), .Y(new_n9142_));
  NOR2  g08757(.A(new_n9142_), .B(new_n833_), .Y(new_n9143_));
  NOR2  g08758(.A(new_n9143_), .B(new_n838_), .Y(new_n9144_));
  NOR2  g08759(.A(new_n9144_), .B(new_n842_), .Y(new_n9145_));
  NOR2  g08760(.A(new_n9145_), .B(new_n847_), .Y(new_n9146_));
  NOR2  g08761(.A(new_n9146_), .B(new_n851_), .Y(new_n9147_));
  NOR2  g08762(.A(new_n9147_), .B(new_n856_), .Y(new_n9148_));
  NOR2  g08763(.A(new_n9148_), .B(new_n860_), .Y(new_n9149_));
  NOR2  g08764(.A(new_n9149_), .B(new_n865_), .Y(new_n9150_));
  NOR2  g08765(.A(new_n9150_), .B(new_n869_), .Y(new_n9151_));
  NOR2  g08766(.A(new_n9151_), .B(new_n874_), .Y(new_n9152_));
  NOR2  g08767(.A(new_n9152_), .B(new_n878_), .Y(new_n9153_));
  NOR2  g08768(.A(new_n9153_), .B(new_n883_), .Y(new_n9154_));
  NOR2  g08769(.A(new_n9154_), .B(new_n887_), .Y(new_n9155_));
  NOR2  g08770(.A(new_n9155_), .B(new_n892_), .Y(new_n9156_));
  NOR2  g08771(.A(new_n9156_), .B(new_n896_), .Y(new_n9157_));
  NOR2  g08772(.A(new_n9157_), .B(new_n901_), .Y(new_n9158_));
  NOR2  g08773(.A(new_n9158_), .B(new_n905_), .Y(new_n9159_));
  NOR2  g08774(.A(new_n9159_), .B(new_n910_), .Y(new_n9160_));
  NOR2  g08775(.A(new_n9160_), .B(new_n914_), .Y(new_n9161_));
  NOR2  g08776(.A(new_n9161_), .B(new_n919_), .Y(new_n9162_));
  NOR2  g08777(.A(new_n9162_), .B(new_n923_), .Y(new_n9163_));
  NOR2  g08778(.A(new_n9163_), .B(new_n928_), .Y(new_n9164_));
  NOR2  g08779(.A(new_n9164_), .B(new_n932_), .Y(new_n9165_));
  NOR2  g08780(.A(new_n9165_), .B(new_n937_), .Y(new_n9166_));
  NOR2  g08781(.A(new_n9166_), .B(new_n941_), .Y(new_n9167_));
  NOR2  g08782(.A(new_n9167_), .B(new_n946_), .Y(new_n9168_));
  NOR2  g08783(.A(new_n9168_), .B(new_n950_), .Y(new_n9169_));
  NOR2  g08784(.A(new_n9169_), .B(new_n955_), .Y(new_n9170_));
  NOR2  g08785(.A(new_n9170_), .B(new_n959_), .Y(new_n9171_));
  NOR2  g08786(.A(new_n9171_), .B(new_n964_), .Y(new_n9172_));
  NOR2  g08787(.A(new_n9172_), .B(new_n968_), .Y(new_n9173_));
  NOR2  g08788(.A(new_n9173_), .B(new_n973_), .Y(new_n9174_));
  NOR2  g08789(.A(new_n9174_), .B(new_n977_), .Y(new_n9175_));
  NOR2  g08790(.A(new_n9175_), .B(new_n982_), .Y(new_n9176_));
  NOR2  g08791(.A(new_n9176_), .B(new_n986_), .Y(new_n9177_));
  NOR2  g08792(.A(new_n9177_), .B(new_n991_), .Y(new_n9178_));
  NOR2  g08793(.A(new_n9178_), .B(new_n995_), .Y(new_n9179_));
  NOR2  g08794(.A(new_n9179_), .B(new_n1000_), .Y(new_n9180_));
  NOR2  g08795(.A(new_n9180_), .B(new_n1004_), .Y(new_n9181_));
  NOR2  g08796(.A(new_n9181_), .B(new_n1009_), .Y(new_n9182_));
  NOR2  g08797(.A(new_n9182_), .B(new_n1013_), .Y(new_n9183_));
  NOR2  g08798(.A(new_n9183_), .B(new_n1018_), .Y(new_n9184_));
  NOR2  g08799(.A(new_n9184_), .B(new_n1022_), .Y(new_n9185_));
  NOR2  g08800(.A(new_n9185_), .B(new_n1027_), .Y(new_n9186_));
  NOR2  g08801(.A(new_n9186_), .B(new_n1031_), .Y(new_n9187_));
  NOR2  g08802(.A(new_n9187_), .B(new_n1036_), .Y(new_n9188_));
  NOR2  g08803(.A(new_n9188_), .B(new_n1040_), .Y(new_n9189_));
  NOR2  g08804(.A(new_n9189_), .B(new_n1045_), .Y(new_n9190_));
  NOR2  g08805(.A(new_n9190_), .B(new_n1049_), .Y(new_n9191_));
  NOR2  g08806(.A(new_n9191_), .B(new_n1054_), .Y(new_n9192_));
  NOR2  g08807(.A(new_n9192_), .B(new_n1058_), .Y(new_n9193_));
  NOR2  g08808(.A(new_n9193_), .B(new_n1063_), .Y(new_n9194_));
  NOR2  g08809(.A(new_n9194_), .B(new_n1067_), .Y(new_n9195_));
  NOR2  g08810(.A(new_n9195_), .B(new_n1072_), .Y(new_n9196_));
  NAND2 g08811(.A(new_n1074_), .B(\req[90] ), .Y(new_n9197_));
  NOR2  g08812(.A(new_n9197_), .B(new_n9196_), .Y(\grant[90] ));
  INV   g08813(.A(new_n1084_), .Y(new_n9199_));
  NOR2  g08814(.A(new_n1430_), .B(new_n9199_), .Y(new_n9200_));
  NOR2  g08815(.A(new_n9200_), .B(new_n1090_), .Y(new_n9201_));
  NOR2  g08816(.A(new_n9201_), .B(new_n1094_), .Y(new_n9202_));
  NOR2  g08817(.A(new_n9202_), .B(new_n1099_), .Y(new_n9203_));
  NOR2  g08818(.A(new_n9203_), .B(new_n1103_), .Y(new_n9204_));
  NOR2  g08819(.A(new_n9204_), .B(new_n1108_), .Y(new_n9205_));
  NOR2  g08820(.A(new_n9205_), .B(new_n1112_), .Y(new_n9206_));
  NOR2  g08821(.A(new_n9206_), .B(new_n1117_), .Y(new_n9207_));
  NOR2  g08822(.A(new_n9207_), .B(new_n1121_), .Y(new_n9208_));
  NOR2  g08823(.A(new_n9208_), .B(new_n1126_), .Y(new_n9209_));
  NOR2  g08824(.A(new_n9209_), .B(new_n1130_), .Y(new_n9210_));
  NOR2  g08825(.A(new_n9210_), .B(new_n1135_), .Y(new_n9211_));
  NOR2  g08826(.A(new_n9211_), .B(new_n1139_), .Y(new_n9212_));
  NOR2  g08827(.A(new_n9212_), .B(new_n1144_), .Y(new_n9213_));
  NOR2  g08828(.A(new_n9213_), .B(new_n1148_), .Y(new_n9214_));
  NOR2  g08829(.A(new_n9214_), .B(new_n1153_), .Y(new_n9215_));
  NOR2  g08830(.A(new_n9215_), .B(new_n1157_), .Y(new_n9216_));
  NOR2  g08831(.A(new_n9216_), .B(new_n1162_), .Y(new_n9217_));
  NOR2  g08832(.A(new_n9217_), .B(new_n1166_), .Y(new_n9218_));
  NOR2  g08833(.A(new_n9218_), .B(new_n1171_), .Y(new_n9219_));
  NOR2  g08834(.A(new_n9219_), .B(new_n1175_), .Y(new_n9220_));
  NOR2  g08835(.A(new_n9220_), .B(new_n1180_), .Y(new_n9221_));
  NOR2  g08836(.A(new_n9221_), .B(new_n1184_), .Y(new_n9222_));
  NOR2  g08837(.A(new_n9222_), .B(new_n1189_), .Y(new_n9223_));
  NOR2  g08838(.A(new_n9223_), .B(new_n1707_), .Y(new_n9224_));
  NOR2  g08839(.A(new_n9224_), .B(new_n1709_), .Y(new_n9225_));
  NOR2  g08840(.A(new_n9225_), .B(new_n1973_), .Y(new_n9226_));
  NOR2  g08841(.A(new_n9226_), .B(new_n1199_), .Y(new_n9227_));
  NOR2  g08842(.A(new_n9227_), .B(new_n1203_), .Y(new_n9228_));
  NOR2  g08843(.A(new_n9228_), .B(new_n1207_), .Y(new_n9229_));
  NOR2  g08844(.A(new_n9229_), .B(new_n1211_), .Y(new_n9230_));
  NOR2  g08845(.A(new_n9230_), .B(new_n1215_), .Y(new_n9231_));
  NOR2  g08846(.A(new_n9231_), .B(new_n1219_), .Y(new_n9232_));
  NOR2  g08847(.A(new_n9232_), .B(new_n1223_), .Y(new_n9233_));
  NOR2  g08848(.A(new_n9233_), .B(new_n1227_), .Y(new_n9234_));
  NOR2  g08849(.A(new_n9234_), .B(new_n1231_), .Y(new_n9235_));
  NOR2  g08850(.A(new_n9235_), .B(new_n1235_), .Y(new_n9236_));
  NOR2  g08851(.A(new_n9236_), .B(new_n1239_), .Y(new_n9237_));
  NOR2  g08852(.A(new_n9237_), .B(new_n1243_), .Y(new_n9238_));
  NOR2  g08853(.A(new_n9238_), .B(new_n1247_), .Y(new_n9239_));
  NOR2  g08854(.A(new_n9239_), .B(new_n1251_), .Y(new_n9240_));
  NOR2  g08855(.A(new_n9240_), .B(new_n1255_), .Y(new_n9241_));
  NOR2  g08856(.A(new_n9241_), .B(new_n1259_), .Y(new_n9242_));
  NOR2  g08857(.A(new_n9242_), .B(new_n1263_), .Y(new_n9243_));
  NOR2  g08858(.A(new_n9243_), .B(new_n1267_), .Y(new_n9244_));
  NOR2  g08859(.A(new_n9244_), .B(new_n1271_), .Y(new_n9245_));
  NOR2  g08860(.A(new_n9245_), .B(new_n1275_), .Y(new_n9246_));
  NOR2  g08861(.A(new_n9246_), .B(new_n1279_), .Y(new_n9247_));
  NOR2  g08862(.A(new_n9247_), .B(new_n1283_), .Y(new_n9248_));
  NOR2  g08863(.A(new_n9248_), .B(new_n1287_), .Y(new_n9249_));
  NOR2  g08864(.A(new_n9249_), .B(new_n1291_), .Y(new_n9250_));
  NOR2  g08865(.A(new_n9250_), .B(new_n1295_), .Y(new_n9251_));
  NOR2  g08866(.A(new_n9251_), .B(new_n1299_), .Y(new_n9252_));
  NOR2  g08867(.A(new_n9252_), .B(new_n1303_), .Y(new_n9253_));
  NOR2  g08868(.A(new_n9253_), .B(new_n1307_), .Y(new_n9254_));
  NOR2  g08869(.A(new_n9254_), .B(new_n1311_), .Y(new_n9255_));
  NOR2  g08870(.A(new_n9255_), .B(new_n1315_), .Y(new_n9256_));
  NOR2  g08871(.A(new_n9256_), .B(new_n1319_), .Y(new_n9257_));
  NOR2  g08872(.A(new_n9257_), .B(new_n1323_), .Y(new_n9258_));
  NOR2  g08873(.A(new_n9258_), .B(new_n1327_), .Y(new_n9259_));
  NOR2  g08874(.A(new_n9259_), .B(new_n1331_), .Y(new_n9260_));
  NOR2  g08875(.A(new_n9260_), .B(new_n1335_), .Y(new_n9261_));
  NOR2  g08876(.A(new_n9261_), .B(new_n1339_), .Y(new_n9262_));
  NOR2  g08877(.A(new_n9262_), .B(new_n1343_), .Y(new_n9263_));
  NOR2  g08878(.A(new_n9263_), .B(new_n1347_), .Y(new_n9264_));
  NOR2  g08879(.A(new_n9264_), .B(new_n1351_), .Y(new_n9265_));
  NOR2  g08880(.A(new_n9265_), .B(new_n1355_), .Y(new_n9266_));
  NOR2  g08881(.A(new_n9266_), .B(new_n1359_), .Y(new_n9267_));
  NOR2  g08882(.A(new_n9267_), .B(new_n1363_), .Y(new_n9268_));
  NOR2  g08883(.A(new_n9268_), .B(new_n1367_), .Y(new_n9269_));
  NOR2  g08884(.A(new_n9269_), .B(new_n1371_), .Y(new_n9270_));
  NOR2  g08885(.A(new_n9270_), .B(new_n1375_), .Y(new_n9271_));
  NOR2  g08886(.A(new_n9271_), .B(new_n1379_), .Y(new_n9272_));
  NOR2  g08887(.A(new_n9272_), .B(new_n1383_), .Y(new_n9273_));
  NOR2  g08888(.A(new_n9273_), .B(new_n1387_), .Y(new_n9274_));
  NOR2  g08889(.A(new_n9274_), .B(new_n1391_), .Y(new_n9275_));
  NOR2  g08890(.A(new_n9275_), .B(new_n1395_), .Y(new_n9276_));
  NOR2  g08891(.A(new_n9276_), .B(new_n1399_), .Y(new_n9277_));
  NOR2  g08892(.A(new_n9277_), .B(new_n1403_), .Y(new_n9278_));
  NOR2  g08893(.A(new_n9278_), .B(new_n1407_), .Y(new_n9279_));
  NOR2  g08894(.A(new_n9279_), .B(new_n1411_), .Y(new_n9280_));
  NOR2  g08895(.A(new_n9280_), .B(new_n1415_), .Y(new_n9281_));
  NOR2  g08896(.A(new_n9281_), .B(new_n1419_), .Y(new_n9282_));
  NOR2  g08897(.A(new_n9282_), .B(new_n1423_), .Y(new_n9283_));
  NAND2 g08898(.A(new_n1425_), .B(\req[91] ), .Y(new_n9284_));
  NOR2  g08899(.A(new_n9284_), .B(new_n9283_), .Y(\grant[91] ));
  INV   g08900(.A(new_n1434_), .Y(new_n9286_));
  NOR2  g08901(.A(new_n9286_), .B(new_n695_), .Y(new_n9287_));
  NOR2  g08902(.A(new_n9287_), .B(new_n1439_), .Y(new_n9288_));
  NOR2  g08903(.A(new_n9288_), .B(new_n1443_), .Y(new_n9289_));
  NOR2  g08904(.A(new_n9289_), .B(new_n1447_), .Y(new_n9290_));
  NOR2  g08905(.A(new_n9290_), .B(new_n1451_), .Y(new_n9291_));
  NOR2  g08906(.A(new_n9291_), .B(new_n1455_), .Y(new_n9292_));
  NOR2  g08907(.A(new_n9292_), .B(new_n1459_), .Y(new_n9293_));
  NOR2  g08908(.A(new_n9293_), .B(new_n1463_), .Y(new_n9294_));
  NOR2  g08909(.A(new_n9294_), .B(new_n1467_), .Y(new_n9295_));
  NOR2  g08910(.A(new_n9295_), .B(new_n1471_), .Y(new_n9296_));
  NOR2  g08911(.A(new_n9296_), .B(new_n1475_), .Y(new_n9297_));
  NOR2  g08912(.A(new_n9297_), .B(new_n1479_), .Y(new_n9298_));
  NOR2  g08913(.A(new_n9298_), .B(new_n1483_), .Y(new_n9299_));
  NOR2  g08914(.A(new_n9299_), .B(new_n1487_), .Y(new_n9300_));
  NOR2  g08915(.A(new_n9300_), .B(new_n1491_), .Y(new_n9301_));
  NOR2  g08916(.A(new_n9301_), .B(new_n1495_), .Y(new_n9302_));
  NOR2  g08917(.A(new_n9302_), .B(new_n1499_), .Y(new_n9303_));
  NOR2  g08918(.A(new_n9303_), .B(new_n1503_), .Y(new_n9304_));
  NOR2  g08919(.A(new_n9304_), .B(new_n1507_), .Y(new_n9305_));
  NOR2  g08920(.A(new_n9305_), .B(new_n1511_), .Y(new_n9306_));
  NOR2  g08921(.A(new_n9306_), .B(new_n1515_), .Y(new_n9307_));
  NOR2  g08922(.A(new_n9307_), .B(new_n1519_), .Y(new_n9308_));
  NOR2  g08923(.A(new_n9308_), .B(new_n1523_), .Y(new_n9309_));
  NOR2  g08924(.A(new_n9309_), .B(new_n1527_), .Y(new_n9310_));
  NOR2  g08925(.A(new_n9310_), .B(new_n1797_), .Y(new_n9311_));
  NOR2  g08926(.A(new_n9311_), .B(new_n396_), .Y(new_n9312_));
  NOR2  g08927(.A(new_n9312_), .B(new_n400_), .Y(new_n9313_));
  NOR2  g08928(.A(new_n9313_), .B(new_n406_), .Y(new_n9314_));
  NOR2  g08929(.A(new_n9314_), .B(new_n410_), .Y(new_n9315_));
  NOR2  g08930(.A(new_n9315_), .B(new_n416_), .Y(new_n9316_));
  NOR2  g08931(.A(new_n9316_), .B(new_n420_), .Y(new_n9317_));
  NOR2  g08932(.A(new_n9317_), .B(new_n426_), .Y(new_n9318_));
  NOR2  g08933(.A(new_n9318_), .B(new_n430_), .Y(new_n9319_));
  NOR2  g08934(.A(new_n9319_), .B(new_n436_), .Y(new_n9320_));
  NOR2  g08935(.A(new_n9320_), .B(new_n440_), .Y(new_n9321_));
  NOR2  g08936(.A(new_n9321_), .B(new_n446_), .Y(new_n9322_));
  NOR2  g08937(.A(new_n9322_), .B(new_n450_), .Y(new_n9323_));
  NOR2  g08938(.A(new_n9323_), .B(new_n456_), .Y(new_n9324_));
  NOR2  g08939(.A(new_n9324_), .B(new_n460_), .Y(new_n9325_));
  NOR2  g08940(.A(new_n9325_), .B(new_n466_), .Y(new_n9326_));
  NOR2  g08941(.A(new_n9326_), .B(new_n470_), .Y(new_n9327_));
  NOR2  g08942(.A(new_n9327_), .B(new_n476_), .Y(new_n9328_));
  NOR2  g08943(.A(new_n9328_), .B(new_n480_), .Y(new_n9329_));
  NOR2  g08944(.A(new_n9329_), .B(new_n486_), .Y(new_n9330_));
  NOR2  g08945(.A(new_n9330_), .B(new_n490_), .Y(new_n9331_));
  NOR2  g08946(.A(new_n9331_), .B(new_n496_), .Y(new_n9332_));
  NOR2  g08947(.A(new_n9332_), .B(new_n500_), .Y(new_n9333_));
  NOR2  g08948(.A(new_n9333_), .B(new_n506_), .Y(new_n9334_));
  NOR2  g08949(.A(new_n9334_), .B(new_n510_), .Y(new_n9335_));
  NOR2  g08950(.A(new_n9335_), .B(new_n516_), .Y(new_n9336_));
  NOR2  g08951(.A(new_n9336_), .B(new_n520_), .Y(new_n9337_));
  NOR2  g08952(.A(new_n9337_), .B(new_n526_), .Y(new_n9338_));
  NOR2  g08953(.A(new_n9338_), .B(new_n530_), .Y(new_n9339_));
  NOR2  g08954(.A(new_n9339_), .B(new_n536_), .Y(new_n9340_));
  NOR2  g08955(.A(new_n9340_), .B(new_n540_), .Y(new_n9341_));
  NOR2  g08956(.A(new_n9341_), .B(new_n546_), .Y(new_n9342_));
  NOR2  g08957(.A(new_n9342_), .B(new_n550_), .Y(new_n9343_));
  NOR2  g08958(.A(new_n9343_), .B(new_n556_), .Y(new_n9344_));
  NOR2  g08959(.A(new_n9344_), .B(new_n560_), .Y(new_n9345_));
  NOR2  g08960(.A(new_n9345_), .B(new_n566_), .Y(new_n9346_));
  NOR2  g08961(.A(new_n9346_), .B(new_n570_), .Y(new_n9347_));
  NOR2  g08962(.A(new_n9347_), .B(new_n576_), .Y(new_n9348_));
  NOR2  g08963(.A(new_n9348_), .B(new_n580_), .Y(new_n9349_));
  NOR2  g08964(.A(new_n9349_), .B(new_n586_), .Y(new_n9350_));
  NOR2  g08965(.A(new_n9350_), .B(new_n590_), .Y(new_n9351_));
  NOR2  g08966(.A(new_n9351_), .B(new_n596_), .Y(new_n9352_));
  NOR2  g08967(.A(new_n9352_), .B(new_n600_), .Y(new_n9353_));
  NOR2  g08968(.A(new_n9353_), .B(new_n606_), .Y(new_n9354_));
  NOR2  g08969(.A(new_n9354_), .B(new_n610_), .Y(new_n9355_));
  NOR2  g08970(.A(new_n9355_), .B(new_n616_), .Y(new_n9356_));
  NOR2  g08971(.A(new_n9356_), .B(new_n620_), .Y(new_n9357_));
  NOR2  g08972(.A(new_n9357_), .B(new_n626_), .Y(new_n9358_));
  NOR2  g08973(.A(new_n9358_), .B(new_n630_), .Y(new_n9359_));
  NOR2  g08974(.A(new_n9359_), .B(new_n636_), .Y(new_n9360_));
  NOR2  g08975(.A(new_n9360_), .B(new_n640_), .Y(new_n9361_));
  NOR2  g08976(.A(new_n9361_), .B(new_n646_), .Y(new_n9362_));
  NOR2  g08977(.A(new_n9362_), .B(new_n650_), .Y(new_n9363_));
  NOR2  g08978(.A(new_n9363_), .B(new_n656_), .Y(new_n9364_));
  NOR2  g08979(.A(new_n9364_), .B(new_n660_), .Y(new_n9365_));
  NOR2  g08980(.A(new_n9365_), .B(new_n666_), .Y(new_n9366_));
  NOR2  g08981(.A(new_n9366_), .B(new_n670_), .Y(new_n9367_));
  NOR2  g08982(.A(new_n9367_), .B(new_n676_), .Y(new_n9368_));
  NOR2  g08983(.A(new_n9368_), .B(new_n680_), .Y(new_n9369_));
  NOR2  g08984(.A(new_n9369_), .B(new_n686_), .Y(new_n9370_));
  NAND2 g08985(.A(new_n688_), .B(\req[92] ), .Y(new_n9371_));
  NOR2  g08986(.A(new_n9371_), .B(new_n9370_), .Y(\grant[92] ));
  INV   g08987(.A(new_n699_), .Y(new_n9373_));
  NOR2  g08988(.A(new_n1089_), .B(new_n9373_), .Y(new_n9374_));
  NOR2  g08989(.A(new_n9374_), .B(new_n706_), .Y(new_n9375_));
  NOR2  g08990(.A(new_n9375_), .B(new_n710_), .Y(new_n9376_));
  NOR2  g08991(.A(new_n9376_), .B(new_n716_), .Y(new_n9377_));
  NOR2  g08992(.A(new_n9377_), .B(new_n720_), .Y(new_n9378_));
  NOR2  g08993(.A(new_n9378_), .B(new_n726_), .Y(new_n9379_));
  NOR2  g08994(.A(new_n9379_), .B(new_n730_), .Y(new_n9380_));
  NOR2  g08995(.A(new_n9380_), .B(new_n736_), .Y(new_n9381_));
  NOR2  g08996(.A(new_n9381_), .B(new_n740_), .Y(new_n9382_));
  NOR2  g08997(.A(new_n9382_), .B(new_n746_), .Y(new_n9383_));
  NOR2  g08998(.A(new_n9383_), .B(new_n750_), .Y(new_n9384_));
  NOR2  g08999(.A(new_n9384_), .B(new_n756_), .Y(new_n9385_));
  NOR2  g09000(.A(new_n9385_), .B(new_n760_), .Y(new_n9386_));
  NOR2  g09001(.A(new_n9386_), .B(new_n766_), .Y(new_n9387_));
  NOR2  g09002(.A(new_n9387_), .B(new_n770_), .Y(new_n9388_));
  NOR2  g09003(.A(new_n9388_), .B(new_n776_), .Y(new_n9389_));
  NOR2  g09004(.A(new_n9389_), .B(new_n780_), .Y(new_n9390_));
  NOR2  g09005(.A(new_n9390_), .B(new_n786_), .Y(new_n9391_));
  NOR2  g09006(.A(new_n9391_), .B(new_n790_), .Y(new_n9392_));
  NOR2  g09007(.A(new_n9392_), .B(new_n796_), .Y(new_n9393_));
  NOR2  g09008(.A(new_n9393_), .B(new_n800_), .Y(new_n9394_));
  NOR2  g09009(.A(new_n9394_), .B(new_n806_), .Y(new_n9395_));
  NOR2  g09010(.A(new_n9395_), .B(new_n1616_), .Y(new_n9396_));
  NOR2  g09011(.A(new_n9396_), .B(new_n1618_), .Y(new_n9397_));
  NOR2  g09012(.A(new_n9397_), .B(new_n1885_), .Y(new_n9398_));
  NOR2  g09013(.A(new_n9398_), .B(new_n820_), .Y(new_n9399_));
  NOR2  g09014(.A(new_n9399_), .B(new_n824_), .Y(new_n9400_));
  NOR2  g09015(.A(new_n9400_), .B(new_n829_), .Y(new_n9401_));
  NOR2  g09016(.A(new_n9401_), .B(new_n833_), .Y(new_n9402_));
  NOR2  g09017(.A(new_n9402_), .B(new_n838_), .Y(new_n9403_));
  NOR2  g09018(.A(new_n9403_), .B(new_n842_), .Y(new_n9404_));
  NOR2  g09019(.A(new_n9404_), .B(new_n847_), .Y(new_n9405_));
  NOR2  g09020(.A(new_n9405_), .B(new_n851_), .Y(new_n9406_));
  NOR2  g09021(.A(new_n9406_), .B(new_n856_), .Y(new_n9407_));
  NOR2  g09022(.A(new_n9407_), .B(new_n860_), .Y(new_n9408_));
  NOR2  g09023(.A(new_n9408_), .B(new_n865_), .Y(new_n9409_));
  NOR2  g09024(.A(new_n9409_), .B(new_n869_), .Y(new_n9410_));
  NOR2  g09025(.A(new_n9410_), .B(new_n874_), .Y(new_n9411_));
  NOR2  g09026(.A(new_n9411_), .B(new_n878_), .Y(new_n9412_));
  NOR2  g09027(.A(new_n9412_), .B(new_n883_), .Y(new_n9413_));
  NOR2  g09028(.A(new_n9413_), .B(new_n887_), .Y(new_n9414_));
  NOR2  g09029(.A(new_n9414_), .B(new_n892_), .Y(new_n9415_));
  NOR2  g09030(.A(new_n9415_), .B(new_n896_), .Y(new_n9416_));
  NOR2  g09031(.A(new_n9416_), .B(new_n901_), .Y(new_n9417_));
  NOR2  g09032(.A(new_n9417_), .B(new_n905_), .Y(new_n9418_));
  NOR2  g09033(.A(new_n9418_), .B(new_n910_), .Y(new_n9419_));
  NOR2  g09034(.A(new_n9419_), .B(new_n914_), .Y(new_n9420_));
  NOR2  g09035(.A(new_n9420_), .B(new_n919_), .Y(new_n9421_));
  NOR2  g09036(.A(new_n9421_), .B(new_n923_), .Y(new_n9422_));
  NOR2  g09037(.A(new_n9422_), .B(new_n928_), .Y(new_n9423_));
  NOR2  g09038(.A(new_n9423_), .B(new_n932_), .Y(new_n9424_));
  NOR2  g09039(.A(new_n9424_), .B(new_n937_), .Y(new_n9425_));
  NOR2  g09040(.A(new_n9425_), .B(new_n941_), .Y(new_n9426_));
  NOR2  g09041(.A(new_n9426_), .B(new_n946_), .Y(new_n9427_));
  NOR2  g09042(.A(new_n9427_), .B(new_n950_), .Y(new_n9428_));
  NOR2  g09043(.A(new_n9428_), .B(new_n955_), .Y(new_n9429_));
  NOR2  g09044(.A(new_n9429_), .B(new_n959_), .Y(new_n9430_));
  NOR2  g09045(.A(new_n9430_), .B(new_n964_), .Y(new_n9431_));
  NOR2  g09046(.A(new_n9431_), .B(new_n968_), .Y(new_n9432_));
  NOR2  g09047(.A(new_n9432_), .B(new_n973_), .Y(new_n9433_));
  NOR2  g09048(.A(new_n9433_), .B(new_n977_), .Y(new_n9434_));
  NOR2  g09049(.A(new_n9434_), .B(new_n982_), .Y(new_n9435_));
  NOR2  g09050(.A(new_n9435_), .B(new_n986_), .Y(new_n9436_));
  NOR2  g09051(.A(new_n9436_), .B(new_n991_), .Y(new_n9437_));
  NOR2  g09052(.A(new_n9437_), .B(new_n995_), .Y(new_n9438_));
  NOR2  g09053(.A(new_n9438_), .B(new_n1000_), .Y(new_n9439_));
  NOR2  g09054(.A(new_n9439_), .B(new_n1004_), .Y(new_n9440_));
  NOR2  g09055(.A(new_n9440_), .B(new_n1009_), .Y(new_n9441_));
  NOR2  g09056(.A(new_n9441_), .B(new_n1013_), .Y(new_n9442_));
  NOR2  g09057(.A(new_n9442_), .B(new_n1018_), .Y(new_n9443_));
  NOR2  g09058(.A(new_n9443_), .B(new_n1022_), .Y(new_n9444_));
  NOR2  g09059(.A(new_n9444_), .B(new_n1027_), .Y(new_n9445_));
  NOR2  g09060(.A(new_n9445_), .B(new_n1031_), .Y(new_n9446_));
  NOR2  g09061(.A(new_n9446_), .B(new_n1036_), .Y(new_n9447_));
  NOR2  g09062(.A(new_n9447_), .B(new_n1040_), .Y(new_n9448_));
  NOR2  g09063(.A(new_n9448_), .B(new_n1045_), .Y(new_n9449_));
  NOR2  g09064(.A(new_n9449_), .B(new_n1049_), .Y(new_n9450_));
  NOR2  g09065(.A(new_n9450_), .B(new_n1054_), .Y(new_n9451_));
  NOR2  g09066(.A(new_n9451_), .B(new_n1058_), .Y(new_n9452_));
  NOR2  g09067(.A(new_n9452_), .B(new_n1063_), .Y(new_n9453_));
  NOR2  g09068(.A(new_n9453_), .B(new_n1067_), .Y(new_n9454_));
  NOR2  g09069(.A(new_n9454_), .B(new_n1072_), .Y(new_n9455_));
  NOR2  g09070(.A(new_n9455_), .B(new_n1076_), .Y(new_n9456_));
  NOR2  g09071(.A(new_n9456_), .B(new_n1081_), .Y(new_n9457_));
  NAND2 g09072(.A(new_n1083_), .B(\req[93] ), .Y(new_n9458_));
  NOR2  g09073(.A(new_n9458_), .B(new_n9457_), .Y(\grant[93] ));
  INV   g09074(.A(new_n1093_), .Y(new_n9460_));
  NOR2  g09075(.A(new_n1438_), .B(new_n9460_), .Y(new_n9461_));
  NOR2  g09076(.A(new_n9461_), .B(new_n1099_), .Y(new_n9462_));
  NOR2  g09077(.A(new_n9462_), .B(new_n1103_), .Y(new_n9463_));
  NOR2  g09078(.A(new_n9463_), .B(new_n1108_), .Y(new_n9464_));
  NOR2  g09079(.A(new_n9464_), .B(new_n1112_), .Y(new_n9465_));
  NOR2  g09080(.A(new_n9465_), .B(new_n1117_), .Y(new_n9466_));
  NOR2  g09081(.A(new_n9466_), .B(new_n1121_), .Y(new_n9467_));
  NOR2  g09082(.A(new_n9467_), .B(new_n1126_), .Y(new_n9468_));
  NOR2  g09083(.A(new_n9468_), .B(new_n1130_), .Y(new_n9469_));
  NOR2  g09084(.A(new_n9469_), .B(new_n1135_), .Y(new_n9470_));
  NOR2  g09085(.A(new_n9470_), .B(new_n1139_), .Y(new_n9471_));
  NOR2  g09086(.A(new_n9471_), .B(new_n1144_), .Y(new_n9472_));
  NOR2  g09087(.A(new_n9472_), .B(new_n1148_), .Y(new_n9473_));
  NOR2  g09088(.A(new_n9473_), .B(new_n1153_), .Y(new_n9474_));
  NOR2  g09089(.A(new_n9474_), .B(new_n1157_), .Y(new_n9475_));
  NOR2  g09090(.A(new_n9475_), .B(new_n1162_), .Y(new_n9476_));
  NOR2  g09091(.A(new_n9476_), .B(new_n1166_), .Y(new_n9477_));
  NOR2  g09092(.A(new_n9477_), .B(new_n1171_), .Y(new_n9478_));
  NOR2  g09093(.A(new_n9478_), .B(new_n1175_), .Y(new_n9479_));
  NOR2  g09094(.A(new_n9479_), .B(new_n1180_), .Y(new_n9480_));
  NOR2  g09095(.A(new_n9480_), .B(new_n1184_), .Y(new_n9481_));
  NOR2  g09096(.A(new_n9481_), .B(new_n1189_), .Y(new_n9482_));
  NOR2  g09097(.A(new_n9482_), .B(new_n1707_), .Y(new_n9483_));
  NOR2  g09098(.A(new_n9483_), .B(new_n1709_), .Y(new_n9484_));
  NOR2  g09099(.A(new_n9484_), .B(new_n1973_), .Y(new_n9485_));
  NOR2  g09100(.A(new_n9485_), .B(new_n1199_), .Y(new_n9486_));
  NOR2  g09101(.A(new_n9486_), .B(new_n1203_), .Y(new_n9487_));
  NOR2  g09102(.A(new_n9487_), .B(new_n1207_), .Y(new_n9488_));
  NOR2  g09103(.A(new_n9488_), .B(new_n1211_), .Y(new_n9489_));
  NOR2  g09104(.A(new_n9489_), .B(new_n1215_), .Y(new_n9490_));
  NOR2  g09105(.A(new_n9490_), .B(new_n1219_), .Y(new_n9491_));
  NOR2  g09106(.A(new_n9491_), .B(new_n1223_), .Y(new_n9492_));
  NOR2  g09107(.A(new_n9492_), .B(new_n1227_), .Y(new_n9493_));
  NOR2  g09108(.A(new_n9493_), .B(new_n1231_), .Y(new_n9494_));
  NOR2  g09109(.A(new_n9494_), .B(new_n1235_), .Y(new_n9495_));
  NOR2  g09110(.A(new_n9495_), .B(new_n1239_), .Y(new_n9496_));
  NOR2  g09111(.A(new_n9496_), .B(new_n1243_), .Y(new_n9497_));
  NOR2  g09112(.A(new_n9497_), .B(new_n1247_), .Y(new_n9498_));
  NOR2  g09113(.A(new_n9498_), .B(new_n1251_), .Y(new_n9499_));
  NOR2  g09114(.A(new_n9499_), .B(new_n1255_), .Y(new_n9500_));
  NOR2  g09115(.A(new_n9500_), .B(new_n1259_), .Y(new_n9501_));
  NOR2  g09116(.A(new_n9501_), .B(new_n1263_), .Y(new_n9502_));
  NOR2  g09117(.A(new_n9502_), .B(new_n1267_), .Y(new_n9503_));
  NOR2  g09118(.A(new_n9503_), .B(new_n1271_), .Y(new_n9504_));
  NOR2  g09119(.A(new_n9504_), .B(new_n1275_), .Y(new_n9505_));
  NOR2  g09120(.A(new_n9505_), .B(new_n1279_), .Y(new_n9506_));
  NOR2  g09121(.A(new_n9506_), .B(new_n1283_), .Y(new_n9507_));
  NOR2  g09122(.A(new_n9507_), .B(new_n1287_), .Y(new_n9508_));
  NOR2  g09123(.A(new_n9508_), .B(new_n1291_), .Y(new_n9509_));
  NOR2  g09124(.A(new_n9509_), .B(new_n1295_), .Y(new_n9510_));
  NOR2  g09125(.A(new_n9510_), .B(new_n1299_), .Y(new_n9511_));
  NOR2  g09126(.A(new_n9511_), .B(new_n1303_), .Y(new_n9512_));
  NOR2  g09127(.A(new_n9512_), .B(new_n1307_), .Y(new_n9513_));
  NOR2  g09128(.A(new_n9513_), .B(new_n1311_), .Y(new_n9514_));
  NOR2  g09129(.A(new_n9514_), .B(new_n1315_), .Y(new_n9515_));
  NOR2  g09130(.A(new_n9515_), .B(new_n1319_), .Y(new_n9516_));
  NOR2  g09131(.A(new_n9516_), .B(new_n1323_), .Y(new_n9517_));
  NOR2  g09132(.A(new_n9517_), .B(new_n1327_), .Y(new_n9518_));
  NOR2  g09133(.A(new_n9518_), .B(new_n1331_), .Y(new_n9519_));
  NOR2  g09134(.A(new_n9519_), .B(new_n1335_), .Y(new_n9520_));
  NOR2  g09135(.A(new_n9520_), .B(new_n1339_), .Y(new_n9521_));
  NOR2  g09136(.A(new_n9521_), .B(new_n1343_), .Y(new_n9522_));
  NOR2  g09137(.A(new_n9522_), .B(new_n1347_), .Y(new_n9523_));
  NOR2  g09138(.A(new_n9523_), .B(new_n1351_), .Y(new_n9524_));
  NOR2  g09139(.A(new_n9524_), .B(new_n1355_), .Y(new_n9525_));
  NOR2  g09140(.A(new_n9525_), .B(new_n1359_), .Y(new_n9526_));
  NOR2  g09141(.A(new_n9526_), .B(new_n1363_), .Y(new_n9527_));
  NOR2  g09142(.A(new_n9527_), .B(new_n1367_), .Y(new_n9528_));
  NOR2  g09143(.A(new_n9528_), .B(new_n1371_), .Y(new_n9529_));
  NOR2  g09144(.A(new_n9529_), .B(new_n1375_), .Y(new_n9530_));
  NOR2  g09145(.A(new_n9530_), .B(new_n1379_), .Y(new_n9531_));
  NOR2  g09146(.A(new_n9531_), .B(new_n1383_), .Y(new_n9532_));
  NOR2  g09147(.A(new_n9532_), .B(new_n1387_), .Y(new_n9533_));
  NOR2  g09148(.A(new_n9533_), .B(new_n1391_), .Y(new_n9534_));
  NOR2  g09149(.A(new_n9534_), .B(new_n1395_), .Y(new_n9535_));
  NOR2  g09150(.A(new_n9535_), .B(new_n1399_), .Y(new_n9536_));
  NOR2  g09151(.A(new_n9536_), .B(new_n1403_), .Y(new_n9537_));
  NOR2  g09152(.A(new_n9537_), .B(new_n1407_), .Y(new_n9538_));
  NOR2  g09153(.A(new_n9538_), .B(new_n1411_), .Y(new_n9539_));
  NOR2  g09154(.A(new_n9539_), .B(new_n1415_), .Y(new_n9540_));
  NOR2  g09155(.A(new_n9540_), .B(new_n1419_), .Y(new_n9541_));
  NOR2  g09156(.A(new_n9541_), .B(new_n1423_), .Y(new_n9542_));
  NOR2  g09157(.A(new_n9542_), .B(new_n1427_), .Y(new_n9543_));
  NOR2  g09158(.A(new_n9543_), .B(new_n1431_), .Y(new_n9544_));
  NAND2 g09159(.A(new_n1433_), .B(\req[94] ), .Y(new_n9545_));
  NOR2  g09160(.A(new_n9545_), .B(new_n9544_), .Y(\grant[94] ));
  INV   g09161(.A(new_n1442_), .Y(new_n9547_));
  NOR2  g09162(.A(new_n9547_), .B(new_n705_), .Y(new_n9548_));
  NOR2  g09163(.A(new_n9548_), .B(new_n1447_), .Y(new_n9549_));
  NOR2  g09164(.A(new_n9549_), .B(new_n1451_), .Y(new_n9550_));
  NOR2  g09165(.A(new_n9550_), .B(new_n1455_), .Y(new_n9551_));
  NOR2  g09166(.A(new_n9551_), .B(new_n1459_), .Y(new_n9552_));
  NOR2  g09167(.A(new_n9552_), .B(new_n1463_), .Y(new_n9553_));
  NOR2  g09168(.A(new_n9553_), .B(new_n1467_), .Y(new_n9554_));
  NOR2  g09169(.A(new_n9554_), .B(new_n1471_), .Y(new_n9555_));
  NOR2  g09170(.A(new_n9555_), .B(new_n1475_), .Y(new_n9556_));
  NOR2  g09171(.A(new_n9556_), .B(new_n1479_), .Y(new_n9557_));
  NOR2  g09172(.A(new_n9557_), .B(new_n1483_), .Y(new_n9558_));
  NOR2  g09173(.A(new_n9558_), .B(new_n1487_), .Y(new_n9559_));
  NOR2  g09174(.A(new_n9559_), .B(new_n1491_), .Y(new_n9560_));
  NOR2  g09175(.A(new_n9560_), .B(new_n1495_), .Y(new_n9561_));
  NOR2  g09176(.A(new_n9561_), .B(new_n1499_), .Y(new_n9562_));
  NOR2  g09177(.A(new_n9562_), .B(new_n1503_), .Y(new_n9563_));
  NOR2  g09178(.A(new_n9563_), .B(new_n1507_), .Y(new_n9564_));
  NOR2  g09179(.A(new_n9564_), .B(new_n1511_), .Y(new_n9565_));
  NOR2  g09180(.A(new_n9565_), .B(new_n1515_), .Y(new_n9566_));
  NOR2  g09181(.A(new_n9566_), .B(new_n1519_), .Y(new_n9567_));
  NOR2  g09182(.A(new_n9567_), .B(new_n1523_), .Y(new_n9568_));
  NOR2  g09183(.A(new_n9568_), .B(new_n1527_), .Y(new_n9569_));
  NOR2  g09184(.A(new_n9569_), .B(new_n1797_), .Y(new_n9570_));
  NOR2  g09185(.A(new_n9570_), .B(new_n396_), .Y(new_n9571_));
  NOR2  g09186(.A(new_n9571_), .B(new_n400_), .Y(new_n9572_));
  NOR2  g09187(.A(new_n9572_), .B(new_n406_), .Y(new_n9573_));
  NOR2  g09188(.A(new_n9573_), .B(new_n410_), .Y(new_n9574_));
  NOR2  g09189(.A(new_n9574_), .B(new_n416_), .Y(new_n9575_));
  NOR2  g09190(.A(new_n9575_), .B(new_n420_), .Y(new_n9576_));
  NOR2  g09191(.A(new_n9576_), .B(new_n426_), .Y(new_n9577_));
  NOR2  g09192(.A(new_n9577_), .B(new_n430_), .Y(new_n9578_));
  NOR2  g09193(.A(new_n9578_), .B(new_n436_), .Y(new_n9579_));
  NOR2  g09194(.A(new_n9579_), .B(new_n440_), .Y(new_n9580_));
  NOR2  g09195(.A(new_n9580_), .B(new_n446_), .Y(new_n9581_));
  NOR2  g09196(.A(new_n9581_), .B(new_n450_), .Y(new_n9582_));
  NOR2  g09197(.A(new_n9582_), .B(new_n456_), .Y(new_n9583_));
  NOR2  g09198(.A(new_n9583_), .B(new_n460_), .Y(new_n9584_));
  NOR2  g09199(.A(new_n9584_), .B(new_n466_), .Y(new_n9585_));
  NOR2  g09200(.A(new_n9585_), .B(new_n470_), .Y(new_n9586_));
  NOR2  g09201(.A(new_n9586_), .B(new_n476_), .Y(new_n9587_));
  NOR2  g09202(.A(new_n9587_), .B(new_n480_), .Y(new_n9588_));
  NOR2  g09203(.A(new_n9588_), .B(new_n486_), .Y(new_n9589_));
  NOR2  g09204(.A(new_n9589_), .B(new_n490_), .Y(new_n9590_));
  NOR2  g09205(.A(new_n9590_), .B(new_n496_), .Y(new_n9591_));
  NOR2  g09206(.A(new_n9591_), .B(new_n500_), .Y(new_n9592_));
  NOR2  g09207(.A(new_n9592_), .B(new_n506_), .Y(new_n9593_));
  NOR2  g09208(.A(new_n9593_), .B(new_n510_), .Y(new_n9594_));
  NOR2  g09209(.A(new_n9594_), .B(new_n516_), .Y(new_n9595_));
  NOR2  g09210(.A(new_n9595_), .B(new_n520_), .Y(new_n9596_));
  NOR2  g09211(.A(new_n9596_), .B(new_n526_), .Y(new_n9597_));
  NOR2  g09212(.A(new_n9597_), .B(new_n530_), .Y(new_n9598_));
  NOR2  g09213(.A(new_n9598_), .B(new_n536_), .Y(new_n9599_));
  NOR2  g09214(.A(new_n9599_), .B(new_n540_), .Y(new_n9600_));
  NOR2  g09215(.A(new_n9600_), .B(new_n546_), .Y(new_n9601_));
  NOR2  g09216(.A(new_n9601_), .B(new_n550_), .Y(new_n9602_));
  NOR2  g09217(.A(new_n9602_), .B(new_n556_), .Y(new_n9603_));
  NOR2  g09218(.A(new_n9603_), .B(new_n560_), .Y(new_n9604_));
  NOR2  g09219(.A(new_n9604_), .B(new_n566_), .Y(new_n9605_));
  NOR2  g09220(.A(new_n9605_), .B(new_n570_), .Y(new_n9606_));
  NOR2  g09221(.A(new_n9606_), .B(new_n576_), .Y(new_n9607_));
  NOR2  g09222(.A(new_n9607_), .B(new_n580_), .Y(new_n9608_));
  NOR2  g09223(.A(new_n9608_), .B(new_n586_), .Y(new_n9609_));
  NOR2  g09224(.A(new_n9609_), .B(new_n590_), .Y(new_n9610_));
  NOR2  g09225(.A(new_n9610_), .B(new_n596_), .Y(new_n9611_));
  NOR2  g09226(.A(new_n9611_), .B(new_n600_), .Y(new_n9612_));
  NOR2  g09227(.A(new_n9612_), .B(new_n606_), .Y(new_n9613_));
  NOR2  g09228(.A(new_n9613_), .B(new_n610_), .Y(new_n9614_));
  NOR2  g09229(.A(new_n9614_), .B(new_n616_), .Y(new_n9615_));
  NOR2  g09230(.A(new_n9615_), .B(new_n620_), .Y(new_n9616_));
  NOR2  g09231(.A(new_n9616_), .B(new_n626_), .Y(new_n9617_));
  NOR2  g09232(.A(new_n9617_), .B(new_n630_), .Y(new_n9618_));
  NOR2  g09233(.A(new_n9618_), .B(new_n636_), .Y(new_n9619_));
  NOR2  g09234(.A(new_n9619_), .B(new_n640_), .Y(new_n9620_));
  NOR2  g09235(.A(new_n9620_), .B(new_n646_), .Y(new_n9621_));
  NOR2  g09236(.A(new_n9621_), .B(new_n650_), .Y(new_n9622_));
  NOR2  g09237(.A(new_n9622_), .B(new_n656_), .Y(new_n9623_));
  NOR2  g09238(.A(new_n9623_), .B(new_n660_), .Y(new_n9624_));
  NOR2  g09239(.A(new_n9624_), .B(new_n666_), .Y(new_n9625_));
  NOR2  g09240(.A(new_n9625_), .B(new_n670_), .Y(new_n9626_));
  NOR2  g09241(.A(new_n9626_), .B(new_n676_), .Y(new_n9627_));
  NOR2  g09242(.A(new_n9627_), .B(new_n680_), .Y(new_n9628_));
  NOR2  g09243(.A(new_n9628_), .B(new_n686_), .Y(new_n9629_));
  NOR2  g09244(.A(new_n9629_), .B(new_n690_), .Y(new_n9630_));
  NOR2  g09245(.A(new_n9630_), .B(new_n696_), .Y(new_n9631_));
  NAND2 g09246(.A(new_n698_), .B(\req[95] ), .Y(new_n9632_));
  NOR2  g09247(.A(new_n9632_), .B(new_n9631_), .Y(\grant[95] ));
  INV   g09248(.A(new_n709_), .Y(new_n9634_));
  NOR2  g09249(.A(new_n1098_), .B(new_n9634_), .Y(new_n9635_));
  NOR2  g09250(.A(new_n9635_), .B(new_n716_), .Y(new_n9636_));
  NOR2  g09251(.A(new_n9636_), .B(new_n720_), .Y(new_n9637_));
  NOR2  g09252(.A(new_n9637_), .B(new_n726_), .Y(new_n9638_));
  NOR2  g09253(.A(new_n9638_), .B(new_n730_), .Y(new_n9639_));
  NOR2  g09254(.A(new_n9639_), .B(new_n736_), .Y(new_n9640_));
  NOR2  g09255(.A(new_n9640_), .B(new_n740_), .Y(new_n9641_));
  NOR2  g09256(.A(new_n9641_), .B(new_n746_), .Y(new_n9642_));
  NOR2  g09257(.A(new_n9642_), .B(new_n750_), .Y(new_n9643_));
  NOR2  g09258(.A(new_n9643_), .B(new_n756_), .Y(new_n9644_));
  NOR2  g09259(.A(new_n9644_), .B(new_n760_), .Y(new_n9645_));
  NOR2  g09260(.A(new_n9645_), .B(new_n766_), .Y(new_n9646_));
  NOR2  g09261(.A(new_n9646_), .B(new_n770_), .Y(new_n9647_));
  NOR2  g09262(.A(new_n9647_), .B(new_n776_), .Y(new_n9648_));
  NOR2  g09263(.A(new_n9648_), .B(new_n780_), .Y(new_n9649_));
  NOR2  g09264(.A(new_n9649_), .B(new_n786_), .Y(new_n9650_));
  NOR2  g09265(.A(new_n9650_), .B(new_n790_), .Y(new_n9651_));
  NOR2  g09266(.A(new_n9651_), .B(new_n796_), .Y(new_n9652_));
  NOR2  g09267(.A(new_n9652_), .B(new_n800_), .Y(new_n9653_));
  NOR2  g09268(.A(new_n9653_), .B(new_n806_), .Y(new_n9654_));
  NOR2  g09269(.A(new_n9654_), .B(new_n1616_), .Y(new_n9655_));
  NOR2  g09270(.A(new_n9655_), .B(new_n1618_), .Y(new_n9656_));
  NOR2  g09271(.A(new_n9656_), .B(new_n1885_), .Y(new_n9657_));
  NOR2  g09272(.A(new_n9657_), .B(new_n820_), .Y(new_n9658_));
  NOR2  g09273(.A(new_n9658_), .B(new_n824_), .Y(new_n9659_));
  NOR2  g09274(.A(new_n9659_), .B(new_n829_), .Y(new_n9660_));
  NOR2  g09275(.A(new_n9660_), .B(new_n833_), .Y(new_n9661_));
  NOR2  g09276(.A(new_n9661_), .B(new_n838_), .Y(new_n9662_));
  NOR2  g09277(.A(new_n9662_), .B(new_n842_), .Y(new_n9663_));
  NOR2  g09278(.A(new_n9663_), .B(new_n847_), .Y(new_n9664_));
  NOR2  g09279(.A(new_n9664_), .B(new_n851_), .Y(new_n9665_));
  NOR2  g09280(.A(new_n9665_), .B(new_n856_), .Y(new_n9666_));
  NOR2  g09281(.A(new_n9666_), .B(new_n860_), .Y(new_n9667_));
  NOR2  g09282(.A(new_n9667_), .B(new_n865_), .Y(new_n9668_));
  NOR2  g09283(.A(new_n9668_), .B(new_n869_), .Y(new_n9669_));
  NOR2  g09284(.A(new_n9669_), .B(new_n874_), .Y(new_n9670_));
  NOR2  g09285(.A(new_n9670_), .B(new_n878_), .Y(new_n9671_));
  NOR2  g09286(.A(new_n9671_), .B(new_n883_), .Y(new_n9672_));
  NOR2  g09287(.A(new_n9672_), .B(new_n887_), .Y(new_n9673_));
  NOR2  g09288(.A(new_n9673_), .B(new_n892_), .Y(new_n9674_));
  NOR2  g09289(.A(new_n9674_), .B(new_n896_), .Y(new_n9675_));
  NOR2  g09290(.A(new_n9675_), .B(new_n901_), .Y(new_n9676_));
  NOR2  g09291(.A(new_n9676_), .B(new_n905_), .Y(new_n9677_));
  NOR2  g09292(.A(new_n9677_), .B(new_n910_), .Y(new_n9678_));
  NOR2  g09293(.A(new_n9678_), .B(new_n914_), .Y(new_n9679_));
  NOR2  g09294(.A(new_n9679_), .B(new_n919_), .Y(new_n9680_));
  NOR2  g09295(.A(new_n9680_), .B(new_n923_), .Y(new_n9681_));
  NOR2  g09296(.A(new_n9681_), .B(new_n928_), .Y(new_n9682_));
  NOR2  g09297(.A(new_n9682_), .B(new_n932_), .Y(new_n9683_));
  NOR2  g09298(.A(new_n9683_), .B(new_n937_), .Y(new_n9684_));
  NOR2  g09299(.A(new_n9684_), .B(new_n941_), .Y(new_n9685_));
  NOR2  g09300(.A(new_n9685_), .B(new_n946_), .Y(new_n9686_));
  NOR2  g09301(.A(new_n9686_), .B(new_n950_), .Y(new_n9687_));
  NOR2  g09302(.A(new_n9687_), .B(new_n955_), .Y(new_n9688_));
  NOR2  g09303(.A(new_n9688_), .B(new_n959_), .Y(new_n9689_));
  NOR2  g09304(.A(new_n9689_), .B(new_n964_), .Y(new_n9690_));
  NOR2  g09305(.A(new_n9690_), .B(new_n968_), .Y(new_n9691_));
  NOR2  g09306(.A(new_n9691_), .B(new_n973_), .Y(new_n9692_));
  NOR2  g09307(.A(new_n9692_), .B(new_n977_), .Y(new_n9693_));
  NOR2  g09308(.A(new_n9693_), .B(new_n982_), .Y(new_n9694_));
  NOR2  g09309(.A(new_n9694_), .B(new_n986_), .Y(new_n9695_));
  NOR2  g09310(.A(new_n9695_), .B(new_n991_), .Y(new_n9696_));
  NOR2  g09311(.A(new_n9696_), .B(new_n995_), .Y(new_n9697_));
  NOR2  g09312(.A(new_n9697_), .B(new_n1000_), .Y(new_n9698_));
  NOR2  g09313(.A(new_n9698_), .B(new_n1004_), .Y(new_n9699_));
  NOR2  g09314(.A(new_n9699_), .B(new_n1009_), .Y(new_n9700_));
  NOR2  g09315(.A(new_n9700_), .B(new_n1013_), .Y(new_n9701_));
  NOR2  g09316(.A(new_n9701_), .B(new_n1018_), .Y(new_n9702_));
  NOR2  g09317(.A(new_n9702_), .B(new_n1022_), .Y(new_n9703_));
  NOR2  g09318(.A(new_n9703_), .B(new_n1027_), .Y(new_n9704_));
  NOR2  g09319(.A(new_n9704_), .B(new_n1031_), .Y(new_n9705_));
  NOR2  g09320(.A(new_n9705_), .B(new_n1036_), .Y(new_n9706_));
  NOR2  g09321(.A(new_n9706_), .B(new_n1040_), .Y(new_n9707_));
  NOR2  g09322(.A(new_n9707_), .B(new_n1045_), .Y(new_n9708_));
  NOR2  g09323(.A(new_n9708_), .B(new_n1049_), .Y(new_n9709_));
  NOR2  g09324(.A(new_n9709_), .B(new_n1054_), .Y(new_n9710_));
  NOR2  g09325(.A(new_n9710_), .B(new_n1058_), .Y(new_n9711_));
  NOR2  g09326(.A(new_n9711_), .B(new_n1063_), .Y(new_n9712_));
  NOR2  g09327(.A(new_n9712_), .B(new_n1067_), .Y(new_n9713_));
  NOR2  g09328(.A(new_n9713_), .B(new_n1072_), .Y(new_n9714_));
  NOR2  g09329(.A(new_n9714_), .B(new_n1076_), .Y(new_n9715_));
  NOR2  g09330(.A(new_n9715_), .B(new_n1081_), .Y(new_n9716_));
  NOR2  g09331(.A(new_n9716_), .B(new_n1085_), .Y(new_n9717_));
  NOR2  g09332(.A(new_n9717_), .B(new_n1090_), .Y(new_n9718_));
  NAND2 g09333(.A(new_n1092_), .B(\req[96] ), .Y(new_n9719_));
  NOR2  g09334(.A(new_n9719_), .B(new_n9718_), .Y(\grant[96] ));
  INV   g09335(.A(new_n1102_), .Y(new_n9721_));
  NOR2  g09336(.A(new_n1446_), .B(new_n9721_), .Y(new_n9722_));
  NOR2  g09337(.A(new_n9722_), .B(new_n1108_), .Y(new_n9723_));
  NOR2  g09338(.A(new_n9723_), .B(new_n1112_), .Y(new_n9724_));
  NOR2  g09339(.A(new_n9724_), .B(new_n1117_), .Y(new_n9725_));
  NOR2  g09340(.A(new_n9725_), .B(new_n1121_), .Y(new_n9726_));
  NOR2  g09341(.A(new_n9726_), .B(new_n1126_), .Y(new_n9727_));
  NOR2  g09342(.A(new_n9727_), .B(new_n1130_), .Y(new_n9728_));
  NOR2  g09343(.A(new_n9728_), .B(new_n1135_), .Y(new_n9729_));
  NOR2  g09344(.A(new_n9729_), .B(new_n1139_), .Y(new_n9730_));
  NOR2  g09345(.A(new_n9730_), .B(new_n1144_), .Y(new_n9731_));
  NOR2  g09346(.A(new_n9731_), .B(new_n1148_), .Y(new_n9732_));
  NOR2  g09347(.A(new_n9732_), .B(new_n1153_), .Y(new_n9733_));
  NOR2  g09348(.A(new_n9733_), .B(new_n1157_), .Y(new_n9734_));
  NOR2  g09349(.A(new_n9734_), .B(new_n1162_), .Y(new_n9735_));
  NOR2  g09350(.A(new_n9735_), .B(new_n1166_), .Y(new_n9736_));
  NOR2  g09351(.A(new_n9736_), .B(new_n1171_), .Y(new_n9737_));
  NOR2  g09352(.A(new_n9737_), .B(new_n1175_), .Y(new_n9738_));
  NOR2  g09353(.A(new_n9738_), .B(new_n1180_), .Y(new_n9739_));
  NOR2  g09354(.A(new_n9739_), .B(new_n1184_), .Y(new_n9740_));
  NOR2  g09355(.A(new_n9740_), .B(new_n1189_), .Y(new_n9741_));
  NOR2  g09356(.A(new_n9741_), .B(new_n1707_), .Y(new_n9742_));
  NOR2  g09357(.A(new_n9742_), .B(new_n1709_), .Y(new_n9743_));
  NOR2  g09358(.A(new_n9743_), .B(new_n1973_), .Y(new_n9744_));
  NOR2  g09359(.A(new_n9744_), .B(new_n1199_), .Y(new_n9745_));
  NOR2  g09360(.A(new_n9745_), .B(new_n1203_), .Y(new_n9746_));
  NOR2  g09361(.A(new_n9746_), .B(new_n1207_), .Y(new_n9747_));
  NOR2  g09362(.A(new_n9747_), .B(new_n1211_), .Y(new_n9748_));
  NOR2  g09363(.A(new_n9748_), .B(new_n1215_), .Y(new_n9749_));
  NOR2  g09364(.A(new_n9749_), .B(new_n1219_), .Y(new_n9750_));
  NOR2  g09365(.A(new_n9750_), .B(new_n1223_), .Y(new_n9751_));
  NOR2  g09366(.A(new_n9751_), .B(new_n1227_), .Y(new_n9752_));
  NOR2  g09367(.A(new_n9752_), .B(new_n1231_), .Y(new_n9753_));
  NOR2  g09368(.A(new_n9753_), .B(new_n1235_), .Y(new_n9754_));
  NOR2  g09369(.A(new_n9754_), .B(new_n1239_), .Y(new_n9755_));
  NOR2  g09370(.A(new_n9755_), .B(new_n1243_), .Y(new_n9756_));
  NOR2  g09371(.A(new_n9756_), .B(new_n1247_), .Y(new_n9757_));
  NOR2  g09372(.A(new_n9757_), .B(new_n1251_), .Y(new_n9758_));
  NOR2  g09373(.A(new_n9758_), .B(new_n1255_), .Y(new_n9759_));
  NOR2  g09374(.A(new_n9759_), .B(new_n1259_), .Y(new_n9760_));
  NOR2  g09375(.A(new_n9760_), .B(new_n1263_), .Y(new_n9761_));
  NOR2  g09376(.A(new_n9761_), .B(new_n1267_), .Y(new_n9762_));
  NOR2  g09377(.A(new_n9762_), .B(new_n1271_), .Y(new_n9763_));
  NOR2  g09378(.A(new_n9763_), .B(new_n1275_), .Y(new_n9764_));
  NOR2  g09379(.A(new_n9764_), .B(new_n1279_), .Y(new_n9765_));
  NOR2  g09380(.A(new_n9765_), .B(new_n1283_), .Y(new_n9766_));
  NOR2  g09381(.A(new_n9766_), .B(new_n1287_), .Y(new_n9767_));
  NOR2  g09382(.A(new_n9767_), .B(new_n1291_), .Y(new_n9768_));
  NOR2  g09383(.A(new_n9768_), .B(new_n1295_), .Y(new_n9769_));
  NOR2  g09384(.A(new_n9769_), .B(new_n1299_), .Y(new_n9770_));
  NOR2  g09385(.A(new_n9770_), .B(new_n1303_), .Y(new_n9771_));
  NOR2  g09386(.A(new_n9771_), .B(new_n1307_), .Y(new_n9772_));
  NOR2  g09387(.A(new_n9772_), .B(new_n1311_), .Y(new_n9773_));
  NOR2  g09388(.A(new_n9773_), .B(new_n1315_), .Y(new_n9774_));
  NOR2  g09389(.A(new_n9774_), .B(new_n1319_), .Y(new_n9775_));
  NOR2  g09390(.A(new_n9775_), .B(new_n1323_), .Y(new_n9776_));
  NOR2  g09391(.A(new_n9776_), .B(new_n1327_), .Y(new_n9777_));
  NOR2  g09392(.A(new_n9777_), .B(new_n1331_), .Y(new_n9778_));
  NOR2  g09393(.A(new_n9778_), .B(new_n1335_), .Y(new_n9779_));
  NOR2  g09394(.A(new_n9779_), .B(new_n1339_), .Y(new_n9780_));
  NOR2  g09395(.A(new_n9780_), .B(new_n1343_), .Y(new_n9781_));
  NOR2  g09396(.A(new_n9781_), .B(new_n1347_), .Y(new_n9782_));
  NOR2  g09397(.A(new_n9782_), .B(new_n1351_), .Y(new_n9783_));
  NOR2  g09398(.A(new_n9783_), .B(new_n1355_), .Y(new_n9784_));
  NOR2  g09399(.A(new_n9784_), .B(new_n1359_), .Y(new_n9785_));
  NOR2  g09400(.A(new_n9785_), .B(new_n1363_), .Y(new_n9786_));
  NOR2  g09401(.A(new_n9786_), .B(new_n1367_), .Y(new_n9787_));
  NOR2  g09402(.A(new_n9787_), .B(new_n1371_), .Y(new_n9788_));
  NOR2  g09403(.A(new_n9788_), .B(new_n1375_), .Y(new_n9789_));
  NOR2  g09404(.A(new_n9789_), .B(new_n1379_), .Y(new_n9790_));
  NOR2  g09405(.A(new_n9790_), .B(new_n1383_), .Y(new_n9791_));
  NOR2  g09406(.A(new_n9791_), .B(new_n1387_), .Y(new_n9792_));
  NOR2  g09407(.A(new_n9792_), .B(new_n1391_), .Y(new_n9793_));
  NOR2  g09408(.A(new_n9793_), .B(new_n1395_), .Y(new_n9794_));
  NOR2  g09409(.A(new_n9794_), .B(new_n1399_), .Y(new_n9795_));
  NOR2  g09410(.A(new_n9795_), .B(new_n1403_), .Y(new_n9796_));
  NOR2  g09411(.A(new_n9796_), .B(new_n1407_), .Y(new_n9797_));
  NOR2  g09412(.A(new_n9797_), .B(new_n1411_), .Y(new_n9798_));
  NOR2  g09413(.A(new_n9798_), .B(new_n1415_), .Y(new_n9799_));
  NOR2  g09414(.A(new_n9799_), .B(new_n1419_), .Y(new_n9800_));
  NOR2  g09415(.A(new_n9800_), .B(new_n1423_), .Y(new_n9801_));
  NOR2  g09416(.A(new_n9801_), .B(new_n1427_), .Y(new_n9802_));
  NOR2  g09417(.A(new_n9802_), .B(new_n1431_), .Y(new_n9803_));
  NOR2  g09418(.A(new_n9803_), .B(new_n1435_), .Y(new_n9804_));
  NOR2  g09419(.A(new_n9804_), .B(new_n1439_), .Y(new_n9805_));
  NAND2 g09420(.A(new_n1441_), .B(\req[97] ), .Y(new_n9806_));
  NOR2  g09421(.A(new_n9806_), .B(new_n9805_), .Y(\grant[97] ));
  INV   g09422(.A(new_n1450_), .Y(new_n9808_));
  NOR2  g09423(.A(new_n9808_), .B(new_n715_), .Y(new_n9809_));
  NOR2  g09424(.A(new_n9809_), .B(new_n1455_), .Y(new_n9810_));
  NOR2  g09425(.A(new_n9810_), .B(new_n1459_), .Y(new_n9811_));
  NOR2  g09426(.A(new_n9811_), .B(new_n1463_), .Y(new_n9812_));
  NOR2  g09427(.A(new_n9812_), .B(new_n1467_), .Y(new_n9813_));
  NOR2  g09428(.A(new_n9813_), .B(new_n1471_), .Y(new_n9814_));
  NOR2  g09429(.A(new_n9814_), .B(new_n1475_), .Y(new_n9815_));
  NOR2  g09430(.A(new_n9815_), .B(new_n1479_), .Y(new_n9816_));
  NOR2  g09431(.A(new_n9816_), .B(new_n1483_), .Y(new_n9817_));
  NOR2  g09432(.A(new_n9817_), .B(new_n1487_), .Y(new_n9818_));
  NOR2  g09433(.A(new_n9818_), .B(new_n1491_), .Y(new_n9819_));
  NOR2  g09434(.A(new_n9819_), .B(new_n1495_), .Y(new_n9820_));
  NOR2  g09435(.A(new_n9820_), .B(new_n1499_), .Y(new_n9821_));
  NOR2  g09436(.A(new_n9821_), .B(new_n1503_), .Y(new_n9822_));
  NOR2  g09437(.A(new_n9822_), .B(new_n1507_), .Y(new_n9823_));
  NOR2  g09438(.A(new_n9823_), .B(new_n1511_), .Y(new_n9824_));
  NOR2  g09439(.A(new_n9824_), .B(new_n1515_), .Y(new_n9825_));
  NOR2  g09440(.A(new_n9825_), .B(new_n1519_), .Y(new_n9826_));
  NOR2  g09441(.A(new_n9826_), .B(new_n1523_), .Y(new_n9827_));
  NOR2  g09442(.A(new_n9827_), .B(new_n1527_), .Y(new_n9828_));
  NOR2  g09443(.A(new_n9828_), .B(new_n1797_), .Y(new_n9829_));
  NOR2  g09444(.A(new_n9829_), .B(new_n396_), .Y(new_n9830_));
  NOR2  g09445(.A(new_n9830_), .B(new_n400_), .Y(new_n9831_));
  NOR2  g09446(.A(new_n9831_), .B(new_n406_), .Y(new_n9832_));
  NOR2  g09447(.A(new_n9832_), .B(new_n410_), .Y(new_n9833_));
  NOR2  g09448(.A(new_n9833_), .B(new_n416_), .Y(new_n9834_));
  NOR2  g09449(.A(new_n9834_), .B(new_n420_), .Y(new_n9835_));
  NOR2  g09450(.A(new_n9835_), .B(new_n426_), .Y(new_n9836_));
  NOR2  g09451(.A(new_n9836_), .B(new_n430_), .Y(new_n9837_));
  NOR2  g09452(.A(new_n9837_), .B(new_n436_), .Y(new_n9838_));
  NOR2  g09453(.A(new_n9838_), .B(new_n440_), .Y(new_n9839_));
  NOR2  g09454(.A(new_n9839_), .B(new_n446_), .Y(new_n9840_));
  NOR2  g09455(.A(new_n9840_), .B(new_n450_), .Y(new_n9841_));
  NOR2  g09456(.A(new_n9841_), .B(new_n456_), .Y(new_n9842_));
  NOR2  g09457(.A(new_n9842_), .B(new_n460_), .Y(new_n9843_));
  NOR2  g09458(.A(new_n9843_), .B(new_n466_), .Y(new_n9844_));
  NOR2  g09459(.A(new_n9844_), .B(new_n470_), .Y(new_n9845_));
  NOR2  g09460(.A(new_n9845_), .B(new_n476_), .Y(new_n9846_));
  NOR2  g09461(.A(new_n9846_), .B(new_n480_), .Y(new_n9847_));
  NOR2  g09462(.A(new_n9847_), .B(new_n486_), .Y(new_n9848_));
  NOR2  g09463(.A(new_n9848_), .B(new_n490_), .Y(new_n9849_));
  NOR2  g09464(.A(new_n9849_), .B(new_n496_), .Y(new_n9850_));
  NOR2  g09465(.A(new_n9850_), .B(new_n500_), .Y(new_n9851_));
  NOR2  g09466(.A(new_n9851_), .B(new_n506_), .Y(new_n9852_));
  NOR2  g09467(.A(new_n9852_), .B(new_n510_), .Y(new_n9853_));
  NOR2  g09468(.A(new_n9853_), .B(new_n516_), .Y(new_n9854_));
  NOR2  g09469(.A(new_n9854_), .B(new_n520_), .Y(new_n9855_));
  NOR2  g09470(.A(new_n9855_), .B(new_n526_), .Y(new_n9856_));
  NOR2  g09471(.A(new_n9856_), .B(new_n530_), .Y(new_n9857_));
  NOR2  g09472(.A(new_n9857_), .B(new_n536_), .Y(new_n9858_));
  NOR2  g09473(.A(new_n9858_), .B(new_n540_), .Y(new_n9859_));
  NOR2  g09474(.A(new_n9859_), .B(new_n546_), .Y(new_n9860_));
  NOR2  g09475(.A(new_n9860_), .B(new_n550_), .Y(new_n9861_));
  NOR2  g09476(.A(new_n9861_), .B(new_n556_), .Y(new_n9862_));
  NOR2  g09477(.A(new_n9862_), .B(new_n560_), .Y(new_n9863_));
  NOR2  g09478(.A(new_n9863_), .B(new_n566_), .Y(new_n9864_));
  NOR2  g09479(.A(new_n9864_), .B(new_n570_), .Y(new_n9865_));
  NOR2  g09480(.A(new_n9865_), .B(new_n576_), .Y(new_n9866_));
  NOR2  g09481(.A(new_n9866_), .B(new_n580_), .Y(new_n9867_));
  NOR2  g09482(.A(new_n9867_), .B(new_n586_), .Y(new_n9868_));
  NOR2  g09483(.A(new_n9868_), .B(new_n590_), .Y(new_n9869_));
  NOR2  g09484(.A(new_n9869_), .B(new_n596_), .Y(new_n9870_));
  NOR2  g09485(.A(new_n9870_), .B(new_n600_), .Y(new_n9871_));
  NOR2  g09486(.A(new_n9871_), .B(new_n606_), .Y(new_n9872_));
  NOR2  g09487(.A(new_n9872_), .B(new_n610_), .Y(new_n9873_));
  NOR2  g09488(.A(new_n9873_), .B(new_n616_), .Y(new_n9874_));
  NOR2  g09489(.A(new_n9874_), .B(new_n620_), .Y(new_n9875_));
  NOR2  g09490(.A(new_n9875_), .B(new_n626_), .Y(new_n9876_));
  NOR2  g09491(.A(new_n9876_), .B(new_n630_), .Y(new_n9877_));
  NOR2  g09492(.A(new_n9877_), .B(new_n636_), .Y(new_n9878_));
  NOR2  g09493(.A(new_n9878_), .B(new_n640_), .Y(new_n9879_));
  NOR2  g09494(.A(new_n9879_), .B(new_n646_), .Y(new_n9880_));
  NOR2  g09495(.A(new_n9880_), .B(new_n650_), .Y(new_n9881_));
  NOR2  g09496(.A(new_n9881_), .B(new_n656_), .Y(new_n9882_));
  NOR2  g09497(.A(new_n9882_), .B(new_n660_), .Y(new_n9883_));
  NOR2  g09498(.A(new_n9883_), .B(new_n666_), .Y(new_n9884_));
  NOR2  g09499(.A(new_n9884_), .B(new_n670_), .Y(new_n9885_));
  NOR2  g09500(.A(new_n9885_), .B(new_n676_), .Y(new_n9886_));
  NOR2  g09501(.A(new_n9886_), .B(new_n680_), .Y(new_n9887_));
  NOR2  g09502(.A(new_n9887_), .B(new_n686_), .Y(new_n9888_));
  NOR2  g09503(.A(new_n9888_), .B(new_n690_), .Y(new_n9889_));
  NOR2  g09504(.A(new_n9889_), .B(new_n696_), .Y(new_n9890_));
  NOR2  g09505(.A(new_n9890_), .B(new_n700_), .Y(new_n9891_));
  NOR2  g09506(.A(new_n9891_), .B(new_n706_), .Y(new_n9892_));
  NAND2 g09507(.A(new_n708_), .B(\req[98] ), .Y(new_n9893_));
  NOR2  g09508(.A(new_n9893_), .B(new_n9892_), .Y(\grant[98] ));
  INV   g09509(.A(new_n719_), .Y(new_n9895_));
  NOR2  g09510(.A(new_n1107_), .B(new_n9895_), .Y(new_n9896_));
  NOR2  g09511(.A(new_n9896_), .B(new_n726_), .Y(new_n9897_));
  NOR2  g09512(.A(new_n9897_), .B(new_n730_), .Y(new_n9898_));
  NOR2  g09513(.A(new_n9898_), .B(new_n736_), .Y(new_n9899_));
  NOR2  g09514(.A(new_n9899_), .B(new_n740_), .Y(new_n9900_));
  NOR2  g09515(.A(new_n9900_), .B(new_n746_), .Y(new_n9901_));
  NOR2  g09516(.A(new_n9901_), .B(new_n750_), .Y(new_n9902_));
  NOR2  g09517(.A(new_n9902_), .B(new_n756_), .Y(new_n9903_));
  NOR2  g09518(.A(new_n9903_), .B(new_n760_), .Y(new_n9904_));
  NOR2  g09519(.A(new_n9904_), .B(new_n766_), .Y(new_n9905_));
  NOR2  g09520(.A(new_n9905_), .B(new_n770_), .Y(new_n9906_));
  NOR2  g09521(.A(new_n9906_), .B(new_n776_), .Y(new_n9907_));
  NOR2  g09522(.A(new_n9907_), .B(new_n780_), .Y(new_n9908_));
  NOR2  g09523(.A(new_n9908_), .B(new_n786_), .Y(new_n9909_));
  NOR2  g09524(.A(new_n9909_), .B(new_n790_), .Y(new_n9910_));
  NOR2  g09525(.A(new_n9910_), .B(new_n796_), .Y(new_n9911_));
  NOR2  g09526(.A(new_n9911_), .B(new_n800_), .Y(new_n9912_));
  NOR2  g09527(.A(new_n9912_), .B(new_n806_), .Y(new_n9913_));
  NOR2  g09528(.A(new_n9913_), .B(new_n1616_), .Y(new_n9914_));
  NOR2  g09529(.A(new_n9914_), .B(new_n1618_), .Y(new_n9915_));
  NOR2  g09530(.A(new_n9915_), .B(new_n1885_), .Y(new_n9916_));
  NOR2  g09531(.A(new_n9916_), .B(new_n820_), .Y(new_n9917_));
  NOR2  g09532(.A(new_n9917_), .B(new_n824_), .Y(new_n9918_));
  NOR2  g09533(.A(new_n9918_), .B(new_n829_), .Y(new_n9919_));
  NOR2  g09534(.A(new_n9919_), .B(new_n833_), .Y(new_n9920_));
  NOR2  g09535(.A(new_n9920_), .B(new_n838_), .Y(new_n9921_));
  NOR2  g09536(.A(new_n9921_), .B(new_n842_), .Y(new_n9922_));
  NOR2  g09537(.A(new_n9922_), .B(new_n847_), .Y(new_n9923_));
  NOR2  g09538(.A(new_n9923_), .B(new_n851_), .Y(new_n9924_));
  NOR2  g09539(.A(new_n9924_), .B(new_n856_), .Y(new_n9925_));
  NOR2  g09540(.A(new_n9925_), .B(new_n860_), .Y(new_n9926_));
  NOR2  g09541(.A(new_n9926_), .B(new_n865_), .Y(new_n9927_));
  NOR2  g09542(.A(new_n9927_), .B(new_n869_), .Y(new_n9928_));
  NOR2  g09543(.A(new_n9928_), .B(new_n874_), .Y(new_n9929_));
  NOR2  g09544(.A(new_n9929_), .B(new_n878_), .Y(new_n9930_));
  NOR2  g09545(.A(new_n9930_), .B(new_n883_), .Y(new_n9931_));
  NOR2  g09546(.A(new_n9931_), .B(new_n887_), .Y(new_n9932_));
  NOR2  g09547(.A(new_n9932_), .B(new_n892_), .Y(new_n9933_));
  NOR2  g09548(.A(new_n9933_), .B(new_n896_), .Y(new_n9934_));
  NOR2  g09549(.A(new_n9934_), .B(new_n901_), .Y(new_n9935_));
  NOR2  g09550(.A(new_n9935_), .B(new_n905_), .Y(new_n9936_));
  NOR2  g09551(.A(new_n9936_), .B(new_n910_), .Y(new_n9937_));
  NOR2  g09552(.A(new_n9937_), .B(new_n914_), .Y(new_n9938_));
  NOR2  g09553(.A(new_n9938_), .B(new_n919_), .Y(new_n9939_));
  NOR2  g09554(.A(new_n9939_), .B(new_n923_), .Y(new_n9940_));
  NOR2  g09555(.A(new_n9940_), .B(new_n928_), .Y(new_n9941_));
  NOR2  g09556(.A(new_n9941_), .B(new_n932_), .Y(new_n9942_));
  NOR2  g09557(.A(new_n9942_), .B(new_n937_), .Y(new_n9943_));
  NOR2  g09558(.A(new_n9943_), .B(new_n941_), .Y(new_n9944_));
  NOR2  g09559(.A(new_n9944_), .B(new_n946_), .Y(new_n9945_));
  NOR2  g09560(.A(new_n9945_), .B(new_n950_), .Y(new_n9946_));
  NOR2  g09561(.A(new_n9946_), .B(new_n955_), .Y(new_n9947_));
  NOR2  g09562(.A(new_n9947_), .B(new_n959_), .Y(new_n9948_));
  NOR2  g09563(.A(new_n9948_), .B(new_n964_), .Y(new_n9949_));
  NOR2  g09564(.A(new_n9949_), .B(new_n968_), .Y(new_n9950_));
  NOR2  g09565(.A(new_n9950_), .B(new_n973_), .Y(new_n9951_));
  NOR2  g09566(.A(new_n9951_), .B(new_n977_), .Y(new_n9952_));
  NOR2  g09567(.A(new_n9952_), .B(new_n982_), .Y(new_n9953_));
  NOR2  g09568(.A(new_n9953_), .B(new_n986_), .Y(new_n9954_));
  NOR2  g09569(.A(new_n9954_), .B(new_n991_), .Y(new_n9955_));
  NOR2  g09570(.A(new_n9955_), .B(new_n995_), .Y(new_n9956_));
  NOR2  g09571(.A(new_n9956_), .B(new_n1000_), .Y(new_n9957_));
  NOR2  g09572(.A(new_n9957_), .B(new_n1004_), .Y(new_n9958_));
  NOR2  g09573(.A(new_n9958_), .B(new_n1009_), .Y(new_n9959_));
  NOR2  g09574(.A(new_n9959_), .B(new_n1013_), .Y(new_n9960_));
  NOR2  g09575(.A(new_n9960_), .B(new_n1018_), .Y(new_n9961_));
  NOR2  g09576(.A(new_n9961_), .B(new_n1022_), .Y(new_n9962_));
  NOR2  g09577(.A(new_n9962_), .B(new_n1027_), .Y(new_n9963_));
  NOR2  g09578(.A(new_n9963_), .B(new_n1031_), .Y(new_n9964_));
  NOR2  g09579(.A(new_n9964_), .B(new_n1036_), .Y(new_n9965_));
  NOR2  g09580(.A(new_n9965_), .B(new_n1040_), .Y(new_n9966_));
  NOR2  g09581(.A(new_n9966_), .B(new_n1045_), .Y(new_n9967_));
  NOR2  g09582(.A(new_n9967_), .B(new_n1049_), .Y(new_n9968_));
  NOR2  g09583(.A(new_n9968_), .B(new_n1054_), .Y(new_n9969_));
  NOR2  g09584(.A(new_n9969_), .B(new_n1058_), .Y(new_n9970_));
  NOR2  g09585(.A(new_n9970_), .B(new_n1063_), .Y(new_n9971_));
  NOR2  g09586(.A(new_n9971_), .B(new_n1067_), .Y(new_n9972_));
  NOR2  g09587(.A(new_n9972_), .B(new_n1072_), .Y(new_n9973_));
  NOR2  g09588(.A(new_n9973_), .B(new_n1076_), .Y(new_n9974_));
  NOR2  g09589(.A(new_n9974_), .B(new_n1081_), .Y(new_n9975_));
  NOR2  g09590(.A(new_n9975_), .B(new_n1085_), .Y(new_n9976_));
  NOR2  g09591(.A(new_n9976_), .B(new_n1090_), .Y(new_n9977_));
  NOR2  g09592(.A(new_n9977_), .B(new_n1094_), .Y(new_n9978_));
  NOR2  g09593(.A(new_n9978_), .B(new_n1099_), .Y(new_n9979_));
  NAND2 g09594(.A(new_n1101_), .B(\req[99] ), .Y(new_n9980_));
  NOR2  g09595(.A(new_n9980_), .B(new_n9979_), .Y(\grant[99] ));
  INV   g09596(.A(new_n1111_), .Y(new_n9982_));
  NOR2  g09597(.A(new_n1454_), .B(new_n9982_), .Y(new_n9983_));
  NOR2  g09598(.A(new_n9983_), .B(new_n1117_), .Y(new_n9984_));
  NOR2  g09599(.A(new_n9984_), .B(new_n1121_), .Y(new_n9985_));
  NOR2  g09600(.A(new_n9985_), .B(new_n1126_), .Y(new_n9986_));
  NOR2  g09601(.A(new_n9986_), .B(new_n1130_), .Y(new_n9987_));
  NOR2  g09602(.A(new_n9987_), .B(new_n1135_), .Y(new_n9988_));
  NOR2  g09603(.A(new_n9988_), .B(new_n1139_), .Y(new_n9989_));
  NOR2  g09604(.A(new_n9989_), .B(new_n1144_), .Y(new_n9990_));
  NOR2  g09605(.A(new_n9990_), .B(new_n1148_), .Y(new_n9991_));
  NOR2  g09606(.A(new_n9991_), .B(new_n1153_), .Y(new_n9992_));
  NOR2  g09607(.A(new_n9992_), .B(new_n1157_), .Y(new_n9993_));
  NOR2  g09608(.A(new_n9993_), .B(new_n1162_), .Y(new_n9994_));
  NOR2  g09609(.A(new_n9994_), .B(new_n1166_), .Y(new_n9995_));
  NOR2  g09610(.A(new_n9995_), .B(new_n1171_), .Y(new_n9996_));
  NOR2  g09611(.A(new_n9996_), .B(new_n1175_), .Y(new_n9997_));
  NOR2  g09612(.A(new_n9997_), .B(new_n1180_), .Y(new_n9998_));
  NOR2  g09613(.A(new_n9998_), .B(new_n1184_), .Y(new_n9999_));
  NOR2  g09614(.A(new_n9999_), .B(new_n1189_), .Y(new_n10000_));
  NOR2  g09615(.A(new_n10000_), .B(new_n1707_), .Y(new_n10001_));
  NOR2  g09616(.A(new_n10001_), .B(new_n1709_), .Y(new_n10002_));
  NOR2  g09617(.A(new_n10002_), .B(new_n1973_), .Y(new_n10003_));
  NOR2  g09618(.A(new_n10003_), .B(new_n1199_), .Y(new_n10004_));
  NOR2  g09619(.A(new_n10004_), .B(new_n1203_), .Y(new_n10005_));
  NOR2  g09620(.A(new_n10005_), .B(new_n1207_), .Y(new_n10006_));
  NOR2  g09621(.A(new_n10006_), .B(new_n1211_), .Y(new_n10007_));
  NOR2  g09622(.A(new_n10007_), .B(new_n1215_), .Y(new_n10008_));
  NOR2  g09623(.A(new_n10008_), .B(new_n1219_), .Y(new_n10009_));
  NOR2  g09624(.A(new_n10009_), .B(new_n1223_), .Y(new_n10010_));
  NOR2  g09625(.A(new_n10010_), .B(new_n1227_), .Y(new_n10011_));
  NOR2  g09626(.A(new_n10011_), .B(new_n1231_), .Y(new_n10012_));
  NOR2  g09627(.A(new_n10012_), .B(new_n1235_), .Y(new_n10013_));
  NOR2  g09628(.A(new_n10013_), .B(new_n1239_), .Y(new_n10014_));
  NOR2  g09629(.A(new_n10014_), .B(new_n1243_), .Y(new_n10015_));
  NOR2  g09630(.A(new_n10015_), .B(new_n1247_), .Y(new_n10016_));
  NOR2  g09631(.A(new_n10016_), .B(new_n1251_), .Y(new_n10017_));
  NOR2  g09632(.A(new_n10017_), .B(new_n1255_), .Y(new_n10018_));
  NOR2  g09633(.A(new_n10018_), .B(new_n1259_), .Y(new_n10019_));
  NOR2  g09634(.A(new_n10019_), .B(new_n1263_), .Y(new_n10020_));
  NOR2  g09635(.A(new_n10020_), .B(new_n1267_), .Y(new_n10021_));
  NOR2  g09636(.A(new_n10021_), .B(new_n1271_), .Y(new_n10022_));
  NOR2  g09637(.A(new_n10022_), .B(new_n1275_), .Y(new_n10023_));
  NOR2  g09638(.A(new_n10023_), .B(new_n1279_), .Y(new_n10024_));
  NOR2  g09639(.A(new_n10024_), .B(new_n1283_), .Y(new_n10025_));
  NOR2  g09640(.A(new_n10025_), .B(new_n1287_), .Y(new_n10026_));
  NOR2  g09641(.A(new_n10026_), .B(new_n1291_), .Y(new_n10027_));
  NOR2  g09642(.A(new_n10027_), .B(new_n1295_), .Y(new_n10028_));
  NOR2  g09643(.A(new_n10028_), .B(new_n1299_), .Y(new_n10029_));
  NOR2  g09644(.A(new_n10029_), .B(new_n1303_), .Y(new_n10030_));
  NOR2  g09645(.A(new_n10030_), .B(new_n1307_), .Y(new_n10031_));
  NOR2  g09646(.A(new_n10031_), .B(new_n1311_), .Y(new_n10032_));
  NOR2  g09647(.A(new_n10032_), .B(new_n1315_), .Y(new_n10033_));
  NOR2  g09648(.A(new_n10033_), .B(new_n1319_), .Y(new_n10034_));
  NOR2  g09649(.A(new_n10034_), .B(new_n1323_), .Y(new_n10035_));
  NOR2  g09650(.A(new_n10035_), .B(new_n1327_), .Y(new_n10036_));
  NOR2  g09651(.A(new_n10036_), .B(new_n1331_), .Y(new_n10037_));
  NOR2  g09652(.A(new_n10037_), .B(new_n1335_), .Y(new_n10038_));
  NOR2  g09653(.A(new_n10038_), .B(new_n1339_), .Y(new_n10039_));
  NOR2  g09654(.A(new_n10039_), .B(new_n1343_), .Y(new_n10040_));
  NOR2  g09655(.A(new_n10040_), .B(new_n1347_), .Y(new_n10041_));
  NOR2  g09656(.A(new_n10041_), .B(new_n1351_), .Y(new_n10042_));
  NOR2  g09657(.A(new_n10042_), .B(new_n1355_), .Y(new_n10043_));
  NOR2  g09658(.A(new_n10043_), .B(new_n1359_), .Y(new_n10044_));
  NOR2  g09659(.A(new_n10044_), .B(new_n1363_), .Y(new_n10045_));
  NOR2  g09660(.A(new_n10045_), .B(new_n1367_), .Y(new_n10046_));
  NOR2  g09661(.A(new_n10046_), .B(new_n1371_), .Y(new_n10047_));
  NOR2  g09662(.A(new_n10047_), .B(new_n1375_), .Y(new_n10048_));
  NOR2  g09663(.A(new_n10048_), .B(new_n1379_), .Y(new_n10049_));
  NOR2  g09664(.A(new_n10049_), .B(new_n1383_), .Y(new_n10050_));
  NOR2  g09665(.A(new_n10050_), .B(new_n1387_), .Y(new_n10051_));
  NOR2  g09666(.A(new_n10051_), .B(new_n1391_), .Y(new_n10052_));
  NOR2  g09667(.A(new_n10052_), .B(new_n1395_), .Y(new_n10053_));
  NOR2  g09668(.A(new_n10053_), .B(new_n1399_), .Y(new_n10054_));
  NOR2  g09669(.A(new_n10054_), .B(new_n1403_), .Y(new_n10055_));
  NOR2  g09670(.A(new_n10055_), .B(new_n1407_), .Y(new_n10056_));
  NOR2  g09671(.A(new_n10056_), .B(new_n1411_), .Y(new_n10057_));
  NOR2  g09672(.A(new_n10057_), .B(new_n1415_), .Y(new_n10058_));
  NOR2  g09673(.A(new_n10058_), .B(new_n1419_), .Y(new_n10059_));
  NOR2  g09674(.A(new_n10059_), .B(new_n1423_), .Y(new_n10060_));
  NOR2  g09675(.A(new_n10060_), .B(new_n1427_), .Y(new_n10061_));
  NOR2  g09676(.A(new_n10061_), .B(new_n1431_), .Y(new_n10062_));
  NOR2  g09677(.A(new_n10062_), .B(new_n1435_), .Y(new_n10063_));
  NOR2  g09678(.A(new_n10063_), .B(new_n1439_), .Y(new_n10064_));
  NOR2  g09679(.A(new_n10064_), .B(new_n1443_), .Y(new_n10065_));
  NOR2  g09680(.A(new_n10065_), .B(new_n1447_), .Y(new_n10066_));
  NAND2 g09681(.A(new_n1449_), .B(\req[100] ), .Y(new_n10067_));
  NOR2  g09682(.A(new_n10067_), .B(new_n10066_), .Y(\grant[100] ));
  INV   g09683(.A(new_n1458_), .Y(new_n10069_));
  NOR2  g09684(.A(new_n10069_), .B(new_n725_), .Y(new_n10070_));
  NOR2  g09685(.A(new_n10070_), .B(new_n1463_), .Y(new_n10071_));
  NOR2  g09686(.A(new_n10071_), .B(new_n1467_), .Y(new_n10072_));
  NOR2  g09687(.A(new_n10072_), .B(new_n1471_), .Y(new_n10073_));
  NOR2  g09688(.A(new_n10073_), .B(new_n1475_), .Y(new_n10074_));
  NOR2  g09689(.A(new_n10074_), .B(new_n1479_), .Y(new_n10075_));
  NOR2  g09690(.A(new_n10075_), .B(new_n1483_), .Y(new_n10076_));
  NOR2  g09691(.A(new_n10076_), .B(new_n1487_), .Y(new_n10077_));
  NOR2  g09692(.A(new_n10077_), .B(new_n1491_), .Y(new_n10078_));
  NOR2  g09693(.A(new_n10078_), .B(new_n1495_), .Y(new_n10079_));
  NOR2  g09694(.A(new_n10079_), .B(new_n1499_), .Y(new_n10080_));
  NOR2  g09695(.A(new_n10080_), .B(new_n1503_), .Y(new_n10081_));
  NOR2  g09696(.A(new_n10081_), .B(new_n1507_), .Y(new_n10082_));
  NOR2  g09697(.A(new_n10082_), .B(new_n1511_), .Y(new_n10083_));
  NOR2  g09698(.A(new_n10083_), .B(new_n1515_), .Y(new_n10084_));
  NOR2  g09699(.A(new_n10084_), .B(new_n1519_), .Y(new_n10085_));
  NOR2  g09700(.A(new_n10085_), .B(new_n1523_), .Y(new_n10086_));
  NOR2  g09701(.A(new_n10086_), .B(new_n1527_), .Y(new_n10087_));
  NOR2  g09702(.A(new_n10087_), .B(new_n1797_), .Y(new_n10088_));
  NOR2  g09703(.A(new_n10088_), .B(new_n396_), .Y(new_n10089_));
  NOR2  g09704(.A(new_n10089_), .B(new_n400_), .Y(new_n10090_));
  NOR2  g09705(.A(new_n10090_), .B(new_n406_), .Y(new_n10091_));
  NOR2  g09706(.A(new_n10091_), .B(new_n410_), .Y(new_n10092_));
  NOR2  g09707(.A(new_n10092_), .B(new_n416_), .Y(new_n10093_));
  NOR2  g09708(.A(new_n10093_), .B(new_n420_), .Y(new_n10094_));
  NOR2  g09709(.A(new_n10094_), .B(new_n426_), .Y(new_n10095_));
  NOR2  g09710(.A(new_n10095_), .B(new_n430_), .Y(new_n10096_));
  NOR2  g09711(.A(new_n10096_), .B(new_n436_), .Y(new_n10097_));
  NOR2  g09712(.A(new_n10097_), .B(new_n440_), .Y(new_n10098_));
  NOR2  g09713(.A(new_n10098_), .B(new_n446_), .Y(new_n10099_));
  NOR2  g09714(.A(new_n10099_), .B(new_n450_), .Y(new_n10100_));
  NOR2  g09715(.A(new_n10100_), .B(new_n456_), .Y(new_n10101_));
  NOR2  g09716(.A(new_n10101_), .B(new_n460_), .Y(new_n10102_));
  NOR2  g09717(.A(new_n10102_), .B(new_n466_), .Y(new_n10103_));
  NOR2  g09718(.A(new_n10103_), .B(new_n470_), .Y(new_n10104_));
  NOR2  g09719(.A(new_n10104_), .B(new_n476_), .Y(new_n10105_));
  NOR2  g09720(.A(new_n10105_), .B(new_n480_), .Y(new_n10106_));
  NOR2  g09721(.A(new_n10106_), .B(new_n486_), .Y(new_n10107_));
  NOR2  g09722(.A(new_n10107_), .B(new_n490_), .Y(new_n10108_));
  NOR2  g09723(.A(new_n10108_), .B(new_n496_), .Y(new_n10109_));
  NOR2  g09724(.A(new_n10109_), .B(new_n500_), .Y(new_n10110_));
  NOR2  g09725(.A(new_n10110_), .B(new_n506_), .Y(new_n10111_));
  NOR2  g09726(.A(new_n10111_), .B(new_n510_), .Y(new_n10112_));
  NOR2  g09727(.A(new_n10112_), .B(new_n516_), .Y(new_n10113_));
  NOR2  g09728(.A(new_n10113_), .B(new_n520_), .Y(new_n10114_));
  NOR2  g09729(.A(new_n10114_), .B(new_n526_), .Y(new_n10115_));
  NOR2  g09730(.A(new_n10115_), .B(new_n530_), .Y(new_n10116_));
  NOR2  g09731(.A(new_n10116_), .B(new_n536_), .Y(new_n10117_));
  NOR2  g09732(.A(new_n10117_), .B(new_n540_), .Y(new_n10118_));
  NOR2  g09733(.A(new_n10118_), .B(new_n546_), .Y(new_n10119_));
  NOR2  g09734(.A(new_n10119_), .B(new_n550_), .Y(new_n10120_));
  NOR2  g09735(.A(new_n10120_), .B(new_n556_), .Y(new_n10121_));
  NOR2  g09736(.A(new_n10121_), .B(new_n560_), .Y(new_n10122_));
  NOR2  g09737(.A(new_n10122_), .B(new_n566_), .Y(new_n10123_));
  NOR2  g09738(.A(new_n10123_), .B(new_n570_), .Y(new_n10124_));
  NOR2  g09739(.A(new_n10124_), .B(new_n576_), .Y(new_n10125_));
  NOR2  g09740(.A(new_n10125_), .B(new_n580_), .Y(new_n10126_));
  NOR2  g09741(.A(new_n10126_), .B(new_n586_), .Y(new_n10127_));
  NOR2  g09742(.A(new_n10127_), .B(new_n590_), .Y(new_n10128_));
  NOR2  g09743(.A(new_n10128_), .B(new_n596_), .Y(new_n10129_));
  NOR2  g09744(.A(new_n10129_), .B(new_n600_), .Y(new_n10130_));
  NOR2  g09745(.A(new_n10130_), .B(new_n606_), .Y(new_n10131_));
  NOR2  g09746(.A(new_n10131_), .B(new_n610_), .Y(new_n10132_));
  NOR2  g09747(.A(new_n10132_), .B(new_n616_), .Y(new_n10133_));
  NOR2  g09748(.A(new_n10133_), .B(new_n620_), .Y(new_n10134_));
  NOR2  g09749(.A(new_n10134_), .B(new_n626_), .Y(new_n10135_));
  NOR2  g09750(.A(new_n10135_), .B(new_n630_), .Y(new_n10136_));
  NOR2  g09751(.A(new_n10136_), .B(new_n636_), .Y(new_n10137_));
  NOR2  g09752(.A(new_n10137_), .B(new_n640_), .Y(new_n10138_));
  NOR2  g09753(.A(new_n10138_), .B(new_n646_), .Y(new_n10139_));
  NOR2  g09754(.A(new_n10139_), .B(new_n650_), .Y(new_n10140_));
  NOR2  g09755(.A(new_n10140_), .B(new_n656_), .Y(new_n10141_));
  NOR2  g09756(.A(new_n10141_), .B(new_n660_), .Y(new_n10142_));
  NOR2  g09757(.A(new_n10142_), .B(new_n666_), .Y(new_n10143_));
  NOR2  g09758(.A(new_n10143_), .B(new_n670_), .Y(new_n10144_));
  NOR2  g09759(.A(new_n10144_), .B(new_n676_), .Y(new_n10145_));
  NOR2  g09760(.A(new_n10145_), .B(new_n680_), .Y(new_n10146_));
  NOR2  g09761(.A(new_n10146_), .B(new_n686_), .Y(new_n10147_));
  NOR2  g09762(.A(new_n10147_), .B(new_n690_), .Y(new_n10148_));
  NOR2  g09763(.A(new_n10148_), .B(new_n696_), .Y(new_n10149_));
  NOR2  g09764(.A(new_n10149_), .B(new_n700_), .Y(new_n10150_));
  NOR2  g09765(.A(new_n10150_), .B(new_n706_), .Y(new_n10151_));
  NOR2  g09766(.A(new_n10151_), .B(new_n710_), .Y(new_n10152_));
  NOR2  g09767(.A(new_n10152_), .B(new_n716_), .Y(new_n10153_));
  NAND2 g09768(.A(new_n718_), .B(\req[101] ), .Y(new_n10154_));
  NOR2  g09769(.A(new_n10154_), .B(new_n10153_), .Y(\grant[101] ));
  INV   g09770(.A(new_n729_), .Y(new_n10156_));
  NOR2  g09771(.A(new_n1116_), .B(new_n10156_), .Y(new_n10157_));
  NOR2  g09772(.A(new_n10157_), .B(new_n736_), .Y(new_n10158_));
  NOR2  g09773(.A(new_n10158_), .B(new_n740_), .Y(new_n10159_));
  NOR2  g09774(.A(new_n10159_), .B(new_n746_), .Y(new_n10160_));
  NOR2  g09775(.A(new_n10160_), .B(new_n750_), .Y(new_n10161_));
  NOR2  g09776(.A(new_n10161_), .B(new_n756_), .Y(new_n10162_));
  NOR2  g09777(.A(new_n10162_), .B(new_n760_), .Y(new_n10163_));
  NOR2  g09778(.A(new_n10163_), .B(new_n766_), .Y(new_n10164_));
  NOR2  g09779(.A(new_n10164_), .B(new_n770_), .Y(new_n10165_));
  NOR2  g09780(.A(new_n10165_), .B(new_n776_), .Y(new_n10166_));
  NOR2  g09781(.A(new_n10166_), .B(new_n780_), .Y(new_n10167_));
  NOR2  g09782(.A(new_n10167_), .B(new_n786_), .Y(new_n10168_));
  NOR2  g09783(.A(new_n10168_), .B(new_n790_), .Y(new_n10169_));
  NOR2  g09784(.A(new_n10169_), .B(new_n796_), .Y(new_n10170_));
  NOR2  g09785(.A(new_n10170_), .B(new_n800_), .Y(new_n10171_));
  NOR2  g09786(.A(new_n10171_), .B(new_n806_), .Y(new_n10172_));
  NOR2  g09787(.A(new_n10172_), .B(new_n1616_), .Y(new_n10173_));
  NOR2  g09788(.A(new_n10173_), .B(new_n1618_), .Y(new_n10174_));
  NOR2  g09789(.A(new_n10174_), .B(new_n1885_), .Y(new_n10175_));
  NOR2  g09790(.A(new_n10175_), .B(new_n820_), .Y(new_n10176_));
  NOR2  g09791(.A(new_n10176_), .B(new_n824_), .Y(new_n10177_));
  NOR2  g09792(.A(new_n10177_), .B(new_n829_), .Y(new_n10178_));
  NOR2  g09793(.A(new_n10178_), .B(new_n833_), .Y(new_n10179_));
  NOR2  g09794(.A(new_n10179_), .B(new_n838_), .Y(new_n10180_));
  NOR2  g09795(.A(new_n10180_), .B(new_n842_), .Y(new_n10181_));
  NOR2  g09796(.A(new_n10181_), .B(new_n847_), .Y(new_n10182_));
  NOR2  g09797(.A(new_n10182_), .B(new_n851_), .Y(new_n10183_));
  NOR2  g09798(.A(new_n10183_), .B(new_n856_), .Y(new_n10184_));
  NOR2  g09799(.A(new_n10184_), .B(new_n860_), .Y(new_n10185_));
  NOR2  g09800(.A(new_n10185_), .B(new_n865_), .Y(new_n10186_));
  NOR2  g09801(.A(new_n10186_), .B(new_n869_), .Y(new_n10187_));
  NOR2  g09802(.A(new_n10187_), .B(new_n874_), .Y(new_n10188_));
  NOR2  g09803(.A(new_n10188_), .B(new_n878_), .Y(new_n10189_));
  NOR2  g09804(.A(new_n10189_), .B(new_n883_), .Y(new_n10190_));
  NOR2  g09805(.A(new_n10190_), .B(new_n887_), .Y(new_n10191_));
  NOR2  g09806(.A(new_n10191_), .B(new_n892_), .Y(new_n10192_));
  NOR2  g09807(.A(new_n10192_), .B(new_n896_), .Y(new_n10193_));
  NOR2  g09808(.A(new_n10193_), .B(new_n901_), .Y(new_n10194_));
  NOR2  g09809(.A(new_n10194_), .B(new_n905_), .Y(new_n10195_));
  NOR2  g09810(.A(new_n10195_), .B(new_n910_), .Y(new_n10196_));
  NOR2  g09811(.A(new_n10196_), .B(new_n914_), .Y(new_n10197_));
  NOR2  g09812(.A(new_n10197_), .B(new_n919_), .Y(new_n10198_));
  NOR2  g09813(.A(new_n10198_), .B(new_n923_), .Y(new_n10199_));
  NOR2  g09814(.A(new_n10199_), .B(new_n928_), .Y(new_n10200_));
  NOR2  g09815(.A(new_n10200_), .B(new_n932_), .Y(new_n10201_));
  NOR2  g09816(.A(new_n10201_), .B(new_n937_), .Y(new_n10202_));
  NOR2  g09817(.A(new_n10202_), .B(new_n941_), .Y(new_n10203_));
  NOR2  g09818(.A(new_n10203_), .B(new_n946_), .Y(new_n10204_));
  NOR2  g09819(.A(new_n10204_), .B(new_n950_), .Y(new_n10205_));
  NOR2  g09820(.A(new_n10205_), .B(new_n955_), .Y(new_n10206_));
  NOR2  g09821(.A(new_n10206_), .B(new_n959_), .Y(new_n10207_));
  NOR2  g09822(.A(new_n10207_), .B(new_n964_), .Y(new_n10208_));
  NOR2  g09823(.A(new_n10208_), .B(new_n968_), .Y(new_n10209_));
  NOR2  g09824(.A(new_n10209_), .B(new_n973_), .Y(new_n10210_));
  NOR2  g09825(.A(new_n10210_), .B(new_n977_), .Y(new_n10211_));
  NOR2  g09826(.A(new_n10211_), .B(new_n982_), .Y(new_n10212_));
  NOR2  g09827(.A(new_n10212_), .B(new_n986_), .Y(new_n10213_));
  NOR2  g09828(.A(new_n10213_), .B(new_n991_), .Y(new_n10214_));
  NOR2  g09829(.A(new_n10214_), .B(new_n995_), .Y(new_n10215_));
  NOR2  g09830(.A(new_n10215_), .B(new_n1000_), .Y(new_n10216_));
  NOR2  g09831(.A(new_n10216_), .B(new_n1004_), .Y(new_n10217_));
  NOR2  g09832(.A(new_n10217_), .B(new_n1009_), .Y(new_n10218_));
  NOR2  g09833(.A(new_n10218_), .B(new_n1013_), .Y(new_n10219_));
  NOR2  g09834(.A(new_n10219_), .B(new_n1018_), .Y(new_n10220_));
  NOR2  g09835(.A(new_n10220_), .B(new_n1022_), .Y(new_n10221_));
  NOR2  g09836(.A(new_n10221_), .B(new_n1027_), .Y(new_n10222_));
  NOR2  g09837(.A(new_n10222_), .B(new_n1031_), .Y(new_n10223_));
  NOR2  g09838(.A(new_n10223_), .B(new_n1036_), .Y(new_n10224_));
  NOR2  g09839(.A(new_n10224_), .B(new_n1040_), .Y(new_n10225_));
  NOR2  g09840(.A(new_n10225_), .B(new_n1045_), .Y(new_n10226_));
  NOR2  g09841(.A(new_n10226_), .B(new_n1049_), .Y(new_n10227_));
  NOR2  g09842(.A(new_n10227_), .B(new_n1054_), .Y(new_n10228_));
  NOR2  g09843(.A(new_n10228_), .B(new_n1058_), .Y(new_n10229_));
  NOR2  g09844(.A(new_n10229_), .B(new_n1063_), .Y(new_n10230_));
  NOR2  g09845(.A(new_n10230_), .B(new_n1067_), .Y(new_n10231_));
  NOR2  g09846(.A(new_n10231_), .B(new_n1072_), .Y(new_n10232_));
  NOR2  g09847(.A(new_n10232_), .B(new_n1076_), .Y(new_n10233_));
  NOR2  g09848(.A(new_n10233_), .B(new_n1081_), .Y(new_n10234_));
  NOR2  g09849(.A(new_n10234_), .B(new_n1085_), .Y(new_n10235_));
  NOR2  g09850(.A(new_n10235_), .B(new_n1090_), .Y(new_n10236_));
  NOR2  g09851(.A(new_n10236_), .B(new_n1094_), .Y(new_n10237_));
  NOR2  g09852(.A(new_n10237_), .B(new_n1099_), .Y(new_n10238_));
  NOR2  g09853(.A(new_n10238_), .B(new_n1103_), .Y(new_n10239_));
  NOR2  g09854(.A(new_n10239_), .B(new_n1108_), .Y(new_n10240_));
  NAND2 g09855(.A(new_n1110_), .B(\req[102] ), .Y(new_n10241_));
  NOR2  g09856(.A(new_n10241_), .B(new_n10240_), .Y(\grant[102] ));
  INV   g09857(.A(new_n1120_), .Y(new_n10243_));
  NOR2  g09858(.A(new_n1462_), .B(new_n10243_), .Y(new_n10244_));
  NOR2  g09859(.A(new_n10244_), .B(new_n1126_), .Y(new_n10245_));
  NOR2  g09860(.A(new_n10245_), .B(new_n1130_), .Y(new_n10246_));
  NOR2  g09861(.A(new_n10246_), .B(new_n1135_), .Y(new_n10247_));
  NOR2  g09862(.A(new_n10247_), .B(new_n1139_), .Y(new_n10248_));
  NOR2  g09863(.A(new_n10248_), .B(new_n1144_), .Y(new_n10249_));
  NOR2  g09864(.A(new_n10249_), .B(new_n1148_), .Y(new_n10250_));
  NOR2  g09865(.A(new_n10250_), .B(new_n1153_), .Y(new_n10251_));
  NOR2  g09866(.A(new_n10251_), .B(new_n1157_), .Y(new_n10252_));
  NOR2  g09867(.A(new_n10252_), .B(new_n1162_), .Y(new_n10253_));
  NOR2  g09868(.A(new_n10253_), .B(new_n1166_), .Y(new_n10254_));
  NOR2  g09869(.A(new_n10254_), .B(new_n1171_), .Y(new_n10255_));
  NOR2  g09870(.A(new_n10255_), .B(new_n1175_), .Y(new_n10256_));
  NOR2  g09871(.A(new_n10256_), .B(new_n1180_), .Y(new_n10257_));
  NOR2  g09872(.A(new_n10257_), .B(new_n1184_), .Y(new_n10258_));
  NOR2  g09873(.A(new_n10258_), .B(new_n1189_), .Y(new_n10259_));
  NOR2  g09874(.A(new_n10259_), .B(new_n1707_), .Y(new_n10260_));
  NOR2  g09875(.A(new_n10260_), .B(new_n1709_), .Y(new_n10261_));
  NOR2  g09876(.A(new_n10261_), .B(new_n1973_), .Y(new_n10262_));
  NOR2  g09877(.A(new_n10262_), .B(new_n1199_), .Y(new_n10263_));
  NOR2  g09878(.A(new_n10263_), .B(new_n1203_), .Y(new_n10264_));
  NOR2  g09879(.A(new_n10264_), .B(new_n1207_), .Y(new_n10265_));
  NOR2  g09880(.A(new_n10265_), .B(new_n1211_), .Y(new_n10266_));
  NOR2  g09881(.A(new_n10266_), .B(new_n1215_), .Y(new_n10267_));
  NOR2  g09882(.A(new_n10267_), .B(new_n1219_), .Y(new_n10268_));
  NOR2  g09883(.A(new_n10268_), .B(new_n1223_), .Y(new_n10269_));
  NOR2  g09884(.A(new_n10269_), .B(new_n1227_), .Y(new_n10270_));
  NOR2  g09885(.A(new_n10270_), .B(new_n1231_), .Y(new_n10271_));
  NOR2  g09886(.A(new_n10271_), .B(new_n1235_), .Y(new_n10272_));
  NOR2  g09887(.A(new_n10272_), .B(new_n1239_), .Y(new_n10273_));
  NOR2  g09888(.A(new_n10273_), .B(new_n1243_), .Y(new_n10274_));
  NOR2  g09889(.A(new_n10274_), .B(new_n1247_), .Y(new_n10275_));
  NOR2  g09890(.A(new_n10275_), .B(new_n1251_), .Y(new_n10276_));
  NOR2  g09891(.A(new_n10276_), .B(new_n1255_), .Y(new_n10277_));
  NOR2  g09892(.A(new_n10277_), .B(new_n1259_), .Y(new_n10278_));
  NOR2  g09893(.A(new_n10278_), .B(new_n1263_), .Y(new_n10279_));
  NOR2  g09894(.A(new_n10279_), .B(new_n1267_), .Y(new_n10280_));
  NOR2  g09895(.A(new_n10280_), .B(new_n1271_), .Y(new_n10281_));
  NOR2  g09896(.A(new_n10281_), .B(new_n1275_), .Y(new_n10282_));
  NOR2  g09897(.A(new_n10282_), .B(new_n1279_), .Y(new_n10283_));
  NOR2  g09898(.A(new_n10283_), .B(new_n1283_), .Y(new_n10284_));
  NOR2  g09899(.A(new_n10284_), .B(new_n1287_), .Y(new_n10285_));
  NOR2  g09900(.A(new_n10285_), .B(new_n1291_), .Y(new_n10286_));
  NOR2  g09901(.A(new_n10286_), .B(new_n1295_), .Y(new_n10287_));
  NOR2  g09902(.A(new_n10287_), .B(new_n1299_), .Y(new_n10288_));
  NOR2  g09903(.A(new_n10288_), .B(new_n1303_), .Y(new_n10289_));
  NOR2  g09904(.A(new_n10289_), .B(new_n1307_), .Y(new_n10290_));
  NOR2  g09905(.A(new_n10290_), .B(new_n1311_), .Y(new_n10291_));
  NOR2  g09906(.A(new_n10291_), .B(new_n1315_), .Y(new_n10292_));
  NOR2  g09907(.A(new_n10292_), .B(new_n1319_), .Y(new_n10293_));
  NOR2  g09908(.A(new_n10293_), .B(new_n1323_), .Y(new_n10294_));
  NOR2  g09909(.A(new_n10294_), .B(new_n1327_), .Y(new_n10295_));
  NOR2  g09910(.A(new_n10295_), .B(new_n1331_), .Y(new_n10296_));
  NOR2  g09911(.A(new_n10296_), .B(new_n1335_), .Y(new_n10297_));
  NOR2  g09912(.A(new_n10297_), .B(new_n1339_), .Y(new_n10298_));
  NOR2  g09913(.A(new_n10298_), .B(new_n1343_), .Y(new_n10299_));
  NOR2  g09914(.A(new_n10299_), .B(new_n1347_), .Y(new_n10300_));
  NOR2  g09915(.A(new_n10300_), .B(new_n1351_), .Y(new_n10301_));
  NOR2  g09916(.A(new_n10301_), .B(new_n1355_), .Y(new_n10302_));
  NOR2  g09917(.A(new_n10302_), .B(new_n1359_), .Y(new_n10303_));
  NOR2  g09918(.A(new_n10303_), .B(new_n1363_), .Y(new_n10304_));
  NOR2  g09919(.A(new_n10304_), .B(new_n1367_), .Y(new_n10305_));
  NOR2  g09920(.A(new_n10305_), .B(new_n1371_), .Y(new_n10306_));
  NOR2  g09921(.A(new_n10306_), .B(new_n1375_), .Y(new_n10307_));
  NOR2  g09922(.A(new_n10307_), .B(new_n1379_), .Y(new_n10308_));
  NOR2  g09923(.A(new_n10308_), .B(new_n1383_), .Y(new_n10309_));
  NOR2  g09924(.A(new_n10309_), .B(new_n1387_), .Y(new_n10310_));
  NOR2  g09925(.A(new_n10310_), .B(new_n1391_), .Y(new_n10311_));
  NOR2  g09926(.A(new_n10311_), .B(new_n1395_), .Y(new_n10312_));
  NOR2  g09927(.A(new_n10312_), .B(new_n1399_), .Y(new_n10313_));
  NOR2  g09928(.A(new_n10313_), .B(new_n1403_), .Y(new_n10314_));
  NOR2  g09929(.A(new_n10314_), .B(new_n1407_), .Y(new_n10315_));
  NOR2  g09930(.A(new_n10315_), .B(new_n1411_), .Y(new_n10316_));
  NOR2  g09931(.A(new_n10316_), .B(new_n1415_), .Y(new_n10317_));
  NOR2  g09932(.A(new_n10317_), .B(new_n1419_), .Y(new_n10318_));
  NOR2  g09933(.A(new_n10318_), .B(new_n1423_), .Y(new_n10319_));
  NOR2  g09934(.A(new_n10319_), .B(new_n1427_), .Y(new_n10320_));
  NOR2  g09935(.A(new_n10320_), .B(new_n1431_), .Y(new_n10321_));
  NOR2  g09936(.A(new_n10321_), .B(new_n1435_), .Y(new_n10322_));
  NOR2  g09937(.A(new_n10322_), .B(new_n1439_), .Y(new_n10323_));
  NOR2  g09938(.A(new_n10323_), .B(new_n1443_), .Y(new_n10324_));
  NOR2  g09939(.A(new_n10324_), .B(new_n1447_), .Y(new_n10325_));
  NOR2  g09940(.A(new_n10325_), .B(new_n1451_), .Y(new_n10326_));
  NOR2  g09941(.A(new_n10326_), .B(new_n1455_), .Y(new_n10327_));
  NAND2 g09942(.A(new_n1457_), .B(\req[103] ), .Y(new_n10328_));
  NOR2  g09943(.A(new_n10328_), .B(new_n10327_), .Y(\grant[103] ));
  INV   g09944(.A(new_n1466_), .Y(new_n10330_));
  NOR2  g09945(.A(new_n10330_), .B(new_n735_), .Y(new_n10331_));
  NOR2  g09946(.A(new_n10331_), .B(new_n1471_), .Y(new_n10332_));
  NOR2  g09947(.A(new_n10332_), .B(new_n1475_), .Y(new_n10333_));
  NOR2  g09948(.A(new_n10333_), .B(new_n1479_), .Y(new_n10334_));
  NOR2  g09949(.A(new_n10334_), .B(new_n1483_), .Y(new_n10335_));
  NOR2  g09950(.A(new_n10335_), .B(new_n1487_), .Y(new_n10336_));
  NOR2  g09951(.A(new_n10336_), .B(new_n1491_), .Y(new_n10337_));
  NOR2  g09952(.A(new_n10337_), .B(new_n1495_), .Y(new_n10338_));
  NOR2  g09953(.A(new_n10338_), .B(new_n1499_), .Y(new_n10339_));
  NOR2  g09954(.A(new_n10339_), .B(new_n1503_), .Y(new_n10340_));
  NOR2  g09955(.A(new_n10340_), .B(new_n1507_), .Y(new_n10341_));
  NOR2  g09956(.A(new_n10341_), .B(new_n1511_), .Y(new_n10342_));
  NOR2  g09957(.A(new_n10342_), .B(new_n1515_), .Y(new_n10343_));
  NOR2  g09958(.A(new_n10343_), .B(new_n1519_), .Y(new_n10344_));
  NOR2  g09959(.A(new_n10344_), .B(new_n1523_), .Y(new_n10345_));
  NOR2  g09960(.A(new_n10345_), .B(new_n1527_), .Y(new_n10346_));
  NOR2  g09961(.A(new_n10346_), .B(new_n1797_), .Y(new_n10347_));
  NOR2  g09962(.A(new_n10347_), .B(new_n396_), .Y(new_n10348_));
  NOR2  g09963(.A(new_n10348_), .B(new_n400_), .Y(new_n10349_));
  NOR2  g09964(.A(new_n10349_), .B(new_n406_), .Y(new_n10350_));
  NOR2  g09965(.A(new_n10350_), .B(new_n410_), .Y(new_n10351_));
  NOR2  g09966(.A(new_n10351_), .B(new_n416_), .Y(new_n10352_));
  NOR2  g09967(.A(new_n10352_), .B(new_n420_), .Y(new_n10353_));
  NOR2  g09968(.A(new_n10353_), .B(new_n426_), .Y(new_n10354_));
  NOR2  g09969(.A(new_n10354_), .B(new_n430_), .Y(new_n10355_));
  NOR2  g09970(.A(new_n10355_), .B(new_n436_), .Y(new_n10356_));
  NOR2  g09971(.A(new_n10356_), .B(new_n440_), .Y(new_n10357_));
  NOR2  g09972(.A(new_n10357_), .B(new_n446_), .Y(new_n10358_));
  NOR2  g09973(.A(new_n10358_), .B(new_n450_), .Y(new_n10359_));
  NOR2  g09974(.A(new_n10359_), .B(new_n456_), .Y(new_n10360_));
  NOR2  g09975(.A(new_n10360_), .B(new_n460_), .Y(new_n10361_));
  NOR2  g09976(.A(new_n10361_), .B(new_n466_), .Y(new_n10362_));
  NOR2  g09977(.A(new_n10362_), .B(new_n470_), .Y(new_n10363_));
  NOR2  g09978(.A(new_n10363_), .B(new_n476_), .Y(new_n10364_));
  NOR2  g09979(.A(new_n10364_), .B(new_n480_), .Y(new_n10365_));
  NOR2  g09980(.A(new_n10365_), .B(new_n486_), .Y(new_n10366_));
  NOR2  g09981(.A(new_n10366_), .B(new_n490_), .Y(new_n10367_));
  NOR2  g09982(.A(new_n10367_), .B(new_n496_), .Y(new_n10368_));
  NOR2  g09983(.A(new_n10368_), .B(new_n500_), .Y(new_n10369_));
  NOR2  g09984(.A(new_n10369_), .B(new_n506_), .Y(new_n10370_));
  NOR2  g09985(.A(new_n10370_), .B(new_n510_), .Y(new_n10371_));
  NOR2  g09986(.A(new_n10371_), .B(new_n516_), .Y(new_n10372_));
  NOR2  g09987(.A(new_n10372_), .B(new_n520_), .Y(new_n10373_));
  NOR2  g09988(.A(new_n10373_), .B(new_n526_), .Y(new_n10374_));
  NOR2  g09989(.A(new_n10374_), .B(new_n530_), .Y(new_n10375_));
  NOR2  g09990(.A(new_n10375_), .B(new_n536_), .Y(new_n10376_));
  NOR2  g09991(.A(new_n10376_), .B(new_n540_), .Y(new_n10377_));
  NOR2  g09992(.A(new_n10377_), .B(new_n546_), .Y(new_n10378_));
  NOR2  g09993(.A(new_n10378_), .B(new_n550_), .Y(new_n10379_));
  NOR2  g09994(.A(new_n10379_), .B(new_n556_), .Y(new_n10380_));
  NOR2  g09995(.A(new_n10380_), .B(new_n560_), .Y(new_n10381_));
  NOR2  g09996(.A(new_n10381_), .B(new_n566_), .Y(new_n10382_));
  NOR2  g09997(.A(new_n10382_), .B(new_n570_), .Y(new_n10383_));
  NOR2  g09998(.A(new_n10383_), .B(new_n576_), .Y(new_n10384_));
  NOR2  g09999(.A(new_n10384_), .B(new_n580_), .Y(new_n10385_));
  NOR2  g10000(.A(new_n10385_), .B(new_n586_), .Y(new_n10386_));
  NOR2  g10001(.A(new_n10386_), .B(new_n590_), .Y(new_n10387_));
  NOR2  g10002(.A(new_n10387_), .B(new_n596_), .Y(new_n10388_));
  NOR2  g10003(.A(new_n10388_), .B(new_n600_), .Y(new_n10389_));
  NOR2  g10004(.A(new_n10389_), .B(new_n606_), .Y(new_n10390_));
  NOR2  g10005(.A(new_n10390_), .B(new_n610_), .Y(new_n10391_));
  NOR2  g10006(.A(new_n10391_), .B(new_n616_), .Y(new_n10392_));
  NOR2  g10007(.A(new_n10392_), .B(new_n620_), .Y(new_n10393_));
  NOR2  g10008(.A(new_n10393_), .B(new_n626_), .Y(new_n10394_));
  NOR2  g10009(.A(new_n10394_), .B(new_n630_), .Y(new_n10395_));
  NOR2  g10010(.A(new_n10395_), .B(new_n636_), .Y(new_n10396_));
  NOR2  g10011(.A(new_n10396_), .B(new_n640_), .Y(new_n10397_));
  NOR2  g10012(.A(new_n10397_), .B(new_n646_), .Y(new_n10398_));
  NOR2  g10013(.A(new_n10398_), .B(new_n650_), .Y(new_n10399_));
  NOR2  g10014(.A(new_n10399_), .B(new_n656_), .Y(new_n10400_));
  NOR2  g10015(.A(new_n10400_), .B(new_n660_), .Y(new_n10401_));
  NOR2  g10016(.A(new_n10401_), .B(new_n666_), .Y(new_n10402_));
  NOR2  g10017(.A(new_n10402_), .B(new_n670_), .Y(new_n10403_));
  NOR2  g10018(.A(new_n10403_), .B(new_n676_), .Y(new_n10404_));
  NOR2  g10019(.A(new_n10404_), .B(new_n680_), .Y(new_n10405_));
  NOR2  g10020(.A(new_n10405_), .B(new_n686_), .Y(new_n10406_));
  NOR2  g10021(.A(new_n10406_), .B(new_n690_), .Y(new_n10407_));
  NOR2  g10022(.A(new_n10407_), .B(new_n696_), .Y(new_n10408_));
  NOR2  g10023(.A(new_n10408_), .B(new_n700_), .Y(new_n10409_));
  NOR2  g10024(.A(new_n10409_), .B(new_n706_), .Y(new_n10410_));
  NOR2  g10025(.A(new_n10410_), .B(new_n710_), .Y(new_n10411_));
  NOR2  g10026(.A(new_n10411_), .B(new_n716_), .Y(new_n10412_));
  NOR2  g10027(.A(new_n10412_), .B(new_n720_), .Y(new_n10413_));
  NOR2  g10028(.A(new_n10413_), .B(new_n726_), .Y(new_n10414_));
  NAND2 g10029(.A(new_n728_), .B(\req[104] ), .Y(new_n10415_));
  NOR2  g10030(.A(new_n10415_), .B(new_n10414_), .Y(\grant[104] ));
  INV   g10031(.A(new_n739_), .Y(new_n10417_));
  NOR2  g10032(.A(new_n1125_), .B(new_n10417_), .Y(new_n10418_));
  NOR2  g10033(.A(new_n10418_), .B(new_n746_), .Y(new_n10419_));
  NOR2  g10034(.A(new_n10419_), .B(new_n750_), .Y(new_n10420_));
  NOR2  g10035(.A(new_n10420_), .B(new_n756_), .Y(new_n10421_));
  NOR2  g10036(.A(new_n10421_), .B(new_n760_), .Y(new_n10422_));
  NOR2  g10037(.A(new_n10422_), .B(new_n766_), .Y(new_n10423_));
  NOR2  g10038(.A(new_n10423_), .B(new_n770_), .Y(new_n10424_));
  NOR2  g10039(.A(new_n10424_), .B(new_n776_), .Y(new_n10425_));
  NOR2  g10040(.A(new_n10425_), .B(new_n780_), .Y(new_n10426_));
  NOR2  g10041(.A(new_n10426_), .B(new_n786_), .Y(new_n10427_));
  NOR2  g10042(.A(new_n10427_), .B(new_n790_), .Y(new_n10428_));
  NOR2  g10043(.A(new_n10428_), .B(new_n796_), .Y(new_n10429_));
  NOR2  g10044(.A(new_n10429_), .B(new_n800_), .Y(new_n10430_));
  NOR2  g10045(.A(new_n10430_), .B(new_n806_), .Y(new_n10431_));
  NOR2  g10046(.A(new_n10431_), .B(new_n1616_), .Y(new_n10432_));
  NOR2  g10047(.A(new_n10432_), .B(new_n1618_), .Y(new_n10433_));
  NOR2  g10048(.A(new_n10433_), .B(new_n1885_), .Y(new_n10434_));
  NOR2  g10049(.A(new_n10434_), .B(new_n820_), .Y(new_n10435_));
  NOR2  g10050(.A(new_n10435_), .B(new_n824_), .Y(new_n10436_));
  NOR2  g10051(.A(new_n10436_), .B(new_n829_), .Y(new_n10437_));
  NOR2  g10052(.A(new_n10437_), .B(new_n833_), .Y(new_n10438_));
  NOR2  g10053(.A(new_n10438_), .B(new_n838_), .Y(new_n10439_));
  NOR2  g10054(.A(new_n10439_), .B(new_n842_), .Y(new_n10440_));
  NOR2  g10055(.A(new_n10440_), .B(new_n847_), .Y(new_n10441_));
  NOR2  g10056(.A(new_n10441_), .B(new_n851_), .Y(new_n10442_));
  NOR2  g10057(.A(new_n10442_), .B(new_n856_), .Y(new_n10443_));
  NOR2  g10058(.A(new_n10443_), .B(new_n860_), .Y(new_n10444_));
  NOR2  g10059(.A(new_n10444_), .B(new_n865_), .Y(new_n10445_));
  NOR2  g10060(.A(new_n10445_), .B(new_n869_), .Y(new_n10446_));
  NOR2  g10061(.A(new_n10446_), .B(new_n874_), .Y(new_n10447_));
  NOR2  g10062(.A(new_n10447_), .B(new_n878_), .Y(new_n10448_));
  NOR2  g10063(.A(new_n10448_), .B(new_n883_), .Y(new_n10449_));
  NOR2  g10064(.A(new_n10449_), .B(new_n887_), .Y(new_n10450_));
  NOR2  g10065(.A(new_n10450_), .B(new_n892_), .Y(new_n10451_));
  NOR2  g10066(.A(new_n10451_), .B(new_n896_), .Y(new_n10452_));
  NOR2  g10067(.A(new_n10452_), .B(new_n901_), .Y(new_n10453_));
  NOR2  g10068(.A(new_n10453_), .B(new_n905_), .Y(new_n10454_));
  NOR2  g10069(.A(new_n10454_), .B(new_n910_), .Y(new_n10455_));
  NOR2  g10070(.A(new_n10455_), .B(new_n914_), .Y(new_n10456_));
  NOR2  g10071(.A(new_n10456_), .B(new_n919_), .Y(new_n10457_));
  NOR2  g10072(.A(new_n10457_), .B(new_n923_), .Y(new_n10458_));
  NOR2  g10073(.A(new_n10458_), .B(new_n928_), .Y(new_n10459_));
  NOR2  g10074(.A(new_n10459_), .B(new_n932_), .Y(new_n10460_));
  NOR2  g10075(.A(new_n10460_), .B(new_n937_), .Y(new_n10461_));
  NOR2  g10076(.A(new_n10461_), .B(new_n941_), .Y(new_n10462_));
  NOR2  g10077(.A(new_n10462_), .B(new_n946_), .Y(new_n10463_));
  NOR2  g10078(.A(new_n10463_), .B(new_n950_), .Y(new_n10464_));
  NOR2  g10079(.A(new_n10464_), .B(new_n955_), .Y(new_n10465_));
  NOR2  g10080(.A(new_n10465_), .B(new_n959_), .Y(new_n10466_));
  NOR2  g10081(.A(new_n10466_), .B(new_n964_), .Y(new_n10467_));
  NOR2  g10082(.A(new_n10467_), .B(new_n968_), .Y(new_n10468_));
  NOR2  g10083(.A(new_n10468_), .B(new_n973_), .Y(new_n10469_));
  NOR2  g10084(.A(new_n10469_), .B(new_n977_), .Y(new_n10470_));
  NOR2  g10085(.A(new_n10470_), .B(new_n982_), .Y(new_n10471_));
  NOR2  g10086(.A(new_n10471_), .B(new_n986_), .Y(new_n10472_));
  NOR2  g10087(.A(new_n10472_), .B(new_n991_), .Y(new_n10473_));
  NOR2  g10088(.A(new_n10473_), .B(new_n995_), .Y(new_n10474_));
  NOR2  g10089(.A(new_n10474_), .B(new_n1000_), .Y(new_n10475_));
  NOR2  g10090(.A(new_n10475_), .B(new_n1004_), .Y(new_n10476_));
  NOR2  g10091(.A(new_n10476_), .B(new_n1009_), .Y(new_n10477_));
  NOR2  g10092(.A(new_n10477_), .B(new_n1013_), .Y(new_n10478_));
  NOR2  g10093(.A(new_n10478_), .B(new_n1018_), .Y(new_n10479_));
  NOR2  g10094(.A(new_n10479_), .B(new_n1022_), .Y(new_n10480_));
  NOR2  g10095(.A(new_n10480_), .B(new_n1027_), .Y(new_n10481_));
  NOR2  g10096(.A(new_n10481_), .B(new_n1031_), .Y(new_n10482_));
  NOR2  g10097(.A(new_n10482_), .B(new_n1036_), .Y(new_n10483_));
  NOR2  g10098(.A(new_n10483_), .B(new_n1040_), .Y(new_n10484_));
  NOR2  g10099(.A(new_n10484_), .B(new_n1045_), .Y(new_n10485_));
  NOR2  g10100(.A(new_n10485_), .B(new_n1049_), .Y(new_n10486_));
  NOR2  g10101(.A(new_n10486_), .B(new_n1054_), .Y(new_n10487_));
  NOR2  g10102(.A(new_n10487_), .B(new_n1058_), .Y(new_n10488_));
  NOR2  g10103(.A(new_n10488_), .B(new_n1063_), .Y(new_n10489_));
  NOR2  g10104(.A(new_n10489_), .B(new_n1067_), .Y(new_n10490_));
  NOR2  g10105(.A(new_n10490_), .B(new_n1072_), .Y(new_n10491_));
  NOR2  g10106(.A(new_n10491_), .B(new_n1076_), .Y(new_n10492_));
  NOR2  g10107(.A(new_n10492_), .B(new_n1081_), .Y(new_n10493_));
  NOR2  g10108(.A(new_n10493_), .B(new_n1085_), .Y(new_n10494_));
  NOR2  g10109(.A(new_n10494_), .B(new_n1090_), .Y(new_n10495_));
  NOR2  g10110(.A(new_n10495_), .B(new_n1094_), .Y(new_n10496_));
  NOR2  g10111(.A(new_n10496_), .B(new_n1099_), .Y(new_n10497_));
  NOR2  g10112(.A(new_n10497_), .B(new_n1103_), .Y(new_n10498_));
  NOR2  g10113(.A(new_n10498_), .B(new_n1108_), .Y(new_n10499_));
  NOR2  g10114(.A(new_n10499_), .B(new_n1112_), .Y(new_n10500_));
  NOR2  g10115(.A(new_n10500_), .B(new_n1117_), .Y(new_n10501_));
  NAND2 g10116(.A(new_n1119_), .B(\req[105] ), .Y(new_n10502_));
  NOR2  g10117(.A(new_n10502_), .B(new_n10501_), .Y(\grant[105] ));
  INV   g10118(.A(new_n1129_), .Y(new_n10504_));
  NOR2  g10119(.A(new_n1470_), .B(new_n10504_), .Y(new_n10505_));
  NOR2  g10120(.A(new_n10505_), .B(new_n1135_), .Y(new_n10506_));
  NOR2  g10121(.A(new_n10506_), .B(new_n1139_), .Y(new_n10507_));
  NOR2  g10122(.A(new_n10507_), .B(new_n1144_), .Y(new_n10508_));
  NOR2  g10123(.A(new_n10508_), .B(new_n1148_), .Y(new_n10509_));
  NOR2  g10124(.A(new_n10509_), .B(new_n1153_), .Y(new_n10510_));
  NOR2  g10125(.A(new_n10510_), .B(new_n1157_), .Y(new_n10511_));
  NOR2  g10126(.A(new_n10511_), .B(new_n1162_), .Y(new_n10512_));
  NOR2  g10127(.A(new_n10512_), .B(new_n1166_), .Y(new_n10513_));
  NOR2  g10128(.A(new_n10513_), .B(new_n1171_), .Y(new_n10514_));
  NOR2  g10129(.A(new_n10514_), .B(new_n1175_), .Y(new_n10515_));
  NOR2  g10130(.A(new_n10515_), .B(new_n1180_), .Y(new_n10516_));
  NOR2  g10131(.A(new_n10516_), .B(new_n1184_), .Y(new_n10517_));
  NOR2  g10132(.A(new_n10517_), .B(new_n1189_), .Y(new_n10518_));
  NOR2  g10133(.A(new_n10518_), .B(new_n1707_), .Y(new_n10519_));
  NOR2  g10134(.A(new_n10519_), .B(new_n1709_), .Y(new_n10520_));
  NOR2  g10135(.A(new_n10520_), .B(new_n1973_), .Y(new_n10521_));
  NOR2  g10136(.A(new_n10521_), .B(new_n1199_), .Y(new_n10522_));
  NOR2  g10137(.A(new_n10522_), .B(new_n1203_), .Y(new_n10523_));
  NOR2  g10138(.A(new_n10523_), .B(new_n1207_), .Y(new_n10524_));
  NOR2  g10139(.A(new_n10524_), .B(new_n1211_), .Y(new_n10525_));
  NOR2  g10140(.A(new_n10525_), .B(new_n1215_), .Y(new_n10526_));
  NOR2  g10141(.A(new_n10526_), .B(new_n1219_), .Y(new_n10527_));
  NOR2  g10142(.A(new_n10527_), .B(new_n1223_), .Y(new_n10528_));
  NOR2  g10143(.A(new_n10528_), .B(new_n1227_), .Y(new_n10529_));
  NOR2  g10144(.A(new_n10529_), .B(new_n1231_), .Y(new_n10530_));
  NOR2  g10145(.A(new_n10530_), .B(new_n1235_), .Y(new_n10531_));
  NOR2  g10146(.A(new_n10531_), .B(new_n1239_), .Y(new_n10532_));
  NOR2  g10147(.A(new_n10532_), .B(new_n1243_), .Y(new_n10533_));
  NOR2  g10148(.A(new_n10533_), .B(new_n1247_), .Y(new_n10534_));
  NOR2  g10149(.A(new_n10534_), .B(new_n1251_), .Y(new_n10535_));
  NOR2  g10150(.A(new_n10535_), .B(new_n1255_), .Y(new_n10536_));
  NOR2  g10151(.A(new_n10536_), .B(new_n1259_), .Y(new_n10537_));
  NOR2  g10152(.A(new_n10537_), .B(new_n1263_), .Y(new_n10538_));
  NOR2  g10153(.A(new_n10538_), .B(new_n1267_), .Y(new_n10539_));
  NOR2  g10154(.A(new_n10539_), .B(new_n1271_), .Y(new_n10540_));
  NOR2  g10155(.A(new_n10540_), .B(new_n1275_), .Y(new_n10541_));
  NOR2  g10156(.A(new_n10541_), .B(new_n1279_), .Y(new_n10542_));
  NOR2  g10157(.A(new_n10542_), .B(new_n1283_), .Y(new_n10543_));
  NOR2  g10158(.A(new_n10543_), .B(new_n1287_), .Y(new_n10544_));
  NOR2  g10159(.A(new_n10544_), .B(new_n1291_), .Y(new_n10545_));
  NOR2  g10160(.A(new_n10545_), .B(new_n1295_), .Y(new_n10546_));
  NOR2  g10161(.A(new_n10546_), .B(new_n1299_), .Y(new_n10547_));
  NOR2  g10162(.A(new_n10547_), .B(new_n1303_), .Y(new_n10548_));
  NOR2  g10163(.A(new_n10548_), .B(new_n1307_), .Y(new_n10549_));
  NOR2  g10164(.A(new_n10549_), .B(new_n1311_), .Y(new_n10550_));
  NOR2  g10165(.A(new_n10550_), .B(new_n1315_), .Y(new_n10551_));
  NOR2  g10166(.A(new_n10551_), .B(new_n1319_), .Y(new_n10552_));
  NOR2  g10167(.A(new_n10552_), .B(new_n1323_), .Y(new_n10553_));
  NOR2  g10168(.A(new_n10553_), .B(new_n1327_), .Y(new_n10554_));
  NOR2  g10169(.A(new_n10554_), .B(new_n1331_), .Y(new_n10555_));
  NOR2  g10170(.A(new_n10555_), .B(new_n1335_), .Y(new_n10556_));
  NOR2  g10171(.A(new_n10556_), .B(new_n1339_), .Y(new_n10557_));
  NOR2  g10172(.A(new_n10557_), .B(new_n1343_), .Y(new_n10558_));
  NOR2  g10173(.A(new_n10558_), .B(new_n1347_), .Y(new_n10559_));
  NOR2  g10174(.A(new_n10559_), .B(new_n1351_), .Y(new_n10560_));
  NOR2  g10175(.A(new_n10560_), .B(new_n1355_), .Y(new_n10561_));
  NOR2  g10176(.A(new_n10561_), .B(new_n1359_), .Y(new_n10562_));
  NOR2  g10177(.A(new_n10562_), .B(new_n1363_), .Y(new_n10563_));
  NOR2  g10178(.A(new_n10563_), .B(new_n1367_), .Y(new_n10564_));
  NOR2  g10179(.A(new_n10564_), .B(new_n1371_), .Y(new_n10565_));
  NOR2  g10180(.A(new_n10565_), .B(new_n1375_), .Y(new_n10566_));
  NOR2  g10181(.A(new_n10566_), .B(new_n1379_), .Y(new_n10567_));
  NOR2  g10182(.A(new_n10567_), .B(new_n1383_), .Y(new_n10568_));
  NOR2  g10183(.A(new_n10568_), .B(new_n1387_), .Y(new_n10569_));
  NOR2  g10184(.A(new_n10569_), .B(new_n1391_), .Y(new_n10570_));
  NOR2  g10185(.A(new_n10570_), .B(new_n1395_), .Y(new_n10571_));
  NOR2  g10186(.A(new_n10571_), .B(new_n1399_), .Y(new_n10572_));
  NOR2  g10187(.A(new_n10572_), .B(new_n1403_), .Y(new_n10573_));
  NOR2  g10188(.A(new_n10573_), .B(new_n1407_), .Y(new_n10574_));
  NOR2  g10189(.A(new_n10574_), .B(new_n1411_), .Y(new_n10575_));
  NOR2  g10190(.A(new_n10575_), .B(new_n1415_), .Y(new_n10576_));
  NOR2  g10191(.A(new_n10576_), .B(new_n1419_), .Y(new_n10577_));
  NOR2  g10192(.A(new_n10577_), .B(new_n1423_), .Y(new_n10578_));
  NOR2  g10193(.A(new_n10578_), .B(new_n1427_), .Y(new_n10579_));
  NOR2  g10194(.A(new_n10579_), .B(new_n1431_), .Y(new_n10580_));
  NOR2  g10195(.A(new_n10580_), .B(new_n1435_), .Y(new_n10581_));
  NOR2  g10196(.A(new_n10581_), .B(new_n1439_), .Y(new_n10582_));
  NOR2  g10197(.A(new_n10582_), .B(new_n1443_), .Y(new_n10583_));
  NOR2  g10198(.A(new_n10583_), .B(new_n1447_), .Y(new_n10584_));
  NOR2  g10199(.A(new_n10584_), .B(new_n1451_), .Y(new_n10585_));
  NOR2  g10200(.A(new_n10585_), .B(new_n1455_), .Y(new_n10586_));
  NOR2  g10201(.A(new_n10586_), .B(new_n1459_), .Y(new_n10587_));
  NOR2  g10202(.A(new_n10587_), .B(new_n1463_), .Y(new_n10588_));
  NAND2 g10203(.A(new_n1465_), .B(\req[106] ), .Y(new_n10589_));
  NOR2  g10204(.A(new_n10589_), .B(new_n10588_), .Y(\grant[106] ));
  INV   g10205(.A(new_n1474_), .Y(new_n10591_));
  NOR2  g10206(.A(new_n10591_), .B(new_n745_), .Y(new_n10592_));
  NOR2  g10207(.A(new_n10592_), .B(new_n1479_), .Y(new_n10593_));
  NOR2  g10208(.A(new_n10593_), .B(new_n1483_), .Y(new_n10594_));
  NOR2  g10209(.A(new_n10594_), .B(new_n1487_), .Y(new_n10595_));
  NOR2  g10210(.A(new_n10595_), .B(new_n1491_), .Y(new_n10596_));
  NOR2  g10211(.A(new_n10596_), .B(new_n1495_), .Y(new_n10597_));
  NOR2  g10212(.A(new_n10597_), .B(new_n1499_), .Y(new_n10598_));
  NOR2  g10213(.A(new_n10598_), .B(new_n1503_), .Y(new_n10599_));
  NOR2  g10214(.A(new_n10599_), .B(new_n1507_), .Y(new_n10600_));
  NOR2  g10215(.A(new_n10600_), .B(new_n1511_), .Y(new_n10601_));
  NOR2  g10216(.A(new_n10601_), .B(new_n1515_), .Y(new_n10602_));
  NOR2  g10217(.A(new_n10602_), .B(new_n1519_), .Y(new_n10603_));
  NOR2  g10218(.A(new_n10603_), .B(new_n1523_), .Y(new_n10604_));
  NOR2  g10219(.A(new_n10604_), .B(new_n1527_), .Y(new_n10605_));
  NOR2  g10220(.A(new_n10605_), .B(new_n1797_), .Y(new_n10606_));
  NOR2  g10221(.A(new_n10606_), .B(new_n396_), .Y(new_n10607_));
  NOR2  g10222(.A(new_n10607_), .B(new_n400_), .Y(new_n10608_));
  NOR2  g10223(.A(new_n10608_), .B(new_n406_), .Y(new_n10609_));
  NOR2  g10224(.A(new_n10609_), .B(new_n410_), .Y(new_n10610_));
  NOR2  g10225(.A(new_n10610_), .B(new_n416_), .Y(new_n10611_));
  NOR2  g10226(.A(new_n10611_), .B(new_n420_), .Y(new_n10612_));
  NOR2  g10227(.A(new_n10612_), .B(new_n426_), .Y(new_n10613_));
  NOR2  g10228(.A(new_n10613_), .B(new_n430_), .Y(new_n10614_));
  NOR2  g10229(.A(new_n10614_), .B(new_n436_), .Y(new_n10615_));
  NOR2  g10230(.A(new_n10615_), .B(new_n440_), .Y(new_n10616_));
  NOR2  g10231(.A(new_n10616_), .B(new_n446_), .Y(new_n10617_));
  NOR2  g10232(.A(new_n10617_), .B(new_n450_), .Y(new_n10618_));
  NOR2  g10233(.A(new_n10618_), .B(new_n456_), .Y(new_n10619_));
  NOR2  g10234(.A(new_n10619_), .B(new_n460_), .Y(new_n10620_));
  NOR2  g10235(.A(new_n10620_), .B(new_n466_), .Y(new_n10621_));
  NOR2  g10236(.A(new_n10621_), .B(new_n470_), .Y(new_n10622_));
  NOR2  g10237(.A(new_n10622_), .B(new_n476_), .Y(new_n10623_));
  NOR2  g10238(.A(new_n10623_), .B(new_n480_), .Y(new_n10624_));
  NOR2  g10239(.A(new_n10624_), .B(new_n486_), .Y(new_n10625_));
  NOR2  g10240(.A(new_n10625_), .B(new_n490_), .Y(new_n10626_));
  NOR2  g10241(.A(new_n10626_), .B(new_n496_), .Y(new_n10627_));
  NOR2  g10242(.A(new_n10627_), .B(new_n500_), .Y(new_n10628_));
  NOR2  g10243(.A(new_n10628_), .B(new_n506_), .Y(new_n10629_));
  NOR2  g10244(.A(new_n10629_), .B(new_n510_), .Y(new_n10630_));
  NOR2  g10245(.A(new_n10630_), .B(new_n516_), .Y(new_n10631_));
  NOR2  g10246(.A(new_n10631_), .B(new_n520_), .Y(new_n10632_));
  NOR2  g10247(.A(new_n10632_), .B(new_n526_), .Y(new_n10633_));
  NOR2  g10248(.A(new_n10633_), .B(new_n530_), .Y(new_n10634_));
  NOR2  g10249(.A(new_n10634_), .B(new_n536_), .Y(new_n10635_));
  NOR2  g10250(.A(new_n10635_), .B(new_n540_), .Y(new_n10636_));
  NOR2  g10251(.A(new_n10636_), .B(new_n546_), .Y(new_n10637_));
  NOR2  g10252(.A(new_n10637_), .B(new_n550_), .Y(new_n10638_));
  NOR2  g10253(.A(new_n10638_), .B(new_n556_), .Y(new_n10639_));
  NOR2  g10254(.A(new_n10639_), .B(new_n560_), .Y(new_n10640_));
  NOR2  g10255(.A(new_n10640_), .B(new_n566_), .Y(new_n10641_));
  NOR2  g10256(.A(new_n10641_), .B(new_n570_), .Y(new_n10642_));
  NOR2  g10257(.A(new_n10642_), .B(new_n576_), .Y(new_n10643_));
  NOR2  g10258(.A(new_n10643_), .B(new_n580_), .Y(new_n10644_));
  NOR2  g10259(.A(new_n10644_), .B(new_n586_), .Y(new_n10645_));
  NOR2  g10260(.A(new_n10645_), .B(new_n590_), .Y(new_n10646_));
  NOR2  g10261(.A(new_n10646_), .B(new_n596_), .Y(new_n10647_));
  NOR2  g10262(.A(new_n10647_), .B(new_n600_), .Y(new_n10648_));
  NOR2  g10263(.A(new_n10648_), .B(new_n606_), .Y(new_n10649_));
  NOR2  g10264(.A(new_n10649_), .B(new_n610_), .Y(new_n10650_));
  NOR2  g10265(.A(new_n10650_), .B(new_n616_), .Y(new_n10651_));
  NOR2  g10266(.A(new_n10651_), .B(new_n620_), .Y(new_n10652_));
  NOR2  g10267(.A(new_n10652_), .B(new_n626_), .Y(new_n10653_));
  NOR2  g10268(.A(new_n10653_), .B(new_n630_), .Y(new_n10654_));
  NOR2  g10269(.A(new_n10654_), .B(new_n636_), .Y(new_n10655_));
  NOR2  g10270(.A(new_n10655_), .B(new_n640_), .Y(new_n10656_));
  NOR2  g10271(.A(new_n10656_), .B(new_n646_), .Y(new_n10657_));
  NOR2  g10272(.A(new_n10657_), .B(new_n650_), .Y(new_n10658_));
  NOR2  g10273(.A(new_n10658_), .B(new_n656_), .Y(new_n10659_));
  NOR2  g10274(.A(new_n10659_), .B(new_n660_), .Y(new_n10660_));
  NOR2  g10275(.A(new_n10660_), .B(new_n666_), .Y(new_n10661_));
  NOR2  g10276(.A(new_n10661_), .B(new_n670_), .Y(new_n10662_));
  NOR2  g10277(.A(new_n10662_), .B(new_n676_), .Y(new_n10663_));
  NOR2  g10278(.A(new_n10663_), .B(new_n680_), .Y(new_n10664_));
  NOR2  g10279(.A(new_n10664_), .B(new_n686_), .Y(new_n10665_));
  NOR2  g10280(.A(new_n10665_), .B(new_n690_), .Y(new_n10666_));
  NOR2  g10281(.A(new_n10666_), .B(new_n696_), .Y(new_n10667_));
  NOR2  g10282(.A(new_n10667_), .B(new_n700_), .Y(new_n10668_));
  NOR2  g10283(.A(new_n10668_), .B(new_n706_), .Y(new_n10669_));
  NOR2  g10284(.A(new_n10669_), .B(new_n710_), .Y(new_n10670_));
  NOR2  g10285(.A(new_n10670_), .B(new_n716_), .Y(new_n10671_));
  NOR2  g10286(.A(new_n10671_), .B(new_n720_), .Y(new_n10672_));
  NOR2  g10287(.A(new_n10672_), .B(new_n726_), .Y(new_n10673_));
  NOR2  g10288(.A(new_n10673_), .B(new_n730_), .Y(new_n10674_));
  NOR2  g10289(.A(new_n10674_), .B(new_n736_), .Y(new_n10675_));
  NAND2 g10290(.A(new_n738_), .B(\req[107] ), .Y(new_n10676_));
  NOR2  g10291(.A(new_n10676_), .B(new_n10675_), .Y(\grant[107] ));
  INV   g10292(.A(new_n749_), .Y(new_n10678_));
  NOR2  g10293(.A(new_n1134_), .B(new_n10678_), .Y(new_n10679_));
  NOR2  g10294(.A(new_n10679_), .B(new_n756_), .Y(new_n10680_));
  NOR2  g10295(.A(new_n10680_), .B(new_n760_), .Y(new_n10681_));
  NOR2  g10296(.A(new_n10681_), .B(new_n766_), .Y(new_n10682_));
  NOR2  g10297(.A(new_n10682_), .B(new_n770_), .Y(new_n10683_));
  NOR2  g10298(.A(new_n10683_), .B(new_n776_), .Y(new_n10684_));
  NOR2  g10299(.A(new_n10684_), .B(new_n780_), .Y(new_n10685_));
  NOR2  g10300(.A(new_n10685_), .B(new_n786_), .Y(new_n10686_));
  NOR2  g10301(.A(new_n10686_), .B(new_n790_), .Y(new_n10687_));
  NOR2  g10302(.A(new_n10687_), .B(new_n796_), .Y(new_n10688_));
  NOR2  g10303(.A(new_n10688_), .B(new_n800_), .Y(new_n10689_));
  NOR2  g10304(.A(new_n10689_), .B(new_n806_), .Y(new_n10690_));
  NOR2  g10305(.A(new_n10690_), .B(new_n1616_), .Y(new_n10691_));
  NOR2  g10306(.A(new_n10691_), .B(new_n1618_), .Y(new_n10692_));
  NOR2  g10307(.A(new_n10692_), .B(new_n1885_), .Y(new_n10693_));
  NOR2  g10308(.A(new_n10693_), .B(new_n820_), .Y(new_n10694_));
  NOR2  g10309(.A(new_n10694_), .B(new_n824_), .Y(new_n10695_));
  NOR2  g10310(.A(new_n10695_), .B(new_n829_), .Y(new_n10696_));
  NOR2  g10311(.A(new_n10696_), .B(new_n833_), .Y(new_n10697_));
  NOR2  g10312(.A(new_n10697_), .B(new_n838_), .Y(new_n10698_));
  NOR2  g10313(.A(new_n10698_), .B(new_n842_), .Y(new_n10699_));
  NOR2  g10314(.A(new_n10699_), .B(new_n847_), .Y(new_n10700_));
  NOR2  g10315(.A(new_n10700_), .B(new_n851_), .Y(new_n10701_));
  NOR2  g10316(.A(new_n10701_), .B(new_n856_), .Y(new_n10702_));
  NOR2  g10317(.A(new_n10702_), .B(new_n860_), .Y(new_n10703_));
  NOR2  g10318(.A(new_n10703_), .B(new_n865_), .Y(new_n10704_));
  NOR2  g10319(.A(new_n10704_), .B(new_n869_), .Y(new_n10705_));
  NOR2  g10320(.A(new_n10705_), .B(new_n874_), .Y(new_n10706_));
  NOR2  g10321(.A(new_n10706_), .B(new_n878_), .Y(new_n10707_));
  NOR2  g10322(.A(new_n10707_), .B(new_n883_), .Y(new_n10708_));
  NOR2  g10323(.A(new_n10708_), .B(new_n887_), .Y(new_n10709_));
  NOR2  g10324(.A(new_n10709_), .B(new_n892_), .Y(new_n10710_));
  NOR2  g10325(.A(new_n10710_), .B(new_n896_), .Y(new_n10711_));
  NOR2  g10326(.A(new_n10711_), .B(new_n901_), .Y(new_n10712_));
  NOR2  g10327(.A(new_n10712_), .B(new_n905_), .Y(new_n10713_));
  NOR2  g10328(.A(new_n10713_), .B(new_n910_), .Y(new_n10714_));
  NOR2  g10329(.A(new_n10714_), .B(new_n914_), .Y(new_n10715_));
  NOR2  g10330(.A(new_n10715_), .B(new_n919_), .Y(new_n10716_));
  NOR2  g10331(.A(new_n10716_), .B(new_n923_), .Y(new_n10717_));
  NOR2  g10332(.A(new_n10717_), .B(new_n928_), .Y(new_n10718_));
  NOR2  g10333(.A(new_n10718_), .B(new_n932_), .Y(new_n10719_));
  NOR2  g10334(.A(new_n10719_), .B(new_n937_), .Y(new_n10720_));
  NOR2  g10335(.A(new_n10720_), .B(new_n941_), .Y(new_n10721_));
  NOR2  g10336(.A(new_n10721_), .B(new_n946_), .Y(new_n10722_));
  NOR2  g10337(.A(new_n10722_), .B(new_n950_), .Y(new_n10723_));
  NOR2  g10338(.A(new_n10723_), .B(new_n955_), .Y(new_n10724_));
  NOR2  g10339(.A(new_n10724_), .B(new_n959_), .Y(new_n10725_));
  NOR2  g10340(.A(new_n10725_), .B(new_n964_), .Y(new_n10726_));
  NOR2  g10341(.A(new_n10726_), .B(new_n968_), .Y(new_n10727_));
  NOR2  g10342(.A(new_n10727_), .B(new_n973_), .Y(new_n10728_));
  NOR2  g10343(.A(new_n10728_), .B(new_n977_), .Y(new_n10729_));
  NOR2  g10344(.A(new_n10729_), .B(new_n982_), .Y(new_n10730_));
  NOR2  g10345(.A(new_n10730_), .B(new_n986_), .Y(new_n10731_));
  NOR2  g10346(.A(new_n10731_), .B(new_n991_), .Y(new_n10732_));
  NOR2  g10347(.A(new_n10732_), .B(new_n995_), .Y(new_n10733_));
  NOR2  g10348(.A(new_n10733_), .B(new_n1000_), .Y(new_n10734_));
  NOR2  g10349(.A(new_n10734_), .B(new_n1004_), .Y(new_n10735_));
  NOR2  g10350(.A(new_n10735_), .B(new_n1009_), .Y(new_n10736_));
  NOR2  g10351(.A(new_n10736_), .B(new_n1013_), .Y(new_n10737_));
  NOR2  g10352(.A(new_n10737_), .B(new_n1018_), .Y(new_n10738_));
  NOR2  g10353(.A(new_n10738_), .B(new_n1022_), .Y(new_n10739_));
  NOR2  g10354(.A(new_n10739_), .B(new_n1027_), .Y(new_n10740_));
  NOR2  g10355(.A(new_n10740_), .B(new_n1031_), .Y(new_n10741_));
  NOR2  g10356(.A(new_n10741_), .B(new_n1036_), .Y(new_n10742_));
  NOR2  g10357(.A(new_n10742_), .B(new_n1040_), .Y(new_n10743_));
  NOR2  g10358(.A(new_n10743_), .B(new_n1045_), .Y(new_n10744_));
  NOR2  g10359(.A(new_n10744_), .B(new_n1049_), .Y(new_n10745_));
  NOR2  g10360(.A(new_n10745_), .B(new_n1054_), .Y(new_n10746_));
  NOR2  g10361(.A(new_n10746_), .B(new_n1058_), .Y(new_n10747_));
  NOR2  g10362(.A(new_n10747_), .B(new_n1063_), .Y(new_n10748_));
  NOR2  g10363(.A(new_n10748_), .B(new_n1067_), .Y(new_n10749_));
  NOR2  g10364(.A(new_n10749_), .B(new_n1072_), .Y(new_n10750_));
  NOR2  g10365(.A(new_n10750_), .B(new_n1076_), .Y(new_n10751_));
  NOR2  g10366(.A(new_n10751_), .B(new_n1081_), .Y(new_n10752_));
  NOR2  g10367(.A(new_n10752_), .B(new_n1085_), .Y(new_n10753_));
  NOR2  g10368(.A(new_n10753_), .B(new_n1090_), .Y(new_n10754_));
  NOR2  g10369(.A(new_n10754_), .B(new_n1094_), .Y(new_n10755_));
  NOR2  g10370(.A(new_n10755_), .B(new_n1099_), .Y(new_n10756_));
  NOR2  g10371(.A(new_n10756_), .B(new_n1103_), .Y(new_n10757_));
  NOR2  g10372(.A(new_n10757_), .B(new_n1108_), .Y(new_n10758_));
  NOR2  g10373(.A(new_n10758_), .B(new_n1112_), .Y(new_n10759_));
  NOR2  g10374(.A(new_n10759_), .B(new_n1117_), .Y(new_n10760_));
  NOR2  g10375(.A(new_n10760_), .B(new_n1121_), .Y(new_n10761_));
  NOR2  g10376(.A(new_n10761_), .B(new_n1126_), .Y(new_n10762_));
  NAND2 g10377(.A(new_n1128_), .B(\req[108] ), .Y(new_n10763_));
  NOR2  g10378(.A(new_n10763_), .B(new_n10762_), .Y(\grant[108] ));
  INV   g10379(.A(new_n1138_), .Y(new_n10765_));
  NOR2  g10380(.A(new_n1478_), .B(new_n10765_), .Y(new_n10766_));
  NOR2  g10381(.A(new_n10766_), .B(new_n1144_), .Y(new_n10767_));
  NOR2  g10382(.A(new_n10767_), .B(new_n1148_), .Y(new_n10768_));
  NOR2  g10383(.A(new_n10768_), .B(new_n1153_), .Y(new_n10769_));
  NOR2  g10384(.A(new_n10769_), .B(new_n1157_), .Y(new_n10770_));
  NOR2  g10385(.A(new_n10770_), .B(new_n1162_), .Y(new_n10771_));
  NOR2  g10386(.A(new_n10771_), .B(new_n1166_), .Y(new_n10772_));
  NOR2  g10387(.A(new_n10772_), .B(new_n1171_), .Y(new_n10773_));
  NOR2  g10388(.A(new_n10773_), .B(new_n1175_), .Y(new_n10774_));
  NOR2  g10389(.A(new_n10774_), .B(new_n1180_), .Y(new_n10775_));
  NOR2  g10390(.A(new_n10775_), .B(new_n1184_), .Y(new_n10776_));
  NOR2  g10391(.A(new_n10776_), .B(new_n1189_), .Y(new_n10777_));
  NOR2  g10392(.A(new_n10777_), .B(new_n1707_), .Y(new_n10778_));
  NOR2  g10393(.A(new_n10778_), .B(new_n1709_), .Y(new_n10779_));
  NOR2  g10394(.A(new_n10779_), .B(new_n1973_), .Y(new_n10780_));
  NOR2  g10395(.A(new_n10780_), .B(new_n1199_), .Y(new_n10781_));
  NOR2  g10396(.A(new_n10781_), .B(new_n1203_), .Y(new_n10782_));
  NOR2  g10397(.A(new_n10782_), .B(new_n1207_), .Y(new_n10783_));
  NOR2  g10398(.A(new_n10783_), .B(new_n1211_), .Y(new_n10784_));
  NOR2  g10399(.A(new_n10784_), .B(new_n1215_), .Y(new_n10785_));
  NOR2  g10400(.A(new_n10785_), .B(new_n1219_), .Y(new_n10786_));
  NOR2  g10401(.A(new_n10786_), .B(new_n1223_), .Y(new_n10787_));
  NOR2  g10402(.A(new_n10787_), .B(new_n1227_), .Y(new_n10788_));
  NOR2  g10403(.A(new_n10788_), .B(new_n1231_), .Y(new_n10789_));
  NOR2  g10404(.A(new_n10789_), .B(new_n1235_), .Y(new_n10790_));
  NOR2  g10405(.A(new_n10790_), .B(new_n1239_), .Y(new_n10791_));
  NOR2  g10406(.A(new_n10791_), .B(new_n1243_), .Y(new_n10792_));
  NOR2  g10407(.A(new_n10792_), .B(new_n1247_), .Y(new_n10793_));
  NOR2  g10408(.A(new_n10793_), .B(new_n1251_), .Y(new_n10794_));
  NOR2  g10409(.A(new_n10794_), .B(new_n1255_), .Y(new_n10795_));
  NOR2  g10410(.A(new_n10795_), .B(new_n1259_), .Y(new_n10796_));
  NOR2  g10411(.A(new_n10796_), .B(new_n1263_), .Y(new_n10797_));
  NOR2  g10412(.A(new_n10797_), .B(new_n1267_), .Y(new_n10798_));
  NOR2  g10413(.A(new_n10798_), .B(new_n1271_), .Y(new_n10799_));
  NOR2  g10414(.A(new_n10799_), .B(new_n1275_), .Y(new_n10800_));
  NOR2  g10415(.A(new_n10800_), .B(new_n1279_), .Y(new_n10801_));
  NOR2  g10416(.A(new_n10801_), .B(new_n1283_), .Y(new_n10802_));
  NOR2  g10417(.A(new_n10802_), .B(new_n1287_), .Y(new_n10803_));
  NOR2  g10418(.A(new_n10803_), .B(new_n1291_), .Y(new_n10804_));
  NOR2  g10419(.A(new_n10804_), .B(new_n1295_), .Y(new_n10805_));
  NOR2  g10420(.A(new_n10805_), .B(new_n1299_), .Y(new_n10806_));
  NOR2  g10421(.A(new_n10806_), .B(new_n1303_), .Y(new_n10807_));
  NOR2  g10422(.A(new_n10807_), .B(new_n1307_), .Y(new_n10808_));
  NOR2  g10423(.A(new_n10808_), .B(new_n1311_), .Y(new_n10809_));
  NOR2  g10424(.A(new_n10809_), .B(new_n1315_), .Y(new_n10810_));
  NOR2  g10425(.A(new_n10810_), .B(new_n1319_), .Y(new_n10811_));
  NOR2  g10426(.A(new_n10811_), .B(new_n1323_), .Y(new_n10812_));
  NOR2  g10427(.A(new_n10812_), .B(new_n1327_), .Y(new_n10813_));
  NOR2  g10428(.A(new_n10813_), .B(new_n1331_), .Y(new_n10814_));
  NOR2  g10429(.A(new_n10814_), .B(new_n1335_), .Y(new_n10815_));
  NOR2  g10430(.A(new_n10815_), .B(new_n1339_), .Y(new_n10816_));
  NOR2  g10431(.A(new_n10816_), .B(new_n1343_), .Y(new_n10817_));
  NOR2  g10432(.A(new_n10817_), .B(new_n1347_), .Y(new_n10818_));
  NOR2  g10433(.A(new_n10818_), .B(new_n1351_), .Y(new_n10819_));
  NOR2  g10434(.A(new_n10819_), .B(new_n1355_), .Y(new_n10820_));
  NOR2  g10435(.A(new_n10820_), .B(new_n1359_), .Y(new_n10821_));
  NOR2  g10436(.A(new_n10821_), .B(new_n1363_), .Y(new_n10822_));
  NOR2  g10437(.A(new_n10822_), .B(new_n1367_), .Y(new_n10823_));
  NOR2  g10438(.A(new_n10823_), .B(new_n1371_), .Y(new_n10824_));
  NOR2  g10439(.A(new_n10824_), .B(new_n1375_), .Y(new_n10825_));
  NOR2  g10440(.A(new_n10825_), .B(new_n1379_), .Y(new_n10826_));
  NOR2  g10441(.A(new_n10826_), .B(new_n1383_), .Y(new_n10827_));
  NOR2  g10442(.A(new_n10827_), .B(new_n1387_), .Y(new_n10828_));
  NOR2  g10443(.A(new_n10828_), .B(new_n1391_), .Y(new_n10829_));
  NOR2  g10444(.A(new_n10829_), .B(new_n1395_), .Y(new_n10830_));
  NOR2  g10445(.A(new_n10830_), .B(new_n1399_), .Y(new_n10831_));
  NOR2  g10446(.A(new_n10831_), .B(new_n1403_), .Y(new_n10832_));
  NOR2  g10447(.A(new_n10832_), .B(new_n1407_), .Y(new_n10833_));
  NOR2  g10448(.A(new_n10833_), .B(new_n1411_), .Y(new_n10834_));
  NOR2  g10449(.A(new_n10834_), .B(new_n1415_), .Y(new_n10835_));
  NOR2  g10450(.A(new_n10835_), .B(new_n1419_), .Y(new_n10836_));
  NOR2  g10451(.A(new_n10836_), .B(new_n1423_), .Y(new_n10837_));
  NOR2  g10452(.A(new_n10837_), .B(new_n1427_), .Y(new_n10838_));
  NOR2  g10453(.A(new_n10838_), .B(new_n1431_), .Y(new_n10839_));
  NOR2  g10454(.A(new_n10839_), .B(new_n1435_), .Y(new_n10840_));
  NOR2  g10455(.A(new_n10840_), .B(new_n1439_), .Y(new_n10841_));
  NOR2  g10456(.A(new_n10841_), .B(new_n1443_), .Y(new_n10842_));
  NOR2  g10457(.A(new_n10842_), .B(new_n1447_), .Y(new_n10843_));
  NOR2  g10458(.A(new_n10843_), .B(new_n1451_), .Y(new_n10844_));
  NOR2  g10459(.A(new_n10844_), .B(new_n1455_), .Y(new_n10845_));
  NOR2  g10460(.A(new_n10845_), .B(new_n1459_), .Y(new_n10846_));
  NOR2  g10461(.A(new_n10846_), .B(new_n1463_), .Y(new_n10847_));
  NOR2  g10462(.A(new_n10847_), .B(new_n1467_), .Y(new_n10848_));
  NOR2  g10463(.A(new_n10848_), .B(new_n1471_), .Y(new_n10849_));
  NAND2 g10464(.A(new_n1473_), .B(\req[109] ), .Y(new_n10850_));
  NOR2  g10465(.A(new_n10850_), .B(new_n10849_), .Y(\grant[109] ));
  INV   g10466(.A(new_n1482_), .Y(new_n10852_));
  NOR2  g10467(.A(new_n10852_), .B(new_n755_), .Y(new_n10853_));
  NOR2  g10468(.A(new_n10853_), .B(new_n1487_), .Y(new_n10854_));
  NOR2  g10469(.A(new_n10854_), .B(new_n1491_), .Y(new_n10855_));
  NOR2  g10470(.A(new_n10855_), .B(new_n1495_), .Y(new_n10856_));
  NOR2  g10471(.A(new_n10856_), .B(new_n1499_), .Y(new_n10857_));
  NOR2  g10472(.A(new_n10857_), .B(new_n1503_), .Y(new_n10858_));
  NOR2  g10473(.A(new_n10858_), .B(new_n1507_), .Y(new_n10859_));
  NOR2  g10474(.A(new_n10859_), .B(new_n1511_), .Y(new_n10860_));
  NOR2  g10475(.A(new_n10860_), .B(new_n1515_), .Y(new_n10861_));
  NOR2  g10476(.A(new_n10861_), .B(new_n1519_), .Y(new_n10862_));
  NOR2  g10477(.A(new_n10862_), .B(new_n1523_), .Y(new_n10863_));
  NOR2  g10478(.A(new_n10863_), .B(new_n1527_), .Y(new_n10864_));
  NOR2  g10479(.A(new_n10864_), .B(new_n1797_), .Y(new_n10865_));
  NOR2  g10480(.A(new_n10865_), .B(new_n396_), .Y(new_n10866_));
  NOR2  g10481(.A(new_n10866_), .B(new_n400_), .Y(new_n10867_));
  NOR2  g10482(.A(new_n10867_), .B(new_n406_), .Y(new_n10868_));
  NOR2  g10483(.A(new_n10868_), .B(new_n410_), .Y(new_n10869_));
  NOR2  g10484(.A(new_n10869_), .B(new_n416_), .Y(new_n10870_));
  NOR2  g10485(.A(new_n10870_), .B(new_n420_), .Y(new_n10871_));
  NOR2  g10486(.A(new_n10871_), .B(new_n426_), .Y(new_n10872_));
  NOR2  g10487(.A(new_n10872_), .B(new_n430_), .Y(new_n10873_));
  NOR2  g10488(.A(new_n10873_), .B(new_n436_), .Y(new_n10874_));
  NOR2  g10489(.A(new_n10874_), .B(new_n440_), .Y(new_n10875_));
  NOR2  g10490(.A(new_n10875_), .B(new_n446_), .Y(new_n10876_));
  NOR2  g10491(.A(new_n10876_), .B(new_n450_), .Y(new_n10877_));
  NOR2  g10492(.A(new_n10877_), .B(new_n456_), .Y(new_n10878_));
  NOR2  g10493(.A(new_n10878_), .B(new_n460_), .Y(new_n10879_));
  NOR2  g10494(.A(new_n10879_), .B(new_n466_), .Y(new_n10880_));
  NOR2  g10495(.A(new_n10880_), .B(new_n470_), .Y(new_n10881_));
  NOR2  g10496(.A(new_n10881_), .B(new_n476_), .Y(new_n10882_));
  NOR2  g10497(.A(new_n10882_), .B(new_n480_), .Y(new_n10883_));
  NOR2  g10498(.A(new_n10883_), .B(new_n486_), .Y(new_n10884_));
  NOR2  g10499(.A(new_n10884_), .B(new_n490_), .Y(new_n10885_));
  NOR2  g10500(.A(new_n10885_), .B(new_n496_), .Y(new_n10886_));
  NOR2  g10501(.A(new_n10886_), .B(new_n500_), .Y(new_n10887_));
  NOR2  g10502(.A(new_n10887_), .B(new_n506_), .Y(new_n10888_));
  NOR2  g10503(.A(new_n10888_), .B(new_n510_), .Y(new_n10889_));
  NOR2  g10504(.A(new_n10889_), .B(new_n516_), .Y(new_n10890_));
  NOR2  g10505(.A(new_n10890_), .B(new_n520_), .Y(new_n10891_));
  NOR2  g10506(.A(new_n10891_), .B(new_n526_), .Y(new_n10892_));
  NOR2  g10507(.A(new_n10892_), .B(new_n530_), .Y(new_n10893_));
  NOR2  g10508(.A(new_n10893_), .B(new_n536_), .Y(new_n10894_));
  NOR2  g10509(.A(new_n10894_), .B(new_n540_), .Y(new_n10895_));
  NOR2  g10510(.A(new_n10895_), .B(new_n546_), .Y(new_n10896_));
  NOR2  g10511(.A(new_n10896_), .B(new_n550_), .Y(new_n10897_));
  NOR2  g10512(.A(new_n10897_), .B(new_n556_), .Y(new_n10898_));
  NOR2  g10513(.A(new_n10898_), .B(new_n560_), .Y(new_n10899_));
  NOR2  g10514(.A(new_n10899_), .B(new_n566_), .Y(new_n10900_));
  NOR2  g10515(.A(new_n10900_), .B(new_n570_), .Y(new_n10901_));
  NOR2  g10516(.A(new_n10901_), .B(new_n576_), .Y(new_n10902_));
  NOR2  g10517(.A(new_n10902_), .B(new_n580_), .Y(new_n10903_));
  NOR2  g10518(.A(new_n10903_), .B(new_n586_), .Y(new_n10904_));
  NOR2  g10519(.A(new_n10904_), .B(new_n590_), .Y(new_n10905_));
  NOR2  g10520(.A(new_n10905_), .B(new_n596_), .Y(new_n10906_));
  NOR2  g10521(.A(new_n10906_), .B(new_n600_), .Y(new_n10907_));
  NOR2  g10522(.A(new_n10907_), .B(new_n606_), .Y(new_n10908_));
  NOR2  g10523(.A(new_n10908_), .B(new_n610_), .Y(new_n10909_));
  NOR2  g10524(.A(new_n10909_), .B(new_n616_), .Y(new_n10910_));
  NOR2  g10525(.A(new_n10910_), .B(new_n620_), .Y(new_n10911_));
  NOR2  g10526(.A(new_n10911_), .B(new_n626_), .Y(new_n10912_));
  NOR2  g10527(.A(new_n10912_), .B(new_n630_), .Y(new_n10913_));
  NOR2  g10528(.A(new_n10913_), .B(new_n636_), .Y(new_n10914_));
  NOR2  g10529(.A(new_n10914_), .B(new_n640_), .Y(new_n10915_));
  NOR2  g10530(.A(new_n10915_), .B(new_n646_), .Y(new_n10916_));
  NOR2  g10531(.A(new_n10916_), .B(new_n650_), .Y(new_n10917_));
  NOR2  g10532(.A(new_n10917_), .B(new_n656_), .Y(new_n10918_));
  NOR2  g10533(.A(new_n10918_), .B(new_n660_), .Y(new_n10919_));
  NOR2  g10534(.A(new_n10919_), .B(new_n666_), .Y(new_n10920_));
  NOR2  g10535(.A(new_n10920_), .B(new_n670_), .Y(new_n10921_));
  NOR2  g10536(.A(new_n10921_), .B(new_n676_), .Y(new_n10922_));
  NOR2  g10537(.A(new_n10922_), .B(new_n680_), .Y(new_n10923_));
  NOR2  g10538(.A(new_n10923_), .B(new_n686_), .Y(new_n10924_));
  NOR2  g10539(.A(new_n10924_), .B(new_n690_), .Y(new_n10925_));
  NOR2  g10540(.A(new_n10925_), .B(new_n696_), .Y(new_n10926_));
  NOR2  g10541(.A(new_n10926_), .B(new_n700_), .Y(new_n10927_));
  NOR2  g10542(.A(new_n10927_), .B(new_n706_), .Y(new_n10928_));
  NOR2  g10543(.A(new_n10928_), .B(new_n710_), .Y(new_n10929_));
  NOR2  g10544(.A(new_n10929_), .B(new_n716_), .Y(new_n10930_));
  NOR2  g10545(.A(new_n10930_), .B(new_n720_), .Y(new_n10931_));
  NOR2  g10546(.A(new_n10931_), .B(new_n726_), .Y(new_n10932_));
  NOR2  g10547(.A(new_n10932_), .B(new_n730_), .Y(new_n10933_));
  NOR2  g10548(.A(new_n10933_), .B(new_n736_), .Y(new_n10934_));
  NOR2  g10549(.A(new_n10934_), .B(new_n740_), .Y(new_n10935_));
  NOR2  g10550(.A(new_n10935_), .B(new_n746_), .Y(new_n10936_));
  NAND2 g10551(.A(new_n748_), .B(\req[110] ), .Y(new_n10937_));
  NOR2  g10552(.A(new_n10937_), .B(new_n10936_), .Y(\grant[110] ));
  INV   g10553(.A(new_n759_), .Y(new_n10939_));
  NOR2  g10554(.A(new_n1143_), .B(new_n10939_), .Y(new_n10940_));
  NOR2  g10555(.A(new_n10940_), .B(new_n766_), .Y(new_n10941_));
  NOR2  g10556(.A(new_n10941_), .B(new_n770_), .Y(new_n10942_));
  NOR2  g10557(.A(new_n10942_), .B(new_n776_), .Y(new_n10943_));
  NOR2  g10558(.A(new_n10943_), .B(new_n780_), .Y(new_n10944_));
  NOR2  g10559(.A(new_n10944_), .B(new_n786_), .Y(new_n10945_));
  NOR2  g10560(.A(new_n10945_), .B(new_n790_), .Y(new_n10946_));
  NOR2  g10561(.A(new_n10946_), .B(new_n796_), .Y(new_n10947_));
  NOR2  g10562(.A(new_n10947_), .B(new_n800_), .Y(new_n10948_));
  NOR2  g10563(.A(new_n10948_), .B(new_n806_), .Y(new_n10949_));
  NOR2  g10564(.A(new_n10949_), .B(new_n1616_), .Y(new_n10950_));
  NOR2  g10565(.A(new_n10950_), .B(new_n1618_), .Y(new_n10951_));
  NOR2  g10566(.A(new_n10951_), .B(new_n1885_), .Y(new_n10952_));
  NOR2  g10567(.A(new_n10952_), .B(new_n820_), .Y(new_n10953_));
  NOR2  g10568(.A(new_n10953_), .B(new_n824_), .Y(new_n10954_));
  NOR2  g10569(.A(new_n10954_), .B(new_n829_), .Y(new_n10955_));
  NOR2  g10570(.A(new_n10955_), .B(new_n833_), .Y(new_n10956_));
  NOR2  g10571(.A(new_n10956_), .B(new_n838_), .Y(new_n10957_));
  NOR2  g10572(.A(new_n10957_), .B(new_n842_), .Y(new_n10958_));
  NOR2  g10573(.A(new_n10958_), .B(new_n847_), .Y(new_n10959_));
  NOR2  g10574(.A(new_n10959_), .B(new_n851_), .Y(new_n10960_));
  NOR2  g10575(.A(new_n10960_), .B(new_n856_), .Y(new_n10961_));
  NOR2  g10576(.A(new_n10961_), .B(new_n860_), .Y(new_n10962_));
  NOR2  g10577(.A(new_n10962_), .B(new_n865_), .Y(new_n10963_));
  NOR2  g10578(.A(new_n10963_), .B(new_n869_), .Y(new_n10964_));
  NOR2  g10579(.A(new_n10964_), .B(new_n874_), .Y(new_n10965_));
  NOR2  g10580(.A(new_n10965_), .B(new_n878_), .Y(new_n10966_));
  NOR2  g10581(.A(new_n10966_), .B(new_n883_), .Y(new_n10967_));
  NOR2  g10582(.A(new_n10967_), .B(new_n887_), .Y(new_n10968_));
  NOR2  g10583(.A(new_n10968_), .B(new_n892_), .Y(new_n10969_));
  NOR2  g10584(.A(new_n10969_), .B(new_n896_), .Y(new_n10970_));
  NOR2  g10585(.A(new_n10970_), .B(new_n901_), .Y(new_n10971_));
  NOR2  g10586(.A(new_n10971_), .B(new_n905_), .Y(new_n10972_));
  NOR2  g10587(.A(new_n10972_), .B(new_n910_), .Y(new_n10973_));
  NOR2  g10588(.A(new_n10973_), .B(new_n914_), .Y(new_n10974_));
  NOR2  g10589(.A(new_n10974_), .B(new_n919_), .Y(new_n10975_));
  NOR2  g10590(.A(new_n10975_), .B(new_n923_), .Y(new_n10976_));
  NOR2  g10591(.A(new_n10976_), .B(new_n928_), .Y(new_n10977_));
  NOR2  g10592(.A(new_n10977_), .B(new_n932_), .Y(new_n10978_));
  NOR2  g10593(.A(new_n10978_), .B(new_n937_), .Y(new_n10979_));
  NOR2  g10594(.A(new_n10979_), .B(new_n941_), .Y(new_n10980_));
  NOR2  g10595(.A(new_n10980_), .B(new_n946_), .Y(new_n10981_));
  NOR2  g10596(.A(new_n10981_), .B(new_n950_), .Y(new_n10982_));
  NOR2  g10597(.A(new_n10982_), .B(new_n955_), .Y(new_n10983_));
  NOR2  g10598(.A(new_n10983_), .B(new_n959_), .Y(new_n10984_));
  NOR2  g10599(.A(new_n10984_), .B(new_n964_), .Y(new_n10985_));
  NOR2  g10600(.A(new_n10985_), .B(new_n968_), .Y(new_n10986_));
  NOR2  g10601(.A(new_n10986_), .B(new_n973_), .Y(new_n10987_));
  NOR2  g10602(.A(new_n10987_), .B(new_n977_), .Y(new_n10988_));
  NOR2  g10603(.A(new_n10988_), .B(new_n982_), .Y(new_n10989_));
  NOR2  g10604(.A(new_n10989_), .B(new_n986_), .Y(new_n10990_));
  NOR2  g10605(.A(new_n10990_), .B(new_n991_), .Y(new_n10991_));
  NOR2  g10606(.A(new_n10991_), .B(new_n995_), .Y(new_n10992_));
  NOR2  g10607(.A(new_n10992_), .B(new_n1000_), .Y(new_n10993_));
  NOR2  g10608(.A(new_n10993_), .B(new_n1004_), .Y(new_n10994_));
  NOR2  g10609(.A(new_n10994_), .B(new_n1009_), .Y(new_n10995_));
  NOR2  g10610(.A(new_n10995_), .B(new_n1013_), .Y(new_n10996_));
  NOR2  g10611(.A(new_n10996_), .B(new_n1018_), .Y(new_n10997_));
  NOR2  g10612(.A(new_n10997_), .B(new_n1022_), .Y(new_n10998_));
  NOR2  g10613(.A(new_n10998_), .B(new_n1027_), .Y(new_n10999_));
  NOR2  g10614(.A(new_n10999_), .B(new_n1031_), .Y(new_n11000_));
  NOR2  g10615(.A(new_n11000_), .B(new_n1036_), .Y(new_n11001_));
  NOR2  g10616(.A(new_n11001_), .B(new_n1040_), .Y(new_n11002_));
  NOR2  g10617(.A(new_n11002_), .B(new_n1045_), .Y(new_n11003_));
  NOR2  g10618(.A(new_n11003_), .B(new_n1049_), .Y(new_n11004_));
  NOR2  g10619(.A(new_n11004_), .B(new_n1054_), .Y(new_n11005_));
  NOR2  g10620(.A(new_n11005_), .B(new_n1058_), .Y(new_n11006_));
  NOR2  g10621(.A(new_n11006_), .B(new_n1063_), .Y(new_n11007_));
  NOR2  g10622(.A(new_n11007_), .B(new_n1067_), .Y(new_n11008_));
  NOR2  g10623(.A(new_n11008_), .B(new_n1072_), .Y(new_n11009_));
  NOR2  g10624(.A(new_n11009_), .B(new_n1076_), .Y(new_n11010_));
  NOR2  g10625(.A(new_n11010_), .B(new_n1081_), .Y(new_n11011_));
  NOR2  g10626(.A(new_n11011_), .B(new_n1085_), .Y(new_n11012_));
  NOR2  g10627(.A(new_n11012_), .B(new_n1090_), .Y(new_n11013_));
  NOR2  g10628(.A(new_n11013_), .B(new_n1094_), .Y(new_n11014_));
  NOR2  g10629(.A(new_n11014_), .B(new_n1099_), .Y(new_n11015_));
  NOR2  g10630(.A(new_n11015_), .B(new_n1103_), .Y(new_n11016_));
  NOR2  g10631(.A(new_n11016_), .B(new_n1108_), .Y(new_n11017_));
  NOR2  g10632(.A(new_n11017_), .B(new_n1112_), .Y(new_n11018_));
  NOR2  g10633(.A(new_n11018_), .B(new_n1117_), .Y(new_n11019_));
  NOR2  g10634(.A(new_n11019_), .B(new_n1121_), .Y(new_n11020_));
  NOR2  g10635(.A(new_n11020_), .B(new_n1126_), .Y(new_n11021_));
  NOR2  g10636(.A(new_n11021_), .B(new_n1130_), .Y(new_n11022_));
  NOR2  g10637(.A(new_n11022_), .B(new_n1135_), .Y(new_n11023_));
  NAND2 g10638(.A(new_n1137_), .B(\req[111] ), .Y(new_n11024_));
  NOR2  g10639(.A(new_n11024_), .B(new_n11023_), .Y(\grant[111] ));
  INV   g10640(.A(new_n1147_), .Y(new_n11026_));
  NOR2  g10641(.A(new_n1486_), .B(new_n11026_), .Y(new_n11027_));
  NOR2  g10642(.A(new_n11027_), .B(new_n1153_), .Y(new_n11028_));
  NOR2  g10643(.A(new_n11028_), .B(new_n1157_), .Y(new_n11029_));
  NOR2  g10644(.A(new_n11029_), .B(new_n1162_), .Y(new_n11030_));
  NOR2  g10645(.A(new_n11030_), .B(new_n1166_), .Y(new_n11031_));
  NOR2  g10646(.A(new_n11031_), .B(new_n1171_), .Y(new_n11032_));
  NOR2  g10647(.A(new_n11032_), .B(new_n1175_), .Y(new_n11033_));
  NOR2  g10648(.A(new_n11033_), .B(new_n1180_), .Y(new_n11034_));
  NOR2  g10649(.A(new_n11034_), .B(new_n1184_), .Y(new_n11035_));
  NOR2  g10650(.A(new_n11035_), .B(new_n1189_), .Y(new_n11036_));
  NOR2  g10651(.A(new_n11036_), .B(new_n1707_), .Y(new_n11037_));
  NOR2  g10652(.A(new_n11037_), .B(new_n1709_), .Y(new_n11038_));
  NOR2  g10653(.A(new_n11038_), .B(new_n1973_), .Y(new_n11039_));
  NOR2  g10654(.A(new_n11039_), .B(new_n1199_), .Y(new_n11040_));
  NOR2  g10655(.A(new_n11040_), .B(new_n1203_), .Y(new_n11041_));
  NOR2  g10656(.A(new_n11041_), .B(new_n1207_), .Y(new_n11042_));
  NOR2  g10657(.A(new_n11042_), .B(new_n1211_), .Y(new_n11043_));
  NOR2  g10658(.A(new_n11043_), .B(new_n1215_), .Y(new_n11044_));
  NOR2  g10659(.A(new_n11044_), .B(new_n1219_), .Y(new_n11045_));
  NOR2  g10660(.A(new_n11045_), .B(new_n1223_), .Y(new_n11046_));
  NOR2  g10661(.A(new_n11046_), .B(new_n1227_), .Y(new_n11047_));
  NOR2  g10662(.A(new_n11047_), .B(new_n1231_), .Y(new_n11048_));
  NOR2  g10663(.A(new_n11048_), .B(new_n1235_), .Y(new_n11049_));
  NOR2  g10664(.A(new_n11049_), .B(new_n1239_), .Y(new_n11050_));
  NOR2  g10665(.A(new_n11050_), .B(new_n1243_), .Y(new_n11051_));
  NOR2  g10666(.A(new_n11051_), .B(new_n1247_), .Y(new_n11052_));
  NOR2  g10667(.A(new_n11052_), .B(new_n1251_), .Y(new_n11053_));
  NOR2  g10668(.A(new_n11053_), .B(new_n1255_), .Y(new_n11054_));
  NOR2  g10669(.A(new_n11054_), .B(new_n1259_), .Y(new_n11055_));
  NOR2  g10670(.A(new_n11055_), .B(new_n1263_), .Y(new_n11056_));
  NOR2  g10671(.A(new_n11056_), .B(new_n1267_), .Y(new_n11057_));
  NOR2  g10672(.A(new_n11057_), .B(new_n1271_), .Y(new_n11058_));
  NOR2  g10673(.A(new_n11058_), .B(new_n1275_), .Y(new_n11059_));
  NOR2  g10674(.A(new_n11059_), .B(new_n1279_), .Y(new_n11060_));
  NOR2  g10675(.A(new_n11060_), .B(new_n1283_), .Y(new_n11061_));
  NOR2  g10676(.A(new_n11061_), .B(new_n1287_), .Y(new_n11062_));
  NOR2  g10677(.A(new_n11062_), .B(new_n1291_), .Y(new_n11063_));
  NOR2  g10678(.A(new_n11063_), .B(new_n1295_), .Y(new_n11064_));
  NOR2  g10679(.A(new_n11064_), .B(new_n1299_), .Y(new_n11065_));
  NOR2  g10680(.A(new_n11065_), .B(new_n1303_), .Y(new_n11066_));
  NOR2  g10681(.A(new_n11066_), .B(new_n1307_), .Y(new_n11067_));
  NOR2  g10682(.A(new_n11067_), .B(new_n1311_), .Y(new_n11068_));
  NOR2  g10683(.A(new_n11068_), .B(new_n1315_), .Y(new_n11069_));
  NOR2  g10684(.A(new_n11069_), .B(new_n1319_), .Y(new_n11070_));
  NOR2  g10685(.A(new_n11070_), .B(new_n1323_), .Y(new_n11071_));
  NOR2  g10686(.A(new_n11071_), .B(new_n1327_), .Y(new_n11072_));
  NOR2  g10687(.A(new_n11072_), .B(new_n1331_), .Y(new_n11073_));
  NOR2  g10688(.A(new_n11073_), .B(new_n1335_), .Y(new_n11074_));
  NOR2  g10689(.A(new_n11074_), .B(new_n1339_), .Y(new_n11075_));
  NOR2  g10690(.A(new_n11075_), .B(new_n1343_), .Y(new_n11076_));
  NOR2  g10691(.A(new_n11076_), .B(new_n1347_), .Y(new_n11077_));
  NOR2  g10692(.A(new_n11077_), .B(new_n1351_), .Y(new_n11078_));
  NOR2  g10693(.A(new_n11078_), .B(new_n1355_), .Y(new_n11079_));
  NOR2  g10694(.A(new_n11079_), .B(new_n1359_), .Y(new_n11080_));
  NOR2  g10695(.A(new_n11080_), .B(new_n1363_), .Y(new_n11081_));
  NOR2  g10696(.A(new_n11081_), .B(new_n1367_), .Y(new_n11082_));
  NOR2  g10697(.A(new_n11082_), .B(new_n1371_), .Y(new_n11083_));
  NOR2  g10698(.A(new_n11083_), .B(new_n1375_), .Y(new_n11084_));
  NOR2  g10699(.A(new_n11084_), .B(new_n1379_), .Y(new_n11085_));
  NOR2  g10700(.A(new_n11085_), .B(new_n1383_), .Y(new_n11086_));
  NOR2  g10701(.A(new_n11086_), .B(new_n1387_), .Y(new_n11087_));
  NOR2  g10702(.A(new_n11087_), .B(new_n1391_), .Y(new_n11088_));
  NOR2  g10703(.A(new_n11088_), .B(new_n1395_), .Y(new_n11089_));
  NOR2  g10704(.A(new_n11089_), .B(new_n1399_), .Y(new_n11090_));
  NOR2  g10705(.A(new_n11090_), .B(new_n1403_), .Y(new_n11091_));
  NOR2  g10706(.A(new_n11091_), .B(new_n1407_), .Y(new_n11092_));
  NOR2  g10707(.A(new_n11092_), .B(new_n1411_), .Y(new_n11093_));
  NOR2  g10708(.A(new_n11093_), .B(new_n1415_), .Y(new_n11094_));
  NOR2  g10709(.A(new_n11094_), .B(new_n1419_), .Y(new_n11095_));
  NOR2  g10710(.A(new_n11095_), .B(new_n1423_), .Y(new_n11096_));
  NOR2  g10711(.A(new_n11096_), .B(new_n1427_), .Y(new_n11097_));
  NOR2  g10712(.A(new_n11097_), .B(new_n1431_), .Y(new_n11098_));
  NOR2  g10713(.A(new_n11098_), .B(new_n1435_), .Y(new_n11099_));
  NOR2  g10714(.A(new_n11099_), .B(new_n1439_), .Y(new_n11100_));
  NOR2  g10715(.A(new_n11100_), .B(new_n1443_), .Y(new_n11101_));
  NOR2  g10716(.A(new_n11101_), .B(new_n1447_), .Y(new_n11102_));
  NOR2  g10717(.A(new_n11102_), .B(new_n1451_), .Y(new_n11103_));
  NOR2  g10718(.A(new_n11103_), .B(new_n1455_), .Y(new_n11104_));
  NOR2  g10719(.A(new_n11104_), .B(new_n1459_), .Y(new_n11105_));
  NOR2  g10720(.A(new_n11105_), .B(new_n1463_), .Y(new_n11106_));
  NOR2  g10721(.A(new_n11106_), .B(new_n1467_), .Y(new_n11107_));
  NOR2  g10722(.A(new_n11107_), .B(new_n1471_), .Y(new_n11108_));
  NOR2  g10723(.A(new_n11108_), .B(new_n1475_), .Y(new_n11109_));
  NOR2  g10724(.A(new_n11109_), .B(new_n1479_), .Y(new_n11110_));
  NAND2 g10725(.A(new_n1481_), .B(\req[112] ), .Y(new_n11111_));
  NOR2  g10726(.A(new_n11111_), .B(new_n11110_), .Y(\grant[112] ));
  INV   g10727(.A(new_n1490_), .Y(new_n11113_));
  NOR2  g10728(.A(new_n11113_), .B(new_n765_), .Y(new_n11114_));
  NOR2  g10729(.A(new_n11114_), .B(new_n1495_), .Y(new_n11115_));
  NOR2  g10730(.A(new_n11115_), .B(new_n1499_), .Y(new_n11116_));
  NOR2  g10731(.A(new_n11116_), .B(new_n1503_), .Y(new_n11117_));
  NOR2  g10732(.A(new_n11117_), .B(new_n1507_), .Y(new_n11118_));
  NOR2  g10733(.A(new_n11118_), .B(new_n1511_), .Y(new_n11119_));
  NOR2  g10734(.A(new_n11119_), .B(new_n1515_), .Y(new_n11120_));
  NOR2  g10735(.A(new_n11120_), .B(new_n1519_), .Y(new_n11121_));
  NOR2  g10736(.A(new_n11121_), .B(new_n1523_), .Y(new_n11122_));
  NOR2  g10737(.A(new_n11122_), .B(new_n1527_), .Y(new_n11123_));
  NOR2  g10738(.A(new_n11123_), .B(new_n1797_), .Y(new_n11124_));
  NOR2  g10739(.A(new_n11124_), .B(new_n396_), .Y(new_n11125_));
  NOR2  g10740(.A(new_n11125_), .B(new_n400_), .Y(new_n11126_));
  NOR2  g10741(.A(new_n11126_), .B(new_n406_), .Y(new_n11127_));
  NOR2  g10742(.A(new_n11127_), .B(new_n410_), .Y(new_n11128_));
  NOR2  g10743(.A(new_n11128_), .B(new_n416_), .Y(new_n11129_));
  NOR2  g10744(.A(new_n11129_), .B(new_n420_), .Y(new_n11130_));
  NOR2  g10745(.A(new_n11130_), .B(new_n426_), .Y(new_n11131_));
  NOR2  g10746(.A(new_n11131_), .B(new_n430_), .Y(new_n11132_));
  NOR2  g10747(.A(new_n11132_), .B(new_n436_), .Y(new_n11133_));
  NOR2  g10748(.A(new_n11133_), .B(new_n440_), .Y(new_n11134_));
  NOR2  g10749(.A(new_n11134_), .B(new_n446_), .Y(new_n11135_));
  NOR2  g10750(.A(new_n11135_), .B(new_n450_), .Y(new_n11136_));
  NOR2  g10751(.A(new_n11136_), .B(new_n456_), .Y(new_n11137_));
  NOR2  g10752(.A(new_n11137_), .B(new_n460_), .Y(new_n11138_));
  NOR2  g10753(.A(new_n11138_), .B(new_n466_), .Y(new_n11139_));
  NOR2  g10754(.A(new_n11139_), .B(new_n470_), .Y(new_n11140_));
  NOR2  g10755(.A(new_n11140_), .B(new_n476_), .Y(new_n11141_));
  NOR2  g10756(.A(new_n11141_), .B(new_n480_), .Y(new_n11142_));
  NOR2  g10757(.A(new_n11142_), .B(new_n486_), .Y(new_n11143_));
  NOR2  g10758(.A(new_n11143_), .B(new_n490_), .Y(new_n11144_));
  NOR2  g10759(.A(new_n11144_), .B(new_n496_), .Y(new_n11145_));
  NOR2  g10760(.A(new_n11145_), .B(new_n500_), .Y(new_n11146_));
  NOR2  g10761(.A(new_n11146_), .B(new_n506_), .Y(new_n11147_));
  NOR2  g10762(.A(new_n11147_), .B(new_n510_), .Y(new_n11148_));
  NOR2  g10763(.A(new_n11148_), .B(new_n516_), .Y(new_n11149_));
  NOR2  g10764(.A(new_n11149_), .B(new_n520_), .Y(new_n11150_));
  NOR2  g10765(.A(new_n11150_), .B(new_n526_), .Y(new_n11151_));
  NOR2  g10766(.A(new_n11151_), .B(new_n530_), .Y(new_n11152_));
  NOR2  g10767(.A(new_n11152_), .B(new_n536_), .Y(new_n11153_));
  NOR2  g10768(.A(new_n11153_), .B(new_n540_), .Y(new_n11154_));
  NOR2  g10769(.A(new_n11154_), .B(new_n546_), .Y(new_n11155_));
  NOR2  g10770(.A(new_n11155_), .B(new_n550_), .Y(new_n11156_));
  NOR2  g10771(.A(new_n11156_), .B(new_n556_), .Y(new_n11157_));
  NOR2  g10772(.A(new_n11157_), .B(new_n560_), .Y(new_n11158_));
  NOR2  g10773(.A(new_n11158_), .B(new_n566_), .Y(new_n11159_));
  NOR2  g10774(.A(new_n11159_), .B(new_n570_), .Y(new_n11160_));
  NOR2  g10775(.A(new_n11160_), .B(new_n576_), .Y(new_n11161_));
  NOR2  g10776(.A(new_n11161_), .B(new_n580_), .Y(new_n11162_));
  NOR2  g10777(.A(new_n11162_), .B(new_n586_), .Y(new_n11163_));
  NOR2  g10778(.A(new_n11163_), .B(new_n590_), .Y(new_n11164_));
  NOR2  g10779(.A(new_n11164_), .B(new_n596_), .Y(new_n11165_));
  NOR2  g10780(.A(new_n11165_), .B(new_n600_), .Y(new_n11166_));
  NOR2  g10781(.A(new_n11166_), .B(new_n606_), .Y(new_n11167_));
  NOR2  g10782(.A(new_n11167_), .B(new_n610_), .Y(new_n11168_));
  NOR2  g10783(.A(new_n11168_), .B(new_n616_), .Y(new_n11169_));
  NOR2  g10784(.A(new_n11169_), .B(new_n620_), .Y(new_n11170_));
  NOR2  g10785(.A(new_n11170_), .B(new_n626_), .Y(new_n11171_));
  NOR2  g10786(.A(new_n11171_), .B(new_n630_), .Y(new_n11172_));
  NOR2  g10787(.A(new_n11172_), .B(new_n636_), .Y(new_n11173_));
  NOR2  g10788(.A(new_n11173_), .B(new_n640_), .Y(new_n11174_));
  NOR2  g10789(.A(new_n11174_), .B(new_n646_), .Y(new_n11175_));
  NOR2  g10790(.A(new_n11175_), .B(new_n650_), .Y(new_n11176_));
  NOR2  g10791(.A(new_n11176_), .B(new_n656_), .Y(new_n11177_));
  NOR2  g10792(.A(new_n11177_), .B(new_n660_), .Y(new_n11178_));
  NOR2  g10793(.A(new_n11178_), .B(new_n666_), .Y(new_n11179_));
  NOR2  g10794(.A(new_n11179_), .B(new_n670_), .Y(new_n11180_));
  NOR2  g10795(.A(new_n11180_), .B(new_n676_), .Y(new_n11181_));
  NOR2  g10796(.A(new_n11181_), .B(new_n680_), .Y(new_n11182_));
  NOR2  g10797(.A(new_n11182_), .B(new_n686_), .Y(new_n11183_));
  NOR2  g10798(.A(new_n11183_), .B(new_n690_), .Y(new_n11184_));
  NOR2  g10799(.A(new_n11184_), .B(new_n696_), .Y(new_n11185_));
  NOR2  g10800(.A(new_n11185_), .B(new_n700_), .Y(new_n11186_));
  NOR2  g10801(.A(new_n11186_), .B(new_n706_), .Y(new_n11187_));
  NOR2  g10802(.A(new_n11187_), .B(new_n710_), .Y(new_n11188_));
  NOR2  g10803(.A(new_n11188_), .B(new_n716_), .Y(new_n11189_));
  NOR2  g10804(.A(new_n11189_), .B(new_n720_), .Y(new_n11190_));
  NOR2  g10805(.A(new_n11190_), .B(new_n726_), .Y(new_n11191_));
  NOR2  g10806(.A(new_n11191_), .B(new_n730_), .Y(new_n11192_));
  NOR2  g10807(.A(new_n11192_), .B(new_n736_), .Y(new_n11193_));
  NOR2  g10808(.A(new_n11193_), .B(new_n740_), .Y(new_n11194_));
  NOR2  g10809(.A(new_n11194_), .B(new_n746_), .Y(new_n11195_));
  NOR2  g10810(.A(new_n11195_), .B(new_n750_), .Y(new_n11196_));
  NOR2  g10811(.A(new_n11196_), .B(new_n756_), .Y(new_n11197_));
  NAND2 g10812(.A(new_n758_), .B(\req[113] ), .Y(new_n11198_));
  NOR2  g10813(.A(new_n11198_), .B(new_n11197_), .Y(\grant[113] ));
  INV   g10814(.A(new_n769_), .Y(new_n11200_));
  NOR2  g10815(.A(new_n1152_), .B(new_n11200_), .Y(new_n11201_));
  NOR2  g10816(.A(new_n11201_), .B(new_n776_), .Y(new_n11202_));
  NOR2  g10817(.A(new_n11202_), .B(new_n780_), .Y(new_n11203_));
  NOR2  g10818(.A(new_n11203_), .B(new_n786_), .Y(new_n11204_));
  NOR2  g10819(.A(new_n11204_), .B(new_n790_), .Y(new_n11205_));
  NOR2  g10820(.A(new_n11205_), .B(new_n796_), .Y(new_n11206_));
  NOR2  g10821(.A(new_n11206_), .B(new_n800_), .Y(new_n11207_));
  NOR2  g10822(.A(new_n11207_), .B(new_n806_), .Y(new_n11208_));
  NOR2  g10823(.A(new_n11208_), .B(new_n1616_), .Y(new_n11209_));
  NOR2  g10824(.A(new_n11209_), .B(new_n1618_), .Y(new_n11210_));
  NOR2  g10825(.A(new_n11210_), .B(new_n1885_), .Y(new_n11211_));
  NOR2  g10826(.A(new_n11211_), .B(new_n820_), .Y(new_n11212_));
  NOR2  g10827(.A(new_n11212_), .B(new_n824_), .Y(new_n11213_));
  NOR2  g10828(.A(new_n11213_), .B(new_n829_), .Y(new_n11214_));
  NOR2  g10829(.A(new_n11214_), .B(new_n833_), .Y(new_n11215_));
  NOR2  g10830(.A(new_n11215_), .B(new_n838_), .Y(new_n11216_));
  NOR2  g10831(.A(new_n11216_), .B(new_n842_), .Y(new_n11217_));
  NOR2  g10832(.A(new_n11217_), .B(new_n847_), .Y(new_n11218_));
  NOR2  g10833(.A(new_n11218_), .B(new_n851_), .Y(new_n11219_));
  NOR2  g10834(.A(new_n11219_), .B(new_n856_), .Y(new_n11220_));
  NOR2  g10835(.A(new_n11220_), .B(new_n860_), .Y(new_n11221_));
  NOR2  g10836(.A(new_n11221_), .B(new_n865_), .Y(new_n11222_));
  NOR2  g10837(.A(new_n11222_), .B(new_n869_), .Y(new_n11223_));
  NOR2  g10838(.A(new_n11223_), .B(new_n874_), .Y(new_n11224_));
  NOR2  g10839(.A(new_n11224_), .B(new_n878_), .Y(new_n11225_));
  NOR2  g10840(.A(new_n11225_), .B(new_n883_), .Y(new_n11226_));
  NOR2  g10841(.A(new_n11226_), .B(new_n887_), .Y(new_n11227_));
  NOR2  g10842(.A(new_n11227_), .B(new_n892_), .Y(new_n11228_));
  NOR2  g10843(.A(new_n11228_), .B(new_n896_), .Y(new_n11229_));
  NOR2  g10844(.A(new_n11229_), .B(new_n901_), .Y(new_n11230_));
  NOR2  g10845(.A(new_n11230_), .B(new_n905_), .Y(new_n11231_));
  NOR2  g10846(.A(new_n11231_), .B(new_n910_), .Y(new_n11232_));
  NOR2  g10847(.A(new_n11232_), .B(new_n914_), .Y(new_n11233_));
  NOR2  g10848(.A(new_n11233_), .B(new_n919_), .Y(new_n11234_));
  NOR2  g10849(.A(new_n11234_), .B(new_n923_), .Y(new_n11235_));
  NOR2  g10850(.A(new_n11235_), .B(new_n928_), .Y(new_n11236_));
  NOR2  g10851(.A(new_n11236_), .B(new_n932_), .Y(new_n11237_));
  NOR2  g10852(.A(new_n11237_), .B(new_n937_), .Y(new_n11238_));
  NOR2  g10853(.A(new_n11238_), .B(new_n941_), .Y(new_n11239_));
  NOR2  g10854(.A(new_n11239_), .B(new_n946_), .Y(new_n11240_));
  NOR2  g10855(.A(new_n11240_), .B(new_n950_), .Y(new_n11241_));
  NOR2  g10856(.A(new_n11241_), .B(new_n955_), .Y(new_n11242_));
  NOR2  g10857(.A(new_n11242_), .B(new_n959_), .Y(new_n11243_));
  NOR2  g10858(.A(new_n11243_), .B(new_n964_), .Y(new_n11244_));
  NOR2  g10859(.A(new_n11244_), .B(new_n968_), .Y(new_n11245_));
  NOR2  g10860(.A(new_n11245_), .B(new_n973_), .Y(new_n11246_));
  NOR2  g10861(.A(new_n11246_), .B(new_n977_), .Y(new_n11247_));
  NOR2  g10862(.A(new_n11247_), .B(new_n982_), .Y(new_n11248_));
  NOR2  g10863(.A(new_n11248_), .B(new_n986_), .Y(new_n11249_));
  NOR2  g10864(.A(new_n11249_), .B(new_n991_), .Y(new_n11250_));
  NOR2  g10865(.A(new_n11250_), .B(new_n995_), .Y(new_n11251_));
  NOR2  g10866(.A(new_n11251_), .B(new_n1000_), .Y(new_n11252_));
  NOR2  g10867(.A(new_n11252_), .B(new_n1004_), .Y(new_n11253_));
  NOR2  g10868(.A(new_n11253_), .B(new_n1009_), .Y(new_n11254_));
  NOR2  g10869(.A(new_n11254_), .B(new_n1013_), .Y(new_n11255_));
  NOR2  g10870(.A(new_n11255_), .B(new_n1018_), .Y(new_n11256_));
  NOR2  g10871(.A(new_n11256_), .B(new_n1022_), .Y(new_n11257_));
  NOR2  g10872(.A(new_n11257_), .B(new_n1027_), .Y(new_n11258_));
  NOR2  g10873(.A(new_n11258_), .B(new_n1031_), .Y(new_n11259_));
  NOR2  g10874(.A(new_n11259_), .B(new_n1036_), .Y(new_n11260_));
  NOR2  g10875(.A(new_n11260_), .B(new_n1040_), .Y(new_n11261_));
  NOR2  g10876(.A(new_n11261_), .B(new_n1045_), .Y(new_n11262_));
  NOR2  g10877(.A(new_n11262_), .B(new_n1049_), .Y(new_n11263_));
  NOR2  g10878(.A(new_n11263_), .B(new_n1054_), .Y(new_n11264_));
  NOR2  g10879(.A(new_n11264_), .B(new_n1058_), .Y(new_n11265_));
  NOR2  g10880(.A(new_n11265_), .B(new_n1063_), .Y(new_n11266_));
  NOR2  g10881(.A(new_n11266_), .B(new_n1067_), .Y(new_n11267_));
  NOR2  g10882(.A(new_n11267_), .B(new_n1072_), .Y(new_n11268_));
  NOR2  g10883(.A(new_n11268_), .B(new_n1076_), .Y(new_n11269_));
  NOR2  g10884(.A(new_n11269_), .B(new_n1081_), .Y(new_n11270_));
  NOR2  g10885(.A(new_n11270_), .B(new_n1085_), .Y(new_n11271_));
  NOR2  g10886(.A(new_n11271_), .B(new_n1090_), .Y(new_n11272_));
  NOR2  g10887(.A(new_n11272_), .B(new_n1094_), .Y(new_n11273_));
  NOR2  g10888(.A(new_n11273_), .B(new_n1099_), .Y(new_n11274_));
  NOR2  g10889(.A(new_n11274_), .B(new_n1103_), .Y(new_n11275_));
  NOR2  g10890(.A(new_n11275_), .B(new_n1108_), .Y(new_n11276_));
  NOR2  g10891(.A(new_n11276_), .B(new_n1112_), .Y(new_n11277_));
  NOR2  g10892(.A(new_n11277_), .B(new_n1117_), .Y(new_n11278_));
  NOR2  g10893(.A(new_n11278_), .B(new_n1121_), .Y(new_n11279_));
  NOR2  g10894(.A(new_n11279_), .B(new_n1126_), .Y(new_n11280_));
  NOR2  g10895(.A(new_n11280_), .B(new_n1130_), .Y(new_n11281_));
  NOR2  g10896(.A(new_n11281_), .B(new_n1135_), .Y(new_n11282_));
  NOR2  g10897(.A(new_n11282_), .B(new_n1139_), .Y(new_n11283_));
  NOR2  g10898(.A(new_n11283_), .B(new_n1144_), .Y(new_n11284_));
  NAND2 g10899(.A(new_n1146_), .B(\req[114] ), .Y(new_n11285_));
  NOR2  g10900(.A(new_n11285_), .B(new_n11284_), .Y(\grant[114] ));
  INV   g10901(.A(new_n1156_), .Y(new_n11287_));
  NOR2  g10902(.A(new_n1494_), .B(new_n11287_), .Y(new_n11288_));
  NOR2  g10903(.A(new_n11288_), .B(new_n1162_), .Y(new_n11289_));
  NOR2  g10904(.A(new_n11289_), .B(new_n1166_), .Y(new_n11290_));
  NOR2  g10905(.A(new_n11290_), .B(new_n1171_), .Y(new_n11291_));
  NOR2  g10906(.A(new_n11291_), .B(new_n1175_), .Y(new_n11292_));
  NOR2  g10907(.A(new_n11292_), .B(new_n1180_), .Y(new_n11293_));
  NOR2  g10908(.A(new_n11293_), .B(new_n1184_), .Y(new_n11294_));
  NOR2  g10909(.A(new_n11294_), .B(new_n1189_), .Y(new_n11295_));
  NOR2  g10910(.A(new_n11295_), .B(new_n1707_), .Y(new_n11296_));
  NOR2  g10911(.A(new_n11296_), .B(new_n1709_), .Y(new_n11297_));
  NOR2  g10912(.A(new_n11297_), .B(new_n1973_), .Y(new_n11298_));
  NOR2  g10913(.A(new_n11298_), .B(new_n1199_), .Y(new_n11299_));
  NOR2  g10914(.A(new_n11299_), .B(new_n1203_), .Y(new_n11300_));
  NOR2  g10915(.A(new_n11300_), .B(new_n1207_), .Y(new_n11301_));
  NOR2  g10916(.A(new_n11301_), .B(new_n1211_), .Y(new_n11302_));
  NOR2  g10917(.A(new_n11302_), .B(new_n1215_), .Y(new_n11303_));
  NOR2  g10918(.A(new_n11303_), .B(new_n1219_), .Y(new_n11304_));
  NOR2  g10919(.A(new_n11304_), .B(new_n1223_), .Y(new_n11305_));
  NOR2  g10920(.A(new_n11305_), .B(new_n1227_), .Y(new_n11306_));
  NOR2  g10921(.A(new_n11306_), .B(new_n1231_), .Y(new_n11307_));
  NOR2  g10922(.A(new_n11307_), .B(new_n1235_), .Y(new_n11308_));
  NOR2  g10923(.A(new_n11308_), .B(new_n1239_), .Y(new_n11309_));
  NOR2  g10924(.A(new_n11309_), .B(new_n1243_), .Y(new_n11310_));
  NOR2  g10925(.A(new_n11310_), .B(new_n1247_), .Y(new_n11311_));
  NOR2  g10926(.A(new_n11311_), .B(new_n1251_), .Y(new_n11312_));
  NOR2  g10927(.A(new_n11312_), .B(new_n1255_), .Y(new_n11313_));
  NOR2  g10928(.A(new_n11313_), .B(new_n1259_), .Y(new_n11314_));
  NOR2  g10929(.A(new_n11314_), .B(new_n1263_), .Y(new_n11315_));
  NOR2  g10930(.A(new_n11315_), .B(new_n1267_), .Y(new_n11316_));
  NOR2  g10931(.A(new_n11316_), .B(new_n1271_), .Y(new_n11317_));
  NOR2  g10932(.A(new_n11317_), .B(new_n1275_), .Y(new_n11318_));
  NOR2  g10933(.A(new_n11318_), .B(new_n1279_), .Y(new_n11319_));
  NOR2  g10934(.A(new_n11319_), .B(new_n1283_), .Y(new_n11320_));
  NOR2  g10935(.A(new_n11320_), .B(new_n1287_), .Y(new_n11321_));
  NOR2  g10936(.A(new_n11321_), .B(new_n1291_), .Y(new_n11322_));
  NOR2  g10937(.A(new_n11322_), .B(new_n1295_), .Y(new_n11323_));
  NOR2  g10938(.A(new_n11323_), .B(new_n1299_), .Y(new_n11324_));
  NOR2  g10939(.A(new_n11324_), .B(new_n1303_), .Y(new_n11325_));
  NOR2  g10940(.A(new_n11325_), .B(new_n1307_), .Y(new_n11326_));
  NOR2  g10941(.A(new_n11326_), .B(new_n1311_), .Y(new_n11327_));
  NOR2  g10942(.A(new_n11327_), .B(new_n1315_), .Y(new_n11328_));
  NOR2  g10943(.A(new_n11328_), .B(new_n1319_), .Y(new_n11329_));
  NOR2  g10944(.A(new_n11329_), .B(new_n1323_), .Y(new_n11330_));
  NOR2  g10945(.A(new_n11330_), .B(new_n1327_), .Y(new_n11331_));
  NOR2  g10946(.A(new_n11331_), .B(new_n1331_), .Y(new_n11332_));
  NOR2  g10947(.A(new_n11332_), .B(new_n1335_), .Y(new_n11333_));
  NOR2  g10948(.A(new_n11333_), .B(new_n1339_), .Y(new_n11334_));
  NOR2  g10949(.A(new_n11334_), .B(new_n1343_), .Y(new_n11335_));
  NOR2  g10950(.A(new_n11335_), .B(new_n1347_), .Y(new_n11336_));
  NOR2  g10951(.A(new_n11336_), .B(new_n1351_), .Y(new_n11337_));
  NOR2  g10952(.A(new_n11337_), .B(new_n1355_), .Y(new_n11338_));
  NOR2  g10953(.A(new_n11338_), .B(new_n1359_), .Y(new_n11339_));
  NOR2  g10954(.A(new_n11339_), .B(new_n1363_), .Y(new_n11340_));
  NOR2  g10955(.A(new_n11340_), .B(new_n1367_), .Y(new_n11341_));
  NOR2  g10956(.A(new_n11341_), .B(new_n1371_), .Y(new_n11342_));
  NOR2  g10957(.A(new_n11342_), .B(new_n1375_), .Y(new_n11343_));
  NOR2  g10958(.A(new_n11343_), .B(new_n1379_), .Y(new_n11344_));
  NOR2  g10959(.A(new_n11344_), .B(new_n1383_), .Y(new_n11345_));
  NOR2  g10960(.A(new_n11345_), .B(new_n1387_), .Y(new_n11346_));
  NOR2  g10961(.A(new_n11346_), .B(new_n1391_), .Y(new_n11347_));
  NOR2  g10962(.A(new_n11347_), .B(new_n1395_), .Y(new_n11348_));
  NOR2  g10963(.A(new_n11348_), .B(new_n1399_), .Y(new_n11349_));
  NOR2  g10964(.A(new_n11349_), .B(new_n1403_), .Y(new_n11350_));
  NOR2  g10965(.A(new_n11350_), .B(new_n1407_), .Y(new_n11351_));
  NOR2  g10966(.A(new_n11351_), .B(new_n1411_), .Y(new_n11352_));
  NOR2  g10967(.A(new_n11352_), .B(new_n1415_), .Y(new_n11353_));
  NOR2  g10968(.A(new_n11353_), .B(new_n1419_), .Y(new_n11354_));
  NOR2  g10969(.A(new_n11354_), .B(new_n1423_), .Y(new_n11355_));
  NOR2  g10970(.A(new_n11355_), .B(new_n1427_), .Y(new_n11356_));
  NOR2  g10971(.A(new_n11356_), .B(new_n1431_), .Y(new_n11357_));
  NOR2  g10972(.A(new_n11357_), .B(new_n1435_), .Y(new_n11358_));
  NOR2  g10973(.A(new_n11358_), .B(new_n1439_), .Y(new_n11359_));
  NOR2  g10974(.A(new_n11359_), .B(new_n1443_), .Y(new_n11360_));
  NOR2  g10975(.A(new_n11360_), .B(new_n1447_), .Y(new_n11361_));
  NOR2  g10976(.A(new_n11361_), .B(new_n1451_), .Y(new_n11362_));
  NOR2  g10977(.A(new_n11362_), .B(new_n1455_), .Y(new_n11363_));
  NOR2  g10978(.A(new_n11363_), .B(new_n1459_), .Y(new_n11364_));
  NOR2  g10979(.A(new_n11364_), .B(new_n1463_), .Y(new_n11365_));
  NOR2  g10980(.A(new_n11365_), .B(new_n1467_), .Y(new_n11366_));
  NOR2  g10981(.A(new_n11366_), .B(new_n1471_), .Y(new_n11367_));
  NOR2  g10982(.A(new_n11367_), .B(new_n1475_), .Y(new_n11368_));
  NOR2  g10983(.A(new_n11368_), .B(new_n1479_), .Y(new_n11369_));
  NOR2  g10984(.A(new_n11369_), .B(new_n1483_), .Y(new_n11370_));
  NOR2  g10985(.A(new_n11370_), .B(new_n1487_), .Y(new_n11371_));
  NAND2 g10986(.A(new_n1489_), .B(\req[115] ), .Y(new_n11372_));
  NOR2  g10987(.A(new_n11372_), .B(new_n11371_), .Y(\grant[115] ));
  INV   g10988(.A(new_n1498_), .Y(new_n11374_));
  NOR2  g10989(.A(new_n11374_), .B(new_n775_), .Y(new_n11375_));
  NOR2  g10990(.A(new_n11375_), .B(new_n1503_), .Y(new_n11376_));
  NOR2  g10991(.A(new_n11376_), .B(new_n1507_), .Y(new_n11377_));
  NOR2  g10992(.A(new_n11377_), .B(new_n1511_), .Y(new_n11378_));
  NOR2  g10993(.A(new_n11378_), .B(new_n1515_), .Y(new_n11379_));
  NOR2  g10994(.A(new_n11379_), .B(new_n1519_), .Y(new_n11380_));
  NOR2  g10995(.A(new_n11380_), .B(new_n1523_), .Y(new_n11381_));
  NOR2  g10996(.A(new_n11381_), .B(new_n1527_), .Y(new_n11382_));
  NOR2  g10997(.A(new_n11382_), .B(new_n1797_), .Y(new_n11383_));
  NOR2  g10998(.A(new_n11383_), .B(new_n396_), .Y(new_n11384_));
  NOR2  g10999(.A(new_n11384_), .B(new_n400_), .Y(new_n11385_));
  NOR2  g11000(.A(new_n11385_), .B(new_n406_), .Y(new_n11386_));
  NOR2  g11001(.A(new_n11386_), .B(new_n410_), .Y(new_n11387_));
  NOR2  g11002(.A(new_n11387_), .B(new_n416_), .Y(new_n11388_));
  NOR2  g11003(.A(new_n11388_), .B(new_n420_), .Y(new_n11389_));
  NOR2  g11004(.A(new_n11389_), .B(new_n426_), .Y(new_n11390_));
  NOR2  g11005(.A(new_n11390_), .B(new_n430_), .Y(new_n11391_));
  NOR2  g11006(.A(new_n11391_), .B(new_n436_), .Y(new_n11392_));
  NOR2  g11007(.A(new_n11392_), .B(new_n440_), .Y(new_n11393_));
  NOR2  g11008(.A(new_n11393_), .B(new_n446_), .Y(new_n11394_));
  NOR2  g11009(.A(new_n11394_), .B(new_n450_), .Y(new_n11395_));
  NOR2  g11010(.A(new_n11395_), .B(new_n456_), .Y(new_n11396_));
  NOR2  g11011(.A(new_n11396_), .B(new_n460_), .Y(new_n11397_));
  NOR2  g11012(.A(new_n11397_), .B(new_n466_), .Y(new_n11398_));
  NOR2  g11013(.A(new_n11398_), .B(new_n470_), .Y(new_n11399_));
  NOR2  g11014(.A(new_n11399_), .B(new_n476_), .Y(new_n11400_));
  NOR2  g11015(.A(new_n11400_), .B(new_n480_), .Y(new_n11401_));
  NOR2  g11016(.A(new_n11401_), .B(new_n486_), .Y(new_n11402_));
  NOR2  g11017(.A(new_n11402_), .B(new_n490_), .Y(new_n11403_));
  NOR2  g11018(.A(new_n11403_), .B(new_n496_), .Y(new_n11404_));
  NOR2  g11019(.A(new_n11404_), .B(new_n500_), .Y(new_n11405_));
  NOR2  g11020(.A(new_n11405_), .B(new_n506_), .Y(new_n11406_));
  NOR2  g11021(.A(new_n11406_), .B(new_n510_), .Y(new_n11407_));
  NOR2  g11022(.A(new_n11407_), .B(new_n516_), .Y(new_n11408_));
  NOR2  g11023(.A(new_n11408_), .B(new_n520_), .Y(new_n11409_));
  NOR2  g11024(.A(new_n11409_), .B(new_n526_), .Y(new_n11410_));
  NOR2  g11025(.A(new_n11410_), .B(new_n530_), .Y(new_n11411_));
  NOR2  g11026(.A(new_n11411_), .B(new_n536_), .Y(new_n11412_));
  NOR2  g11027(.A(new_n11412_), .B(new_n540_), .Y(new_n11413_));
  NOR2  g11028(.A(new_n11413_), .B(new_n546_), .Y(new_n11414_));
  NOR2  g11029(.A(new_n11414_), .B(new_n550_), .Y(new_n11415_));
  NOR2  g11030(.A(new_n11415_), .B(new_n556_), .Y(new_n11416_));
  NOR2  g11031(.A(new_n11416_), .B(new_n560_), .Y(new_n11417_));
  NOR2  g11032(.A(new_n11417_), .B(new_n566_), .Y(new_n11418_));
  NOR2  g11033(.A(new_n11418_), .B(new_n570_), .Y(new_n11419_));
  NOR2  g11034(.A(new_n11419_), .B(new_n576_), .Y(new_n11420_));
  NOR2  g11035(.A(new_n11420_), .B(new_n580_), .Y(new_n11421_));
  NOR2  g11036(.A(new_n11421_), .B(new_n586_), .Y(new_n11422_));
  NOR2  g11037(.A(new_n11422_), .B(new_n590_), .Y(new_n11423_));
  NOR2  g11038(.A(new_n11423_), .B(new_n596_), .Y(new_n11424_));
  NOR2  g11039(.A(new_n11424_), .B(new_n600_), .Y(new_n11425_));
  NOR2  g11040(.A(new_n11425_), .B(new_n606_), .Y(new_n11426_));
  NOR2  g11041(.A(new_n11426_), .B(new_n610_), .Y(new_n11427_));
  NOR2  g11042(.A(new_n11427_), .B(new_n616_), .Y(new_n11428_));
  NOR2  g11043(.A(new_n11428_), .B(new_n620_), .Y(new_n11429_));
  NOR2  g11044(.A(new_n11429_), .B(new_n626_), .Y(new_n11430_));
  NOR2  g11045(.A(new_n11430_), .B(new_n630_), .Y(new_n11431_));
  NOR2  g11046(.A(new_n11431_), .B(new_n636_), .Y(new_n11432_));
  NOR2  g11047(.A(new_n11432_), .B(new_n640_), .Y(new_n11433_));
  NOR2  g11048(.A(new_n11433_), .B(new_n646_), .Y(new_n11434_));
  NOR2  g11049(.A(new_n11434_), .B(new_n650_), .Y(new_n11435_));
  NOR2  g11050(.A(new_n11435_), .B(new_n656_), .Y(new_n11436_));
  NOR2  g11051(.A(new_n11436_), .B(new_n660_), .Y(new_n11437_));
  NOR2  g11052(.A(new_n11437_), .B(new_n666_), .Y(new_n11438_));
  NOR2  g11053(.A(new_n11438_), .B(new_n670_), .Y(new_n11439_));
  NOR2  g11054(.A(new_n11439_), .B(new_n676_), .Y(new_n11440_));
  NOR2  g11055(.A(new_n11440_), .B(new_n680_), .Y(new_n11441_));
  NOR2  g11056(.A(new_n11441_), .B(new_n686_), .Y(new_n11442_));
  NOR2  g11057(.A(new_n11442_), .B(new_n690_), .Y(new_n11443_));
  NOR2  g11058(.A(new_n11443_), .B(new_n696_), .Y(new_n11444_));
  NOR2  g11059(.A(new_n11444_), .B(new_n700_), .Y(new_n11445_));
  NOR2  g11060(.A(new_n11445_), .B(new_n706_), .Y(new_n11446_));
  NOR2  g11061(.A(new_n11446_), .B(new_n710_), .Y(new_n11447_));
  NOR2  g11062(.A(new_n11447_), .B(new_n716_), .Y(new_n11448_));
  NOR2  g11063(.A(new_n11448_), .B(new_n720_), .Y(new_n11449_));
  NOR2  g11064(.A(new_n11449_), .B(new_n726_), .Y(new_n11450_));
  NOR2  g11065(.A(new_n11450_), .B(new_n730_), .Y(new_n11451_));
  NOR2  g11066(.A(new_n11451_), .B(new_n736_), .Y(new_n11452_));
  NOR2  g11067(.A(new_n11452_), .B(new_n740_), .Y(new_n11453_));
  NOR2  g11068(.A(new_n11453_), .B(new_n746_), .Y(new_n11454_));
  NOR2  g11069(.A(new_n11454_), .B(new_n750_), .Y(new_n11455_));
  NOR2  g11070(.A(new_n11455_), .B(new_n756_), .Y(new_n11456_));
  NOR2  g11071(.A(new_n11456_), .B(new_n760_), .Y(new_n11457_));
  NOR2  g11072(.A(new_n11457_), .B(new_n766_), .Y(new_n11458_));
  NAND2 g11073(.A(new_n768_), .B(\req[116] ), .Y(new_n11459_));
  NOR2  g11074(.A(new_n11459_), .B(new_n11458_), .Y(\grant[116] ));
  INV   g11075(.A(new_n779_), .Y(new_n11461_));
  NOR2  g11076(.A(new_n1161_), .B(new_n11461_), .Y(new_n11462_));
  NOR2  g11077(.A(new_n11462_), .B(new_n786_), .Y(new_n11463_));
  NOR2  g11078(.A(new_n11463_), .B(new_n790_), .Y(new_n11464_));
  NOR2  g11079(.A(new_n11464_), .B(new_n796_), .Y(new_n11465_));
  NOR2  g11080(.A(new_n11465_), .B(new_n800_), .Y(new_n11466_));
  NOR2  g11081(.A(new_n11466_), .B(new_n806_), .Y(new_n11467_));
  NOR2  g11082(.A(new_n11467_), .B(new_n1616_), .Y(new_n11468_));
  NOR2  g11083(.A(new_n11468_), .B(new_n1618_), .Y(new_n11469_));
  NOR2  g11084(.A(new_n11469_), .B(new_n1885_), .Y(new_n11470_));
  NOR2  g11085(.A(new_n11470_), .B(new_n820_), .Y(new_n11471_));
  NOR2  g11086(.A(new_n11471_), .B(new_n824_), .Y(new_n11472_));
  NOR2  g11087(.A(new_n11472_), .B(new_n829_), .Y(new_n11473_));
  NOR2  g11088(.A(new_n11473_), .B(new_n833_), .Y(new_n11474_));
  NOR2  g11089(.A(new_n11474_), .B(new_n838_), .Y(new_n11475_));
  NOR2  g11090(.A(new_n11475_), .B(new_n842_), .Y(new_n11476_));
  NOR2  g11091(.A(new_n11476_), .B(new_n847_), .Y(new_n11477_));
  NOR2  g11092(.A(new_n11477_), .B(new_n851_), .Y(new_n11478_));
  NOR2  g11093(.A(new_n11478_), .B(new_n856_), .Y(new_n11479_));
  NOR2  g11094(.A(new_n11479_), .B(new_n860_), .Y(new_n11480_));
  NOR2  g11095(.A(new_n11480_), .B(new_n865_), .Y(new_n11481_));
  NOR2  g11096(.A(new_n11481_), .B(new_n869_), .Y(new_n11482_));
  NOR2  g11097(.A(new_n11482_), .B(new_n874_), .Y(new_n11483_));
  NOR2  g11098(.A(new_n11483_), .B(new_n878_), .Y(new_n11484_));
  NOR2  g11099(.A(new_n11484_), .B(new_n883_), .Y(new_n11485_));
  NOR2  g11100(.A(new_n11485_), .B(new_n887_), .Y(new_n11486_));
  NOR2  g11101(.A(new_n11486_), .B(new_n892_), .Y(new_n11487_));
  NOR2  g11102(.A(new_n11487_), .B(new_n896_), .Y(new_n11488_));
  NOR2  g11103(.A(new_n11488_), .B(new_n901_), .Y(new_n11489_));
  NOR2  g11104(.A(new_n11489_), .B(new_n905_), .Y(new_n11490_));
  NOR2  g11105(.A(new_n11490_), .B(new_n910_), .Y(new_n11491_));
  NOR2  g11106(.A(new_n11491_), .B(new_n914_), .Y(new_n11492_));
  NOR2  g11107(.A(new_n11492_), .B(new_n919_), .Y(new_n11493_));
  NOR2  g11108(.A(new_n11493_), .B(new_n923_), .Y(new_n11494_));
  NOR2  g11109(.A(new_n11494_), .B(new_n928_), .Y(new_n11495_));
  NOR2  g11110(.A(new_n11495_), .B(new_n932_), .Y(new_n11496_));
  NOR2  g11111(.A(new_n11496_), .B(new_n937_), .Y(new_n11497_));
  NOR2  g11112(.A(new_n11497_), .B(new_n941_), .Y(new_n11498_));
  NOR2  g11113(.A(new_n11498_), .B(new_n946_), .Y(new_n11499_));
  NOR2  g11114(.A(new_n11499_), .B(new_n950_), .Y(new_n11500_));
  NOR2  g11115(.A(new_n11500_), .B(new_n955_), .Y(new_n11501_));
  NOR2  g11116(.A(new_n11501_), .B(new_n959_), .Y(new_n11502_));
  NOR2  g11117(.A(new_n11502_), .B(new_n964_), .Y(new_n11503_));
  NOR2  g11118(.A(new_n11503_), .B(new_n968_), .Y(new_n11504_));
  NOR2  g11119(.A(new_n11504_), .B(new_n973_), .Y(new_n11505_));
  NOR2  g11120(.A(new_n11505_), .B(new_n977_), .Y(new_n11506_));
  NOR2  g11121(.A(new_n11506_), .B(new_n982_), .Y(new_n11507_));
  NOR2  g11122(.A(new_n11507_), .B(new_n986_), .Y(new_n11508_));
  NOR2  g11123(.A(new_n11508_), .B(new_n991_), .Y(new_n11509_));
  NOR2  g11124(.A(new_n11509_), .B(new_n995_), .Y(new_n11510_));
  NOR2  g11125(.A(new_n11510_), .B(new_n1000_), .Y(new_n11511_));
  NOR2  g11126(.A(new_n11511_), .B(new_n1004_), .Y(new_n11512_));
  NOR2  g11127(.A(new_n11512_), .B(new_n1009_), .Y(new_n11513_));
  NOR2  g11128(.A(new_n11513_), .B(new_n1013_), .Y(new_n11514_));
  NOR2  g11129(.A(new_n11514_), .B(new_n1018_), .Y(new_n11515_));
  NOR2  g11130(.A(new_n11515_), .B(new_n1022_), .Y(new_n11516_));
  NOR2  g11131(.A(new_n11516_), .B(new_n1027_), .Y(new_n11517_));
  NOR2  g11132(.A(new_n11517_), .B(new_n1031_), .Y(new_n11518_));
  NOR2  g11133(.A(new_n11518_), .B(new_n1036_), .Y(new_n11519_));
  NOR2  g11134(.A(new_n11519_), .B(new_n1040_), .Y(new_n11520_));
  NOR2  g11135(.A(new_n11520_), .B(new_n1045_), .Y(new_n11521_));
  NOR2  g11136(.A(new_n11521_), .B(new_n1049_), .Y(new_n11522_));
  NOR2  g11137(.A(new_n11522_), .B(new_n1054_), .Y(new_n11523_));
  NOR2  g11138(.A(new_n11523_), .B(new_n1058_), .Y(new_n11524_));
  NOR2  g11139(.A(new_n11524_), .B(new_n1063_), .Y(new_n11525_));
  NOR2  g11140(.A(new_n11525_), .B(new_n1067_), .Y(new_n11526_));
  NOR2  g11141(.A(new_n11526_), .B(new_n1072_), .Y(new_n11527_));
  NOR2  g11142(.A(new_n11527_), .B(new_n1076_), .Y(new_n11528_));
  NOR2  g11143(.A(new_n11528_), .B(new_n1081_), .Y(new_n11529_));
  NOR2  g11144(.A(new_n11529_), .B(new_n1085_), .Y(new_n11530_));
  NOR2  g11145(.A(new_n11530_), .B(new_n1090_), .Y(new_n11531_));
  NOR2  g11146(.A(new_n11531_), .B(new_n1094_), .Y(new_n11532_));
  NOR2  g11147(.A(new_n11532_), .B(new_n1099_), .Y(new_n11533_));
  NOR2  g11148(.A(new_n11533_), .B(new_n1103_), .Y(new_n11534_));
  NOR2  g11149(.A(new_n11534_), .B(new_n1108_), .Y(new_n11535_));
  NOR2  g11150(.A(new_n11535_), .B(new_n1112_), .Y(new_n11536_));
  NOR2  g11151(.A(new_n11536_), .B(new_n1117_), .Y(new_n11537_));
  NOR2  g11152(.A(new_n11537_), .B(new_n1121_), .Y(new_n11538_));
  NOR2  g11153(.A(new_n11538_), .B(new_n1126_), .Y(new_n11539_));
  NOR2  g11154(.A(new_n11539_), .B(new_n1130_), .Y(new_n11540_));
  NOR2  g11155(.A(new_n11540_), .B(new_n1135_), .Y(new_n11541_));
  NOR2  g11156(.A(new_n11541_), .B(new_n1139_), .Y(new_n11542_));
  NOR2  g11157(.A(new_n11542_), .B(new_n1144_), .Y(new_n11543_));
  NOR2  g11158(.A(new_n11543_), .B(new_n1148_), .Y(new_n11544_));
  NOR2  g11159(.A(new_n11544_), .B(new_n1153_), .Y(new_n11545_));
  NAND2 g11160(.A(new_n1155_), .B(\req[117] ), .Y(new_n11546_));
  NOR2  g11161(.A(new_n11546_), .B(new_n11545_), .Y(\grant[117] ));
  INV   g11162(.A(new_n1165_), .Y(new_n11548_));
  NOR2  g11163(.A(new_n1502_), .B(new_n11548_), .Y(new_n11549_));
  NOR2  g11164(.A(new_n11549_), .B(new_n1171_), .Y(new_n11550_));
  NOR2  g11165(.A(new_n11550_), .B(new_n1175_), .Y(new_n11551_));
  NOR2  g11166(.A(new_n11551_), .B(new_n1180_), .Y(new_n11552_));
  NOR2  g11167(.A(new_n11552_), .B(new_n1184_), .Y(new_n11553_));
  NOR2  g11168(.A(new_n11553_), .B(new_n1189_), .Y(new_n11554_));
  NOR2  g11169(.A(new_n11554_), .B(new_n1707_), .Y(new_n11555_));
  NOR2  g11170(.A(new_n11555_), .B(new_n1709_), .Y(new_n11556_));
  NOR2  g11171(.A(new_n11556_), .B(new_n1973_), .Y(new_n11557_));
  NOR2  g11172(.A(new_n11557_), .B(new_n1199_), .Y(new_n11558_));
  NOR2  g11173(.A(new_n11558_), .B(new_n1203_), .Y(new_n11559_));
  NOR2  g11174(.A(new_n11559_), .B(new_n1207_), .Y(new_n11560_));
  NOR2  g11175(.A(new_n11560_), .B(new_n1211_), .Y(new_n11561_));
  NOR2  g11176(.A(new_n11561_), .B(new_n1215_), .Y(new_n11562_));
  NOR2  g11177(.A(new_n11562_), .B(new_n1219_), .Y(new_n11563_));
  NOR2  g11178(.A(new_n11563_), .B(new_n1223_), .Y(new_n11564_));
  NOR2  g11179(.A(new_n11564_), .B(new_n1227_), .Y(new_n11565_));
  NOR2  g11180(.A(new_n11565_), .B(new_n1231_), .Y(new_n11566_));
  NOR2  g11181(.A(new_n11566_), .B(new_n1235_), .Y(new_n11567_));
  NOR2  g11182(.A(new_n11567_), .B(new_n1239_), .Y(new_n11568_));
  NOR2  g11183(.A(new_n11568_), .B(new_n1243_), .Y(new_n11569_));
  NOR2  g11184(.A(new_n11569_), .B(new_n1247_), .Y(new_n11570_));
  NOR2  g11185(.A(new_n11570_), .B(new_n1251_), .Y(new_n11571_));
  NOR2  g11186(.A(new_n11571_), .B(new_n1255_), .Y(new_n11572_));
  NOR2  g11187(.A(new_n11572_), .B(new_n1259_), .Y(new_n11573_));
  NOR2  g11188(.A(new_n11573_), .B(new_n1263_), .Y(new_n11574_));
  NOR2  g11189(.A(new_n11574_), .B(new_n1267_), .Y(new_n11575_));
  NOR2  g11190(.A(new_n11575_), .B(new_n1271_), .Y(new_n11576_));
  NOR2  g11191(.A(new_n11576_), .B(new_n1275_), .Y(new_n11577_));
  NOR2  g11192(.A(new_n11577_), .B(new_n1279_), .Y(new_n11578_));
  NOR2  g11193(.A(new_n11578_), .B(new_n1283_), .Y(new_n11579_));
  NOR2  g11194(.A(new_n11579_), .B(new_n1287_), .Y(new_n11580_));
  NOR2  g11195(.A(new_n11580_), .B(new_n1291_), .Y(new_n11581_));
  NOR2  g11196(.A(new_n11581_), .B(new_n1295_), .Y(new_n11582_));
  NOR2  g11197(.A(new_n11582_), .B(new_n1299_), .Y(new_n11583_));
  NOR2  g11198(.A(new_n11583_), .B(new_n1303_), .Y(new_n11584_));
  NOR2  g11199(.A(new_n11584_), .B(new_n1307_), .Y(new_n11585_));
  NOR2  g11200(.A(new_n11585_), .B(new_n1311_), .Y(new_n11586_));
  NOR2  g11201(.A(new_n11586_), .B(new_n1315_), .Y(new_n11587_));
  NOR2  g11202(.A(new_n11587_), .B(new_n1319_), .Y(new_n11588_));
  NOR2  g11203(.A(new_n11588_), .B(new_n1323_), .Y(new_n11589_));
  NOR2  g11204(.A(new_n11589_), .B(new_n1327_), .Y(new_n11590_));
  NOR2  g11205(.A(new_n11590_), .B(new_n1331_), .Y(new_n11591_));
  NOR2  g11206(.A(new_n11591_), .B(new_n1335_), .Y(new_n11592_));
  NOR2  g11207(.A(new_n11592_), .B(new_n1339_), .Y(new_n11593_));
  NOR2  g11208(.A(new_n11593_), .B(new_n1343_), .Y(new_n11594_));
  NOR2  g11209(.A(new_n11594_), .B(new_n1347_), .Y(new_n11595_));
  NOR2  g11210(.A(new_n11595_), .B(new_n1351_), .Y(new_n11596_));
  NOR2  g11211(.A(new_n11596_), .B(new_n1355_), .Y(new_n11597_));
  NOR2  g11212(.A(new_n11597_), .B(new_n1359_), .Y(new_n11598_));
  NOR2  g11213(.A(new_n11598_), .B(new_n1363_), .Y(new_n11599_));
  NOR2  g11214(.A(new_n11599_), .B(new_n1367_), .Y(new_n11600_));
  NOR2  g11215(.A(new_n11600_), .B(new_n1371_), .Y(new_n11601_));
  NOR2  g11216(.A(new_n11601_), .B(new_n1375_), .Y(new_n11602_));
  NOR2  g11217(.A(new_n11602_), .B(new_n1379_), .Y(new_n11603_));
  NOR2  g11218(.A(new_n11603_), .B(new_n1383_), .Y(new_n11604_));
  NOR2  g11219(.A(new_n11604_), .B(new_n1387_), .Y(new_n11605_));
  NOR2  g11220(.A(new_n11605_), .B(new_n1391_), .Y(new_n11606_));
  NOR2  g11221(.A(new_n11606_), .B(new_n1395_), .Y(new_n11607_));
  NOR2  g11222(.A(new_n11607_), .B(new_n1399_), .Y(new_n11608_));
  NOR2  g11223(.A(new_n11608_), .B(new_n1403_), .Y(new_n11609_));
  NOR2  g11224(.A(new_n11609_), .B(new_n1407_), .Y(new_n11610_));
  NOR2  g11225(.A(new_n11610_), .B(new_n1411_), .Y(new_n11611_));
  NOR2  g11226(.A(new_n11611_), .B(new_n1415_), .Y(new_n11612_));
  NOR2  g11227(.A(new_n11612_), .B(new_n1419_), .Y(new_n11613_));
  NOR2  g11228(.A(new_n11613_), .B(new_n1423_), .Y(new_n11614_));
  NOR2  g11229(.A(new_n11614_), .B(new_n1427_), .Y(new_n11615_));
  NOR2  g11230(.A(new_n11615_), .B(new_n1431_), .Y(new_n11616_));
  NOR2  g11231(.A(new_n11616_), .B(new_n1435_), .Y(new_n11617_));
  NOR2  g11232(.A(new_n11617_), .B(new_n1439_), .Y(new_n11618_));
  NOR2  g11233(.A(new_n11618_), .B(new_n1443_), .Y(new_n11619_));
  NOR2  g11234(.A(new_n11619_), .B(new_n1447_), .Y(new_n11620_));
  NOR2  g11235(.A(new_n11620_), .B(new_n1451_), .Y(new_n11621_));
  NOR2  g11236(.A(new_n11621_), .B(new_n1455_), .Y(new_n11622_));
  NOR2  g11237(.A(new_n11622_), .B(new_n1459_), .Y(new_n11623_));
  NOR2  g11238(.A(new_n11623_), .B(new_n1463_), .Y(new_n11624_));
  NOR2  g11239(.A(new_n11624_), .B(new_n1467_), .Y(new_n11625_));
  NOR2  g11240(.A(new_n11625_), .B(new_n1471_), .Y(new_n11626_));
  NOR2  g11241(.A(new_n11626_), .B(new_n1475_), .Y(new_n11627_));
  NOR2  g11242(.A(new_n11627_), .B(new_n1479_), .Y(new_n11628_));
  NOR2  g11243(.A(new_n11628_), .B(new_n1483_), .Y(new_n11629_));
  NOR2  g11244(.A(new_n11629_), .B(new_n1487_), .Y(new_n11630_));
  NOR2  g11245(.A(new_n11630_), .B(new_n1491_), .Y(new_n11631_));
  NOR2  g11246(.A(new_n11631_), .B(new_n1495_), .Y(new_n11632_));
  NAND2 g11247(.A(new_n1497_), .B(\req[118] ), .Y(new_n11633_));
  NOR2  g11248(.A(new_n11633_), .B(new_n11632_), .Y(\grant[118] ));
  INV   g11249(.A(new_n1506_), .Y(new_n11635_));
  NOR2  g11250(.A(new_n11635_), .B(new_n785_), .Y(new_n11636_));
  NOR2  g11251(.A(new_n11636_), .B(new_n1511_), .Y(new_n11637_));
  NOR2  g11252(.A(new_n11637_), .B(new_n1515_), .Y(new_n11638_));
  NOR2  g11253(.A(new_n11638_), .B(new_n1519_), .Y(new_n11639_));
  NOR2  g11254(.A(new_n11639_), .B(new_n1523_), .Y(new_n11640_));
  NOR2  g11255(.A(new_n11640_), .B(new_n1527_), .Y(new_n11641_));
  NOR2  g11256(.A(new_n11641_), .B(new_n1797_), .Y(new_n11642_));
  NOR2  g11257(.A(new_n11642_), .B(new_n396_), .Y(new_n11643_));
  NOR2  g11258(.A(new_n11643_), .B(new_n400_), .Y(new_n11644_));
  NOR2  g11259(.A(new_n11644_), .B(new_n406_), .Y(new_n11645_));
  NOR2  g11260(.A(new_n11645_), .B(new_n410_), .Y(new_n11646_));
  NOR2  g11261(.A(new_n11646_), .B(new_n416_), .Y(new_n11647_));
  NOR2  g11262(.A(new_n11647_), .B(new_n420_), .Y(new_n11648_));
  NOR2  g11263(.A(new_n11648_), .B(new_n426_), .Y(new_n11649_));
  NOR2  g11264(.A(new_n11649_), .B(new_n430_), .Y(new_n11650_));
  NOR2  g11265(.A(new_n11650_), .B(new_n436_), .Y(new_n11651_));
  NOR2  g11266(.A(new_n11651_), .B(new_n440_), .Y(new_n11652_));
  NOR2  g11267(.A(new_n11652_), .B(new_n446_), .Y(new_n11653_));
  NOR2  g11268(.A(new_n11653_), .B(new_n450_), .Y(new_n11654_));
  NOR2  g11269(.A(new_n11654_), .B(new_n456_), .Y(new_n11655_));
  NOR2  g11270(.A(new_n11655_), .B(new_n460_), .Y(new_n11656_));
  NOR2  g11271(.A(new_n11656_), .B(new_n466_), .Y(new_n11657_));
  NOR2  g11272(.A(new_n11657_), .B(new_n470_), .Y(new_n11658_));
  NOR2  g11273(.A(new_n11658_), .B(new_n476_), .Y(new_n11659_));
  NOR2  g11274(.A(new_n11659_), .B(new_n480_), .Y(new_n11660_));
  NOR2  g11275(.A(new_n11660_), .B(new_n486_), .Y(new_n11661_));
  NOR2  g11276(.A(new_n11661_), .B(new_n490_), .Y(new_n11662_));
  NOR2  g11277(.A(new_n11662_), .B(new_n496_), .Y(new_n11663_));
  NOR2  g11278(.A(new_n11663_), .B(new_n500_), .Y(new_n11664_));
  NOR2  g11279(.A(new_n11664_), .B(new_n506_), .Y(new_n11665_));
  NOR2  g11280(.A(new_n11665_), .B(new_n510_), .Y(new_n11666_));
  NOR2  g11281(.A(new_n11666_), .B(new_n516_), .Y(new_n11667_));
  NOR2  g11282(.A(new_n11667_), .B(new_n520_), .Y(new_n11668_));
  NOR2  g11283(.A(new_n11668_), .B(new_n526_), .Y(new_n11669_));
  NOR2  g11284(.A(new_n11669_), .B(new_n530_), .Y(new_n11670_));
  NOR2  g11285(.A(new_n11670_), .B(new_n536_), .Y(new_n11671_));
  NOR2  g11286(.A(new_n11671_), .B(new_n540_), .Y(new_n11672_));
  NOR2  g11287(.A(new_n11672_), .B(new_n546_), .Y(new_n11673_));
  NOR2  g11288(.A(new_n11673_), .B(new_n550_), .Y(new_n11674_));
  NOR2  g11289(.A(new_n11674_), .B(new_n556_), .Y(new_n11675_));
  NOR2  g11290(.A(new_n11675_), .B(new_n560_), .Y(new_n11676_));
  NOR2  g11291(.A(new_n11676_), .B(new_n566_), .Y(new_n11677_));
  NOR2  g11292(.A(new_n11677_), .B(new_n570_), .Y(new_n11678_));
  NOR2  g11293(.A(new_n11678_), .B(new_n576_), .Y(new_n11679_));
  NOR2  g11294(.A(new_n11679_), .B(new_n580_), .Y(new_n11680_));
  NOR2  g11295(.A(new_n11680_), .B(new_n586_), .Y(new_n11681_));
  NOR2  g11296(.A(new_n11681_), .B(new_n590_), .Y(new_n11682_));
  NOR2  g11297(.A(new_n11682_), .B(new_n596_), .Y(new_n11683_));
  NOR2  g11298(.A(new_n11683_), .B(new_n600_), .Y(new_n11684_));
  NOR2  g11299(.A(new_n11684_), .B(new_n606_), .Y(new_n11685_));
  NOR2  g11300(.A(new_n11685_), .B(new_n610_), .Y(new_n11686_));
  NOR2  g11301(.A(new_n11686_), .B(new_n616_), .Y(new_n11687_));
  NOR2  g11302(.A(new_n11687_), .B(new_n620_), .Y(new_n11688_));
  NOR2  g11303(.A(new_n11688_), .B(new_n626_), .Y(new_n11689_));
  NOR2  g11304(.A(new_n11689_), .B(new_n630_), .Y(new_n11690_));
  NOR2  g11305(.A(new_n11690_), .B(new_n636_), .Y(new_n11691_));
  NOR2  g11306(.A(new_n11691_), .B(new_n640_), .Y(new_n11692_));
  NOR2  g11307(.A(new_n11692_), .B(new_n646_), .Y(new_n11693_));
  NOR2  g11308(.A(new_n11693_), .B(new_n650_), .Y(new_n11694_));
  NOR2  g11309(.A(new_n11694_), .B(new_n656_), .Y(new_n11695_));
  NOR2  g11310(.A(new_n11695_), .B(new_n660_), .Y(new_n11696_));
  NOR2  g11311(.A(new_n11696_), .B(new_n666_), .Y(new_n11697_));
  NOR2  g11312(.A(new_n11697_), .B(new_n670_), .Y(new_n11698_));
  NOR2  g11313(.A(new_n11698_), .B(new_n676_), .Y(new_n11699_));
  NOR2  g11314(.A(new_n11699_), .B(new_n680_), .Y(new_n11700_));
  NOR2  g11315(.A(new_n11700_), .B(new_n686_), .Y(new_n11701_));
  NOR2  g11316(.A(new_n11701_), .B(new_n690_), .Y(new_n11702_));
  NOR2  g11317(.A(new_n11702_), .B(new_n696_), .Y(new_n11703_));
  NOR2  g11318(.A(new_n11703_), .B(new_n700_), .Y(new_n11704_));
  NOR2  g11319(.A(new_n11704_), .B(new_n706_), .Y(new_n11705_));
  NOR2  g11320(.A(new_n11705_), .B(new_n710_), .Y(new_n11706_));
  NOR2  g11321(.A(new_n11706_), .B(new_n716_), .Y(new_n11707_));
  NOR2  g11322(.A(new_n11707_), .B(new_n720_), .Y(new_n11708_));
  NOR2  g11323(.A(new_n11708_), .B(new_n726_), .Y(new_n11709_));
  NOR2  g11324(.A(new_n11709_), .B(new_n730_), .Y(new_n11710_));
  NOR2  g11325(.A(new_n11710_), .B(new_n736_), .Y(new_n11711_));
  NOR2  g11326(.A(new_n11711_), .B(new_n740_), .Y(new_n11712_));
  NOR2  g11327(.A(new_n11712_), .B(new_n746_), .Y(new_n11713_));
  NOR2  g11328(.A(new_n11713_), .B(new_n750_), .Y(new_n11714_));
  NOR2  g11329(.A(new_n11714_), .B(new_n756_), .Y(new_n11715_));
  NOR2  g11330(.A(new_n11715_), .B(new_n760_), .Y(new_n11716_));
  NOR2  g11331(.A(new_n11716_), .B(new_n766_), .Y(new_n11717_));
  NOR2  g11332(.A(new_n11717_), .B(new_n770_), .Y(new_n11718_));
  NOR2  g11333(.A(new_n11718_), .B(new_n776_), .Y(new_n11719_));
  NAND2 g11334(.A(new_n778_), .B(\req[119] ), .Y(new_n11720_));
  NOR2  g11335(.A(new_n11720_), .B(new_n11719_), .Y(\grant[119] ));
  INV   g11336(.A(new_n789_), .Y(new_n11722_));
  NOR2  g11337(.A(new_n1170_), .B(new_n11722_), .Y(new_n11723_));
  NOR2  g11338(.A(new_n11723_), .B(new_n796_), .Y(new_n11724_));
  NOR2  g11339(.A(new_n11724_), .B(new_n800_), .Y(new_n11725_));
  NOR2  g11340(.A(new_n11725_), .B(new_n806_), .Y(new_n11726_));
  NOR2  g11341(.A(new_n11726_), .B(new_n1616_), .Y(new_n11727_));
  NOR2  g11342(.A(new_n11727_), .B(new_n1618_), .Y(new_n11728_));
  NOR2  g11343(.A(new_n11728_), .B(new_n1885_), .Y(new_n11729_));
  NOR2  g11344(.A(new_n11729_), .B(new_n820_), .Y(new_n11730_));
  NOR2  g11345(.A(new_n11730_), .B(new_n824_), .Y(new_n11731_));
  NOR2  g11346(.A(new_n11731_), .B(new_n829_), .Y(new_n11732_));
  NOR2  g11347(.A(new_n11732_), .B(new_n833_), .Y(new_n11733_));
  NOR2  g11348(.A(new_n11733_), .B(new_n838_), .Y(new_n11734_));
  NOR2  g11349(.A(new_n11734_), .B(new_n842_), .Y(new_n11735_));
  NOR2  g11350(.A(new_n11735_), .B(new_n847_), .Y(new_n11736_));
  NOR2  g11351(.A(new_n11736_), .B(new_n851_), .Y(new_n11737_));
  NOR2  g11352(.A(new_n11737_), .B(new_n856_), .Y(new_n11738_));
  NOR2  g11353(.A(new_n11738_), .B(new_n860_), .Y(new_n11739_));
  NOR2  g11354(.A(new_n11739_), .B(new_n865_), .Y(new_n11740_));
  NOR2  g11355(.A(new_n11740_), .B(new_n869_), .Y(new_n11741_));
  NOR2  g11356(.A(new_n11741_), .B(new_n874_), .Y(new_n11742_));
  NOR2  g11357(.A(new_n11742_), .B(new_n878_), .Y(new_n11743_));
  NOR2  g11358(.A(new_n11743_), .B(new_n883_), .Y(new_n11744_));
  NOR2  g11359(.A(new_n11744_), .B(new_n887_), .Y(new_n11745_));
  NOR2  g11360(.A(new_n11745_), .B(new_n892_), .Y(new_n11746_));
  NOR2  g11361(.A(new_n11746_), .B(new_n896_), .Y(new_n11747_));
  NOR2  g11362(.A(new_n11747_), .B(new_n901_), .Y(new_n11748_));
  NOR2  g11363(.A(new_n11748_), .B(new_n905_), .Y(new_n11749_));
  NOR2  g11364(.A(new_n11749_), .B(new_n910_), .Y(new_n11750_));
  NOR2  g11365(.A(new_n11750_), .B(new_n914_), .Y(new_n11751_));
  NOR2  g11366(.A(new_n11751_), .B(new_n919_), .Y(new_n11752_));
  NOR2  g11367(.A(new_n11752_), .B(new_n923_), .Y(new_n11753_));
  NOR2  g11368(.A(new_n11753_), .B(new_n928_), .Y(new_n11754_));
  NOR2  g11369(.A(new_n11754_), .B(new_n932_), .Y(new_n11755_));
  NOR2  g11370(.A(new_n11755_), .B(new_n937_), .Y(new_n11756_));
  NOR2  g11371(.A(new_n11756_), .B(new_n941_), .Y(new_n11757_));
  NOR2  g11372(.A(new_n11757_), .B(new_n946_), .Y(new_n11758_));
  NOR2  g11373(.A(new_n11758_), .B(new_n950_), .Y(new_n11759_));
  NOR2  g11374(.A(new_n11759_), .B(new_n955_), .Y(new_n11760_));
  NOR2  g11375(.A(new_n11760_), .B(new_n959_), .Y(new_n11761_));
  NOR2  g11376(.A(new_n11761_), .B(new_n964_), .Y(new_n11762_));
  NOR2  g11377(.A(new_n11762_), .B(new_n968_), .Y(new_n11763_));
  NOR2  g11378(.A(new_n11763_), .B(new_n973_), .Y(new_n11764_));
  NOR2  g11379(.A(new_n11764_), .B(new_n977_), .Y(new_n11765_));
  NOR2  g11380(.A(new_n11765_), .B(new_n982_), .Y(new_n11766_));
  NOR2  g11381(.A(new_n11766_), .B(new_n986_), .Y(new_n11767_));
  NOR2  g11382(.A(new_n11767_), .B(new_n991_), .Y(new_n11768_));
  NOR2  g11383(.A(new_n11768_), .B(new_n995_), .Y(new_n11769_));
  NOR2  g11384(.A(new_n11769_), .B(new_n1000_), .Y(new_n11770_));
  NOR2  g11385(.A(new_n11770_), .B(new_n1004_), .Y(new_n11771_));
  NOR2  g11386(.A(new_n11771_), .B(new_n1009_), .Y(new_n11772_));
  NOR2  g11387(.A(new_n11772_), .B(new_n1013_), .Y(new_n11773_));
  NOR2  g11388(.A(new_n11773_), .B(new_n1018_), .Y(new_n11774_));
  NOR2  g11389(.A(new_n11774_), .B(new_n1022_), .Y(new_n11775_));
  NOR2  g11390(.A(new_n11775_), .B(new_n1027_), .Y(new_n11776_));
  NOR2  g11391(.A(new_n11776_), .B(new_n1031_), .Y(new_n11777_));
  NOR2  g11392(.A(new_n11777_), .B(new_n1036_), .Y(new_n11778_));
  NOR2  g11393(.A(new_n11778_), .B(new_n1040_), .Y(new_n11779_));
  NOR2  g11394(.A(new_n11779_), .B(new_n1045_), .Y(new_n11780_));
  NOR2  g11395(.A(new_n11780_), .B(new_n1049_), .Y(new_n11781_));
  NOR2  g11396(.A(new_n11781_), .B(new_n1054_), .Y(new_n11782_));
  NOR2  g11397(.A(new_n11782_), .B(new_n1058_), .Y(new_n11783_));
  NOR2  g11398(.A(new_n11783_), .B(new_n1063_), .Y(new_n11784_));
  NOR2  g11399(.A(new_n11784_), .B(new_n1067_), .Y(new_n11785_));
  NOR2  g11400(.A(new_n11785_), .B(new_n1072_), .Y(new_n11786_));
  NOR2  g11401(.A(new_n11786_), .B(new_n1076_), .Y(new_n11787_));
  NOR2  g11402(.A(new_n11787_), .B(new_n1081_), .Y(new_n11788_));
  NOR2  g11403(.A(new_n11788_), .B(new_n1085_), .Y(new_n11789_));
  NOR2  g11404(.A(new_n11789_), .B(new_n1090_), .Y(new_n11790_));
  NOR2  g11405(.A(new_n11790_), .B(new_n1094_), .Y(new_n11791_));
  NOR2  g11406(.A(new_n11791_), .B(new_n1099_), .Y(new_n11792_));
  NOR2  g11407(.A(new_n11792_), .B(new_n1103_), .Y(new_n11793_));
  NOR2  g11408(.A(new_n11793_), .B(new_n1108_), .Y(new_n11794_));
  NOR2  g11409(.A(new_n11794_), .B(new_n1112_), .Y(new_n11795_));
  NOR2  g11410(.A(new_n11795_), .B(new_n1117_), .Y(new_n11796_));
  NOR2  g11411(.A(new_n11796_), .B(new_n1121_), .Y(new_n11797_));
  NOR2  g11412(.A(new_n11797_), .B(new_n1126_), .Y(new_n11798_));
  NOR2  g11413(.A(new_n11798_), .B(new_n1130_), .Y(new_n11799_));
  NOR2  g11414(.A(new_n11799_), .B(new_n1135_), .Y(new_n11800_));
  NOR2  g11415(.A(new_n11800_), .B(new_n1139_), .Y(new_n11801_));
  NOR2  g11416(.A(new_n11801_), .B(new_n1144_), .Y(new_n11802_));
  NOR2  g11417(.A(new_n11802_), .B(new_n1148_), .Y(new_n11803_));
  NOR2  g11418(.A(new_n11803_), .B(new_n1153_), .Y(new_n11804_));
  NOR2  g11419(.A(new_n11804_), .B(new_n1157_), .Y(new_n11805_));
  NOR2  g11420(.A(new_n11805_), .B(new_n1162_), .Y(new_n11806_));
  NAND2 g11421(.A(new_n1164_), .B(\req[120] ), .Y(new_n11807_));
  NOR2  g11422(.A(new_n11807_), .B(new_n11806_), .Y(\grant[120] ));
  INV   g11423(.A(new_n1174_), .Y(new_n11809_));
  NOR2  g11424(.A(new_n1510_), .B(new_n11809_), .Y(new_n11810_));
  NOR2  g11425(.A(new_n11810_), .B(new_n1180_), .Y(new_n11811_));
  NOR2  g11426(.A(new_n11811_), .B(new_n1184_), .Y(new_n11812_));
  NOR2  g11427(.A(new_n11812_), .B(new_n1189_), .Y(new_n11813_));
  NOR2  g11428(.A(new_n11813_), .B(new_n1707_), .Y(new_n11814_));
  NOR2  g11429(.A(new_n11814_), .B(new_n1709_), .Y(new_n11815_));
  NOR2  g11430(.A(new_n11815_), .B(new_n1973_), .Y(new_n11816_));
  NOR2  g11431(.A(new_n11816_), .B(new_n1199_), .Y(new_n11817_));
  NOR2  g11432(.A(new_n11817_), .B(new_n1203_), .Y(new_n11818_));
  NOR2  g11433(.A(new_n11818_), .B(new_n1207_), .Y(new_n11819_));
  NOR2  g11434(.A(new_n11819_), .B(new_n1211_), .Y(new_n11820_));
  NOR2  g11435(.A(new_n11820_), .B(new_n1215_), .Y(new_n11821_));
  NOR2  g11436(.A(new_n11821_), .B(new_n1219_), .Y(new_n11822_));
  NOR2  g11437(.A(new_n11822_), .B(new_n1223_), .Y(new_n11823_));
  NOR2  g11438(.A(new_n11823_), .B(new_n1227_), .Y(new_n11824_));
  NOR2  g11439(.A(new_n11824_), .B(new_n1231_), .Y(new_n11825_));
  NOR2  g11440(.A(new_n11825_), .B(new_n1235_), .Y(new_n11826_));
  NOR2  g11441(.A(new_n11826_), .B(new_n1239_), .Y(new_n11827_));
  NOR2  g11442(.A(new_n11827_), .B(new_n1243_), .Y(new_n11828_));
  NOR2  g11443(.A(new_n11828_), .B(new_n1247_), .Y(new_n11829_));
  NOR2  g11444(.A(new_n11829_), .B(new_n1251_), .Y(new_n11830_));
  NOR2  g11445(.A(new_n11830_), .B(new_n1255_), .Y(new_n11831_));
  NOR2  g11446(.A(new_n11831_), .B(new_n1259_), .Y(new_n11832_));
  NOR2  g11447(.A(new_n11832_), .B(new_n1263_), .Y(new_n11833_));
  NOR2  g11448(.A(new_n11833_), .B(new_n1267_), .Y(new_n11834_));
  NOR2  g11449(.A(new_n11834_), .B(new_n1271_), .Y(new_n11835_));
  NOR2  g11450(.A(new_n11835_), .B(new_n1275_), .Y(new_n11836_));
  NOR2  g11451(.A(new_n11836_), .B(new_n1279_), .Y(new_n11837_));
  NOR2  g11452(.A(new_n11837_), .B(new_n1283_), .Y(new_n11838_));
  NOR2  g11453(.A(new_n11838_), .B(new_n1287_), .Y(new_n11839_));
  NOR2  g11454(.A(new_n11839_), .B(new_n1291_), .Y(new_n11840_));
  NOR2  g11455(.A(new_n11840_), .B(new_n1295_), .Y(new_n11841_));
  NOR2  g11456(.A(new_n11841_), .B(new_n1299_), .Y(new_n11842_));
  NOR2  g11457(.A(new_n11842_), .B(new_n1303_), .Y(new_n11843_));
  NOR2  g11458(.A(new_n11843_), .B(new_n1307_), .Y(new_n11844_));
  NOR2  g11459(.A(new_n11844_), .B(new_n1311_), .Y(new_n11845_));
  NOR2  g11460(.A(new_n11845_), .B(new_n1315_), .Y(new_n11846_));
  NOR2  g11461(.A(new_n11846_), .B(new_n1319_), .Y(new_n11847_));
  NOR2  g11462(.A(new_n11847_), .B(new_n1323_), .Y(new_n11848_));
  NOR2  g11463(.A(new_n11848_), .B(new_n1327_), .Y(new_n11849_));
  NOR2  g11464(.A(new_n11849_), .B(new_n1331_), .Y(new_n11850_));
  NOR2  g11465(.A(new_n11850_), .B(new_n1335_), .Y(new_n11851_));
  NOR2  g11466(.A(new_n11851_), .B(new_n1339_), .Y(new_n11852_));
  NOR2  g11467(.A(new_n11852_), .B(new_n1343_), .Y(new_n11853_));
  NOR2  g11468(.A(new_n11853_), .B(new_n1347_), .Y(new_n11854_));
  NOR2  g11469(.A(new_n11854_), .B(new_n1351_), .Y(new_n11855_));
  NOR2  g11470(.A(new_n11855_), .B(new_n1355_), .Y(new_n11856_));
  NOR2  g11471(.A(new_n11856_), .B(new_n1359_), .Y(new_n11857_));
  NOR2  g11472(.A(new_n11857_), .B(new_n1363_), .Y(new_n11858_));
  NOR2  g11473(.A(new_n11858_), .B(new_n1367_), .Y(new_n11859_));
  NOR2  g11474(.A(new_n11859_), .B(new_n1371_), .Y(new_n11860_));
  NOR2  g11475(.A(new_n11860_), .B(new_n1375_), .Y(new_n11861_));
  NOR2  g11476(.A(new_n11861_), .B(new_n1379_), .Y(new_n11862_));
  NOR2  g11477(.A(new_n11862_), .B(new_n1383_), .Y(new_n11863_));
  NOR2  g11478(.A(new_n11863_), .B(new_n1387_), .Y(new_n11864_));
  NOR2  g11479(.A(new_n11864_), .B(new_n1391_), .Y(new_n11865_));
  NOR2  g11480(.A(new_n11865_), .B(new_n1395_), .Y(new_n11866_));
  NOR2  g11481(.A(new_n11866_), .B(new_n1399_), .Y(new_n11867_));
  NOR2  g11482(.A(new_n11867_), .B(new_n1403_), .Y(new_n11868_));
  NOR2  g11483(.A(new_n11868_), .B(new_n1407_), .Y(new_n11869_));
  NOR2  g11484(.A(new_n11869_), .B(new_n1411_), .Y(new_n11870_));
  NOR2  g11485(.A(new_n11870_), .B(new_n1415_), .Y(new_n11871_));
  NOR2  g11486(.A(new_n11871_), .B(new_n1419_), .Y(new_n11872_));
  NOR2  g11487(.A(new_n11872_), .B(new_n1423_), .Y(new_n11873_));
  NOR2  g11488(.A(new_n11873_), .B(new_n1427_), .Y(new_n11874_));
  NOR2  g11489(.A(new_n11874_), .B(new_n1431_), .Y(new_n11875_));
  NOR2  g11490(.A(new_n11875_), .B(new_n1435_), .Y(new_n11876_));
  NOR2  g11491(.A(new_n11876_), .B(new_n1439_), .Y(new_n11877_));
  NOR2  g11492(.A(new_n11877_), .B(new_n1443_), .Y(new_n11878_));
  NOR2  g11493(.A(new_n11878_), .B(new_n1447_), .Y(new_n11879_));
  NOR2  g11494(.A(new_n11879_), .B(new_n1451_), .Y(new_n11880_));
  NOR2  g11495(.A(new_n11880_), .B(new_n1455_), .Y(new_n11881_));
  NOR2  g11496(.A(new_n11881_), .B(new_n1459_), .Y(new_n11882_));
  NOR2  g11497(.A(new_n11882_), .B(new_n1463_), .Y(new_n11883_));
  NOR2  g11498(.A(new_n11883_), .B(new_n1467_), .Y(new_n11884_));
  NOR2  g11499(.A(new_n11884_), .B(new_n1471_), .Y(new_n11885_));
  NOR2  g11500(.A(new_n11885_), .B(new_n1475_), .Y(new_n11886_));
  NOR2  g11501(.A(new_n11886_), .B(new_n1479_), .Y(new_n11887_));
  NOR2  g11502(.A(new_n11887_), .B(new_n1483_), .Y(new_n11888_));
  NOR2  g11503(.A(new_n11888_), .B(new_n1487_), .Y(new_n11889_));
  NOR2  g11504(.A(new_n11889_), .B(new_n1491_), .Y(new_n11890_));
  NOR2  g11505(.A(new_n11890_), .B(new_n1495_), .Y(new_n11891_));
  NOR2  g11506(.A(new_n11891_), .B(new_n1499_), .Y(new_n11892_));
  NOR2  g11507(.A(new_n11892_), .B(new_n1503_), .Y(new_n11893_));
  NAND2 g11508(.A(new_n1505_), .B(\req[121] ), .Y(new_n11894_));
  NOR2  g11509(.A(new_n11894_), .B(new_n11893_), .Y(\grant[121] ));
  INV   g11510(.A(new_n1514_), .Y(new_n11896_));
  NOR2  g11511(.A(new_n11896_), .B(new_n795_), .Y(new_n11897_));
  NOR2  g11512(.A(new_n11897_), .B(new_n1519_), .Y(new_n11898_));
  NOR2  g11513(.A(new_n11898_), .B(new_n1523_), .Y(new_n11899_));
  NOR2  g11514(.A(new_n11899_), .B(new_n1527_), .Y(new_n11900_));
  NOR2  g11515(.A(new_n11900_), .B(new_n1797_), .Y(new_n11901_));
  NOR2  g11516(.A(new_n11901_), .B(new_n396_), .Y(new_n11902_));
  NOR2  g11517(.A(new_n11902_), .B(new_n400_), .Y(new_n11903_));
  NOR2  g11518(.A(new_n11903_), .B(new_n406_), .Y(new_n11904_));
  NOR2  g11519(.A(new_n11904_), .B(new_n410_), .Y(new_n11905_));
  NOR2  g11520(.A(new_n11905_), .B(new_n416_), .Y(new_n11906_));
  NOR2  g11521(.A(new_n11906_), .B(new_n420_), .Y(new_n11907_));
  NOR2  g11522(.A(new_n11907_), .B(new_n426_), .Y(new_n11908_));
  NOR2  g11523(.A(new_n11908_), .B(new_n430_), .Y(new_n11909_));
  NOR2  g11524(.A(new_n11909_), .B(new_n436_), .Y(new_n11910_));
  NOR2  g11525(.A(new_n11910_), .B(new_n440_), .Y(new_n11911_));
  NOR2  g11526(.A(new_n11911_), .B(new_n446_), .Y(new_n11912_));
  NOR2  g11527(.A(new_n11912_), .B(new_n450_), .Y(new_n11913_));
  NOR2  g11528(.A(new_n11913_), .B(new_n456_), .Y(new_n11914_));
  NOR2  g11529(.A(new_n11914_), .B(new_n460_), .Y(new_n11915_));
  NOR2  g11530(.A(new_n11915_), .B(new_n466_), .Y(new_n11916_));
  NOR2  g11531(.A(new_n11916_), .B(new_n470_), .Y(new_n11917_));
  NOR2  g11532(.A(new_n11917_), .B(new_n476_), .Y(new_n11918_));
  NOR2  g11533(.A(new_n11918_), .B(new_n480_), .Y(new_n11919_));
  NOR2  g11534(.A(new_n11919_), .B(new_n486_), .Y(new_n11920_));
  NOR2  g11535(.A(new_n11920_), .B(new_n490_), .Y(new_n11921_));
  NOR2  g11536(.A(new_n11921_), .B(new_n496_), .Y(new_n11922_));
  NOR2  g11537(.A(new_n11922_), .B(new_n500_), .Y(new_n11923_));
  NOR2  g11538(.A(new_n11923_), .B(new_n506_), .Y(new_n11924_));
  NOR2  g11539(.A(new_n11924_), .B(new_n510_), .Y(new_n11925_));
  NOR2  g11540(.A(new_n11925_), .B(new_n516_), .Y(new_n11926_));
  NOR2  g11541(.A(new_n11926_), .B(new_n520_), .Y(new_n11927_));
  NOR2  g11542(.A(new_n11927_), .B(new_n526_), .Y(new_n11928_));
  NOR2  g11543(.A(new_n11928_), .B(new_n530_), .Y(new_n11929_));
  NOR2  g11544(.A(new_n11929_), .B(new_n536_), .Y(new_n11930_));
  NOR2  g11545(.A(new_n11930_), .B(new_n540_), .Y(new_n11931_));
  NOR2  g11546(.A(new_n11931_), .B(new_n546_), .Y(new_n11932_));
  NOR2  g11547(.A(new_n11932_), .B(new_n550_), .Y(new_n11933_));
  NOR2  g11548(.A(new_n11933_), .B(new_n556_), .Y(new_n11934_));
  NOR2  g11549(.A(new_n11934_), .B(new_n560_), .Y(new_n11935_));
  NOR2  g11550(.A(new_n11935_), .B(new_n566_), .Y(new_n11936_));
  NOR2  g11551(.A(new_n11936_), .B(new_n570_), .Y(new_n11937_));
  NOR2  g11552(.A(new_n11937_), .B(new_n576_), .Y(new_n11938_));
  NOR2  g11553(.A(new_n11938_), .B(new_n580_), .Y(new_n11939_));
  NOR2  g11554(.A(new_n11939_), .B(new_n586_), .Y(new_n11940_));
  NOR2  g11555(.A(new_n11940_), .B(new_n590_), .Y(new_n11941_));
  NOR2  g11556(.A(new_n11941_), .B(new_n596_), .Y(new_n11942_));
  NOR2  g11557(.A(new_n11942_), .B(new_n600_), .Y(new_n11943_));
  NOR2  g11558(.A(new_n11943_), .B(new_n606_), .Y(new_n11944_));
  NOR2  g11559(.A(new_n11944_), .B(new_n610_), .Y(new_n11945_));
  NOR2  g11560(.A(new_n11945_), .B(new_n616_), .Y(new_n11946_));
  NOR2  g11561(.A(new_n11946_), .B(new_n620_), .Y(new_n11947_));
  NOR2  g11562(.A(new_n11947_), .B(new_n626_), .Y(new_n11948_));
  NOR2  g11563(.A(new_n11948_), .B(new_n630_), .Y(new_n11949_));
  NOR2  g11564(.A(new_n11949_), .B(new_n636_), .Y(new_n11950_));
  NOR2  g11565(.A(new_n11950_), .B(new_n640_), .Y(new_n11951_));
  NOR2  g11566(.A(new_n11951_), .B(new_n646_), .Y(new_n11952_));
  NOR2  g11567(.A(new_n11952_), .B(new_n650_), .Y(new_n11953_));
  NOR2  g11568(.A(new_n11953_), .B(new_n656_), .Y(new_n11954_));
  NOR2  g11569(.A(new_n11954_), .B(new_n660_), .Y(new_n11955_));
  NOR2  g11570(.A(new_n11955_), .B(new_n666_), .Y(new_n11956_));
  NOR2  g11571(.A(new_n11956_), .B(new_n670_), .Y(new_n11957_));
  NOR2  g11572(.A(new_n11957_), .B(new_n676_), .Y(new_n11958_));
  NOR2  g11573(.A(new_n11958_), .B(new_n680_), .Y(new_n11959_));
  NOR2  g11574(.A(new_n11959_), .B(new_n686_), .Y(new_n11960_));
  NOR2  g11575(.A(new_n11960_), .B(new_n690_), .Y(new_n11961_));
  NOR2  g11576(.A(new_n11961_), .B(new_n696_), .Y(new_n11962_));
  NOR2  g11577(.A(new_n11962_), .B(new_n700_), .Y(new_n11963_));
  NOR2  g11578(.A(new_n11963_), .B(new_n706_), .Y(new_n11964_));
  NOR2  g11579(.A(new_n11964_), .B(new_n710_), .Y(new_n11965_));
  NOR2  g11580(.A(new_n11965_), .B(new_n716_), .Y(new_n11966_));
  NOR2  g11581(.A(new_n11966_), .B(new_n720_), .Y(new_n11967_));
  NOR2  g11582(.A(new_n11967_), .B(new_n726_), .Y(new_n11968_));
  NOR2  g11583(.A(new_n11968_), .B(new_n730_), .Y(new_n11969_));
  NOR2  g11584(.A(new_n11969_), .B(new_n736_), .Y(new_n11970_));
  NOR2  g11585(.A(new_n11970_), .B(new_n740_), .Y(new_n11971_));
  NOR2  g11586(.A(new_n11971_), .B(new_n746_), .Y(new_n11972_));
  NOR2  g11587(.A(new_n11972_), .B(new_n750_), .Y(new_n11973_));
  NOR2  g11588(.A(new_n11973_), .B(new_n756_), .Y(new_n11974_));
  NOR2  g11589(.A(new_n11974_), .B(new_n760_), .Y(new_n11975_));
  NOR2  g11590(.A(new_n11975_), .B(new_n766_), .Y(new_n11976_));
  NOR2  g11591(.A(new_n11976_), .B(new_n770_), .Y(new_n11977_));
  NOR2  g11592(.A(new_n11977_), .B(new_n776_), .Y(new_n11978_));
  NOR2  g11593(.A(new_n11978_), .B(new_n780_), .Y(new_n11979_));
  NOR2  g11594(.A(new_n11979_), .B(new_n786_), .Y(new_n11980_));
  NAND2 g11595(.A(new_n788_), .B(\req[122] ), .Y(new_n11981_));
  NOR2  g11596(.A(new_n11981_), .B(new_n11980_), .Y(\grant[122] ));
  INV   g11597(.A(new_n799_), .Y(new_n11983_));
  NOR2  g11598(.A(new_n1179_), .B(new_n11983_), .Y(new_n11984_));
  NOR2  g11599(.A(new_n11984_), .B(new_n806_), .Y(new_n11985_));
  NOR2  g11600(.A(new_n11985_), .B(new_n1616_), .Y(new_n11986_));
  NOR2  g11601(.A(new_n11986_), .B(new_n1618_), .Y(new_n11987_));
  NOR2  g11602(.A(new_n11987_), .B(new_n1885_), .Y(new_n11988_));
  NOR2  g11603(.A(new_n11988_), .B(new_n820_), .Y(new_n11989_));
  NOR2  g11604(.A(new_n11989_), .B(new_n824_), .Y(new_n11990_));
  NOR2  g11605(.A(new_n11990_), .B(new_n829_), .Y(new_n11991_));
  NOR2  g11606(.A(new_n11991_), .B(new_n833_), .Y(new_n11992_));
  NOR2  g11607(.A(new_n11992_), .B(new_n838_), .Y(new_n11993_));
  NOR2  g11608(.A(new_n11993_), .B(new_n842_), .Y(new_n11994_));
  NOR2  g11609(.A(new_n11994_), .B(new_n847_), .Y(new_n11995_));
  NOR2  g11610(.A(new_n11995_), .B(new_n851_), .Y(new_n11996_));
  NOR2  g11611(.A(new_n11996_), .B(new_n856_), .Y(new_n11997_));
  NOR2  g11612(.A(new_n11997_), .B(new_n860_), .Y(new_n11998_));
  NOR2  g11613(.A(new_n11998_), .B(new_n865_), .Y(new_n11999_));
  NOR2  g11614(.A(new_n11999_), .B(new_n869_), .Y(new_n12000_));
  NOR2  g11615(.A(new_n12000_), .B(new_n874_), .Y(new_n12001_));
  NOR2  g11616(.A(new_n12001_), .B(new_n878_), .Y(new_n12002_));
  NOR2  g11617(.A(new_n12002_), .B(new_n883_), .Y(new_n12003_));
  NOR2  g11618(.A(new_n12003_), .B(new_n887_), .Y(new_n12004_));
  NOR2  g11619(.A(new_n12004_), .B(new_n892_), .Y(new_n12005_));
  NOR2  g11620(.A(new_n12005_), .B(new_n896_), .Y(new_n12006_));
  NOR2  g11621(.A(new_n12006_), .B(new_n901_), .Y(new_n12007_));
  NOR2  g11622(.A(new_n12007_), .B(new_n905_), .Y(new_n12008_));
  NOR2  g11623(.A(new_n12008_), .B(new_n910_), .Y(new_n12009_));
  NOR2  g11624(.A(new_n12009_), .B(new_n914_), .Y(new_n12010_));
  NOR2  g11625(.A(new_n12010_), .B(new_n919_), .Y(new_n12011_));
  NOR2  g11626(.A(new_n12011_), .B(new_n923_), .Y(new_n12012_));
  NOR2  g11627(.A(new_n12012_), .B(new_n928_), .Y(new_n12013_));
  NOR2  g11628(.A(new_n12013_), .B(new_n932_), .Y(new_n12014_));
  NOR2  g11629(.A(new_n12014_), .B(new_n937_), .Y(new_n12015_));
  NOR2  g11630(.A(new_n12015_), .B(new_n941_), .Y(new_n12016_));
  NOR2  g11631(.A(new_n12016_), .B(new_n946_), .Y(new_n12017_));
  NOR2  g11632(.A(new_n12017_), .B(new_n950_), .Y(new_n12018_));
  NOR2  g11633(.A(new_n12018_), .B(new_n955_), .Y(new_n12019_));
  NOR2  g11634(.A(new_n12019_), .B(new_n959_), .Y(new_n12020_));
  NOR2  g11635(.A(new_n12020_), .B(new_n964_), .Y(new_n12021_));
  NOR2  g11636(.A(new_n12021_), .B(new_n968_), .Y(new_n12022_));
  NOR2  g11637(.A(new_n12022_), .B(new_n973_), .Y(new_n12023_));
  NOR2  g11638(.A(new_n12023_), .B(new_n977_), .Y(new_n12024_));
  NOR2  g11639(.A(new_n12024_), .B(new_n982_), .Y(new_n12025_));
  NOR2  g11640(.A(new_n12025_), .B(new_n986_), .Y(new_n12026_));
  NOR2  g11641(.A(new_n12026_), .B(new_n991_), .Y(new_n12027_));
  NOR2  g11642(.A(new_n12027_), .B(new_n995_), .Y(new_n12028_));
  NOR2  g11643(.A(new_n12028_), .B(new_n1000_), .Y(new_n12029_));
  NOR2  g11644(.A(new_n12029_), .B(new_n1004_), .Y(new_n12030_));
  NOR2  g11645(.A(new_n12030_), .B(new_n1009_), .Y(new_n12031_));
  NOR2  g11646(.A(new_n12031_), .B(new_n1013_), .Y(new_n12032_));
  NOR2  g11647(.A(new_n12032_), .B(new_n1018_), .Y(new_n12033_));
  NOR2  g11648(.A(new_n12033_), .B(new_n1022_), .Y(new_n12034_));
  NOR2  g11649(.A(new_n12034_), .B(new_n1027_), .Y(new_n12035_));
  NOR2  g11650(.A(new_n12035_), .B(new_n1031_), .Y(new_n12036_));
  NOR2  g11651(.A(new_n12036_), .B(new_n1036_), .Y(new_n12037_));
  NOR2  g11652(.A(new_n12037_), .B(new_n1040_), .Y(new_n12038_));
  NOR2  g11653(.A(new_n12038_), .B(new_n1045_), .Y(new_n12039_));
  NOR2  g11654(.A(new_n12039_), .B(new_n1049_), .Y(new_n12040_));
  NOR2  g11655(.A(new_n12040_), .B(new_n1054_), .Y(new_n12041_));
  NOR2  g11656(.A(new_n12041_), .B(new_n1058_), .Y(new_n12042_));
  NOR2  g11657(.A(new_n12042_), .B(new_n1063_), .Y(new_n12043_));
  NOR2  g11658(.A(new_n12043_), .B(new_n1067_), .Y(new_n12044_));
  NOR2  g11659(.A(new_n12044_), .B(new_n1072_), .Y(new_n12045_));
  NOR2  g11660(.A(new_n12045_), .B(new_n1076_), .Y(new_n12046_));
  NOR2  g11661(.A(new_n12046_), .B(new_n1081_), .Y(new_n12047_));
  NOR2  g11662(.A(new_n12047_), .B(new_n1085_), .Y(new_n12048_));
  NOR2  g11663(.A(new_n12048_), .B(new_n1090_), .Y(new_n12049_));
  NOR2  g11664(.A(new_n12049_), .B(new_n1094_), .Y(new_n12050_));
  NOR2  g11665(.A(new_n12050_), .B(new_n1099_), .Y(new_n12051_));
  NOR2  g11666(.A(new_n12051_), .B(new_n1103_), .Y(new_n12052_));
  NOR2  g11667(.A(new_n12052_), .B(new_n1108_), .Y(new_n12053_));
  NOR2  g11668(.A(new_n12053_), .B(new_n1112_), .Y(new_n12054_));
  NOR2  g11669(.A(new_n12054_), .B(new_n1117_), .Y(new_n12055_));
  NOR2  g11670(.A(new_n12055_), .B(new_n1121_), .Y(new_n12056_));
  NOR2  g11671(.A(new_n12056_), .B(new_n1126_), .Y(new_n12057_));
  NOR2  g11672(.A(new_n12057_), .B(new_n1130_), .Y(new_n12058_));
  NOR2  g11673(.A(new_n12058_), .B(new_n1135_), .Y(new_n12059_));
  NOR2  g11674(.A(new_n12059_), .B(new_n1139_), .Y(new_n12060_));
  NOR2  g11675(.A(new_n12060_), .B(new_n1144_), .Y(new_n12061_));
  NOR2  g11676(.A(new_n12061_), .B(new_n1148_), .Y(new_n12062_));
  NOR2  g11677(.A(new_n12062_), .B(new_n1153_), .Y(new_n12063_));
  NOR2  g11678(.A(new_n12063_), .B(new_n1157_), .Y(new_n12064_));
  NOR2  g11679(.A(new_n12064_), .B(new_n1162_), .Y(new_n12065_));
  NOR2  g11680(.A(new_n12065_), .B(new_n1166_), .Y(new_n12066_));
  NOR2  g11681(.A(new_n12066_), .B(new_n1171_), .Y(new_n12067_));
  NAND2 g11682(.A(new_n1173_), .B(\req[123] ), .Y(new_n12068_));
  NOR2  g11683(.A(new_n12068_), .B(new_n12067_), .Y(\grant[123] ));
  INV   g11684(.A(new_n1183_), .Y(new_n12070_));
  NOR2  g11685(.A(new_n1518_), .B(new_n12070_), .Y(new_n12071_));
  NOR2  g11686(.A(new_n12071_), .B(new_n1189_), .Y(new_n12072_));
  NOR2  g11687(.A(new_n12072_), .B(new_n1707_), .Y(new_n12073_));
  NOR2  g11688(.A(new_n12073_), .B(new_n1709_), .Y(new_n12074_));
  NOR2  g11689(.A(new_n12074_), .B(new_n1973_), .Y(new_n12075_));
  NOR2  g11690(.A(new_n12075_), .B(new_n1199_), .Y(new_n12076_));
  NOR2  g11691(.A(new_n12076_), .B(new_n1203_), .Y(new_n12077_));
  NOR2  g11692(.A(new_n12077_), .B(new_n1207_), .Y(new_n12078_));
  NOR2  g11693(.A(new_n12078_), .B(new_n1211_), .Y(new_n12079_));
  NOR2  g11694(.A(new_n12079_), .B(new_n1215_), .Y(new_n12080_));
  NOR2  g11695(.A(new_n12080_), .B(new_n1219_), .Y(new_n12081_));
  NOR2  g11696(.A(new_n12081_), .B(new_n1223_), .Y(new_n12082_));
  NOR2  g11697(.A(new_n12082_), .B(new_n1227_), .Y(new_n12083_));
  NOR2  g11698(.A(new_n12083_), .B(new_n1231_), .Y(new_n12084_));
  NOR2  g11699(.A(new_n12084_), .B(new_n1235_), .Y(new_n12085_));
  NOR2  g11700(.A(new_n12085_), .B(new_n1239_), .Y(new_n12086_));
  NOR2  g11701(.A(new_n12086_), .B(new_n1243_), .Y(new_n12087_));
  NOR2  g11702(.A(new_n12087_), .B(new_n1247_), .Y(new_n12088_));
  NOR2  g11703(.A(new_n12088_), .B(new_n1251_), .Y(new_n12089_));
  NOR2  g11704(.A(new_n12089_), .B(new_n1255_), .Y(new_n12090_));
  NOR2  g11705(.A(new_n12090_), .B(new_n1259_), .Y(new_n12091_));
  NOR2  g11706(.A(new_n12091_), .B(new_n1263_), .Y(new_n12092_));
  NOR2  g11707(.A(new_n12092_), .B(new_n1267_), .Y(new_n12093_));
  NOR2  g11708(.A(new_n12093_), .B(new_n1271_), .Y(new_n12094_));
  NOR2  g11709(.A(new_n12094_), .B(new_n1275_), .Y(new_n12095_));
  NOR2  g11710(.A(new_n12095_), .B(new_n1279_), .Y(new_n12096_));
  NOR2  g11711(.A(new_n12096_), .B(new_n1283_), .Y(new_n12097_));
  NOR2  g11712(.A(new_n12097_), .B(new_n1287_), .Y(new_n12098_));
  NOR2  g11713(.A(new_n12098_), .B(new_n1291_), .Y(new_n12099_));
  NOR2  g11714(.A(new_n12099_), .B(new_n1295_), .Y(new_n12100_));
  NOR2  g11715(.A(new_n12100_), .B(new_n1299_), .Y(new_n12101_));
  NOR2  g11716(.A(new_n12101_), .B(new_n1303_), .Y(new_n12102_));
  NOR2  g11717(.A(new_n12102_), .B(new_n1307_), .Y(new_n12103_));
  NOR2  g11718(.A(new_n12103_), .B(new_n1311_), .Y(new_n12104_));
  NOR2  g11719(.A(new_n12104_), .B(new_n1315_), .Y(new_n12105_));
  NOR2  g11720(.A(new_n12105_), .B(new_n1319_), .Y(new_n12106_));
  NOR2  g11721(.A(new_n12106_), .B(new_n1323_), .Y(new_n12107_));
  NOR2  g11722(.A(new_n12107_), .B(new_n1327_), .Y(new_n12108_));
  NOR2  g11723(.A(new_n12108_), .B(new_n1331_), .Y(new_n12109_));
  NOR2  g11724(.A(new_n12109_), .B(new_n1335_), .Y(new_n12110_));
  NOR2  g11725(.A(new_n12110_), .B(new_n1339_), .Y(new_n12111_));
  NOR2  g11726(.A(new_n12111_), .B(new_n1343_), .Y(new_n12112_));
  NOR2  g11727(.A(new_n12112_), .B(new_n1347_), .Y(new_n12113_));
  NOR2  g11728(.A(new_n12113_), .B(new_n1351_), .Y(new_n12114_));
  NOR2  g11729(.A(new_n12114_), .B(new_n1355_), .Y(new_n12115_));
  NOR2  g11730(.A(new_n12115_), .B(new_n1359_), .Y(new_n12116_));
  NOR2  g11731(.A(new_n12116_), .B(new_n1363_), .Y(new_n12117_));
  NOR2  g11732(.A(new_n12117_), .B(new_n1367_), .Y(new_n12118_));
  NOR2  g11733(.A(new_n12118_), .B(new_n1371_), .Y(new_n12119_));
  NOR2  g11734(.A(new_n12119_), .B(new_n1375_), .Y(new_n12120_));
  NOR2  g11735(.A(new_n12120_), .B(new_n1379_), .Y(new_n12121_));
  NOR2  g11736(.A(new_n12121_), .B(new_n1383_), .Y(new_n12122_));
  NOR2  g11737(.A(new_n12122_), .B(new_n1387_), .Y(new_n12123_));
  NOR2  g11738(.A(new_n12123_), .B(new_n1391_), .Y(new_n12124_));
  NOR2  g11739(.A(new_n12124_), .B(new_n1395_), .Y(new_n12125_));
  NOR2  g11740(.A(new_n12125_), .B(new_n1399_), .Y(new_n12126_));
  NOR2  g11741(.A(new_n12126_), .B(new_n1403_), .Y(new_n12127_));
  NOR2  g11742(.A(new_n12127_), .B(new_n1407_), .Y(new_n12128_));
  NOR2  g11743(.A(new_n12128_), .B(new_n1411_), .Y(new_n12129_));
  NOR2  g11744(.A(new_n12129_), .B(new_n1415_), .Y(new_n12130_));
  NOR2  g11745(.A(new_n12130_), .B(new_n1419_), .Y(new_n12131_));
  NOR2  g11746(.A(new_n12131_), .B(new_n1423_), .Y(new_n12132_));
  NOR2  g11747(.A(new_n12132_), .B(new_n1427_), .Y(new_n12133_));
  NOR2  g11748(.A(new_n12133_), .B(new_n1431_), .Y(new_n12134_));
  NOR2  g11749(.A(new_n12134_), .B(new_n1435_), .Y(new_n12135_));
  NOR2  g11750(.A(new_n12135_), .B(new_n1439_), .Y(new_n12136_));
  NOR2  g11751(.A(new_n12136_), .B(new_n1443_), .Y(new_n12137_));
  NOR2  g11752(.A(new_n12137_), .B(new_n1447_), .Y(new_n12138_));
  NOR2  g11753(.A(new_n12138_), .B(new_n1451_), .Y(new_n12139_));
  NOR2  g11754(.A(new_n12139_), .B(new_n1455_), .Y(new_n12140_));
  NOR2  g11755(.A(new_n12140_), .B(new_n1459_), .Y(new_n12141_));
  NOR2  g11756(.A(new_n12141_), .B(new_n1463_), .Y(new_n12142_));
  NOR2  g11757(.A(new_n12142_), .B(new_n1467_), .Y(new_n12143_));
  NOR2  g11758(.A(new_n12143_), .B(new_n1471_), .Y(new_n12144_));
  NOR2  g11759(.A(new_n12144_), .B(new_n1475_), .Y(new_n12145_));
  NOR2  g11760(.A(new_n12145_), .B(new_n1479_), .Y(new_n12146_));
  NOR2  g11761(.A(new_n12146_), .B(new_n1483_), .Y(new_n12147_));
  NOR2  g11762(.A(new_n12147_), .B(new_n1487_), .Y(new_n12148_));
  NOR2  g11763(.A(new_n12148_), .B(new_n1491_), .Y(new_n12149_));
  NOR2  g11764(.A(new_n12149_), .B(new_n1495_), .Y(new_n12150_));
  NOR2  g11765(.A(new_n12150_), .B(new_n1499_), .Y(new_n12151_));
  NOR2  g11766(.A(new_n12151_), .B(new_n1503_), .Y(new_n12152_));
  NOR2  g11767(.A(new_n12152_), .B(new_n1507_), .Y(new_n12153_));
  NOR2  g11768(.A(new_n12153_), .B(new_n1511_), .Y(new_n12154_));
  NAND2 g11769(.A(new_n1513_), .B(\req[124] ), .Y(new_n12155_));
  NOR2  g11770(.A(new_n12155_), .B(new_n12154_), .Y(\grant[124] ));
  INV   g11771(.A(new_n1522_), .Y(new_n12157_));
  NOR2  g11772(.A(new_n12157_), .B(new_n805_), .Y(new_n12158_));
  NOR2  g11773(.A(new_n12158_), .B(new_n1527_), .Y(new_n12159_));
  NOR2  g11774(.A(new_n12159_), .B(new_n1797_), .Y(new_n12160_));
  NOR2  g11775(.A(new_n12160_), .B(new_n396_), .Y(new_n12161_));
  NOR2  g11776(.A(new_n12161_), .B(new_n400_), .Y(new_n12162_));
  NOR2  g11777(.A(new_n12162_), .B(new_n406_), .Y(new_n12163_));
  NOR2  g11778(.A(new_n12163_), .B(new_n410_), .Y(new_n12164_));
  NOR2  g11779(.A(new_n12164_), .B(new_n416_), .Y(new_n12165_));
  NOR2  g11780(.A(new_n12165_), .B(new_n420_), .Y(new_n12166_));
  NOR2  g11781(.A(new_n12166_), .B(new_n426_), .Y(new_n12167_));
  NOR2  g11782(.A(new_n12167_), .B(new_n430_), .Y(new_n12168_));
  NOR2  g11783(.A(new_n12168_), .B(new_n436_), .Y(new_n12169_));
  NOR2  g11784(.A(new_n12169_), .B(new_n440_), .Y(new_n12170_));
  NOR2  g11785(.A(new_n12170_), .B(new_n446_), .Y(new_n12171_));
  NOR2  g11786(.A(new_n12171_), .B(new_n450_), .Y(new_n12172_));
  NOR2  g11787(.A(new_n12172_), .B(new_n456_), .Y(new_n12173_));
  NOR2  g11788(.A(new_n12173_), .B(new_n460_), .Y(new_n12174_));
  NOR2  g11789(.A(new_n12174_), .B(new_n466_), .Y(new_n12175_));
  NOR2  g11790(.A(new_n12175_), .B(new_n470_), .Y(new_n12176_));
  NOR2  g11791(.A(new_n12176_), .B(new_n476_), .Y(new_n12177_));
  NOR2  g11792(.A(new_n12177_), .B(new_n480_), .Y(new_n12178_));
  NOR2  g11793(.A(new_n12178_), .B(new_n486_), .Y(new_n12179_));
  NOR2  g11794(.A(new_n12179_), .B(new_n490_), .Y(new_n12180_));
  NOR2  g11795(.A(new_n12180_), .B(new_n496_), .Y(new_n12181_));
  NOR2  g11796(.A(new_n12181_), .B(new_n500_), .Y(new_n12182_));
  NOR2  g11797(.A(new_n12182_), .B(new_n506_), .Y(new_n12183_));
  NOR2  g11798(.A(new_n12183_), .B(new_n510_), .Y(new_n12184_));
  NOR2  g11799(.A(new_n12184_), .B(new_n516_), .Y(new_n12185_));
  NOR2  g11800(.A(new_n12185_), .B(new_n520_), .Y(new_n12186_));
  NOR2  g11801(.A(new_n12186_), .B(new_n526_), .Y(new_n12187_));
  NOR2  g11802(.A(new_n12187_), .B(new_n530_), .Y(new_n12188_));
  NOR2  g11803(.A(new_n12188_), .B(new_n536_), .Y(new_n12189_));
  NOR2  g11804(.A(new_n12189_), .B(new_n540_), .Y(new_n12190_));
  NOR2  g11805(.A(new_n12190_), .B(new_n546_), .Y(new_n12191_));
  NOR2  g11806(.A(new_n12191_), .B(new_n550_), .Y(new_n12192_));
  NOR2  g11807(.A(new_n12192_), .B(new_n556_), .Y(new_n12193_));
  NOR2  g11808(.A(new_n12193_), .B(new_n560_), .Y(new_n12194_));
  NOR2  g11809(.A(new_n12194_), .B(new_n566_), .Y(new_n12195_));
  NOR2  g11810(.A(new_n12195_), .B(new_n570_), .Y(new_n12196_));
  NOR2  g11811(.A(new_n12196_), .B(new_n576_), .Y(new_n12197_));
  NOR2  g11812(.A(new_n12197_), .B(new_n580_), .Y(new_n12198_));
  NOR2  g11813(.A(new_n12198_), .B(new_n586_), .Y(new_n12199_));
  NOR2  g11814(.A(new_n12199_), .B(new_n590_), .Y(new_n12200_));
  NOR2  g11815(.A(new_n12200_), .B(new_n596_), .Y(new_n12201_));
  NOR2  g11816(.A(new_n12201_), .B(new_n600_), .Y(new_n12202_));
  NOR2  g11817(.A(new_n12202_), .B(new_n606_), .Y(new_n12203_));
  NOR2  g11818(.A(new_n12203_), .B(new_n610_), .Y(new_n12204_));
  NOR2  g11819(.A(new_n12204_), .B(new_n616_), .Y(new_n12205_));
  NOR2  g11820(.A(new_n12205_), .B(new_n620_), .Y(new_n12206_));
  NOR2  g11821(.A(new_n12206_), .B(new_n626_), .Y(new_n12207_));
  NOR2  g11822(.A(new_n12207_), .B(new_n630_), .Y(new_n12208_));
  NOR2  g11823(.A(new_n12208_), .B(new_n636_), .Y(new_n12209_));
  NOR2  g11824(.A(new_n12209_), .B(new_n640_), .Y(new_n12210_));
  NOR2  g11825(.A(new_n12210_), .B(new_n646_), .Y(new_n12211_));
  NOR2  g11826(.A(new_n12211_), .B(new_n650_), .Y(new_n12212_));
  NOR2  g11827(.A(new_n12212_), .B(new_n656_), .Y(new_n12213_));
  NOR2  g11828(.A(new_n12213_), .B(new_n660_), .Y(new_n12214_));
  NOR2  g11829(.A(new_n12214_), .B(new_n666_), .Y(new_n12215_));
  NOR2  g11830(.A(new_n12215_), .B(new_n670_), .Y(new_n12216_));
  NOR2  g11831(.A(new_n12216_), .B(new_n676_), .Y(new_n12217_));
  NOR2  g11832(.A(new_n12217_), .B(new_n680_), .Y(new_n12218_));
  NOR2  g11833(.A(new_n12218_), .B(new_n686_), .Y(new_n12219_));
  NOR2  g11834(.A(new_n12219_), .B(new_n690_), .Y(new_n12220_));
  NOR2  g11835(.A(new_n12220_), .B(new_n696_), .Y(new_n12221_));
  NOR2  g11836(.A(new_n12221_), .B(new_n700_), .Y(new_n12222_));
  NOR2  g11837(.A(new_n12222_), .B(new_n706_), .Y(new_n12223_));
  NOR2  g11838(.A(new_n12223_), .B(new_n710_), .Y(new_n12224_));
  NOR2  g11839(.A(new_n12224_), .B(new_n716_), .Y(new_n12225_));
  NOR2  g11840(.A(new_n12225_), .B(new_n720_), .Y(new_n12226_));
  NOR2  g11841(.A(new_n12226_), .B(new_n726_), .Y(new_n12227_));
  NOR2  g11842(.A(new_n12227_), .B(new_n730_), .Y(new_n12228_));
  NOR2  g11843(.A(new_n12228_), .B(new_n736_), .Y(new_n12229_));
  NOR2  g11844(.A(new_n12229_), .B(new_n740_), .Y(new_n12230_));
  NOR2  g11845(.A(new_n12230_), .B(new_n746_), .Y(new_n12231_));
  NOR2  g11846(.A(new_n12231_), .B(new_n750_), .Y(new_n12232_));
  NOR2  g11847(.A(new_n12232_), .B(new_n756_), .Y(new_n12233_));
  NOR2  g11848(.A(new_n12233_), .B(new_n760_), .Y(new_n12234_));
  NOR2  g11849(.A(new_n12234_), .B(new_n766_), .Y(new_n12235_));
  NOR2  g11850(.A(new_n12235_), .B(new_n770_), .Y(new_n12236_));
  NOR2  g11851(.A(new_n12236_), .B(new_n776_), .Y(new_n12237_));
  NOR2  g11852(.A(new_n12237_), .B(new_n780_), .Y(new_n12238_));
  NOR2  g11853(.A(new_n12238_), .B(new_n786_), .Y(new_n12239_));
  NOR2  g11854(.A(new_n12239_), .B(new_n790_), .Y(new_n12240_));
  NOR2  g11855(.A(new_n12240_), .B(new_n796_), .Y(new_n12241_));
  NAND2 g11856(.A(new_n798_), .B(\req[125] ), .Y(new_n12242_));
  NOR2  g11857(.A(new_n12242_), .B(new_n12241_), .Y(\grant[125] ));
  INV   g11858(.A(new_n1615_), .Y(new_n12244_));
  NOR2  g11859(.A(new_n12244_), .B(new_n1188_), .Y(new_n12245_));
  NOR2  g11860(.A(new_n12245_), .B(new_n1618_), .Y(new_n12246_));
  NOR2  g11861(.A(new_n12246_), .B(new_n1885_), .Y(new_n12247_));
  NOR2  g11862(.A(new_n12247_), .B(new_n820_), .Y(new_n12248_));
  NOR2  g11863(.A(new_n12248_), .B(new_n824_), .Y(new_n12249_));
  NOR2  g11864(.A(new_n12249_), .B(new_n829_), .Y(new_n12250_));
  NOR2  g11865(.A(new_n12250_), .B(new_n833_), .Y(new_n12251_));
  NOR2  g11866(.A(new_n12251_), .B(new_n838_), .Y(new_n12252_));
  NOR2  g11867(.A(new_n12252_), .B(new_n842_), .Y(new_n12253_));
  NOR2  g11868(.A(new_n12253_), .B(new_n847_), .Y(new_n12254_));
  NOR2  g11869(.A(new_n12254_), .B(new_n851_), .Y(new_n12255_));
  NOR2  g11870(.A(new_n12255_), .B(new_n856_), .Y(new_n12256_));
  NOR2  g11871(.A(new_n12256_), .B(new_n860_), .Y(new_n12257_));
  NOR2  g11872(.A(new_n12257_), .B(new_n865_), .Y(new_n12258_));
  NOR2  g11873(.A(new_n12258_), .B(new_n869_), .Y(new_n12259_));
  NOR2  g11874(.A(new_n12259_), .B(new_n874_), .Y(new_n12260_));
  NOR2  g11875(.A(new_n12260_), .B(new_n878_), .Y(new_n12261_));
  NOR2  g11876(.A(new_n12261_), .B(new_n883_), .Y(new_n12262_));
  NOR2  g11877(.A(new_n12262_), .B(new_n887_), .Y(new_n12263_));
  NOR2  g11878(.A(new_n12263_), .B(new_n892_), .Y(new_n12264_));
  NOR2  g11879(.A(new_n12264_), .B(new_n896_), .Y(new_n12265_));
  NOR2  g11880(.A(new_n12265_), .B(new_n901_), .Y(new_n12266_));
  NOR2  g11881(.A(new_n12266_), .B(new_n905_), .Y(new_n12267_));
  NOR2  g11882(.A(new_n12267_), .B(new_n910_), .Y(new_n12268_));
  NOR2  g11883(.A(new_n12268_), .B(new_n914_), .Y(new_n12269_));
  NOR2  g11884(.A(new_n12269_), .B(new_n919_), .Y(new_n12270_));
  NOR2  g11885(.A(new_n12270_), .B(new_n923_), .Y(new_n12271_));
  NOR2  g11886(.A(new_n12271_), .B(new_n928_), .Y(new_n12272_));
  NOR2  g11887(.A(new_n12272_), .B(new_n932_), .Y(new_n12273_));
  NOR2  g11888(.A(new_n12273_), .B(new_n937_), .Y(new_n12274_));
  NOR2  g11889(.A(new_n12274_), .B(new_n941_), .Y(new_n12275_));
  NOR2  g11890(.A(new_n12275_), .B(new_n946_), .Y(new_n12276_));
  NOR2  g11891(.A(new_n12276_), .B(new_n950_), .Y(new_n12277_));
  NOR2  g11892(.A(new_n12277_), .B(new_n955_), .Y(new_n12278_));
  NOR2  g11893(.A(new_n12278_), .B(new_n959_), .Y(new_n12279_));
  NOR2  g11894(.A(new_n12279_), .B(new_n964_), .Y(new_n12280_));
  NOR2  g11895(.A(new_n12280_), .B(new_n968_), .Y(new_n12281_));
  NOR2  g11896(.A(new_n12281_), .B(new_n973_), .Y(new_n12282_));
  NOR2  g11897(.A(new_n12282_), .B(new_n977_), .Y(new_n12283_));
  NOR2  g11898(.A(new_n12283_), .B(new_n982_), .Y(new_n12284_));
  NOR2  g11899(.A(new_n12284_), .B(new_n986_), .Y(new_n12285_));
  NOR2  g11900(.A(new_n12285_), .B(new_n991_), .Y(new_n12286_));
  NOR2  g11901(.A(new_n12286_), .B(new_n995_), .Y(new_n12287_));
  NOR2  g11902(.A(new_n12287_), .B(new_n1000_), .Y(new_n12288_));
  NOR2  g11903(.A(new_n12288_), .B(new_n1004_), .Y(new_n12289_));
  NOR2  g11904(.A(new_n12289_), .B(new_n1009_), .Y(new_n12290_));
  NOR2  g11905(.A(new_n12290_), .B(new_n1013_), .Y(new_n12291_));
  NOR2  g11906(.A(new_n12291_), .B(new_n1018_), .Y(new_n12292_));
  NOR2  g11907(.A(new_n12292_), .B(new_n1022_), .Y(new_n12293_));
  NOR2  g11908(.A(new_n12293_), .B(new_n1027_), .Y(new_n12294_));
  NOR2  g11909(.A(new_n12294_), .B(new_n1031_), .Y(new_n12295_));
  NOR2  g11910(.A(new_n12295_), .B(new_n1036_), .Y(new_n12296_));
  NOR2  g11911(.A(new_n12296_), .B(new_n1040_), .Y(new_n12297_));
  NOR2  g11912(.A(new_n12297_), .B(new_n1045_), .Y(new_n12298_));
  NOR2  g11913(.A(new_n12298_), .B(new_n1049_), .Y(new_n12299_));
  NOR2  g11914(.A(new_n12299_), .B(new_n1054_), .Y(new_n12300_));
  NOR2  g11915(.A(new_n12300_), .B(new_n1058_), .Y(new_n12301_));
  NOR2  g11916(.A(new_n12301_), .B(new_n1063_), .Y(new_n12302_));
  NOR2  g11917(.A(new_n12302_), .B(new_n1067_), .Y(new_n12303_));
  NOR2  g11918(.A(new_n12303_), .B(new_n1072_), .Y(new_n12304_));
  NOR2  g11919(.A(new_n12304_), .B(new_n1076_), .Y(new_n12305_));
  NOR2  g11920(.A(new_n12305_), .B(new_n1081_), .Y(new_n12306_));
  NOR2  g11921(.A(new_n12306_), .B(new_n1085_), .Y(new_n12307_));
  NOR2  g11922(.A(new_n12307_), .B(new_n1090_), .Y(new_n12308_));
  NOR2  g11923(.A(new_n12308_), .B(new_n1094_), .Y(new_n12309_));
  NOR2  g11924(.A(new_n12309_), .B(new_n1099_), .Y(new_n12310_));
  NOR2  g11925(.A(new_n12310_), .B(new_n1103_), .Y(new_n12311_));
  NOR2  g11926(.A(new_n12311_), .B(new_n1108_), .Y(new_n12312_));
  NOR2  g11927(.A(new_n12312_), .B(new_n1112_), .Y(new_n12313_));
  NOR2  g11928(.A(new_n12313_), .B(new_n1117_), .Y(new_n12314_));
  NOR2  g11929(.A(new_n12314_), .B(new_n1121_), .Y(new_n12315_));
  NOR2  g11930(.A(new_n12315_), .B(new_n1126_), .Y(new_n12316_));
  NOR2  g11931(.A(new_n12316_), .B(new_n1130_), .Y(new_n12317_));
  NOR2  g11932(.A(new_n12317_), .B(new_n1135_), .Y(new_n12318_));
  NOR2  g11933(.A(new_n12318_), .B(new_n1139_), .Y(new_n12319_));
  NOR2  g11934(.A(new_n12319_), .B(new_n1144_), .Y(new_n12320_));
  NOR2  g11935(.A(new_n12320_), .B(new_n1148_), .Y(new_n12321_));
  NOR2  g11936(.A(new_n12321_), .B(new_n1153_), .Y(new_n12322_));
  NOR2  g11937(.A(new_n12322_), .B(new_n1157_), .Y(new_n12323_));
  NOR2  g11938(.A(new_n12323_), .B(new_n1162_), .Y(new_n12324_));
  NOR2  g11939(.A(new_n12324_), .B(new_n1166_), .Y(new_n12325_));
  NOR2  g11940(.A(new_n12325_), .B(new_n1171_), .Y(new_n12326_));
  NOR2  g11941(.A(new_n12326_), .B(new_n1175_), .Y(new_n12327_));
  NOR2  g11942(.A(new_n12327_), .B(new_n1180_), .Y(new_n12328_));
  NAND2 g11943(.A(new_n1182_), .B(\req[126] ), .Y(new_n12329_));
  NOR2  g11944(.A(new_n12329_), .B(new_n12328_), .Y(\grant[126] ));
  INV   g11945(.A(new_n1706_), .Y(new_n12331_));
  NOR2  g11946(.A(new_n12331_), .B(new_n1526_), .Y(new_n12332_));
  NOR2  g11947(.A(new_n12332_), .B(new_n1709_), .Y(new_n12333_));
  NOR2  g11948(.A(new_n12333_), .B(new_n1973_), .Y(new_n12334_));
  NOR2  g11949(.A(new_n12334_), .B(new_n1199_), .Y(new_n12335_));
  NOR2  g11950(.A(new_n12335_), .B(new_n1203_), .Y(new_n12336_));
  NOR2  g11951(.A(new_n12336_), .B(new_n1207_), .Y(new_n12337_));
  NOR2  g11952(.A(new_n12337_), .B(new_n1211_), .Y(new_n12338_));
  NOR2  g11953(.A(new_n12338_), .B(new_n1215_), .Y(new_n12339_));
  NOR2  g11954(.A(new_n12339_), .B(new_n1219_), .Y(new_n12340_));
  NOR2  g11955(.A(new_n12340_), .B(new_n1223_), .Y(new_n12341_));
  NOR2  g11956(.A(new_n12341_), .B(new_n1227_), .Y(new_n12342_));
  NOR2  g11957(.A(new_n12342_), .B(new_n1231_), .Y(new_n12343_));
  NOR2  g11958(.A(new_n12343_), .B(new_n1235_), .Y(new_n12344_));
  NOR2  g11959(.A(new_n12344_), .B(new_n1239_), .Y(new_n12345_));
  NOR2  g11960(.A(new_n12345_), .B(new_n1243_), .Y(new_n12346_));
  NOR2  g11961(.A(new_n12346_), .B(new_n1247_), .Y(new_n12347_));
  NOR2  g11962(.A(new_n12347_), .B(new_n1251_), .Y(new_n12348_));
  NOR2  g11963(.A(new_n12348_), .B(new_n1255_), .Y(new_n12349_));
  NOR2  g11964(.A(new_n12349_), .B(new_n1259_), .Y(new_n12350_));
  NOR2  g11965(.A(new_n12350_), .B(new_n1263_), .Y(new_n12351_));
  NOR2  g11966(.A(new_n12351_), .B(new_n1267_), .Y(new_n12352_));
  NOR2  g11967(.A(new_n12352_), .B(new_n1271_), .Y(new_n12353_));
  NOR2  g11968(.A(new_n12353_), .B(new_n1275_), .Y(new_n12354_));
  NOR2  g11969(.A(new_n12354_), .B(new_n1279_), .Y(new_n12355_));
  NOR2  g11970(.A(new_n12355_), .B(new_n1283_), .Y(new_n12356_));
  NOR2  g11971(.A(new_n12356_), .B(new_n1287_), .Y(new_n12357_));
  NOR2  g11972(.A(new_n12357_), .B(new_n1291_), .Y(new_n12358_));
  NOR2  g11973(.A(new_n12358_), .B(new_n1295_), .Y(new_n12359_));
  NOR2  g11974(.A(new_n12359_), .B(new_n1299_), .Y(new_n12360_));
  NOR2  g11975(.A(new_n12360_), .B(new_n1303_), .Y(new_n12361_));
  NOR2  g11976(.A(new_n12361_), .B(new_n1307_), .Y(new_n12362_));
  NOR2  g11977(.A(new_n12362_), .B(new_n1311_), .Y(new_n12363_));
  NOR2  g11978(.A(new_n12363_), .B(new_n1315_), .Y(new_n12364_));
  NOR2  g11979(.A(new_n12364_), .B(new_n1319_), .Y(new_n12365_));
  NOR2  g11980(.A(new_n12365_), .B(new_n1323_), .Y(new_n12366_));
  NOR2  g11981(.A(new_n12366_), .B(new_n1327_), .Y(new_n12367_));
  NOR2  g11982(.A(new_n12367_), .B(new_n1331_), .Y(new_n12368_));
  NOR2  g11983(.A(new_n12368_), .B(new_n1335_), .Y(new_n12369_));
  NOR2  g11984(.A(new_n12369_), .B(new_n1339_), .Y(new_n12370_));
  NOR2  g11985(.A(new_n12370_), .B(new_n1343_), .Y(new_n12371_));
  NOR2  g11986(.A(new_n12371_), .B(new_n1347_), .Y(new_n12372_));
  NOR2  g11987(.A(new_n12372_), .B(new_n1351_), .Y(new_n12373_));
  NOR2  g11988(.A(new_n12373_), .B(new_n1355_), .Y(new_n12374_));
  NOR2  g11989(.A(new_n12374_), .B(new_n1359_), .Y(new_n12375_));
  NOR2  g11990(.A(new_n12375_), .B(new_n1363_), .Y(new_n12376_));
  NOR2  g11991(.A(new_n12376_), .B(new_n1367_), .Y(new_n12377_));
  NOR2  g11992(.A(new_n12377_), .B(new_n1371_), .Y(new_n12378_));
  NOR2  g11993(.A(new_n12378_), .B(new_n1375_), .Y(new_n12379_));
  NOR2  g11994(.A(new_n12379_), .B(new_n1379_), .Y(new_n12380_));
  NOR2  g11995(.A(new_n12380_), .B(new_n1383_), .Y(new_n12381_));
  NOR2  g11996(.A(new_n12381_), .B(new_n1387_), .Y(new_n12382_));
  NOR2  g11997(.A(new_n12382_), .B(new_n1391_), .Y(new_n12383_));
  NOR2  g11998(.A(new_n12383_), .B(new_n1395_), .Y(new_n12384_));
  NOR2  g11999(.A(new_n12384_), .B(new_n1399_), .Y(new_n12385_));
  NOR2  g12000(.A(new_n12385_), .B(new_n1403_), .Y(new_n12386_));
  NOR2  g12001(.A(new_n12386_), .B(new_n1407_), .Y(new_n12387_));
  NOR2  g12002(.A(new_n12387_), .B(new_n1411_), .Y(new_n12388_));
  NOR2  g12003(.A(new_n12388_), .B(new_n1415_), .Y(new_n12389_));
  NOR2  g12004(.A(new_n12389_), .B(new_n1419_), .Y(new_n12390_));
  NOR2  g12005(.A(new_n12390_), .B(new_n1423_), .Y(new_n12391_));
  NOR2  g12006(.A(new_n12391_), .B(new_n1427_), .Y(new_n12392_));
  NOR2  g12007(.A(new_n12392_), .B(new_n1431_), .Y(new_n12393_));
  NOR2  g12008(.A(new_n12393_), .B(new_n1435_), .Y(new_n12394_));
  NOR2  g12009(.A(new_n12394_), .B(new_n1439_), .Y(new_n12395_));
  NOR2  g12010(.A(new_n12395_), .B(new_n1443_), .Y(new_n12396_));
  NOR2  g12011(.A(new_n12396_), .B(new_n1447_), .Y(new_n12397_));
  NOR2  g12012(.A(new_n12397_), .B(new_n1451_), .Y(new_n12398_));
  NOR2  g12013(.A(new_n12398_), .B(new_n1455_), .Y(new_n12399_));
  NOR2  g12014(.A(new_n12399_), .B(new_n1459_), .Y(new_n12400_));
  NOR2  g12015(.A(new_n12400_), .B(new_n1463_), .Y(new_n12401_));
  NOR2  g12016(.A(new_n12401_), .B(new_n1467_), .Y(new_n12402_));
  NOR2  g12017(.A(new_n12402_), .B(new_n1471_), .Y(new_n12403_));
  NOR2  g12018(.A(new_n12403_), .B(new_n1475_), .Y(new_n12404_));
  NOR2  g12019(.A(new_n12404_), .B(new_n1479_), .Y(new_n12405_));
  NOR2  g12020(.A(new_n12405_), .B(new_n1483_), .Y(new_n12406_));
  NOR2  g12021(.A(new_n12406_), .B(new_n1487_), .Y(new_n12407_));
  NOR2  g12022(.A(new_n12407_), .B(new_n1491_), .Y(new_n12408_));
  NOR2  g12023(.A(new_n12408_), .B(new_n1495_), .Y(new_n12409_));
  NOR2  g12024(.A(new_n12409_), .B(new_n1499_), .Y(new_n12410_));
  NOR2  g12025(.A(new_n12410_), .B(new_n1503_), .Y(new_n12411_));
  NOR2  g12026(.A(new_n12411_), .B(new_n1507_), .Y(new_n12412_));
  NOR2  g12027(.A(new_n12412_), .B(new_n1511_), .Y(new_n12413_));
  NOR2  g12028(.A(new_n12413_), .B(new_n1515_), .Y(new_n12414_));
  NOR2  g12029(.A(new_n12414_), .B(new_n1519_), .Y(new_n12415_));
  NAND2 g12030(.A(new_n1521_), .B(\req[127] ), .Y(new_n12416_));
  NOR2  g12031(.A(new_n12416_), .B(new_n12415_), .Y(\grant[127] ));
  NOR2  g12032(.A(new_n1623_), .B(new_n11722_), .Y(new_n12418_));
  NOR2  g12033(.A(new_n2674_), .B(new_n2152_), .Y(new_n12419_));
  NAND2 g12034(.A(new_n12419_), .B(new_n12418_), .Y(new_n12420_));
  NOR2  g12035(.A(new_n10156_), .B(new_n9634_), .Y(new_n12421_));
  NOR2  g12036(.A(new_n11200_), .B(new_n10678_), .Y(new_n12422_));
  NAND2 g12037(.A(new_n12422_), .B(new_n12421_), .Y(new_n12423_));
  NOR2  g12038(.A(new_n12423_), .B(new_n12420_), .Y(new_n12424_));
  NOR2  g12039(.A(new_n5806_), .B(new_n5284_), .Y(new_n12425_));
  NOR2  g12040(.A(new_n6850_), .B(new_n6328_), .Y(new_n12426_));
  NAND2 g12041(.A(new_n12426_), .B(new_n12425_), .Y(new_n12427_));
  NOR2  g12042(.A(new_n3718_), .B(new_n3196_), .Y(new_n12428_));
  NOR2  g12043(.A(new_n4762_), .B(new_n4240_), .Y(new_n12429_));
  NAND2 g12044(.A(new_n12429_), .B(new_n12428_), .Y(new_n12430_));
  NOR2  g12045(.A(new_n12430_), .B(new_n12427_), .Y(new_n12431_));
  NAND2 g12046(.A(new_n12431_), .B(new_n12424_), .Y(new_n12432_));
  NOR2  g12047(.A(new_n3892_), .B(new_n3370_), .Y(new_n12433_));
  NOR2  g12048(.A(new_n4936_), .B(new_n4414_), .Y(new_n12434_));
  NAND2 g12049(.A(new_n12434_), .B(new_n12433_), .Y(new_n12435_));
  NOR2  g12050(.A(new_n1802_), .B(new_n390_), .Y(new_n12436_));
  NOR2  g12051(.A(new_n2848_), .B(new_n2326_), .Y(new_n12437_));
  NAND2 g12052(.A(new_n12437_), .B(new_n12436_), .Y(new_n12438_));
  NOR2  g12053(.A(new_n12438_), .B(new_n12435_), .Y(new_n12439_));
  NOR2  g12054(.A(new_n8068_), .B(new_n7546_), .Y(new_n12440_));
  NOR2  g12055(.A(new_n9112_), .B(new_n8590_), .Y(new_n12441_));
  NAND2 g12056(.A(new_n12441_), .B(new_n12440_), .Y(new_n12442_));
  NOR2  g12057(.A(new_n5980_), .B(new_n5458_), .Y(new_n12443_));
  NOR2  g12058(.A(new_n7024_), .B(new_n6502_), .Y(new_n12444_));
  NAND2 g12059(.A(new_n12444_), .B(new_n12443_), .Y(new_n12445_));
  NOR2  g12060(.A(new_n12445_), .B(new_n12442_), .Y(new_n12446_));
  NAND2 g12061(.A(new_n12446_), .B(new_n12439_), .Y(new_n12447_));
  NOR2  g12062(.A(new_n12447_), .B(new_n12432_), .Y(new_n12448_));
  NOR2  g12063(.A(new_n7198_), .B(new_n6676_), .Y(new_n12449_));
  NOR2  g12064(.A(new_n8242_), .B(new_n7720_), .Y(new_n12450_));
  NAND2 g12065(.A(new_n12450_), .B(new_n12449_), .Y(new_n12451_));
  NOR2  g12066(.A(new_n5110_), .B(new_n4588_), .Y(new_n12452_));
  NOR2  g12067(.A(new_n6154_), .B(new_n5632_), .Y(new_n12453_));
  NAND2 g12068(.A(new_n12453_), .B(new_n12452_), .Y(new_n12454_));
  NOR2  g12069(.A(new_n12454_), .B(new_n12451_), .Y(new_n12455_));
  NOR2  g12070(.A(new_n11374_), .B(new_n10852_), .Y(new_n12456_));
  NOR2  g12071(.A(new_n12244_), .B(new_n11896_), .Y(new_n12457_));
  NAND2 g12072(.A(new_n12457_), .B(new_n12456_), .Y(new_n12458_));
  NOR2  g12073(.A(new_n9286_), .B(new_n8764_), .Y(new_n12459_));
  NOR2  g12074(.A(new_n10330_), .B(new_n9808_), .Y(new_n12460_));
  NAND2 g12075(.A(new_n12460_), .B(new_n12459_), .Y(new_n12461_));
  NOR2  g12076(.A(new_n12461_), .B(new_n12458_), .Y(new_n12462_));
  NAND2 g12077(.A(new_n12462_), .B(new_n12455_), .Y(new_n12463_));
  NOR2  g12078(.A(new_n9982_), .B(new_n9460_), .Y(new_n12464_));
  NOR2  g12079(.A(new_n11026_), .B(new_n10504_), .Y(new_n12465_));
  NAND2 g12080(.A(new_n12465_), .B(new_n12464_), .Y(new_n12466_));
  NOR2  g12081(.A(new_n7894_), .B(new_n7372_), .Y(new_n12467_));
  NOR2  g12082(.A(new_n8938_), .B(new_n8416_), .Y(new_n12468_));
  NAND2 g12083(.A(new_n12468_), .B(new_n12467_), .Y(new_n12469_));
  NOR2  g12084(.A(new_n12469_), .B(new_n12466_), .Y(new_n12470_));
  NOR2  g12085(.A(new_n3022_), .B(new_n2500_), .Y(new_n12471_));
  NOR2  g12086(.A(new_n4066_), .B(new_n3544_), .Y(new_n12472_));
  NAND2 g12087(.A(new_n12472_), .B(new_n12471_), .Y(new_n12473_));
  NOR2  g12088(.A(new_n12070_), .B(new_n11548_), .Y(new_n12474_));
  NOR2  g12089(.A(new_n1978_), .B(new_n1195_), .Y(new_n12475_));
  NAND2 g12090(.A(new_n12475_), .B(new_n12474_), .Y(new_n12476_));
  NOR2  g12091(.A(new_n12476_), .B(new_n12473_), .Y(new_n12477_));
  NAND2 g12092(.A(new_n12477_), .B(new_n12470_), .Y(new_n12478_));
  NOR2  g12093(.A(new_n12478_), .B(new_n12463_), .Y(new_n12479_));
  NAND2 g12094(.A(new_n12479_), .B(new_n12448_), .Y(anyGrant));
endmodule


