//Converted to Combinational (Partial output: n60) , Module name: s1488_n60 , Timestamp: 2018-12-03T15:51:02.597894 
module s1488_n60 ( v1, CLR, v7, v10, v8, v11, v2, v9, v12, v3, v6, v0, v5, v4, n60 );
input CLR, v1, v7, v10, v8, v11, v2, v9, v12, v3, v6, v0, v5, v4;
output n60;
wire n267, n308, n315, n45, n299, n307, n311, n314, n72, n294, n298, n190, n302, n306, n103, n309, n310, n313, n204, n312, n82, n293, n297, n68, n295, n296, n135, n301, n305, n48, n304, n79, n63, n64, n57, n217, n109, n74, n203, n213, n110, n90, n259, n123, n300, n142, n251, n154, n58, n303, n104, n47;
AOI21X1  g271(.A0(n315), .A1(n308), .B0(n267), .Y(n60));
INVX1    g222(.A(CLR), .Y(n267));
OAI21X1  g263(.A0(n307), .A1(n299), .B0(n45), .Y(n308));
NOR2X1   g270(.A(n314), .B(n311), .Y(n315));
INVX1    g000(.A(v7), .Y(n45));
AOI21X1  g254(.A0(n298), .A1(n294), .B0(n72), .Y(n299));
NAND3X1  g262(.A(n306), .B(n302), .C(n190), .Y(n307));
AOI21X1  g266(.A0(n310), .A1(n309), .B0(n103), .Y(n311));
OAI22X1  g269(.A0(n312), .A1(n204), .B0(v10), .B1(n313), .Y(n314));
INVX1    g027(.A(v8), .Y(n72));
NAND3X1  g249(.A(n293), .B(n82), .C(n103), .Y(n294));
AOI22X1  g253(.A0(n296), .A1(n295), .B0(n68), .B1(n297), .Y(n298));
OR2X1    g145(.A(n135), .B(v11), .Y(n190));
NAND3X1  g257(.A(n301), .B(n72), .C(n82), .Y(n302));
AOI21X1  g261(.A0(n304), .A1(n48), .B0(n305), .Y(n306));
INVX1    g058(.A(v2), .Y(n103));
NAND4X1  g264(.A(n64), .B(n63), .C(v10), .D(n79), .Y(n309));
NAND3X1  g265(.A(n57), .B(n45), .C(v9), .Y(n310));
AOI22X1  g268(.A0(n74), .A1(n109), .B0(n217), .B1(v12), .Y(n313));
INVX1    g159(.A(n203), .Y(n204));
AOI22X1  g267(.A0(n110), .A1(v11), .B0(n217), .B1(n213), .Y(n312));
INVX1    g037(.A(v12), .Y(n82));
MX2X1    g248(.A(v10), .B(n90), .S0(v9), .Y(n293));
OAI21X1  g252(.A0(v9), .A1(v3), .B0(n109), .Y(n297));
INVX1    g023(.A(v10), .Y(n68));
NAND3X1  g250(.A(v0), .B(n259), .C(v6), .Y(n295));
AND2X1   g251(.A(n123), .B(v3), .Y(n296));
NAND2X1  g090(.A(v10), .B(v12), .Y(n135));
OAI21X1  g256(.A0(n142), .A1(v9), .B0(n300), .Y(n301));
NOR2X1   g260(.A(n251), .B(n63), .Y(n305));
INVX1    g003(.A(v6), .Y(n48));
OAI22X1  g259(.A0(n303), .A1(n58), .B0(v11), .B1(n154), .Y(n304));
AND2X1   g034(.A(v7), .B(v8), .Y(n79));
INVX1    g018(.A(v9), .Y(n63));
AND2X1   g019(.A(v11), .B(v12), .Y(n64));
NOR2X1   g012(.A(v10), .B(v12), .Y(n57));
NOR2X1   g172(.A(n72), .B(v11), .Y(n217));
NOR2X1   g064(.A(n104), .B(v12), .Y(n109));
NOR2X1   g029(.A(v8), .B(n63), .Y(n74));
NOR2X1   g158(.A(n45), .B(v12), .Y(n203));
NOR2X1   g168(.A(v9), .B(n68), .Y(n213));
NOR2X1   g065(.A(v8), .B(v10), .Y(n110));
AND2X1   g045(.A(v4), .B(v5), .Y(n90));
INVX1    g214(.A(v1), .Y(n259));
AND2X1   g078(.A(v9), .B(v12), .Y(n123));
NAND3X1  g255(.A(v9), .B(n68), .C(n259), .Y(n300));
NAND2X1  g097(.A(v10), .B(v11), .Y(n142));
MX2X1    g206(.A(v11), .B(n47), .S0(n68), .Y(n251));
NAND2X1  g109(.A(n63), .B(v12), .Y(n154));
INVX1    g013(.A(n57), .Y(n58));
NAND2X1  g258(.A(n72), .B(v9), .Y(n303));
INVX1    g059(.A(v11), .Y(n104));
NAND2X1  g002(.A(v11), .B(v12), .Y(n47));

endmodule
