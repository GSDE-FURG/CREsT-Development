//Converted to Combinational , Module name: s1494 , Timestamp: 2018-12-03T15:51:02.629875 
module s1494 ( CLR, v6, v5, v4, v3, v2, v1, v0, v12, v11, v10, v9, v8, v7, v13_D_24, v13_D_23, v13_D_22, v13_D_21, v13_D_20, v13_D_19, v13_D_18, v13_D_17, v13_D_16, v13_D_15, v13_D_14, v13_D_13, v13_D_12, v13_D_11, v13_D_10, v13_D_9, v13_D_8, v13_D_7, v13_D_6, n55, n60, n65, n70, n75, n80 );
input CLR, v6, v5, v4, v3, v2, v1, v0, v12, v11, v10, v9, v8, v7;
output v13_D_24, v13_D_23, v13_D_22, v13_D_21, v13_D_20, v13_D_19, v13_D_18, v13_D_17, v13_D_16, v13_D_15, v13_D_14, v13_D_13, v13_D_12, v13_D_11, v13_D_10, v13_D_9, v13_D_8, v13_D_7, v13_D_6, n55, n60, n65, n70, n75, n80;
wire n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55_1, n56, n57, n58, n59, n60_1, n61, n62, n63, n64, n65_1, n66, n67, n68, n69, n70_1, n71, n72, n73, n74, n75_1, n76, n77, n78, n79, n81, n82, n83, n84, n85, n86, n87, n88, n89, n91, n92, n93, n94, n95, n96, n97, n98, n100, n101, n102, n103, n104, n106, n107, n108, n109, n111, n112, n113, n114, n115, n116, n118, n119, n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n146, n147, n148, n150, n151, n152, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n196, n197, n198, n199, n200, n201, n202, n203, n204, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n220, n221, n222, n223, n224, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n244, n245, n246, n247, n248, n249, n250, n251, n252, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420;
INVX1    g000(.A(v10), .Y(n45));
NOR3X1   g001(.A(n45), .B(v11), .C(v12), .Y(n46));
AND2X1   g002(.A(v8), .B(v9), .Y(n47));
AND2X1   g003(.A(v3), .B(v6), .Y(n48));
AND2X1   g004(.A(n48), .B(n47), .Y(n49));
NAND2X1  g005(.A(v10), .B(v12), .Y(n50));
OR2X1    g006(.A(n50), .B(v11), .Y(n51));
INVX1    g007(.A(v5), .Y(n52));
AND2X1   g008(.A(v11), .B(v12), .Y(n53));
NOR2X1   g009(.A(v11), .B(v12), .Y(n54));
AOI21X1  g010(.A0(n54), .A1(n52), .B0(n53), .Y(n55_1));
OAI21X1  g011(.A0(n55_1), .A1(v10), .B0(n51), .Y(n56));
OR2X1    g012(.A(v8), .B(v9), .Y(n57));
INVX1    g013(.A(n57), .Y(n58));
AOI22X1  g014(.A0(n56), .A1(n58), .B0(n49), .B1(n46), .Y(n59));
NOR2X1   g015(.A(v7), .B(v8), .Y(n60_1));
NAND4X1  g016(.A(v10), .B(v11), .C(n52), .D(n60_1), .Y(n61));
INVX1    g017(.A(v2), .Y(n62));
NAND4X1  g018(.A(v8), .B(n45), .C(n62), .D(v7), .Y(n63));
OR2X1    g019(.A(v9), .B(v12), .Y(n64));
OR2X1    g020(.A(n64), .B(v0), .Y(n65_1));
AOI21X1  g021(.A0(n63), .A1(n61), .B0(n65_1), .Y(n66));
INVX1    g022(.A(v12), .Y(n67));
INVX1    g023(.A(v7), .Y(n68));
NOR4X1   g024(.A(v9), .B(n45), .C(n67), .D(n68), .Y(n69));
INVX1    g025(.A(v9), .Y(n70_1));
NOR2X1   g026(.A(n68), .B(v10), .Y(n71));
NOR4X1   g027(.A(n70_1), .B(v12), .C(v5), .D(n71), .Y(n72));
NOR2X1   g028(.A(n72), .B(n69), .Y(n73));
NAND2X1  g029(.A(v8), .B(n62), .Y(n74));
XOR2X1   g030(.A(n47), .B(v10), .Y(n75_1));
NOR2X1   g031(.A(n68), .B(v12), .Y(n76));
INVX1    g032(.A(n76), .Y(n77));
OAI22X1  g033(.A0(n75_1), .A1(n77), .B0(n74), .B1(n73), .Y(n78));
AOI21X1  g034(.A0(n78), .A1(v11), .B0(n66), .Y(n79));
OAI21X1  g035(.A0(n59), .A1(v7), .B0(n79), .Y(v13_D_24));
INVX1    g036(.A(n60_1), .Y(n81));
NAND4X1  g037(.A(v10), .B(v11), .C(v12), .D(v9), .Y(n82));
INVX1    g038(.A(v0), .Y(n83));
INVX1    g039(.A(v11), .Y(n84));
NOR4X1   g040(.A(n84), .B(v12), .C(n83), .D(n45), .Y(n85));
INVX1    g041(.A(v6), .Y(n86));
OR2X1    g042(.A(v10), .B(v11), .Y(n87));
NOR3X1   g043(.A(n87), .B(n67), .C(n86), .Y(n88));
OAI21X1  g044(.A0(n88), .A1(n85), .B0(n70_1), .Y(n89));
AOI21X1  g045(.A0(n89), .A1(n82), .B0(n81), .Y(v13_D_23));
INVX1    g046(.A(n46), .Y(n91));
NAND3X1  g047(.A(v7), .B(v8), .C(v9), .Y(n92));
INVX1    g048(.A(v8), .Y(n93));
NOR2X1   g049(.A(n93), .B(v11), .Y(n94));
NOR2X1   g050(.A(v12), .B(v2), .Y(n95));
NOR2X1   g051(.A(v8), .B(n70_1), .Y(n96));
AOI22X1  g052(.A0(n95), .A1(n94), .B0(v12), .B1(n96), .Y(n97));
OR2X1    g053(.A(v7), .B(v10), .Y(n98));
OAI22X1  g054(.A0(n97), .A1(n98), .B0(n92), .B1(n91), .Y(v13_D_22));
NAND2X1  g055(.A(v4), .B(v5), .Y(n100));
NOR3X1   g056(.A(n100), .B(n57), .C(v11), .Y(n101));
AOI21X1  g057(.A0(n47), .A1(v2), .B0(n101), .Y(n102));
NOR2X1   g058(.A(v10), .B(v12), .Y(n103));
INVX1    g059(.A(n103), .Y(n104));
NOR3X1   g060(.A(n104), .B(n102), .C(v7), .Y(v13_D_21));
INVX1    g061(.A(n47), .Y(n106));
NAND2X1  g062(.A(v11), .B(v12), .Y(n107));
NAND3X1  g063(.A(n68), .B(v10), .C(v3), .Y(n108));
NOR2X1   g064(.A(v1), .B(n86), .Y(n109));
NOR4X1   g065(.A(n108), .B(n107), .C(n106), .D(n109), .Y(v13_D_20));
AND2X1   g066(.A(v10), .B(v2), .Y(n111));
NAND2X1  g067(.A(v7), .B(v8), .Y(n112));
INVX1    g068(.A(n112), .Y(n113));
NAND4X1  g069(.A(n111), .B(n53), .C(n70_1), .D(n113), .Y(n114));
NOR4X1   g070(.A(n45), .B(v12), .C(n86), .D(n106), .Y(n115));
NOR2X1   g071(.A(v9), .B(v10), .Y(n116));
NOR4X1   g072(.A(v8), .B(n67), .C(v6), .D(n169), .Y(n118));
INVX1    g073(.A(v3), .Y(n119));
NOR3X1   g074(.A(v7), .B(v11), .C(n119), .Y(n120));
OAI21X1  g075(.A0(n118), .A1(n115), .B0(n120), .Y(n121));
NAND2X1  g076(.A(n121), .B(n114), .Y(v13_D_19));
NOR2X1   g077(.A(v10), .B(v11), .Y(n123));
AND2X1   g078(.A(v4), .B(v5), .Y(n124));
NAND4X1  g079(.A(n123), .B(n93), .C(n70_1), .D(n124), .Y(n125));
NOR3X1   g080(.A(n57), .B(n45), .C(v0), .Y(n126));
NOR3X1   g081(.A(n93), .B(n70_1), .C(v2), .Y(n127));
INVX1    g082(.A(v4), .Y(n128));
AOI21X1  g083(.A0(n128), .A1(n52), .B0(n84), .Y(n129));
OAI21X1  g084(.A0(n127), .A1(n126), .B0(n129), .Y(n130));
OR2X1    g085(.A(v7), .B(v12), .Y(n131));
AOI21X1  g086(.A0(n130), .A1(n125), .B0(n131), .Y(v13_D_18));
OR4X1    g087(.A(n87), .B(n64), .C(n81), .D(n100), .Y(n133));
MX2X1    g088(.A(n83), .B(n70_1), .S0(n84), .Y(n134));
AOI22X1  g089(.A0(n68), .A1(n134), .B0(v9), .B1(v11), .Y(n135));
AND2X1   g090(.A(v8), .B(v11), .Y(n136));
INVX1    g091(.A(n136), .Y(n137));
OAI22X1  g092(.A0(n135), .A1(n45), .B0(n116), .B1(n137), .Y(n138));
NAND2X1  g093(.A(v11), .B(n67), .Y(n139));
NAND2X1  g094(.A(v10), .B(v11), .Y(n140));
INVX1    g095(.A(n140), .Y(n141));
AOI21X1  g096(.A0(n141), .A1(n70_1), .B0(n67), .Y(n142));
OAI22X1  g097(.A0(n139), .A1(v10), .B0(n93), .B1(n142), .Y(n143));
AOI22X1  g098(.A0(n138), .A1(n67), .B0(v7), .B1(n143), .Y(n144));
OAI21X1  g099(.A0(n144), .A1(n62), .B0(n133), .Y(v13_D_17));
NAND4X1  g100(.A(n48), .B(n68), .C(v9), .D(n54), .Y(n146));
NAND4X1  g101(.A(v7), .B(n70_1), .C(v2), .D(n53), .Y(n147));
NAND2X1  g102(.A(v8), .B(v10), .Y(n148));
AOI21X1  g103(.A0(n147), .A1(n146), .B0(n148), .Y(v13_D_16));
NOR4X1   g104(.A(n70_1), .B(n84), .C(v2), .D(n93), .Y(n150));
OAI21X1  g105(.A0(n140), .A1(v0), .B0(n87), .Y(n151));
AOI21X1  g106(.A0(n151), .A1(n58), .B0(n150), .Y(n152));
NOR4X1   g107(.A(n131), .B(n128), .C(v5), .D(n152), .Y(v13_D_15));
AOI21X1  g108(.A0(v10), .A1(n83), .B0(n84), .Y(n154));
OAI21X1  g109(.A0(n154), .A1(v9), .B0(n93), .Y(n155));
AOI21X1  g110(.A0(v11), .A1(n62), .B0(n93), .Y(n156));
OAI22X1  g111(.A0(v11), .A1(n45), .B0(v4), .B1(v5), .Y(n157));
NOR4X1   g112(.A(n156), .B(n124), .C(v12), .D(n157), .Y(n158));
AND2X1   g113(.A(n158), .B(n155), .Y(n159));
NOR2X1   g114(.A(v9), .B(n45), .Y(n160));
OAI21X1  g115(.A0(n160), .A1(n84), .B0(n93), .Y(n161));
AOI21X1  g116(.A0(n87), .A1(v9), .B0(n93), .Y(n162));
AOI21X1  g117(.A0(n161), .A1(n76), .B0(n162), .Y(n163));
OAI21X1  g118(.A0(n159), .A1(v7), .B0(n163), .Y(v13_D_14));
MX2X1    g119(.A(v11), .B(n107), .S0(n45), .Y(n165));
OAI21X1  g120(.A0(n165), .A1(v8), .B0(n91), .Y(n166));
NOR3X1   g121(.A(n154), .B(v8), .C(v9), .Y(n167));
OAI21X1  g122(.A0(n167), .A1(n150), .B0(n124), .Y(n168));
OR2X1    g123(.A(v9), .B(v10), .Y(n169));
NAND3X1  g124(.A(n169), .B(n136), .C(v2), .Y(n170));
AOI21X1  g125(.A0(n170), .A1(n168), .B0(v12), .Y(n171));
AOI21X1  g126(.A0(n166), .A1(n70_1), .B0(n171), .Y(n172));
NAND4X1  g127(.A(v11), .B(n67), .C(v1), .D(v9), .Y(n173));
INVX1    g128(.A(v1), .Y(n174));
OAI21X1  g129(.A0(n93), .A1(n84), .B0(n131), .Y(n175));
AOI22X1  g130(.A0(n53), .A1(v8), .B0(n174), .B1(n175), .Y(n176));
OAI21X1  g131(.A0(n176), .A1(v9), .B0(n173), .Y(n177));
NOR2X1   g132(.A(v8), .B(v10), .Y(n178));
INVX1    g133(.A(n178), .Y(n179));
AOI22X1  g134(.A0(n107), .A1(n116), .B0(n46), .B1(v9), .Y(n180));
OAI22X1  g135(.A0(n179), .A1(n139), .B0(n93), .B1(n180), .Y(n181));
AOI22X1  g136(.A0(n177), .A1(v10), .B0(v7), .B1(n181), .Y(n182));
OAI21X1  g137(.A0(n172), .A1(v7), .B0(n182), .Y(v13_D_13));
NAND2X1  g138(.A(v9), .B(v10), .Y(n184));
NOR3X1   g139(.A(n184), .B(n84), .C(v12), .Y(n185));
AOI22X1  g140(.A0(n45), .A1(n124), .B0(v11), .B1(v0), .Y(n186));
OAI21X1  g141(.A0(n186), .A1(v12), .B0(n51), .Y(n187));
AOI21X1  g142(.A0(n187), .A1(n70_1), .B0(n185), .Y(n188));
OAI22X1  g143(.A0(n169), .A1(n139), .B0(v7), .B1(n188), .Y(n189));
NAND2X1  g144(.A(n70_1), .B(v12), .Y(n190));
INVX1    g145(.A(n190), .Y(n191));
NOR2X1   g146(.A(v12), .B(n62), .Y(n192));
AOI22X1  g147(.A0(n169), .A1(n192), .B0(n191), .B1(v10), .Y(n193));
OAI21X1  g148(.A0(n193), .A1(n84), .B0(n77), .Y(n194));
MX2X1    g149(.A(n189), .B(n194), .S0(v8), .Y(v13_D_12));
MX2X1    g150(.A(v10), .B(v0), .S0(v11), .Y(n196));
NOR2X1   g151(.A(n196), .B(v9), .Y(n197));
NOR2X1   g152(.A(n197), .B(v8), .Y(n198));
MX2X1    g153(.A(n62), .B(n48), .S0(n84), .Y(n199));
NOR2X1   g154(.A(n199), .B(n93), .Y(n200));
AOI21X1  g155(.A0(v8), .A1(n84), .B0(n100), .Y(n201));
NOR4X1   g156(.A(n200), .B(n198), .C(v12), .D(n201), .Y(n202));
INVX1    g157(.A(n139), .Y(n203));
AOI21X1  g158(.A0(n178), .A1(n203), .B0(n162), .Y(n204));
OAI21X1  g159(.A0(n202), .A1(v7), .B0(n204), .Y(v13_D_11));
NOR2X1   g160(.A(v7), .B(v2), .Y(n206));
OR2X1    g161(.A(n116), .B(v12), .Y(n207));
OAI22X1  g162(.A0(n206), .A1(n207), .B0(n190), .B1(n45), .Y(n208));
AOI21X1  g163(.A0(n50), .A1(n70_1), .B0(n103), .Y(n209));
NOR3X1   g164(.A(n209), .B(n68), .C(v11), .Y(n210));
AOI21X1  g165(.A0(n208), .A1(v11), .B0(n210), .Y(n211));
AOI22X1  g166(.A0(n111), .A1(n84), .B0(n93), .B1(n196), .Y(n212));
NOR3X1   g167(.A(n212), .B(v7), .C(v9), .Y(n213));
XOR2X1   g168(.A(v9), .B(v10), .Y(n214));
NAND2X1  g169(.A(n93), .B(v11), .Y(n215));
AOI22X1  g170(.A0(n47), .A1(v11), .B0(n70_1), .B1(n60_1), .Y(n216));
OAI22X1  g171(.A0(n215), .A1(n214), .B0(n100), .B1(n216), .Y(n217));
OAI21X1  g172(.A0(n217), .A1(n213), .B0(n67), .Y(n218));
OAI21X1  g173(.A0(n211), .A1(n93), .B0(n218), .Y(v13_D_10));
OAI21X1  g174(.A0(n123), .A1(n93), .B0(n140), .Y(n220));
AOI22X1  g175(.A0(n141), .A1(n93), .B0(v7), .B1(n220), .Y(n221));
OR2X1    g176(.A(n221), .B(n70_1), .Y(n222));
OAI22X1  g177(.A0(n74), .A1(v9), .B0(n83), .B1(n215), .Y(n223));
NAND3X1  g178(.A(n223), .B(n68), .C(v10), .Y(n224));
AOI21X1  g179(.A0(n224), .A1(n222), .B0(v12), .Y(v13_D_9));
OAI21X1  g180(.A0(v12), .A1(v0), .B0(v11), .Y(n226));
AND2X1   g181(.A(n226), .B(n70_1), .Y(n227));
AOI21X1  g182(.A0(n227), .A1(n91), .B0(v8), .Y(n228));
NAND2X1  g183(.A(n111), .B(n67), .Y(n229));
OAI21X1  g184(.A0(n45), .A1(v12), .B0(v8), .Y(n230));
AOI21X1  g185(.A0(n230), .A1(n229), .B0(v11), .Y(n231));
AOI21X1  g186(.A0(n70_1), .A1(v11), .B0(v12), .Y(n232));
NOR2X1   g187(.A(n232), .B(v10), .Y(n233));
AOI22X1  g188(.A0(v9), .A1(n62), .B0(v11), .B1(n93), .Y(n234));
NOR2X1   g189(.A(v4), .B(n52), .Y(n235));
OAI22X1  g190(.A0(n234), .A1(n235), .B0(n203), .B1(n70_1), .Y(n236));
NOR4X1   g191(.A(n233), .B(n231), .C(n228), .D(n236), .Y(n237));
NOR2X1   g192(.A(n93), .B(v10), .Y(n238));
MX2X1    g193(.A(v12), .B(n84), .S0(v9), .Y(n239));
AOI21X1  g194(.A0(n107), .A1(n70_1), .B0(n54), .Y(n240));
OAI22X1  g195(.A0(n179), .A1(n139), .B0(n148), .B1(n240), .Y(n241));
AOI22X1  g196(.A0(n239), .A1(n238), .B0(v7), .B1(n241), .Y(n242));
OAI21X1  g197(.A0(n237), .A1(v7), .B0(n242), .Y(v13_D_8));
INVX1    g198(.A(n94), .Y(n244));
AOI22X1  g199(.A0(n191), .A1(n45), .B0(n67), .B1(n169), .Y(n245));
OR4X1    g200(.A(n70_1), .B(n84), .C(v12), .D(n238), .Y(n246));
OAI21X1  g201(.A0(n245), .A1(n244), .B0(n246), .Y(n247));
OAI21X1  g202(.A0(n107), .A1(v10), .B0(n91), .Y(n248));
AOI22X1  g203(.A0(n111), .A1(n54), .B0(n93), .B1(n248), .Y(n249));
AOI21X1  g204(.A0(n128), .A1(v5), .B0(v12), .Y(n250));
OAI21X1  g205(.A0(n150), .A1(n126), .B0(n250), .Y(n251));
OAI21X1  g206(.A0(n249), .A1(v9), .B0(n251), .Y(n252));
MX2X1    g207(.A(n247), .B(n252), .S0(n68), .Y(v13_D_7));
AND2X1   g208(.A(v9), .B(v12), .Y(n254));
MX2X1    g209(.A(n71), .B(n87), .S0(v12), .Y(n255));
AOI22X1  g210(.A0(n254), .A1(n123), .B0(n70_1), .B1(n255), .Y(n256));
INVX1    g211(.A(n50), .Y(n257));
OR2X1    g212(.A(n111), .B(v11), .Y(n258));
AOI21X1  g213(.A0(v9), .A1(n62), .B0(n84), .Y(n259));
NOR2X1   g214(.A(n259), .B(v12), .Y(n260));
AOI21X1  g215(.A0(n260), .A1(n258), .B0(n93), .Y(n261));
OAI21X1  g216(.A0(v4), .A1(n52), .B0(n45), .Y(n262));
AOI21X1  g217(.A0(n262), .A1(n67), .B0(v11), .Y(n263));
AOI21X1  g218(.A0(n179), .A1(n203), .B0(n70_1), .Y(n264));
NOR4X1   g219(.A(n263), .B(n261), .C(n257), .D(n264), .Y(n265));
OAI22X1  g220(.A0(n256), .A1(n93), .B0(v7), .B1(n265), .Y(v13_D_6));
INVX1    g221(.A(CLR), .Y(n267));
NAND4X1  g222(.A(n45), .B(v11), .C(n67), .D(v9), .Y(n268));
AOI21X1  g223(.A0(n100), .A1(n62), .B0(n139), .Y(n269));
OAI21X1  g224(.A0(n269), .A1(n70_1), .B0(v10), .Y(n270));
AOI21X1  g225(.A0(n270), .A1(n268), .B0(n93), .Y(n271));
NOR3X1   g226(.A(v9), .B(v11), .C(v12), .Y(n272));
NAND4X1  g227(.A(n174), .B(v3), .C(v6), .D(v8), .Y(n273));
OAI22X1  g228(.A0(n100), .A1(n64), .B0(n107), .B1(n273), .Y(n274));
AOI21X1  g229(.A0(n274), .A1(n83), .B0(n272), .Y(n275));
NAND4X1  g230(.A(n70_1), .B(v12), .C(v6), .D(n123), .Y(n276));
OAI21X1  g231(.A0(n140), .A1(n70_1), .B0(n276), .Y(n277));
NAND4X1  g232(.A(v10), .B(v11), .C(v0), .D(v8), .Y(n278));
OAI22X1  g233(.A0(n109), .A1(n278), .B0(n87), .B1(n57), .Y(n279));
AND2X1   g234(.A(v12), .B(v3), .Y(n280));
AOI22X1  g235(.A0(n279), .A1(n280), .B0(n277), .B1(n93), .Y(n281));
OAI21X1  g236(.A0(n275), .A1(n45), .B0(n281), .Y(n282));
OAI21X1  g237(.A0(n282), .A1(n271), .B0(n68), .Y(n283));
AOI22X1  g238(.A0(n203), .A1(n93), .B0(n64), .B1(n94), .Y(n284));
OAI22X1  g239(.A0(n139), .A1(n184), .B0(v10), .B1(n284), .Y(n285));
NOR3X1   g240(.A(n140), .B(n93), .C(v9), .Y(n286));
NOR3X1   g241(.A(n131), .B(n174), .C(n86), .Y(n287));
NOR3X1   g242(.A(n87), .B(v8), .C(n70_1), .Y(n288));
AOI21X1  g243(.A0(n288), .A1(n287), .B0(n286), .Y(n289));
OAI22X1  g244(.A0(n148), .A1(n64), .B0(v2), .B1(n289), .Y(n290));
AOI21X1  g245(.A0(n285), .A1(v7), .B0(n290), .Y(n291));
AOI21X1  g246(.A0(n291), .A1(n283), .B0(n267), .Y(n55));
NOR3X1   g247(.A(n83), .B(v1), .C(n86), .Y(n293));
NOR3X1   g248(.A(n293), .B(n67), .C(n119), .Y(n294));
OAI21X1  g249(.A0(n294), .A1(n84), .B0(v9), .Y(n295));
MX2X1    g250(.A(v10), .B(n124), .S0(v9), .Y(n296));
AOI21X1  g251(.A0(n70_1), .A1(n119), .B0(n139), .Y(n297));
OAI22X1  g252(.A0(v10), .A1(n297), .B0(v11), .B1(n67), .Y(n298));
AOI21X1  g253(.A0(n296), .A1(n95), .B0(n298), .Y(n299));
AOI21X1  g254(.A0(n299), .A1(n295), .B0(n93), .Y(n300));
NAND3X1  g255(.A(v9), .B(n45), .C(n174), .Y(n301));
OAI21X1  g256(.A0(n140), .A1(v9), .B0(n301), .Y(n302));
NAND3X1  g257(.A(n302), .B(n93), .C(n67), .Y(n303));
NAND2X1  g258(.A(n93), .B(v9), .Y(n304));
OAI22X1  g259(.A0(n304), .A1(n104), .B0(n190), .B1(v11), .Y(n305));
NOR2X1   g260(.A(n165), .B(n70_1), .Y(n306));
AOI21X1  g261(.A0(n305), .A1(n86), .B0(n306), .Y(n307));
NAND3X1  g262(.A(n307), .B(n303), .C(n51), .Y(n308));
OAI21X1  g263(.A0(n308), .A1(n300), .B0(n68), .Y(n309));
OR4X1    g264(.A(n107), .B(v9), .C(n45), .D(n112), .Y(n310));
NAND3X1  g265(.A(n103), .B(n68), .C(v9), .Y(n311));
AOI21X1  g266(.A0(n311), .A1(n310), .B0(n62), .Y(n312));
AOI22X1  g267(.A0(n160), .A1(n94), .B0(v11), .B1(n178), .Y(n313));
AOI22X1  g268(.A0(n94), .A1(v12), .B0(n203), .B1(n96), .Y(n314));
OAI22X1  g269(.A0(n313), .A1(n77), .B0(v10), .B1(n314), .Y(n315));
NOR2X1   g270(.A(n315), .B(n312), .Y(n316));
AOI21X1  g271(.A0(n316), .A1(n309), .B0(n267), .Y(n60));
NOR3X1   g272(.A(n293), .B(n107), .C(n119), .Y(n318));
NOR3X1   g273(.A(v11), .B(v12), .C(v6), .Y(n319));
OAI21X1  g274(.A0(n319), .A1(n318), .B0(v9), .Y(n320));
MX2X1    g275(.A(v11), .B(n100), .S0(n67), .Y(n321));
OAI21X1  g276(.A0(n192), .A1(v11), .B0(n104), .Y(n322));
AOI22X1  g277(.A0(n321), .A1(n45), .B0(n70_1), .B1(n322), .Y(n323));
AOI21X1  g278(.A0(n323), .A1(n320), .B0(n93), .Y(n324));
NOR2X1   g279(.A(n100), .B(v12), .Y(n325));
MX2X1    g280(.A(n47), .B(n178), .S0(v12), .Y(n326));
AOI22X1  g281(.A0(n325), .A1(n116), .B0(n119), .B1(n326), .Y(n327));
NOR2X1   g282(.A(v8), .B(n67), .Y(n328));
AOI21X1  g283(.A0(n84), .A1(v6), .B0(v9), .Y(n329));
OAI22X1  g284(.A0(n140), .A1(v9), .B0(v10), .B1(n329), .Y(n330));
MX2X1    g285(.A(v8), .B(n96), .S0(v10), .Y(n331));
AOI22X1  g286(.A0(n330), .A1(n328), .B0(n192), .B1(n331), .Y(n332));
OAI21X1  g287(.A0(n327), .A1(v11), .B0(n332), .Y(n333));
OAI21X1  g288(.A0(n333), .A1(n324), .B0(n68), .Y(n334));
NAND3X1  g289(.A(n70_1), .B(v10), .C(v12), .Y(n335));
OAI21X1  g290(.A0(n191), .A1(v10), .B0(n335), .Y(n336));
AOI21X1  g291(.A0(v8), .A1(n45), .B0(v11), .Y(n337));
NOR4X1   g292(.A(n68), .B(n70_1), .C(v12), .D(n337), .Y(n338));
AOI21X1  g293(.A0(n336), .A1(n94), .B0(n338), .Y(n339));
AOI21X1  g294(.A0(n339), .A1(n334), .B0(n267), .Y(n65));
NAND4X1  g295(.A(v10), .B(n84), .C(n67), .D(n70_1), .Y(n341));
NAND2X1  g296(.A(v12), .B(v1), .Y(n342));
AOI21X1  g297(.A0(n342), .A1(n70_1), .B0(n137), .Y(n343));
NOR4X1   g298(.A(n70_1), .B(v11), .C(v12), .D(v8), .Y(n344));
OAI21X1  g299(.A0(n344), .A1(n343), .B0(n45), .Y(n345));
AOI21X1  g300(.A0(n345), .A1(n341), .B0(n62), .Y(n346));
INVX1    g301(.A(n54), .Y(n347));
OAI22X1  g302(.A0(n74), .A1(n107), .B0(n347), .B1(n304), .Y(n348));
AOI22X1  g303(.A0(n272), .A1(n124), .B0(n174), .B1(n348), .Y(n349));
NAND4X1  g304(.A(v9), .B(n67), .C(n86), .D(n123), .Y(n350));
NOR2X1   g305(.A(n45), .B(v12), .Y(n351));
NAND2X1  g306(.A(v11), .B(n83), .Y(n352));
AOI22X1  g307(.A0(n53), .A1(n45), .B0(n351), .B1(n352), .Y(n353));
OAI21X1  g308(.A0(n353), .A1(v9), .B0(n350), .Y(n354));
NOR3X1   g309(.A(n64), .B(v8), .C(n45), .Y(n355));
NOR4X1   g310(.A(n70_1), .B(v10), .C(n84), .D(n93), .Y(n356));
OAI21X1  g311(.A0(n356), .A1(n355), .B0(n100), .Y(n357));
NOR3X1   g312(.A(n87), .B(v12), .C(n119), .Y(n358));
AND2X1   g313(.A(n254), .B(n140), .Y(n359));
OAI21X1  g314(.A0(n359), .A1(n358), .B0(v8), .Y(n360));
NAND4X1  g315(.A(v10), .B(n84), .C(v12), .D(v9), .Y(n361));
NAND3X1  g316(.A(n361), .B(n360), .C(n357), .Y(n362));
AOI21X1  g317(.A0(n354), .A1(n93), .B0(n362), .Y(n363));
OAI21X1  g318(.A0(n349), .A1(v10), .B0(n363), .Y(n364));
OAI21X1  g319(.A0(n364), .A1(n346), .B0(n68), .Y(n365));
NOR4X1   g320(.A(v8), .B(n67), .C(v6), .D(v7), .Y(n366));
NOR2X1   g321(.A(n93), .B(v12), .Y(n367));
OAI21X1  g322(.A0(n367), .A1(n366), .B0(n119), .Y(n368));
OAI21X1  g323(.A0(n244), .A1(v12), .B0(n368), .Y(n369));
AOI21X1  g324(.A0(v10), .A1(n84), .B0(n67), .Y(n370));
OAI21X1  g325(.A0(n111), .A1(n84), .B0(n370), .Y(n371));
AOI22X1  g326(.A0(n87), .A1(n67), .B0(n70_1), .B1(n371), .Y(n372));
OAI22X1  g327(.A0(n160), .A1(n139), .B0(n93), .B1(n372), .Y(n373));
AOI22X1  g328(.A0(n369), .A1(n116), .B0(v7), .B1(n373), .Y(n374));
AOI21X1  g329(.A0(n374), .A1(n365), .B0(n267), .Y(n70));
NOR2X1   g330(.A(n45), .B(v11), .Y(n376));
OR2X1    g331(.A(v3), .B(v6), .Y(n377));
AOI21X1  g332(.A0(n377), .A1(n84), .B0(v10), .Y(n378));
OAI21X1  g333(.A0(n378), .A1(n376), .B0(v12), .Y(n379));
AOI22X1  g334(.A0(n151), .A1(n325), .B0(n91), .B1(v9), .Y(n380));
AOI21X1  g335(.A0(n380), .A1(n379), .B0(v8), .Y(n381));
NOR3X1   g336(.A(n107), .B(v10), .C(v1), .Y(n382));
OAI21X1  g337(.A0(n50), .A1(v3), .B0(n70_1), .Y(n383));
AOI21X1  g338(.A0(n383), .A1(n93), .B0(n382), .Y(n384));
AOI22X1  g339(.A0(n116), .A1(n367), .B0(n53), .B1(v9), .Y(n385));
OAI21X1  g340(.A0(n384), .A1(n62), .B0(n385), .Y(n386));
OAI21X1  g341(.A0(n386), .A1(n381), .B0(n68), .Y(n387));
MX2X1    g342(.A(n70_1), .B(v8), .S0(n45), .Y(n388));
AOI21X1  g343(.A0(n70_1), .A1(v12), .B0(n84), .Y(n389));
MX2X1    g344(.A(n139), .B(n389), .S0(n45), .Y(n390));
OAI22X1  g345(.A0(n388), .A1(n139), .B0(n93), .B1(n390), .Y(n391));
OAI22X1  g346(.A0(n190), .A1(n68), .B0(n45), .B1(n139), .Y(n392));
NAND3X1  g347(.A(n124), .B(v8), .C(n67), .Y(n393));
OAI21X1  g348(.A0(n342), .A1(v10), .B0(n393), .Y(n394));
NOR2X1   g349(.A(v7), .B(n84), .Y(n395));
AOI22X1  g350(.A0(n394), .A1(n395), .B0(n392), .B1(v8), .Y(n396));
AOI22X1  g351(.A0(n70_1), .A1(v12), .B0(v3), .B1(n103), .Y(n397));
OAI22X1  g352(.A0(n396), .A1(v2), .B0(n244), .B1(n397), .Y(n398));
AOI21X1  g353(.A0(n391), .A1(v7), .B0(n398), .Y(n399));
AOI21X1  g354(.A0(n399), .A1(n387), .B0(n267), .Y(n75));
NOR3X1   g355(.A(v8), .B(v11), .C(v12), .Y(n401));
AOI21X1  g356(.A0(n53), .A1(v6), .B0(n401), .Y(n402));
OR2X1    g357(.A(n402), .B(v1), .Y(n403));
OAI21X1  g358(.A0(n93), .A1(v11), .B0(v10), .Y(n404));
OR2X1    g359(.A(n401), .B(n53), .Y(n405));
AOI22X1  g360(.A0(n404), .A1(v12), .B0(n119), .B1(n405), .Y(n406));
AOI21X1  g361(.A0(n406), .A1(n403), .B0(n70_1), .Y(n407));
NOR3X1   g362(.A(v9), .B(n45), .C(v0), .Y(n408));
NAND4X1  g363(.A(n124), .B(v11), .C(n67), .D(n408), .Y(n409));
AOI21X1  g364(.A0(v10), .A1(n67), .B0(n84), .Y(n410));
AOI21X1  g365(.A0(n45), .A1(v6), .B0(n347), .Y(n411));
OAI21X1  g366(.A0(n411), .A1(n410), .B0(v9), .Y(n412));
AOI21X1  g367(.A0(n412), .A1(n409), .B0(v8), .Y(n413));
OAI21X1  g368(.A0(n413), .A1(n407), .B0(n68), .Y(n414));
OAI22X1  g369(.A0(n190), .A1(n141), .B0(n70_1), .B1(n87), .Y(n415));
NOR2X1   g370(.A(v8), .B(v11), .Y(n416));
AOI21X1  g371(.A0(n136), .A1(n124), .B0(n416), .Y(n417));
NAND3X1  g372(.A(n68), .B(v9), .C(n67), .Y(n418));
OAI22X1  g373(.A0(n417), .A1(n418), .B0(n112), .B1(n190), .Y(n419));
AOI22X1  g374(.A0(n415), .A1(n113), .B0(n62), .B1(n419), .Y(n420));
AOI21X1  g375(.A0(n420), .A1(n414), .B0(n267), .Y(n80));
endmodule
