//Converted to Combinational (Partial output: n80) , Module name: s1494_n80 , Timestamp: 2018-12-03T15:51:02.662855 
module s1494_n80 ( v1, CLR, v7, v8, v2, v9, v1, v12, v11, v10, v6, v3, v0, v5, v4, n80 );
input v1, CLR, v7, v8, v2, v9, v1, v12, v11, v10, v6, v3, v0, v5, v4;
output n80;
wire n267, n414, n420, n68, n407, n413, n419, n62, n113, n415, n70_1, n403, n406, n409, n412, n190, n112, n418, n417, n87, n141, n402, n405, n119, n404, n408, n67, n124, n410, n411, n416, n136, n140, n401, n53, n93, n45, n84, n347, n54;
AOI21X1  g375(.A0(n420), .A1(n414), .B0(n267), .Y(n80));
INVX1    g221(.A(CLR), .Y(n267));
OAI21X1  g368(.A0(n413), .A1(n407), .B0(n68), .Y(n414));
AOI22X1  g374(.A0(n415), .A1(n113), .B0(n62), .B1(n419), .Y(n420));
INVX1    g023(.A(v7), .Y(n68));
AOI21X1  g361(.A0(n406), .A1(n403), .B0(n70_1), .Y(n407));
AOI21X1  g367(.A0(n412), .A1(n409), .B0(v8), .Y(n413));
OAI22X1  g373(.A0(n417), .A1(n418), .B0(n112), .B1(n190), .Y(n419));
INVX1    g017(.A(v2), .Y(n62));
INVX1    g068(.A(n112), .Y(n113));
OAI22X1  g369(.A0(n190), .A1(n141), .B0(n70_1), .B1(n87), .Y(n415));
INVX1    g025(.A(v9), .Y(n70_1));
OR2X1    g357(.A(n402), .B(v1), .Y(n403));
AOI22X1  g360(.A0(n404), .A1(v12), .B0(n119), .B1(n405), .Y(n406));
NAND4X1  g363(.A(n124), .B(v11), .C(n67), .D(n408), .Y(n409));
OAI21X1  g366(.A0(n411), .A1(n410), .B0(v9), .Y(n412));
NAND2X1  g144(.A(n70_1), .B(v12), .Y(n190));
NAND2X1  g067(.A(v7), .B(v8), .Y(n112));
NAND3X1  g372(.A(n68), .B(v9), .C(n67), .Y(n418));
AOI21X1  g371(.A0(n136), .A1(n124), .B0(n416), .Y(n417));
OR2X1    g042(.A(v10), .B(v11), .Y(n87));
INVX1    g095(.A(n140), .Y(n141));
AOI21X1  g356(.A0(n53), .A1(v6), .B0(n401), .Y(n402));
OR2X1    g359(.A(n401), .B(n53), .Y(n405));
INVX1    g073(.A(v3), .Y(n119));
OAI21X1  g358(.A0(n93), .A1(v11), .B0(v10), .Y(n404));
NOR3X1   g362(.A(v9), .B(n45), .C(v0), .Y(n408));
INVX1    g022(.A(v12), .Y(n67));
AND2X1   g078(.A(v4), .B(v5), .Y(n124));
AOI21X1  g364(.A0(v10), .A1(n67), .B0(n84), .Y(n410));
AOI21X1  g365(.A0(n45), .A1(v6), .B0(n347), .Y(n411));
NOR2X1   g370(.A(v8), .B(v11), .Y(n416));
AND2X1   g090(.A(v8), .B(v11), .Y(n136));
NAND2X1  g094(.A(v10), .B(v11), .Y(n140));
NOR3X1   g355(.A(v8), .B(v11), .C(v12), .Y(n401));
AND2X1   g008(.A(v11), .B(v12), .Y(n53));
INVX1    g048(.A(v8), .Y(n93));
INVX1    g000(.A(v10), .Y(n45));
INVX1    g039(.A(v11), .Y(n84));
INVX1    g301(.A(n54), .Y(n347));
NOR2X1   g009(.A(v11), .B(v12), .Y(n54));

endmodule
