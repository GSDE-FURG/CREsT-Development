//Converted to Combinational (Partial output: G542) , Module name: s1196_G542
module s1196_G542 ( G4, G1, G3, G10, G7, G8, G9, G13, G6, G34, G46, G12, G11, G5, G31, G30, G2, G0, G542 );
input G4, G3, G1, G10, G7, G8, G9, G13, G6, G34, G46, G12, G11, G5, G31, G30, G2, G0;
output G542;
wire n285, n293, n283, n284, n292, n286, n157, n287, n86, n115, n209, n87_1, n112_1, n256, n288, n290, n291, n130, n205, n111, n137_1, n289, n116, n129, n121, n125, n106, n110, n126, n88, n128, n118, n120, n122_1, n123, n124, n105, n109, n85, n94, n127_1, n117_1, n114, n119, n108, n113, n107_1;
NAND2X1  g212(.A(n293), .B(n285), .Y(G542));
NAND2X1  g203(.A(n284), .B(n283), .Y(n285));
AOI22X1  g211(.A0(n287), .A1(n157), .B0(n286), .B1(n292), .Y(n293));
NOR3X1   g201(.A(G10), .B(n115), .C(n86), .Y(n283));
OAI22X1  g202(.A0(n256), .A1(n112_1), .B0(n87_1), .B1(n209), .Y(n284));
NAND3X1  g210(.A(n291), .B(n290), .C(n288), .Y(n292));
NOR2X1   g204(.A(n209), .B(n87_1), .Y(n286));
AND2X1   g075(.A(G10), .B(G7), .Y(n157));
AOI21X1  g205(.A0(G9), .A1(G8), .B0(n256), .Y(n287));
INVX1    g004(.A(G7), .Y(n86));
INVX1    g033(.A(G9), .Y(n115));
OR4X1    g127(.A(n111), .B(G13), .C(n205), .D(n130), .Y(n209));
INVX1    g005(.A(G6), .Y(n87_1));
INVX1    g030(.A(G8), .Y(n112_1));
INVX1    g174(.A(G34), .Y(n256));
INVX1    g206(.A(n137_1), .Y(n288));
NAND2X1  g208(.A(n289), .B(n115), .Y(n290));
OAI21X1  g209(.A0(n115), .A1(n86), .B0(n116), .Y(n291));
NAND4X1  g048(.A(n125), .B(n121), .C(G46), .D(n129), .Y(n130));
INVX1    g123(.A(G12), .Y(n205));
NOR2X1   g029(.A(n110), .B(n106), .Y(n111));
NOR4X1   g055(.A(n88), .B(n115), .C(G8), .D(n126), .Y(n137_1));
OAI21X1  g207(.A0(G8), .A1(n86), .B0(n88), .Y(n289));
AND2X1   g034(.A(G10), .B(G8), .Y(n116));
NAND4X1  g047(.A(n126), .B(G9), .C(n86), .D(n128), .Y(n129));
OAI21X1  g039(.A0(n120), .A1(n118), .B0(G11), .Y(n121));
NAND3X1  g043(.A(n124), .B(n123), .C(n122_1), .Y(n125));
NOR2X1   g024(.A(G5), .B(n105), .Y(n106));
AOI22X1  g028(.A0(n94), .A1(G3), .B0(n85), .B1(n109), .Y(n110));
INVX1    g044(.A(G11), .Y(n126));
INVX1    g006(.A(G10), .Y(n88));
MX2X1    g046(.A(G10), .B(n127_1), .S0(G8), .Y(n128));
NOR4X1   g036(.A(n114), .B(G31), .C(n112_1), .D(n117_1), .Y(n118));
OAI22X1  g038(.A0(G30), .A1(G6), .B0(G9), .B1(n119), .Y(n120));
NAND3X1  g040(.A(G30), .B(G7), .C(n87_1), .Y(n122_1));
NOR3X1   g041(.A(G11), .B(G10), .C(G9), .Y(n123));
NAND2X1  g042(.A(G31), .B(G8), .Y(n124));
INVX1    g023(.A(G4), .Y(n105));
AOI21X1  g027(.A0(n108), .A1(G2), .B0(G3), .Y(n109));
INVX1    g003(.A(G5), .Y(n85));
NOR2X1   g012(.A(G4), .B(G0), .Y(n94));
INVX1    g045(.A(G31), .Y(n127_1));
NOR2X1   g035(.A(n116), .B(n115), .Y(n117_1));
NOR3X1   g032(.A(n113), .B(n86), .C(G6), .Y(n114));
OR2X1    g037(.A(G8), .B(G7), .Y(n119));
OAI22X1  g026(.A0(n85), .A1(G1), .B0(n105), .B1(n107_1), .Y(n108));
INVX1    g031(.A(G30), .Y(n113));
AND2X1   g025(.A(G5), .B(G3), .Y(n107_1));

endmodule
