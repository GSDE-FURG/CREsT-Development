//Converted to Combinational (Partial output: g9299) , Module name: s13207_g9299 , Timestamp: 2018-12-03T15:51:04.657357 
module s13207_g9299 ( g2, g71, g77, g62, g619, g764, g772, g756, g702, g465, g677, g718, g68, g41, g45, g86, g52, g83, g74, g158, g181, g432, g384, g547, g598, g134, g100, g622, g630, g270, g222, g303, g351, g606, g611, g80, g42, g55, g44, g846, g863, g652, g513, g9299 );
input g2, g71, g77, g62, g619, g764, g772, g756, g702, g465, g677, g718, g68, g41, g45, g86, g52, g83, g74, g158, g181, g432, g384, g547, g598, g134, g100, g622, g630, g270, g222, g303, g351, g606, g611, g80, g42, g55, g44, g846, g863, g652, g513;
output g9299;
wire n2464, n2463, n2338, n2448, n2362_1, n2462_1, n2337_1, n2323, n2328, n2331, n2286, n2447_1, n2441, n2361, n2339, n2340, n2345, n2461, n2452_1, n2453, n2456, n2333, n2336, n2320, n2321, n2322_1, n2325, n2327_1, n2329, n2330, n2275, n2277, n2285, n2314, n2445, n2446, n2440, n2434, n2438, n2439, n2350, n2355, n2360, n2248, n2238, n2240, n2206, n2344, n2341, n2342_1, n2343, n2460, n2457_1, n2458, n2459, n2449, n2450, n2451, n2349, n2454, n2455, n2332_1, n2335, n2250, n2334, n2319, n2230, n2274, n2235, n2264, n2266_1, n2276, n2200, n2324, n2268, n2326, n2191, n2263, n2293_1, n2233_1, n2279, n2281, n2284, n2313, n2290, n2304, n2306, n2307_1, n2296, n2444, n2311, n2309, n2251_1, n2246, n2254, n2237_1, n2243, n2245, n2437_1, n2253, n2386, n2346, n2347_1, n2348, n2354, n2351, n2352_1, n2353, n2359, n2356, n2357_1, n2358, n2232, n2229, n2247_1, n2227, n2226, n2239, n2283_1, n2280, n2282, n1899, n2241, n2190, n2273_1, n2278_1, n2252, n2312_1, n2310, n2289, n2303, n2300, n2287, n2288_1, n2299, n2305, n2295, n2442_1, n2443, n2188, n2249, n2231, n2234, n2236, n2242_1, n2244, n2435, n2436, n2298, n2291, n2292, n2294, n2189_1;
NAND2X1  g0335(.A(n2464), .B(g62), .Y(g9299));
AOI21X1  g0334(.A0(n2448), .A1(n2338), .B0(n2463), .Y(n2464));
AOI21X1  g0333(.A0(n2462_1), .A1(n2362_1), .B0(n2338), .Y(n2463));
NOR4X1   g0210(.A(n2331), .B(n2328), .C(n2323), .D(n2337_1), .Y(n2338));
MX2X1    g0318(.A(n2441), .B(n2447_1), .S0(n2286), .Y(n2448));
OR4X1    g0234(.A(n2345), .B(n2340), .C(n2339), .D(n2361), .Y(n2362_1));
NOR4X1   g0332(.A(n2456), .B(n2453), .C(n2452_1), .D(n2461), .Y(n2462_1));
OR2X1    g0209(.A(n2336), .B(n2333), .Y(n2337_1));
NAND3X1  g0195(.A(n2322_1), .B(n2321), .C(n2320), .Y(n2323));
NAND2X1  g0200(.A(n2327_1), .B(n2325), .Y(n2328));
NAND2X1  g0203(.A(n2330), .B(n2329), .Y(n2331));
NAND3X1  g0158(.A(n2285), .B(n2277), .C(n2275), .Y(n2286));
NAND3X1  g0317(.A(n2446), .B(n2445), .C(n2314), .Y(n2447_1));
NAND4X1  g0311(.A(n2439), .B(n2438), .C(n2434), .D(n2440), .Y(n2441));
NAND3X1  g0233(.A(n2360), .B(n2355), .C(n2350), .Y(n2361));
NOR3X1   g0211(.A(n2240), .B(n2238), .C(n2248), .Y(n2339));
NOR3X1   g0212(.A(n2240), .B(n2238), .C(n2206), .Y(n2340));
OR4X1    g0217(.A(n2343), .B(n2342_1), .C(n2341), .D(n2344), .Y(n2345));
NAND4X1  g0331(.A(n2459), .B(n2458), .C(n2457_1), .D(n2460), .Y(n2461));
NAND3X1  g0322(.A(n2451), .B(n2450), .C(n2449), .Y(n2452_1));
AND2X1   g0323(.A(n2349), .B(g619), .Y(n2453));
NAND2X1  g0326(.A(n2455), .B(n2454), .Y(n2456));
OAI21X1  g0205(.A0(n2240), .A1(n2206), .B0(n2332_1), .Y(n2333));
OAI21X1  g0208(.A0(n2334), .A1(n2250), .B0(n2335), .Y(n2336));
OAI21X1  g0192(.A0(n2274), .A1(n2230), .B0(n2319), .Y(n2320));
OAI21X1  g0193(.A0(n2264), .A1(n2235), .B0(n2319), .Y(n2321));
OAI21X1  g0194(.A0(n2276), .A1(n2266_1), .B0(n2319), .Y(n2322_1));
OAI21X1  g0197(.A0(n2324), .A1(n2200), .B0(n2319), .Y(n2325));
OAI21X1  g0199(.A0(n2326), .A1(n2268), .B0(n2319), .Y(n2327_1));
AOI22X1  g0201(.A0(n2293_1), .A1(n2319), .B0(n2263), .B1(n2191), .Y(n2329));
OAI21X1  g0202(.A0(n2233_1), .A1(n2191), .B0(n2319), .Y(n2330));
OAI21X1  g0147(.A0(n2274), .A1(n2235), .B0(n2263), .Y(n2275));
OAI21X1  g0149(.A0(n2276), .A1(n2230), .B0(n2263), .Y(n2277));
NOR3X1   g0157(.A(n2284), .B(n2281), .C(n2279), .Y(n2285));
OR4X1    g0186(.A(n2306), .B(n2304), .C(n2290), .D(n2313), .Y(n2314));
OAI21X1  g0315(.A0(n2444), .A1(n2296), .B0(n2307_1), .Y(n2445));
AOI22X1  g0316(.A0(n2309), .A1(g772), .B0(g764), .B1(n2311), .Y(n2446));
AOI22X1  g0310(.A0(n2246), .A1(g702), .B0(g756), .B1(n2251_1), .Y(n2440));
OR4X1    g0304(.A(n2245), .B(n2243), .C(n2237_1), .D(n2254), .Y(n2434));
AOI21X1  g0308(.A0(n2243), .A1(g465), .B0(n2437_1), .Y(n2438));
AOI22X1  g0309(.A0(n2386), .A1(g718), .B0(g677), .B1(n2253), .Y(n2439));
NOR4X1   g0222(.A(n2348), .B(n2347_1), .C(n2346), .D(n2349), .Y(n2350));
NOR4X1   g0227(.A(n2353), .B(n2352_1), .C(n2351), .D(n2354), .Y(n2355));
NOR4X1   g0232(.A(n2358), .B(n2357_1), .C(n2356), .D(n2359), .Y(n2360));
NAND4X1  g0120(.A(g68), .B(n2247_1), .C(n2229), .D(n2232), .Y(n2248));
OR4X1    g0110(.A(n2226), .B(g45), .C(g41), .D(n2227), .Y(n2238));
OR4X1    g0112(.A(g83), .B(g52), .C(n2239), .D(g86), .Y(n2240));
OR4X1    g0078(.A(g68), .B(g74), .C(g77), .D(g71), .Y(n2206));
NOR3X1   g0216(.A(n2334), .B(n2250), .C(n2238), .Y(n2344));
NOR3X1   g0213(.A(n2334), .B(n2283_1), .C(n2238), .Y(n2341));
NOR3X1   g0214(.A(n2334), .B(n2280), .C(n2238), .Y(n2342_1));
NOR3X1   g0215(.A(n2334), .B(n2282), .C(n2238), .Y(n2343));
AOI22X1  g0330(.A0(n2358), .A1(g181), .B0(g158), .B1(n2359), .Y(n2460));
AOI22X1  g0327(.A0(n2351), .A1(g384), .B0(g432), .B1(n2352_1), .Y(n2457_1));
AOI22X1  g0328(.A0(n2346), .A1(g598), .B0(g547), .B1(n2353), .Y(n2458));
AOI22X1  g0329(.A0(n2356), .A1(g100), .B0(g134), .B1(n2357_1), .Y(n2459));
AOI22X1  g0319(.A0(n2339), .A1(g630), .B0(g622), .B1(n2340), .Y(n2449));
AOI22X1  g0320(.A0(n2341), .A1(g222), .B0(g270), .B1(n2342_1), .Y(n2450));
AOI22X1  g0321(.A0(n2343), .A1(g351), .B0(g303), .B1(n2344), .Y(n2451));
NOR2X1   g0221(.A(n2332_1), .B(n2238), .Y(n2349));
NAND4X1  g0324(.A(n2266_1), .B(n1899), .C(g606), .D(n2319), .Y(n2454));
NAND2X1  g0325(.A(n2348), .B(g611), .Y(n2455));
NAND4X1  g0204(.A(n2241), .B(g71), .C(g68), .D(n2319), .Y(n2332_1));
NAND4X1  g0207(.A(n2241), .B(g71), .C(n2190), .D(n2319), .Y(n2335));
NAND4X1  g0122(.A(n2190), .B(g74), .C(n2229), .D(g71), .Y(n2250));
OR4X1    g0206(.A(g83), .B(g52), .C(g80), .D(g86), .Y(n2334));
NOR4X1   g0191(.A(g83), .B(g52), .C(g80), .D(g86), .Y(n2319));
NOR4X1   g0102(.A(n2190), .B(g74), .C(n2229), .D(g71), .Y(n2230));
INVX1    g0146(.A(n2273_1), .Y(n2274));
NOR4X1   g0107(.A(g68), .B(g74), .C(n2229), .D(g71), .Y(n2235));
NOR4X1   g0136(.A(g68), .B(n2247_1), .C(n2229), .D(g71), .Y(n2264));
NOR4X1   g0138(.A(n2190), .B(n2247_1), .C(n2229), .D(g71), .Y(n2266_1));
NOR4X1   g0148(.A(n2190), .B(g74), .C(n2229), .D(n2232), .Y(n2276));
NOR4X1   g0072(.A(g68), .B(g74), .C(g77), .D(g71), .Y(n2200));
NOR4X1   g0196(.A(g68), .B(n2247_1), .C(g77), .D(g71), .Y(n2324));
NOR4X1   g0140(.A(n2190), .B(g74), .C(g77), .D(n2232), .Y(n2268));
NOR4X1   g0198(.A(n2190), .B(n2247_1), .C(g77), .D(g71), .Y(n2326));
NOR4X1   g0063(.A(n2190), .B(g74), .C(g77), .D(g71), .Y(n2191));
NOR4X1   g0135(.A(g83), .B(g52), .C(n2239), .D(g86), .Y(n2263));
NOR4X1   g0165(.A(n2190), .B(n2247_1), .C(g77), .D(n2232), .Y(n2293_1));
NOR4X1   g0105(.A(g68), .B(g74), .C(g77), .D(n2232), .Y(n2233_1));
AOI21X1  g0151(.A0(n2252), .A1(n2278_1), .B0(n2240), .Y(n2279));
AOI21X1  g0153(.A0(n2280), .A1(n2250), .B0(n2240), .Y(n2281));
AOI21X1  g0156(.A0(n2283_1), .A1(n2282), .B0(n2240), .Y(n2284));
OR4X1    g0185(.A(n2311), .B(n2310), .C(n2309), .D(n2312_1), .Y(n2313));
NOR3X1   g0162(.A(n2240), .B(n2289), .C(n2238), .Y(n2290));
NOR3X1   g0176(.A(n2303), .B(n2240), .C(n2238), .Y(n2304));
OR4X1    g0178(.A(n2299), .B(n2288_1), .C(n2287), .D(n2300), .Y(n2306));
OR2X1    g0179(.A(n2306), .B(n2305), .Y(n2307_1));
NOR4X1   g0168(.A(n2290), .B(n2288_1), .C(n2287), .D(n2295), .Y(n2296));
NAND2X1  g0314(.A(n2443), .B(n2442_1), .Y(n2444));
NOR3X1   g0183(.A(n2252), .B(n2240), .C(n2238), .Y(n2311));
NOR3X1   g0181(.A(n2280), .B(n2240), .C(n2238), .Y(n2309));
NOR3X1   g0123(.A(n2250), .B(n2238), .C(n2188), .Y(n2251_1));
NOR3X1   g0118(.A(n2238), .B(n2206), .C(n2188), .Y(n2246));
OR4X1    g0126(.A(n2251_1), .B(n2249), .C(n2246), .D(n2253), .Y(n2254));
NAND3X1  g0109(.A(n2236), .B(n2234), .C(n2231), .Y(n2237_1));
NOR3X1   g0115(.A(n2242_1), .B(n2240), .C(n2238), .Y(n2243));
NOR3X1   g0117(.A(n2244), .B(n2240), .C(n2238), .Y(n2245));
NAND2X1  g0307(.A(n2436), .B(n2435), .Y(n2437_1));
NOR3X1   g0125(.A(n2252), .B(n2238), .C(n2188), .Y(n2253));
NOR3X1   g0258(.A(n2278_1), .B(n2238), .C(n2188), .Y(n2386));
NOR3X1   g0218(.A(n2334), .B(n2242_1), .C(n2238), .Y(n2346));
NOR3X1   g0219(.A(n2334), .B(n2244), .C(n2238), .Y(n2347_1));
NOR2X1   g0220(.A(n2335), .B(n2238), .Y(n2348));
NOR3X1   g0226(.A(n2334), .B(n2273_1), .C(n2238), .Y(n2354));
NOR3X1   g0223(.A(n2334), .B(n2289), .C(n2238), .Y(n2351));
NOR3X1   g0224(.A(n2334), .B(n2298), .C(n2238), .Y(n2352_1));
NOR3X1   g0225(.A(n2334), .B(n2303), .C(n2238), .Y(n2353));
NOR3X1   g0231(.A(n2334), .B(n2238), .C(n2206), .Y(n2359));
NOR3X1   g0228(.A(n2334), .B(n2278_1), .C(n2238), .Y(n2356));
NOR3X1   g0229(.A(n2334), .B(n2252), .C(n2238), .Y(n2357_1));
NOR3X1   g0230(.A(n2334), .B(n2238), .C(n2248), .Y(n2358));
INVX1    g0104(.A(g71), .Y(n2232));
INVX1    g0101(.A(g77), .Y(n2229));
INVX1    g0119(.A(g74), .Y(n2247_1));
OR2X1    g0099(.A(g55), .B(g42), .Y(n2227));
INVX1    g0098(.A(g44), .Y(n2226));
INVX1    g0111(.A(g80), .Y(n2239));
NAND4X1  g0155(.A(n2190), .B(g74), .C(n2229), .D(n2232), .Y(n2283_1));
NAND4X1  g0152(.A(g68), .B(g74), .C(n2229), .D(n2232), .Y(n2280));
NAND4X1  g0154(.A(g68), .B(g74), .C(n2229), .D(g71), .Y(n2282));
NOR4X1   g0100(.A(n2226), .B(g45), .C(g41), .D(n2227), .Y(n1899));
AND2X1   g0113(.A(g74), .B(g77), .Y(n2241));
INVX1    g0062(.A(g68), .Y(n2190));
NAND4X1  g0145(.A(n2190), .B(n2247_1), .C(g77), .D(g71), .Y(n2273_1));
NAND4X1  g0150(.A(n2190), .B(n2247_1), .C(n2229), .D(g71), .Y(n2278_1));
NAND4X1  g0124(.A(g68), .B(n2247_1), .C(n2229), .D(g71), .Y(n2252));
NOR3X1   g0184(.A(n2240), .B(n2278_1), .C(n2238), .Y(n2312_1));
NOR3X1   g0182(.A(n2283_1), .B(n2240), .C(n2238), .Y(n2310));
NAND4X1  g0161(.A(n2190), .B(n2247_1), .C(g77), .D(n2232), .Y(n2289));
NAND4X1  g0175(.A(g68), .B(n2247_1), .C(g77), .D(g71), .Y(n2303));
NOR3X1   g0172(.A(n2282), .B(n2240), .C(n2238), .Y(n2300));
NOR3X1   g0159(.A(n2273_1), .B(n2240), .C(n2238), .Y(n2287));
NOR3X1   g0160(.A(n2250), .B(n2240), .C(n2238), .Y(n2288_1));
NOR3X1   g0171(.A(n2240), .B(n2298), .C(n2238), .Y(n2299));
OR2X1    g0177(.A(n2304), .B(n2290), .Y(n2305));
NAND3X1  g0167(.A(n2294), .B(n2292), .C(n2291), .Y(n2295));
NAND4X1  g0312(.A(n2263), .B(n1899), .C(g846), .D(n2276), .Y(n2442_1));
AOI22X1  g0313(.A0(n2299), .A1(g2), .B0(g863), .B1(n2300), .Y(n2443));
NAND4X1  g0060(.A(g83), .B(g52), .C(g80), .D(g86), .Y(n2188));
NOR3X1   g0121(.A(n2238), .B(n2248), .C(n2188), .Y(n2249));
NAND3X1  g0103(.A(n2230), .B(n1899), .C(n2189_1), .Y(n2231));
NAND3X1  g0106(.A(n2233_1), .B(n1899), .C(n2189_1), .Y(n2234));
NAND3X1  g0108(.A(n2235), .B(n1899), .C(n2189_1), .Y(n2236));
NAND3X1  g0114(.A(n2241), .B(n2232), .C(n2190), .Y(n2242_1));
NAND3X1  g0116(.A(n2241), .B(n2232), .C(g68), .Y(n2244));
NAND4X1  g0305(.A(n2191), .B(n2189_1), .C(g652), .D(n1899), .Y(n2435));
NAND4X1  g0306(.A(n2263), .B(n1899), .C(g513), .D(n2266_1), .Y(n2436));
NAND4X1  g0170(.A(g68), .B(n2247_1), .C(g77), .D(n2232), .Y(n2298));
NAND3X1  g0163(.A(n2276), .B(n2263), .C(n1899), .Y(n2291));
NAND3X1  g0164(.A(n2263), .B(n2230), .C(n1899), .Y(n2292));
NAND3X1  g0166(.A(n2293_1), .B(n2263), .C(n1899), .Y(n2294));
INVX1    g0061(.A(n2188), .Y(n2189_1));

endmodule
