//Converted to Combinational (Partial output: n901) , Module name: s9234_n901 , Timestamp: 2018-12-03T15:51:03.518331 
module s9234_n901 ( g314, g301, g306, g310, g54, g319, g79, g84, g374, g323, g332, g361, g49, g345, g349, g338, g341, g357, g353, g59, g69, g74, g64, n901 );
input g314, g301, g306, g310, g54, g319, g79, g84, g374, g323, g332, g361, g49, g345, g349, g338, g341, g357, g353, g59, g69, g74, g64;
output n901;
wire n1055, n1051_1, n1655, n1054, n755, n1050, n1026_1, n1654, n1649, n1034, n1053, n1022, n1046_1, n1049, n1025, n1653, n1016_1, n1052, n1014, n1018, n1021_1, n1033, n1045, n1048, n1013, n1047, n1037, n1024, n1652, n1478, n751_1, n1017, n1015, n1019, n1020, n1032, n1036_1, n1035, n1039, n1023, n1650, n1651, n750, n748, n749, n1031_1, n1028, n1029, n1030, n1038;
OAI21X1  g0946(.A0(n1655), .A1(n1051_1), .B0(n1055), .Y(n901));
OAI21X1  g0346(.A0(n1050), .A1(n755), .B0(n1054), .Y(n1055));
OR2X1    g0342(.A(n1050), .B(n755), .Y(n1051_1));
MX2X1    g0945(.A(n1649), .B(n1654), .S0(n1026_1), .Y(n1655));
NOR3X1   g0345(.A(n1053), .B(n755), .C(n1034), .Y(n1054));
NOR4X1   g0047(.A(g310), .B(g306), .C(g301), .D(g314), .Y(n755));
AOI21X1  g0341(.A0(n1049), .A1(n1046_1), .B0(n1022), .Y(n1050));
NAND2X1  g0317(.A(n1025), .B(n1022), .Y(n1026_1));
XOR2X1   g0944(.A(n1653), .B(g54), .Y(n1654));
INVX1    g0939(.A(g54), .Y(n1649));
NOR3X1   g0325(.A(g314), .B(n1016_1), .C(g306), .Y(n1034));
INVX1    g0344(.A(n1052), .Y(n1053));
OAI21X1  g0313(.A0(n1021_1), .A1(n1018), .B0(n1014), .Y(n1022));
OR2X1    g0337(.A(n1045), .B(n1033), .Y(n1046_1));
OR4X1    g0340(.A(n1037), .B(n1047), .C(n1013), .D(n1048), .Y(n1049));
OAI21X1  g0316(.A0(n1024), .A1(g319), .B0(n1014), .Y(n1025));
MX2X1    g0943(.A(n1478), .B(n1652), .S0(n1025), .Y(n1653));
INVX1    g0307(.A(g310), .Y(n1016_1));
AOI21X1  g0343(.A0(n1016_1), .A1(g306), .B0(n1021_1), .Y(n1052));
INVX1    g0305(.A(n751_1), .Y(n1014));
AOI21X1  g0309(.A0(n1016_1), .A1(n1015), .B0(n1017), .Y(n1018));
NOR3X1   g0312(.A(g319), .B(n1020), .C(n1019), .Y(n1021_1));
OR2X1    g0324(.A(n1032), .B(g79), .Y(n1033));
OR4X1    g0336(.A(n1035), .B(n1034), .C(g84), .D(n1036_1), .Y(n1045));
INVX1    g0339(.A(n1039), .Y(n1048));
INVX1    g0304(.A(g84), .Y(n1013));
INVX1    g0338(.A(g79), .Y(n1047));
NOR3X1   g0328(.A(n1036_1), .B(n1035), .C(n1034), .Y(n1037));
NOR4X1   g0315(.A(g319), .B(n1020), .C(g306), .D(n1023), .Y(n1024));
MX2X1    g0942(.A(n1651), .B(n1650), .S0(n1037), .Y(n1652));
INVX1    g0768(.A(g374), .Y(n1478));
NAND4X1  g0043(.A(n749), .B(n748), .C(g323), .D(n750), .Y(n751_1));
INVX1    g0308(.A(g332), .Y(n1017));
INVX1    g0306(.A(g306), .Y(n1015));
INVX1    g0310(.A(g301), .Y(n1019));
INVX1    g0311(.A(g314), .Y(n1020));
NAND4X1  g0323(.A(n1030), .B(n1029), .C(n1028), .D(n1031_1), .Y(n1032));
NOR3X1   g0327(.A(g314), .B(g310), .C(n1015), .Y(n1036_1));
NOR2X1   g0326(.A(n1020), .B(g306), .Y(n1035));
NOR4X1   g0330(.A(n1030), .B(n1029), .C(n1028), .D(n1038), .Y(n1039));
OR2X1    g0314(.A(g310), .B(g301), .Y(n1023));
OR2X1    g0940(.A(g49), .B(g361), .Y(n1650));
NAND2X1  g0941(.A(g49), .B(g361), .Y(n1651));
NOR4X1   g0042(.A(g341), .B(g338), .C(g349), .D(g345), .Y(n750));
INVX1    g0040(.A(g357), .Y(n748));
INVX1    g0041(.A(g353), .Y(n749));
NOR4X1   g0322(.A(g49), .B(g54), .C(g361), .D(g59), .Y(n1031_1));
INVX1    g0319(.A(g69), .Y(n1028));
INVX1    g0320(.A(g74), .Y(n1029));
INVX1    g0321(.A(g64), .Y(n1030));
NAND4X1  g0329(.A(g49), .B(g54), .C(g361), .D(g59), .Y(n1038));

endmodule
