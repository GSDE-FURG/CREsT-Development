//Converted to Combinational (Partial output: n117) , Module name: s1238_n117
module s1238_n117 ( G1, G3, G4, G10, G34, G13, G7, G9, G6, G8, G12, G11, G46, G5, G31, G0, G2, G30, n117 );
input G1, G3, G4, G10, G34, G13, G7, G9, G6, G8, G12, G11, G46, G5, G31, G0, G2, G30;
output n117;
wire n394, n214, n216, n393, n120, n392, n101, n104, n130, n100, n215, n105, n223, n119, n82_1, n97_1, n125, n387, n118, n98, n111, n115, n84, n86, n96, n117_1, n99, n107_1, n110, n103, n113, n114, n83, n85, n87_1, n88, n95, n116, n106, n108, n109, n102_1, n112_1, n94, n90, n89, n93, n92_1, n91;
AOI21X1  g313(.A0(n216), .A1(n214), .B0(n394), .Y(n117));
OAI21X1  g312(.A0(n392), .A1(n120), .B0(n393), .Y(n394));
NOR3X1   g132(.A(G10), .B(n104), .C(n101), .Y(n214));
OAI22X1  g134(.A0(n215), .A1(n100), .B0(n130), .B1(n120), .Y(n216));
NAND3X1  g311(.A(n223), .B(n105), .C(G34), .Y(n393));
OR4X1    g038(.A(n97_1), .B(G13), .C(n82_1), .D(n119), .Y(n120));
OR2X1    g310(.A(n387), .B(n125), .Y(n392));
INVX1    g019(.A(G7), .Y(n101));
INVX1    g022(.A(G9), .Y(n104));
INVX1    g048(.A(G6), .Y(n130));
INVX1    g018(.A(G8), .Y(n100));
INVX1    g133(.A(G34), .Y(n215));
AND2X1   g023(.A(G10), .B(G8), .Y(n105));
NAND2X1  g141(.A(G9), .B(G7), .Y(n223));
OR4X1    g037(.A(n115), .B(n111), .C(n98), .D(n118), .Y(n119));
INVX1    g000(.A(G12), .Y(n82_1));
AOI21X1  g015(.A0(n96), .A1(n86), .B0(n84), .Y(n97_1));
NAND2X1  g043(.A(G10), .B(G7), .Y(n125));
AND2X1   g305(.A(G9), .B(G6), .Y(n387));
NOR4X1   g036(.A(G11), .B(n104), .C(G7), .D(n117_1), .Y(n118));
INVX1    g016(.A(G46), .Y(n98));
AOI21X1  g029(.A0(n110), .A1(n107_1), .B0(n99), .Y(n111));
NOR3X1   g033(.A(n114), .B(n113), .C(n103), .Y(n115));
NOR2X1   g002(.A(G5), .B(n83), .Y(n84));
NAND3X1  g004(.A(n83), .B(G3), .C(n85), .Y(n86));
OAI21X1  g014(.A0(n95), .A1(n88), .B0(n87_1), .Y(n96));
MX2X1    g035(.A(n116), .B(G31), .S0(G8), .Y(n117_1));
INVX1    g017(.A(G11), .Y(n99));
OR4X1    g025(.A(n103), .B(G31), .C(n100), .D(n106), .Y(n107_1));
NOR2X1   g028(.A(n109), .B(n108), .Y(n110));
NOR3X1   g021(.A(n102_1), .B(n101), .C(G6), .Y(n103));
NAND2X1  g031(.A(n112_1), .B(n104), .Y(n113));
AND2X1   g032(.A(G31), .B(G8), .Y(n114));
INVX1    g001(.A(G4), .Y(n83));
INVX1    g003(.A(G0), .Y(n85));
INVX1    g005(.A(G5), .Y(n87_1));
NOR3X1   g006(.A(G3), .B(G2), .C(n85), .Y(n88));
AOI21X1  g013(.A0(n94), .A1(G0), .B0(G4), .Y(n95));
INVX1    g034(.A(G10), .Y(n116));
NOR2X1   g024(.A(n105), .B(n104), .Y(n106));
NOR3X1   g026(.A(G9), .B(G8), .C(G7), .Y(n108));
NOR2X1   g027(.A(G30), .B(G6), .Y(n109));
INVX1    g020(.A(G30), .Y(n102_1));
NOR2X1   g030(.A(G11), .B(G10), .Y(n112_1));
OAI21X1  g012(.A0(n93), .A1(n89), .B0(n90), .Y(n94));
INVX1    g008(.A(G3), .Y(n90));
INVX1    g007(.A(G2), .Y(n89));
AOI22X1  g011(.A0(G5), .A1(n91), .B0(G4), .B1(n92_1), .Y(n93));
NAND2X1  g010(.A(G5), .B(G3), .Y(n92_1));
INVX1    g009(.A(G1), .Y(n91));

endmodule
