//Converted to Combinational (Partial output: n1243) , Module name: s38584_n1243 , Timestamp: 2018-12-03T15:51:16.137127 
module s38584_n1243 ( g35, g671, g703, g676, g504, g499, g650, g661, g728, g718, g655, g645, g528, g681, g699, g490, g482, g385, g358, g370, g376, n1243 );
input g35, g671, g703, g676, g504, g499, g650, g661, g728, g718, g655, g645, g528, g681, g699, g490, g482, g385, g358, g370, g376;
output n1243;
wire n6243, n6238, n6240, n6242, n6237, n6239, n6241_1, n6236_1, n6233, n5879, n6234, n6235, n6232, n6227, n6228, n6230, n5878, n5688, n6231_1, n6229, n5132, n5130_1, n5600, n5598, n5687, n5599;
MX2X1    g1604(.A(g671), .B(n6243), .S0(g35), .Y(n1243));
AOI21X1  g1603(.A0(n6242), .A1(n6240), .B0(n6238), .Y(n6243));
NAND2X1  g1598(.A(n6237), .B(g703), .Y(n6238));
NAND2X1  g1600(.A(n6239), .B(g676), .Y(n6240));
NAND3X1  g1602(.A(n6236_1), .B(g671), .C(n6241_1), .Y(n6242));
NAND2X1  g1597(.A(n6236_1), .B(n6233), .Y(n6237));
NAND2X1  g1599(.A(n6236_1), .B(g671), .Y(n6239));
INVX1    g1601(.A(g676), .Y(n6241_1));
NOR4X1   g1596(.A(n6235), .B(n6234), .C(g504), .D(n5879), .Y(n6236_1));
NOR4X1   g1593(.A(n6230), .B(n6228), .C(n6227), .D(n6232), .Y(n6233));
INVX1    g1239(.A(n5878), .Y(n5879));
INVX1    g1594(.A(g499), .Y(n6234));
INVX1    g1595(.A(n5688), .Y(n6235));
OR2X1    g1592(.A(g650), .B(n6231_1), .Y(n6232));
XOR2X1   g1587(.A(g728), .B(g661), .Y(n6227));
XOR2X1   g1588(.A(g655), .B(g718), .Y(n6228));
OR2X1    g1590(.A(n6229), .B(g645), .Y(n6230));
NOR3X1   g1238(.A(n5130_1), .B(g528), .C(n5132), .Y(n5878));
NOR4X1   g1048(.A(n5599), .B(n5687), .C(n5598), .D(n5600), .Y(n5688));
INVX1    g1591(.A(g681), .Y(n6231_1));
INVX1    g1589(.A(g699), .Y(n6229));
INVX1    g0500(.A(g490), .Y(n5132));
INVX1    g0498(.A(g482), .Y(n5130_1));
INVX1    g0960(.A(g385), .Y(n5600));
INVX1    g0958(.A(g358), .Y(n5598));
INVX1    g1047(.A(g370), .Y(n5687));
INVX1    g0959(.A(g376), .Y(n5599));

endmodule
