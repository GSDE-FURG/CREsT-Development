//Converted to Combinational (Partial output: n65) , Module name: s1488_n65 , Timestamp: 2018-12-03T15:51:02.598893 
module s1488_n65 ( v1, CLR, v7, v11, v10, v12, v9, v8, v3, v6, v0, v5, v4, v2, n65 );
input v1, CLR, v7, v11, v10, v12, v9, v8, v3, v6, v0, v5, v4, v2;
output n65;
wire n267, n333, n336, n45, n323, n332, n335, n217, n203, n232, n72, n319, n322, n331, n326, n334, n219, n63, n318, n320, n321, n330, n247, n327, n329, n325, n86, n83, n324, n154, n48, n61, n317, n295, n47, n90, n74, n103, n82, n328, n142, n50, n68, n54, n259, n104;
AOI21X1  g292(.A0(n336), .A1(n333), .B0(n267), .Y(n65));
INVX1    g222(.A(CLR), .Y(n267));
OAI21X1  g288(.A0(n332), .A1(n323), .B0(n45), .Y(n333));
AOI22X1  g291(.A0(n232), .A1(n203), .B0(n217), .B1(n335), .Y(n336));
INVX1    g000(.A(v7), .Y(n45));
AOI21X1  g278(.A0(n322), .A1(n319), .B0(n72), .Y(n323));
OAI21X1  g287(.A0(n326), .A1(v11), .B0(n331), .Y(n332));
OAI21X1  g290(.A0(n219), .A1(v10), .B0(n334), .Y(n335));
NOR2X1   g172(.A(n72), .B(v11), .Y(n217));
NOR2X1   g158(.A(n45), .B(v12), .Y(n203));
AND2X1   g187(.A(v9), .B(v11), .Y(n232));
INVX1    g027(.A(v8), .Y(n72));
OR2X1    g274(.A(n318), .B(n63), .Y(n319));
AOI21X1  g277(.A0(n321), .A1(n63), .B0(n320), .Y(n322));
AOI22X1  g286(.A0(n329), .A1(n327), .B0(n247), .B1(n330), .Y(n331));
AOI22X1  g281(.A0(n324), .A1(n83), .B0(n86), .B1(n325), .Y(n326));
NAND3X1  g289(.A(n63), .B(v10), .C(v12), .Y(n334));
INVX1    g174(.A(n154), .Y(n219));
INVX1    g018(.A(v9), .Y(n63));
AOI22X1  g273(.A0(n295), .A1(n317), .B0(n61), .B1(n48), .Y(n318));
AOI21X1  g275(.A0(n90), .A1(n47), .B0(v10), .Y(n320));
OAI21X1  g276(.A0(n247), .A1(v11), .B0(v10), .Y(n321));
MX2X1    g285(.A(v8), .B(n74), .S0(v10), .Y(n330));
NOR2X1   g202(.A(v12), .B(n103), .Y(n247));
NOR2X1   g282(.A(v8), .B(n82), .Y(n327));
OAI22X1  g284(.A0(n142), .A1(v9), .B0(v10), .B1(n328), .Y(n329));
MX2X1    g280(.A(n68), .B(n50), .S0(n82), .Y(n325));
INVX1    g041(.A(v3), .Y(n86));
NOR2X1   g038(.A(v9), .B(v10), .Y(n83));
NOR2X1   g279(.A(n54), .B(v12), .Y(n324));
NAND2X1  g109(.A(n63), .B(v12), .Y(n154));
INVX1    g003(.A(v6), .Y(n48));
NOR2X1   g016(.A(v11), .B(v12), .Y(n61));
NOR2X1   g272(.A(n47), .B(n86), .Y(n317));
NAND3X1  g250(.A(v0), .B(n259), .C(v6), .Y(n295));
NAND2X1  g002(.A(v11), .B(v12), .Y(n47));
AND2X1   g045(.A(v4), .B(v5), .Y(n90));
NOR2X1   g029(.A(v8), .B(n63), .Y(n74));
INVX1    g058(.A(v2), .Y(n103));
INVX1    g037(.A(v12), .Y(n82));
AOI21X1  g283(.A0(n104), .A1(v6), .B0(v9), .Y(n328));
NAND2X1  g097(.A(v10), .B(v11), .Y(n142));
AND2X1   g005(.A(v8), .B(v9), .Y(n50));
INVX1    g023(.A(v10), .Y(n68));
NAND2X1  g009(.A(v4), .B(v5), .Y(n54));
INVX1    g214(.A(v1), .Y(n259));
INVX1    g059(.A(v11), .Y(n104));

endmodule
