//Converted to Combinational (Partial output: n4583) , Module name: s35932_n4583 , Timestamp: 2018-12-03T15:51:09.384768 
module s35932_n4583 ( RESET, TM1, TM0, WX5657, WX5881, WX6009, WX7174, WX7302, WX5817, WX5945, WX7110, WX7238, WX6011, WX6013, WX6015, WX6017, WX6019, WX6021, WX6023, WX6025, WX6027, WX6029, WX6031, WX6033, WX6035, WX6037, WX6039, WX6041, WX6043, WX6045, WX6047, WX6049, WX6051, WX6053, WX6055, WX6057, WX6059, WX6061, WX6063, WX6065, WX6067, WX6069, WX6071, n4583 );
input RESET, TM1, TM0, WX5657, WX5881, WX6009, WX7174, WX7302, WX5817, WX5945, WX7110, WX7238, WX6011, WX6013, WX6015, WX6017, WX6019, WX6021, WX6023, WX6025, WX6027, WX6029, WX6031, WX6033, WX6035, WX6037, WX6039, WX6041, WX6043, WX6045, WX6047, WX6049, WX6051, WX6053, WX6055, WX6057, WX6059, WX6061, WX6063, WX6065, WX6067, WX6069, WX6071;
output n4583;
wire n5827, n8155_1, n8154, n8152, n5539, n7571, n8153, n8150_1, n8145_1, n7568, n7570, n8147, n8149, CRC_OUT_5_31, n7567_1, n7569, n8146, n8148, n8690_1, CRC_OUT_5_30, n8688, CRC_OUT_5_29, n8686, CRC_OUT_5_28, n8684, CRC_OUT_5_27, n8682, CRC_OUT_5_26, n8680_1, CRC_OUT_5_25, n8678, CRC_OUT_5_24, n8676, CRC_OUT_5_23, n8674, CRC_OUT_5_22, n8672, CRC_OUT_5_21, n8670_1, CRC_OUT_5_20, n8668, CRC_OUT_5_19, n8666, CRC_OUT_5_18, n8664, CRC_OUT_5_17, n8662, CRC_OUT_5_16, n8660_1, CRC_OUT_5_15, n8659, n8657, CRC_OUT_5_14, n8655_1, CRC_OUT_5_13, n8653, CRC_OUT_5_12, n8651, CRC_OUT_5_11, n8649, CRC_OUT_5_10, n8648, n8646, CRC_OUT_5_9, n8644, CRC_OUT_5_8, n8642, CRC_OUT_5_7, n8640_1, CRC_OUT_5_6, n8638, CRC_OUT_5_5, n8636, CRC_OUT_5_4, n8634, CRC_OUT_5_3, n8633, n8631, CRC_OUT_5_2, n8629, CRC_OUT_5_1, n8627, CRC_OUT_5_0, n8625_1;
NOR2X1   g2488(.A(n8155_1), .B(n5827), .Y(n4583));
INVX1    g0288(.A(RESET), .Y(n5827));
MX2X1    g2487(.A(n8152), .B(n8154), .S0(TM1), .Y(n8155_1));
MX2X1    g2486(.A(n8153), .B(n7571), .S0(n5539), .Y(n8154));
MX2X1    g2484(.A(n8145_1), .B(n8150_1), .S0(n5539), .Y(n8152));
INVX1    g0000(.A(TM0), .Y(n5539));
XOR2X1   g1936(.A(n7570), .B(n7568), .Y(n7571));
INVX1    g2485(.A(WX5657), .Y(n8153));
XOR2X1   g2483(.A(n8149), .B(n8147), .Y(n8150_1));
INVX1    g2478(.A(CRC_OUT_5_31), .Y(n8145_1));
XOR2X1   g1933(.A(n7567_1), .B(WX5881), .Y(n7568));
XOR2X1   g1935(.A(WX6009), .B(n7569), .Y(n7570));
XOR2X1   g2480(.A(n8146), .B(WX7174), .Y(n8147));
XOR2X1   g2482(.A(WX7302), .B(n8148), .Y(n8149));
NOR2X1   g2992(.A(n8690_1), .B(n5827), .Y(CRC_OUT_5_31));
XOR2X1   g1932(.A(WX5817), .B(TM1), .Y(n7567_1));
INVX1    g1934(.A(WX5945), .Y(n7569));
XOR2X1   g2479(.A(WX7110), .B(TM1), .Y(n8146));
INVX1    g2481(.A(WX7238), .Y(n8148));
XOR2X1   g2991(.A(CRC_OUT_5_30), .B(WX6009), .Y(n8690_1));
NOR2X1   g2990(.A(n8688), .B(n5827), .Y(CRC_OUT_5_30));
XOR2X1   g2989(.A(CRC_OUT_5_29), .B(WX6011), .Y(n8688));
NOR2X1   g2988(.A(n8686), .B(n5827), .Y(CRC_OUT_5_29));
XOR2X1   g2987(.A(CRC_OUT_5_28), .B(WX6013), .Y(n8686));
NOR2X1   g2986(.A(n8684), .B(n5827), .Y(CRC_OUT_5_28));
XOR2X1   g2985(.A(CRC_OUT_5_27), .B(WX6015), .Y(n8684));
NOR2X1   g2984(.A(n8682), .B(n5827), .Y(CRC_OUT_5_27));
XOR2X1   g2983(.A(CRC_OUT_5_26), .B(WX6017), .Y(n8682));
NOR2X1   g2982(.A(n8680_1), .B(n5827), .Y(CRC_OUT_5_26));
XOR2X1   g2981(.A(CRC_OUT_5_25), .B(WX6019), .Y(n8680_1));
NOR2X1   g2980(.A(n8678), .B(n5827), .Y(CRC_OUT_5_25));
XOR2X1   g2979(.A(CRC_OUT_5_24), .B(WX6021), .Y(n8678));
NOR2X1   g2978(.A(n8676), .B(n5827), .Y(CRC_OUT_5_24));
XOR2X1   g2977(.A(CRC_OUT_5_23), .B(WX6023), .Y(n8676));
NOR2X1   g2976(.A(n8674), .B(n5827), .Y(CRC_OUT_5_23));
XOR2X1   g2975(.A(CRC_OUT_5_22), .B(WX6025), .Y(n8674));
NOR2X1   g2974(.A(n8672), .B(n5827), .Y(CRC_OUT_5_22));
XOR2X1   g2973(.A(CRC_OUT_5_21), .B(WX6027), .Y(n8672));
NOR2X1   g2972(.A(n8670_1), .B(n5827), .Y(CRC_OUT_5_21));
XOR2X1   g2971(.A(CRC_OUT_5_20), .B(WX6029), .Y(n8670_1));
NOR2X1   g2970(.A(n8668), .B(n5827), .Y(CRC_OUT_5_20));
XOR2X1   g2969(.A(CRC_OUT_5_19), .B(WX6031), .Y(n8668));
NOR2X1   g2968(.A(n8666), .B(n5827), .Y(CRC_OUT_5_19));
XOR2X1   g2967(.A(CRC_OUT_5_18), .B(WX6033), .Y(n8666));
NOR2X1   g2966(.A(n8664), .B(n5827), .Y(CRC_OUT_5_18));
XOR2X1   g2965(.A(CRC_OUT_5_17), .B(WX6035), .Y(n8664));
NOR2X1   g2964(.A(n8662), .B(n5827), .Y(CRC_OUT_5_17));
XOR2X1   g2963(.A(CRC_OUT_5_16), .B(WX6037), .Y(n8662));
NOR2X1   g2962(.A(n8660_1), .B(n5827), .Y(CRC_OUT_5_16));
XOR2X1   g2961(.A(n8659), .B(CRC_OUT_5_15), .Y(n8660_1));
NOR2X1   g2959(.A(n8657), .B(n5827), .Y(CRC_OUT_5_15));
XOR2X1   g2960(.A(CRC_OUT_5_31), .B(WX6039), .Y(n8659));
XOR2X1   g2958(.A(CRC_OUT_5_14), .B(WX6041), .Y(n8657));
NOR2X1   g2957(.A(n8655_1), .B(n5827), .Y(CRC_OUT_5_14));
XOR2X1   g2956(.A(CRC_OUT_5_13), .B(WX6043), .Y(n8655_1));
NOR2X1   g2955(.A(n8653), .B(n5827), .Y(CRC_OUT_5_13));
XOR2X1   g2954(.A(CRC_OUT_5_12), .B(WX6045), .Y(n8653));
NOR2X1   g2953(.A(n8651), .B(n5827), .Y(CRC_OUT_5_12));
XOR2X1   g2952(.A(CRC_OUT_5_11), .B(WX6047), .Y(n8651));
NOR2X1   g2951(.A(n8649), .B(n5827), .Y(CRC_OUT_5_11));
XOR2X1   g2950(.A(n8648), .B(CRC_OUT_5_10), .Y(n8649));
NOR2X1   g2948(.A(n8646), .B(n5827), .Y(CRC_OUT_5_10));
XOR2X1   g2949(.A(CRC_OUT_5_31), .B(WX6049), .Y(n8648));
XOR2X1   g2947(.A(CRC_OUT_5_9), .B(WX6051), .Y(n8646));
NOR2X1   g2946(.A(n8644), .B(n5827), .Y(CRC_OUT_5_9));
XOR2X1   g2945(.A(CRC_OUT_5_8), .B(WX6053), .Y(n8644));
NOR2X1   g2944(.A(n8642), .B(n5827), .Y(CRC_OUT_5_8));
XOR2X1   g2943(.A(CRC_OUT_5_7), .B(WX6055), .Y(n8642));
NOR2X1   g2942(.A(n8640_1), .B(n5827), .Y(CRC_OUT_5_7));
XOR2X1   g2941(.A(CRC_OUT_5_6), .B(WX6057), .Y(n8640_1));
NOR2X1   g2940(.A(n8638), .B(n5827), .Y(CRC_OUT_5_6));
XOR2X1   g2939(.A(CRC_OUT_5_5), .B(WX6059), .Y(n8638));
NOR2X1   g2938(.A(n8636), .B(n5827), .Y(CRC_OUT_5_5));
XOR2X1   g2937(.A(CRC_OUT_5_4), .B(WX6061), .Y(n8636));
NOR2X1   g2936(.A(n8634), .B(n5827), .Y(CRC_OUT_5_4));
XOR2X1   g2935(.A(n8633), .B(CRC_OUT_5_3), .Y(n8634));
NOR2X1   g2933(.A(n8631), .B(n5827), .Y(CRC_OUT_5_3));
XOR2X1   g2934(.A(CRC_OUT_5_31), .B(WX6063), .Y(n8633));
XOR2X1   g2932(.A(CRC_OUT_5_2), .B(WX6065), .Y(n8631));
NOR2X1   g2931(.A(n8629), .B(n5827), .Y(CRC_OUT_5_2));
XOR2X1   g2930(.A(CRC_OUT_5_1), .B(WX6067), .Y(n8629));
NOR2X1   g2929(.A(n8627), .B(n5827), .Y(CRC_OUT_5_1));
XOR2X1   g2928(.A(CRC_OUT_5_0), .B(WX6069), .Y(n8627));
NOR2X1   g2927(.A(n8625_1), .B(n5827), .Y(CRC_OUT_5_0));
XOR2X1   g2926(.A(CRC_OUT_5_31), .B(WX6071), .Y(n8625_1));

endmodule
