// Benchmark "b13_C" written by ABC on Wed Aug 05 14:40:28 2020

module b13_C ( 
    EOC, DATA_OUT_REG_SCAN_IN, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_,
    DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_, DSR,
    TX_END_REG_SCAN_IN, S2_REG_0__SCAN_IN, S2_REG_1__SCAN_IN,
    CANALE_REG_3__SCAN_IN, CANALE_REG_2__SCAN_IN, CANALE_REG_1__SCAN_IN,
    CANALE_REG_0__SCAN_IN, CONTA_TMP_REG_3__SCAN_IN,
    CONTA_TMP_REG_2__SCAN_IN, CONTA_TMP_REG_1__SCAN_IN,
    CONTA_TMP_REG_0__SCAN_IN, ITFC_STATE_REG_1__SCAN_IN,
    ITFC_STATE_REG_0__SCAN_IN, OUT_REG_REG_7__SCAN_IN,
    OUT_REG_REG_6__SCAN_IN, OUT_REG_REG_5__SCAN_IN, OUT_REG_REG_4__SCAN_IN,
    OUT_REG_REG_3__SCAN_IN, OUT_REG_REG_2__SCAN_IN, OUT_REG_REG_1__SCAN_IN,
    OUT_REG_REG_0__SCAN_IN, NEXT_BIT_REG_3__SCAN_IN,
    NEXT_BIT_REG_2__SCAN_IN, NEXT_BIT_REG_1__SCAN_IN,
    NEXT_BIT_REG_0__SCAN_IN, TX_CONTA_REG_9__SCAN_IN,
    TX_CONTA_REG_8__SCAN_IN, TX_CONTA_REG_7__SCAN_IN,
    TX_CONTA_REG_6__SCAN_IN, TX_CONTA_REG_5__SCAN_IN,
    TX_CONTA_REG_4__SCAN_IN, TX_CONTA_REG_3__SCAN_IN,
    TX_CONTA_REG_2__SCAN_IN, TX_CONTA_REG_1__SCAN_IN,
    TX_CONTA_REG_0__SCAN_IN, LOAD_REG_SCAN_IN, SEND_DATA_REG_SCAN_IN,
    SEND_EN_REG_SCAN_IN, MUX_EN_REG_SCAN_IN, TRE_REG_SCAN_IN,
    LOAD_DATO_REG_SCAN_IN, SOC_REG_SCAN_IN, SEND_REG_SCAN_IN,
    MPX_REG_SCAN_IN, CONFIRM_REG_SCAN_IN, SHOT_REG_SCAN_IN,
    ADD_MPX2_REG_SCAN_IN, RDY_REG_SCAN_IN, ERROR_REG_SCAN_IN,
    S1_REG_2__SCAN_IN, S1_REG_1__SCAN_IN, S1_REG_0__SCAN_IN,
    U416, U415, U414, U413, U417, U412, U411, U410, U452, U409, U453, U454,
    U455, U456, U457, U458, U459, U460, U461, U408, U407, U462, U406, U405,
    U404, U403, U402, U401, U400, U399, U398, U397, U396, U395, U394, U393,
    U392, U391, U450, U390, U389, U388, U387, U386, U385, U451, U383, U464,
    U384, U463, U382, U381, U380  );
  input  EOC, DATA_OUT_REG_SCAN_IN, DATA_IN_7_, DATA_IN_6_, DATA_IN_5_,
    DATA_IN_4_, DATA_IN_3_, DATA_IN_2_, DATA_IN_1_, DATA_IN_0_, DSR,
    TX_END_REG_SCAN_IN, S2_REG_0__SCAN_IN, S2_REG_1__SCAN_IN,
    CANALE_REG_3__SCAN_IN, CANALE_REG_2__SCAN_IN, CANALE_REG_1__SCAN_IN,
    CANALE_REG_0__SCAN_IN, CONTA_TMP_REG_3__SCAN_IN,
    CONTA_TMP_REG_2__SCAN_IN, CONTA_TMP_REG_1__SCAN_IN,
    CONTA_TMP_REG_0__SCAN_IN, ITFC_STATE_REG_1__SCAN_IN,
    ITFC_STATE_REG_0__SCAN_IN, OUT_REG_REG_7__SCAN_IN,
    OUT_REG_REG_6__SCAN_IN, OUT_REG_REG_5__SCAN_IN, OUT_REG_REG_4__SCAN_IN,
    OUT_REG_REG_3__SCAN_IN, OUT_REG_REG_2__SCAN_IN, OUT_REG_REG_1__SCAN_IN,
    OUT_REG_REG_0__SCAN_IN, NEXT_BIT_REG_3__SCAN_IN,
    NEXT_BIT_REG_2__SCAN_IN, NEXT_BIT_REG_1__SCAN_IN,
    NEXT_BIT_REG_0__SCAN_IN, TX_CONTA_REG_9__SCAN_IN,
    TX_CONTA_REG_8__SCAN_IN, TX_CONTA_REG_7__SCAN_IN,
    TX_CONTA_REG_6__SCAN_IN, TX_CONTA_REG_5__SCAN_IN,
    TX_CONTA_REG_4__SCAN_IN, TX_CONTA_REG_3__SCAN_IN,
    TX_CONTA_REG_2__SCAN_IN, TX_CONTA_REG_1__SCAN_IN,
    TX_CONTA_REG_0__SCAN_IN, LOAD_REG_SCAN_IN, SEND_DATA_REG_SCAN_IN,
    SEND_EN_REG_SCAN_IN, MUX_EN_REG_SCAN_IN, TRE_REG_SCAN_IN,
    LOAD_DATO_REG_SCAN_IN, SOC_REG_SCAN_IN, SEND_REG_SCAN_IN,
    MPX_REG_SCAN_IN, CONFIRM_REG_SCAN_IN, SHOT_REG_SCAN_IN,
    ADD_MPX2_REG_SCAN_IN, RDY_REG_SCAN_IN, ERROR_REG_SCAN_IN,
    S1_REG_2__SCAN_IN, S1_REG_1__SCAN_IN, S1_REG_0__SCAN_IN;
  output U416, U415, U414, U413, U417, U412, U411, U410, U452, U409, U453,
    U454, U455, U456, U457, U458, U459, U460, U461, U408, U407, U462, U406,
    U405, U404, U403, U402, U401, U400, U399, U398, U397, U396, U395, U394,
    U393, U392, U391, U450, U390, U389, U388, U387, U386, U385, U451, U383,
    U464, U384, U463, U382, U381, U380;
  wire n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
    n137, n138, n140, n141, n143, n144, n145, n146, n148, n149, n151, n153,
    n155, n158, n159, n160, n162, n163, n164, n166, n167, n168, n169, n171,
    n172, n174, n175, n177, n178, n180, n181, n183, n184, n186, n187, n189,
    n190, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
    n203, n204, n205, n206, n207, n208, n210, n211, n212, n213, n214, n215,
    n217, n218, n219, n221, n222, n224, n225, n226, n227, n228, n230, n231,
    n233, n235, n236, n238, n239, n241, n243, n244, n246, n247, n248, n250,
    n251, n253, n255, n256, n257, n258, n260, n261, n262, n264, n266, n267,
    n268, n269, n272, n274, n276, n278, n279, n280, n282, n284, n285, n286,
    n288, n290, n291, n292, n294, n295, n296, n297, n300, n301, n303, n304,
    n306, n307, n310, n312, n313, n314, n315, n316, n317, n318, n319, n320,
    n321, n322, n323;
  INVX1   g000(.A(CONTA_TMP_REG_3__SCAN_IN), .Y(n126));
  INVX1   g001(.A(S1_REG_2__SCAN_IN), .Y(n127));
  INVX1   g002(.A(S1_REG_0__SCAN_IN), .Y(n128));
  NAND2X1 g003(.A(n128), .B(S1_REG_1__SCAN_IN), .Y(n129));
  OAI21X1 g004(.A0(n129), .A1(n127), .B0(CANALE_REG_3__SCAN_IN), .Y(n130));
  INVX1   g005(.A(S1_REG_1__SCAN_IN), .Y(n131));
  NOR3X1  g006(.A(S1_REG_0__SCAN_IN), .B(n131), .C(n127), .Y(n132));
  INVX1   g007(.A(n132), .Y(n133));
  INVX1   g008(.A(CONTA_TMP_REG_1__SCAN_IN), .Y(n134));
  INVX1   g009(.A(CONTA_TMP_REG_0__SCAN_IN), .Y(n135));
  NOR2X1  g010(.A(n135), .B(n134), .Y(n136));
  AOI21X1 g011(.A0(n136), .A1(CONTA_TMP_REG_2__SCAN_IN), .B0(n133), .Y(n137));
  INVX1   g012(.A(n137), .Y(n138));
  OAI21X1 g013(.A0(n138), .A1(n126), .B0(n130), .Y(U416));
  INVX1   g014(.A(CONTA_TMP_REG_2__SCAN_IN), .Y(n140));
  AOI22X1 g015(.A0(n136), .A1(n137), .B0(n133), .B1(CANALE_REG_2__SCAN_IN), .Y(n141));
  OAI21X1 g016(.A0(n138), .A1(n140), .B0(n141), .Y(U415));
  NAND3X1 g017(.A(CONTA_TMP_REG_0__SCAN_IN), .B(CONTA_TMP_REG_1__SCAN_IN), .C(CONTA_TMP_REG_2__SCAN_IN), .Y(n143));
  NAND4X1 g018(.A(n132), .B(n135), .C(CONTA_TMP_REG_1__SCAN_IN), .D(n143), .Y(n144));
  OAI21X1 g019(.A0(n129), .A1(n127), .B0(CANALE_REG_1__SCAN_IN), .Y(n145));
  NAND4X1 g020(.A(n132), .B(CONTA_TMP_REG_0__SCAN_IN), .C(n134), .D(n143), .Y(n146));
  NAND3X1 g021(.A(n146), .B(n145), .C(n144), .Y(U414));
  NAND3X1 g022(.A(n143), .B(n132), .C(n135), .Y(n148));
  OAI21X1 g023(.A0(n129), .A1(n127), .B0(CANALE_REG_0__SCAN_IN), .Y(n149));
  NAND2X1 g024(.A(n149), .B(n148), .Y(U413));
  NOR4X1  g025(.A(n127), .B(n135), .C(n134), .D(n129), .Y(n151));
  AOI21X1 g026(.A0(n151), .A1(CONTA_TMP_REG_2__SCAN_IN), .B0(n126), .Y(U417));
  NAND3X1 g027(.A(n143), .B(n136), .C(n132), .Y(n153));
  OAI21X1 g028(.A0(n151), .A1(n140), .B0(n153), .Y(U412));
  NOR4X1  g029(.A(n131), .B(n127), .C(n135), .D(S1_REG_0__SCAN_IN), .Y(n155));
  OAI21X1 g030(.A0(n155), .A1(n134), .B0(n146), .Y(U411));
  OAI21X1 g031(.A0(n132), .A1(n135), .B0(n148), .Y(U410));
  INVX1   g032(.A(ITFC_STATE_REG_1__SCAN_IN), .Y(n158));
  INVX1   g033(.A(TX_END_REG_SCAN_IN), .Y(n159));
  OAI21X1 g034(.A0(n158), .A1(n159), .B0(ITFC_STATE_REG_0__SCAN_IN), .Y(n160));
  OAI21X1 g035(.A0(ITFC_STATE_REG_0__SCAN_IN), .A1(n158), .B0(n160), .Y(U452));
  INVX1   g036(.A(SHOT_REG_SCAN_IN), .Y(n162));
  NAND2X1 g037(.A(ITFC_STATE_REG_0__SCAN_IN), .B(TX_END_REG_SCAN_IN), .Y(n163));
  NAND2X1 g038(.A(n163), .B(ITFC_STATE_REG_1__SCAN_IN), .Y(n164));
  OAI21X1 g039(.A0(n162), .A1(ITFC_STATE_REG_0__SCAN_IN), .B0(n164), .Y(U409));
  INVX1   g040(.A(TRE_REG_SCAN_IN), .Y(n166));
  NAND3X1 g041(.A(n166), .B(LOAD_REG_SCAN_IN), .C(DATA_IN_7_), .Y(n167));
  INVX1   g042(.A(LOAD_REG_SCAN_IN), .Y(n168));
  OAI21X1 g043(.A0(TRE_REG_SCAN_IN), .A1(n168), .B0(OUT_REG_REG_7__SCAN_IN), .Y(n169));
  NAND2X1 g044(.A(n169), .B(n167), .Y(U453));
  NAND3X1 g045(.A(n166), .B(LOAD_REG_SCAN_IN), .C(DATA_IN_6_), .Y(n171));
  OAI21X1 g046(.A0(TRE_REG_SCAN_IN), .A1(n168), .B0(OUT_REG_REG_6__SCAN_IN), .Y(n172));
  NAND2X1 g047(.A(n172), .B(n171), .Y(U454));
  NAND3X1 g048(.A(n166), .B(LOAD_REG_SCAN_IN), .C(DATA_IN_5_), .Y(n174));
  OAI21X1 g049(.A0(TRE_REG_SCAN_IN), .A1(n168), .B0(OUT_REG_REG_5__SCAN_IN), .Y(n175));
  NAND2X1 g050(.A(n175), .B(n174), .Y(U455));
  NAND3X1 g051(.A(n166), .B(LOAD_REG_SCAN_IN), .C(DATA_IN_4_), .Y(n177));
  OAI21X1 g052(.A0(TRE_REG_SCAN_IN), .A1(n168), .B0(OUT_REG_REG_4__SCAN_IN), .Y(n178));
  NAND2X1 g053(.A(n178), .B(n177), .Y(U456));
  NAND3X1 g054(.A(n166), .B(LOAD_REG_SCAN_IN), .C(DATA_IN_3_), .Y(n180));
  OAI21X1 g055(.A0(TRE_REG_SCAN_IN), .A1(n168), .B0(OUT_REG_REG_3__SCAN_IN), .Y(n181));
  NAND2X1 g056(.A(n181), .B(n180), .Y(U457));
  NAND3X1 g057(.A(n166), .B(LOAD_REG_SCAN_IN), .C(DATA_IN_2_), .Y(n183));
  OAI21X1 g058(.A0(TRE_REG_SCAN_IN), .A1(n168), .B0(OUT_REG_REG_2__SCAN_IN), .Y(n184));
  NAND2X1 g059(.A(n184), .B(n183), .Y(U458));
  NAND3X1 g060(.A(n166), .B(LOAD_REG_SCAN_IN), .C(DATA_IN_1_), .Y(n186));
  OAI21X1 g061(.A0(TRE_REG_SCAN_IN), .A1(n168), .B0(OUT_REG_REG_1__SCAN_IN), .Y(n187));
  NAND2X1 g062(.A(n187), .B(n186), .Y(U459));
  NAND3X1 g063(.A(n166), .B(LOAD_REG_SCAN_IN), .C(DATA_IN_0_), .Y(n189));
  OAI21X1 g064(.A0(TRE_REG_SCAN_IN), .A1(n168), .B0(OUT_REG_REG_0__SCAN_IN), .Y(n190));
  NAND2X1 g065(.A(n190), .B(n189), .Y(U460));
  INVX1   g066(.A(NEXT_BIT_REG_3__SCAN_IN), .Y(n192));
  INVX1   g067(.A(NEXT_BIT_REG_0__SCAN_IN), .Y(n193));
  INVX1   g068(.A(SEND_EN_REG_SCAN_IN), .Y(n194));
  INVX1   g069(.A(TX_CONTA_REG_4__SCAN_IN), .Y(n195));
  INVX1   g070(.A(TX_CONTA_REG_3__SCAN_IN), .Y(n196));
  NOR3X1  g071(.A(TX_CONTA_REG_0__SCAN_IN), .B(TX_CONTA_REG_1__SCAN_IN), .C(TX_CONTA_REG_2__SCAN_IN), .Y(n197));
  OAI21X1 g072(.A0(n197), .A1(n196), .B0(n195), .Y(n198));
  INVX1   g073(.A(TX_CONTA_REG_6__SCAN_IN), .Y(n199));
  INVX1   g074(.A(TX_CONTA_REG_5__SCAN_IN), .Y(n200));
  NOR2X1  g075(.A(n200), .B(n199), .Y(n201));
  INVX1   g076(.A(TX_CONTA_REG_9__SCAN_IN), .Y(n202));
  INVX1   g077(.A(TX_CONTA_REG_8__SCAN_IN), .Y(n203));
  INVX1   g078(.A(TX_CONTA_REG_7__SCAN_IN), .Y(n204));
  NAND3X1 g079(.A(n204), .B(n203), .C(n202), .Y(n205));
  AOI21X1 g080(.A0(n201), .A1(n198), .B0(n205), .Y(n206));
  NOR3X1  g081(.A(n206), .B(n194), .C(n193), .Y(n207));
  NAND3X1 g082(.A(n207), .B(NEXT_BIT_REG_1__SCAN_IN), .C(NEXT_BIT_REG_2__SCAN_IN), .Y(n208));
  OAI21X1 g083(.A0(n207), .A1(n192), .B0(n208), .Y(U461));
  INVX1   g084(.A(NEXT_BIT_REG_2__SCAN_IN), .Y(n210));
  NAND3X1 g085(.A(n207), .B(NEXT_BIT_REG_1__SCAN_IN), .C(n210), .Y(n211));
  INVX1   g086(.A(NEXT_BIT_REG_1__SCAN_IN), .Y(n212));
  NOR2X1  g087(.A(n206), .B(n194), .Y(n213));
  NAND2X1 g088(.A(n213), .B(NEXT_BIT_REG_0__SCAN_IN), .Y(n214));
  OAI21X1 g089(.A0(n214), .A1(n212), .B0(NEXT_BIT_REG_2__SCAN_IN), .Y(n215));
  NAND2X1 g090(.A(n215), .B(n211), .Y(U408));
  OAI21X1 g091(.A0(NEXT_BIT_REG_2__SCAN_IN), .A1(NEXT_BIT_REG_3__SCAN_IN), .B0(n193), .Y(n217));
  OAI21X1 g092(.A0(NEXT_BIT_REG_1__SCAN_IN), .A1(n210), .B0(NEXT_BIT_REG_0__SCAN_IN), .Y(n218));
  NAND3X1 g093(.A(n218), .B(n217), .C(n213), .Y(n219));
  OAI21X1 g094(.A0(n207), .A1(n212), .B0(n219), .Y(U407));
  AOI21X1 g095(.A0(n212), .A1(n210), .B0(NEXT_BIT_REG_0__SCAN_IN), .Y(n221));
  OAI21X1 g096(.A0(n221), .A1(NEXT_BIT_REG_3__SCAN_IN), .B0(n213), .Y(n222));
  OAI21X1 g097(.A0(n213), .A1(n193), .B0(n222), .Y(U462));
  NAND4X1 g098(.A(TX_CONTA_REG_1__SCAN_IN), .B(TX_CONTA_REG_2__SCAN_IN), .C(TX_CONTA_REG_3__SCAN_IN), .D(TX_CONTA_REG_0__SCAN_IN), .Y(n224));
  NOR4X1  g099(.A(n195), .B(n200), .C(n199), .D(n224), .Y(n225));
  NAND3X1 g100(.A(n225), .B(TX_CONTA_REG_7__SCAN_IN), .C(TX_CONTA_REG_8__SCAN_IN), .Y(n226));
  XOR2X1  g101(.A(n226), .B(TX_CONTA_REG_9__SCAN_IN), .Y(n227));
  NAND2X1 g102(.A(n206), .B(SEND_EN_REG_SCAN_IN), .Y(n228));
  OAI22X1 g103(.A0(n227), .A1(n228), .B0(SEND_EN_REG_SCAN_IN), .B1(n202), .Y(U406));
  NAND2X1 g104(.A(n225), .B(TX_CONTA_REG_7__SCAN_IN), .Y(n230));
  XOR2X1  g105(.A(n230), .B(TX_CONTA_REG_8__SCAN_IN), .Y(n231));
  OAI22X1 g106(.A0(n228), .A1(n231), .B0(SEND_EN_REG_SCAN_IN), .B1(n203), .Y(U405));
  XOR2X1  g107(.A(n225), .B(n204), .Y(n233));
  OAI22X1 g108(.A0(n228), .A1(n233), .B0(SEND_EN_REG_SCAN_IN), .B1(n204), .Y(U404));
  NOR3X1  g109(.A(n224), .B(n195), .C(n200), .Y(n235));
  XOR2X1  g110(.A(n235), .B(n199), .Y(n236));
  OAI22X1 g111(.A0(n228), .A1(n236), .B0(SEND_EN_REG_SCAN_IN), .B1(n199), .Y(U403));
  NOR2X1  g112(.A(n224), .B(n195), .Y(n238));
  XOR2X1  g113(.A(n238), .B(n200), .Y(n239));
  OAI22X1 g114(.A0(n228), .A1(n239), .B0(SEND_EN_REG_SCAN_IN), .B1(n200), .Y(U402));
  XOR2X1  g115(.A(n224), .B(TX_CONTA_REG_4__SCAN_IN), .Y(n241));
  OAI22X1 g116(.A0(n228), .A1(n241), .B0(SEND_EN_REG_SCAN_IN), .B1(n195), .Y(U401));
  NAND3X1 g117(.A(TX_CONTA_REG_0__SCAN_IN), .B(TX_CONTA_REG_1__SCAN_IN), .C(TX_CONTA_REG_2__SCAN_IN), .Y(n243));
  XOR2X1  g118(.A(n243), .B(TX_CONTA_REG_3__SCAN_IN), .Y(n244));
  OAI22X1 g119(.A0(n228), .A1(n244), .B0(SEND_EN_REG_SCAN_IN), .B1(n196), .Y(U400));
  NAND2X1 g120(.A(n194), .B(TX_CONTA_REG_2__SCAN_IN), .Y(n246));
  NAND2X1 g121(.A(TX_CONTA_REG_0__SCAN_IN), .B(TX_CONTA_REG_1__SCAN_IN), .Y(n247));
  XOR2X1  g122(.A(n247), .B(TX_CONTA_REG_2__SCAN_IN), .Y(n248));
  OAI21X1 g123(.A0(n248), .A1(n228), .B0(n246), .Y(U399));
  INVX1   g124(.A(TX_CONTA_REG_1__SCAN_IN), .Y(n250));
  XOR2X1  g125(.A(TX_CONTA_REG_0__SCAN_IN), .B(n250), .Y(n251));
  OAI22X1 g126(.A0(n228), .A1(n251), .B0(SEND_EN_REG_SCAN_IN), .B1(n250), .Y(U398));
  NAND2X1 g127(.A(n194), .B(TX_CONTA_REG_0__SCAN_IN), .Y(n253));
  OAI21X1 g128(.A0(n228), .A1(TX_CONTA_REG_0__SCAN_IN), .B0(n253), .Y(U397));
  INVX1   g129(.A(ITFC_STATE_REG_0__SCAN_IN), .Y(n255));
  OAI21X1 g130(.A0(n255), .A1(ITFC_STATE_REG_1__SCAN_IN), .B0(LOAD_REG_SCAN_IN), .Y(n256));
  NOR2X1  g131(.A(ITFC_STATE_REG_0__SCAN_IN), .B(ITFC_STATE_REG_1__SCAN_IN), .Y(n257));
  NAND2X1 g132(.A(n257), .B(SHOT_REG_SCAN_IN), .Y(n258));
  NAND2X1 g133(.A(n258), .B(n256), .Y(U396));
  NAND3X1 g134(.A(S1_REG_0__SCAN_IN), .B(S1_REG_1__SCAN_IN), .C(RDY_REG_SCAN_IN), .Y(n260));
  NAND2X1 g135(.A(n260), .B(SEND_DATA_REG_SCAN_IN), .Y(n261));
  NAND3X1 g136(.A(S1_REG_0__SCAN_IN), .B(S1_REG_1__SCAN_IN), .C(S1_REG_2__SCAN_IN), .Y(n262));
  NAND2X1 g137(.A(n262), .B(n261), .Y(U395));
  NAND3X1 g138(.A(SEND_REG_SCAN_IN), .B(TRE_REG_SCAN_IN), .C(DSR), .Y(n264));
  OAI21X1 g139(.A0(n194), .A1(TX_END_REG_SCAN_IN), .B0(n264), .Y(U394));
  NOR2X1  g140(.A(S1_REG_1__SCAN_IN), .B(EOC), .Y(n266));
  NAND3X1 g141(.A(n266), .B(S1_REG_0__SCAN_IN), .C(S1_REG_2__SCAN_IN), .Y(n267));
  NAND2X1 g142(.A(n267), .B(MUX_EN_REG_SCAN_IN), .Y(n268));
  NAND3X1 g143(.A(n128), .B(n131), .C(n127), .Y(n269));
  NAND2X1 g144(.A(n269), .B(n268), .Y(U393));
  NAND3X1 g145(.A(n166), .B(n168), .C(n159), .Y(U392));
  INVX1   g146(.A(LOAD_DATO_REG_SCAN_IN), .Y(n272));
  OAI21X1 g147(.A0(n132), .A1(n272), .B0(n267), .Y(U391));
  OAI21X1 g148(.A0(S1_REG_0__SCAN_IN), .A1(n131), .B0(SOC_REG_SCAN_IN), .Y(n274));
  OAI21X1 g149(.A0(n129), .A1(S1_REG_2__SCAN_IN), .B0(n274), .Y(U450));
  OAI21X1 g150(.A0(ITFC_STATE_REG_0__SCAN_IN), .A1(n158), .B0(SEND_REG_SCAN_IN), .Y(n276));
  OAI21X1 g151(.A0(n255), .A1(ITFC_STATE_REG_1__SCAN_IN), .B0(n276), .Y(U390));
  INVX1   g152(.A(MPX_REG_SCAN_IN), .Y(n278));
  INVX1   g153(.A(S2_REG_0__SCAN_IN), .Y(n279));
  NAND3X1 g154(.A(CONFIRM_REG_SCAN_IN), .B(S2_REG_1__SCAN_IN), .C(n279), .Y(n280));
  XOR2X1  g155(.A(n280), .B(n278), .Y(U389));
  INVX1   g156(.A(CONFIRM_REG_SCAN_IN), .Y(n282));
  OAI22X1 g157(.A0(n163), .A1(n158), .B0(n282), .B1(n257), .Y(U388));
  INVX1   g158(.A(S2_REG_1__SCAN_IN), .Y(n284));
  NAND2X1 g159(.A(n284), .B(S2_REG_0__SCAN_IN), .Y(n285));
  NOR3X1  g160(.A(CONFIRM_REG_SCAN_IN), .B(n284), .C(S2_REG_0__SCAN_IN), .Y(n286));
  OAI21X1 g161(.A0(n286), .A1(n162), .B0(n285), .Y(U387));
  INVX1   g162(.A(ADD_MPX2_REG_SCAN_IN), .Y(n288));
  OAI21X1 g163(.A0(n280), .A1(MPX_REG_SCAN_IN), .B0(n288), .Y(U386));
  INVX1   g164(.A(RDY_REG_SCAN_IN), .Y(n290));
  NAND3X1 g165(.A(SEND_DATA_REG_SCAN_IN), .B(n284), .C(n279), .Y(n291));
  NOR4X1  g166(.A(n278), .B(n284), .C(S2_REG_0__SCAN_IN), .D(n282), .Y(n292));
  OAI21X1 g167(.A0(n292), .A1(n290), .B0(n291), .Y(U385));
  NOR2X1  g168(.A(n166), .B(n168), .Y(n294));
  AOI21X1 g169(.A0(ERROR_REG_SCAN_IN), .A1(n168), .B0(n294), .Y(n295));
  NAND2X1 g170(.A(TRE_REG_SCAN_IN), .B(DSR), .Y(n296));
  NAND2X1 g171(.A(n296), .B(SEND_REG_SCAN_IN), .Y(n297));
  OAI21X1 g172(.A0(n295), .A1(SEND_REG_SCAN_IN), .B0(n297), .Y(U451));
  OAI21X1 g173(.A0(n128), .A1(n127), .B0(n129), .Y(U383));
  AOI21X1 g174(.A0(S1_REG_1__SCAN_IN), .A1(RDY_REG_SCAN_IN), .B0(S1_REG_2__SCAN_IN), .Y(n300));
  OAI21X1 g175(.A0(n300), .A1(n266), .B0(S1_REG_0__SCAN_IN), .Y(n301));
  OAI21X1 g176(.A0(S1_REG_0__SCAN_IN), .A1(n127), .B0(n301), .Y(U464));
  NAND3X1 g177(.A(S1_REG_1__SCAN_IN), .B(n127), .C(n290), .Y(n303));
  NAND3X1 g178(.A(n131), .B(S1_REG_2__SCAN_IN), .C(EOC), .Y(n304));
  NAND3X1 g179(.A(n304), .B(n303), .C(S1_REG_0__SCAN_IN), .Y(U384));
  NOR2X1  g180(.A(n282), .B(MPX_REG_SCAN_IN), .Y(n306));
  NAND2X1 g181(.A(S2_REG_1__SCAN_IN), .B(n279), .Y(n307));
  OAI21X1 g182(.A0(n307), .A1(n306), .B0(n285), .Y(U463));
  NAND2X1 g183(.A(n291), .B(n280), .Y(U382));
  NAND3X1 g184(.A(n212), .B(n210), .C(n192), .Y(n310));
  NOR4X1  g185(.A(n206), .B(n194), .C(n193), .D(n310), .Y(U381));
  NAND3X1 g186(.A(NEXT_BIT_REG_1__SCAN_IN), .B(n210), .C(OUT_REG_REG_7__SCAN_IN), .Y(n312));
  NAND2X1 g187(.A(NEXT_BIT_REG_3__SCAN_IN), .B(OUT_REG_REG_1__SCAN_IN), .Y(n313));
  NAND3X1 g188(.A(NEXT_BIT_REG_1__SCAN_IN), .B(NEXT_BIT_REG_2__SCAN_IN), .C(OUT_REG_REG_3__SCAN_IN), .Y(n314));
  NAND3X1 g189(.A(n212), .B(NEXT_BIT_REG_2__SCAN_IN), .C(OUT_REG_REG_5__SCAN_IN), .Y(n315));
  NAND4X1 g190(.A(n314), .B(n313), .C(n312), .D(n315), .Y(n316));
  NAND2X1 g191(.A(n316), .B(n193), .Y(n317));
  NOR2X1  g192(.A(NEXT_BIT_REG_1__SCAN_IN), .B(n210), .Y(n318));
  AOI22X1 g193(.A0(NEXT_BIT_REG_3__SCAN_IN), .A1(OUT_REG_REG_0__SCAN_IN), .B0(OUT_REG_REG_4__SCAN_IN), .B1(n318), .Y(n319));
  NAND3X1 g194(.A(NEXT_BIT_REG_1__SCAN_IN), .B(n210), .C(OUT_REG_REG_6__SCAN_IN), .Y(n320));
  NAND3X1 g195(.A(NEXT_BIT_REG_1__SCAN_IN), .B(NEXT_BIT_REG_2__SCAN_IN), .C(OUT_REG_REG_2__SCAN_IN), .Y(n321));
  NAND4X1 g196(.A(n320), .B(n319), .C(n310), .D(n321), .Y(n322));
  NAND2X1 g197(.A(n322), .B(NEXT_BIT_REG_0__SCAN_IN), .Y(n323));
  NAND3X1 g198(.A(n323), .B(n317), .C(n213), .Y(U380));
endmodule


