//Converted to Combinational (Partial output: n485) , Module name: s15850_n485 , Timestamp: 2018-12-03T15:51:04.842243 
module s15850_n485 ( g599, g591, g605, g611, g713, g617, g731, g718, g722, g627, g639, g654, g646, g650, g643, g695, g704, g677, g686, g668, g658, n485 );
input g599, g591, g605, g611, g713, g617, g731, g718, g722, g627, g639, g654, g646, g650, g643, g695, g704, g677, g686, g668, g658;
output n485;
wire n2478, n2461, n2473, n2477, n2474, n2462, n2475_1, n2446, n2460_1, n2430, n2472, n2476, n2437, n2442, n2445_1, n2459, n2465_1, n2471, n2441, n2434, n2438, n2444, n2458, n2447, n2464, n2452, n2453, n2470_1, n2466, n2467, n2454, n2439, n2440_1, n2433, n2435, n2436_1, n2443, n2451, n2457, n2463, n2469, n2431_1, n2432, n2448, n2449, n2450_1, n2456, n2455_1, n2468;
OAI21X1  g0639(.A0(n2473), .A1(n2461), .B0(n2478), .Y(n485));
OR4X1    g0638(.A(n2475_1), .B(n2462), .C(n2474), .D(n2477), .Y(n2478));
MX2X1    g0621(.A(n2430), .B(n2460_1), .S0(n2446), .Y(n2461));
OR2X1    g0633(.A(n2472), .B(n2462), .Y(n2473));
INVX1    g0637(.A(n2476), .Y(n2477));
NOR3X1   g0634(.A(n2437), .B(g591), .C(g599), .Y(n2474));
NOR4X1   g0622(.A(g591), .B(g599), .C(g611), .D(g605), .Y(n2462));
INVX1    g0635(.A(n2472), .Y(n2475_1));
NAND2X1  g0606(.A(n2445_1), .B(n2442), .Y(n2446));
XOR2X1   g0620(.A(n2459), .B(g713), .Y(n2460_1));
INVX1    g0590(.A(g713), .Y(n2430));
AOI21X1  g0632(.A0(n2471), .A1(n2465_1), .B0(n2442), .Y(n2472));
AOI21X1  g0636(.A0(n2437), .A1(g599), .B0(n2441), .Y(n2476));
INVX1    g0597(.A(g605), .Y(n2437));
OAI21X1  g0602(.A0(n2441), .A1(n2438), .B0(n2434), .Y(n2442));
OAI21X1  g0605(.A0(n2444), .A1(g617), .B0(n2434), .Y(n2445_1));
MX2X1    g0619(.A(n2447), .B(n2458), .S0(n2445_1), .Y(n2459));
OR4X1    g0625(.A(n2453), .B(n2452), .C(g731), .D(n2464), .Y(n2465_1));
OR4X1    g0631(.A(n2454), .B(n2467), .C(n2466), .D(n2470_1), .Y(n2471));
NOR3X1   g0601(.A(n2440_1), .B(g617), .C(n2439), .Y(n2441));
INVX1    g0594(.A(n2433), .Y(n2434));
AOI21X1  g0598(.A0(n2437), .A1(n2436_1), .B0(n2435), .Y(n2438));
NOR4X1   g0604(.A(n2440_1), .B(g599), .C(g617), .D(n2443), .Y(n2444));
MX2X1    g0618(.A(n2457), .B(n2451), .S0(n2454), .Y(n2458));
INVX1    g0607(.A(g718), .Y(n2447));
OR2X1    g0624(.A(n2463), .B(g722), .Y(n2464));
NOR3X1   g0612(.A(g605), .B(g591), .C(n2436_1), .Y(n2452));
AOI21X1  g0613(.A0(n2437), .A1(n2440_1), .B0(g599), .Y(n2453));
INVX1    g0630(.A(n2469), .Y(n2470_1));
INVX1    g0626(.A(g722), .Y(n2466));
INVX1    g0627(.A(g731), .Y(n2467));
NOR2X1   g0614(.A(n2453), .B(n2452), .Y(n2454));
INVX1    g0599(.A(g611), .Y(n2439));
INVX1    g0600(.A(g591), .Y(n2440_1));
NAND3X1  g0593(.A(n2432), .B(n2431_1), .C(g627), .Y(n2433));
INVX1    g0595(.A(g639), .Y(n2435));
INVX1    g0596(.A(g599), .Y(n2436_1));
OR2X1    g0603(.A(g605), .B(g611), .Y(n2443));
NAND3X1  g0611(.A(n2450_1), .B(n2449), .C(n2448), .Y(n2451));
OR4X1    g0617(.A(n2455_1), .B(n2449), .C(n2448), .D(n2456), .Y(n2457));
NAND4X1  g0623(.A(n2449), .B(n2448), .C(n2430), .D(n2450_1), .Y(n2463));
NOR4X1   g0629(.A(n2449), .B(n2448), .C(n2430), .D(n2468), .Y(n2469));
INVX1    g0591(.A(g654), .Y(n2431_1));
NOR3X1   g0592(.A(g643), .B(g650), .C(g646), .Y(n2432));
INVX1    g0608(.A(g695), .Y(n2448));
INVX1    g0609(.A(g704), .Y(n2449));
NOR4X1   g0610(.A(g658), .B(g668), .C(g686), .D(g677), .Y(n2450_1));
NAND3X1  g0616(.A(g677), .B(g658), .C(g668), .Y(n2456));
INVX1    g0615(.A(g686), .Y(n2455_1));
NAND4X1  g0628(.A(g658), .B(g668), .C(g686), .D(g677), .Y(n2468));

endmodule
