//Converted to Combinational (Partial output: CRC_OUT_2_20) , Module name: s35932_CRC_OUT_2_20 , Timestamp: 2018-12-03T15:51:11.038754 
module s35932_CRC_OUT_2_20 ( RESET, WX9910, WX9912, WX9914, WX9916, WX9918, WX9920, WX9888, WX9922, WX9890, WX9924, WX9892, WX9926, WX9894, WX9928, WX9896, WX9930, WX9898, WX9932, WX9900, WX9934, WX9902, WX9936, WX9904, WX9938, WX9906, WX9940, WX9908, WX9942, WX9944, WX9946, WX9948, WX9950, CRC_OUT_2_20 );
input RESET, WX9910, WX9912, WX9914, WX9916, WX9918, WX9920, WX9888, WX9922, WX9890, WX9924, WX9892, WX9926, WX9894, WX9928, WX9896, WX9930, WX9898, WX9932, WX9900, WX9934, WX9902, WX9936, WX9904, WX9938, WX9906, WX9940, WX9908, WX9942, WX9944, WX9946, WX9948, WX9950;
output CRC_OUT_2_20;
wire n5827, n10405, CRC_OUT_2_19, n10403, CRC_OUT_2_18, n10401, CRC_OUT_2_17, n10399, CRC_OUT_2_16, n10397, CRC_OUT_2_15, n10396, n10394, CRC_OUT_2_31, CRC_OUT_2_14, n10427, n10392, CRC_OUT_2_30, CRC_OUT_2_13, n10425, n10390, CRC_OUT_2_29, CRC_OUT_2_12, n10423, n10388, CRC_OUT_2_28, CRC_OUT_2_11, n10421, n10386, CRC_OUT_2_27, CRC_OUT_2_10, n10385, n10419, n10383, CRC_OUT_2_26, CRC_OUT_2_9, n10417, n10381, CRC_OUT_2_25, CRC_OUT_2_8, n10415, n10379, CRC_OUT_2_24, CRC_OUT_2_7, n10413, n10377, CRC_OUT_2_23, CRC_OUT_2_6, n10411, n10375, CRC_OUT_2_22, CRC_OUT_2_5, n10409, n10373, CRC_OUT_2_21, CRC_OUT_2_4, n10407, n10371, CRC_OUT_2_3, n10370, n10368, CRC_OUT_2_2, n10366, CRC_OUT_2_1, n10364, CRC_OUT_2_0, n10362;
NOR2X1   g4611(.A(n10405), .B(n5827), .Y(CRC_OUT_2_20));
INVX1    g0288(.A(RESET), .Y(n5827));
XOR2X1   g4610(.A(CRC_OUT_2_19), .B(WX9910), .Y(n10405));
NOR2X1   g4609(.A(n10403), .B(n5827), .Y(CRC_OUT_2_19));
XOR2X1   g4608(.A(CRC_OUT_2_18), .B(WX9912), .Y(n10403));
NOR2X1   g4607(.A(n10401), .B(n5827), .Y(CRC_OUT_2_18));
XOR2X1   g4606(.A(CRC_OUT_2_17), .B(WX9914), .Y(n10401));
NOR2X1   g4605(.A(n10399), .B(n5827), .Y(CRC_OUT_2_17));
XOR2X1   g4604(.A(CRC_OUT_2_16), .B(WX9916), .Y(n10399));
NOR2X1   g4603(.A(n10397), .B(n5827), .Y(CRC_OUT_2_16));
XOR2X1   g4602(.A(n10396), .B(CRC_OUT_2_15), .Y(n10397));
NOR2X1   g4600(.A(n10394), .B(n5827), .Y(CRC_OUT_2_15));
XOR2X1   g4601(.A(CRC_OUT_2_31), .B(WX9918), .Y(n10396));
XOR2X1   g4599(.A(CRC_OUT_2_14), .B(WX9920), .Y(n10394));
NOR2X1   g4633(.A(n10427), .B(n5827), .Y(CRC_OUT_2_31));
NOR2X1   g4598(.A(n10392), .B(n5827), .Y(CRC_OUT_2_14));
XOR2X1   g4632(.A(CRC_OUT_2_30), .B(WX9888), .Y(n10427));
XOR2X1   g4597(.A(CRC_OUT_2_13), .B(WX9922), .Y(n10392));
NOR2X1   g4631(.A(n10425), .B(n5827), .Y(CRC_OUT_2_30));
NOR2X1   g4596(.A(n10390), .B(n5827), .Y(CRC_OUT_2_13));
XOR2X1   g4630(.A(CRC_OUT_2_29), .B(WX9890), .Y(n10425));
XOR2X1   g4595(.A(CRC_OUT_2_12), .B(WX9924), .Y(n10390));
NOR2X1   g4629(.A(n10423), .B(n5827), .Y(CRC_OUT_2_29));
NOR2X1   g4594(.A(n10388), .B(n5827), .Y(CRC_OUT_2_12));
XOR2X1   g4628(.A(CRC_OUT_2_28), .B(WX9892), .Y(n10423));
XOR2X1   g4593(.A(CRC_OUT_2_11), .B(WX9926), .Y(n10388));
NOR2X1   g4627(.A(n10421), .B(n5827), .Y(CRC_OUT_2_28));
NOR2X1   g4592(.A(n10386), .B(n5827), .Y(CRC_OUT_2_11));
XOR2X1   g4626(.A(CRC_OUT_2_27), .B(WX9894), .Y(n10421));
XOR2X1   g4591(.A(n10385), .B(CRC_OUT_2_10), .Y(n10386));
NOR2X1   g4625(.A(n10419), .B(n5827), .Y(CRC_OUT_2_27));
NOR2X1   g4589(.A(n10383), .B(n5827), .Y(CRC_OUT_2_10));
XOR2X1   g4590(.A(CRC_OUT_2_31), .B(WX9928), .Y(n10385));
XOR2X1   g4624(.A(CRC_OUT_2_26), .B(WX9896), .Y(n10419));
XOR2X1   g4588(.A(CRC_OUT_2_9), .B(WX9930), .Y(n10383));
NOR2X1   g4623(.A(n10417), .B(n5827), .Y(CRC_OUT_2_26));
NOR2X1   g4587(.A(n10381), .B(n5827), .Y(CRC_OUT_2_9));
XOR2X1   g4622(.A(CRC_OUT_2_25), .B(WX9898), .Y(n10417));
XOR2X1   g4586(.A(CRC_OUT_2_8), .B(WX9932), .Y(n10381));
NOR2X1   g4621(.A(n10415), .B(n5827), .Y(CRC_OUT_2_25));
NOR2X1   g4585(.A(n10379), .B(n5827), .Y(CRC_OUT_2_8));
XOR2X1   g4620(.A(CRC_OUT_2_24), .B(WX9900), .Y(n10415));
XOR2X1   g4584(.A(CRC_OUT_2_7), .B(WX9934), .Y(n10379));
NOR2X1   g4619(.A(n10413), .B(n5827), .Y(CRC_OUT_2_24));
NOR2X1   g4583(.A(n10377), .B(n5827), .Y(CRC_OUT_2_7));
XOR2X1   g4618(.A(CRC_OUT_2_23), .B(WX9902), .Y(n10413));
XOR2X1   g4582(.A(CRC_OUT_2_6), .B(WX9936), .Y(n10377));
NOR2X1   g4617(.A(n10411), .B(n5827), .Y(CRC_OUT_2_23));
NOR2X1   g4581(.A(n10375), .B(n5827), .Y(CRC_OUT_2_6));
XOR2X1   g4616(.A(CRC_OUT_2_22), .B(WX9904), .Y(n10411));
XOR2X1   g4580(.A(CRC_OUT_2_5), .B(WX9938), .Y(n10375));
NOR2X1   g4615(.A(n10409), .B(n5827), .Y(CRC_OUT_2_22));
NOR2X1   g4579(.A(n10373), .B(n5827), .Y(CRC_OUT_2_5));
XOR2X1   g4614(.A(CRC_OUT_2_21), .B(WX9906), .Y(n10409));
XOR2X1   g4578(.A(CRC_OUT_2_4), .B(WX9940), .Y(n10373));
NOR2X1   g4613(.A(n10407), .B(n5827), .Y(CRC_OUT_2_21));
NOR2X1   g4577(.A(n10371), .B(n5827), .Y(CRC_OUT_2_4));
XOR2X1   g4612(.A(CRC_OUT_2_20), .B(WX9908), .Y(n10407));
XOR2X1   g4576(.A(n10370), .B(CRC_OUT_2_3), .Y(n10371));
NOR2X1   g4574(.A(n10368), .B(n5827), .Y(CRC_OUT_2_3));
XOR2X1   g4575(.A(CRC_OUT_2_31), .B(WX9942), .Y(n10370));
XOR2X1   g4573(.A(CRC_OUT_2_2), .B(WX9944), .Y(n10368));
NOR2X1   g4572(.A(n10366), .B(n5827), .Y(CRC_OUT_2_2));
XOR2X1   g4571(.A(CRC_OUT_2_1), .B(WX9946), .Y(n10366));
NOR2X1   g4570(.A(n10364), .B(n5827), .Y(CRC_OUT_2_1));
XOR2X1   g4569(.A(CRC_OUT_2_0), .B(WX9948), .Y(n10364));
NOR2X1   g4568(.A(n10362), .B(n5827), .Y(CRC_OUT_2_0));
XOR2X1   g4567(.A(CRC_OUT_2_31), .B(WX9950), .Y(n10362));

endmodule
