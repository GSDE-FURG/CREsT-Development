// Benchmark "b09_C" written by ABC on Wed Aug 05 14:39:26 2020

module b09_C ( 
    D_IN_REG_0__SCAN_IN, X, D_OUT_REG_7__SCAN_IN, D_OUT_REG_6__SCAN_IN,
    D_OUT_REG_5__SCAN_IN, D_OUT_REG_4__SCAN_IN, D_OUT_REG_3__SCAN_IN,
    D_OUT_REG_2__SCAN_IN, D_OUT_REG_1__SCAN_IN, D_OUT_REG_0__SCAN_IN,
    OLD_REG_7__SCAN_IN, OLD_REG_6__SCAN_IN, OLD_REG_5__SCAN_IN,
    OLD_REG_4__SCAN_IN, OLD_REG_3__SCAN_IN, OLD_REG_2__SCAN_IN,
    OLD_REG_1__SCAN_IN, OLD_REG_0__SCAN_IN, Y_REG_SCAN_IN,
    STATO_REG_1__SCAN_IN, STATO_REG_0__SCAN_IN, D_IN_REG_8__SCAN_IN,
    D_IN_REG_7__SCAN_IN, D_IN_REG_6__SCAN_IN, D_IN_REG_5__SCAN_IN,
    D_IN_REG_4__SCAN_IN, D_IN_REG_3__SCAN_IN, D_IN_REG_2__SCAN_IN,
    D_IN_REG_1__SCAN_IN,
    U118, U117, U116, U115, U114, U113, U112, U111, U110, U109, U108, U107,
    U106, U105, U104, U103, U102, U92, U91, U101, U100, U99, U98, U97, U96,
    U95, U94, U93  );
  input  D_IN_REG_0__SCAN_IN, X, D_OUT_REG_7__SCAN_IN,
    D_OUT_REG_6__SCAN_IN, D_OUT_REG_5__SCAN_IN, D_OUT_REG_4__SCAN_IN,
    D_OUT_REG_3__SCAN_IN, D_OUT_REG_2__SCAN_IN, D_OUT_REG_1__SCAN_IN,
    D_OUT_REG_0__SCAN_IN, OLD_REG_7__SCAN_IN, OLD_REG_6__SCAN_IN,
    OLD_REG_5__SCAN_IN, OLD_REG_4__SCAN_IN, OLD_REG_3__SCAN_IN,
    OLD_REG_2__SCAN_IN, OLD_REG_1__SCAN_IN, OLD_REG_0__SCAN_IN,
    Y_REG_SCAN_IN, STATO_REG_1__SCAN_IN, STATO_REG_0__SCAN_IN,
    D_IN_REG_8__SCAN_IN, D_IN_REG_7__SCAN_IN, D_IN_REG_6__SCAN_IN,
    D_IN_REG_5__SCAN_IN, D_IN_REG_4__SCAN_IN, D_IN_REG_3__SCAN_IN,
    D_IN_REG_2__SCAN_IN, D_IN_REG_1__SCAN_IN;
  output U118, U117, U116, U115, U114, U113, U112, U111, U110, U109, U108,
    U107, U106, U105, U104, U103, U102, U92, U91, U101, U100, U99, U98,
    U97, U96, U95, U94, U93;
  wire n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
    n72, n73, n74, n75, n76, n78, n79, n80, n82, n83, n85, n86, n88, n89,
    n91, n92, n94, n95, n97, n98, n100, n101, n102, n103, n105, n107, n109,
    n111, n113, n115, n117, n119, n120, n121, n122, n123, n126, n127, n128,
    n130, n131, n132, n133;
  INVX1   g00(.A(D_IN_REG_8__SCAN_IN), .Y(n58));
  NAND2X1 g01(.A(STATO_REG_0__SCAN_IN), .B(D_IN_REG_0__SCAN_IN), .Y(n59));
  XOR2X1  g02(.A(D_IN_REG_7__SCAN_IN), .B(OLD_REG_6__SCAN_IN), .Y(n60));
  XOR2X1  g03(.A(D_IN_REG_8__SCAN_IN), .B(OLD_REG_7__SCAN_IN), .Y(n61));
  XOR2X1  g04(.A(D_IN_REG_6__SCAN_IN), .B(OLD_REG_5__SCAN_IN), .Y(n62));
  XOR2X1  g05(.A(D_IN_REG_5__SCAN_IN), .B(OLD_REG_4__SCAN_IN), .Y(n63));
  NOR4X1  g06(.A(n62), .B(n61), .C(n60), .D(n63), .Y(n64));
  XOR2X1  g07(.A(D_IN_REG_2__SCAN_IN), .B(OLD_REG_1__SCAN_IN), .Y(n65));
  XOR2X1  g08(.A(D_IN_REG_1__SCAN_IN), .B(OLD_REG_0__SCAN_IN), .Y(n66));
  XOR2X1  g09(.A(D_IN_REG_4__SCAN_IN), .B(OLD_REG_3__SCAN_IN), .Y(n67));
  XOR2X1  g10(.A(D_IN_REG_3__SCAN_IN), .B(OLD_REG_2__SCAN_IN), .Y(n68));
  NOR4X1  g11(.A(n67), .B(n66), .C(n65), .D(n68), .Y(n69));
  AOI21X1 g12(.A0(n69), .A1(n64), .B0(n59), .Y(n70));
  INVX1   g13(.A(STATO_REG_1__SCAN_IN), .Y(n71));
  NAND2X1 g14(.A(n71), .B(D_IN_REG_0__SCAN_IN), .Y(n72));
  OAI21X1 g15(.A0(STATO_REG_0__SCAN_IN), .A1(D_IN_REG_0__SCAN_IN), .B0(n72), .Y(n73));
  NOR2X1  g16(.A(n73), .B(n70), .Y(n74));
  NAND2X1 g17(.A(n74), .B(D_OUT_REG_7__SCAN_IN), .Y(n75));
  OAI21X1 g18(.A0(n73), .A1(n70), .B0(STATO_REG_0__SCAN_IN), .Y(n76));
  OAI21X1 g19(.A0(n76), .A1(n58), .B0(n75), .Y(U118));
  INVX1   g20(.A(D_IN_REG_7__SCAN_IN), .Y(n78));
  NOR3X1  g21(.A(STATO_REG_0__SCAN_IN), .B(n71), .C(D_IN_REG_0__SCAN_IN), .Y(n79));
  AOI22X1 g22(.A0(n74), .A1(D_OUT_REG_6__SCAN_IN), .B0(D_OUT_REG_7__SCAN_IN), .B1(n79), .Y(n80));
  OAI21X1 g23(.A0(n76), .A1(n78), .B0(n80), .Y(U117));
  INVX1   g24(.A(D_IN_REG_6__SCAN_IN), .Y(n82));
  AOI22X1 g25(.A0(n74), .A1(D_OUT_REG_5__SCAN_IN), .B0(D_OUT_REG_6__SCAN_IN), .B1(n79), .Y(n83));
  OAI21X1 g26(.A0(n76), .A1(n82), .B0(n83), .Y(U116));
  INVX1   g27(.A(D_IN_REG_5__SCAN_IN), .Y(n85));
  AOI22X1 g28(.A0(n74), .A1(D_OUT_REG_4__SCAN_IN), .B0(D_OUT_REG_5__SCAN_IN), .B1(n79), .Y(n86));
  OAI21X1 g29(.A0(n76), .A1(n85), .B0(n86), .Y(U115));
  INVX1   g30(.A(D_IN_REG_4__SCAN_IN), .Y(n88));
  AOI22X1 g31(.A0(n74), .A1(D_OUT_REG_3__SCAN_IN), .B0(D_OUT_REG_4__SCAN_IN), .B1(n79), .Y(n89));
  OAI21X1 g32(.A0(n76), .A1(n88), .B0(n89), .Y(U114));
  INVX1   g33(.A(D_IN_REG_3__SCAN_IN), .Y(n91));
  AOI22X1 g34(.A0(n74), .A1(D_OUT_REG_2__SCAN_IN), .B0(D_OUT_REG_3__SCAN_IN), .B1(n79), .Y(n92));
  OAI21X1 g35(.A0(n76), .A1(n91), .B0(n92), .Y(U113));
  INVX1   g36(.A(D_IN_REG_2__SCAN_IN), .Y(n94));
  AOI22X1 g37(.A0(n74), .A1(D_OUT_REG_1__SCAN_IN), .B0(D_OUT_REG_2__SCAN_IN), .B1(n79), .Y(n95));
  OAI21X1 g38(.A0(n76), .A1(n94), .B0(n95), .Y(U112));
  INVX1   g39(.A(D_IN_REG_1__SCAN_IN), .Y(n97));
  AOI22X1 g40(.A0(n74), .A1(D_OUT_REG_0__SCAN_IN), .B0(D_OUT_REG_1__SCAN_IN), .B1(n79), .Y(n98));
  OAI21X1 g41(.A0(n76), .A1(n97), .B0(n98), .Y(U111));
  INVX1   g42(.A(OLD_REG_7__SCAN_IN), .Y(n100));
  INVX1   g43(.A(D_IN_REG_0__SCAN_IN), .Y(n101));
  NOR2X1  g44(.A(STATO_REG_0__SCAN_IN), .B(n71), .Y(n102));
  AOI21X1 g45(.A0(STATO_REG_0__SCAN_IN), .A1(n101), .B0(n102), .Y(n103));
  OAI22X1 g46(.A0(n59), .A1(n58), .B0(n100), .B1(n103), .Y(U110));
  INVX1   g47(.A(OLD_REG_6__SCAN_IN), .Y(n105));
  OAI22X1 g48(.A0(n59), .A1(n78), .B0(n105), .B1(n103), .Y(U109));
  INVX1   g49(.A(OLD_REG_5__SCAN_IN), .Y(n107));
  OAI22X1 g50(.A0(n59), .A1(n82), .B0(n107), .B1(n103), .Y(U108));
  INVX1   g51(.A(OLD_REG_4__SCAN_IN), .Y(n109));
  OAI22X1 g52(.A0(n59), .A1(n85), .B0(n109), .B1(n103), .Y(U107));
  INVX1   g53(.A(OLD_REG_3__SCAN_IN), .Y(n111));
  OAI22X1 g54(.A0(n59), .A1(n88), .B0(n111), .B1(n103), .Y(U106));
  INVX1   g55(.A(OLD_REG_2__SCAN_IN), .Y(n113));
  OAI22X1 g56(.A0(n59), .A1(n91), .B0(n113), .B1(n103), .Y(U105));
  INVX1   g57(.A(OLD_REG_1__SCAN_IN), .Y(n115));
  OAI22X1 g58(.A0(n59), .A1(n94), .B0(n115), .B1(n103), .Y(U104));
  INVX1   g59(.A(OLD_REG_0__SCAN_IN), .Y(n117));
  OAI22X1 g60(.A0(n59), .A1(n97), .B0(n117), .B1(n103), .Y(U103));
  INVX1   g61(.A(n70), .Y(n119));
  INVX1   g62(.A(STATO_REG_0__SCAN_IN), .Y(n120));
  NAND4X1 g63(.A(STATO_REG_1__SCAN_IN), .B(D_OUT_REG_0__SCAN_IN), .C(n101), .D(n120), .Y(n121));
  NOR2X1  g64(.A(n120), .B(STATO_REG_1__SCAN_IN), .Y(n122));
  OAI21X1 g65(.A0(Y_REG_SCAN_IN), .A1(D_IN_REG_0__SCAN_IN), .B0(n122), .Y(n123));
  NAND3X1 g66(.A(n123), .B(n121), .C(n119), .Y(U102));
  NAND2X1 g67(.A(n59), .B(n71), .Y(U92));
  NAND4X1 g68(.A(n64), .B(STATO_REG_0__SCAN_IN), .C(STATO_REG_1__SCAN_IN), .D(n69), .Y(n126));
  AOI21X1 g69(.A0(STATO_REG_1__SCAN_IN), .A1(n101), .B0(STATO_REG_0__SCAN_IN), .Y(n127));
  AOI21X1 g70(.A0(STATO_REG_0__SCAN_IN), .A1(n101), .B0(n127), .Y(n128));
  NAND2X1 g71(.A(n128), .B(n126), .Y(U91));
  NAND2X1 g72(.A(n69), .B(n64), .Y(n130));
  OAI21X1 g73(.A0(n130), .A1(n71), .B0(STATO_REG_0__SCAN_IN), .Y(n131));
  AOI21X1 g74(.A0(STATO_REG_0__SCAN_IN), .A1(D_IN_REG_0__SCAN_IN), .B0(n71), .Y(n132));
  OAI21X1 g75(.A0(n132), .A1(n122), .B0(X), .Y(n133));
  OAI21X1 g76(.A0(n131), .A1(n101), .B0(n133), .Y(U101));
  NOR2X1  g77(.A(n103), .B(n58), .Y(U100));
  NOR2X1  g78(.A(n103), .B(n78), .Y(U99));
  NOR2X1  g79(.A(n103), .B(n82), .Y(U98));
  NOR2X1  g80(.A(n103), .B(n85), .Y(U97));
  NOR2X1  g81(.A(n103), .B(n88), .Y(U96));
  NOR2X1  g82(.A(n103), .B(n91), .Y(U95));
  NOR2X1  g83(.A(n103), .B(n94), .Y(U94));
  NOR2X1  g84(.A(n103), .B(n97), .Y(U93));
endmodule


