//Converted to Combinational , Module name: s1196 , Timestamp: 2018-12-03T15:51:02.215802 
module s1196 ( G0, G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42, G43, G44, G46, G546, G539, G550, G551, G552, G547, G548, G549, G530, G45, G542, G532, G535, G537, n57, n62, n67, n72, n77, n82, n87, n92, n97, n102, n107, n112, n117, n122, n127, n132, n141 );
input G0, G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G29, G30, G31, G32, G33, G34, G35, G36, G37, G38, G39, G40, G41, G42, G43, G44, G46;
output G546, G539, G550, G551, G552, G547, G548, G549, G530, G45, G542, G532, G535, G537, n57, n62, n67, n72, n77, n82, n87, n92, n97, n102, n107, n112, n117, n122, n127, n132, n141;
wire n83, n84, n85, n86, n87_1, n88, n89, n90, n91, n92_1, n93, n94, n95, n96, n97_1, n98, n99, n100, n101, n102_1, n103, n104, n105, n106, n107_1, n108, n109, n110, n111, n112_1, n113, n114, n115, n116, n117_1, n118, n119, n120, n121, n122_1, n123, n124, n125, n126, n127_1, n128, n129, n130, n131, n132_1, n133, n134, n135, n136, n137_1, n138, n139, n140, n141_1, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n236, n237, n238, n239, n240, n241, n242, n243, n244, n246, n247, n248, n249, n250, n251, n252, n253, n254, n256, n257, n258, n259, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n273, n274, n275, n276, n277, n278, n279, n280, n281, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n348, n349, n353, n355, n356, n358, n360, n361, n363, n368, n369, n370, n371, n373, n374, n376, n377, n378, n379, n381, n382, n383, n384, n386, n387, n388, n390, n391, n393, n394, n395, n396, n397, n398, n399, n400, n401;
INVX1    g000(.A(G41), .Y(G546));
INVX1    g001(.A(G13), .Y(n83));
INVX1    g002(.A(G3), .Y(n84));
INVX1    g003(.A(G5), .Y(n85));
INVX1    g004(.A(G7), .Y(n86));
INVX1    g005(.A(G6), .Y(n87_1));
INVX1    g006(.A(G10), .Y(n88));
NOR4X1   g007(.A(G9), .B(G8), .C(n87_1), .D(n88), .Y(n89));
NAND4X1  g008(.A(n86), .B(n85), .C(n84), .D(n89), .Y(n90));
NAND2X1  g009(.A(G5), .B(G3), .Y(n91));
NAND2X1  g010(.A(G37), .B(G8), .Y(n92_1));
OR4X1    g011(.A(n91), .B(G10), .C(n86), .D(n92_1), .Y(n93));
NOR2X1   g012(.A(G4), .B(G0), .Y(n94));
NAND2X1  g013(.A(n94), .B(G11), .Y(n95));
AOI21X1  g014(.A0(n93), .A1(n90), .B0(n95), .Y(n96));
INVX1    g015(.A(G0), .Y(n97_1));
NAND3X1  g016(.A(G11), .B(G9), .C(G8), .Y(n98));
NAND2X1  g017(.A(G10), .B(G7), .Y(n99));
NAND2X1  g018(.A(G6), .B(G4), .Y(n100));
OR4X1    g019(.A(n99), .B(n98), .C(n91), .D(n100), .Y(n101));
NOR2X1   g020(.A(n101), .B(n97_1), .Y(n102_1));
AND2X1   g021(.A(G2), .B(G1), .Y(n103));
OAI21X1  g022(.A0(n102_1), .A1(n96), .B0(n103), .Y(n104));
INVX1    g023(.A(G4), .Y(n105));
NOR2X1   g024(.A(G5), .B(n105), .Y(n106));
AND2X1   g025(.A(G5), .B(G3), .Y(n107_1));
OAI22X1  g026(.A0(n85), .A1(G1), .B0(n105), .B1(n107_1), .Y(n108));
AOI21X1  g027(.A0(n108), .A1(G2), .B0(G3), .Y(n109));
AOI22X1  g028(.A0(n94), .A1(G3), .B0(n85), .B1(n109), .Y(n110));
NOR2X1   g029(.A(n110), .B(n106), .Y(n111));
INVX1    g030(.A(G8), .Y(n112_1));
INVX1    g031(.A(G30), .Y(n113));
NOR3X1   g032(.A(n113), .B(n86), .C(G6), .Y(n114));
INVX1    g033(.A(G9), .Y(n115));
AND2X1   g034(.A(G10), .B(G8), .Y(n116));
NOR2X1   g035(.A(n116), .B(n115), .Y(n117_1));
NOR4X1   g036(.A(n114), .B(G31), .C(n112_1), .D(n117_1), .Y(n118));
OR2X1    g037(.A(G8), .B(G7), .Y(n119));
OAI22X1  g038(.A0(G30), .A1(G6), .B0(G9), .B1(n119), .Y(n120));
OAI21X1  g039(.A0(n120), .A1(n118), .B0(G11), .Y(n121));
NAND3X1  g040(.A(G30), .B(G7), .C(n87_1), .Y(n122_1));
NOR3X1   g041(.A(G11), .B(G10), .C(G9), .Y(n123));
NAND2X1  g042(.A(G31), .B(G8), .Y(n124));
NAND3X1  g043(.A(n124), .B(n123), .C(n122_1), .Y(n125));
INVX1    g044(.A(G11), .Y(n126));
INVX1    g045(.A(G31), .Y(n127_1));
MX2X1    g046(.A(G10), .B(n127_1), .S0(G8), .Y(n128));
NAND4X1  g047(.A(n126), .B(G9), .C(n86), .D(n128), .Y(n129));
NAND4X1  g048(.A(n125), .B(n121), .C(G46), .D(n129), .Y(n130));
OR2X1    g049(.A(n130), .B(n111), .Y(n131));
NAND4X1  g050(.A(n104), .B(n83), .C(G12), .D(n131), .Y(n132_1));
INVX1    g051(.A(G1), .Y(n133));
NOR4X1   g052(.A(G4), .B(n84), .C(n133), .D(n87_1), .Y(n134));
NAND3X1  g053(.A(G6), .B(G4), .C(G3), .Y(n135));
NOR2X1   g054(.A(n135), .B(G1), .Y(n136));
NOR4X1   g055(.A(n88), .B(n115), .C(G8), .D(n126), .Y(n137_1));
OAI21X1  g056(.A0(n136), .A1(n134), .B0(n137_1), .Y(n138));
OR4X1    g057(.A(n98), .B(G10), .C(G1), .D(n135), .Y(n139));
AOI21X1  g058(.A0(n139), .A1(n138), .B0(G7), .Y(n140));
OR2X1    g059(.A(G6), .B(G4), .Y(n141_1));
OR4X1    g060(.A(G8), .B(n84), .C(G1), .D(n141_1), .Y(n142));
OAI21X1  g061(.A0(n136), .A1(n134), .B0(G8), .Y(n143));
NAND4X1  g062(.A(n88), .B(n115), .C(G7), .D(G11), .Y(n144));
AOI21X1  g063(.A0(n143), .A1(n142), .B0(n144), .Y(n145));
INVX1    g064(.A(G2), .Y(n146));
NOR2X1   g065(.A(G5), .B(n146), .Y(n147));
OAI21X1  g066(.A0(n145), .A1(n140), .B0(n147), .Y(n148));
OR2X1    g067(.A(n99), .B(n98), .Y(n149));
NAND2X1  g068(.A(n88), .B(G9), .Y(n150));
NOR3X1   g069(.A(G11), .B(G8), .C(G7), .Y(n151));
INVX1    g070(.A(n151), .Y(n152));
OAI21X1  g071(.A0(n152), .A1(n150), .B0(n149), .Y(n153));
NOR4X1   g072(.A(n91), .B(n146), .C(n133), .D(n100), .Y(n154));
NAND2X1  g073(.A(n154), .B(n153), .Y(n155));
AND2X1   g074(.A(n155), .B(n148), .Y(n156));
AND2X1   g075(.A(G10), .B(G7), .Y(n157));
AND2X1   g076(.A(n157), .B(n98), .Y(n158));
NAND2X1  g077(.A(G8), .B(n86), .Y(n159));
OAI22X1  g078(.A0(n150), .A1(n86), .B0(n113), .B1(n159), .Y(n160));
XOR2X1   g079(.A(G3), .B(G2), .Y(n161));
AOI21X1  g080(.A0(n91), .A1(G4), .B0(n161), .Y(n162));
OR2X1    g081(.A(n162), .B(n87_1), .Y(n163));
AND2X1   g082(.A(G6), .B(G4), .Y(n164));
OAI21X1  g083(.A0(n164), .A1(n84), .B0(n141_1), .Y(n165));
AOI22X1  g084(.A0(n106), .A1(n84), .B0(G5), .B1(n165), .Y(n166));
AOI21X1  g085(.A0(n166), .A1(n163), .B0(n133), .Y(n167));
OAI21X1  g086(.A0(n87_1), .A1(G4), .B0(n85), .Y(n168));
NOR2X1   g087(.A(n146), .B(G1), .Y(n169));
NAND2X1  g088(.A(n169), .B(n168), .Y(n170));
AND2X1   g089(.A(G4), .B(G1), .Y(n171));
NAND3X1  g090(.A(n171), .B(n87_1), .C(G2), .Y(n172));
NAND2X1  g091(.A(n172), .B(n170), .Y(n173));
OAI22X1  g092(.A0(n167), .A1(n173), .B0(n160), .B1(n158), .Y(n174));
NOR2X1   g093(.A(n83), .B(G12), .Y(n175));
AND2X1   g094(.A(n175), .B(n174), .Y(n176));
NAND2X1  g095(.A(G36), .B(n87_1), .Y(n177));
NOR4X1   g096(.A(n115), .B(G8), .C(G7), .D(n88), .Y(n178));
NOR4X1   g097(.A(G9), .B(n112_1), .C(n86), .D(G10), .Y(n179));
NOR3X1   g098(.A(n100), .B(n126), .C(n85), .Y(n180));
OAI21X1  g099(.A0(n179), .A1(n178), .B0(n180), .Y(n181));
AOI21X1  g100(.A0(n181), .A1(n177), .B0(G3), .Y(n182));
NAND2X1  g101(.A(n182), .B(n146), .Y(n183));
NOR2X1   g102(.A(n179), .B(n178), .Y(n184));
OAI21X1  g103(.A0(n159), .A1(n150), .B0(n184), .Y(n185));
NOR4X1   g104(.A(n126), .B(G5), .C(G2), .D(n135), .Y(n186));
NAND4X1  g105(.A(n88), .B(G9), .C(G5), .D(n151), .Y(n187));
NOR2X1   g106(.A(n187), .B(n135), .Y(n188));
NAND2X1  g107(.A(G35), .B(G3), .Y(n189));
OR4X1    g108(.A(n126), .B(G5), .C(G4), .D(n189), .Y(n190));
NAND2X1  g109(.A(n190), .B(n101), .Y(n191));
OR2X1    g110(.A(n191), .B(n188), .Y(n192));
AOI22X1  g111(.A0(n186), .A1(n185), .B0(G2), .B1(n192), .Y(n193));
AND2X1   g112(.A(n193), .B(n183), .Y(n194));
INVX1    g113(.A(G32), .Y(n195));
NOR2X1   g114(.A(n160), .B(n158), .Y(n196));
OAI21X1  g115(.A0(n196), .A1(n195), .B0(n83), .Y(n197));
NOR2X1   g116(.A(n197), .B(G12), .Y(n198));
AOI22X1  g117(.A0(n194), .A1(n198), .B0(n176), .B1(n156), .Y(n199));
NAND2X1  g118(.A(n199), .B(n132_1), .Y(G539));
NOR3X1   g119(.A(n174), .B(n171), .C(n85), .Y(n201));
INVX1    g120(.A(n171), .Y(n202));
NOR3X1   g121(.A(n174), .B(n202), .C(G5), .Y(n203));
NOR2X1   g122(.A(n203), .B(n201), .Y(n204));
INVX1    g123(.A(G12), .Y(n205));
NAND3X1  g124(.A(G13), .B(n205), .C(G2), .Y(n206));
NAND3X1  g125(.A(n171), .B(G3), .C(n97_1), .Y(n207));
OAI21X1  g126(.A0(G29), .A1(n97_1), .B0(n207), .Y(n208));
OR4X1    g127(.A(n111), .B(G13), .C(n205), .D(n130), .Y(n209));
INVX1    g128(.A(n209), .Y(n210));
NOR2X1   g129(.A(G33), .B(G13), .Y(n211));
NAND2X1  g130(.A(n211), .B(G3), .Y(n212));
NOR4X1   g131(.A(n195), .B(G13), .C(G12), .D(n196), .Y(n213));
INVX1    g132(.A(n213), .Y(n214));
OAI21X1  g133(.A0(n105), .A1(n146), .B0(n107_1), .Y(n215));
OAI21X1  g134(.A0(n215), .A1(n214), .B0(n212), .Y(n216));
AOI21X1  g135(.A0(n210), .A1(n208), .B0(n216), .Y(n217));
OAI21X1  g136(.A0(n206), .A1(n204), .B0(n217), .Y(G550));
INVX1    g137(.A(n175), .Y(n219));
NOR4X1   g138(.A(n202), .B(n84), .C(G2), .D(n174), .Y(n220));
NOR4X1   g139(.A(n105), .B(n146), .C(G1), .D(n174), .Y(n221));
NOR4X1   g140(.A(G5), .B(n84), .C(G2), .D(n87_1), .Y(n222));
OAI22X1  g141(.A0(G5), .A1(n105), .B0(G3), .B1(n100), .Y(n223));
NOR2X1   g142(.A(n223), .B(n222), .Y(n224));
NOR3X1   g143(.A(n224), .B(n174), .C(n133), .Y(n225));
NOR3X1   g144(.A(n225), .B(n221), .C(n220), .Y(n226));
AND2X1   g145(.A(G39), .B(G4), .Y(n227));
AND2X1   g146(.A(G2), .B(G0), .Y(n228));
MX2X1    g147(.A(G1), .B(G4), .S0(n228), .Y(n229));
AND2X1   g148(.A(G3), .B(G0), .Y(n230));
MX2X1    g149(.A(n230), .B(n97_1), .S0(n171), .Y(n231));
AOI21X1  g150(.A0(n229), .A1(n84), .B0(n231), .Y(n232));
NOR3X1   g151(.A(n232), .B(n209), .C(n85), .Y(n233));
AOI21X1  g152(.A0(n227), .A1(n213), .B0(n233), .Y(n234));
OAI21X1  g153(.A0(n226), .A1(n219), .B0(n234), .Y(G551));
NAND3X1  g154(.A(G6), .B(G3), .C(n146), .Y(n236));
XOR2X1   g155(.A(G5), .B(G4), .Y(n237));
AOI22X1  g156(.A0(n164), .A1(n84), .B0(G6), .B1(n237), .Y(n238));
OAI22X1  g157(.A0(n236), .A1(n106), .B0(n146), .B1(n238), .Y(n239));
NAND2X1  g158(.A(G5), .B(G2), .Y(n240));
OAI21X1  g159(.A0(n171), .A1(n146), .B0(n91), .Y(n241));
AOI22X1  g160(.A0(n240), .A1(n164), .B0(G6), .B1(n241), .Y(n242));
NOR3X1   g161(.A(n242), .B(n219), .C(n174), .Y(n243));
AOI21X1  g162(.A0(n239), .A1(n213), .B0(n243), .Y(n244));
OAI21X1  g163(.A0(n209), .A1(G40), .B0(n244), .Y(G552));
XOR2X1   g164(.A(n116), .B(G7), .Y(n246));
NAND3X1  g165(.A(n246), .B(G34), .C(G9), .Y(n247));
NOR3X1   g166(.A(n99), .B(n115), .C(G6), .Y(n248));
MX2X1    g167(.A(n115), .B(n126), .S0(n88), .Y(n249));
AND2X1   g168(.A(G11), .B(G9), .Y(n250));
INVX1    g169(.A(n150), .Y(n251));
AOI22X1  g170(.A0(n251), .A1(n159), .B0(n250), .B1(n112_1), .Y(n252));
OAI21X1  g171(.A0(n249), .A1(n159), .B0(n252), .Y(n253));
AOI21X1  g172(.A0(n253), .A1(G6), .B0(n248), .Y(n254));
OAI21X1  g173(.A0(n254), .A1(n209), .B0(n247), .Y(G547));
INVX1    g174(.A(G34), .Y(n256));
NOR4X1   g175(.A(n126), .B(n115), .C(n86), .D(n116), .Y(n257));
OAI22X1  g176(.A0(n251), .A1(n159), .B0(n99), .B1(G9), .Y(n258));
AOI21X1  g177(.A0(n258), .A1(G11), .B0(n257), .Y(n259));
OAI22X1  g178(.A0(n209), .A1(G42), .B0(n256), .B1(n259), .Y(G548));
OR4X1    g179(.A(n209), .B(n105), .C(n133), .D(n230), .Y(n261));
NOR2X1   g180(.A(n173), .B(n167), .Y(n262));
MX2X1    g181(.A(G2), .B(n100), .S0(n84), .Y(n263));
OAI21X1  g182(.A0(G3), .A1(n146), .B0(n85), .Y(n264));
NOR3X1   g183(.A(G5), .B(n105), .C(n146), .Y(n265));
AOI21X1  g184(.A0(n264), .A1(n105), .B0(n265), .Y(n266));
OAI21X1  g185(.A0(n263), .A1(n85), .B0(n266), .Y(n267));
NAND2X1  g186(.A(n267), .B(n175), .Y(n268));
OR4X1    g187(.A(n262), .B(n196), .C(n133), .D(n268), .Y(n269));
NAND2X1  g188(.A(G4), .B(G3), .Y(n270));
NAND4X1  g189(.A(n213), .B(G5), .C(G2), .D(n270), .Y(n271));
NAND4X1  g190(.A(n269), .B(n261), .C(n212), .D(n271), .Y(G549));
NOR3X1   g191(.A(n130), .B(n111), .C(n205), .Y(n273));
AND2X1   g192(.A(G3), .B(G1), .Y(n274));
INVX1    g193(.A(n274), .Y(n275));
OAI22X1  g194(.A0(n91), .A1(G4), .B0(G5), .B1(n275), .Y(n276));
OR2X1    g195(.A(n276), .B(n108), .Y(n277));
MX2X1    g196(.A(G1), .B(n277), .S0(G0), .Y(n278));
NAND4X1  g197(.A(n273), .B(n83), .C(G2), .D(n278), .Y(n279));
AOI21X1  g198(.A0(n193), .A1(n183), .B0(n197), .Y(n280));
NAND3X1  g199(.A(n280), .B(n182), .C(n205), .Y(n281));
NAND2X1  g200(.A(n281), .B(n279), .Y(G530));
NOR3X1   g201(.A(G10), .B(n115), .C(n86), .Y(n283));
OAI22X1  g202(.A0(n256), .A1(n112_1), .B0(n87_1), .B1(n209), .Y(n284));
NAND2X1  g203(.A(n284), .B(n283), .Y(n285));
NOR2X1   g204(.A(n209), .B(n87_1), .Y(n286));
AOI21X1  g205(.A0(G9), .A1(G8), .B0(n256), .Y(n287));
INVX1    g206(.A(n137_1), .Y(n288));
OAI21X1  g207(.A0(G8), .A1(n86), .B0(n88), .Y(n289));
NAND2X1  g208(.A(n289), .B(n115), .Y(n290));
OAI21X1  g209(.A0(n115), .A1(n86), .B0(n116), .Y(n291));
NAND3X1  g210(.A(n291), .B(n290), .C(n288), .Y(n292));
AOI22X1  g211(.A0(n287), .A1(n157), .B0(n286), .B1(n292), .Y(n293));
NAND2X1  g212(.A(n293), .B(n285), .Y(G542));
OR2X1    g213(.A(n274), .B(n146), .Y(n295));
NOR2X1   g214(.A(G5), .B(G3), .Y(n296));
AOI21X1  g215(.A0(n107_1), .A1(n146), .B0(n296), .Y(n297));
AOI21X1  g216(.A0(n297), .A1(n295), .B0(n105), .Y(n298));
OR2X1    g217(.A(G3), .B(G2), .Y(n299));
OAI22X1  g218(.A0(n275), .A1(G4), .B0(n133), .B1(n299), .Y(n300));
OAI21X1  g219(.A0(n300), .A1(n298), .B0(G0), .Y(n301));
NAND2X1  g220(.A(n155), .B(n148), .Y(n302));
NAND2X1  g221(.A(n302), .B(G13), .Y(n303));
INVX1    g222(.A(n135), .Y(n304));
NAND2X1  g223(.A(n280), .B(n304), .Y(n305));
AOI21X1  g224(.A0(n305), .A1(n303), .B0(n288), .Y(n306));
AOI21X1  g225(.A0(n155), .A1(n148), .B0(n83), .Y(n307));
NOR2X1   g226(.A(n307), .B(n280), .Y(n308));
OAI21X1  g227(.A0(n184), .A1(G4), .B0(n187), .Y(n309));
NAND2X1  g228(.A(n309), .B(G6), .Y(n310));
OR4X1    g229(.A(n87_1), .B(n85), .C(n105), .D(n144), .Y(n311));
AOI21X1  g230(.A0(n311), .A1(n141_1), .B0(G3), .Y(n312));
NOR3X1   g231(.A(n174), .B(G43), .C(n83), .Y(n313));
AOI21X1  g232(.A0(n312), .A1(n280), .B0(n313), .Y(n314));
OAI21X1  g233(.A0(n310), .A1(n308), .B0(n314), .Y(n315));
OAI21X1  g234(.A0(n315), .A1(n306), .B0(n205), .Y(n316));
OAI21X1  g235(.A0(n301), .A1(n209), .B0(n316), .Y(G532));
INVX1    g236(.A(n106), .Y(n318));
OAI21X1  g237(.A0(G9), .A1(G7), .B0(n88), .Y(n319));
NOR4X1   g238(.A(n156), .B(n318), .C(n83), .D(n319), .Y(n320));
NOR3X1   g239(.A(n308), .B(n184), .C(G4), .Y(n321));
NOR2X1   g240(.A(n321), .B(n320), .Y(n322));
NAND2X1  g241(.A(n205), .B(G6), .Y(n323));
AND2X1   g242(.A(n280), .B(n205), .Y(n324));
NAND3X1  g243(.A(n131), .B(n83), .C(G12), .Y(n325));
NOR4X1   g244(.A(n104), .B(n91), .C(n133), .D(n325), .Y(n326));
AND2X1   g245(.A(G38), .B(G37), .Y(n327));
NAND4X1  g246(.A(G11), .B(n85), .C(G3), .D(n164), .Y(n328));
OAI22X1  g247(.A0(n328), .A1(n319), .B0(G44), .B1(G3), .Y(n329));
AOI22X1  g248(.A0(n327), .A1(n326), .B0(n324), .B1(n329), .Y(n330));
OAI21X1  g249(.A0(n323), .A1(n322), .B0(n330), .Y(G535));
NOR4X1   g250(.A(G9), .B(n86), .C(n87_1), .D(G10), .Y(n332));
OAI21X1  g251(.A0(n332), .A1(n107_1), .B0(G8), .Y(n333));
OAI21X1  g252(.A0(n179), .A1(n178), .B0(n304), .Y(n334));
OAI22X1  g253(.A0(n333), .A1(n308), .B0(n303), .B1(n334), .Y(n335));
NAND3X1  g254(.A(G38), .B(n115), .C(G6), .Y(n336));
NAND2X1  g255(.A(n336), .B(n99), .Y(n337));
AOI22X1  g256(.A0(n335), .A1(n205), .B0(n326), .B1(n337), .Y(n338));
INVX1    g257(.A(n334), .Y(n339));
NOR3X1   g258(.A(G6), .B(G5), .C(G4), .Y(n340));
NAND3X1  g259(.A(n340), .B(n126), .C(n88), .Y(n341));
NAND4X1  g260(.A(n250), .B(G10), .C(G5), .D(n164), .Y(n342));
AOI21X1  g261(.A0(n342), .A1(n341), .B0(n119), .Y(n343));
NOR4X1   g262(.A(n99), .B(n98), .C(G6), .D(n318), .Y(n344));
NOR3X1   g263(.A(n344), .B(n343), .C(n339), .Y(n345));
OR4X1    g264(.A(n197), .B(n194), .C(G12), .D(n345), .Y(n346));
OAI21X1  g265(.A0(n338), .A1(n146), .B0(n346), .Y(G537));
NOR2X1   g266(.A(n84), .B(G2), .Y(n348));
MX2X1    g267(.A(G5), .B(G3), .S0(G4), .Y(n349));
AOI22X1  g268(.A0(n169), .A1(n349), .B0(n348), .B1(n318), .Y(n57));
OAI21X1  g269(.A0(n126), .A1(G9), .B0(n88), .Y(n62));
OAI22X1  g270(.A0(n126), .A1(G7), .B0(n88), .B1(n250), .Y(n67));
AOI21X1  g271(.A0(n168), .A1(n348), .B0(n265), .Y(n353));
OAI21X1  g272(.A0(n240), .A1(n304), .B0(n353), .Y(n72));
NOR3X1   g273(.A(n196), .B(n195), .C(G12), .Y(n355));
NOR3X1   g274(.A(G4), .B(n133), .C(n97_1), .Y(n356));
AOI22X1  g275(.A0(n265), .A1(n355), .B0(n273), .B1(n356), .Y(n77));
MX2X1    g276(.A(n195), .B(n262), .S0(G13), .Y(n358));
NOR3X1   g277(.A(n358), .B(n196), .C(G12), .Y(n82));
OR2X1    g278(.A(G8), .B(G6), .Y(n360));
OR4X1    g279(.A(G10), .B(G9), .C(n86), .D(n360), .Y(n361));
OAI21X1  g280(.A0(n184), .A1(n87_1), .B0(n361), .Y(n87));
OR4X1    g281(.A(G10), .B(G8), .C(G7), .D(G11), .Y(n363));
AOI21X1  g282(.A0(n363), .A1(n149), .B0(G5), .Y(n92));
XOR2X1   g283(.A(G9), .B(G6), .Y(n97));
NOR4X1   g284(.A(n86), .B(G4), .C(G0), .D(G10), .Y(n102));
XOR2X1   g285(.A(n107_1), .B(G2), .Y(n107));
AND2X1   g286(.A(G9), .B(G6), .Y(n368));
AOI22X1  g287(.A0(G30), .A1(n87_1), .B0(n126), .B1(n368), .Y(n369));
OAI22X1  g288(.A0(n127_1), .A1(n87_1), .B0(n86), .B1(n369), .Y(n370));
NOR3X1   g289(.A(n98), .B(G10), .C(n87_1), .Y(n371));
AOI21X1  g290(.A0(n370), .A1(G8), .B0(n371), .Y(n112));
OR2X1    g291(.A(n368), .B(n99), .Y(n373));
OAI22X1  g292(.A0(n291), .A1(n256), .B0(n209), .B1(n373), .Y(n374));
AOI21X1  g293(.A0(n284), .A1(n283), .B0(n374), .Y(n117));
NOR4X1   g294(.A(n126), .B(n115), .C(n87_1), .D(n157), .Y(n376));
NAND3X1  g295(.A(n150), .B(G7), .C(n87_1), .Y(n377));
AOI22X1  g296(.A0(n112_1), .A1(G7), .B0(G6), .B1(n116), .Y(n378));
OAI21X1  g297(.A0(n378), .A1(G9), .B0(n377), .Y(n379));
AOI21X1  g298(.A0(n379), .A1(G11), .B0(n376), .Y(n122));
NAND3X1  g299(.A(n87_1), .B(G4), .C(G2), .Y(n381));
AOI22X1  g300(.A0(n100), .A1(G5), .B0(G6), .B1(n106), .Y(n382));
AOI21X1  g301(.A0(n382), .A1(n381), .B0(n275), .Y(n383));
OAI22X1  g302(.A0(n170), .A1(n84), .B0(n133), .B1(n236), .Y(n384));
NOR2X1   g303(.A(n384), .B(n383), .Y(n127));
NOR4X1   g304(.A(n99), .B(n98), .C(G5), .D(n141_1), .Y(n386));
NAND3X1  g305(.A(n123), .B(n87_1), .C(n85), .Y(n387));
AOI21X1  g306(.A0(n387), .A1(n342), .B0(n119), .Y(n388));
NOR2X1   g307(.A(n388), .B(n386), .Y(n132));
NAND2X1  g308(.A(n176), .B(n302), .Y(n390));
OAI21X1  g309(.A0(n325), .A1(n104), .B0(n390), .Y(n391));
OR2X1    g310(.A(n391), .B(n324), .Y(G45));
NAND2X1  g311(.A(n109), .B(n318), .Y(n393));
AOI21X1  g312(.A0(n348), .A1(n106), .B0(n97_1), .Y(n394));
AOI21X1  g313(.A0(n394), .A1(n393), .B0(G1), .Y(n395));
NOR2X1   g314(.A(n84), .B(G1), .Y(n396));
AOI21X1  g315(.A0(n105), .A1(G3), .B0(n97_1), .Y(n397));
OAI21X1  g316(.A0(n397), .A1(n396), .B0(G2), .Y(n398));
NOR3X1   g317(.A(G30), .B(G10), .C(G6), .Y(n399));
AOI21X1  g318(.A0(n86), .A1(n87_1), .B0(n399), .Y(n400));
OAI21X1  g319(.A0(n398), .A1(n108), .B0(n400), .Y(n401));
NOR2X1   g320(.A(n401), .B(n395), .Y(n141));
endmodule
