// Benchmark "b17_C" written by ABC on Wed Aug 05 14:42:11 2020

module b17_C ( 
    P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
    DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
    DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
    DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
    DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
    DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
    P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
    P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
    P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
    P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
    P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
    P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
    P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
    P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
    P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
    P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
    P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
    P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
    P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
    P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
    P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
    P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
    P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
    P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN,
    P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
    P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN,
    P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
    P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN,
    P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
    P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN,
    P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
    P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN,
    P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
    P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
    P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
    P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
    P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
    P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN,
    P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
    P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN,
    P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
    P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN,
    P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
    P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN,
    P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN,
    P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN,
    P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN,
    P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN,
    P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
    P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
    P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
    P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
    P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
    P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
    P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
    P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
    P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
    P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
    P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
    P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
    P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
    P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
    P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
    P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN,
    P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN,
    P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN,
    P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN,
    P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN,
    P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN,
    P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN,
    P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN,
    P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN,
    P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN,
    P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN,
    P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN,
    P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN,
    P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN,
    P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN,
    P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN,
    P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN,
    P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN,
    P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN,
    P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN,
    P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN,
    P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN,
    P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN,
    P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN,
    P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN,
    P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN,
    P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN,
    P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN,
    P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN,
    P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN,
    P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN,
    P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN,
    P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN,
    P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN,
    P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN,
    P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN,
    P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN,
    P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN,
    P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN,
    P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN,
    P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN,
    P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN,
    P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN,
    P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN,
    P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN,
    P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN,
    P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN,
    P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN,
    P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
    P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
    P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
    P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
    P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
    P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN,
    P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN,
    P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN,
    P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN,
    P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN,
    P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN,
    P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN,
    P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN,
    P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN,
    P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN,
    P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN,
    P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN,
    P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN,
    P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN,
    P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN,
    P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN,
    P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN,
    BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN,
    BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN,
    BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN,
    BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN,
    BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN,
    BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN,
    BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN,
    BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN,
    BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN,
    BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN,
    BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN,
    BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN,
    BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN,
    BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN,
    BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN,
    BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN,
    BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN,
    BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN,
    BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN,
    BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN,
    BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN,
    READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN,
    READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN,
    P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN,
    P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN,
    P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN,
    P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN,
    P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN,
    P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN,
    P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN,
    P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN,
    P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN,
    P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN,
    P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN,
    P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN,
    P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN,
    P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN,
    P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN,
    P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN,
    P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN,
    P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN,
    P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN,
    P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN,
    P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN,
    P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN,
    P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN,
    P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN,
    P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN,
    P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN,
    P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN,
    P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN,
    P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN,
    P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN,
    P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN,
    P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN,
    P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN,
    P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN,
    P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN,
    P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN,
    P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN,
    P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN,
    P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN,
    P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN,
    P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN,
    P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN,
    P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN,
    P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN,
    P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN,
    P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN,
    P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN,
    P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN,
    P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN,
    P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN,
    P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN,
    P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN,
    P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN,
    P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN,
    P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN,
    P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN,
    P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN,
    P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN,
    P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN,
    P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN,
    P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN,
    P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN,
    P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN,
    P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN,
    P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN,
    P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN,
    P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN,
    P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN,
    P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN,
    P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN,
    P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN,
    P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN,
    P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN,
    P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN,
    P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN,
    P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN,
    P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN,
    P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN,
    P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN,
    P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN,
    P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN,
    P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN,
    P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN,
    P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN,
    P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN,
    P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN,
    P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN,
    P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN,
    P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN,
    P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN,
    P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN,
    P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN,
    P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN,
    P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN,
    P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN,
    P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN,
    P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN,
    P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN,
    P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN,
    P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
    P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
    P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
    P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
    P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
    P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
    P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
    P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
    P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
    P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
    P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
    P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN,
    P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN,
    P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN,
    P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN,
    P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN,
    P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN,
    P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN,
    P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN,
    P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN,
    P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN,
    P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
    P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
    P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
    P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
    P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
    P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
    P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
    P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
    P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
    P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
    P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
    P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
    P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
    P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
    P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
    P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
    P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
    P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
    P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
    P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
    P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
    P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
    P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
    P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
    P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
    P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
    P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
    P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
    P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
    P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
    P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
    P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
    P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
    P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
    P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
    P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
    P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
    P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
    P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
    P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
    P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
    P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
    P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
    P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
    P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
    P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
    P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
    P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
    P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
    P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
    P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
    P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
    P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN,
    P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
    P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN,
    P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
    P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN,
    P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
    P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
    P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
    P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
    P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
    P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN,
    P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
    P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN,
    P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
    P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN,
    P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
    P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN,
    P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
    P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN,
    P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
    P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
    P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
    P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
    P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
    P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
    P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
    P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
    P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
    P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
    P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
    P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
    P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
    P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
    P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
    P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
    P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
    P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
    P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
    P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
    P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN,
    P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN,
    P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN,
    P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN,
    P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN,
    P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN,
    P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN,
    P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN,
    P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN,
    P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN,
    P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN,
    P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN,
    P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN,
    P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN,
    P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN,
    P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN,
    P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN,
    P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN,
    P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN,
    P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN,
    P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN,
    P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN,
    P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN,
    P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN,
    P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN,
    P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN,
    P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN,
    P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN,
    P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN,
    P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN,
    P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN,
    P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN,
    P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN,
    P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN,
    P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN,
    P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN,
    P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN,
    P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN,
    P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN,
    P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN,
    P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN,
    P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN,
    P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN,
    P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN,
    P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN,
    P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN,
    P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN,
    P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN,
    P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN,
    P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN,
    P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN,
    P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN,
    P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN,
    P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN,
    P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN,
    P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN,
    P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN,
    P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN,
    P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN,
    P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN,
    P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN,
    P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN,
    P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN,
    P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN,
    P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN,
    P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN,
    P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN,
    P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN,
    P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN,
    P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN,
    P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN,
    P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN,
    P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN,
    P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN,
    P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN,
    P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN,
    P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN,
    P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN,
    P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN,
    P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN,
    P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN,
    P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN,
    P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN,
    P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN,
    P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN,
    P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN,
    P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN,
    P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN,
    P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN,
    P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN,
    P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN,
    P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN,
    P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN,
    P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN,
    P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN,
    P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN,
    P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN,
    P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN,
    P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN,
    P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
    P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
    P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
    P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
    P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
    P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
    P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
    P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
    P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
    P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
    P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
    P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN,
    P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN,
    P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN,
    P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN,
    P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN,
    P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN,
    P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN,
    P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN,
    P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN,
    P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN,
    P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
    P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
    P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
    P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
    P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
    P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
    P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
    P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
    P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
    P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
    P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
    P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
    P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
    P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
    P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
    P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
    P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
    P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
    P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
    P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
    P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
    P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
    P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
    P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
    P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
    P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
    P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
    P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
    P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
    P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
    P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
    P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
    P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
    P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
    P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
    P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
    P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
    P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
    P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
    P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
    P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
    P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
    P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
    P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
    P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
    P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
    P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
    P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
    P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
    P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
    P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
    P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
    P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN,
    P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
    P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN,
    P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
    P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN,
    P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
    P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
    P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
    P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
    P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
    P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN,
    P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
    P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN,
    P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
    P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN,
    P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
    P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN,
    P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
    P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN,
    P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
    P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
    P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
    P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
    P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
    P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
    P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
    P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
    P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
    P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
    P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
    P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
    P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
    P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
    P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
    P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
    P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
    P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
    P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
    P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
    P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN,
    P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN,
    P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN,
    P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN,
    P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN,
    P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN,
    P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN,
    P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN,
    P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN,
    P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN,
    P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN,
    P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN,
    P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN,
    P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN,
    P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN,
    P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN,
    P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN,
    P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN,
    P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN,
    P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN,
    P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN,
    P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN,
    P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN,
    P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN,
    P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN,
    P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN,
    P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN,
    P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN,
    P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN,
    P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN,
    P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN,
    P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN,
    P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN,
    P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN,
    P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN,
    P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN,
    P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN,
    P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN,
    P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN,
    P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN,
    P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN,
    P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN,
    P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN,
    P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN,
    P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN,
    P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN,
    P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN,
    P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN,
    P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN,
    P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN,
    P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN,
    P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN,
    P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN,
    P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN,
    P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN,
    P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN,
    P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN,
    P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN,
    P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN,
    P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN,
    P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN,
    P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN,
    P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN,
    P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN,
    P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN,
    P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN,
    P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN,
    P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN,
    P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN,
    P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN,
    P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN,
    P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN,
    P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN,
    P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN,
    P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN,
    P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN,
    P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN,
    P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN,
    P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN,
    P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN,
    P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN,
    P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN,
    P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN,
    U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367,
    U368, U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350,
    U351, U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242,
    U241, U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230,
    U229, U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218,
    U217, U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260,
    U261, U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272,
    U273, U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215,
    U213, U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060,
    P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053,
    P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046,
    P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039,
    P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032,
    P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027,
    P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020,
    P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013,
    P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006,
    P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999,
    P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993,
    P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986,
    P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979,
    P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972,
    P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965,
    P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958,
    P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951,
    P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944,
    P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937,
    P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930,
    P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923,
    P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916,
    P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909,
    P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902,
    P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895,
    P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888,
    P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881,
    P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874,
    P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284,
    P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865,
    P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858,
    P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851,
    P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844,
    P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837,
    P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830,
    P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823,
    P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816,
    P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809,
    P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802,
    P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795,
    P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788,
    P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781,
    P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774,
    P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767,
    P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760,
    P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753,
    P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746,
    P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739,
    P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732,
    P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725,
    P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718,
    P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711,
    P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704,
    P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697,
    P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690,
    P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683,
    P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676,
    P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669,
    P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662,
    P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655,
    P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648,
    P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641,
    P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637,
    P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633,
    P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241,
    P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
    P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
    P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
    P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213,
    P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208,
    P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201,
    P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194,
    P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187,
    P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180,
    P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174,
    P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167,
    P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160,
    P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153,
    P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146,
    P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139,
    P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132,
    P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125,
    P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118,
    P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111,
    P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104,
    P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097,
    P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090,
    P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083,
    P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076,
    P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069,
    P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062,
    P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055,
    P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048,
    P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602,
    P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043,
    P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036,
    P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029,
    P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022,
    P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015,
    P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008,
    P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001,
    P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994,
    P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987,
    P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980,
    P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973,
    P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966,
    P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959,
    P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952,
    P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945,
    P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938,
    P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931,
    P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924,
    P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917,
    P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910,
    P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903,
    P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896,
    P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889,
    P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882,
    P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875,
    P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868,
    P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861,
    P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854,
    P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847,
    P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840,
    P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833,
    P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826,
    P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608,
    P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816,
    P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461,
    P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220,
    P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213,
    P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206,
    P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199,
    P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465,
    P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187,
    P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180,
    P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173,
    P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166,
    P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160,
    P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153,
    P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146,
    P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139,
    P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132,
    P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125,
    P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118,
    P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111,
    P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104,
    P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097,
    P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090,
    P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083,
    P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076,
    P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069,
    P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062,
    P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055,
    P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048,
    P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041,
    P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034,
    P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032,
    P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029,
    P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022,
    P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015,
    P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008,
    P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001,
    P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994,
    P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987,
    P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980,
    P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973,
    P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966,
    P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959,
    P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952,
    P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945,
    P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938,
    P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931,
    P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924,
    P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917,
    P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910,
    P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903,
    P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896,
    P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889,
    P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882,
    P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875,
    P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868,
    P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861,
    P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854,
    P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847,
    P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840,
    P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833,
    P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826,
    P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819,
    P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812,
    P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482,
    P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486,
    P1_U2803, P1_U2802, P1_U3487, P1_U2801  );
  input  P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_,
    DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_,
    DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_,
    DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_,
    DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_,
    DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
    P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
    P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
    P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
    P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
    P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
    P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
    P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
    P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
    P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
    P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
    P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
    P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
    P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
    P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
    P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
    P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
    P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
    P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN,
    P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
    P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN,
    P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
    P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN,
    P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
    P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN,
    P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
    P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN,
    P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
    P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
    P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
    P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
    P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
    P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN,
    P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
    P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN,
    P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
    P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN,
    P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
    P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN,
    P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN,
    P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN,
    P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN,
    P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN,
    P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
    P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
    P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
    P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
    P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
    P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
    P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
    P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
    P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
    P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
    P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
    P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
    P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
    P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
    P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
    P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN,
    P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN,
    P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN,
    P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN,
    P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN,
    P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN,
    P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN,
    P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN,
    P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN,
    P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN,
    P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN,
    P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN,
    P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN,
    P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN,
    P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN,
    P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN,
    P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN,
    P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN,
    P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN,
    P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN,
    P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN,
    P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN,
    P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN,
    P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN,
    P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN,
    P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN,
    P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN,
    P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN,
    P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN,
    P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN,
    P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN,
    P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN,
    P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN,
    P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN,
    P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN,
    P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN,
    P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN,
    P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN,
    P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN,
    P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN,
    P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN,
    P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN,
    P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN,
    P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN,
    P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN,
    P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN,
    P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN,
    P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN,
    P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
    P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
    P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
    P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
    P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
    P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN,
    P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN,
    P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN,
    P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN,
    P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN,
    P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN,
    P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN,
    P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN,
    P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN,
    P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN,
    P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN,
    P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN,
    P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN,
    P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN,
    P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN,
    P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN,
    P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN,
    BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN,
    BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN,
    BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN,
    BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN,
    BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN,
    BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN,
    BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN,
    BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN,
    BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN,
    BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN,
    BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN,
    BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN,
    BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN,
    BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN,
    BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN,
    BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN,
    BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN,
    BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN,
    BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN,
    BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN,
    BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN,
    READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN,
    READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN,
    P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN,
    P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN,
    P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN,
    P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN,
    P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN,
    P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN,
    P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN,
    P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN,
    P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN,
    P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN,
    P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN,
    P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN,
    P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN,
    P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN,
    P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN,
    P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN,
    P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN,
    P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN,
    P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN,
    P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN,
    P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN,
    P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN,
    P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN,
    P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN,
    P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN,
    P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN,
    P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN,
    P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN,
    P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN,
    P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN,
    P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN,
    P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN,
    P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN,
    P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN,
    P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN,
    P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN,
    P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN,
    P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN,
    P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN,
    P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN,
    P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN,
    P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN,
    P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN,
    P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN,
    P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN,
    P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN,
    P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN,
    P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN,
    P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN,
    P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN,
    P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN,
    P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN,
    P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN,
    P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN,
    P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN,
    P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN,
    P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN,
    P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN,
    P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN,
    P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN,
    P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN,
    P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN,
    P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN,
    P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN,
    P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN,
    P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN,
    P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN,
    P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN,
    P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN,
    P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN,
    P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN,
    P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN,
    P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN,
    P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN,
    P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN,
    P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN,
    P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN,
    P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN,
    P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN,
    P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN,
    P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN,
    P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN,
    P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN,
    P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN,
    P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN,
    P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN,
    P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN,
    P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN,
    P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN,
    P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN,
    P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN,
    P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN,
    P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN,
    P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN,
    P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN,
    P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN,
    P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN,
    P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN,
    P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN,
    P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
    P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
    P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
    P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
    P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
    P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
    P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
    P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
    P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
    P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
    P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
    P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN,
    P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN,
    P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN,
    P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN,
    P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN,
    P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN,
    P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN,
    P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN,
    P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN,
    P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN,
    P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
    P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
    P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
    P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
    P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
    P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
    P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
    P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
    P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
    P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
    P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
    P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
    P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
    P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
    P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
    P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
    P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
    P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
    P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
    P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
    P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
    P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
    P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
    P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
    P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
    P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
    P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
    P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
    P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
    P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
    P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
    P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
    P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
    P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
    P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
    P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
    P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
    P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
    P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
    P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
    P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
    P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
    P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
    P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
    P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
    P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
    P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
    P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
    P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
    P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
    P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
    P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
    P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN,
    P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
    P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN,
    P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
    P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN,
    P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
    P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
    P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
    P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
    P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
    P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN,
    P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
    P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN,
    P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
    P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN,
    P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
    P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN,
    P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
    P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN,
    P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
    P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
    P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
    P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
    P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
    P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
    P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
    P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
    P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
    P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
    P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
    P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
    P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
    P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
    P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
    P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
    P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
    P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
    P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
    P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
    P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN,
    P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN,
    P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN,
    P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN,
    P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN,
    P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN,
    P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN,
    P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN,
    P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN,
    P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN,
    P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN,
    P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN,
    P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN,
    P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN,
    P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN,
    P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN,
    P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN,
    P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN,
    P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN,
    P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN,
    P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN,
    P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN,
    P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN,
    P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN,
    P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN,
    P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN,
    P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN,
    P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN,
    P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN,
    P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN,
    P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN,
    P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN,
    P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN,
    P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN,
    P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN,
    P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN,
    P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN,
    P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN,
    P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN,
    P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN,
    P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN,
    P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN,
    P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN,
    P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN,
    P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN,
    P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN,
    P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN,
    P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN,
    P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN,
    P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN,
    P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN,
    P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN,
    P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN,
    P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN,
    P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN,
    P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN,
    P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN,
    P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN,
    P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN,
    P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN,
    P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN,
    P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN,
    P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN,
    P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN,
    P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN,
    P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN,
    P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN,
    P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN,
    P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN,
    P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN,
    P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN,
    P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN,
    P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN,
    P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN,
    P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN,
    P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN,
    P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN,
    P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN,
    P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN,
    P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN,
    P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN,
    P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN,
    P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN,
    P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN,
    P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN,
    P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN,
    P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN,
    P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN,
    P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN,
    P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN,
    P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN,
    P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN,
    P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN,
    P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN,
    P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN,
    P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN,
    P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN,
    P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN,
    P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN,
    P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
    P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
    P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
    P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
    P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
    P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
    P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
    P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
    P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
    P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
    P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
    P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN,
    P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN,
    P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN,
    P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN,
    P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN,
    P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN,
    P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN,
    P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN,
    P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN,
    P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN,
    P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
    P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
    P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
    P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
    P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
    P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
    P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
    P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
    P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
    P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
    P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
    P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
    P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
    P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
    P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
    P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
    P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
    P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
    P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
    P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
    P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
    P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
    P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
    P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
    P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
    P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
    P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
    P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
    P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
    P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
    P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
    P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
    P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
    P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
    P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
    P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
    P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
    P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
    P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
    P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
    P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
    P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
    P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
    P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
    P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
    P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
    P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
    P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
    P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
    P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
    P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
    P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
    P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN,
    P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
    P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN,
    P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
    P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN,
    P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
    P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
    P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
    P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
    P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
    P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN,
    P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
    P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN,
    P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
    P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN,
    P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
    P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN,
    P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
    P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN,
    P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
    P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
    P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
    P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
    P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
    P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
    P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
    P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
    P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
    P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
    P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
    P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
    P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
    P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
    P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
    P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
    P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
    P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
    P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
    P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
    P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN,
    P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN,
    P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN,
    P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN,
    P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN,
    P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN,
    P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN,
    P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN,
    P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN,
    P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN,
    P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN,
    P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN,
    P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN,
    P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN,
    P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN,
    P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN,
    P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN,
    P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN,
    P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN,
    P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN,
    P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN,
    P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN,
    P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN,
    P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN,
    P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN,
    P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN,
    P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN,
    P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN,
    P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN,
    P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN,
    P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN,
    P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN,
    P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN,
    P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN,
    P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN,
    P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN,
    P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN,
    P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN,
    P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN,
    P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN,
    P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN,
    P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN,
    P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN,
    P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN,
    P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN,
    P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN,
    P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN,
    P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN,
    P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN,
    P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN,
    P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN,
    P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN,
    P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN,
    P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN,
    P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN,
    P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN,
    P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN,
    P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN,
    P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN,
    P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN,
    P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN,
    P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN,
    P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN,
    P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN,
    P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN,
    P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN,
    P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN,
    P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN,
    P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN,
    P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN,
    P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN,
    P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN,
    P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN,
    P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN,
    P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN,
    P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN,
    P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN,
    P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN,
    P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN,
    P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN,
    P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN,
    P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN,
    P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
    U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348, U349,
    U350, U351, U352, U353, U354, U365, U376, U247, U246, U245, U244, U243,
    U242, U241, U240, U239, U238, U237, U236, U235, U234, U233, U232, U231,
    U230, U229, U228, U227, U226, U225, U224, U223, U222, U221, U220, U219,
    U218, U217, U216, U251, U252, U253, U254, U255, U256, U257, U258, U259,
    U260, U261, U262, U263, U264, U265, U266, U267, U268, U269, U270, U271,
    U272, U273, U274, U275, U276, U277, U278, U279, U280, U281, U282, U212,
    U215, U213, U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061,
    P3_U3060, P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054,
    P3_U3053, P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047,
    P3_U3046, P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040,
    P3_U3039, P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033,
    P3_U3032, P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028,
    P3_U3027, P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021,
    P3_U3020, P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014,
    P3_U3013, P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007,
    P3_U3006, P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000,
    P3_U2999, P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994,
    P3_U2993, P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987,
    P3_U2986, P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980,
    P3_U2979, P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973,
    P3_U2972, P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966,
    P3_U2965, P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959,
    P3_U2958, P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952,
    P3_U2951, P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945,
    P3_U2944, P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938,
    P3_U2937, P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931,
    P3_U2930, P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924,
    P3_U2923, P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917,
    P3_U2916, P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910,
    P3_U2909, P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903,
    P3_U2902, P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896,
    P3_U2895, P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889,
    P3_U2888, P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882,
    P3_U2881, P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875,
    P3_U2874, P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868,
    P3_U3284, P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866,
    P3_U2865, P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859,
    P3_U2858, P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852,
    P3_U2851, P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845,
    P3_U2844, P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838,
    P3_U2837, P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831,
    P3_U2830, P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824,
    P3_U2823, P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817,
    P3_U2816, P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810,
    P3_U2809, P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803,
    P3_U2802, P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796,
    P3_U2795, P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789,
    P3_U2788, P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782,
    P3_U2781, P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775,
    P3_U2774, P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768,
    P3_U2767, P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761,
    P3_U2760, P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754,
    P3_U2753, P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747,
    P3_U2746, P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740,
    P3_U2739, P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733,
    P3_U2732, P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726,
    P3_U2725, P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719,
    P3_U2718, P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712,
    P3_U2711, P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705,
    P3_U2704, P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698,
    P3_U2697, P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691,
    P3_U2690, P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684,
    P3_U2683, P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677,
    P3_U2676, P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670,
    P3_U2669, P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663,
    P3_U2662, P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656,
    P3_U2655, P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649,
    P3_U2648, P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642,
    P3_U2641, P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294,
    P3_U2637, P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634,
    P3_U2633, P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588,
    P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
    P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
    P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
    P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214,
    P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592,
    P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202,
    P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195,
    P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188,
    P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181,
    P2_U3180, P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175,
    P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168,
    P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161,
    P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154,
    P2_U3153, P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147,
    P2_U3146, P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140,
    P2_U3139, P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133,
    P2_U3132, P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126,
    P2_U3125, P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119,
    P2_U3118, P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112,
    P2_U3111, P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105,
    P2_U3104, P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098,
    P2_U3097, P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091,
    P2_U3090, P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084,
    P2_U3083, P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077,
    P2_U3076, P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070,
    P2_U3069, P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063,
    P2_U3062, P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056,
    P2_U3055, P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049,
    P2_U3048, P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047,
    P2_U3602, P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044,
    P2_U3043, P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037,
    P2_U3036, P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030,
    P2_U3029, P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023,
    P2_U3022, P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016,
    P2_U3015, P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009,
    P2_U3008, P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002,
    P2_U3001, P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995,
    P2_U2994, P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988,
    P2_U2987, P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981,
    P2_U2980, P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974,
    P2_U2973, P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967,
    P2_U2966, P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960,
    P2_U2959, P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953,
    P2_U2952, P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946,
    P2_U2945, P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939,
    P2_U2938, P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932,
    P2_U2931, P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925,
    P2_U2924, P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918,
    P2_U2917, P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911,
    P2_U2910, P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904,
    P2_U2903, P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897,
    P2_U2896, P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890,
    P2_U2889, P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883,
    P2_U2882, P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876,
    P2_U2875, P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869,
    P2_U2868, P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862,
    P2_U2861, P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855,
    P2_U2854, P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848,
    P2_U2847, P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841,
    P2_U2840, P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834,
    P2_U2833, P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827,
    P2_U2826, P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820,
    P2_U3608, P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611,
    P2_U2816, P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460,
    P1_U3461, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221,
    P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214,
    P1_U3213, P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207,
    P1_U3206, P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200,
    P1_U3199, P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464,
    P1_U3465, P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188,
    P1_U3187, P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181,
    P1_U3180, P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174,
    P1_U3173, P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167,
    P1_U3166, P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161,
    P1_U3160, P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154,
    P1_U3153, P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147,
    P1_U3146, P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140,
    P1_U3139, P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133,
    P1_U3132, P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126,
    P1_U3125, P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119,
    P1_U3118, P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112,
    P1_U3111, P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105,
    P1_U3104, P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098,
    P1_U3097, P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091,
    P1_U3090, P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084,
    P1_U3083, P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077,
    P1_U3076, P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070,
    P1_U3069, P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063,
    P1_U3062, P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056,
    P1_U3055, P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049,
    P1_U3048, P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042,
    P1_U3041, P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035,
    P1_U3034, P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474,
    P1_U3032, P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030,
    P1_U3029, P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023,
    P1_U3022, P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016,
    P1_U3015, P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009,
    P1_U3008, P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002,
    P1_U3001, P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995,
    P1_U2994, P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988,
    P1_U2987, P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981,
    P1_U2980, P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974,
    P1_U2973, P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967,
    P1_U2966, P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960,
    P1_U2959, P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953,
    P1_U2952, P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946,
    P1_U2945, P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939,
    P1_U2938, P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932,
    P1_U2931, P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925,
    P1_U2924, P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918,
    P1_U2917, P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911,
    P1_U2910, P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904,
    P1_U2903, P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897,
    P1_U2896, P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890,
    P1_U2889, P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883,
    P1_U2882, P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876,
    P1_U2875, P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869,
    P1_U2868, P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862,
    P1_U2861, P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855,
    P1_U2854, P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848,
    P1_U2847, P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841,
    P1_U2840, P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834,
    P1_U2833, P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827,
    P1_U2826, P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820,
    P1_U2819, P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813,
    P1_U2812, P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807,
    P1_U3482, P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804,
    P1_U3486, P1_U2803, P1_U2802, P1_U3487, P1_U2801;
  wire n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2973, n2974,
    n2976, n2977, n2979, n2980, n2982, n2983, n2985, n2986, n2988, n2989,
    n2991, n2992, n2994, n2995, n2997, n2998, n3000, n3001, n3003, n3004,
    n3006, n3007, n3009, n3010, n3012, n3013, n3015, n3016, n3018, n3019,
    n3021, n3022, n3024, n3025, n3027, n3028, n3030, n3031, n3033, n3034,
    n3036, n3037, n3039, n3040, n3042, n3043, n3045, n3046, n3048, n3049,
    n3051, n3052, n3054, n3055, n3057, n3058, n3060, n3061, n3062, n3063,
    n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
    n3074, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
    n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
    n3095, n3097, n3098, n3100, n3101, n3103, n3104, n3106, n3107, n3109,
    n3110, n3112, n3113, n3115, n3116, n3118, n3119, n3121, n3122, n3124,
    n3125, n3127, n3128, n3130, n3131, n3133, n3134, n3136, n3137, n3139,
    n3140, n3142, n3143, n3145, n3146, n3148, n3149, n3151, n3152, n3154,
    n3155, n3157, n3158, n3160, n3161, n3163, n3164, n3166, n3167, n3169,
    n3170, n3172, n3173, n3175, n3176, n3178, n3179, n3181, n3182, n3184,
    n3185, n3187, n3188, n3190, n3191, n3192, n3194, n3195, n3197, n3198,
    n3200, n3201, n3203, n3204, n3206, n3207, n3209, n3210, n3212, n3213,
    n3215, n3216, n3218, n3219, n3221, n3222, n3224, n3225, n3227, n3228,
    n3230, n3231, n3233, n3234, n3236, n3237, n3239, n3240, n3242, n3243,
    n3245, n3246, n3248, n3249, n3251, n3252, n3254, n3255, n3257, n3258,
    n3260, n3261, n3263, n3264, n3266, n3267, n3269, n3270, n3272, n3273,
    n3275, n3276, n3278, n3279, n3281, n3282, n3284, n3285, n3287, n3290,
    n3291, n3292, n3294, n3295, n3296, n3297, n3299, n3300, n3301, n3302,
    n3304, n3305, n3307, n3308, n3310, n3311, n3312, n3313, n3315, n3316,
    n3318, n3319, n3321, n3322, n3324, n3325, n3327, n3328, n3330, n3331,
    n3333, n3334, n3336, n3337, n3339, n3340, n3342, n3343, n3345, n3346,
    n3348, n3349, n3351, n3352, n3354, n3355, n3357, n3358, n3360, n3361,
    n3363, n3364, n3366, n3367, n3369, n3370, n3372, n3373, n3375, n3376,
    n3378, n3379, n3381, n3382, n3384, n3385, n3387, n3388, n3390, n3391,
    n3393, n3394, n3396, n3397, n3399, n3400, n3402, n3403, n3404, n3405,
    n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
    n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3424, n3425, n3426,
    n3427, n3428, n3429, n3430, n3431, n3432, n3434, n3435, n3436, n3437,
    n3439, n3440, n3441, n3442, n3443, n3445, n3446, n3447, n3449, n3451,
    n3453, n3455, n3457, n3459, n3461, n3463, n3465, n3467, n3469, n3471,
    n3473, n3475, n3477, n3479, n3481, n3483, n3485, n3487, n3489, n3491,
    n3493, n3495, n3497, n3499, n3501, n3503, n3505, n3507, n3509, n3510,
    n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
    n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
    n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
    n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3549, n3550, n3551,
    n3552, n3553, n3554, n3555, n3557, n3559, n3560, n3561, n3562, n3563,
    n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
    n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
    n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
    n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
    n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
    n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
    n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
    n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
    n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
    n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
    n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
    n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
    n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
    n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
    n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
    n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
    n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
    n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
    n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
    n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
    n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
    n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
    n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
    n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
    n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
    n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
    n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
    n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
    n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
    n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
    n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
    n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
    n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
    n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
    n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
    n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
    n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
    n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3943, n3944,
    n3945, n3946, n3947, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
    n3956, n3958, n3959, n3960, n3961, n3962, n3963, n3965, n3966, n3967,
    n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977,
    n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3987, n3988,
    n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
    n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
    n4009, n4010, n4011, n4013, n4014, n4015, n4016, n4017, n4018, n4020,
    n4021, n4022, n4023, n4024, n4025, n4027, n4028, n4029, n4030, n4031,
    n4032, n4034, n4035, n4036, n4037, n4038, n4039, n4041, n4042, n4043,
    n4044, n4045, n4046, n4048, n4049, n4050, n4051, n4052, n4053, n4055,
    n4056, n4057, n4058, n4059, n4060, n4062, n4063, n4065, n4066, n4068,
    n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
    n4079, n4080, n4081, n4082, n4083, n4085, n4086, n4087, n4088, n4089,
    n4090, n4091, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4101,
    n4102, n4103, n4104, n4105, n4106, n4107, n4109, n4110, n4111, n4112,
    n4113, n4114, n4115, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
    n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4133, n4134, n4135,
    n4136, n4137, n4138, n4139, n4142, n4143, n4144, n4145, n4146, n4147,
    n4148, n4149, n4150, n4151, n4152, n4153, n4156, n4158, n4159, n4160,
    n4161, n4163, n4164, n4165, n4166, n4168, n4169, n4170, n4171, n4173,
    n4174, n4175, n4176, n4178, n4179, n4180, n4181, n4183, n4184, n4185,
    n4186, n4188, n4189, n4190, n4191, n4193, n4194, n4195, n4196, n4197,
    n4199, n4200, n4201, n4203, n4204, n4205, n4207, n4208, n4209, n4210,
    n4211, n4212, n4214, n4215, n4217, n4218, n4219, n4220, n4221, n4223,
    n4224, n4225, n4226, n4227, n4229, n4230, n4231, n4232, n4233, n4235,
    n4236, n4237, n4238, n4239, n4241, n4242, n4243, n4244, n4245, n4247,
    n4248, n4249, n4250, n4251, n4253, n4254, n4255, n4256, n4257, n4260,
    n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270,
    n4273, n4275, n4276, n4277, n4278, n4280, n4281, n4282, n4283, n4285,
    n4286, n4287, n4288, n4290, n4291, n4292, n4293, n4295, n4296, n4297,
    n4298, n4300, n4301, n4302, n4303, n4305, n4306, n4307, n4308, n4310,
    n4313, n4314, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
    n4324, n4326, n4327, n4329, n4330, n4331, n4332, n4333, n4335, n4336,
    n4337, n4338, n4339, n4341, n4342, n4343, n4344, n4345, n4347, n4348,
    n4349, n4350, n4351, n4353, n4354, n4355, n4356, n4357, n4359, n4360,
    n4361, n4362, n4363, n4365, n4366, n4367, n4368, n4369, n4372, n4373,
    n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4385,
    n4387, n4388, n4389, n4390, n4392, n4393, n4394, n4395, n4397, n4398,
    n4399, n4400, n4402, n4403, n4404, n4405, n4407, n4408, n4409, n4410,
    n4412, n4413, n4414, n4415, n4417, n4418, n4419, n4420, n4422, n4423,
    n4424, n4425, n4426, n4428, n4429, n4430, n4432, n4433, n4434, n4435,
    n4436, n4437, n4439, n4440, n4442, n4443, n4444, n4445, n4446, n4448,
    n4449, n4450, n4451, n4452, n4454, n4455, n4456, n4457, n4458, n4460,
    n4461, n4462, n4463, n4464, n4466, n4467, n4468, n4469, n4470, n4472,
    n4473, n4474, n4475, n4476, n4478, n4479, n4480, n4481, n4482, n4485,
    n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4497,
    n4499, n4500, n4501, n4502, n4504, n4505, n4506, n4507, n4509, n4510,
    n4511, n4512, n4514, n4515, n4516, n4517, n4519, n4520, n4521, n4522,
    n4524, n4525, n4526, n4527, n4529, n4530, n4531, n4532, n4534, n4537,
    n4538, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
    n4550, n4551, n4553, n4554, n4555, n4556, n4557, n4559, n4560, n4561,
    n4562, n4563, n4565, n4566, n4567, n4568, n4569, n4571, n4572, n4573,
    n4574, n4575, n4577, n4578, n4579, n4580, n4581, n4583, n4584, n4585,
    n4586, n4587, n4589, n4590, n4591, n4592, n4593, n4596, n4597, n4598,
    n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4609, n4611,
    n4612, n4613, n4614, n4616, n4617, n4618, n4619, n4621, n4622, n4623,
    n4624, n4626, n4627, n4628, n4629, n4631, n4632, n4633, n4634, n4636,
    n4637, n4638, n4639, n4641, n4642, n4643, n4644, n4646, n4648, n4649,
    n4650, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
    n4662, n4664, n4665, n4666, n4667, n4668, n4670, n4671, n4672, n4673,
    n4674, n4676, n4677, n4678, n4679, n4680, n4682, n4683, n4684, n4685,
    n4686, n4688, n4689, n4690, n4691, n4692, n4694, n4695, n4696, n4697,
    n4698, n4700, n4701, n4702, n4703, n4704, n4708, n4709, n4710, n4711,
    n4712, n4713, n4714, n4715, n4717, n4718, n4719, n4721, n4722, n4723,
    n4724, n4726, n4727, n4728, n4729, n4731, n4732, n4733, n4734, n4736,
    n4737, n4738, n4739, n4741, n4742, n4743, n4744, n4746, n4747, n4748,
    n4749, n4751, n4752, n4753, n4754, n4757, n4758, n4761, n4762, n4763,
    n4764, n4765, n4766, n4767, n4768, n4769, n4771, n4772, n4773, n4774,
    n4776, n4777, n4778, n4779, n4781, n4782, n4783, n4784, n4786, n4787,
    n4788, n4789, n4791, n4792, n4793, n4794, n4796, n4797, n4798, n4799,
    n4801, n4802, n4803, n4804, n4806, n4809, n4810, n4811, n4812, n4813,
    n4814, n4816, n4817, n4818, n4820, n4821, n4822, n4823, n4825, n4826,
    n4827, n4828, n4830, n4831, n4832, n4833, n4835, n4836, n4837, n4838,
    n4840, n4841, n4842, n4843, n4845, n4846, n4847, n4848, n4850, n4851,
    n4852, n4853, n4855, n4858, n4859, n4861, n4862, n4863, n4864, n4865,
    n4866, n4867, n4868, n4870, n4871, n4872, n4873, n4875, n4876, n4877,
    n4878, n4880, n4881, n4882, n4883, n4885, n4886, n4887, n4888, n4890,
    n4891, n4892, n4893, n4895, n4896, n4897, n4898, n4900, n4901, n4902,
    n4903, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4913, n4914,
    n4915, n4916, n4918, n4919, n4920, n4921, n4922, n4923, n4925, n4926,
    n4927, n4928, n4929, n4931, n4932, n4933, n4935, n4936, n4938, n4939,
    n4940, n4942, n4943, n4944, n4945, n4946, n4947, n4952, n4953, n4954,
    n4955, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4965, n4966,
    n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
    n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4988, n4991,
    n4994, n4997, n4998, n5001, n5004, n5007, n5010, n5011, n5012, n5013,
    n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
    n5024, n5025, n5026, n5027, n5029, n5030, n5031, n5032, n5033, n5034,
    n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
    n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
    n5055, n5056, n5058, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
    n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
    n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
    n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
    n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5106, n5107, n5108,
    n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
    n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5127, n5128, n5129,
    n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5140,
    n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5151,
    n5152, n5153, n5156, n5159, n5162, n5163, n5164, n5165, n5167, n5168,
    n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
    n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
    n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
    n5199, n5200, n5201, n5202, n5203, n5204, n5207, n5213, n5214, n5215,
    n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
    n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
    n5236, n5237, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246,
    n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256,
    n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5266, n5267,
    n5268, n5271, n5272, n5275, n5276, n5281, n5282, n5283, n5284, n5285,
    n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
    n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
    n5306, n5307, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316,
    n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326,
    n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336,
    n5337, n5338, n5339, n5340, n5342, n5343, n5344, n5345, n5346, n5347,
    n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5357, n5358, n5359,
    n5360, n5361, n5362, n5363, n5364, n5366, n5368, n5369, n5370, n5371,
    n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
    n5382, n5383, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
    n5397, n5398, n5399, n5400, n5401, n5404, n5405, n5406, n5407, n5408,
    n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
    n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
    n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5439, n5440,
    n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
    n5451, n5452, n5453, n5455, n5459, n5460, n5461, n5463, n5466, n5467,
    n5468, n5470, n5471, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
    n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
    n5491, n5492, n5493, n5494, n5498, n5499, n5500, n5501, n5502, n5503,
    n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5517,
    n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
    n5528, n5529, n5530, n5531, n5532, n5535, n5536, n5537, n5538, n5539,
    n5540, n5541, n5542, n5543, n5545, n5547, n5548, n5549, n5550, n5551,
    n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
    n5562, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
    n5573, n5574, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
    n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
    n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
    n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5614, n5615, n5616,
    n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5625, n5626, n5627,
    n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
    n5638, n5639, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
    n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5659, n5660,
    n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
    n5671, n5672, n5673, n5674, n5675, n5676, n5679, n5680, n5681, n5682,
    n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
    n5693, n5694, n5695, n5696, n5698, n5699, n5700, n5701, n5702, n5703,
    n5704, n5705, n5706, n5707, n5708, n5709, n5711, n5712, n5713, n5714,
    n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
    n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
    n5737, n5738, n5739, n5740, n5742, n5743, n5744, n5745, n5746, n5747,
    n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
    n5758, n5759, n5760, n5761, n5764, n5765, n5766, n5767, n5768, n5769,
    n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
    n5780, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
    n5791, n5792, n5793, n5794, n5797, n5798, n5799, n5800, n5801, n5802,
    n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
    n5813, n5814, n5815, n5816, n5817, n5818, n5820, n5821, n5822, n5823,
    n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
    n5834, n5835, n5836, n5837, n5838, n5839, n5842, n5843, n5844, n5845,
    n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
    n5856, n5857, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
    n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5877, n5878,
    n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
    n5889, n5890, n5891, n5892, n5894, n5895, n5896, n5897, n5898, n5899,
    n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
    n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5921, n5922,
    n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
    n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5941, n5942, n5943,
    n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
    n5954, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
    n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5976,
    n5977, n5978, n5979, n5980, n5981, n5984, n5985, n5986, n5987, n5988,
    n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
    n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
    n6012, n6013, n6014, n6015, n6016, n6017, n6019, n6020, n6021, n6022,
    n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
    n6033, n6034, n6035, n6036, n6037, n6040, n6041, n6042, n6043, n6044,
    n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
    n6055, n6056, n6057, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
    n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
    n6076, n6077, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
    n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6097, n6098,
    n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
    n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6119, n6120,
    n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
    n6131, n6132, n6133, n6134, n6135, n6136, n6138, n6139, n6140, n6141,
    n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
    n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6163,
    n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
    n6174, n6175, n6176, n6177, n6178, n6180, n6181, n6182, n6183, n6184,
    n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
    n6195, n6196, n6197, n6200, n6201, n6202, n6203, n6204, n6205, n6206,
    n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6217,
    n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227,
    n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237,
    n6238, n6239, n6240, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
    n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6260,
    n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
    n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6281, n6282,
    n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
    n6293, n6294, n6295, n6296, n6298, n6299, n6300, n6301, n6302, n6303,
    n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
    n6314, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
    n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6334, n6335, n6336,
    n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
    n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
    n6357, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
    n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6379,
    n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
    n6390, n6391, n6392, n6393, n6394, n6395, n6398, n6399, n6400, n6401,
    n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
    n6412, n6413, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
    n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
    n6433, n6434, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
    n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6454, n6455,
    n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
    n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
    n6476, n6477, n6478, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
    n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
    n6498, n6499, n6500, n6502, n6503, n6504, n6505, n6507, n6508, n6509,
    n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6518, n6519, n6520,
    n6521, n6522, n6524, n6525, n6526, n6527, n6528, n6529, n6531, n6532,
    n6533, n6534, n6535, n6536, n6537, n6539, n6540, n6541, n6543, n6544,
    n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
    n6555, n6556, n6557, n6558, n6560, n6561, n6562, n6563, n6564, n6565,
    n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6575, n6576,
    n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586,
    n6587, n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597,
    n6598, n6599, n6600, n6601, n6603, n6604, n6605, n6606, n6607, n6608,
    n6609, n6610, n6611, n6612, n6613, n6614, n6616, n6617, n6618, n6619,
    n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6630,
    n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
    n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
    n6652, n6653, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
    n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6671, n6672, n6673,
    n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
    n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
    n6695, n6696, n6697, n6698, n6700, n6701, n6702, n6703, n6704, n6705,
    n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6715, n6716,
    n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6727,
    n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737,
    n6738, n6739, n6740, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
    n6749, n6750, n6751, n6752, n6753, n6754, n6756, n6757, n6758, n6759,
    n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6768, n6769, n6770,
    n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
    n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
    n6792, n6793, n6794, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
    n6803, n6804, n6805, n6806, n6807, n6808, n6810, n6811, n6812, n6813,
    n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
    n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
    n6835, n6836, n6837, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
    n6846, n6847, n6848, n6849, n6850, n6851, n6853, n6854, n6855, n6856,
    n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6867,
    n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877,
    n6878, n6879, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
    n6889, n6890, n6891, n6892, n6893, n6895, n6896, n6897, n6898, n6899,
    n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6909, n6910,
    n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
    n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
    n6932, n6933, n6934, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
    n6944, n6946, n6948, n6950, n6952, n6954, n6956, n6958, n6960, n6962,
    n6964, n6966, n6968, n6970, n6972, n6974, n6976, n6978, n6980, n6982,
    n6984, n6986, n6988, n6990, n6992, n6994, n6996, n6998, n7000, n7002,
    n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7013, n7014,
    n7016, n7017, n7019, n7020, n7022, n7023, n7025, n7026, n7028, n7029,
    n7031, n7032, n7034, n7035, n7037, n7038, n7040, n7041, n7043, n7044,
    n7046, n7047, n7049, n7050, n7052, n7053, n7055, n7056, n7058, n7059,
    n7060, n7062, n7063, n7065, n7066, n7068, n7069, n7071, n7072, n7074,
    n7075, n7077, n7078, n7080, n7081, n7083, n7084, n7086, n7087, n7089,
    n7090, n7092, n7093, n7095, n7096, n7098, n7099, n7101, n7102, n7105,
    n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7114, n7115, n7116,
    n7117, n7119, n7120, n7121, n7122, n7123, n7125, n7126, n7127, n7128,
    n7129, n7131, n7132, n7133, n7134, n7135, n7137, n7138, n7139, n7140,
    n7141, n7143, n7144, n7145, n7146, n7147, n7149, n7150, n7151, n7152,
    n7153, n7154, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
    n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
    n7174, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
    n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
    n7195, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
    n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
    n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7224, n7225, n7226,
    n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236,
    n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246,
    n7247, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257,
    n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267,
    n7268, n7269, n7270, n7271, n7272, n7274, n7275, n7276, n7277, n7278,
    n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
    n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7299,
    n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
    n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
    n7320, n7321, n7322, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
    n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
    n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7349, n7350, n7351,
    n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361,
    n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371,
    n7372, n7378, n7383, n7388, n7393, n7394, n7399, n7404, n7409, n7414,
    n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7425,
    n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
    n7436, n7437, n7438, n7439, n7440, n7441, n7443, n7444, n7445, n7446,
    n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456,
    n7457, n7458, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467,
    n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7477, n7478,
    n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
    n7489, n7490, n7491, n7492, n7494, n7495, n7496, n7497, n7498, n7499,
    n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
    n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
    n7521, n7522, n7523, n7524, n7525, n7526, n7530, n7533, n7534, n7537,
    n7540, n7541, n7544, n7547, n7550, n7553, n7554, n7555, n7556, n7557,
    n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567,
    n7568, n7569, n7570, n7571, n7572, n7574, n7575, n7576, n7577, n7578,
    n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
    n7589, n7590, n7591, n7592, n7593, n7594, n7596, n7597, n7598, n7599,
    n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
    n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7618, n7619, n7620,
    n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
    n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7639, n7640, n7641,
    n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
    n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7660, n7661, n7662,
    n7663, n7664, n7667, n7670, n7671, n7672, n7673, n7674, n7675, n7676,
    n7677, n7678, n7679, n7680, n7681, n7682, n7684, n7685, n7686, n7687,
    n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697,
    n7698, n7699, n7700, n7701, n7702, n7704, n7705, n7706, n7707, n7708,
    n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
    n7719, n7720, n7721, n7723, n7724, n7725, n7726, n7728, n7729, n7730,
    n7731, n7732, n7733, n7735, n7736, n7737, n7739, n7740, n7741, n7743,
    n7744, n7745, n7746, n7747, n7749, n7750, n7751, n7753, n7754, n7755,
    n7756, n7757, n7759, n7760, n7761, n7763, n7764, n7765, n7766, n7767,
    n7768, n7770, n7771, n7772, n7774, n7775, n7776, n7778, n7779, n7780,
    n7781, n7782, n7784, n7785, n7786, n7787, n7788, n7790, n7791, n7792,
    n7793, n7794, n7796, n7797, n7798, n7799, n7800, n7802, n7803, n7804,
    n7805, n7806, n7808, n7809, n7810, n7811, n7813, n7814, n7815, n7816,
    n7817, n7819, n7820, n7821, n7822, n7823, n7825, n7826, n7827, n7828,
    n7829, n7830, n7832, n7833, n7834, n7835, n7836, n7838, n7839, n7840,
    n7841, n7842, n7844, n7845, n7846, n7847, n7849, n7850, n7851, n7852,
    n7853, n7855, n7856, n7857, n7858, n7859, n7861, n7862, n7863, n7864,
    n7865, n7867, n7868, n7869, n7870, n7872, n7873, n7874, n7875, n7876,
    n7878, n7879, n7880, n7881, n7882, n7884, n7885, n7886, n7887, n7888,
    n7890, n7891, n7892, n7893, n7895, n7896, n7897, n7898, n7899, n7901,
    n7902, n7903, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7913,
    n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
    n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
    n7935, n7936, n7937, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
    n7946, n7947, n7948, n7949, n7950, n7952, n7953, n7954, n7955, n7956,
    n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7967,
    n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977,
    n7978, n7979, n7980, n7981, n7982, n7983, n7985, n7986, n7987, n7988,
    n7989, n7990, n7991, n7993, n7994, n7995, n7996, n7997, n7999, n8000,
    n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8009, n8010, n8011,
    n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021,
    n8022, n8023, n8024, n8025, n8027, n8028, n8029, n8030, n8031, n8032,
    n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
    n8043, n8044, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
    n8054, n8055, n8056, n8057, n8058, n8060, n8061, n8062, n8063, n8064,
    n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
    n8075, n8076, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
    n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8094, n8095, n8096,
    n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106,
    n8107, n8108, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117,
    n8118, n8119, n8120, n8121, n8122, n8123, n8125, n8126, n8127, n8128,
    n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
    n8139, n8140, n8141, n8142, n8144, n8145, n8146, n8147, n8148, n8149,
    n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8158, n8159, n8160,
    n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170,
    n8171, n8172, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181,
    n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8190, n8191, n8192,
    n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
    n8203, n8204, n8205, n8206, n8208, n8209, n8210, n8211, n8212, n8213,
    n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8223, n8224,
    n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
    n8235, n8236, n8237, n8238, n8239, n8240, n8242, n8243, n8244, n8245,
    n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
    n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266,
    n8267, n8268, n8269, n8270, n8271, n8273, n8274, n8275, n8276, n8277,
    n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
    n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
    n8299, n8300, n8301, n8302, n8303, n8304, n8306, n8307, n8308, n8309,
    n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
    n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330,
    n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8339, n8340, n8341,
    n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8351, n8352,
    n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
    n8363, n8364, n8365, n8366, n8368, n8369, n8370, n8371, n8372, n8373,
    n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8383, n8384,
    n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
    n8395, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
    n8406, n8407, n8408, n8409, n8411, n8412, n8413, n8414, n8415, n8416,
    n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8426, n8427,
    n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437,
    n8438, n8439, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
    n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8459,
    n8460, n8461, n8462, n8464, n8465, n8467, n8469, n8471, n8472, n8474,
    n8475, n8477, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486,
    n8487, n8489, n8490, n8491, n8493, n8497, n8499, n8500, n8501, n8503,
    n8504, n8506, n8507, n8508, n8509, n8511, n8512, n8513, n8514, n8516,
    n8517, n8519, n8520, n8522, n8523, n8524, n8525, n8527, n8528, n8530,
    n8531, n8533, n8534, n8536, n8537, n8539, n8540, n8542, n8543, n8545,
    n8546, n8548, n8549, n8551, n8552, n8554, n8555, n8557, n8558, n8560,
    n8561, n8563, n8564, n8566, n8567, n8569, n8570, n8572, n8573, n8575,
    n8576, n8578, n8579, n8581, n8582, n8584, n8585, n8587, n8588, n8590,
    n8591, n8593, n8594, n8596, n8597, n8599, n8600, n8602, n8603, n8605,
    n8606, n8608, n8609, n8611, n8612, n8614, n8615, n8616, n8617, n8618,
    n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
    n8629, n8630, n8631, n8632, n8633, n8635, n8636, n8637, n8638, n8639,
    n8640, n8641, n8642, n8644, n8645, n8646, n8647, n8648, n8650, n8651,
    n8652, n8653, n8655, n8656, n8657, n8659, n8661, n8663, n8665, n8667,
    n8669, n8671, n8673, n8675, n8677, n8679, n8681, n8683, n8685, n8687,
    n8689, n8691, n8693, n8695, n8697, n8699, n8701, n8703, n8705, n8707,
    n8709, n8711, n8713, n8715, n8717, n8719, n8720, n8721, n8722, n8723,
    n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
    n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743,
    n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753,
    n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763,
    n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773,
    n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783,
    n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793,
    n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
    n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
    n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
    n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
    n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843,
    n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853,
    n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863,
    n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873,
    n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883,
    n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893,
    n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903,
    n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913,
    n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923,
    n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933,
    n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943,
    n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
    n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963,
    n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973,
    n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
    n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
    n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
    n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
    n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9024,
    n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
    n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
    n9045, n9046, n9047, n9048, n9049, n9051, n9052, n9053, n9054, n9055,
    n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
    n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
    n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
    n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
    n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
    n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
    n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
    n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9137,
    n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
    n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
    n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
    n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
    n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
    n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
    n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
    n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
    n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
    n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
    n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
    n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
    n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
    n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
    n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
    n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
    n9298, n9299, n9300, n9301, n9303, n9304, n9305, n9307, n9308, n9309,
    n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
    n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
    n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
    n9340, n9341, n9342, n9343, n9347, n9348, n9349, n9350, n9354, n9355,
    n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
    n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
    n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
    n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
    n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
    n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
    n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
    n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
    n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
    n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
    n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
    n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
    n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
    n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
    n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
    n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
    n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
    n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
    n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
    n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
    n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
    n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
    n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
    n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
    n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
    n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
    n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
    n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
    n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
    n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
    n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
    n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
    n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9687,
    n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
    n9703, n9704, n9705, n9706, n9707, n9708, n9710, n9711, n9712, n9713,
    n9714, n9715, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
    n9725, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
    n9736, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
    n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
    n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
    n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
    n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787,
    n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797,
    n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
    n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
    n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
    n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
    n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
    n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9858,
    n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
    n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9877, n9878, n9879,
    n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
    n9890, n9891, n9892, n9893, n9894, n9896, n9897, n9898, n9899, n9900,
    n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
    n9911, n9912, n9913, n9915, n9916, n9917, n9918, n9919, n9920, n9921,
    n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931,
    n9932, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
    n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9953,
    n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
    n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9972, n9973, n9974,
    n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
    n9985, n9986, n9987, n9988, n9989, n9991, n9992, n9993, n9994, n9995,
    n9996, n9997, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
    n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
    n10016, n10017, n10018, n10019, n10021, n10022, n10023, n10024, n10026,
    n10027, n10028, n10029, n10031, n10032, n10033, n10034, n10036, n10037,
    n10038, n10039, n10041, n10042, n10043, n10044, n10046, n10047, n10048,
    n10049, n10051, n10052, n10053, n10054, n10055, n10056, n10058, n10059,
    n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
    n10069, n10070, n10071, n10073, n10074, n10075, n10076, n10078, n10079,
    n10080, n10081, n10083, n10084, n10085, n10086, n10088, n10089, n10090,
    n10091, n10093, n10094, n10095, n10096, n10098, n10099, n10100, n10101,
    n10103, n10104, n10105, n10106, n10108, n10109, n10110, n10111, n10112,
    n10113, n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
    n10123, n10124, n10125, n10126, n10127, n10128, n10130, n10131, n10132,
    n10133, n10135, n10136, n10137, n10138, n10140, n10141, n10142, n10143,
    n10145, n10146, n10147, n10148, n10150, n10151, n10152, n10153, n10155,
    n10156, n10157, n10158, n10160, n10161, n10162, n10163, n10165, n10166,
    n10167, n10168, n10169, n10170, n10171, n10173, n10174, n10175, n10176,
    n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
    n10186, n10188, n10189, n10190, n10191, n10193, n10194, n10195, n10196,
    n10198, n10199, n10200, n10201, n10203, n10204, n10205, n10206, n10208,
    n10209, n10210, n10211, n10213, n10214, n10215, n10216, n10218, n10219,
    n10220, n10221, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
    n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
    n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10248, n10249,
    n10250, n10251, n10253, n10254, n10255, n10256, n10258, n10259, n10260,
    n10261, n10263, n10264, n10265, n10266, n10268, n10269, n10270, n10271,
    n10273, n10274, n10275, n10276, n10278, n10279, n10280, n10281, n10283,
    n10284, n10285, n10286, n10287, n10288, n10289, n10291, n10292, n10293,
    n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302,
    n10303, n10304, n10306, n10307, n10308, n10309, n10311, n10312, n10313,
    n10314, n10316, n10317, n10318, n10319, n10321, n10322, n10323, n10324,
    n10326, n10327, n10328, n10329, n10331, n10332, n10333, n10334, n10336,
    n10337, n10338, n10339, n10341, n10342, n10343, n10344, n10345, n10346,
    n10347, n10349, n10350, n10353, n10354, n10355, n10356, n10357, n10358,
    n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10368,
    n10369, n10370, n10371, n10373, n10374, n10375, n10376, n10378, n10379,
    n10380, n10381, n10383, n10384, n10385, n10386, n10388, n10389, n10390,
    n10391, n10393, n10394, n10395, n10396, n10398, n10399, n10400, n10401,
    n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
    n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420,
    n10421, n10423, n10424, n10425, n10426, n10428, n10429, n10430, n10431,
    n10433, n10434, n10435, n10436, n10438, n10439, n10440, n10441, n10443,
    n10444, n10445, n10446, n10448, n10449, n10450, n10451, n10453, n10454,
    n10455, n10456, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
    n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
    n10475, n10476, n10477, n10478, n10479, n10481, n10482, n10483, n10484,
    n10486, n10487, n10488, n10489, n10491, n10492, n10493, n10494, n10496,
    n10497, n10498, n10499, n10501, n10502, n10503, n10504, n10506, n10507,
    n10508, n10509, n10511, n10512, n10513, n10514, n10516, n10517, n10518,
    n10519, n10520, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
    n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10537, n10538,
    n10539, n10540, n10542, n10543, n10544, n10545, n10547, n10548, n10549,
    n10550, n10552, n10553, n10554, n10555, n10557, n10558, n10559, n10560,
    n10562, n10563, n10564, n10565, n10567, n10568, n10569, n10570, n10572,
    n10573, n10574, n10575, n10576, n10578, n10579, n10580, n10581, n10582,
    n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
    n10593, n10594, n10595, n10596, n10598, n10599, n10600, n10601, n10603,
    n10604, n10605, n10606, n10608, n10609, n10610, n10611, n10613, n10614,
    n10615, n10616, n10618, n10619, n10620, n10621, n10623, n10624, n10625,
    n10626, n10628, n10629, n10630, n10631, n10632, n10634, n10635, n10636,
    n10637, n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645,
    n10646, n10647, n10649, n10650, n10651, n10652, n10654, n10655, n10656,
    n10657, n10659, n10660, n10661, n10662, n10664, n10665, n10666, n10667,
    n10669, n10670, n10671, n10672, n10674, n10675, n10676, n10677, n10679,
    n10680, n10681, n10682, n10684, n10685, n10686, n10687, n10688, n10690,
    n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699,
    n10700, n10701, n10702, n10703, n10704, n10705, n10707, n10708, n10709,
    n10710, n10712, n10713, n10714, n10715, n10717, n10718, n10719, n10720,
    n10722, n10723, n10724, n10725, n10727, n10728, n10729, n10730, n10732,
    n10733, n10734, n10735, n10737, n10738, n10739, n10740, n10742, n10743,
    n10744, n10745, n10746, n10748, n10749, n10750, n10751, n10752, n10753,
    n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10763,
    n10764, n10765, n10766, n10768, n10769, n10770, n10771, n10773, n10774,
    n10775, n10776, n10778, n10779, n10780, n10781, n10783, n10784, n10785,
    n10786, n10788, n10789, n10790, n10791, n10793, n10794, n10795, n10796,
    n10798, n10799, n10800, n10801, n10804, n10805, n10806, n10807, n10808,
    n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
    n10819, n10820, n10821, n10822, n10824, n10825, n10826, n10827, n10829,
    n10830, n10831, n10832, n10834, n10835, n10836, n10837, n10839, n10840,
    n10841, n10842, n10844, n10845, n10846, n10847, n10849, n10850, n10851,
    n10852, n10854, n10855, n10856, n10857, n10858, n10859, n10861, n10862,
    n10863, n10865, n10866, n10867, n10869, n10870, n10871, n10873, n10874,
    n10875, n10877, n10879, n10880, n10882, n10883, n10884, n10885, n10886,
    n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
    n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
    n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
    n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922,
    n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931,
    n10932, n10933, n10934, n10935, n10937, n10938, n10939, n10940, n10941,
    n10942, n10943, n10944, n10946, n10947, n10948, n10949, n10950, n10951,
    n10952, n10953, n10954, n10955, n10956, n10958, n10959, n10960, n10961,
    n10962, n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971,
    n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980,
    n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989,
    n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998,
    n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
    n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
    n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
    n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034,
    n11035, n11036, n11037, n11039, n11040, n11041, n11042, n11044, n11045,
    n11046, n11048, n11049, n11050, n11051, n11052, n11054, n11055, n11056,
    n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
    n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
    n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
    n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11093,
    n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102,
    n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
    n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
    n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
    n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11138, n11139,
    n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148,
    n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157,
    n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
    n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
    n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
    n11185, n11186, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
    n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
    n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212,
    n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221,
    n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230,
    n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
    n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
    n11249, n11250, n11251, n11252, n11253, n11254, n11256, n11257, n11258,
    n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
    n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276,
    n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285,
    n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294,
    n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
    n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
    n11313, n11314, n11315, n11316, n11317, n11318, n11320, n11321, n11322,
    n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
    n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340,
    n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349,
    n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
    n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
    n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
    n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11386,
    n11387, n11388, n11389, n11390, n11391, n11392, n11395, n11396, n11397,
    n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406,
    n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
    n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
    n11425, n11426, n11427, n11428, n11429, n11430, n11432, n11433, n11434,
    n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
    n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452,
    n11453, n11454, n11456, n11457, n11458, n11459, n11460, n11461, n11462,
    n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
    n11472, n11473, n11474, n11477, n11478, n11479, n11480, n11481, n11482,
    n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
    n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500,
    n11501, n11504, n11507, n11510, n11513, n11514, n11517, n11520, n11523,
    n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534,
    n11535, n11536, n11537, n11539, n11540, n11541, n11542, n11543, n11544,
    n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
    n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
    n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
    n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580,
    n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589,
    n11590, n11591, n11592, n11594, n11595, n11596, n11597, n11598, n11599,
    n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
    n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
    n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
    n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
    n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11645,
    n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654,
    n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
    n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
    n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
    n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
    n11691, n11692, n11693, n11695, n11696, n11697, n11698, n11699, n11700,
    n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709,
    n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718,
    n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
    n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
    n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
    n11746, n11747, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
    n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764,
    n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773,
    n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782,
    n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
    n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
    n11801, n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
    n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819,
    n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828,
    n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837,
    n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846,
    n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11855, n11856,
    n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
    n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
    n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883,
    n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892,
    n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901,
    n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
    n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
    n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
    n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
    n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
    n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957,
    n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966,
    n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
    n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
    n11985, n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
    n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
    n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012,
    n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021,
    n12022, n12023, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
    n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
    n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
    n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
    n12059, n12060, n12061, n12062, n12063, n12065, n12066, n12067, n12068,
    n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077,
    n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086,
    n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
    n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12105,
    n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
    n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123,
    n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132,
    n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141,
    n12142, n12143, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
    n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
    n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
    n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
    n12179, n12180, n12181, n12183, n12184, n12185, n12186, n12187, n12188,
    n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197,
    n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206,
    n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
    n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
    n12225, n12226, n12227, n12229, n12230, n12231, n12232, n12233, n12234,
    n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243,
    n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252,
    n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261,
    n12262, n12263, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
    n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
    n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
    n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
    n12299, n12300, n12301, n12302, n12304, n12305, n12306, n12307, n12308,
    n12309, n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317,
    n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326,
    n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
    n12336, n12337, n12338, n12339, n12341, n12342, n12343, n12344, n12345,
    n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
    n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
    n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372,
    n12373, n12374, n12375, n12377, n12378, n12379, n12380, n12381, n12382,
    n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
    n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
    n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
    n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12418, n12419,
    n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427, n12428,
    n12429, n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437,
    n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446,
    n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
    n12456, n12457, n12458, n12459, n12461, n12462, n12463, n12464, n12465,
    n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
    n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
    n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492,
    n12493, n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502,
    n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
    n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
    n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
    n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12539,
    n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548,
    n12549, n12551, n12553, n12554, n12555, n12556, n12557, n12559, n12560,
    n12561, n12562, n12564, n12565, n12566, n12567, n12568, n12569, n12571,
    n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580,
    n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12590, n12591,
    n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12600, n12601,
    n12602, n12603, n12604, n12605, n12606, n12609, n12610, n12611, n12612,
    n12613, n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12624,
    n12625, n12626, n12627, n12628, n12629, n12630, n12632, n12633, n12634,
    n12635, n12636, n12637, n12639, n12640, n12641, n12642, n12643, n12644,
    n12645, n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12655,
    n12656, n12657, n12658, n12659, n12661, n12662, n12663, n12664, n12665,
    n12666, n12667, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
    n12677, n12678, n12679, n12680, n12681, n12682, n12684, n12685, n12686,
    n12687, n12688, n12689, n12690, n12692, n12693, n12694, n12695, n12696,
    n12697, n12698, n12700, n12701, n12702, n12703, n12704, n12706, n12707,
    n12708, n12709, n12710, n12711, n12712, n12714, n12715, n12716, n12717,
    n12718, n12719, n12720, n12722, n12723, n12724, n12725, n12726, n12727,
    n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12737, n12738,
    n12739, n12740, n12741, n12742, n12743, n12745, n12746, n12747, n12748,
    n12749, n12750, n12751, n12753, n12755, n12756, n12757, n12758, n12759,
    n12760, n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12770,
    n12771, n12772, n12773, n12774, n12776, n12777, n12778, n12779, n12780,
    n12781, n12783, n12784, n12785, n12786, n12788, n12789, n12790, n12791,
    n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
    n12802, n12803, n12804, n12805, n12806, n12807, n12809, n12810, n12811,
    n12812, n12813, n12814, n12816, n12817, n12818, n12819, n12820, n12822,
    n12823, n12824, n12825, n12826, n12828, n12829, n12830, n12831, n12832,
    n12834, n12835, n12836, n12837, n12838, n12840, n12841, n12842, n12843,
    n12844, n12846, n12848, n12850, n12852, n12854, n12856, n12858, n12860,
    n12862, n12864, n12866, n12868, n12870, n12872, n12874, n12876, n12878,
    n12880, n12882, n12884, n12886, n12888, n12890, n12892, n12893, n12894,
    n12895, n12896, n12897, n12898, n12899, n12900, n12902, n12903, n12905,
    n12906, n12908, n12909, n12911, n12912, n12914, n12915, n12917, n12918,
    n12920, n12921, n12923, n12924, n12926, n12927, n12929, n12930, n12932,
    n12933, n12935, n12936, n12938, n12939, n12941, n12942, n12944, n12945,
    n12947, n12948, n12949, n12951, n12952, n12954, n12955, n12957, n12958,
    n12960, n12961, n12963, n12964, n12966, n12967, n12969, n12970, n12972,
    n12973, n12975, n12976, n12978, n12979, n12981, n12982, n12984, n12985,
    n12987, n12988, n12990, n12991, n12994, n12995, n12996, n12997, n12998,
    n12999, n13000, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
    n13009, n13010, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
    n13019, n13021, n13022, n13023, n13024, n13025, n13026, n13027, n13028,
    n13030, n13031, n13032, n13033, n13034, n13036, n13037, n13038, n13039,
    n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
    n13049, n13050, n13052, n13053, n13054, n13055, n13056, n13057, n13059,
    n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067, n13068,
    n13069, n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077,
    n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086,
    n13087, n13088, n13089, n13090, n13092, n13093, n13094, n13095, n13096,
    n13097, n13098, n13100, n13101, n13102, n13103, n13104, n13106, n13107,
    n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116,
    n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125,
    n13126, n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
    n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
    n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
    n13155, n13156, n13157, n13158, n13159, n13161, n13162, n13163, n13164,
    n13165, n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173,
    n13174, n13175, n13176, n13177, n13178, n13179, n13181, n13182, n13183,
    n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
    n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13202,
    n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211,
    n13213, n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221,
    n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230,
    n13231, n13232, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
    n13242, n13243, n13244, n13245, n13246, n13248, n13249, n13250, n13251,
    n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260,
    n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13269, n13270,
    n13271, n13274, n13277, n13280, n13283, n13284, n13287, n13290, n13293,
    n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
    n13305, n13306, n13307, n13309, n13310, n13311, n13312, n13313, n13314,
    n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323,
    n13324, n13325, n13326, n13327, n13328, n13329, n13331, n13332, n13333,
    n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342,
    n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
    n13352, n13353, n13354, n13356, n13357, n13358, n13359, n13360, n13361,
    n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
    n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13380,
    n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389,
    n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398,
    n13399, n13400, n13401, n13402, n13404, n13405, n13406, n13407, n13408,
    n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
    n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
    n13427, n13429, n13430, n13431, n13432, n13433, n13434, n13435, n13436,
    n13437, n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445,
    n13446, n13447, n13448, n13449, n13450, n13451, n13453, n13454, n13455,
    n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
    n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
    n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
    n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491,
    n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499, n13500,
    n13501, n13502, n13503, n13504, n13506, n13507, n13508, n13509, n13510,
    n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
    n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
    n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
    n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
    n13547, n13548, n13550, n13551, n13552, n13553, n13554, n13555, n13557,
    n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566,
    n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
    n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
    n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13594,
    n13595, n13596, n13597, n13598, n13599, n13600, n13602, n13603, n13604,
    n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613,
    n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622,
    n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
    n13632, n13633, n13634, n13635, n13636, n13638, n13639, n13640, n13641,
    n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
    n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659,
    n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667, n13668,
    n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677,
    n13678, n13680, n13681, n13682, n13683, n13684, n13685, n13687, n13688,
    n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
    n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
    n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715,
    n13716, n13717, n13718, n13719, n13720, n13722, n13723, n13724, n13725,
    n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734,
    n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
    n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
    n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
    n13762, n13763, n13764, n13766, n13767, n13768, n13769, n13771, n13772,
    n13773, n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781,
    n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790,
    n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
    n13800, n13801, n13802, n13803, n13806, n13807, n13808, n13809, n13810,
    n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819,
    n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828,
    n13829, n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837,
    n13838, n13839, n13840, n13841, n13843, n13844, n13846, n13847, n13848,
    n13849, n13850, n13852, n13854, n13856, n13858, n13860, n13862, n13863,
    n13865, n13867, n13869, n13871, n13873, n13875, n13877, n13879, n13881,
    n13883, n13885, n13887, n13889, n13891, n13893, n13895, n13897, n13899,
    n13901, n13903, n13905, n13907, n13909, n13910, n13912, n13913, n13914,
    n13916, n13918, n13919, n13920, n13921, n13922, n13924, n13925, n13926,
    n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
    n13936, n13937, n13938, n13940, n13941, n13942, n13943, n13944, n13945,
    n13946, n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955,
    n13956, n13957, n13959, n13960, n13961, n13962, n13963, n13964, n13965,
    n13966, n13967, n13968, n13969, n13970, n13972, n13973, n13974, n13975,
    n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13985,
    n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
    n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14004, n14005,
    n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014,
    n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
    n14025, n14026, n14027, n14028, n14029, n14031, n14032, n14033, n14034,
    n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14043, n14044,
    n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053,
    n14054, n14055, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
    n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14072, n14073,
    n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
    n14083, n14084, n14085, n14087, n14088, n14089, n14090, n14091, n14092,
    n14093, n14094, n14095, n14096, n14097, n14098, n14100, n14101, n14102,
    n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
    n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
    n14122, n14123, n14124, n14125, n14126, n14127, n14129, n14130, n14131,
    n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140,
    n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150,
    n14151, n14152, n14153, n14154, n14155, n14156, n14158, n14159, n14160,
    n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
    n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179,
    n14180, n14181, n14182, n14184, n14185, n14186, n14187, n14188, n14189,
    n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14198, n14199,
    n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
    n14209, n14210, n14211, n14212, n14214, n14215, n14216, n14217, n14218,
    n14219, n14220, n14221, n14222, n14223, n14224, n14226, n14227, n14228,
    n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237,
    n14238, n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
    n14248, n14249, n14250, n14252, n14253, n14254, n14255, n14256, n14257,
    n14258, n14259, n14260, n14261, n14262, n14263, n14265, n14266, n14267,
    n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14277,
    n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286,
    n14287, n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
    n14297, n14298, n14299, n14300, n14302, n14303, n14304, n14305, n14306,
    n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14315, n14316,
    n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325,
    n14326, n14327, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
    n14336, n14337, n14338, n14339, n14340, n14342, n14343, n14344, n14345,
    n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14355,
    n14356, n14358, n14359, n14360, n14361, n14362, n14363, n14365, n14366,
    n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
    n14376, n14377, n14378, n14379, n14380, n14382, n14383, n14384, n14385,
    n14386, n14388, n14390, n14391, n14393, n14394, n14396, n14397, n14398,
    n14399, n14401, n14402, n14404, n14406, n14407, n14408, n14409, n14410,
    n14411, n14412, n14413, n14414, n14415, n14417, n14418, n14419, n14421,
    n14423, n14425, n14427, n14428, n14430, n14431, n14432, n14433, n14434,
    n14436, n14437, n14438, n14439, n14441, n14442, n14443, n14444, n14446,
    n14447, n14449, n14450, n14452, n14453, n14454, n14455, n14457, n14458,
    n14460, n14461, n14463, n14464, n14466, n14467, n14469, n14470, n14472,
    n14473, n14475, n14476, n14478, n14479, n14481, n14482, n14484, n14485,
    n14487, n14488, n14490, n14491, n14493, n14494, n14496, n14497, n14499,
    n14500, n14502, n14503, n14505, n14506, n14508, n14509, n14511, n14512,
    n14514, n14515, n14517, n14518, n14520, n14521, n14523, n14524, n14526,
    n14527, n14529, n14530, n14532, n14533, n14535, n14536, n14538, n14539,
    n14541, n14542, n14544, n14545, n14546, n14547, n14548, n14549, n14550,
    n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559,
    n14560, n14561, n14562, n14563, n14564, n14566, n14567, n14568, n14569,
    n14570, n14571, n14572, n14574, n14575, n14576, n14577, n14578, n14580,
    n14581, n14582, n14583, n14585, n14586, n14587, n14589, n14591, n14593,
    n14595, n14597, n14599, n14601, n14603, n14605, n14607, n14609, n14611,
    n14613, n14615, n14617, n14619, n14621, n14623, n14625, n14627, n14629,
    n14631, n14633, n14635, n14637, n14639, n14641, n14643, n14645, n14647,
    n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
    n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
    n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675,
    n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684,
    n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693,
    n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702,
    n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711,
    n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
    n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
    n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
    n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
    n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756,
    n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765,
    n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774,
    n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783,
    n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
    n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
    n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
    n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
    n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828,
    n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837,
    n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846,
    n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855,
    n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
    n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
    n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
    n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
    n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900,
    n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909,
    n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918,
    n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927,
    n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
    n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
    n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
    n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
    n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972,
    n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981,
    n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990,
    n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999,
    n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
    n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
    n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
    n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
    n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044,
    n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053,
    n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062,
    n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071,
    n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
    n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
    n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
    n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107,
    n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116,
    n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125,
    n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134,
    n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143,
    n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
    n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
    n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,
    n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179,
    n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188,
    n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197,
    n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206,
    n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215,
    n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
    n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
    n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242,
    n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251,
    n15252, n15253, n15255, n15256, n15257, n15258, n15259, n15260, n15261,
    n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270,
    n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279,
    n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
    n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
    n15298, n15299, n15300, n15301, n15302, n15304, n15305, n15306, n15307,
    n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317,
    n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327,
    n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
    n15337, n15338, n15339, n15340, n15341, n15342, n15344, n15345, n15346,
    n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
    n15357, n15359, n15360, n15361, n15362, n15363, n15365, n15366, n15367,
    n15370, n15372, n15373, n15375, n15376, n15378, n15379, n15380, n15381,
    n15382, n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391,
    n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
    n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15411,
    n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420,
    n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429,
    n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438,
    n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447,
    n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
    n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
    n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474,
    n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483,
    n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492,
    n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501,
    n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509, n15510,
    n15511, n15512, n15513, n15514, n15515, n15517, n15518, n15519, n15520,
    n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
    n15530, n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539,
    n15540, n15541, n15542, n15543, n15544, n15545, n15547, n15548, n15549,
    n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558,
    n15559, n15560, n15562, n15563, n15564, n15565, n15566, n15567, n15568,
    n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15578,
    n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587,
    n15588, n15589, n15590, n15591, n15592, n15594, n15595, n15596, n15597,
    n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606,
    n15607, n15608, n15610, n15611, n15612, n15613, n15614, n15615, n15616,
    n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15626,
    n15627, n15628, n15629, n15630, n15631, n15634, n15635, n15636, n15637,
    n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645, n15646,
    n15647, n15648, n15650, n15651, n15652, n15653, n15655, n15656, n15657,
    n15658, n15660, n15661, n15662, n15663, n15665, n15666, n15667, n15668,
    n15670, n15671, n15672, n15673, n15675, n15676, n15677, n15678, n15680,
    n15681, n15682, n15683, n15685, n15686, n15687, n15688, n15692, n15693,
    n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701, n15702,
    n15703, n15704, n15705, n15706, n15708, n15709, n15710, n15711, n15713,
    n15714, n15715, n15716, n15718, n15719, n15720, n15721, n15723, n15724,
    n15725, n15726, n15728, n15729, n15730, n15731, n15733, n15734, n15735,
    n15736, n15738, n15739, n15740, n15741, n15743, n15744, n15745, n15746,
    n15747, n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15758,
    n15759, n15760, n15761, n15762, n15763, n15764, n15766, n15767, n15768,
    n15769, n15771, n15772, n15773, n15774, n15776, n15777, n15778, n15779,
    n15781, n15782, n15783, n15784, n15786, n15787, n15788, n15789, n15791,
    n15792, n15793, n15794, n15796, n15797, n15798, n15799, n15801, n15802,
    n15803, n15804, n15805, n15807, n15808, n15809, n15810, n15811, n15812,
    n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821,
    n15822, n15824, n15825, n15826, n15827, n15829, n15830, n15831, n15832,
    n15834, n15835, n15836, n15837, n15839, n15840, n15841, n15842, n15844,
    n15845, n15846, n15847, n15849, n15850, n15851, n15852, n15854, n15855,
    n15856, n15857, n15859, n15860, n15861, n15863, n15864, n15865, n15866,
    n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875,
    n15876, n15877, n15879, n15880, n15881, n15882, n15884, n15885, n15886,
    n15887, n15889, n15890, n15891, n15892, n15894, n15895, n15896, n15897,
    n15899, n15900, n15901, n15902, n15904, n15905, n15906, n15907, n15909,
    n15910, n15911, n15912, n15914, n15915, n15916, n15918, n15919, n15920,
    n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
    n15930, n15931, n15933, n15934, n15935, n15936, n15938, n15939, n15940,
    n15941, n15943, n15944, n15945, n15946, n15948, n15949, n15950, n15951,
    n15953, n15954, n15955, n15956, n15958, n15959, n15960, n15961, n15963,
    n15964, n15965, n15966, n15968, n15969, n15970, n15972, n15973, n15974,
    n15975, n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983,
    n15984, n15985, n15987, n15988, n15989, n15990, n15992, n15993, n15994,
    n15995, n15997, n15998, n15999, n16000, n16002, n16003, n16004, n16005,
    n16007, n16008, n16009, n16010, n16012, n16013, n16014, n16015, n16017,
    n16018, n16019, n16020, n16022, n16023, n16025, n16026, n16027, n16028,
    n16029, n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037,
    n16038, n16039, n16040, n16042, n16043, n16044, n16045, n16047, n16048,
    n16049, n16050, n16052, n16053, n16054, n16055, n16057, n16058, n16059,
    n16060, n16062, n16063, n16064, n16065, n16067, n16068, n16069, n16070,
    n16072, n16073, n16074, n16075, n16077, n16078, n16079, n16081, n16082,
    n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091,
    n16092, n16093, n16094, n16096, n16097, n16098, n16099, n16101, n16102,
    n16103, n16104, n16106, n16107, n16108, n16109, n16111, n16112, n16113,
    n16114, n16116, n16117, n16118, n16119, n16121, n16122, n16123, n16124,
    n16126, n16127, n16128, n16129, n16131, n16132, n16133, n16135, n16136,
    n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
    n16146, n16147, n16148, n16150, n16151, n16152, n16153, n16155, n16156,
    n16157, n16158, n16160, n16161, n16162, n16163, n16165, n16166, n16167,
    n16168, n16170, n16171, n16172, n16173, n16175, n16176, n16177, n16178,
    n16180, n16181, n16182, n16183, n16185, n16186, n16187, n16189, n16190,
    n16191, n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199,
    n16200, n16201, n16202, n16204, n16205, n16206, n16207, n16209, n16210,
    n16211, n16212, n16214, n16215, n16216, n16217, n16219, n16220, n16221,
    n16222, n16224, n16225, n16226, n16227, n16229, n16230, n16231, n16232,
    n16234, n16235, n16236, n16237, n16239, n16240, n16241, n16242, n16244,
    n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253,
    n16254, n16255, n16256, n16257, n16258, n16260, n16261, n16262, n16263,
    n16265, n16266, n16267, n16268, n16270, n16271, n16272, n16273, n16275,
    n16276, n16277, n16278, n16280, n16281, n16282, n16283, n16285, n16286,
    n16287, n16288, n16290, n16291, n16292, n16293, n16295, n16296, n16297,
    n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307,
    n16308, n16309, n16310, n16311, n16312, n16314, n16315, n16316, n16317,
    n16319, n16320, n16321, n16322, n16324, n16325, n16326, n16327, n16329,
    n16330, n16331, n16332, n16334, n16335, n16336, n16337, n16339, n16340,
    n16341, n16342, n16344, n16345, n16346, n16347, n16349, n16350, n16351,
    n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
    n16362, n16363, n16364, n16365, n16366, n16368, n16369, n16370, n16371,
    n16373, n16374, n16375, n16376, n16378, n16379, n16380, n16381, n16383,
    n16384, n16385, n16386, n16388, n16389, n16390, n16391, n16393, n16394,
    n16395, n16396, n16398, n16399, n16400, n16401, n16403, n16404, n16407,
    n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416,
    n16417, n16418, n16419, n16420, n16422, n16423, n16424, n16425, n16427,
    n16428, n16429, n16430, n16432, n16433, n16434, n16435, n16437, n16438,
    n16439, n16440, n16442, n16443, n16444, n16445, n16447, n16448, n16449,
    n16450, n16452, n16453, n16454, n16455, n16457, n16458, n16459, n16460,
    n16461, n16463, n16464, n16465, n16467, n16468, n16469, n16471, n16472,
    n16473, n16474, n16476, n16477, n16478, n16480, n16481, n16483, n16484,
    n16486, n16487, n16488, n16489, n16490, n16491, n16492, n16493, n16496,
    n16497, n16498, n16499, n16500, n16502, n16503, n16504, n16505, n16506,
    n16508, n16509, n16510, n16511, n16513, n16514, n16515, n16516, n16517,
    n16518, n16519, n16520, n16521, n16522, n16523, n16524, n16525, n16526,
    n16527, n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535,
    n16536, n16537, n16538, n16540, n16541, n16542, n16543, n16544, n16545,
    n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554,
    n16555, n16556, n16557, n16558, n16559, n16560, n16562, n16563, n16564,
    n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572, n16573,
    n16574, n16575, n16576, n16577, n16578, n16579, n16580, n16581, n16582,
    n16583, n16584, n16585, n16586, n16587, n16588, n16590, n16591, n16592,
    n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
    n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610,
    n16611, n16612, n16613, n16614, n16616, n16617, n16618, n16619, n16620,
    n16621, n16622, n16623, n16624, n16625, n16627, n16628, n16629, n16630,
    n16631, n16632, n16633, n16634, n16635, n16636, n16637, n16638, n16639,
    n16640, n16641, n16642, n16643, n16645, n16646, n16647, n16648, n16649,
    n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658,
    n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666, n16667,
    n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675, n16676,
    n16677, n16678, n16679, n16680, n16681, n16682, n16683, n16684, n16685,
    n16686, n16687, n16688, n16689, n16690, n16691, n16692, n16693, n16695,
    n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704,
    n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
    n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722,
    n16723, n16724, n16725, n16728, n16729, n16730, n16731, n16732, n16733,
    n16734, n16735, n16736, n16737, n16738, n16739, n16740, n16741, n16742,
    n16743, n16744, n16745, n16746, n16747, n16748, n16749, n16750, n16751,
    n16752, n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
    n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770,
    n16771, n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779,
    n16780, n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788,
    n16789, n16790, n16791, n16792, n16793, n16794, n16795, n16796, n16797,
    n16798, n16799, n16800, n16801, n16802, n16803, n16804, n16805, n16806,
    n16808, n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816,
    n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16827,
    n16828, n16829, n16830, n16831, n16832, n16833, n16834, n16835, n16836,
    n16837, n16838, n16839, n16840, n16841, n16842, n16843, n16844, n16845,
    n16846, n16847, n16848, n16849, n16850, n16851, n16852, n16853, n16854,
    n16856, n16857, n16858, n16859, n16862, n16865, n16868, n16871, n16872,
    n16875, n16878, n16881, n16884, n16885, n16886, n16887, n16888, n16889,
    n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897, n16898,
    n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907,
    n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915, n16916,
    n16917, n16918, n16919, n16920, n16921, n16923, n16924, n16925, n16926,
    n16927, n16928, n16929, n16930, n16931, n16932, n16933, n16934, n16935,
    n16936, n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944,
    n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
    n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16962, n16963,
    n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971, n16972,
    n16973, n16974, n16975, n16976, n16977, n16978, n16979, n16980, n16981,
    n16982, n16983, n16984, n16985, n16986, n16988, n16989, n16990, n16991,
    n16992, n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000,
    n17001, n17002, n17003, n17005, n17006, n17007, n17008, n17009, n17010,
    n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019,
    n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027, n17028,
    n17029, n17030, n17031, n17032, n17033, n17034, n17035, n17036, n17037,
    n17038, n17039, n17040, n17041, n17042, n17043, n17044, n17045, n17046,
    n17047, n17048, n17049, n17050, n17052, n17053, n17054, n17055, n17056,
    n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
    n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074,
    n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082, n17083,
    n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091, n17092,
    n17093, n17094, n17096, n17097, n17098, n17099, n17100, n17101, n17102,
    n17103, n17104, n17105, n17106, n17107, n17108, n17109, n17110, n17111,
    n17112, n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
    n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130,
    n17131, n17133, n17134, n17135, n17136, n17137, n17138, n17139, n17140,
    n17141, n17142, n17143, n17144, n17145, n17146, n17147, n17148, n17149,
    n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17158, n17159,
    n17160, n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168,
    n17169, n17170, n17171, n17172, n17173, n17175, n17176, n17177, n17178,
    n17179, n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187,
    n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195, n17196,
    n17197, n17198, n17199, n17200, n17201, n17202, n17203, n17204, n17205,
    n17206, n17207, n17208, n17209, n17210, n17211, n17212, n17213, n17214,
    n17215, n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224,
    n17225, n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
    n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242,
    n17243, n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251,
    n17253, n17254, n17255, n17256, n17257, n17259, n17260, n17261, n17262,
    n17263, n17264, n17265, n17266, n17267, n17268, n17269, n17270, n17271,
    n17272, n17273, n17274, n17275, n17276, n17278, n17279, n17280, n17281,
    n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17290,
    n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299,
    n17300, n17303, n17304, n17305, n17306, n17307, n17308, n17309, n17310,
    n17311, n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319,
    n17320, n17321, n17322, n17323, n17324, n17325, n17326, n17328, n17329,
    n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338,
    n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347,
    n17348, n17350, n17351, n17352, n17353, n17354, n17355, n17356, n17357,
    n17358, n17359, n17360, n17361, n17362, n17363, n17364, n17365, n17366,
    n17367, n17368, n17369, n17370, n17371, n17374, n17375, n17376, n17377,
    n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386,
    n17387, n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395,
    n17396, n17397, n17399, n17400, n17401, n17405, n17406, n17407, n17408,
    n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
    n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425, n17426,
    n17427, n17429, n17430, n17431, n17432, n17433, n17434, n17435, n17436,
    n17437, n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445,
    n17446, n17447, n17448, n17450, n17451, n17452, n17453, n17454, n17455,
    n17456, n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464,
    n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17473, n17474,
    n17477, n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485,
    n17486, n17487, n17488, n17489, n17490, n17491, n17492, n17493, n17494,
    n17495, n17496, n17497, n17498, n17500, n17501, n17502, n17503, n17504,
    n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
    n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522,
    n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531, n17532,
    n17533, n17534, n17535, n17536, n17537, n17538, n17539, n17540, n17541,
    n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17550, n17551,
    n17552, n17553, n17554, n17555, n17556, n17558, n17559, n17561, n17563,
    n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578,
    n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587,
    n17588, n17589, n17590, n17591, n17593, n17594, n17595, n17596, n17597,
    n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605, n17606,
    n17607, n17608, n17609, n17610, n17611, n17612, n17613, n17614, n17615,
    n17616, n17617, n17618, n17619, n17621, n17622, n17623, n17628, n17633,
    n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17642,
    n17643, n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651,
    n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659, n17660,
    n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669, n17670,
    n17671, n17672, n17673, n17674, n17675, n17676, n17677, n17678, n17679,
    n17680, n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688,
    n17690, n17693, n17694, n17695, n17696, n17697, n17699, n17700, n17701,
    n17702, n17703, n17704, n17705, n17706, n17707, n17708, n17709, n17710,
    n17711, n17712, n17713, n17714, n17715, n17716, n17717, n17718, n17719,
    n17720, n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
    n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738,
    n17739, n17740, n17741, n17742, n17743, n17744, n17747, n17748, n17749,
    n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758,
    n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766, n17768,
    n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
    n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17786,
    n17787, n17788, n17789, n17790, n17792, n17793, n17794, n17795, n17796,
    n17797, n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805,
    n17806, n17807, n17808, n17809, n17810, n17811, n17812, n17813, n17814,
    n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824,
    n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
    n17834, n17835, n17836, n17838, n17839, n17840, n17841, n17842, n17843,
    n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851, n17852,
    n17853, n17854, n17856, n17857, n17858, n17859, n17860, n17861, n17862,
    n17863, n17864, n17865, n17866, n17867, n17868, n17869, n17870, n17871,
    n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879, n17880,
    n17881, n17883, n17884, n17885, n17886, n17887, n17888, n17889, n17890,
    n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899,
    n17900, n17902, n17903, n17904, n17905, n17906, n17907, n17908, n17909,
    n17910, n17911, n17912, n17913, n17914, n17915, n17916, n17917, n17918,
    n17919, n17920, n17921, n17922, n17924, n17925, n17926, n17927, n17928,
    n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
    n17938, n17939, n17940, n17942, n17943, n17944, n17945, n17946, n17947,
    n17948, n17949, n17950, n17951, n17952, n17953, n17954, n17955, n17956,
    n17957, n17958, n17959, n17960, n17961, n17962, n17963, n17964, n17965,
    n17966, n17968, n17969, n17970, n17971, n17972, n17973, n17974, n17975,
    n17976, n17977, n17978, n17979, n17980, n17981, n17982, n17983, n17984,
    n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994,
    n17995, n17996, n17997, n17998, n17999, n18000, n18001, n18002, n18003,
    n18004, n18005, n18006, n18007, n18009, n18010, n18011, n18012, n18013,
    n18014, n18015, n18016, n18017, n18018, n18019, n18020, n18021, n18022,
    n18023, n18024, n18025, n18026, n18027, n18028, n18030, n18031, n18032,
    n18033, n18034, n18037, n18040, n18043, n18046, n18047, n18050, n18053,
    n18056, n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066,
    n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074, n18075,
    n18076, n18077, n18078, n18079, n18080, n18081, n18082, n18083, n18084,
    n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093, n18094,
    n18095, n18096, n18097, n18098, n18099, n18100, n18101, n18102, n18103,
    n18104, n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112,
    n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121, n18122,
    n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130, n18131,
    n18132, n18133, n18134, n18135, n18136, n18137, n18138, n18139, n18140,
    n18141, n18142, n18143, n18144, n18146, n18147, n18148, n18149, n18150,
    n18151, n18152, n18153, n18154, n18155, n18156, n18157, n18158, n18159,
    n18160, n18161, n18162, n18163, n18164, n18165, n18166, n18167, n18168,
    n18169, n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
    n18179, n18180, n18181, n18182, n18183, n18184, n18185, n18186, n18187,
    n18188, n18189, n18190, n18191, n18192, n18193, n18194, n18195, n18196,
    n18197, n18198, n18199, n18200, n18201, n18202, n18203, n18204, n18205,
    n18206, n18208, n18209, n18210, n18211, n18212, n18213, n18215, n18216,
    n18217, n18220, n18221, n18223, n18224, n18225, n18226, n18227, n18228,
    n18229, n18230, n18231, n18232, n18233, n18234, n18235, n18236, n18237,
    n18238, n18239, n18240, n18241, n18242, n18243, n18244, n18245, n18246,
    n18247, n18248, n18249, n18250, n18252, n18253, n18254, n18255, n18256,
    n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
    n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273, n18274,
    n18275, n18276, n18277, n18278, n18279, n18280, n18281, n18282, n18283,
    n18284, n18285, n18286, n18287, n18288, n18290, n18291, n18292, n18293,
    n18296, n18299, n18300, n18303, n18306, n18307, n18310, n18313, n18316,
    n18319, n18320, n18321, n18322, n18323, n18324, n18325, n18326, n18327,
    n18328, n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336,
    n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
    n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18354, n18355,
    n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363, n18364,
    n18365, n18366, n18367, n18368, n18369, n18370, n18371, n18372, n18373,
    n18374, n18375, n18376, n18377, n18378, n18379, n18380, n18381, n18382,
    n18383, n18384, n18385, n18387, n18388, n18389, n18390, n18391, n18392,
    n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
    n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409, n18410,
    n18411, n18412, n18413, n18414, n18415, n18416, n18418, n18419, n18420,
    n18421, n18422, n18423, n18424, n18425, n18426, n18427, n18428, n18429,
    n18430, n18431, n18432, n18433, n18434, n18435, n18436, n18437, n18438,
    n18439, n18440, n18441, n18442, n18443, n18444, n18445, n18446, n18447,
    n18448, n18449, n18450, n18451, n18452, n18453, n18455, n18456, n18457,
    n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465, n18466,
    n18467, n18468, n18469, n18470, n18471, n18472, n18473, n18474, n18475,
    n18476, n18477, n18478, n18479, n18481, n18482, n18483, n18484, n18485,
    n18486, n18487, n18488, n18490, n18491, n18492, n18493, n18494, n18495,
    n18496, n18497, n18498, n18499, n18500, n18501, n18502, n18503, n18504,
    n18505, n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
    n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521, n18522,
    n18523, n18524, n18525, n18526, n18527, n18529, n18530, n18531, n18532,
    n18533, n18534, n18535, n18536, n18537, n18538, n18539, n18540, n18541,
    n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549, n18550,
    n18551, n18552, n18553, n18554, n18555, n18556, n18557, n18558, n18559,
    n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
    n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577, n18578,
    n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587,
    n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595, n18596,
    n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605, n18606,
    n18607, n18608, n18609, n18610, n18611, n18612, n18613, n18614, n18615,
    n18616, n18617, n18618, n18619, n18620, n18621, n18622, n18624, n18625,
    n18626, n18627, n18628, n18629, n18630, n18631, n18633, n18634, n18635,
    n18636, n18638, n18639, n18640, n18641, n18643, n18644, n18645, n18646,
    n18648, n18649, n18650, n18651, n18653, n18654, n18655, n18656, n18658,
    n18659, n18660, n18661, n18663, n18664, n18665, n18666, n18668, n18669,
    n18670, n18672, n18673, n18674, n18676, n18677, n18678, n18680, n18681,
    n18682, n18684, n18685, n18686, n18688, n18689, n18690, n18692, n18693,
    n18694, n18696, n18697, n18698, n18700, n18701, n18703, n18704, n18706,
    n18707, n18709, n18710, n18712, n18713, n18715, n18716, n18718, n18719,
    n18721, n18722, n18724, n18725, n18727, n18728, n18730, n18731, n18733,
    n18734, n18736, n18737, n18739, n18740, n18742, n18743, n18745, n18746,
    n18747, n18748, n18749, n18750, n18751, n18752, n18753, n18755, n18757,
    n18759, n18760, n18762, n18764, n18765, n18767, n18768, n18770, n18771,
    n18773, n18774, n18776, n18778, n18780, n18782, n18784, n18786, n18788,
    n18790, n18791, n18792, n18794, n18795, n18797, n18798, n18800, n18801,
    n18803, n18804, n18806, n18808, n18810, n18812, n18814, n18815, n18817,
    n18818, n18820, n18821, n18823, n18824, n18826, n18827, n18829, n18831,
    n18833, n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
    n18842, n18843, n18845, n18847, n18849, n18850, n18852, n18854, n18856,
    n18858, n18860, n18862, n18864, n18866, n18867, n18869, n18871, n18873,
    n18875, n18876, n18878, n18879, n18880, n18881, n18882, n18884, n18885,
    n18887, n18888, n18889, n18891, n18892, n18894, n18895, n18897, n18898,
    n18900, n18901, n18903, n18904, n18906, n18907, n18909, n18910, n18912,
    n18913, n18915, n18916, n18917, n18919, n18920, n18922, n18923, n18925,
    n18926, n18928, n18929, n18930, n18932, n18933, n18934, n18935, n18936,
    n18937, n18938, n18939, n18940, n18942, n18944, n18946, n18947, n18949,
    n18950, n18952, n18953, n18955, n18956, n18958, n18959, n18961, n18962,
    n18964, n18965, n18967, n18968, n18970, n18971, n18973, n18974, n18976,
    n18977, n18979, n18980, n18982, n18983, n18985, n18986, n18988, n18989,
    n18991, n18992, n18994, n18995, n18997, n18998, n19000, n19001, n19003,
    n19004, n19006, n19007, n19009, n19010, n19012, n19013, n19015, n19016,
    n19018, n19019, n19021, n19022, n19023, n19025, n19026, n19028, n19029,
    n19031, n19033, n19034, n19035, n19036, n19037, n19038, n19039, n19040,
    n19041, n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
    n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057, n19058,
    n19059, n19061, n19062, n19063, n19064, n19065, n19066, n19067, n19068,
    n19069, n19071, n19072, n19073, n19074, n19075, n19076, n19077, n19078,
    n19080, n19081, n19082, n19083, n19084, n19085, n19086, n19087, n19088,
    n19089, n19090, n19092, n19093, n19094, n19095, n19096, n19098, n19099,
    n19100, n19101, n19102, n19104, n19105, n19106, n19107, n19108, n19109,
    n19110, n19111, n19112, n19114, n19115, n19116, n19117, n19118, n19119,
    n19120, n19121, n19122, n19123, n19125, n19126, n19127, n19128, n19129,
    n19130, n19131, n19132, n19133, n19135, n19136, n19137, n19138, n19139,
    n19140, n19141, n19142, n19143, n19145, n19146, n19147, n19148, n19149,
    n19150, n19151, n19152, n19153, n19155, n19156, n19157, n19158, n19159,
    n19160, n19161, n19162, n19163, n19165, n19166, n19167, n19168, n19169,
    n19170, n19171, n19172, n19173, n19175, n19176, n19177, n19178, n19179,
    n19180, n19181, n19182, n19183, n19185, n19186, n19187, n19188, n19189,
    n19190, n19191, n19192, n19193, n19195, n19196, n19197, n19198, n19199,
    n19200, n19201, n19202, n19203, n19205, n19206, n19207, n19208, n19209,
    n19210, n19211, n19212, n19213, n19215, n19216, n19217, n19218, n19219,
    n19220, n19221, n19222, n19223, n19225, n19226, n19227, n19228, n19229,
    n19230, n19231, n19232, n19233, n19235, n19236, n19237, n19238, n19239,
    n19240, n19241, n19242, n19243, n19245, n19246, n19247, n19248, n19249,
    n19250, n19251, n19252, n19253, n19255, n19256, n19257, n19258, n19259,
    n19260, n19261, n19262, n19263, n19265, n19266, n19267, n19268, n19269,
    n19270, n19271, n19272, n19274, n19275, n19276, n19277, n19278, n19279,
    n19280, n19281, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
    n19290, n19292, n19293, n19294, n19295, n19296, n19297, n19298, n19299,
    n19301, n19302, n19303, n19304, n19305, n19306, n19307, n19308, n19310,
    n19311, n19312, n19313, n19314, n19315, n19316, n19317, n19319, n19320,
    n19321, n19322, n19323, n19324, n19325, n19326, n19328, n19329, n19330,
    n19331, n19332, n19333, n19334, n19335, n19336, n19338, n19339, n19340,
    n19341, n19342, n19343, n19344, n19345, n19346, n19348, n19349, n19350,
    n19351, n19352, n19353, n19354, n19355, n19356, n19358, n19359, n19360,
    n19361, n19362, n19363, n19364, n19365, n19367, n19368, n19369, n19370,
    n19371, n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379,
    n19380, n19381, n19382, n19383, n19385, n19386, n19387, n19388, n19390,
    n19391, n19393, n19395, n19397, n19399, n19400, n19402, n19404, n19405,
    n19406, n19407, n19408, n19409, n19410, n19412, n19413, n19414, n19416,
    n19417, n19419, n19420, n19422, n19424, n19425, n19426, n19428, n19429,
    n19430;
  INVX1   g00000(.A(P3_DATAO_REG_31__SCAN_IN), .Y(n2964));
  NAND2X1 g00001(.A(n2964), .B(P3_DATAO_REG_30__SCAN_IN), .Y(n2965));
  INVX1   g00002(.A(P1_DATAO_REG_31__SCAN_IN), .Y(n2966));
  INVX1   g00003(.A(P2_DATAO_REG_31__SCAN_IN), .Y(n2967));
  AOI22X1 g00004(.A0(P2_DATAO_REG_30__SCAN_IN), .A1(n2967), .B0(P1_DATAO_REG_30__SCAN_IN), .B1(n2966), .Y(n2968));
  NAND3X1 g00005(.A(n2968), .B(n2965), .C(P3_ADDRESS_REG_29__SCAN_IN), .Y(n2969));
  NAND2X1 g00006(.A(n2968), .B(n2965), .Y(n2970));
  NAND2X1 g00007(.A(n2970), .B(P2_ADDRESS_REG_29__SCAN_IN), .Y(n2971));
  NAND2X1 g00008(.A(n2971), .B(n2969), .Y(U355));
  NAND3X1 g00009(.A(n2968), .B(n2965), .C(P3_ADDRESS_REG_28__SCAN_IN), .Y(n2973));
  NAND2X1 g00010(.A(n2970), .B(P2_ADDRESS_REG_28__SCAN_IN), .Y(n2974));
  NAND2X1 g00011(.A(n2974), .B(n2973), .Y(U356));
  NAND3X1 g00012(.A(n2968), .B(n2965), .C(P3_ADDRESS_REG_27__SCAN_IN), .Y(n2976));
  NAND2X1 g00013(.A(n2970), .B(P2_ADDRESS_REG_27__SCAN_IN), .Y(n2977));
  NAND2X1 g00014(.A(n2977), .B(n2976), .Y(U357));
  NAND3X1 g00015(.A(n2968), .B(n2965), .C(P3_ADDRESS_REG_26__SCAN_IN), .Y(n2979));
  NAND2X1 g00016(.A(n2970), .B(P2_ADDRESS_REG_26__SCAN_IN), .Y(n2980));
  NAND2X1 g00017(.A(n2980), .B(n2979), .Y(U358));
  NAND3X1 g00018(.A(n2968), .B(n2965), .C(P3_ADDRESS_REG_25__SCAN_IN), .Y(n2982));
  NAND2X1 g00019(.A(n2970), .B(P2_ADDRESS_REG_25__SCAN_IN), .Y(n2983));
  NAND2X1 g00020(.A(n2983), .B(n2982), .Y(U359));
  NAND3X1 g00021(.A(n2968), .B(n2965), .C(P3_ADDRESS_REG_24__SCAN_IN), .Y(n2985));
  NAND2X1 g00022(.A(n2970), .B(P2_ADDRESS_REG_24__SCAN_IN), .Y(n2986));
  NAND2X1 g00023(.A(n2986), .B(n2985), .Y(U360));
  NAND3X1 g00024(.A(n2968), .B(n2965), .C(P3_ADDRESS_REG_23__SCAN_IN), .Y(n2988));
  NAND2X1 g00025(.A(n2970), .B(P2_ADDRESS_REG_23__SCAN_IN), .Y(n2989));
  NAND2X1 g00026(.A(n2989), .B(n2988), .Y(U361));
  NAND3X1 g00027(.A(n2968), .B(n2965), .C(P3_ADDRESS_REG_22__SCAN_IN), .Y(n2991));
  NAND2X1 g00028(.A(n2970), .B(P2_ADDRESS_REG_22__SCAN_IN), .Y(n2992));
  NAND2X1 g00029(.A(n2992), .B(n2991), .Y(U362));
  NAND3X1 g00030(.A(n2968), .B(n2965), .C(P3_ADDRESS_REG_21__SCAN_IN), .Y(n2994));
  NAND2X1 g00031(.A(n2970), .B(P2_ADDRESS_REG_21__SCAN_IN), .Y(n2995));
  NAND2X1 g00032(.A(n2995), .B(n2994), .Y(U363));
  NAND3X1 g00033(.A(n2968), .B(n2965), .C(P3_ADDRESS_REG_20__SCAN_IN), .Y(n2997));
  NAND2X1 g00034(.A(n2970), .B(P2_ADDRESS_REG_20__SCAN_IN), .Y(n2998));
  NAND2X1 g00035(.A(n2998), .B(n2997), .Y(U364));
  NAND3X1 g00036(.A(n2968), .B(n2965), .C(P3_ADDRESS_REG_19__SCAN_IN), .Y(n3000));
  NAND2X1 g00037(.A(n2970), .B(P2_ADDRESS_REG_19__SCAN_IN), .Y(n3001));
  NAND2X1 g00038(.A(n3001), .B(n3000), .Y(U366));
  NAND3X1 g00039(.A(n2968), .B(n2965), .C(P3_ADDRESS_REG_18__SCAN_IN), .Y(n3003));
  NAND2X1 g00040(.A(n2970), .B(P2_ADDRESS_REG_18__SCAN_IN), .Y(n3004));
  NAND2X1 g00041(.A(n3004), .B(n3003), .Y(U367));
  NAND3X1 g00042(.A(n2968), .B(n2965), .C(P3_ADDRESS_REG_17__SCAN_IN), .Y(n3006));
  NAND2X1 g00043(.A(n2970), .B(P2_ADDRESS_REG_17__SCAN_IN), .Y(n3007));
  NAND2X1 g00044(.A(n3007), .B(n3006), .Y(U368));
  NAND3X1 g00045(.A(n2968), .B(n2965), .C(P3_ADDRESS_REG_16__SCAN_IN), .Y(n3009));
  NAND2X1 g00046(.A(n2970), .B(P2_ADDRESS_REG_16__SCAN_IN), .Y(n3010));
  NAND2X1 g00047(.A(n3010), .B(n3009), .Y(U369));
  NAND3X1 g00048(.A(n2968), .B(n2965), .C(P3_ADDRESS_REG_15__SCAN_IN), .Y(n3012));
  NAND2X1 g00049(.A(n2970), .B(P2_ADDRESS_REG_15__SCAN_IN), .Y(n3013));
  NAND2X1 g00050(.A(n3013), .B(n3012), .Y(U370));
  NAND3X1 g00051(.A(n2968), .B(n2965), .C(P3_ADDRESS_REG_14__SCAN_IN), .Y(n3015));
  NAND2X1 g00052(.A(n2970), .B(P2_ADDRESS_REG_14__SCAN_IN), .Y(n3016));
  NAND2X1 g00053(.A(n3016), .B(n3015), .Y(U371));
  NAND3X1 g00054(.A(n2968), .B(n2965), .C(P3_ADDRESS_REG_13__SCAN_IN), .Y(n3018));
  NAND2X1 g00055(.A(n2970), .B(P2_ADDRESS_REG_13__SCAN_IN), .Y(n3019));
  NAND2X1 g00056(.A(n3019), .B(n3018), .Y(U372));
  NAND3X1 g00057(.A(n2968), .B(n2965), .C(P3_ADDRESS_REG_12__SCAN_IN), .Y(n3021));
  NAND2X1 g00058(.A(n2970), .B(P2_ADDRESS_REG_12__SCAN_IN), .Y(n3022));
  NAND2X1 g00059(.A(n3022), .B(n3021), .Y(U373));
  NAND3X1 g00060(.A(n2968), .B(n2965), .C(P3_ADDRESS_REG_11__SCAN_IN), .Y(n3024));
  NAND2X1 g00061(.A(n2970), .B(P2_ADDRESS_REG_11__SCAN_IN), .Y(n3025));
  NAND2X1 g00062(.A(n3025), .B(n3024), .Y(U374));
  NAND3X1 g00063(.A(n2968), .B(n2965), .C(P3_ADDRESS_REG_10__SCAN_IN), .Y(n3027));
  NAND2X1 g00064(.A(n2970), .B(P2_ADDRESS_REG_10__SCAN_IN), .Y(n3028));
  NAND2X1 g00065(.A(n3028), .B(n3027), .Y(U375));
  NAND3X1 g00066(.A(n2968), .B(n2965), .C(P3_ADDRESS_REG_9__SCAN_IN), .Y(n3030));
  NAND2X1 g00067(.A(n2970), .B(P2_ADDRESS_REG_9__SCAN_IN), .Y(n3031));
  NAND2X1 g00068(.A(n3031), .B(n3030), .Y(U347));
  NAND3X1 g00069(.A(n2968), .B(n2965), .C(P3_ADDRESS_REG_8__SCAN_IN), .Y(n3033));
  NAND2X1 g00070(.A(n2970), .B(P2_ADDRESS_REG_8__SCAN_IN), .Y(n3034));
  NAND2X1 g00071(.A(n3034), .B(n3033), .Y(U348));
  NAND3X1 g00072(.A(n2968), .B(n2965), .C(P3_ADDRESS_REG_7__SCAN_IN), .Y(n3036));
  NAND2X1 g00073(.A(n2970), .B(P2_ADDRESS_REG_7__SCAN_IN), .Y(n3037));
  NAND2X1 g00074(.A(n3037), .B(n3036), .Y(U349));
  NAND3X1 g00075(.A(n2968), .B(n2965), .C(P3_ADDRESS_REG_6__SCAN_IN), .Y(n3039));
  NAND2X1 g00076(.A(n2970), .B(P2_ADDRESS_REG_6__SCAN_IN), .Y(n3040));
  NAND2X1 g00077(.A(n3040), .B(n3039), .Y(U350));
  NAND3X1 g00078(.A(n2968), .B(n2965), .C(P3_ADDRESS_REG_5__SCAN_IN), .Y(n3042));
  NAND2X1 g00079(.A(n2970), .B(P2_ADDRESS_REG_5__SCAN_IN), .Y(n3043));
  NAND2X1 g00080(.A(n3043), .B(n3042), .Y(U351));
  NAND3X1 g00081(.A(n2968), .B(n2965), .C(P3_ADDRESS_REG_4__SCAN_IN), .Y(n3045));
  NAND2X1 g00082(.A(n2970), .B(P2_ADDRESS_REG_4__SCAN_IN), .Y(n3046));
  NAND2X1 g00083(.A(n3046), .B(n3045), .Y(U352));
  NAND3X1 g00084(.A(n2968), .B(n2965), .C(P3_ADDRESS_REG_3__SCAN_IN), .Y(n3048));
  NAND2X1 g00085(.A(n2970), .B(P2_ADDRESS_REG_3__SCAN_IN), .Y(n3049));
  NAND2X1 g00086(.A(n3049), .B(n3048), .Y(U353));
  NAND3X1 g00087(.A(n2968), .B(n2965), .C(P3_ADDRESS_REG_2__SCAN_IN), .Y(n3051));
  NAND2X1 g00088(.A(n2970), .B(P2_ADDRESS_REG_2__SCAN_IN), .Y(n3052));
  NAND2X1 g00089(.A(n3052), .B(n3051), .Y(U354));
  NAND3X1 g00090(.A(n2968), .B(n2965), .C(P3_ADDRESS_REG_1__SCAN_IN), .Y(n3054));
  NAND2X1 g00091(.A(n2970), .B(P2_ADDRESS_REG_1__SCAN_IN), .Y(n3055));
  NAND2X1 g00092(.A(n3055), .B(n3054), .Y(U365));
  NAND3X1 g00093(.A(n2968), .B(n2965), .C(P3_ADDRESS_REG_0__SCAN_IN), .Y(n3057));
  NAND2X1 g00094(.A(n2970), .B(P2_ADDRESS_REG_0__SCAN_IN), .Y(n3058));
  NAND2X1 g00095(.A(n3058), .B(n3057), .Y(U376));
  NOR4X1  g00096(.A(P1_ADDRESS_REG_11__SCAN_IN), .B(P1_ADDRESS_REG_17__SCAN_IN), .C(P1_ADDRESS_REG_23__SCAN_IN), .D(P1_ADDRESS_REG_1__SCAN_IN), .Y(n3060));
  NOR4X1  g00097(.A(P1_ADDRESS_REG_8__SCAN_IN), .B(P1_ADDRESS_REG_16__SCAN_IN), .C(P1_ADDRESS_REG_18__SCAN_IN), .D(P1_ADDRESS_REG_0__SCAN_IN), .Y(n3061));
  NOR3X1  g00098(.A(P1_ADDRESS_REG_10__SCAN_IN), .B(P1_ADDRESS_REG_19__SCAN_IN), .C(P1_ADDRESS_REG_24__SCAN_IN), .Y(n3062));
  NOR4X1  g00099(.A(P1_ADDRESS_REG_9__SCAN_IN), .B(P1_ADDRESS_REG_22__SCAN_IN), .C(P1_ADDRESS_REG_25__SCAN_IN), .D(P1_ADDRESS_REG_7__SCAN_IN), .Y(n3063));
  NAND4X1 g00100(.A(n3062), .B(n3061), .C(n3060), .D(n3063), .Y(n3064));
  NOR2X1  g00101(.A(P1_ADDRESS_REG_26__SCAN_IN), .B(P1_ADDRESS_REG_28__SCAN_IN), .Y(n3065));
  NOR4X1  g00102(.A(P1_ADDRESS_REG_12__SCAN_IN), .B(P1_ADDRESS_REG_14__SCAN_IN), .C(P1_ADDRESS_REG_21__SCAN_IN), .D(P1_ADDRESS_REG_6__SCAN_IN), .Y(n3066));
  NOR4X1  g00103(.A(P1_ADDRESS_REG_3__SCAN_IN), .B(P1_ADDRESS_REG_5__SCAN_IN), .C(P1_ADDRESS_REG_15__SCAN_IN), .D(P1_ADDRESS_REG_2__SCAN_IN), .Y(n3067));
  NOR4X1  g00104(.A(P1_ADDRESS_REG_13__SCAN_IN), .B(P1_ADDRESS_REG_20__SCAN_IN), .C(P1_ADDRESS_REG_27__SCAN_IN), .D(P1_ADDRESS_REG_4__SCAN_IN), .Y(n3068));
  NAND4X1 g00105(.A(n3067), .B(n3066), .C(n3065), .D(n3068), .Y(n3069));
  OAI21X1 g00106(.A0(n3069), .A1(n3064), .B0(P1_ADDRESS_REG_29__SCAN_IN), .Y(n3070));
  NOR2X1  g00107(.A(P1_BE_N_REG_2__SCAN_IN), .B(P1_ADS_N_REG_SCAN_IN), .Y(n3071));
  NOR4X1  g00108(.A(P1_BE_N_REG_1__SCAN_IN), .B(P1_BE_N_REG_3__SCAN_IN), .C(P1_D_C_N_REG_SCAN_IN), .D(P1_BE_N_REG_0__SCAN_IN), .Y(n3072));
  NAND4X1 g00109(.A(n3071), .B(P1_W_R_N_REG_SCAN_IN), .C(P1_M_IO_N_REG_SCAN_IN), .D(n3072), .Y(n3073));
  NOR2X1  g00110(.A(n3073), .B(n3070), .Y(n3074));
  INVX1   g00111(.A(n3074), .Y(U214));
  NOR4X1  g00112(.A(P2_ADDRESS_REG_11__SCAN_IN), .B(P2_ADDRESS_REG_17__SCAN_IN), .C(P2_ADDRESS_REG_23__SCAN_IN), .D(P2_ADDRESS_REG_1__SCAN_IN), .Y(n3076));
  NOR4X1  g00113(.A(P2_ADDRESS_REG_8__SCAN_IN), .B(P2_ADDRESS_REG_16__SCAN_IN), .C(P2_ADDRESS_REG_18__SCAN_IN), .D(P2_ADDRESS_REG_0__SCAN_IN), .Y(n3077));
  NOR3X1  g00114(.A(P2_ADDRESS_REG_10__SCAN_IN), .B(P2_ADDRESS_REG_19__SCAN_IN), .C(P2_ADDRESS_REG_24__SCAN_IN), .Y(n3078));
  NOR4X1  g00115(.A(P2_ADDRESS_REG_9__SCAN_IN), .B(P2_ADDRESS_REG_22__SCAN_IN), .C(P2_ADDRESS_REG_25__SCAN_IN), .D(P2_ADDRESS_REG_7__SCAN_IN), .Y(n3079));
  NAND4X1 g00116(.A(n3078), .B(n3077), .C(n3076), .D(n3079), .Y(n3080));
  NOR2X1  g00117(.A(P2_ADDRESS_REG_26__SCAN_IN), .B(P2_ADDRESS_REG_28__SCAN_IN), .Y(n3081));
  NOR4X1  g00118(.A(P2_ADDRESS_REG_12__SCAN_IN), .B(P2_ADDRESS_REG_14__SCAN_IN), .C(P2_ADDRESS_REG_21__SCAN_IN), .D(P2_ADDRESS_REG_6__SCAN_IN), .Y(n3082));
  NOR4X1  g00119(.A(P2_ADDRESS_REG_3__SCAN_IN), .B(P2_ADDRESS_REG_5__SCAN_IN), .C(P2_ADDRESS_REG_15__SCAN_IN), .D(P2_ADDRESS_REG_2__SCAN_IN), .Y(n3083));
  NOR4X1  g00120(.A(P2_ADDRESS_REG_13__SCAN_IN), .B(P2_ADDRESS_REG_20__SCAN_IN), .C(P2_ADDRESS_REG_27__SCAN_IN), .D(P2_ADDRESS_REG_4__SCAN_IN), .Y(n3084));
  NAND4X1 g00121(.A(n3083), .B(n3082), .C(n3081), .D(n3084), .Y(n3085));
  OAI21X1 g00122(.A0(n3085), .A1(n3080), .B0(P2_ADDRESS_REG_29__SCAN_IN), .Y(n3086));
  INVX1   g00123(.A(P2_W_R_N_REG_SCAN_IN), .Y(n3087));
  NOR4X1  g00124(.A(P2_D_C_N_REG_SCAN_IN), .B(n3087), .C(P2_BE_N_REG_3__SCAN_IN), .D(P2_ADS_N_REG_SCAN_IN), .Y(n3088));
  INVX1   g00125(.A(P2_M_IO_N_REG_SCAN_IN), .Y(n3089));
  NOR4X1  g00126(.A(P2_BE_N_REG_0__SCAN_IN), .B(P2_BE_N_REG_1__SCAN_IN), .C(P2_BE_N_REG_2__SCAN_IN), .D(n3089), .Y(n3090));
  NAND2X1 g00127(.A(n3090), .B(n3088), .Y(n3091));
  OAI22X1 g00128(.A0(n3086), .A1(n3091), .B0(n3073), .B1(n3070), .Y(n3092));
  NAND3X1 g00129(.A(n3092), .B(U214), .C(P2_DATAO_REG_0__SCAN_IN), .Y(n3093));
  INVX1   g00130(.A(n3092), .Y(n3094));
  AOI22X1 g00131(.A0(n3074), .A1(P1_DATAO_REG_0__SCAN_IN), .B0(BUF1_REG_0__SCAN_IN), .B1(n3094), .Y(n3095));
  NAND2X1 g00132(.A(n3095), .B(n3093), .Y(U247));
  NAND3X1 g00133(.A(n3092), .B(U214), .C(P2_DATAO_REG_1__SCAN_IN), .Y(n3097));
  AOI22X1 g00134(.A0(n3074), .A1(P1_DATAO_REG_1__SCAN_IN), .B0(BUF1_REG_1__SCAN_IN), .B1(n3094), .Y(n3098));
  NAND2X1 g00135(.A(n3098), .B(n3097), .Y(U246));
  NAND3X1 g00136(.A(n3092), .B(U214), .C(P2_DATAO_REG_2__SCAN_IN), .Y(n3100));
  AOI22X1 g00137(.A0(n3074), .A1(P1_DATAO_REG_2__SCAN_IN), .B0(BUF1_REG_2__SCAN_IN), .B1(n3094), .Y(n3101));
  NAND2X1 g00138(.A(n3101), .B(n3100), .Y(U245));
  NAND3X1 g00139(.A(n3092), .B(U214), .C(P2_DATAO_REG_3__SCAN_IN), .Y(n3103));
  AOI22X1 g00140(.A0(n3074), .A1(P1_DATAO_REG_3__SCAN_IN), .B0(BUF1_REG_3__SCAN_IN), .B1(n3094), .Y(n3104));
  NAND2X1 g00141(.A(n3104), .B(n3103), .Y(U244));
  NAND3X1 g00142(.A(n3092), .B(U214), .C(P2_DATAO_REG_4__SCAN_IN), .Y(n3106));
  AOI22X1 g00143(.A0(n3074), .A1(P1_DATAO_REG_4__SCAN_IN), .B0(BUF1_REG_4__SCAN_IN), .B1(n3094), .Y(n3107));
  NAND2X1 g00144(.A(n3107), .B(n3106), .Y(U243));
  NAND3X1 g00145(.A(n3092), .B(U214), .C(P2_DATAO_REG_5__SCAN_IN), .Y(n3109));
  AOI22X1 g00146(.A0(n3074), .A1(P1_DATAO_REG_5__SCAN_IN), .B0(BUF1_REG_5__SCAN_IN), .B1(n3094), .Y(n3110));
  NAND2X1 g00147(.A(n3110), .B(n3109), .Y(U242));
  NAND3X1 g00148(.A(n3092), .B(U214), .C(P2_DATAO_REG_6__SCAN_IN), .Y(n3112));
  AOI22X1 g00149(.A0(n3074), .A1(P1_DATAO_REG_6__SCAN_IN), .B0(BUF1_REG_6__SCAN_IN), .B1(n3094), .Y(n3113));
  NAND2X1 g00150(.A(n3113), .B(n3112), .Y(U241));
  NAND3X1 g00151(.A(n3092), .B(U214), .C(P2_DATAO_REG_7__SCAN_IN), .Y(n3115));
  AOI22X1 g00152(.A0(n3074), .A1(P1_DATAO_REG_7__SCAN_IN), .B0(BUF1_REG_7__SCAN_IN), .B1(n3094), .Y(n3116));
  NAND2X1 g00153(.A(n3116), .B(n3115), .Y(U240));
  NAND3X1 g00154(.A(n3092), .B(U214), .C(P2_DATAO_REG_8__SCAN_IN), .Y(n3118));
  AOI22X1 g00155(.A0(n3074), .A1(P1_DATAO_REG_8__SCAN_IN), .B0(BUF1_REG_8__SCAN_IN), .B1(n3094), .Y(n3119));
  NAND2X1 g00156(.A(n3119), .B(n3118), .Y(U239));
  NAND3X1 g00157(.A(n3092), .B(U214), .C(P2_DATAO_REG_9__SCAN_IN), .Y(n3121));
  AOI22X1 g00158(.A0(n3074), .A1(P1_DATAO_REG_9__SCAN_IN), .B0(BUF1_REG_9__SCAN_IN), .B1(n3094), .Y(n3122));
  NAND2X1 g00159(.A(n3122), .B(n3121), .Y(U238));
  NAND3X1 g00160(.A(n3092), .B(U214), .C(P2_DATAO_REG_10__SCAN_IN), .Y(n3124));
  AOI22X1 g00161(.A0(n3074), .A1(P1_DATAO_REG_10__SCAN_IN), .B0(BUF1_REG_10__SCAN_IN), .B1(n3094), .Y(n3125));
  NAND2X1 g00162(.A(n3125), .B(n3124), .Y(U237));
  NAND3X1 g00163(.A(n3092), .B(U214), .C(P2_DATAO_REG_11__SCAN_IN), .Y(n3127));
  AOI22X1 g00164(.A0(n3074), .A1(P1_DATAO_REG_11__SCAN_IN), .B0(BUF1_REG_11__SCAN_IN), .B1(n3094), .Y(n3128));
  NAND2X1 g00165(.A(n3128), .B(n3127), .Y(U236));
  NAND3X1 g00166(.A(n3092), .B(U214), .C(P2_DATAO_REG_12__SCAN_IN), .Y(n3130));
  AOI22X1 g00167(.A0(n3074), .A1(P1_DATAO_REG_12__SCAN_IN), .B0(BUF1_REG_12__SCAN_IN), .B1(n3094), .Y(n3131));
  NAND2X1 g00168(.A(n3131), .B(n3130), .Y(U235));
  NAND3X1 g00169(.A(n3092), .B(U214), .C(P2_DATAO_REG_13__SCAN_IN), .Y(n3133));
  AOI22X1 g00170(.A0(n3074), .A1(P1_DATAO_REG_13__SCAN_IN), .B0(BUF1_REG_13__SCAN_IN), .B1(n3094), .Y(n3134));
  NAND2X1 g00171(.A(n3134), .B(n3133), .Y(U234));
  NAND3X1 g00172(.A(n3092), .B(U214), .C(P2_DATAO_REG_14__SCAN_IN), .Y(n3136));
  AOI22X1 g00173(.A0(n3074), .A1(P1_DATAO_REG_14__SCAN_IN), .B0(BUF1_REG_14__SCAN_IN), .B1(n3094), .Y(n3137));
  NAND2X1 g00174(.A(n3137), .B(n3136), .Y(U233));
  NAND3X1 g00175(.A(n3092), .B(U214), .C(P2_DATAO_REG_15__SCAN_IN), .Y(n3139));
  AOI22X1 g00176(.A0(n3074), .A1(P1_DATAO_REG_15__SCAN_IN), .B0(BUF1_REG_15__SCAN_IN), .B1(n3094), .Y(n3140));
  NAND2X1 g00177(.A(n3140), .B(n3139), .Y(U232));
  NAND3X1 g00178(.A(n3092), .B(U214), .C(P2_DATAO_REG_16__SCAN_IN), .Y(n3142));
  AOI22X1 g00179(.A0(n3074), .A1(P1_DATAO_REG_16__SCAN_IN), .B0(BUF1_REG_16__SCAN_IN), .B1(n3094), .Y(n3143));
  NAND2X1 g00180(.A(n3143), .B(n3142), .Y(U231));
  NAND3X1 g00181(.A(n3092), .B(U214), .C(P2_DATAO_REG_17__SCAN_IN), .Y(n3145));
  AOI22X1 g00182(.A0(n3074), .A1(P1_DATAO_REG_17__SCAN_IN), .B0(BUF1_REG_17__SCAN_IN), .B1(n3094), .Y(n3146));
  NAND2X1 g00183(.A(n3146), .B(n3145), .Y(U230));
  NAND3X1 g00184(.A(n3092), .B(U214), .C(P2_DATAO_REG_18__SCAN_IN), .Y(n3148));
  AOI22X1 g00185(.A0(n3074), .A1(P1_DATAO_REG_18__SCAN_IN), .B0(BUF1_REG_18__SCAN_IN), .B1(n3094), .Y(n3149));
  NAND2X1 g00186(.A(n3149), .B(n3148), .Y(U229));
  NAND3X1 g00187(.A(n3092), .B(U214), .C(P2_DATAO_REG_19__SCAN_IN), .Y(n3151));
  AOI22X1 g00188(.A0(n3074), .A1(P1_DATAO_REG_19__SCAN_IN), .B0(BUF1_REG_19__SCAN_IN), .B1(n3094), .Y(n3152));
  NAND2X1 g00189(.A(n3152), .B(n3151), .Y(U228));
  NAND3X1 g00190(.A(n3092), .B(U214), .C(P2_DATAO_REG_20__SCAN_IN), .Y(n3154));
  AOI22X1 g00191(.A0(n3074), .A1(P1_DATAO_REG_20__SCAN_IN), .B0(BUF1_REG_20__SCAN_IN), .B1(n3094), .Y(n3155));
  NAND2X1 g00192(.A(n3155), .B(n3154), .Y(U227));
  NAND3X1 g00193(.A(n3092), .B(U214), .C(P2_DATAO_REG_21__SCAN_IN), .Y(n3157));
  AOI22X1 g00194(.A0(n3074), .A1(P1_DATAO_REG_21__SCAN_IN), .B0(BUF1_REG_21__SCAN_IN), .B1(n3094), .Y(n3158));
  NAND2X1 g00195(.A(n3158), .B(n3157), .Y(U226));
  NAND3X1 g00196(.A(n3092), .B(U214), .C(P2_DATAO_REG_22__SCAN_IN), .Y(n3160));
  AOI22X1 g00197(.A0(n3074), .A1(P1_DATAO_REG_22__SCAN_IN), .B0(BUF1_REG_22__SCAN_IN), .B1(n3094), .Y(n3161));
  NAND2X1 g00198(.A(n3161), .B(n3160), .Y(U225));
  NAND3X1 g00199(.A(n3092), .B(U214), .C(P2_DATAO_REG_23__SCAN_IN), .Y(n3163));
  AOI22X1 g00200(.A0(n3074), .A1(P1_DATAO_REG_23__SCAN_IN), .B0(BUF1_REG_23__SCAN_IN), .B1(n3094), .Y(n3164));
  NAND2X1 g00201(.A(n3164), .B(n3163), .Y(U224));
  NAND3X1 g00202(.A(n3092), .B(U214), .C(P2_DATAO_REG_24__SCAN_IN), .Y(n3166));
  AOI22X1 g00203(.A0(n3074), .A1(P1_DATAO_REG_24__SCAN_IN), .B0(BUF1_REG_24__SCAN_IN), .B1(n3094), .Y(n3167));
  NAND2X1 g00204(.A(n3167), .B(n3166), .Y(U223));
  NAND3X1 g00205(.A(n3092), .B(U214), .C(P2_DATAO_REG_25__SCAN_IN), .Y(n3169));
  AOI22X1 g00206(.A0(n3074), .A1(P1_DATAO_REG_25__SCAN_IN), .B0(BUF1_REG_25__SCAN_IN), .B1(n3094), .Y(n3170));
  NAND2X1 g00207(.A(n3170), .B(n3169), .Y(U222));
  NAND3X1 g00208(.A(n3092), .B(U214), .C(P2_DATAO_REG_26__SCAN_IN), .Y(n3172));
  AOI22X1 g00209(.A0(n3074), .A1(P1_DATAO_REG_26__SCAN_IN), .B0(BUF1_REG_26__SCAN_IN), .B1(n3094), .Y(n3173));
  NAND2X1 g00210(.A(n3173), .B(n3172), .Y(U221));
  NAND3X1 g00211(.A(n3092), .B(U214), .C(P2_DATAO_REG_27__SCAN_IN), .Y(n3175));
  AOI22X1 g00212(.A0(n3074), .A1(P1_DATAO_REG_27__SCAN_IN), .B0(BUF1_REG_27__SCAN_IN), .B1(n3094), .Y(n3176));
  NAND2X1 g00213(.A(n3176), .B(n3175), .Y(U220));
  NAND3X1 g00214(.A(n3092), .B(U214), .C(P2_DATAO_REG_28__SCAN_IN), .Y(n3178));
  AOI22X1 g00215(.A0(n3074), .A1(P1_DATAO_REG_28__SCAN_IN), .B0(BUF1_REG_28__SCAN_IN), .B1(n3094), .Y(n3179));
  NAND2X1 g00216(.A(n3179), .B(n3178), .Y(U219));
  NAND3X1 g00217(.A(n3092), .B(U214), .C(P2_DATAO_REG_29__SCAN_IN), .Y(n3181));
  AOI22X1 g00218(.A0(n3074), .A1(P1_DATAO_REG_29__SCAN_IN), .B0(BUF1_REG_29__SCAN_IN), .B1(n3094), .Y(n3182));
  NAND2X1 g00219(.A(n3182), .B(n3181), .Y(U218));
  NAND3X1 g00220(.A(n3092), .B(U214), .C(P2_DATAO_REG_30__SCAN_IN), .Y(n3184));
  AOI22X1 g00221(.A0(n3074), .A1(P1_DATAO_REG_30__SCAN_IN), .B0(BUF1_REG_30__SCAN_IN), .B1(n3094), .Y(n3185));
  NAND2X1 g00222(.A(n3185), .B(n3184), .Y(U217));
  NAND3X1 g00223(.A(n3092), .B(U214), .C(P2_DATAO_REG_31__SCAN_IN), .Y(n3187));
  AOI22X1 g00224(.A0(n3074), .A1(P1_DATAO_REG_31__SCAN_IN), .B0(BUF1_REG_31__SCAN_IN), .B1(n3094), .Y(n3188));
  NAND2X1 g00225(.A(n3188), .B(n3187), .Y(U216));
  INVX1   g00226(.A(BUF2_REG_0__SCAN_IN), .Y(n3190));
  NOR2X1  g00227(.A(n3091), .B(P2_ADDRESS_REG_29__SCAN_IN), .Y(n3191));
  NAND2X1 g00228(.A(n3191), .B(P2_DATAO_REG_0__SCAN_IN), .Y(n3192));
  OAI21X1 g00229(.A0(n3191), .A1(n3190), .B0(n3192), .Y(U251));
  INVX1   g00230(.A(BUF2_REG_1__SCAN_IN), .Y(n3194));
  NAND2X1 g00231(.A(n3191), .B(P2_DATAO_REG_1__SCAN_IN), .Y(n3195));
  OAI21X1 g00232(.A0(n3191), .A1(n3194), .B0(n3195), .Y(U252));
  INVX1   g00233(.A(BUF2_REG_2__SCAN_IN), .Y(n3197));
  NAND2X1 g00234(.A(n3191), .B(P2_DATAO_REG_2__SCAN_IN), .Y(n3198));
  OAI21X1 g00235(.A0(n3191), .A1(n3197), .B0(n3198), .Y(U253));
  INVX1   g00236(.A(BUF2_REG_3__SCAN_IN), .Y(n3200));
  NAND2X1 g00237(.A(n3191), .B(P2_DATAO_REG_3__SCAN_IN), .Y(n3201));
  OAI21X1 g00238(.A0(n3191), .A1(n3200), .B0(n3201), .Y(U254));
  INVX1   g00239(.A(BUF2_REG_4__SCAN_IN), .Y(n3203));
  NAND2X1 g00240(.A(n3191), .B(P2_DATAO_REG_4__SCAN_IN), .Y(n3204));
  OAI21X1 g00241(.A0(n3191), .A1(n3203), .B0(n3204), .Y(U255));
  INVX1   g00242(.A(BUF2_REG_5__SCAN_IN), .Y(n3206));
  NAND2X1 g00243(.A(n3191), .B(P2_DATAO_REG_5__SCAN_IN), .Y(n3207));
  OAI21X1 g00244(.A0(n3191), .A1(n3206), .B0(n3207), .Y(U256));
  INVX1   g00245(.A(BUF2_REG_6__SCAN_IN), .Y(n3209));
  NAND2X1 g00246(.A(n3191), .B(P2_DATAO_REG_6__SCAN_IN), .Y(n3210));
  OAI21X1 g00247(.A0(n3191), .A1(n3209), .B0(n3210), .Y(U257));
  INVX1   g00248(.A(BUF2_REG_7__SCAN_IN), .Y(n3212));
  NAND2X1 g00249(.A(n3191), .B(P2_DATAO_REG_7__SCAN_IN), .Y(n3213));
  OAI21X1 g00250(.A0(n3191), .A1(n3212), .B0(n3213), .Y(U258));
  INVX1   g00251(.A(BUF2_REG_8__SCAN_IN), .Y(n3215));
  NAND2X1 g00252(.A(n3191), .B(P2_DATAO_REG_8__SCAN_IN), .Y(n3216));
  OAI21X1 g00253(.A0(n3191), .A1(n3215), .B0(n3216), .Y(U259));
  INVX1   g00254(.A(BUF2_REG_9__SCAN_IN), .Y(n3218));
  NAND2X1 g00255(.A(n3191), .B(P2_DATAO_REG_9__SCAN_IN), .Y(n3219));
  OAI21X1 g00256(.A0(n3191), .A1(n3218), .B0(n3219), .Y(U260));
  INVX1   g00257(.A(BUF2_REG_10__SCAN_IN), .Y(n3221));
  NAND2X1 g00258(.A(n3191), .B(P2_DATAO_REG_10__SCAN_IN), .Y(n3222));
  OAI21X1 g00259(.A0(n3191), .A1(n3221), .B0(n3222), .Y(U261));
  INVX1   g00260(.A(BUF2_REG_11__SCAN_IN), .Y(n3224));
  NAND2X1 g00261(.A(n3191), .B(P2_DATAO_REG_11__SCAN_IN), .Y(n3225));
  OAI21X1 g00262(.A0(n3191), .A1(n3224), .B0(n3225), .Y(U262));
  INVX1   g00263(.A(BUF2_REG_12__SCAN_IN), .Y(n3227));
  NAND2X1 g00264(.A(n3191), .B(P2_DATAO_REG_12__SCAN_IN), .Y(n3228));
  OAI21X1 g00265(.A0(n3191), .A1(n3227), .B0(n3228), .Y(U263));
  INVX1   g00266(.A(BUF2_REG_13__SCAN_IN), .Y(n3230));
  NAND2X1 g00267(.A(n3191), .B(P2_DATAO_REG_13__SCAN_IN), .Y(n3231));
  OAI21X1 g00268(.A0(n3191), .A1(n3230), .B0(n3231), .Y(U264));
  INVX1   g00269(.A(BUF2_REG_14__SCAN_IN), .Y(n3233));
  NAND2X1 g00270(.A(n3191), .B(P2_DATAO_REG_14__SCAN_IN), .Y(n3234));
  OAI21X1 g00271(.A0(n3191), .A1(n3233), .B0(n3234), .Y(U265));
  INVX1   g00272(.A(BUF2_REG_15__SCAN_IN), .Y(n3236));
  NAND2X1 g00273(.A(n3191), .B(P2_DATAO_REG_15__SCAN_IN), .Y(n3237));
  OAI21X1 g00274(.A0(n3191), .A1(n3236), .B0(n3237), .Y(U266));
  INVX1   g00275(.A(BUF2_REG_16__SCAN_IN), .Y(n3239));
  NAND2X1 g00276(.A(n3191), .B(P2_DATAO_REG_16__SCAN_IN), .Y(n3240));
  OAI21X1 g00277(.A0(n3191), .A1(n3239), .B0(n3240), .Y(U267));
  INVX1   g00278(.A(BUF2_REG_17__SCAN_IN), .Y(n3242));
  NAND2X1 g00279(.A(n3191), .B(P2_DATAO_REG_17__SCAN_IN), .Y(n3243));
  OAI21X1 g00280(.A0(n3191), .A1(n3242), .B0(n3243), .Y(U268));
  INVX1   g00281(.A(BUF2_REG_18__SCAN_IN), .Y(n3245));
  NAND2X1 g00282(.A(n3191), .B(P2_DATAO_REG_18__SCAN_IN), .Y(n3246));
  OAI21X1 g00283(.A0(n3191), .A1(n3245), .B0(n3246), .Y(U269));
  INVX1   g00284(.A(BUF2_REG_19__SCAN_IN), .Y(n3248));
  NAND2X1 g00285(.A(n3191), .B(P2_DATAO_REG_19__SCAN_IN), .Y(n3249));
  OAI21X1 g00286(.A0(n3191), .A1(n3248), .B0(n3249), .Y(U270));
  INVX1   g00287(.A(BUF2_REG_20__SCAN_IN), .Y(n3251));
  NAND2X1 g00288(.A(n3191), .B(P2_DATAO_REG_20__SCAN_IN), .Y(n3252));
  OAI21X1 g00289(.A0(n3191), .A1(n3251), .B0(n3252), .Y(U271));
  INVX1   g00290(.A(BUF2_REG_21__SCAN_IN), .Y(n3254));
  NAND2X1 g00291(.A(n3191), .B(P2_DATAO_REG_21__SCAN_IN), .Y(n3255));
  OAI21X1 g00292(.A0(n3191), .A1(n3254), .B0(n3255), .Y(U272));
  INVX1   g00293(.A(BUF2_REG_22__SCAN_IN), .Y(n3257));
  NAND2X1 g00294(.A(n3191), .B(P2_DATAO_REG_22__SCAN_IN), .Y(n3258));
  OAI21X1 g00295(.A0(n3191), .A1(n3257), .B0(n3258), .Y(U273));
  INVX1   g00296(.A(BUF2_REG_23__SCAN_IN), .Y(n3260));
  NAND2X1 g00297(.A(n3191), .B(P2_DATAO_REG_23__SCAN_IN), .Y(n3261));
  OAI21X1 g00298(.A0(n3191), .A1(n3260), .B0(n3261), .Y(U274));
  INVX1   g00299(.A(BUF2_REG_24__SCAN_IN), .Y(n3263));
  NAND2X1 g00300(.A(n3191), .B(P2_DATAO_REG_24__SCAN_IN), .Y(n3264));
  OAI21X1 g00301(.A0(n3191), .A1(n3263), .B0(n3264), .Y(U275));
  INVX1   g00302(.A(BUF2_REG_25__SCAN_IN), .Y(n3266));
  NAND2X1 g00303(.A(n3191), .B(P2_DATAO_REG_25__SCAN_IN), .Y(n3267));
  OAI21X1 g00304(.A0(n3191), .A1(n3266), .B0(n3267), .Y(U276));
  INVX1   g00305(.A(BUF2_REG_26__SCAN_IN), .Y(n3269));
  NAND2X1 g00306(.A(n3191), .B(P2_DATAO_REG_26__SCAN_IN), .Y(n3270));
  OAI21X1 g00307(.A0(n3191), .A1(n3269), .B0(n3270), .Y(U277));
  INVX1   g00308(.A(BUF2_REG_27__SCAN_IN), .Y(n3272));
  NAND2X1 g00309(.A(n3191), .B(P2_DATAO_REG_27__SCAN_IN), .Y(n3273));
  OAI21X1 g00310(.A0(n3191), .A1(n3272), .B0(n3273), .Y(U278));
  INVX1   g00311(.A(BUF2_REG_28__SCAN_IN), .Y(n3275));
  NAND2X1 g00312(.A(n3191), .B(P2_DATAO_REG_28__SCAN_IN), .Y(n3276));
  OAI21X1 g00313(.A0(n3191), .A1(n3275), .B0(n3276), .Y(U279));
  INVX1   g00314(.A(BUF2_REG_29__SCAN_IN), .Y(n3278));
  NAND2X1 g00315(.A(n3191), .B(P2_DATAO_REG_29__SCAN_IN), .Y(n3279));
  OAI21X1 g00316(.A0(n3191), .A1(n3278), .B0(n3279), .Y(U280));
  INVX1   g00317(.A(BUF2_REG_30__SCAN_IN), .Y(n3281));
  NAND2X1 g00318(.A(n3191), .B(P2_DATAO_REG_30__SCAN_IN), .Y(n3282));
  OAI21X1 g00319(.A0(n3191), .A1(n3281), .B0(n3282), .Y(U281));
  INVX1   g00320(.A(BUF2_REG_31__SCAN_IN), .Y(n3284));
  NAND2X1 g00321(.A(n3191), .B(P2_DATAO_REG_31__SCAN_IN), .Y(n3285));
  OAI21X1 g00322(.A0(n3191), .A1(n3284), .B0(n3285), .Y(U282));
  NOR2X1  g00323(.A(n3091), .B(n3086), .Y(n3287));
  OAI21X1 g00324(.A0(n3073), .A1(n3070), .B0(n3287), .Y(U212));
  INVX1   g00325(.A(n3191), .Y(U215));
  INVX1   g00326(.A(P3_M_IO_N_REG_SCAN_IN), .Y(n3290));
  NOR4X1  g00327(.A(n3290), .B(P3_BE_N_REG_2__SCAN_IN), .C(P3_BE_N_REG_3__SCAN_IN), .D(P3_ADS_N_REG_SCAN_IN), .Y(n3291));
  NOR4X1  g00328(.A(P3_W_R_N_REG_SCAN_IN), .B(P3_BE_N_REG_0__SCAN_IN), .C(P3_BE_N_REG_1__SCAN_IN), .D(P3_D_C_N_REG_SCAN_IN), .Y(n3292));
  NAND3X1 g00329(.A(n3292), .B(n3291), .C(U215), .Y(U213));
  INVX1   g00330(.A(P3_STATE_REG_0__SCAN_IN), .Y(n3294));
  NAND3X1 g00331(.A(P3_BYTEENABLE_REG_3__SCAN_IN), .B(n3294), .C(P3_STATE_REG_1__SCAN_IN), .Y(n3295));
  INVX1   g00332(.A(P3_STATE_REG_1__SCAN_IN), .Y(n3296));
  OAI21X1 g00333(.A0(P3_STATE_REG_0__SCAN_IN), .A1(n3296), .B0(P3_BE_N_REG_3__SCAN_IN), .Y(n3297));
  NAND2X1 g00334(.A(n3297), .B(n3295), .Y(P3_U3274));
  INVX1   g00335(.A(P3_BYTEENABLE_REG_2__SCAN_IN), .Y(n3299));
  NOR2X1  g00336(.A(P3_STATE_REG_0__SCAN_IN), .B(n3296), .Y(n3300));
  INVX1   g00337(.A(n3300), .Y(n3301));
  OAI21X1 g00338(.A0(P3_STATE_REG_0__SCAN_IN), .A1(n3296), .B0(P3_BE_N_REG_2__SCAN_IN), .Y(n3302));
  OAI21X1 g00339(.A0(n3301), .A1(n3299), .B0(n3302), .Y(P3_U3275));
  NAND3X1 g00340(.A(P3_BYTEENABLE_REG_1__SCAN_IN), .B(n3294), .C(P3_STATE_REG_1__SCAN_IN), .Y(n3304));
  OAI21X1 g00341(.A0(P3_STATE_REG_0__SCAN_IN), .A1(n3296), .B0(P3_BE_N_REG_1__SCAN_IN), .Y(n3305));
  NAND2X1 g00342(.A(n3305), .B(n3304), .Y(P3_U3276));
  INVX1   g00343(.A(P3_BYTEENABLE_REG_0__SCAN_IN), .Y(n3307));
  OAI21X1 g00344(.A0(P3_STATE_REG_0__SCAN_IN), .A1(n3296), .B0(P3_BE_N_REG_0__SCAN_IN), .Y(n3308));
  OAI21X1 g00345(.A0(n3301), .A1(n3307), .B0(n3308), .Y(P3_U3277));
  INVX1   g00346(.A(P3_REIP_REG_30__SCAN_IN), .Y(n3310));
  NAND3X1 g00347(.A(n3294), .B(P3_STATE_REG_1__SCAN_IN), .C(P3_STATE_REG_2__SCAN_IN), .Y(n3311));
  NOR3X1  g00348(.A(P3_STATE_REG_0__SCAN_IN), .B(n3296), .C(P3_STATE_REG_2__SCAN_IN), .Y(n3312));
  AOI22X1 g00349(.A0(n3301), .A1(P3_ADDRESS_REG_29__SCAN_IN), .B0(P3_REIP_REG_31__SCAN_IN), .B1(n3312), .Y(n3313));
  OAI21X1 g00350(.A0(n3311), .A1(n3310), .B0(n3313), .Y(P3_U3061));
  INVX1   g00351(.A(P3_REIP_REG_29__SCAN_IN), .Y(n3315));
  AOI22X1 g00352(.A0(n3301), .A1(P3_ADDRESS_REG_28__SCAN_IN), .B0(P3_REIP_REG_30__SCAN_IN), .B1(n3312), .Y(n3316));
  OAI21X1 g00353(.A0(n3311), .A1(n3315), .B0(n3316), .Y(P3_U3060));
  NAND4X1 g00354(.A(n3294), .B(P3_STATE_REG_1__SCAN_IN), .C(P3_STATE_REG_2__SCAN_IN), .D(P3_REIP_REG_28__SCAN_IN), .Y(n3318));
  AOI22X1 g00355(.A0(n3301), .A1(P3_ADDRESS_REG_27__SCAN_IN), .B0(P3_REIP_REG_29__SCAN_IN), .B1(n3312), .Y(n3319));
  NAND2X1 g00356(.A(n3319), .B(n3318), .Y(P3_U3059));
  INVX1   g00357(.A(P3_REIP_REG_27__SCAN_IN), .Y(n3321));
  AOI22X1 g00358(.A0(n3301), .A1(P3_ADDRESS_REG_26__SCAN_IN), .B0(P3_REIP_REG_28__SCAN_IN), .B1(n3312), .Y(n3322));
  OAI21X1 g00359(.A0(n3311), .A1(n3321), .B0(n3322), .Y(P3_U3058));
  INVX1   g00360(.A(P3_REIP_REG_26__SCAN_IN), .Y(n3324));
  AOI22X1 g00361(.A0(n3301), .A1(P3_ADDRESS_REG_25__SCAN_IN), .B0(P3_REIP_REG_27__SCAN_IN), .B1(n3312), .Y(n3325));
  OAI21X1 g00362(.A0(n3311), .A1(n3324), .B0(n3325), .Y(P3_U3057));
  INVX1   g00363(.A(P3_REIP_REG_25__SCAN_IN), .Y(n3327));
  AOI22X1 g00364(.A0(n3301), .A1(P3_ADDRESS_REG_24__SCAN_IN), .B0(P3_REIP_REG_26__SCAN_IN), .B1(n3312), .Y(n3328));
  OAI21X1 g00365(.A0(n3311), .A1(n3327), .B0(n3328), .Y(P3_U3056));
  INVX1   g00366(.A(P3_REIP_REG_24__SCAN_IN), .Y(n3330));
  AOI22X1 g00367(.A0(n3301), .A1(P3_ADDRESS_REG_23__SCAN_IN), .B0(P3_REIP_REG_25__SCAN_IN), .B1(n3312), .Y(n3331));
  OAI21X1 g00368(.A0(n3311), .A1(n3330), .B0(n3331), .Y(P3_U3055));
  INVX1   g00369(.A(P3_REIP_REG_23__SCAN_IN), .Y(n3333));
  AOI22X1 g00370(.A0(n3301), .A1(P3_ADDRESS_REG_22__SCAN_IN), .B0(P3_REIP_REG_24__SCAN_IN), .B1(n3312), .Y(n3334));
  OAI21X1 g00371(.A0(n3311), .A1(n3333), .B0(n3334), .Y(P3_U3054));
  INVX1   g00372(.A(P3_REIP_REG_22__SCAN_IN), .Y(n3336));
  AOI22X1 g00373(.A0(n3301), .A1(P3_ADDRESS_REG_21__SCAN_IN), .B0(P3_REIP_REG_23__SCAN_IN), .B1(n3312), .Y(n3337));
  OAI21X1 g00374(.A0(n3311), .A1(n3336), .B0(n3337), .Y(P3_U3053));
  INVX1   g00375(.A(P3_REIP_REG_21__SCAN_IN), .Y(n3339));
  AOI22X1 g00376(.A0(n3301), .A1(P3_ADDRESS_REG_20__SCAN_IN), .B0(P3_REIP_REG_22__SCAN_IN), .B1(n3312), .Y(n3340));
  OAI21X1 g00377(.A0(n3311), .A1(n3339), .B0(n3340), .Y(P3_U3052));
  INVX1   g00378(.A(P3_REIP_REG_20__SCAN_IN), .Y(n3342));
  AOI22X1 g00379(.A0(n3301), .A1(P3_ADDRESS_REG_19__SCAN_IN), .B0(P3_REIP_REG_21__SCAN_IN), .B1(n3312), .Y(n3343));
  OAI21X1 g00380(.A0(n3311), .A1(n3342), .B0(n3343), .Y(P3_U3051));
  INVX1   g00381(.A(P3_REIP_REG_19__SCAN_IN), .Y(n3345));
  AOI22X1 g00382(.A0(n3301), .A1(P3_ADDRESS_REG_18__SCAN_IN), .B0(P3_REIP_REG_20__SCAN_IN), .B1(n3312), .Y(n3346));
  OAI21X1 g00383(.A0(n3311), .A1(n3345), .B0(n3346), .Y(P3_U3050));
  INVX1   g00384(.A(P3_REIP_REG_18__SCAN_IN), .Y(n3348));
  AOI22X1 g00385(.A0(n3301), .A1(P3_ADDRESS_REG_17__SCAN_IN), .B0(P3_REIP_REG_19__SCAN_IN), .B1(n3312), .Y(n3349));
  OAI21X1 g00386(.A0(n3311), .A1(n3348), .B0(n3349), .Y(P3_U3049));
  INVX1   g00387(.A(P3_REIP_REG_17__SCAN_IN), .Y(n3351));
  AOI22X1 g00388(.A0(n3301), .A1(P3_ADDRESS_REG_16__SCAN_IN), .B0(P3_REIP_REG_18__SCAN_IN), .B1(n3312), .Y(n3352));
  OAI21X1 g00389(.A0(n3311), .A1(n3351), .B0(n3352), .Y(P3_U3048));
  INVX1   g00390(.A(P3_REIP_REG_16__SCAN_IN), .Y(n3354));
  AOI22X1 g00391(.A0(n3301), .A1(P3_ADDRESS_REG_15__SCAN_IN), .B0(P3_REIP_REG_17__SCAN_IN), .B1(n3312), .Y(n3355));
  OAI21X1 g00392(.A0(n3311), .A1(n3354), .B0(n3355), .Y(P3_U3047));
  INVX1   g00393(.A(P3_REIP_REG_15__SCAN_IN), .Y(n3357));
  AOI22X1 g00394(.A0(n3301), .A1(P3_ADDRESS_REG_14__SCAN_IN), .B0(P3_REIP_REG_16__SCAN_IN), .B1(n3312), .Y(n3358));
  OAI21X1 g00395(.A0(n3311), .A1(n3357), .B0(n3358), .Y(P3_U3046));
  INVX1   g00396(.A(P3_REIP_REG_14__SCAN_IN), .Y(n3360));
  AOI22X1 g00397(.A0(n3301), .A1(P3_ADDRESS_REG_13__SCAN_IN), .B0(P3_REIP_REG_15__SCAN_IN), .B1(n3312), .Y(n3361));
  OAI21X1 g00398(.A0(n3311), .A1(n3360), .B0(n3361), .Y(P3_U3045));
  INVX1   g00399(.A(P3_REIP_REG_13__SCAN_IN), .Y(n3363));
  AOI22X1 g00400(.A0(n3301), .A1(P3_ADDRESS_REG_12__SCAN_IN), .B0(P3_REIP_REG_14__SCAN_IN), .B1(n3312), .Y(n3364));
  OAI21X1 g00401(.A0(n3311), .A1(n3363), .B0(n3364), .Y(P3_U3044));
  INVX1   g00402(.A(P3_REIP_REG_12__SCAN_IN), .Y(n3366));
  AOI22X1 g00403(.A0(n3301), .A1(P3_ADDRESS_REG_11__SCAN_IN), .B0(P3_REIP_REG_13__SCAN_IN), .B1(n3312), .Y(n3367));
  OAI21X1 g00404(.A0(n3311), .A1(n3366), .B0(n3367), .Y(P3_U3043));
  INVX1   g00405(.A(P3_REIP_REG_11__SCAN_IN), .Y(n3369));
  AOI22X1 g00406(.A0(n3301), .A1(P3_ADDRESS_REG_10__SCAN_IN), .B0(P3_REIP_REG_12__SCAN_IN), .B1(n3312), .Y(n3370));
  OAI21X1 g00407(.A0(n3311), .A1(n3369), .B0(n3370), .Y(P3_U3042));
  INVX1   g00408(.A(P3_REIP_REG_10__SCAN_IN), .Y(n3372));
  AOI22X1 g00409(.A0(n3301), .A1(P3_ADDRESS_REG_9__SCAN_IN), .B0(P3_REIP_REG_11__SCAN_IN), .B1(n3312), .Y(n3373));
  OAI21X1 g00410(.A0(n3311), .A1(n3372), .B0(n3373), .Y(P3_U3041));
  INVX1   g00411(.A(P3_REIP_REG_9__SCAN_IN), .Y(n3375));
  AOI22X1 g00412(.A0(n3301), .A1(P3_ADDRESS_REG_8__SCAN_IN), .B0(P3_REIP_REG_10__SCAN_IN), .B1(n3312), .Y(n3376));
  OAI21X1 g00413(.A0(n3311), .A1(n3375), .B0(n3376), .Y(P3_U3040));
  INVX1   g00414(.A(P3_REIP_REG_8__SCAN_IN), .Y(n3378));
  AOI22X1 g00415(.A0(n3301), .A1(P3_ADDRESS_REG_7__SCAN_IN), .B0(P3_REIP_REG_9__SCAN_IN), .B1(n3312), .Y(n3379));
  OAI21X1 g00416(.A0(n3311), .A1(n3378), .B0(n3379), .Y(P3_U3039));
  INVX1   g00417(.A(P3_REIP_REG_7__SCAN_IN), .Y(n3381));
  AOI22X1 g00418(.A0(n3301), .A1(P3_ADDRESS_REG_6__SCAN_IN), .B0(P3_REIP_REG_8__SCAN_IN), .B1(n3312), .Y(n3382));
  OAI21X1 g00419(.A0(n3311), .A1(n3381), .B0(n3382), .Y(P3_U3038));
  INVX1   g00420(.A(P3_REIP_REG_6__SCAN_IN), .Y(n3384));
  AOI22X1 g00421(.A0(n3301), .A1(P3_ADDRESS_REG_5__SCAN_IN), .B0(P3_REIP_REG_7__SCAN_IN), .B1(n3312), .Y(n3385));
  OAI21X1 g00422(.A0(n3311), .A1(n3384), .B0(n3385), .Y(P3_U3037));
  INVX1   g00423(.A(P3_REIP_REG_5__SCAN_IN), .Y(n3387));
  AOI22X1 g00424(.A0(n3301), .A1(P3_ADDRESS_REG_4__SCAN_IN), .B0(P3_REIP_REG_6__SCAN_IN), .B1(n3312), .Y(n3388));
  OAI21X1 g00425(.A0(n3311), .A1(n3387), .B0(n3388), .Y(P3_U3036));
  INVX1   g00426(.A(P3_REIP_REG_4__SCAN_IN), .Y(n3390));
  AOI22X1 g00427(.A0(n3301), .A1(P3_ADDRESS_REG_3__SCAN_IN), .B0(P3_REIP_REG_5__SCAN_IN), .B1(n3312), .Y(n3391));
  OAI21X1 g00428(.A0(n3311), .A1(n3390), .B0(n3391), .Y(P3_U3035));
  INVX1   g00429(.A(P3_REIP_REG_3__SCAN_IN), .Y(n3393));
  AOI22X1 g00430(.A0(n3301), .A1(P3_ADDRESS_REG_2__SCAN_IN), .B0(P3_REIP_REG_4__SCAN_IN), .B1(n3312), .Y(n3394));
  OAI21X1 g00431(.A0(n3311), .A1(n3393), .B0(n3394), .Y(P3_U3034));
  INVX1   g00432(.A(P3_REIP_REG_2__SCAN_IN), .Y(n3396));
  AOI22X1 g00433(.A0(n3301), .A1(P3_ADDRESS_REG_1__SCAN_IN), .B0(P3_REIP_REG_3__SCAN_IN), .B1(n3312), .Y(n3397));
  OAI21X1 g00434(.A0(n3311), .A1(n3396), .B0(n3397), .Y(P3_U3033));
  INVX1   g00435(.A(P3_REIP_REG_1__SCAN_IN), .Y(n3399));
  AOI22X1 g00436(.A0(n3301), .A1(P3_ADDRESS_REG_0__SCAN_IN), .B0(P3_REIP_REG_2__SCAN_IN), .B1(n3312), .Y(n3400));
  OAI21X1 g00437(.A0(n3311), .A1(n3399), .B0(n3400), .Y(P3_U3032));
  INVX1   g00438(.A(P3_STATE_REG_2__SCAN_IN), .Y(n3402));
  INVX1   g00439(.A(READY2), .Y(n3403));
  INVX1   g00440(.A(READY22_REG_SCAN_IN), .Y(n3404));
  NOR2X1  g00441(.A(P3_REQUESTPENDING_REG_SCAN_IN), .B(HOLD), .Y(n3405));
  OAI21X1 g00442(.A0(n3404), .A1(n3403), .B0(n3405), .Y(n3406));
  NOR2X1  g00443(.A(n3404), .B(n3403), .Y(n3407));
  INVX1   g00444(.A(n3407), .Y(n3408));
  INVX1   g00445(.A(P3_REQUESTPENDING_REG_SCAN_IN), .Y(n3409));
  NOR2X1  g00446(.A(n3409), .B(HOLD), .Y(n3410));
  AOI21X1 g00447(.A0(n3410), .A1(n3408), .B0(n3296), .Y(n3411));
  NAND2X1 g00448(.A(P3_STATE_REG_0__SCAN_IN), .B(HOLD), .Y(n3412));
  OAI21X1 g00449(.A0(P3_STATE_REG_0__SCAN_IN), .A1(NA), .B0(n3412), .Y(n3413));
  AOI21X1 g00450(.A0(n3411), .A1(n3406), .B0(n3413), .Y(n3414));
  NAND4X1 g00451(.A(n3402), .B(READY22_REG_SCAN_IN), .C(READY2), .D(P3_STATE_REG_1__SCAN_IN), .Y(n3415));
  NOR2X1  g00452(.A(P3_STATE_REG_1__SCAN_IN), .B(P3_STATE_REG_2__SCAN_IN), .Y(n3416));
  NAND3X1 g00453(.A(n3416), .B(n3409), .C(HOLD), .Y(n3417));
  OAI21X1 g00454(.A0(n3415), .A1(n3405), .B0(n3417), .Y(n3418));
  INVX1   g00455(.A(NA), .Y(n3419));
  NOR3X1  g00456(.A(n3296), .B(P3_STATE_REG_2__SCAN_IN), .C(n3419), .Y(n3420));
  NOR2X1  g00457(.A(n3420), .B(n3294), .Y(n3421));
  AOI22X1 g00458(.A0(n3418), .A1(n3421), .B0(n3300), .B1(P3_STATE_REG_2__SCAN_IN), .Y(n3422));
  OAI21X1 g00459(.A0(n3414), .A1(n3402), .B0(n3422), .Y(P3_U3031));
  OAI21X1 g00460(.A0(n3410), .A1(n3294), .B0(P3_STATE_REG_2__SCAN_IN), .Y(n3424));
  NAND2X1 g00461(.A(P3_REQUESTPENDING_REG_SCAN_IN), .B(P3_STATE_REG_0__SCAN_IN), .Y(n3425));
  OAI21X1 g00462(.A0(n3425), .A1(P3_STATE_REG_2__SCAN_IN), .B0(n3424), .Y(n3426));
  NAND2X1 g00463(.A(n3426), .B(n3296), .Y(n3427));
  INVX1   g00464(.A(HOLD), .Y(n3428));
  AOI21X1 g00465(.A0(READY22_REG_SCAN_IN), .A1(READY2), .B0(n3428), .Y(n3429));
  OAI21X1 g00466(.A0(n3429), .A1(n3294), .B0(P3_STATE_REG_2__SCAN_IN), .Y(n3430));
  NAND3X1 g00467(.A(n3430), .B(n3406), .C(P3_STATE_REG_1__SCAN_IN), .Y(n3431));
  OAI21X1 g00468(.A0(n3407), .A1(n3402), .B0(n3300), .Y(n3432));
  NAND3X1 g00469(.A(n3432), .B(n3431), .C(n3427), .Y(P3_U3030));
  OAI21X1 g00470(.A0(n3425), .A1(n3411), .B0(n3402), .Y(n3434));
  OAI22X1 g00471(.A0(P3_STATE_REG_0__SCAN_IN), .A1(n3419), .B0(n3402), .B1(n3410), .Y(n3435));
  NOR3X1  g00472(.A(n3410), .B(n3294), .C(n3402), .Y(n3436));
  AOI21X1 g00473(.A0(n3435), .A1(n3296), .B0(n3436), .Y(n3437));
  NAND2X1 g00474(.A(n3437), .B(n3434), .Y(P3_U3029));
  INVX1   g00475(.A(BS16), .Y(n3439));
  OAI21X1 g00476(.A0(P3_STATE_REG_1__SCAN_IN), .A1(P3_STATE_REG_2__SCAN_IN), .B0(n3439), .Y(n3440));
  NOR3X1  g00477(.A(n3294), .B(n3296), .C(P3_STATE_REG_2__SCAN_IN), .Y(n3441));
  AOI21X1 g00478(.A0(n3294), .A1(n3296), .B0(n3441), .Y(n3442));
  NAND2X1 g00479(.A(n3442), .B(P3_DATAWIDTH_REG_0__SCAN_IN), .Y(n3443));
  OAI21X1 g00480(.A0(n3442), .A1(n3440), .B0(n3443), .Y(P3_U3280));
  INVX1   g00481(.A(P3_DATAWIDTH_REG_1__SCAN_IN), .Y(n3445));
  INVX1   g00482(.A(n3442), .Y(n3446));
  NAND2X1 g00483(.A(n3446), .B(n3440), .Y(n3447));
  OAI21X1 g00484(.A0(n3446), .A1(n3445), .B0(n3447), .Y(P3_U3281));
  INVX1   g00485(.A(P3_DATAWIDTH_REG_2__SCAN_IN), .Y(n3449));
  NOR2X1  g00486(.A(n3446), .B(n3449), .Y(P3_U3028));
  INVX1   g00487(.A(P3_DATAWIDTH_REG_3__SCAN_IN), .Y(n3451));
  NOR2X1  g00488(.A(n3446), .B(n3451), .Y(P3_U3027));
  INVX1   g00489(.A(P3_DATAWIDTH_REG_4__SCAN_IN), .Y(n3453));
  NOR2X1  g00490(.A(n3446), .B(n3453), .Y(P3_U3026));
  INVX1   g00491(.A(P3_DATAWIDTH_REG_5__SCAN_IN), .Y(n3455));
  NOR2X1  g00492(.A(n3446), .B(n3455), .Y(P3_U3025));
  INVX1   g00493(.A(P3_DATAWIDTH_REG_6__SCAN_IN), .Y(n3457));
  NOR2X1  g00494(.A(n3446), .B(n3457), .Y(P3_U3024));
  INVX1   g00495(.A(P3_DATAWIDTH_REG_7__SCAN_IN), .Y(n3459));
  NOR2X1  g00496(.A(n3446), .B(n3459), .Y(P3_U3023));
  INVX1   g00497(.A(P3_DATAWIDTH_REG_8__SCAN_IN), .Y(n3461));
  NOR2X1  g00498(.A(n3446), .B(n3461), .Y(P3_U3022));
  INVX1   g00499(.A(P3_DATAWIDTH_REG_9__SCAN_IN), .Y(n3463));
  NOR2X1  g00500(.A(n3446), .B(n3463), .Y(P3_U3021));
  INVX1   g00501(.A(P3_DATAWIDTH_REG_10__SCAN_IN), .Y(n3465));
  NOR2X1  g00502(.A(n3446), .B(n3465), .Y(P3_U3020));
  INVX1   g00503(.A(P3_DATAWIDTH_REG_11__SCAN_IN), .Y(n3467));
  NOR2X1  g00504(.A(n3446), .B(n3467), .Y(P3_U3019));
  INVX1   g00505(.A(P3_DATAWIDTH_REG_12__SCAN_IN), .Y(n3469));
  NOR2X1  g00506(.A(n3446), .B(n3469), .Y(P3_U3018));
  INVX1   g00507(.A(P3_DATAWIDTH_REG_13__SCAN_IN), .Y(n3471));
  NOR2X1  g00508(.A(n3446), .B(n3471), .Y(P3_U3017));
  INVX1   g00509(.A(P3_DATAWIDTH_REG_14__SCAN_IN), .Y(n3473));
  NOR2X1  g00510(.A(n3446), .B(n3473), .Y(P3_U3016));
  INVX1   g00511(.A(P3_DATAWIDTH_REG_15__SCAN_IN), .Y(n3475));
  NOR2X1  g00512(.A(n3446), .B(n3475), .Y(P3_U3015));
  INVX1   g00513(.A(P3_DATAWIDTH_REG_16__SCAN_IN), .Y(n3477));
  NOR2X1  g00514(.A(n3446), .B(n3477), .Y(P3_U3014));
  INVX1   g00515(.A(P3_DATAWIDTH_REG_17__SCAN_IN), .Y(n3479));
  NOR2X1  g00516(.A(n3446), .B(n3479), .Y(P3_U3013));
  INVX1   g00517(.A(P3_DATAWIDTH_REG_18__SCAN_IN), .Y(n3481));
  NOR2X1  g00518(.A(n3446), .B(n3481), .Y(P3_U3012));
  INVX1   g00519(.A(P3_DATAWIDTH_REG_19__SCAN_IN), .Y(n3483));
  NOR2X1  g00520(.A(n3446), .B(n3483), .Y(P3_U3011));
  INVX1   g00521(.A(P3_DATAWIDTH_REG_20__SCAN_IN), .Y(n3485));
  NOR2X1  g00522(.A(n3446), .B(n3485), .Y(P3_U3010));
  INVX1   g00523(.A(P3_DATAWIDTH_REG_21__SCAN_IN), .Y(n3487));
  NOR2X1  g00524(.A(n3446), .B(n3487), .Y(P3_U3009));
  INVX1   g00525(.A(P3_DATAWIDTH_REG_22__SCAN_IN), .Y(n3489));
  NOR2X1  g00526(.A(n3446), .B(n3489), .Y(P3_U3008));
  INVX1   g00527(.A(P3_DATAWIDTH_REG_23__SCAN_IN), .Y(n3491));
  NOR2X1  g00528(.A(n3446), .B(n3491), .Y(P3_U3007));
  INVX1   g00529(.A(P3_DATAWIDTH_REG_24__SCAN_IN), .Y(n3493));
  NOR2X1  g00530(.A(n3446), .B(n3493), .Y(P3_U3006));
  INVX1   g00531(.A(P3_DATAWIDTH_REG_25__SCAN_IN), .Y(n3495));
  NOR2X1  g00532(.A(n3446), .B(n3495), .Y(P3_U3005));
  INVX1   g00533(.A(P3_DATAWIDTH_REG_26__SCAN_IN), .Y(n3497));
  NOR2X1  g00534(.A(n3446), .B(n3497), .Y(P3_U3004));
  INVX1   g00535(.A(P3_DATAWIDTH_REG_27__SCAN_IN), .Y(n3499));
  NOR2X1  g00536(.A(n3446), .B(n3499), .Y(P3_U3003));
  INVX1   g00537(.A(P3_DATAWIDTH_REG_28__SCAN_IN), .Y(n3501));
  NOR2X1  g00538(.A(n3446), .B(n3501), .Y(P3_U3002));
  INVX1   g00539(.A(P3_DATAWIDTH_REG_29__SCAN_IN), .Y(n3503));
  NOR2X1  g00540(.A(n3446), .B(n3503), .Y(P3_U3001));
  INVX1   g00541(.A(P3_DATAWIDTH_REG_30__SCAN_IN), .Y(n3505));
  NOR2X1  g00542(.A(n3446), .B(n3505), .Y(P3_U3000));
  INVX1   g00543(.A(P3_DATAWIDTH_REG_31__SCAN_IN), .Y(n3507));
  NOR2X1  g00544(.A(n3446), .B(n3507), .Y(P3_U2999));
  INVX1   g00545(.A(P3_STATE2_REG_3__SCAN_IN), .Y(n3509));
  INVX1   g00546(.A(P3_STATE2_REG_0__SCAN_IN), .Y(n3510));
  INVX1   g00547(.A(P3_STATE2_REG_2__SCAN_IN), .Y(n3511));
  INVX1   g00548(.A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .Y(n3512));
  INVX1   g00549(.A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .Y(n3513));
  NOR2X1  g00550(.A(n3513), .B(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n3514));
  INVX1   g00551(.A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Y(n3515));
  INVX1   g00552(.A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .Y(n3516));
  INVX1   g00553(.A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Y(n3517));
  INVX1   g00554(.A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Y(n3518));
  INVX1   g00555(.A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Y(n3519));
  AOI21X1 g00556(.A0(n3519), .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B0(n3518), .Y(n3520));
  NAND3X1 g00557(.A(n3519), .B(n3518), .C(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n3521));
  AOI21X1 g00558(.A0(n3521), .A1(n3517), .B0(n3520), .Y(n3522));
  AOI21X1 g00559(.A0(n3516), .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B0(n3522), .Y(n3523));
  AOI21X1 g00560(.A0(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A1(n3515), .B0(n3523), .Y(n3524));
  AOI21X1 g00561(.A0(n3513), .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B0(n3524), .Y(n3525));
  NOR2X1  g00562(.A(n3512), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .Y(n3526));
  NOR3X1  g00563(.A(n3526), .B(n3525), .C(n3514), .Y(n3527));
  AOI21X1 g00564(.A0(n3512), .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B0(n3527), .Y(n3528));
  INVX1   g00565(.A(n3528), .Y(n3529));
  NOR2X1  g00566(.A(n3525), .B(n3514), .Y(n3530));
  INVX1   g00567(.A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .Y(n3531));
  XOR2X1  g00568(.A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B(n3531), .Y(n3532));
  XOR2X1  g00569(.A(n3532), .B(n3530), .Y(n3533));
  INVX1   g00570(.A(n3533), .Y(n3534));
  INVX1   g00571(.A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n3535));
  XOR2X1  g00572(.A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n3535), .Y(n3536));
  XOR2X1  g00573(.A(n3536), .B(n3524), .Y(n3537));
  INVX1   g00574(.A(n3537), .Y(n3538));
  XOR2X1  g00575(.A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n3515), .Y(n3539));
  XOR2X1  g00576(.A(n3539), .B(n3522), .Y(n3540));
  INVX1   g00577(.A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n3541));
  NOR2X1  g00578(.A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n3541), .Y(n3542));
  XOR2X1  g00579(.A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n3517), .Y(n3543));
  XOR2X1  g00580(.A(n3543), .B(n3542), .Y(n3544));
  XOR2X1  g00581(.A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n3541), .Y(n3545));
  AOI21X1 g00582(.A0(n3545), .A1(n3544), .B0(n3540), .Y(n3546));
  NOR3X1  g00583(.A(n3546), .B(n3538), .C(n3534), .Y(n3547));
  INVX1   g00584(.A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .Y(n3549));
  NOR4X1  g00585(.A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .D(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n3550));
  INVX1   g00586(.A(n3550), .Y(n3551));
  NOR2X1  g00587(.A(n3551), .B(n3549), .Y(n3552));
  INVX1   g00588(.A(P3_INSTQUEUE_REG_9__2__SCAN_IN), .Y(n3553));
  INVX1   g00589(.A(P3_INSTQUEUE_REG_3__2__SCAN_IN), .Y(n3554));
  NOR4X1  g00590(.A(n3517), .B(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .D(n3541), .Y(n3555));
  NOR4X1  g00591(.A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(n3535), .D(n3541), .Y(n3557));
  OAI22X1 g00592(.A0(n7188), .A1(n3554), .B0(n3553), .B1(n7166), .Y(n3559));
  NOR4X1  g00593(.A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(n3535), .D(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n3560));
  NAND2X1 g00594(.A(n3560), .B(P3_INSTQUEUE_REG_8__2__SCAN_IN), .Y(n3561));
  NOR4X1  g00595(.A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .D(n3541), .Y(n3562));
  NOR4X1  g00596(.A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n3515), .C(n3535), .D(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n3563));
  AOI22X1 g00597(.A0(n3562), .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B0(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3563), .Y(n3564));
  NOR4X1  g00598(.A(n3517), .B(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(n3535), .D(n3541), .Y(n3565));
  NOR4X1  g00599(.A(n3517), .B(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(n3535), .D(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n3566));
  AOI22X1 g00600(.A0(n3565), .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B0(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3566), .Y(n3567));
  NOR4X1  g00601(.A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n3515), .C(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .D(n3541), .Y(n3568));
  NOR4X1  g00602(.A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n3515), .C(n3535), .D(n3541), .Y(n3569));
  AOI22X1 g00603(.A0(n3568), .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B0(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3569), .Y(n3570));
  NOR4X1  g00604(.A(n3517), .B(n3515), .C(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .D(n3541), .Y(n3571));
  NOR4X1  g00605(.A(n3517), .B(n3515), .C(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .D(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n3572));
  AOI22X1 g00606(.A0(n3571), .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B0(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3572), .Y(n3573));
  NOR4X1  g00607(.A(n3517), .B(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .D(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n3574));
  NOR4X1  g00608(.A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n3515), .C(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .D(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n3575));
  AOI22X1 g00609(.A0(n3574), .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B0(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3575), .Y(n3576));
  NOR4X1  g00610(.A(n3517), .B(n3515), .C(n3535), .D(n3541), .Y(n3577));
  NOR4X1  g00611(.A(n3517), .B(n3515), .C(n3535), .D(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n3578));
  AOI22X1 g00612(.A0(n3577), .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B0(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3578), .Y(n3579));
  NAND4X1 g00613(.A(n3576), .B(n3573), .C(n3570), .D(n3579), .Y(n3580));
  INVX1   g00614(.A(n3580), .Y(n3581));
  NAND4X1 g00615(.A(n3567), .B(n3564), .C(n3561), .D(n3581), .Y(n3582));
  NOR3X1  g00616(.A(n3582), .B(n3559), .C(n3552), .Y(n3583));
  INVX1   g00617(.A(n3583), .Y(n3584));
  INVX1   g00618(.A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .Y(n3585));
  NOR2X1  g00619(.A(n3551), .B(n3585), .Y(n3586));
  INVX1   g00620(.A(P3_INSTQUEUE_REG_9__7__SCAN_IN), .Y(n3587));
  INVX1   g00621(.A(P3_INSTQUEUE_REG_3__7__SCAN_IN), .Y(n3588));
  OAI22X1 g00622(.A0(n7188), .A1(n3588), .B0(n3587), .B1(n7166), .Y(n3589));
  NAND2X1 g00623(.A(n3560), .B(P3_INSTQUEUE_REG_8__7__SCAN_IN), .Y(n3590));
  AOI22X1 g00624(.A0(n3562), .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B0(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3563), .Y(n3591));
  AOI22X1 g00625(.A0(n3565), .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B0(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3566), .Y(n3592));
  AOI22X1 g00626(.A0(n3568), .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B0(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3569), .Y(n3593));
  AOI22X1 g00627(.A0(n3571), .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B0(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3572), .Y(n3594));
  AOI22X1 g00628(.A0(n3574), .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B0(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3575), .Y(n3595));
  AOI22X1 g00629(.A0(n3577), .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B0(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3578), .Y(n3596));
  NAND4X1 g00630(.A(n3595), .B(n3594), .C(n3593), .D(n3596), .Y(n3597));
  INVX1   g00631(.A(n3597), .Y(n3598));
  NAND4X1 g00632(.A(n3592), .B(n3591), .C(n3590), .D(n3598), .Y(n3599));
  NOR3X1  g00633(.A(n3599), .B(n3589), .C(n3586), .Y(n3600));
  INVX1   g00634(.A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .Y(n3601));
  NOR2X1  g00635(.A(n3551), .B(n3601), .Y(n3602));
  INVX1   g00636(.A(P3_INSTQUEUE_REG_9__3__SCAN_IN), .Y(n3603));
  INVX1   g00637(.A(P3_INSTQUEUE_REG_3__3__SCAN_IN), .Y(n3604));
  OAI22X1 g00638(.A0(n7188), .A1(n3604), .B0(n3603), .B1(n7166), .Y(n3605));
  NAND2X1 g00639(.A(n3560), .B(P3_INSTQUEUE_REG_8__3__SCAN_IN), .Y(n3606));
  AOI22X1 g00640(.A0(n3562), .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B0(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3563), .Y(n3607));
  AOI22X1 g00641(.A0(n3565), .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B0(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3566), .Y(n3608));
  AOI22X1 g00642(.A0(n3568), .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B0(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3569), .Y(n3609));
  AOI22X1 g00643(.A0(n3571), .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B0(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3572), .Y(n3610));
  AOI22X1 g00644(.A0(n3574), .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B0(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3575), .Y(n3611));
  AOI22X1 g00645(.A0(n3577), .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B0(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3578), .Y(n3612));
  NAND4X1 g00646(.A(n3611), .B(n3610), .C(n3609), .D(n3612), .Y(n3613));
  INVX1   g00647(.A(n3613), .Y(n3614));
  NAND4X1 g00648(.A(n3608), .B(n3607), .C(n3606), .D(n3614), .Y(n3615));
  NOR3X1  g00649(.A(n3615), .B(n3605), .C(n3602), .Y(n3616));
  NOR3X1  g00650(.A(n3616), .B(n3600), .C(n3584), .Y(n3617));
  INVX1   g00651(.A(n3617), .Y(n3618));
  INVX1   g00652(.A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .Y(n3619));
  NOR2X1  g00653(.A(n3551), .B(n3619), .Y(n3620));
  INVX1   g00654(.A(P3_INSTQUEUE_REG_9__4__SCAN_IN), .Y(n3621));
  INVX1   g00655(.A(P3_INSTQUEUE_REG_3__4__SCAN_IN), .Y(n3622));
  OAI22X1 g00656(.A0(n7188), .A1(n3622), .B0(n3621), .B1(n7166), .Y(n3623));
  NAND2X1 g00657(.A(n3560), .B(P3_INSTQUEUE_REG_8__4__SCAN_IN), .Y(n3624));
  AOI22X1 g00658(.A0(n3562), .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B0(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3563), .Y(n3625));
  AOI22X1 g00659(.A0(n3565), .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B0(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3566), .Y(n3626));
  AOI22X1 g00660(.A0(n3568), .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B0(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3569), .Y(n3627));
  AOI22X1 g00661(.A0(n3571), .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B0(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3572), .Y(n3628));
  AOI22X1 g00662(.A0(n3574), .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B0(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3575), .Y(n3629));
  AOI22X1 g00663(.A0(n3577), .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B0(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3578), .Y(n3630));
  NAND4X1 g00664(.A(n3629), .B(n3628), .C(n3627), .D(n3630), .Y(n3631));
  INVX1   g00665(.A(n3631), .Y(n3632));
  NAND4X1 g00666(.A(n3626), .B(n3625), .C(n3624), .D(n3632), .Y(n3633));
  NOR3X1  g00667(.A(n3633), .B(n3623), .C(n3620), .Y(n3634));
  INVX1   g00668(.A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .Y(n3635));
  NOR2X1  g00669(.A(n3551), .B(n3635), .Y(n3636));
  INVX1   g00670(.A(P3_INSTQUEUE_REG_9__5__SCAN_IN), .Y(n3637));
  INVX1   g00671(.A(P3_INSTQUEUE_REG_3__5__SCAN_IN), .Y(n3638));
  OAI22X1 g00672(.A0(n7188), .A1(n3638), .B0(n3637), .B1(n7166), .Y(n3639));
  NAND2X1 g00673(.A(n3560), .B(P3_INSTQUEUE_REG_8__5__SCAN_IN), .Y(n3640));
  AOI22X1 g00674(.A0(n3562), .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B0(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3563), .Y(n3641));
  AOI22X1 g00675(.A0(n3565), .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B0(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3566), .Y(n3642));
  AOI22X1 g00676(.A0(n3568), .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B0(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3569), .Y(n3643));
  AOI22X1 g00677(.A0(n3571), .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B0(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3572), .Y(n3644));
  AOI22X1 g00678(.A0(n3574), .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B0(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3575), .Y(n3645));
  AOI22X1 g00679(.A0(n3577), .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B0(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3578), .Y(n3646));
  NAND4X1 g00680(.A(n3645), .B(n3644), .C(n3643), .D(n3646), .Y(n3647));
  INVX1   g00681(.A(n3647), .Y(n3648));
  NAND4X1 g00682(.A(n3642), .B(n3641), .C(n3640), .D(n3648), .Y(n3649));
  NOR3X1  g00683(.A(n3649), .B(n3639), .C(n3636), .Y(n3650));
  INVX1   g00684(.A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .Y(n3651));
  NOR2X1  g00685(.A(n3551), .B(n3651), .Y(n3652));
  INVX1   g00686(.A(P3_INSTQUEUE_REG_9__6__SCAN_IN), .Y(n3653));
  INVX1   g00687(.A(P3_INSTQUEUE_REG_3__6__SCAN_IN), .Y(n3654));
  OAI22X1 g00688(.A0(n7188), .A1(n3654), .B0(n3653), .B1(n7166), .Y(n3655));
  NAND2X1 g00689(.A(n3560), .B(P3_INSTQUEUE_REG_8__6__SCAN_IN), .Y(n3656));
  AOI22X1 g00690(.A0(n3562), .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B0(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3563), .Y(n3657));
  AOI22X1 g00691(.A0(n3565), .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B0(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3566), .Y(n3658));
  AOI22X1 g00692(.A0(n3568), .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B0(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3569), .Y(n3659));
  AOI22X1 g00693(.A0(n3571), .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B0(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3572), .Y(n3660));
  AOI22X1 g00694(.A0(n3574), .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B0(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3575), .Y(n3661));
  AOI22X1 g00695(.A0(n3577), .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B0(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3578), .Y(n3662));
  NAND4X1 g00696(.A(n3661), .B(n3660), .C(n3659), .D(n3662), .Y(n3663));
  INVX1   g00697(.A(n3663), .Y(n3664));
  NAND4X1 g00698(.A(n3658), .B(n3657), .C(n3656), .D(n3664), .Y(n3665));
  NOR4X1  g00699(.A(n3655), .B(n3652), .C(n3650), .D(n3665), .Y(n3666));
  INVX1   g00700(.A(n3666), .Y(n3667));
  INVX1   g00701(.A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .Y(n3668));
  AOI22X1 g00702(.A0(n3555), .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B0(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3557), .Y(n3669));
  OAI21X1 g00703(.A0(n3551), .A1(n3668), .B0(n3669), .Y(n3670));
  NAND2X1 g00704(.A(n3560), .B(P3_INSTQUEUE_REG_8__1__SCAN_IN), .Y(n3671));
  AOI22X1 g00705(.A0(n3562), .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B0(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3563), .Y(n3672));
  AOI22X1 g00706(.A0(n3565), .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B0(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3566), .Y(n3673));
  AOI22X1 g00707(.A0(n3568), .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B0(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3569), .Y(n3674));
  AOI22X1 g00708(.A0(n3571), .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B0(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3572), .Y(n3675));
  AOI22X1 g00709(.A0(n3574), .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B0(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3575), .Y(n3676));
  AOI22X1 g00710(.A0(n3577), .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B0(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3578), .Y(n3677));
  NAND4X1 g00711(.A(n3676), .B(n3675), .C(n3674), .D(n3677), .Y(n3678));
  INVX1   g00712(.A(n3678), .Y(n3679));
  NAND4X1 g00713(.A(n3673), .B(n3672), .C(n3671), .D(n3679), .Y(n3680));
  NOR2X1  g00714(.A(n3680), .B(n3670), .Y(n3681));
  INVX1   g00715(.A(n3681), .Y(n3682));
  INVX1   g00716(.A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .Y(n3683));
  NOR2X1  g00717(.A(n3551), .B(n3683), .Y(n3684));
  INVX1   g00718(.A(P3_INSTQUEUE_REG_9__0__SCAN_IN), .Y(n3685));
  INVX1   g00719(.A(P3_INSTQUEUE_REG_3__0__SCAN_IN), .Y(n3686));
  OAI22X1 g00720(.A0(n7188), .A1(n3686), .B0(n3685), .B1(n7166), .Y(n3687));
  NAND2X1 g00721(.A(n3560), .B(P3_INSTQUEUE_REG_8__0__SCAN_IN), .Y(n3688));
  AOI22X1 g00722(.A0(n3562), .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B0(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3563), .Y(n3689));
  AOI22X1 g00723(.A0(n3565), .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B0(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3566), .Y(n3690));
  AOI22X1 g00724(.A0(n3568), .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B0(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3569), .Y(n3691));
  AOI22X1 g00725(.A0(n3571), .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B0(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3572), .Y(n3692));
  AOI22X1 g00726(.A0(n3574), .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B0(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3575), .Y(n3693));
  AOI22X1 g00727(.A0(n3577), .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B0(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3578), .Y(n3694));
  NAND4X1 g00728(.A(n3693), .B(n3692), .C(n3691), .D(n3694), .Y(n3695));
  INVX1   g00729(.A(n3695), .Y(n3696));
  NAND4X1 g00730(.A(n3690), .B(n3689), .C(n3688), .D(n3696), .Y(n3697));
  NOR3X1  g00731(.A(n3697), .B(n3687), .C(n3684), .Y(n3698));
  INVX1   g00732(.A(n3698), .Y(n3699));
  NOR2X1  g00733(.A(n3699), .B(n3682), .Y(n3700));
  INVX1   g00734(.A(n3700), .Y(n3701));
  NOR4X1  g00735(.A(n3667), .B(n3634), .C(n3618), .D(n3701), .Y(n3702));
  NAND2X1 g00736(.A(n3544), .B(n3540), .Y(n3703));
  NOR3X1  g00737(.A(n3703), .B(n3538), .C(n3534), .Y(n3704));
  NOR2X1  g00738(.A(n3704), .B(n3529), .Y(n3705));
  INVX1   g00739(.A(n3616), .Y(n3706));
  INVX1   g00740(.A(n3634), .Y(n3707));
  NOR3X1  g00741(.A(n3665), .B(n3655), .C(n3652), .Y(n3708));
  NOR2X1  g00742(.A(n3708), .B(n3650), .Y(n3709));
  INVX1   g00743(.A(n3709), .Y(n3710));
  NOR4X1  g00744(.A(n3707), .B(n3706), .C(n3600), .D(n3710), .Y(n3711));
  INVX1   g00745(.A(n3711), .Y(n3712));
  NOR3X1  g00746(.A(n3712), .B(n3701), .C(n3583), .Y(n3713));
  INVX1   g00747(.A(n3650), .Y(n3714));
  INVX1   g00748(.A(n3708), .Y(n3715));
  NOR3X1  g00749(.A(n3715), .B(n3714), .C(n3707), .Y(n3716));
  INVX1   g00750(.A(n3716), .Y(n3717));
  NOR2X1  g00751(.A(n3698), .B(n3681), .Y(n3718));
  INVX1   g00752(.A(n3718), .Y(n3719));
  NOR3X1  g00753(.A(n3719), .B(n3717), .C(n3618), .Y(n3720));
  OAI21X1 g00754(.A0(n3720), .A1(n3713), .B0(n3705), .Y(n3721));
  NOR2X1  g00755(.A(n3721), .B(n3407), .Y(n3722));
  AOI21X1 g00756(.A0(n3702), .A1(n3893), .B0(n3722), .Y(n3723));
  XOR2X1  g00757(.A(P3_STATE_REG_1__SCAN_IN), .B(n3402), .Y(n3724));
  NOR2X1  g00758(.A(n3724), .B(P3_STATE_REG_0__SCAN_IN), .Y(n3725));
  INVX1   g00759(.A(n3725), .Y(n3726));
  NOR4X1  g00760(.A(n3687), .B(n3684), .C(n3681), .D(n3697), .Y(n3727));
  INVX1   g00761(.A(n3727), .Y(n3728));
  NOR3X1  g00762(.A(n3728), .B(n3712), .C(n3583), .Y(n3729));
  NOR3X1  g00763(.A(n3698), .B(n3680), .C(n3670), .Y(n3730));
  INVX1   g00764(.A(n3730), .Y(n3731));
  NOR3X1  g00765(.A(n3731), .B(n3717), .C(n3618), .Y(n3732));
  OAI21X1 g00766(.A0(n3732), .A1(n3729), .B0(n3705), .Y(n3733));
  NOR3X1  g00767(.A(n3733), .B(n3726), .C(n3407), .Y(n3734));
  AOI21X1 g00768(.A0(n3698), .A1(n3634), .B0(n3616), .Y(n3735));
  OAI21X1 g00769(.A0(n3699), .A1(n3681), .B0(n3735), .Y(n3736));
  NOR4X1  g00770(.A(n3649), .B(n3639), .C(n3636), .D(n3708), .Y(n3737));
  NOR4X1  g00771(.A(n3715), .B(n3650), .C(n3707), .D(n3681), .Y(n3738));
  NOR4X1  g00772(.A(n3737), .B(n3736), .C(n3600), .D(n3738), .Y(n3739));
  NOR3X1  g00773(.A(n3737), .B(n3666), .C(n3600), .Y(n3740));
  NOR2X1  g00774(.A(n3740), .B(n3731), .Y(n3741));
  AOI21X1 g00775(.A0(n3711), .A1(n3698), .B0(n3583), .Y(n3742));
  NOR2X1  g00776(.A(n3742), .B(n3741), .Y(n3743));
  OAI21X1 g00777(.A0(n3739), .A1(n3584), .B0(n3743), .Y(n3744));
  NOR4X1  g00778(.A(n3667), .B(n3634), .C(n3618), .D(n3719), .Y(n3745));
  NAND2X1 g00779(.A(n3745), .B(n3893), .Y(n3746));
  NOR4X1  g00780(.A(n3582), .B(n3559), .C(n3552), .D(n3634), .Y(n3747));
  INVX1   g00781(.A(n3747), .Y(n3748));
  OAI21X1 g00782(.A0(n3748), .A1(n3666), .B0(n3746), .Y(n3749));
  NOR3X1  g00783(.A(n3749), .B(n3744), .C(n3734), .Y(n3750));
  NAND2X1 g00784(.A(n3750), .B(n3723), .Y(n3751));
  INVX1   g00785(.A(n3751), .Y(n3752));
  INVX1   g00786(.A(n3713), .Y(n3753));
  NAND3X1 g00787(.A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n3754));
  XOR2X1  g00788(.A(n3754), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .Y(n3755));
  NOR3X1  g00789(.A(n3755), .B(n3752), .C(n3753), .Y(n3756));
  AOI21X1 g00790(.A0(n3752), .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B0(n3756), .Y(n3757));
  NOR3X1  g00791(.A(n3717), .B(n3698), .C(n3618), .Y(n3758));
  NOR4X1  g00792(.A(n3714), .B(n3706), .C(n3584), .D(n3708), .Y(n3759));
  NAND2X1 g00793(.A(n3759), .B(n3700), .Y(n3760));
  NOR2X1  g00794(.A(n3760), .B(n3600), .Y(n3761));
  NOR3X1  g00795(.A(n3761), .B(n3758), .C(n3729), .Y(n3762));
  INVX1   g00796(.A(n3762), .Y(n3763));
  AOI21X1 g00797(.A0(n3740), .A1(n3706), .B0(n3731), .Y(n3764));
  INVX1   g00798(.A(n3764), .Y(n3765));
  NOR2X1  g00799(.A(n3616), .B(n3600), .Y(n3766));
  INVX1   g00800(.A(n3766), .Y(n3767));
  AOI21X1 g00801(.A0(n3650), .A1(n3600), .B0(n3681), .Y(n3768));
  NOR2X1  g00802(.A(n3715), .B(n3707), .Y(n3769));
  AOI22X1 g00803(.A0(n3709), .A1(n3700), .B0(n3698), .B1(n3769), .Y(n3770));
  INVX1   g00804(.A(n3770), .Y(n3771));
  AOI21X1 g00805(.A0(n3768), .A1(n3767), .B0(n3771), .Y(n3772));
  AOI21X1 g00806(.A0(n3772), .A1(n3765), .B0(n3584), .Y(n3773));
  INVX1   g00807(.A(n3600), .Y(n3774));
  OAI21X1 g00808(.A0(n3682), .A1(n3774), .B0(n3698), .Y(n3775));
  NAND3X1 g00809(.A(n3775), .B(n3714), .C(n3616), .Y(n3776));
  NAND3X1 g00810(.A(n3682), .B(n3708), .C(n3600), .Y(n3777));
  OAI21X1 g00811(.A0(n3728), .A1(n3709), .B0(n3777), .Y(n3778));
  NOR3X1  g00812(.A(n3769), .B(n3714), .C(n3616), .Y(n3779));
  NOR3X1  g00813(.A(n3779), .B(n3778), .C(n3738), .Y(n3780));
  NAND2X1 g00814(.A(n3780), .B(n3776), .Y(n3781));
  NOR3X1  g00815(.A(n3730), .B(n3709), .C(n3600), .Y(n3782));
  NOR4X1  g00816(.A(n3655), .B(n3652), .C(n3600), .D(n3665), .Y(n3783));
  NOR3X1  g00817(.A(n3783), .B(n3737), .C(n3706), .Y(n3784));
  OAI22X1 g00818(.A0(n3782), .A1(n3634), .B0(n3583), .B1(n3784), .Y(n3785));
  NOR3X1  g00819(.A(n3785), .B(n3781), .C(n3773), .Y(n3786));
  INVX1   g00820(.A(n3786), .Y(n3787));
  NOR2X1  g00821(.A(n3715), .B(n3706), .Y(n3788));
  INVX1   g00822(.A(n3788), .Y(n3789));
  NOR4X1  g00823(.A(n3699), .B(n3682), .C(n3600), .D(n3748), .Y(n3790));
  INVX1   g00824(.A(n3790), .Y(n3791));
  NOR4X1  g00825(.A(n3707), .B(n3774), .C(n3583), .D(n3714), .Y(n3792));
  INVX1   g00826(.A(n3792), .Y(n3793));
  AOI21X1 g00827(.A0(n3793), .A1(n3791), .B0(n3789), .Y(n3794));
  NOR3X1  g00828(.A(n3708), .B(n3650), .C(n3707), .Y(n3795));
  NOR3X1  g00829(.A(n3706), .B(n3774), .C(n3583), .Y(n3796));
  NAND3X1 g00830(.A(n3796), .B(n3727), .C(n3795), .Y(n3797));
  INVX1   g00831(.A(n3797), .Y(n3798));
  NOR4X1  g00832(.A(n3707), .B(n3767), .C(n3584), .D(n3710), .Y(n3799));
  AOI21X1 g00833(.A0(n3799), .A1(n3682), .B0(n3798), .Y(n3800));
  INVX1   g00834(.A(n3800), .Y(n3801));
  INVX1   g00835(.A(n3759), .Y(n3802));
  NOR2X1  g00836(.A(n3707), .B(n3774), .Y(n3803));
  INVX1   g00837(.A(n3803), .Y(n3804));
  NOR3X1  g00838(.A(n3804), .B(n3802), .C(n3719), .Y(n3805));
  NOR4X1  g00839(.A(n3801), .B(n3794), .C(n3787), .D(n3805), .Y(n3806));
  NAND2X1 g00840(.A(n3806), .B(n3760), .Y(n3807));
  AOI21X1 g00841(.A0(n3807), .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B0(n3763), .Y(n3808));
  NOR3X1  g00842(.A(n3808), .B(n3517), .C(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Y(n3809));
  AOI21X1 g00843(.A0(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B0(n3515), .Y(n3810));
  NOR3X1  g00844(.A(n3682), .B(n3715), .C(n3706), .Y(n3811));
  OAI21X1 g00845(.A0(n3792), .A1(n3747), .B0(n3811), .Y(n3812));
  XOR2X1  g00846(.A(n3698), .B(n3681), .Y(n3813));
  NAND2X1 g00847(.A(n3803), .B(n3759), .Y(n3814));
  OAI21X1 g00848(.A0(n3814), .A1(n3813), .B0(n3812), .Y(n3815));
  NOR2X1  g00849(.A(n3815), .B(n3801), .Y(n3816));
  INVX1   g00850(.A(n3816), .Y(n3817));
  OAI21X1 g00851(.A0(n3817), .A1(n3787), .B0(n3810), .Y(n3818));
  NOR2X1  g00852(.A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n3515), .Y(n3819));
  NAND2X1 g00853(.A(n3819), .B(n3763), .Y(n3820));
  NOR2X1  g00854(.A(n3517), .B(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Y(n3821));
  OAI21X1 g00855(.A0(n3819), .A1(n3821), .B0(n3713), .Y(n3822));
  NOR2X1  g00856(.A(n3541), .B(n3517), .Y(n3823));
  XOR2X1  g00857(.A(n3823), .B(n3515), .Y(n3824));
  INVX1   g00858(.A(n3824), .Y(n3825));
  NOR2X1  g00859(.A(n3825), .B(n3813), .Y(n3826));
  NAND4X1 g00860(.A(n3666), .B(n3707), .C(n3617), .D(n3826), .Y(n3827));
  NAND4X1 g00861(.A(n3822), .B(n3820), .C(n3818), .D(n3827), .Y(n3828));
  NOR2X1  g00862(.A(n3828), .B(n3809), .Y(n3829));
  INVX1   g00863(.A(n3829), .Y(n3830));
  NOR2X1  g00864(.A(n3751), .B(n3515), .Y(n3831));
  AOI21X1 g00865(.A0(n3830), .A1(n3751), .B0(n3831), .Y(n3832));
  NOR2X1  g00866(.A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(n3517), .Y(n3833));
  NOR2X1  g00867(.A(n3804), .B(n3760), .Y(n3834));
  INVX1   g00868(.A(n3834), .Y(n3835));
  NAND2X1 g00869(.A(n3835), .B(n3806), .Y(n3836));
  NOR4X1  g00870(.A(n3634), .B(n3767), .C(n3584), .D(n3667), .Y(n3837));
  AOI22X1 g00871(.A0(n3718), .A1(n3837), .B0(n3666), .B1(n3790), .Y(n3838));
  XOR2X1  g00872(.A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(n3517), .Y(n3839));
  OAI22X1 g00873(.A0(n3838), .A1(n3839), .B0(n3753), .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Y(n3840));
  AOI21X1 g00874(.A0(n3836), .A1(n3833), .B0(n3840), .Y(n3841));
  OAI21X1 g00875(.A0(n3808), .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B0(n3841), .Y(n3842));
  NOR2X1  g00876(.A(n3751), .B(n3517), .Y(n3843));
  AOI21X1 g00877(.A0(n3842), .A1(n3751), .B0(n3843), .Y(n3844));
  NAND3X1 g00878(.A(n3838), .B(n3835), .C(n3806), .Y(n3845));
  NAND2X1 g00879(.A(n3845), .B(n3541), .Y(n3846));
  OAI21X1 g00880(.A0(n3763), .A1(n3713), .B0(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n3847));
  NAND2X1 g00881(.A(n3847), .B(n3846), .Y(n3848));
  OAI21X1 g00882(.A0(n3751), .A1(n3541), .B0(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Y(n3849));
  AOI21X1 g00883(.A0(n3848), .A1(n3751), .B0(n3849), .Y(n3850));
  AOI21X1 g00884(.A0(n3850), .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B0(n3844), .Y(n3851));
  NOR2X1  g00885(.A(n3850), .B(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Y(n3852));
  NOR2X1  g00886(.A(n3852), .B(n3851), .Y(n3853));
  OAI21X1 g00887(.A0(n3832), .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B0(n3853), .Y(n3854));
  NOR4X1  g00888(.A(n3517), .B(n3515), .C(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .D(n3808), .Y(n3855));
  NAND2X1 g00889(.A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Y(n3856));
  NOR3X1  g00890(.A(n3732), .B(n3729), .C(n3720), .Y(n3857));
  NOR3X1  g00891(.A(n3760), .B(n3634), .C(n3600), .Y(n3858));
  INVX1   g00892(.A(n3858), .Y(n3859));
  NOR3X1  g00893(.A(n3760), .B(n3707), .C(n3600), .Y(n3860));
  INVX1   g00894(.A(n3860), .Y(n3861));
  NAND4X1 g00895(.A(n3859), .B(n3857), .C(n3786), .D(n3861), .Y(n3862));
  NAND3X1 g00896(.A(n3862), .B(n3856), .C(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n3863));
  NOR3X1  g00897(.A(n3786), .B(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C(n3535), .Y(n3864));
  INVX1   g00898(.A(n3864), .Y(n3865));
  NOR3X1  g00899(.A(n3541), .B(n3517), .C(n3515), .Y(n3866));
  NOR2X1  g00900(.A(n3866), .B(n3535), .Y(n3867));
  NAND2X1 g00901(.A(n3515), .B(n3535), .Y(n3868));
  OAI21X1 g00902(.A0(n3823), .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B0(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n3869));
  OAI21X1 g00903(.A0(n3868), .A1(n3823), .B0(n3869), .Y(n3870));
  NOR2X1  g00904(.A(n3870), .B(n3813), .Y(n3871));
  XOR2X1  g00905(.A(n3856), .B(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n3872));
  NOR4X1  g00906(.A(n3712), .B(n3701), .C(n3583), .D(n3872), .Y(n3873));
  AOI21X1 g00907(.A0(n3871), .A1(n3837), .B0(n3873), .Y(n3874));
  INVX1   g00908(.A(n3874), .Y(n3875));
  AOI21X1 g00909(.A0(n3867), .A1(n3817), .B0(n3875), .Y(n3876));
  NAND3X1 g00910(.A(n3876), .B(n3865), .C(n3863), .Y(n3877));
  NOR2X1  g00911(.A(n3877), .B(n3855), .Y(n3878));
  INVX1   g00912(.A(n3878), .Y(n3879));
  NOR2X1  g00913(.A(n3751), .B(n3535), .Y(n3880));
  AOI21X1 g00914(.A0(n3879), .A1(n3751), .B0(n3880), .Y(n3881));
  AOI22X1 g00915(.A0(n3832), .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B0(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B1(n3881), .Y(n3882));
  OAI22X1 g00916(.A0(n3881), .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B0(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B1(n3757), .Y(n3883));
  AOI21X1 g00917(.A0(n3882), .A1(n3854), .B0(n3883), .Y(n3884));
  AOI21X1 g00918(.A0(n3757), .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B0(n3884), .Y(n3885));
  NOR2X1  g00919(.A(n3751), .B(n3531), .Y(n3886));
  NOR2X1  g00920(.A(n3538), .B(n3534), .Y(n3887));
  OAI21X1 g00921(.A0(n3545), .A1(n3544), .B0(n3540), .Y(n3888));
  INVX1   g00922(.A(n3888), .Y(n3889));
  AOI21X1 g00923(.A0(n3889), .A1(n3887), .B0(n3529), .Y(n3890));
  INVX1   g00924(.A(n3890), .Y(n3891));
  NOR2X1  g00925(.A(n3546), .B(n3538), .Y(n3892));
  AOI21X1 g00926(.A0(n3892), .A1(n3533), .B0(n3529), .Y(n3893));
  INVX1   g00927(.A(n3795), .Y(n3894));
  NOR3X1  g00928(.A(n3894), .B(n3698), .C(n3618), .Y(n3895));
  OAI21X1 g00929(.A0(n3893), .A1(n3682), .B0(n3895), .Y(n3896));
  AOI21X1 g00930(.A0(n3891), .A1(n3682), .B0(n3896), .Y(n3897));
  NOR2X1  g00931(.A(n3705), .B(n3682), .Y(n3898));
  OAI21X1 g00932(.A0(n3704), .A1(n3529), .B0(n3682), .Y(n3899));
  NAND3X1 g00933(.A(n3899), .B(n3711), .C(n3698), .Y(n3900));
  NOR2X1  g00934(.A(n3900), .B(n3898), .Y(n3901));
  NOR2X1  g00935(.A(n3901), .B(n3583), .Y(n3902));
  NOR4X1  g00936(.A(n3717), .B(n3698), .C(n3767), .D(n3898), .Y(n3903));
  AOI21X1 g00937(.A0(n3903), .A1(n3899), .B0(n3584), .Y(n3904));
  NOR4X1  g00938(.A(n3670), .B(n3583), .C(n3407), .D(n3680), .Y(n3905));
  NOR3X1  g00939(.A(n3724), .B(n3407), .C(P3_STATE_REG_0__SCAN_IN), .Y(n3906));
  NOR4X1  g00940(.A(n3559), .B(n3552), .C(n3407), .D(n3582), .Y(n3907));
  OAI21X1 g00941(.A0(n3906), .A1(n3682), .B0(n3907), .Y(n3908));
  NOR4X1  g00942(.A(n3681), .B(n3583), .C(n3407), .D(n3726), .Y(n3909));
  INVX1   g00943(.A(n3909), .Y(n3910));
  NAND2X1 g00944(.A(n3910), .B(n3908), .Y(n3911));
  NOR4X1  g00945(.A(n3905), .B(n3904), .C(n3902), .D(n3911), .Y(n3912));
  OAI21X1 g00946(.A0(P3_MORE_REG_SCAN_IN), .A1(P3_FLUSH_REG_SCAN_IN), .B0(n3912), .Y(n3913));
  NOR3X1  g00947(.A(n3719), .B(n3894), .C(n3618), .Y(n3914));
  NAND2X1 g00948(.A(n3914), .B(n3891), .Y(n3915));
  OAI21X1 g00949(.A0(n3753), .A1(n3705), .B0(n3915), .Y(n3916));
  INVX1   g00950(.A(n3729), .Y(n3917));
  INVX1   g00951(.A(n3732), .Y(n3918));
  AOI21X1 g00952(.A0(n3918), .A1(n3917), .B0(n3705), .Y(n3919));
  INVX1   g00953(.A(n3720), .Y(n3920));
  NOR3X1  g00954(.A(n3731), .B(n3894), .C(n3618), .Y(n3921));
  INVX1   g00955(.A(n3921), .Y(n3922));
  OAI22X1 g00956(.A0(n3893), .A1(n3922), .B0(n3920), .B1(n3705), .Y(n3923));
  INVX1   g00957(.A(n3702), .Y(n3924));
  INVX1   g00958(.A(n3745), .Y(n3925));
  AOI21X1 g00959(.A0(n3925), .A1(n3924), .B0(n3893), .Y(n3926));
  NOR4X1  g00960(.A(n3923), .B(n3919), .C(n3916), .D(n3926), .Y(n3927));
  OAI21X1 g00961(.A0(n3927), .A1(n3912), .B0(n3913), .Y(n3928));
  NOR4X1  g00962(.A(n3897), .B(n3756), .C(n3886), .D(n3928), .Y(n3929));
  OAI21X1 g00963(.A0(n3881), .A1(n3832), .B0(n3929), .Y(n3930));
  AOI21X1 g00964(.A0(READY22_REG_SCAN_IN), .A1(READY2), .B0(P3_STATEBS16_REG_SCAN_IN), .Y(n3931));
  INVX1   g00965(.A(n3931), .Y(n3932));
  NOR3X1  g00966(.A(n3932), .B(n3918), .C(n3726), .Y(n3933));
  NOR4X1  g00967(.A(n3930), .B(n3885), .C(P3_STATE2_REG_1__SCAN_IN), .D(n3933), .Y(n3934));
  NOR2X1  g00968(.A(n3934), .B(n3510), .Y(n3935));
  AOI21X1 g00969(.A0(n3407), .A1(P3_STATE2_REG_1__SCAN_IN), .B0(P3_STATE2_REG_0__SCAN_IN), .Y(n3936));
  NOR3X1  g00970(.A(n3936), .B(n3935), .C(n3511), .Y(n3937));
  NOR2X1  g00971(.A(n3937), .B(n3510), .Y(n3938));
  INVX1   g00972(.A(P3_STATE2_REG_1__SCAN_IN), .Y(n3939));
  NOR2X1  g00973(.A(n3939), .B(n3511), .Y(n3940));
  NAND2X1 g00974(.A(n3938), .B(n3940), .Y(n3941));
  OAI21X1 g00975(.A0(n3938), .A1(n3509), .B0(n3941), .Y(P3_U3282));
  OAI21X1 g00976(.A0(n3407), .A1(P3_STATE2_REG_2__SCAN_IN), .B0(P3_STATE2_REG_0__SCAN_IN), .Y(n3943));
  INVX1   g00977(.A(P3_STATEBS16_REG_SCAN_IN), .Y(n3944));
  AOI21X1 g00978(.A0(n3944), .A1(n3510), .B0(n3939), .Y(n3945));
  NOR2X1  g00979(.A(P3_STATE2_REG_1__SCAN_IN), .B(n3511), .Y(n3946));
  AOI21X1 g00980(.A0(n3945), .A1(n3943), .B0(n3946), .Y(n3947));
  OAI21X1 g00981(.A0(n3938), .A1(n3511), .B0(n3947), .Y(P3_U2998));
  NOR2X1  g00982(.A(P3_STATE2_REG_1__SCAN_IN), .B(P3_STATE2_REG_3__SCAN_IN), .Y(n3949));
  NAND3X1 g00983(.A(n3949), .B(n3938), .C(n3408), .Y(n3950));
  NOR4X1  g00984(.A(P3_STATE2_REG_2__SCAN_IN), .B(n3404), .C(n3403), .D(n3510), .Y(n3951));
  OAI21X1 g00985(.A0(n3951), .A1(n3937), .B0(P3_STATE2_REG_1__SCAN_IN), .Y(n3952));
  INVX1   g00986(.A(n3937), .Y(n3953));
  NOR4X1  g00987(.A(P3_STATE2_REG_0__SCAN_IN), .B(n3939), .C(P3_STATE2_REG_2__SCAN_IN), .D(P3_STATEBS16_REG_SCAN_IN), .Y(n3954));
  NOR3X1  g00988(.A(n3510), .B(P3_STATE2_REG_1__SCAN_IN), .C(n3511), .Y(n3955));
  AOI21X1 g00989(.A0(n3955), .A1(n3953), .B0(n3954), .Y(n3956));
  NAND3X1 g00990(.A(n3956), .B(n3952), .C(n3950), .Y(P3_U2997));
  INVX1   g00991(.A(n3940), .Y(n3958));
  INVX1   g00992(.A(P3_FLUSH_REG_SCAN_IN), .Y(n3959));
  INVX1   g00993(.A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .Y(n3960));
  INVX1   g00994(.A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .Y(n3961));
  NOR2X1  g00995(.A(n3961), .B(n3960), .Y(n3962));
  NOR2X1  g00996(.A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n3960), .Y(n3963));
  XOR2X1  g00997(.A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n3960), .Y(n3965));
  NOR2X1  g00998(.A(n3965), .B(n3961), .Y(n3966));
  INVX1   g00999(.A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .Y(n3967));
  NOR2X1  g01000(.A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n3967), .Y(n3968));
  NOR4X1  g01001(.A(n3966), .B(n3960), .C(n3959), .D(n3968), .Y(n3969));
  NOR3X1  g01002(.A(n3963), .B(n3962), .C(n3959), .Y(n3970));
  AOI21X1 g01003(.A0(n3541), .A1(n3517), .B0(P3_FLUSH_REG_SCAN_IN), .Y(n3971));
  NOR3X1  g01004(.A(n3971), .B(n3970), .C(n3969), .Y(n3972));
  INVX1   g01005(.A(n3965), .Y(n3973));
  AOI21X1 g01006(.A0(n3973), .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B0(n3968), .Y(n3974));
  NAND3X1 g01007(.A(n3959), .B(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n3975));
  OAI22X1 g01008(.A0(n3972), .A1(n3975), .B0(P3_FLUSH_REG_SCAN_IN), .B1(n3531), .Y(n3976));
  NOR2X1  g01009(.A(n3976), .B(n3958), .Y(n3977));
  OAI21X1 g01010(.A0(n3977), .A1(n3937), .B0(P3_STATE2_REG_0__SCAN_IN), .Y(n3978));
  NOR2X1  g01011(.A(P3_STATE2_REG_1__SCAN_IN), .B(P3_STATE2_REG_2__SCAN_IN), .Y(n3979));
  NOR2X1  g01012(.A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n3509), .Y(n3980));
  AOI21X1 g01013(.A0(n3980), .A1(n3979), .B0(P3_STATE2_REG_0__SCAN_IN), .Y(n3981));
  NAND2X1 g01014(.A(n3981), .B(n3953), .Y(n3982));
  OAI21X1 g01015(.A0(n3930), .A1(n3885), .B0(n3955), .Y(n3983));
  NOR4X1  g01016(.A(P3_STATE2_REG_1__SCAN_IN), .B(P3_STATE2_REG_2__SCAN_IN), .C(n3509), .D(n3510), .Y(n3984));
  NOR2X1  g01017(.A(n3984), .B(n3951), .Y(n3985));
  NAND4X1 g01018(.A(n3983), .B(n3982), .C(n3978), .D(n3985), .Y(P3_U2996));
  NAND3X1 g01019(.A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .Y(n3987));
  AOI21X1 g01020(.A0(n3944), .A1(n3509), .B0(P3_STATE2_REG_2__SCAN_IN), .Y(n3988));
  INVX1   g01021(.A(n3988), .Y(n3989));
  NAND3X1 g01022(.A(n3518), .B(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .Y(n3990));
  OAI21X1 g01023(.A0(n3990), .A1(n3989), .B0(n3987), .Y(n3991));
  INVX1   g01024(.A(n3946), .Y(n3992));
  AOI22X1 g01025(.A0(P3_STATE2_REG_1__SCAN_IN), .A1(n3511), .B0(P3_STATE2_REG_3__SCAN_IN), .B1(n3531), .Y(n3993));
  AOI21X1 g01026(.A0(n3993), .A1(n3992), .B0(P3_STATE2_REG_0__SCAN_IN), .Y(n3994));
  NAND3X1 g01027(.A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .Y(n3995));
  OAI21X1 g01028(.A0(n3995), .A1(n3513), .B0(P3_STATE2_REG_3__SCAN_IN), .Y(n3996));
  NAND3X1 g01029(.A(n3996), .B(n3994), .C(n3991), .Y(n3997));
  NAND2X1 g01030(.A(n3997), .B(P3_INSTQUEUE_REG_15__7__SCAN_IN), .Y(n3998));
  NOR3X1  g01031(.A(n3944), .B(P3_STATE2_REG_2__SCAN_IN), .C(P3_STATE2_REG_3__SCAN_IN), .Y(n3999));
  NAND2X1 g01032(.A(n3999), .B(n3990), .Y(n4000));
  AOI21X1 g01033(.A0(n4000), .A1(n3988), .B0(n3987), .Y(n4001));
  NAND3X1 g01034(.A(n4001), .B(n3994), .C(BUF2_REG_7__SCAN_IN), .Y(n4002));
  NOR4X1  g01035(.A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n3516), .C(n3513), .D(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Y(n4003));
  NAND4X1 g01036(.A(n3994), .B(n4003), .C(BUF2_REG_31__SCAN_IN), .D(n3999), .Y(n4004));
  NOR2X1  g01037(.A(n3995), .B(n3513), .Y(n4005));
  NOR4X1  g01038(.A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n3516), .C(n3513), .D(n3519), .Y(n4006));
  INVX1   g01039(.A(n3994), .Y(n4007));
  INVX1   g01040(.A(n3999), .Y(n4008));
  NOR3X1  g01041(.A(n4008), .B(n4007), .C(n3260), .Y(n4009));
  NOR3X1  g01042(.A(n4007), .B(n3600), .C(n3509), .Y(n4010));
  AOI22X1 g01043(.A0(n4009), .A1(n4006), .B0(n4005), .B1(n4010), .Y(n4011));
  NAND4X1 g01044(.A(n4004), .B(n4002), .C(n3998), .D(n4011), .Y(P3_U2995));
  NAND2X1 g01045(.A(n3997), .B(P3_INSTQUEUE_REG_15__6__SCAN_IN), .Y(n4013));
  NAND3X1 g01046(.A(n4001), .B(n3994), .C(BUF2_REG_6__SCAN_IN), .Y(n4014));
  NAND4X1 g01047(.A(n3994), .B(n4003), .C(BUF2_REG_30__SCAN_IN), .D(n3999), .Y(n4015));
  NOR3X1  g01048(.A(n4008), .B(n4007), .C(n3257), .Y(n4016));
  NOR3X1  g01049(.A(n4007), .B(n3708), .C(n3509), .Y(n4017));
  AOI22X1 g01050(.A0(n4016), .A1(n4006), .B0(n4005), .B1(n4017), .Y(n4018));
  NAND4X1 g01051(.A(n4015), .B(n4014), .C(n4013), .D(n4018), .Y(P3_U2994));
  NAND2X1 g01052(.A(n3997), .B(P3_INSTQUEUE_REG_15__5__SCAN_IN), .Y(n4020));
  NAND3X1 g01053(.A(n4001), .B(n3994), .C(BUF2_REG_5__SCAN_IN), .Y(n4021));
  NAND4X1 g01054(.A(n3994), .B(n4003), .C(BUF2_REG_29__SCAN_IN), .D(n3999), .Y(n4022));
  NOR3X1  g01055(.A(n4008), .B(n4007), .C(n3254), .Y(n4023));
  NOR3X1  g01056(.A(n4007), .B(n3650), .C(n3509), .Y(n4024));
  AOI22X1 g01057(.A0(n4023), .A1(n4006), .B0(n4005), .B1(n4024), .Y(n4025));
  NAND4X1 g01058(.A(n4022), .B(n4021), .C(n4020), .D(n4025), .Y(P3_U2993));
  NAND2X1 g01059(.A(n3997), .B(P3_INSTQUEUE_REG_15__4__SCAN_IN), .Y(n4027));
  NAND3X1 g01060(.A(n4001), .B(n3994), .C(BUF2_REG_4__SCAN_IN), .Y(n4028));
  NAND4X1 g01061(.A(n3994), .B(n4003), .C(BUF2_REG_28__SCAN_IN), .D(n3999), .Y(n4029));
  NOR3X1  g01062(.A(n4008), .B(n4007), .C(n3251), .Y(n4030));
  NOR3X1  g01063(.A(n4007), .B(n3634), .C(n3509), .Y(n4031));
  AOI22X1 g01064(.A0(n4030), .A1(n4006), .B0(n4005), .B1(n4031), .Y(n4032));
  NAND4X1 g01065(.A(n4029), .B(n4028), .C(n4027), .D(n4032), .Y(P3_U2992));
  NAND2X1 g01066(.A(n3997), .B(P3_INSTQUEUE_REG_15__3__SCAN_IN), .Y(n4034));
  NAND3X1 g01067(.A(n4001), .B(n3994), .C(BUF2_REG_3__SCAN_IN), .Y(n4035));
  NAND4X1 g01068(.A(n3994), .B(n4003), .C(BUF2_REG_27__SCAN_IN), .D(n3999), .Y(n4036));
  NOR3X1  g01069(.A(n4008), .B(n4007), .C(n3248), .Y(n4037));
  NOR3X1  g01070(.A(n4007), .B(n3616), .C(n3509), .Y(n4038));
  AOI22X1 g01071(.A0(n4037), .A1(n4006), .B0(n4005), .B1(n4038), .Y(n4039));
  NAND4X1 g01072(.A(n4036), .B(n4035), .C(n4034), .D(n4039), .Y(P3_U2991));
  NAND2X1 g01073(.A(n3997), .B(P3_INSTQUEUE_REG_15__2__SCAN_IN), .Y(n4041));
  NAND3X1 g01074(.A(n4001), .B(n3994), .C(BUF2_REG_2__SCAN_IN), .Y(n4042));
  NAND4X1 g01075(.A(n3994), .B(n4003), .C(BUF2_REG_26__SCAN_IN), .D(n3999), .Y(n4043));
  NOR3X1  g01076(.A(n4008), .B(n4007), .C(n3245), .Y(n4044));
  NOR3X1  g01077(.A(n4007), .B(n3583), .C(n3509), .Y(n4045));
  AOI22X1 g01078(.A0(n4044), .A1(n4006), .B0(n4005), .B1(n4045), .Y(n4046));
  NAND4X1 g01079(.A(n4043), .B(n4042), .C(n4041), .D(n4046), .Y(P3_U2990));
  NAND2X1 g01080(.A(n3997), .B(P3_INSTQUEUE_REG_15__1__SCAN_IN), .Y(n4048));
  NAND3X1 g01081(.A(n4001), .B(n3994), .C(BUF2_REG_1__SCAN_IN), .Y(n4049));
  NAND4X1 g01082(.A(n3994), .B(n4003), .C(BUF2_REG_25__SCAN_IN), .D(n3999), .Y(n4050));
  NOR3X1  g01083(.A(n4008), .B(n4007), .C(n3242), .Y(n4051));
  NOR3X1  g01084(.A(n4007), .B(n3681), .C(n3509), .Y(n4052));
  AOI22X1 g01085(.A0(n4051), .A1(n4006), .B0(n4005), .B1(n4052), .Y(n4053));
  NAND4X1 g01086(.A(n4050), .B(n4049), .C(n4048), .D(n4053), .Y(P3_U2989));
  NAND2X1 g01087(.A(n3997), .B(P3_INSTQUEUE_REG_15__0__SCAN_IN), .Y(n4055));
  NAND3X1 g01088(.A(n4001), .B(n3994), .C(BUF2_REG_0__SCAN_IN), .Y(n4056));
  NAND4X1 g01089(.A(n3994), .B(n4003), .C(BUF2_REG_24__SCAN_IN), .D(n3999), .Y(n4057));
  NOR3X1  g01090(.A(n4008), .B(n4007), .C(n3239), .Y(n4058));
  NOR3X1  g01091(.A(n4007), .B(n3698), .C(n3509), .Y(n4059));
  AOI22X1 g01092(.A0(n4058), .A1(n4006), .B0(n4005), .B1(n4059), .Y(n4060));
  NAND4X1 g01093(.A(n4057), .B(n4056), .C(n4055), .D(n4060), .Y(P3_U2988));
  INVX1   g01094(.A(P3_INSTQUEUE_REG_14__7__SCAN_IN), .Y(n4062));
  NOR4X1  g01095(.A(n3518), .B(n3516), .C(n3513), .D(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Y(n4063));
  NOR4X1  g01096(.A(n3518), .B(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C(n3513), .D(n3519), .Y(n4065));
  INVX1   g01097(.A(n4065), .Y(n4066));
  INVX1   g01098(.A(n4003), .Y(n4068));
  AOI21X1 g01099(.A0(n4068), .A1(n4066), .B0(n3989), .Y(n4069));
  NOR3X1  g01100(.A(n4069), .B(n4006), .C(n4063), .Y(n4070));
  OAI21X1 g01101(.A0(n4063), .A1(n3509), .B0(n3994), .Y(n4071));
  NOR2X1  g01102(.A(n4071), .B(n4070), .Y(n4072));
  NOR2X1  g01103(.A(P3_STATE2_REG_2__SCAN_IN), .B(P3_STATE2_REG_3__SCAN_IN), .Y(n4073));
  INVX1   g01104(.A(n4073), .Y(n4074));
  NOR4X1  g01105(.A(n4065), .B(n4074), .C(n3944), .D(n4003), .Y(n4075));
  OAI22X1 g01106(.A0(n4006), .A1(n4063), .B0(n3989), .B1(n4075), .Y(n4076));
  NOR3X1  g01107(.A(n4076), .B(n4007), .C(n3212), .Y(n4077));
  NOR4X1  g01108(.A(n4008), .B(n4007), .C(n3284), .D(n4066), .Y(n4078));
  INVX1   g01109(.A(n4009), .Y(n4079));
  INVX1   g01110(.A(n4010), .Y(n4080));
  INVX1   g01111(.A(n4063), .Y(n4081));
  OAI22X1 g01112(.A0(n4081), .A1(n4080), .B0(n4079), .B1(n4068), .Y(n4082));
  NOR3X1  g01113(.A(n4082), .B(n4078), .C(n4077), .Y(n4083));
  OAI21X1 g01114(.A0(n4072), .A1(n4062), .B0(n4083), .Y(P3_U2987));
  INVX1   g01115(.A(P3_INSTQUEUE_REG_14__6__SCAN_IN), .Y(n4085));
  NOR3X1  g01116(.A(n4076), .B(n4007), .C(n3209), .Y(n4086));
  NOR4X1  g01117(.A(n4008), .B(n4007), .C(n3281), .D(n4066), .Y(n4087));
  INVX1   g01118(.A(n4016), .Y(n4088));
  INVX1   g01119(.A(n4017), .Y(n4089));
  OAI22X1 g01120(.A0(n4081), .A1(n4089), .B0(n4088), .B1(n4068), .Y(n4090));
  NOR3X1  g01121(.A(n4090), .B(n4087), .C(n4086), .Y(n4091));
  OAI21X1 g01122(.A0(n4072), .A1(n4085), .B0(n4091), .Y(P3_U2986));
  INVX1   g01123(.A(P3_INSTQUEUE_REG_14__5__SCAN_IN), .Y(n4093));
  NOR3X1  g01124(.A(n4076), .B(n4007), .C(n3206), .Y(n4094));
  NOR4X1  g01125(.A(n4008), .B(n4007), .C(n3278), .D(n4066), .Y(n4095));
  INVX1   g01126(.A(n4023), .Y(n4096));
  INVX1   g01127(.A(n4024), .Y(n4097));
  OAI22X1 g01128(.A0(n4081), .A1(n4097), .B0(n4096), .B1(n4068), .Y(n4098));
  NOR3X1  g01129(.A(n4098), .B(n4095), .C(n4094), .Y(n4099));
  OAI21X1 g01130(.A0(n4072), .A1(n4093), .B0(n4099), .Y(P3_U2985));
  INVX1   g01131(.A(P3_INSTQUEUE_REG_14__4__SCAN_IN), .Y(n4101));
  NOR3X1  g01132(.A(n4076), .B(n4007), .C(n3203), .Y(n4102));
  NOR4X1  g01133(.A(n4008), .B(n4007), .C(n3275), .D(n4066), .Y(n4103));
  INVX1   g01134(.A(n4030), .Y(n4104));
  INVX1   g01135(.A(n4031), .Y(n4105));
  OAI22X1 g01136(.A0(n4081), .A1(n4105), .B0(n4104), .B1(n4068), .Y(n4106));
  NOR3X1  g01137(.A(n4106), .B(n4103), .C(n4102), .Y(n4107));
  OAI21X1 g01138(.A0(n4072), .A1(n4101), .B0(n4107), .Y(P3_U2984));
  INVX1   g01139(.A(P3_INSTQUEUE_REG_14__3__SCAN_IN), .Y(n4109));
  NOR3X1  g01140(.A(n4076), .B(n4007), .C(n3200), .Y(n4110));
  NOR4X1  g01141(.A(n4008), .B(n4007), .C(n3272), .D(n4066), .Y(n4111));
  INVX1   g01142(.A(n4037), .Y(n4112));
  INVX1   g01143(.A(n4038), .Y(n4113));
  OAI22X1 g01144(.A0(n4081), .A1(n4113), .B0(n4112), .B1(n4068), .Y(n4114));
  NOR3X1  g01145(.A(n4114), .B(n4111), .C(n4110), .Y(n4115));
  OAI21X1 g01146(.A0(n4072), .A1(n4109), .B0(n4115), .Y(P3_U2983));
  INVX1   g01147(.A(P3_INSTQUEUE_REG_14__2__SCAN_IN), .Y(n4117));
  NOR3X1  g01148(.A(n4076), .B(n4007), .C(n3197), .Y(n4118));
  NOR4X1  g01149(.A(n4008), .B(n4007), .C(n3269), .D(n4066), .Y(n4119));
  INVX1   g01150(.A(n4044), .Y(n4120));
  INVX1   g01151(.A(n4045), .Y(n4121));
  OAI22X1 g01152(.A0(n4081), .A1(n4121), .B0(n4120), .B1(n4068), .Y(n4122));
  NOR3X1  g01153(.A(n4122), .B(n4119), .C(n4118), .Y(n4123));
  OAI21X1 g01154(.A0(n4072), .A1(n4117), .B0(n4123), .Y(P3_U2982));
  INVX1   g01155(.A(P3_INSTQUEUE_REG_14__1__SCAN_IN), .Y(n4125));
  NOR3X1  g01156(.A(n4076), .B(n4007), .C(n3194), .Y(n4126));
  NOR4X1  g01157(.A(n4008), .B(n4007), .C(n3266), .D(n4066), .Y(n4127));
  INVX1   g01158(.A(n4051), .Y(n4128));
  INVX1   g01159(.A(n4052), .Y(n4129));
  OAI22X1 g01160(.A0(n4081), .A1(n4129), .B0(n4128), .B1(n4068), .Y(n4130));
  NOR3X1  g01161(.A(n4130), .B(n4127), .C(n4126), .Y(n4131));
  OAI21X1 g01162(.A0(n4072), .A1(n4125), .B0(n4131), .Y(P3_U2981));
  INVX1   g01163(.A(P3_INSTQUEUE_REG_14__0__SCAN_IN), .Y(n4133));
  NOR3X1  g01164(.A(n4076), .B(n4007), .C(n3190), .Y(n4134));
  NOR4X1  g01165(.A(n4008), .B(n4007), .C(n3263), .D(n4066), .Y(n4135));
  INVX1   g01166(.A(n4058), .Y(n4136));
  INVX1   g01167(.A(n4059), .Y(n4137));
  OAI22X1 g01168(.A0(n4081), .A1(n4137), .B0(n4136), .B1(n4068), .Y(n4138));
  NOR3X1  g01169(.A(n4138), .B(n4135), .C(n4134), .Y(n4139));
  OAI21X1 g01170(.A0(n4072), .A1(n4133), .B0(n4139), .Y(P3_U2980));
  NAND3X1 g01171(.A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n3516), .C(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .Y(n4142));
  OAI21X1 g01172(.A0(n4142), .A1(n3989), .B0(n3990), .Y(n4143));
  NAND2X1 g01173(.A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n3518), .Y(n4144));
  NAND2X1 g01174(.A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .Y(n4145));
  OAI21X1 g01175(.A0(n4145), .A1(n4144), .B0(P3_STATE2_REG_3__SCAN_IN), .Y(n4146));
  NAND3X1 g01176(.A(n4146), .B(n4143), .C(n3994), .Y(n4147));
  NAND2X1 g01177(.A(n4147), .B(P3_INSTQUEUE_REG_13__7__SCAN_IN), .Y(n4148));
  NAND2X1 g01178(.A(n4142), .B(n3999), .Y(n4149));
  AOI21X1 g01179(.A0(n4149), .A1(n3988), .B0(n3990), .Y(n4150));
  NAND3X1 g01180(.A(n4150), .B(n3994), .C(BUF2_REG_7__SCAN_IN), .Y(n4151));
  NOR4X1  g01181(.A(n3518), .B(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C(n3513), .D(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Y(n4152));
  NAND4X1 g01182(.A(n3999), .B(n3994), .C(BUF2_REG_31__SCAN_IN), .D(n4152), .Y(n4153));
  AOI22X1 g01183(.A0(n4006), .A1(n4010), .B0(n4009), .B1(n4065), .Y(n4156));
  NAND4X1 g01184(.A(n4153), .B(n4151), .C(n4148), .D(n4156), .Y(P3_U2979));
  NAND2X1 g01185(.A(n4147), .B(P3_INSTQUEUE_REG_13__6__SCAN_IN), .Y(n4158));
  NAND3X1 g01186(.A(n4150), .B(n3994), .C(BUF2_REG_6__SCAN_IN), .Y(n4159));
  NAND4X1 g01187(.A(n3999), .B(n3994), .C(BUF2_REG_30__SCAN_IN), .D(n4152), .Y(n4160));
  AOI22X1 g01188(.A0(n4006), .A1(n4017), .B0(n4016), .B1(n4065), .Y(n4161));
  NAND4X1 g01189(.A(n4160), .B(n4159), .C(n4158), .D(n4161), .Y(P3_U2978));
  NAND2X1 g01190(.A(n4147), .B(P3_INSTQUEUE_REG_13__5__SCAN_IN), .Y(n4163));
  NAND3X1 g01191(.A(n4150), .B(n3994), .C(BUF2_REG_5__SCAN_IN), .Y(n4164));
  NAND4X1 g01192(.A(n3999), .B(n3994), .C(BUF2_REG_29__SCAN_IN), .D(n4152), .Y(n4165));
  AOI22X1 g01193(.A0(n4006), .A1(n4024), .B0(n4023), .B1(n4065), .Y(n4166));
  NAND4X1 g01194(.A(n4165), .B(n4164), .C(n4163), .D(n4166), .Y(P3_U2977));
  NAND2X1 g01195(.A(n4147), .B(P3_INSTQUEUE_REG_13__4__SCAN_IN), .Y(n4168));
  NAND3X1 g01196(.A(n4150), .B(n3994), .C(BUF2_REG_4__SCAN_IN), .Y(n4169));
  NAND4X1 g01197(.A(n3999), .B(n3994), .C(BUF2_REG_28__SCAN_IN), .D(n4152), .Y(n4170));
  AOI22X1 g01198(.A0(n4006), .A1(n4031), .B0(n4030), .B1(n4065), .Y(n4171));
  NAND4X1 g01199(.A(n4170), .B(n4169), .C(n4168), .D(n4171), .Y(P3_U2976));
  NAND2X1 g01200(.A(n4147), .B(P3_INSTQUEUE_REG_13__3__SCAN_IN), .Y(n4173));
  NAND3X1 g01201(.A(n4150), .B(n3994), .C(BUF2_REG_3__SCAN_IN), .Y(n4174));
  NAND4X1 g01202(.A(n3999), .B(n3994), .C(BUF2_REG_27__SCAN_IN), .D(n4152), .Y(n4175));
  AOI22X1 g01203(.A0(n4006), .A1(n4038), .B0(n4037), .B1(n4065), .Y(n4176));
  NAND4X1 g01204(.A(n4175), .B(n4174), .C(n4173), .D(n4176), .Y(P3_U2975));
  NAND2X1 g01205(.A(n4147), .B(P3_INSTQUEUE_REG_13__2__SCAN_IN), .Y(n4178));
  NAND3X1 g01206(.A(n4150), .B(n3994), .C(BUF2_REG_2__SCAN_IN), .Y(n4179));
  NAND4X1 g01207(.A(n3999), .B(n3994), .C(BUF2_REG_26__SCAN_IN), .D(n4152), .Y(n4180));
  AOI22X1 g01208(.A0(n4006), .A1(n4045), .B0(n4044), .B1(n4065), .Y(n4181));
  NAND4X1 g01209(.A(n4180), .B(n4179), .C(n4178), .D(n4181), .Y(P3_U2974));
  NAND2X1 g01210(.A(n4147), .B(P3_INSTQUEUE_REG_13__1__SCAN_IN), .Y(n4183));
  NAND3X1 g01211(.A(n4150), .B(n3994), .C(BUF2_REG_1__SCAN_IN), .Y(n4184));
  NAND4X1 g01212(.A(n3999), .B(n3994), .C(BUF2_REG_25__SCAN_IN), .D(n4152), .Y(n4185));
  AOI22X1 g01213(.A0(n4006), .A1(n4052), .B0(n4051), .B1(n4065), .Y(n4186));
  NAND4X1 g01214(.A(n4185), .B(n4184), .C(n4183), .D(n4186), .Y(P3_U2973));
  NAND2X1 g01215(.A(n4147), .B(P3_INSTQUEUE_REG_13__0__SCAN_IN), .Y(n4188));
  NAND3X1 g01216(.A(n4150), .B(n3994), .C(BUF2_REG_0__SCAN_IN), .Y(n4189));
  NAND4X1 g01217(.A(n3999), .B(n3994), .C(BUF2_REG_24__SCAN_IN), .D(n4152), .Y(n4190));
  AOI22X1 g01218(.A0(n4006), .A1(n4059), .B0(n4058), .B1(n4065), .Y(n4191));
  NAND4X1 g01219(.A(n4190), .B(n4189), .C(n4188), .D(n4191), .Y(P3_U2972));
  INVX1   g01220(.A(P3_INSTQUEUE_REG_12__7__SCAN_IN), .Y(n4193));
  NAND2X1 g01221(.A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Y(n4194));
  XOR2X1  g01222(.A(n4194), .B(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .Y(n4195));
  XOR2X1  g01223(.A(n3995), .B(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .Y(n4196));
  XOR2X1  g01224(.A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n3518), .Y(n4197));
  NOR3X1  g01225(.A(n4957), .B(n4196), .C(n4195), .Y(n4199));
  NOR4X1  g01226(.A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C(n3513), .D(n3519), .Y(n4200));
  INVX1   g01227(.A(n4200), .Y(n4201));
  INVX1   g01228(.A(n4152), .Y(n4203));
  AOI21X1 g01229(.A0(n4203), .A1(n4201), .B0(n3989), .Y(n4204));
  NOR2X1  g01230(.A(n4204), .B(n4199), .Y(n4205));
  OAI21X1 g01231(.A0(n4003), .A1(n3509), .B0(n3994), .Y(n4207));
  NOR2X1  g01232(.A(n4207), .B(n4205), .Y(n4208));
  NOR4X1  g01233(.A(n4200), .B(n4074), .C(n3944), .D(n4152), .Y(n4209));
  OAI21X1 g01234(.A0(n4209), .A1(n3989), .B0(n4199), .Y(n4210));
  NOR3X1  g01235(.A(n4210), .B(n4007), .C(n3212), .Y(n4211));
  NOR4X1  g01236(.A(n4008), .B(n4007), .C(n3284), .D(n4201), .Y(n4212));
  OAI22X1 g01237(.A0(n4203), .A1(n4079), .B0(n4080), .B1(n4068), .Y(n4214));
  NOR3X1  g01238(.A(n4214), .B(n4212), .C(n4211), .Y(n4215));
  OAI21X1 g01239(.A0(n4208), .A1(n4193), .B0(n4215), .Y(P3_U2971));
  INVX1   g01240(.A(P3_INSTQUEUE_REG_12__6__SCAN_IN), .Y(n4217));
  NOR3X1  g01241(.A(n4210), .B(n4007), .C(n3209), .Y(n4218));
  NOR4X1  g01242(.A(n4008), .B(n4007), .C(n3281), .D(n4201), .Y(n4219));
  OAI22X1 g01243(.A0(n4203), .A1(n4088), .B0(n4089), .B1(n4068), .Y(n4220));
  NOR3X1  g01244(.A(n4220), .B(n4219), .C(n4218), .Y(n4221));
  OAI21X1 g01245(.A0(n4208), .A1(n4217), .B0(n4221), .Y(P3_U2970));
  INVX1   g01246(.A(P3_INSTQUEUE_REG_12__5__SCAN_IN), .Y(n4223));
  NOR3X1  g01247(.A(n4210), .B(n4007), .C(n3206), .Y(n4224));
  NOR4X1  g01248(.A(n4008), .B(n4007), .C(n3278), .D(n4201), .Y(n4225));
  OAI22X1 g01249(.A0(n4203), .A1(n4096), .B0(n4097), .B1(n4068), .Y(n4226));
  NOR3X1  g01250(.A(n4226), .B(n4225), .C(n4224), .Y(n4227));
  OAI21X1 g01251(.A0(n4208), .A1(n4223), .B0(n4227), .Y(P3_U2969));
  INVX1   g01252(.A(P3_INSTQUEUE_REG_12__4__SCAN_IN), .Y(n4229));
  NOR3X1  g01253(.A(n4210), .B(n4007), .C(n3203), .Y(n4230));
  NOR4X1  g01254(.A(n4008), .B(n4007), .C(n3275), .D(n4201), .Y(n4231));
  OAI22X1 g01255(.A0(n4203), .A1(n4104), .B0(n4105), .B1(n4068), .Y(n4232));
  NOR3X1  g01256(.A(n4232), .B(n4231), .C(n4230), .Y(n4233));
  OAI21X1 g01257(.A0(n4208), .A1(n4229), .B0(n4233), .Y(P3_U2968));
  INVX1   g01258(.A(P3_INSTQUEUE_REG_12__3__SCAN_IN), .Y(n4235));
  NOR3X1  g01259(.A(n4210), .B(n4007), .C(n3200), .Y(n4236));
  NOR4X1  g01260(.A(n4008), .B(n4007), .C(n3272), .D(n4201), .Y(n4237));
  OAI22X1 g01261(.A0(n4203), .A1(n4112), .B0(n4113), .B1(n4068), .Y(n4238));
  NOR3X1  g01262(.A(n4238), .B(n4237), .C(n4236), .Y(n4239));
  OAI21X1 g01263(.A0(n4208), .A1(n4235), .B0(n4239), .Y(P3_U2967));
  INVX1   g01264(.A(P3_INSTQUEUE_REG_12__2__SCAN_IN), .Y(n4241));
  NOR3X1  g01265(.A(n4210), .B(n4007), .C(n3197), .Y(n4242));
  NOR4X1  g01266(.A(n4008), .B(n4007), .C(n3269), .D(n4201), .Y(n4243));
  OAI22X1 g01267(.A0(n4203), .A1(n4120), .B0(n4121), .B1(n4068), .Y(n4244));
  NOR3X1  g01268(.A(n4244), .B(n4243), .C(n4242), .Y(n4245));
  OAI21X1 g01269(.A0(n4208), .A1(n4241), .B0(n4245), .Y(P3_U2966));
  INVX1   g01270(.A(P3_INSTQUEUE_REG_12__1__SCAN_IN), .Y(n4247));
  NOR3X1  g01271(.A(n4210), .B(n4007), .C(n3194), .Y(n4248));
  NOR4X1  g01272(.A(n4008), .B(n4007), .C(n3266), .D(n4201), .Y(n4249));
  OAI22X1 g01273(.A0(n4203), .A1(n4128), .B0(n4129), .B1(n4068), .Y(n4250));
  NOR3X1  g01274(.A(n4250), .B(n4249), .C(n4248), .Y(n4251));
  OAI21X1 g01275(.A0(n4208), .A1(n4247), .B0(n4251), .Y(P3_U2965));
  INVX1   g01276(.A(P3_INSTQUEUE_REG_12__0__SCAN_IN), .Y(n4253));
  NOR3X1  g01277(.A(n4210), .B(n4007), .C(n3190), .Y(n4254));
  NOR4X1  g01278(.A(n4008), .B(n4007), .C(n3263), .D(n4201), .Y(n4255));
  OAI22X1 g01279(.A0(n4203), .A1(n4136), .B0(n4137), .B1(n4068), .Y(n4256));
  NOR3X1  g01280(.A(n4256), .B(n4255), .C(n4254), .Y(n4257));
  OAI21X1 g01281(.A0(n4208), .A1(n4253), .B0(n4257), .Y(P3_U2964));
  NAND3X1 g01282(.A(n3518), .B(n3516), .C(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .Y(n4260));
  OAI21X1 g01283(.A0(n4260), .A1(n3989), .B0(n4142), .Y(n4261));
  NAND3X1 g01284(.A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C(n3516), .Y(n4262));
  OAI21X1 g01285(.A0(n4262), .A1(n3513), .B0(P3_STATE2_REG_3__SCAN_IN), .Y(n4263));
  NAND3X1 g01286(.A(n4263), .B(n4261), .C(n3994), .Y(n4264));
  NAND2X1 g01287(.A(n4264), .B(P3_INSTQUEUE_REG_11__7__SCAN_IN), .Y(n4265));
  NAND2X1 g01288(.A(n4260), .B(n3999), .Y(n4266));
  AOI21X1 g01289(.A0(n4266), .A1(n3988), .B0(n4142), .Y(n4267));
  NAND3X1 g01290(.A(n4267), .B(n3994), .C(BUF2_REG_7__SCAN_IN), .Y(n4268));
  NOR4X1  g01291(.A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C(n3513), .D(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Y(n4269));
  NAND4X1 g01292(.A(n3999), .B(n3994), .C(BUF2_REG_31__SCAN_IN), .D(n4269), .Y(n4270));
  AOI22X1 g01293(.A0(n4065), .A1(n4010), .B0(n4009), .B1(n4200), .Y(n4273));
  NAND4X1 g01294(.A(n4270), .B(n4268), .C(n4265), .D(n4273), .Y(P3_U2963));
  NAND2X1 g01295(.A(n4264), .B(P3_INSTQUEUE_REG_11__6__SCAN_IN), .Y(n4275));
  NAND3X1 g01296(.A(n4267), .B(n3994), .C(BUF2_REG_6__SCAN_IN), .Y(n4276));
  NAND4X1 g01297(.A(n3999), .B(n3994), .C(BUF2_REG_30__SCAN_IN), .D(n4269), .Y(n4277));
  AOI22X1 g01298(.A0(n4065), .A1(n4017), .B0(n4016), .B1(n4200), .Y(n4278));
  NAND4X1 g01299(.A(n4277), .B(n4276), .C(n4275), .D(n4278), .Y(P3_U2962));
  NAND2X1 g01300(.A(n4264), .B(P3_INSTQUEUE_REG_11__5__SCAN_IN), .Y(n4280));
  NAND3X1 g01301(.A(n4267), .B(n3994), .C(BUF2_REG_5__SCAN_IN), .Y(n4281));
  NAND4X1 g01302(.A(n3999), .B(n3994), .C(BUF2_REG_29__SCAN_IN), .D(n4269), .Y(n4282));
  AOI22X1 g01303(.A0(n4065), .A1(n4024), .B0(n4023), .B1(n4200), .Y(n4283));
  NAND4X1 g01304(.A(n4282), .B(n4281), .C(n4280), .D(n4283), .Y(P3_U2961));
  NAND2X1 g01305(.A(n4264), .B(P3_INSTQUEUE_REG_11__4__SCAN_IN), .Y(n4285));
  NAND3X1 g01306(.A(n4267), .B(n3994), .C(BUF2_REG_4__SCAN_IN), .Y(n4286));
  NAND4X1 g01307(.A(n3999), .B(n3994), .C(BUF2_REG_28__SCAN_IN), .D(n4269), .Y(n4287));
  AOI22X1 g01308(.A0(n4065), .A1(n4031), .B0(n4030), .B1(n4200), .Y(n4288));
  NAND4X1 g01309(.A(n4287), .B(n4286), .C(n4285), .D(n4288), .Y(P3_U2960));
  NAND2X1 g01310(.A(n4264), .B(P3_INSTQUEUE_REG_11__3__SCAN_IN), .Y(n4290));
  NAND3X1 g01311(.A(n4267), .B(n3994), .C(BUF2_REG_3__SCAN_IN), .Y(n4291));
  NAND4X1 g01312(.A(n3999), .B(n3994), .C(BUF2_REG_27__SCAN_IN), .D(n4269), .Y(n4292));
  AOI22X1 g01313(.A0(n4065), .A1(n4038), .B0(n4037), .B1(n4200), .Y(n4293));
  NAND4X1 g01314(.A(n4292), .B(n4291), .C(n4290), .D(n4293), .Y(P3_U2959));
  NAND2X1 g01315(.A(n4264), .B(P3_INSTQUEUE_REG_11__2__SCAN_IN), .Y(n4295));
  NAND3X1 g01316(.A(n4267), .B(n3994), .C(BUF2_REG_2__SCAN_IN), .Y(n4296));
  NAND4X1 g01317(.A(n3999), .B(n3994), .C(BUF2_REG_26__SCAN_IN), .D(n4269), .Y(n4297));
  AOI22X1 g01318(.A0(n4065), .A1(n4045), .B0(n4044), .B1(n4200), .Y(n4298));
  NAND4X1 g01319(.A(n4297), .B(n4296), .C(n4295), .D(n4298), .Y(P3_U2958));
  NAND2X1 g01320(.A(n4264), .B(P3_INSTQUEUE_REG_11__1__SCAN_IN), .Y(n4300));
  NAND3X1 g01321(.A(n4267), .B(n3994), .C(BUF2_REG_1__SCAN_IN), .Y(n4301));
  NAND4X1 g01322(.A(n3999), .B(n3994), .C(BUF2_REG_25__SCAN_IN), .D(n4269), .Y(n4302));
  AOI22X1 g01323(.A0(n4065), .A1(n4052), .B0(n4051), .B1(n4200), .Y(n4303));
  NAND4X1 g01324(.A(n4302), .B(n4301), .C(n4300), .D(n4303), .Y(P3_U2957));
  NAND2X1 g01325(.A(n4264), .B(P3_INSTQUEUE_REG_11__0__SCAN_IN), .Y(n4305));
  NAND3X1 g01326(.A(n4267), .B(n3994), .C(BUF2_REG_0__SCAN_IN), .Y(n4306));
  NAND4X1 g01327(.A(n3999), .B(n3994), .C(BUF2_REG_24__SCAN_IN), .D(n4269), .Y(n4307));
  AOI22X1 g01328(.A0(n4065), .A1(n4059), .B0(n4058), .B1(n4200), .Y(n4308));
  NAND4X1 g01329(.A(n4307), .B(n4306), .C(n4305), .D(n4308), .Y(P3_U2956));
  INVX1   g01330(.A(P3_INSTQUEUE_REG_10__7__SCAN_IN), .Y(n4310));
  NOR4X1  g01331(.A(n3518), .B(n3516), .C(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .D(n3519), .Y(n4313));
  INVX1   g01332(.A(n4313), .Y(n4314));
  INVX1   g01333(.A(n4269), .Y(n4316));
  AOI21X1 g01334(.A0(n4316), .A1(n4314), .B0(n3989), .Y(n4317));
  NOR3X1  g01335(.A(n4317), .B(n4200), .C(n4152), .Y(n4318));
  OAI21X1 g01336(.A0(n4152), .A1(n3509), .B0(n3994), .Y(n4319));
  NOR2X1  g01337(.A(n4319), .B(n4318), .Y(n4320));
  NOR4X1  g01338(.A(n4313), .B(n4074), .C(n3944), .D(n4269), .Y(n4321));
  OAI22X1 g01339(.A0(n4200), .A1(n4152), .B0(n3989), .B1(n4321), .Y(n4322));
  NOR3X1  g01340(.A(n4322), .B(n4007), .C(n3212), .Y(n4323));
  NOR4X1  g01341(.A(n4008), .B(n4007), .C(n3284), .D(n4314), .Y(n4324));
  OAI22X1 g01342(.A0(n4203), .A1(n4080), .B0(n4079), .B1(n4316), .Y(n4326));
  NOR3X1  g01343(.A(n4326), .B(n4324), .C(n4323), .Y(n4327));
  OAI21X1 g01344(.A0(n4320), .A1(n4310), .B0(n4327), .Y(P3_U2955));
  INVX1   g01345(.A(P3_INSTQUEUE_REG_10__6__SCAN_IN), .Y(n4329));
  NOR3X1  g01346(.A(n4322), .B(n4007), .C(n3209), .Y(n4330));
  NOR4X1  g01347(.A(n4008), .B(n4007), .C(n3281), .D(n4314), .Y(n4331));
  OAI22X1 g01348(.A0(n4203), .A1(n4089), .B0(n4088), .B1(n4316), .Y(n4332));
  NOR3X1  g01349(.A(n4332), .B(n4331), .C(n4330), .Y(n4333));
  OAI21X1 g01350(.A0(n4320), .A1(n4329), .B0(n4333), .Y(P3_U2954));
  INVX1   g01351(.A(P3_INSTQUEUE_REG_10__5__SCAN_IN), .Y(n4335));
  NOR3X1  g01352(.A(n4322), .B(n4007), .C(n3206), .Y(n4336));
  NOR4X1  g01353(.A(n4008), .B(n4007), .C(n3278), .D(n4314), .Y(n4337));
  OAI22X1 g01354(.A0(n4203), .A1(n4097), .B0(n4096), .B1(n4316), .Y(n4338));
  NOR3X1  g01355(.A(n4338), .B(n4337), .C(n4336), .Y(n4339));
  OAI21X1 g01356(.A0(n4320), .A1(n4335), .B0(n4339), .Y(P3_U2953));
  INVX1   g01357(.A(P3_INSTQUEUE_REG_10__4__SCAN_IN), .Y(n4341));
  NOR3X1  g01358(.A(n4322), .B(n4007), .C(n3203), .Y(n4342));
  NOR4X1  g01359(.A(n4008), .B(n4007), .C(n3275), .D(n4314), .Y(n4343));
  OAI22X1 g01360(.A0(n4203), .A1(n4105), .B0(n4104), .B1(n4316), .Y(n4344));
  NOR3X1  g01361(.A(n4344), .B(n4343), .C(n4342), .Y(n4345));
  OAI21X1 g01362(.A0(n4320), .A1(n4341), .B0(n4345), .Y(P3_U2952));
  INVX1   g01363(.A(P3_INSTQUEUE_REG_10__3__SCAN_IN), .Y(n4347));
  NOR3X1  g01364(.A(n4322), .B(n4007), .C(n3200), .Y(n4348));
  NOR4X1  g01365(.A(n4008), .B(n4007), .C(n3272), .D(n4314), .Y(n4349));
  OAI22X1 g01366(.A0(n4203), .A1(n4113), .B0(n4112), .B1(n4316), .Y(n4350));
  NOR3X1  g01367(.A(n4350), .B(n4349), .C(n4348), .Y(n4351));
  OAI21X1 g01368(.A0(n4320), .A1(n4347), .B0(n4351), .Y(P3_U2951));
  INVX1   g01369(.A(P3_INSTQUEUE_REG_10__2__SCAN_IN), .Y(n4353));
  NOR3X1  g01370(.A(n4322), .B(n4007), .C(n3197), .Y(n4354));
  NOR4X1  g01371(.A(n4008), .B(n4007), .C(n3269), .D(n4314), .Y(n4355));
  OAI22X1 g01372(.A0(n4203), .A1(n4121), .B0(n4120), .B1(n4316), .Y(n4356));
  NOR3X1  g01373(.A(n4356), .B(n4355), .C(n4354), .Y(n4357));
  OAI21X1 g01374(.A0(n4320), .A1(n4353), .B0(n4357), .Y(P3_U2950));
  INVX1   g01375(.A(P3_INSTQUEUE_REG_10__1__SCAN_IN), .Y(n4359));
  NOR3X1  g01376(.A(n4322), .B(n4007), .C(n3194), .Y(n4360));
  NOR4X1  g01377(.A(n4008), .B(n4007), .C(n3266), .D(n4314), .Y(n4361));
  OAI22X1 g01378(.A0(n4203), .A1(n4129), .B0(n4128), .B1(n4316), .Y(n4362));
  NOR3X1  g01379(.A(n4362), .B(n4361), .C(n4360), .Y(n4363));
  OAI21X1 g01380(.A0(n4320), .A1(n4359), .B0(n4363), .Y(P3_U2949));
  INVX1   g01381(.A(P3_INSTQUEUE_REG_10__0__SCAN_IN), .Y(n4365));
  NOR3X1  g01382(.A(n4322), .B(n4007), .C(n3190), .Y(n4366));
  NOR4X1  g01383(.A(n4008), .B(n4007), .C(n3263), .D(n4314), .Y(n4367));
  OAI22X1 g01384(.A0(n4203), .A1(n4137), .B0(n4136), .B1(n4316), .Y(n4368));
  NOR3X1  g01385(.A(n4368), .B(n4367), .C(n4366), .Y(n4369));
  OAI21X1 g01386(.A0(n4320), .A1(n4365), .B0(n4369), .Y(P3_U2948));
  NAND3X1 g01387(.A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C(n3513), .Y(n4372));
  OAI21X1 g01388(.A0(n4372), .A1(n3989), .B0(n4260), .Y(n4373));
  NAND2X1 g01389(.A(n3516), .B(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .Y(n4374));
  OAI21X1 g01390(.A0(n4374), .A1(n4144), .B0(P3_STATE2_REG_3__SCAN_IN), .Y(n4375));
  NAND3X1 g01391(.A(n4375), .B(n4373), .C(n3994), .Y(n4376));
  NAND2X1 g01392(.A(n4376), .B(P3_INSTQUEUE_REG_9__7__SCAN_IN), .Y(n4377));
  NAND2X1 g01393(.A(n4372), .B(n3999), .Y(n4378));
  AOI21X1 g01394(.A0(n4378), .A1(n3988), .B0(n4260), .Y(n4379));
  NAND3X1 g01395(.A(n4379), .B(n3994), .C(BUF2_REG_7__SCAN_IN), .Y(n4380));
  NOR4X1  g01396(.A(n3518), .B(n3516), .C(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .D(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Y(n4381));
  NAND4X1 g01397(.A(n3999), .B(n3994), .C(BUF2_REG_31__SCAN_IN), .D(n4381), .Y(n4382));
  AOI22X1 g01398(.A0(n4200), .A1(n4010), .B0(n4009), .B1(n4313), .Y(n4385));
  NAND4X1 g01399(.A(n4382), .B(n4380), .C(n4377), .D(n4385), .Y(P3_U2947));
  NAND2X1 g01400(.A(n4376), .B(P3_INSTQUEUE_REG_9__6__SCAN_IN), .Y(n4387));
  NAND3X1 g01401(.A(n4379), .B(n3994), .C(BUF2_REG_6__SCAN_IN), .Y(n4388));
  NAND4X1 g01402(.A(n3999), .B(n3994), .C(BUF2_REG_30__SCAN_IN), .D(n4381), .Y(n4389));
  AOI22X1 g01403(.A0(n4200), .A1(n4017), .B0(n4016), .B1(n4313), .Y(n4390));
  NAND4X1 g01404(.A(n4389), .B(n4388), .C(n4387), .D(n4390), .Y(P3_U2946));
  NAND2X1 g01405(.A(n4376), .B(P3_INSTQUEUE_REG_9__5__SCAN_IN), .Y(n4392));
  NAND3X1 g01406(.A(n4379), .B(n3994), .C(BUF2_REG_5__SCAN_IN), .Y(n4393));
  NAND4X1 g01407(.A(n3999), .B(n3994), .C(BUF2_REG_29__SCAN_IN), .D(n4381), .Y(n4394));
  AOI22X1 g01408(.A0(n4200), .A1(n4024), .B0(n4023), .B1(n4313), .Y(n4395));
  NAND4X1 g01409(.A(n4394), .B(n4393), .C(n4392), .D(n4395), .Y(P3_U2945));
  NAND2X1 g01410(.A(n4376), .B(P3_INSTQUEUE_REG_9__4__SCAN_IN), .Y(n4397));
  NAND3X1 g01411(.A(n4379), .B(n3994), .C(BUF2_REG_4__SCAN_IN), .Y(n4398));
  NAND4X1 g01412(.A(n3999), .B(n3994), .C(BUF2_REG_28__SCAN_IN), .D(n4381), .Y(n4399));
  AOI22X1 g01413(.A0(n4200), .A1(n4031), .B0(n4030), .B1(n4313), .Y(n4400));
  NAND4X1 g01414(.A(n4399), .B(n4398), .C(n4397), .D(n4400), .Y(P3_U2944));
  NAND2X1 g01415(.A(n4376), .B(P3_INSTQUEUE_REG_9__3__SCAN_IN), .Y(n4402));
  NAND3X1 g01416(.A(n4379), .B(n3994), .C(BUF2_REG_3__SCAN_IN), .Y(n4403));
  NAND4X1 g01417(.A(n3999), .B(n3994), .C(BUF2_REG_27__SCAN_IN), .D(n4381), .Y(n4404));
  AOI22X1 g01418(.A0(n4200), .A1(n4038), .B0(n4037), .B1(n4313), .Y(n4405));
  NAND4X1 g01419(.A(n4404), .B(n4403), .C(n4402), .D(n4405), .Y(P3_U2943));
  NAND2X1 g01420(.A(n4376), .B(P3_INSTQUEUE_REG_9__2__SCAN_IN), .Y(n4407));
  NAND3X1 g01421(.A(n4379), .B(n3994), .C(BUF2_REG_2__SCAN_IN), .Y(n4408));
  NAND4X1 g01422(.A(n3999), .B(n3994), .C(BUF2_REG_26__SCAN_IN), .D(n4381), .Y(n4409));
  AOI22X1 g01423(.A0(n4200), .A1(n4045), .B0(n4044), .B1(n4313), .Y(n4410));
  NAND4X1 g01424(.A(n4409), .B(n4408), .C(n4407), .D(n4410), .Y(P3_U2942));
  NAND2X1 g01425(.A(n4376), .B(P3_INSTQUEUE_REG_9__1__SCAN_IN), .Y(n4412));
  NAND3X1 g01426(.A(n4379), .B(n3994), .C(BUF2_REG_1__SCAN_IN), .Y(n4413));
  NAND4X1 g01427(.A(n3999), .B(n3994), .C(BUF2_REG_25__SCAN_IN), .D(n4381), .Y(n4414));
  AOI22X1 g01428(.A0(n4200), .A1(n4052), .B0(n4051), .B1(n4313), .Y(n4415));
  NAND4X1 g01429(.A(n4414), .B(n4413), .C(n4412), .D(n4415), .Y(P3_U2941));
  NAND2X1 g01430(.A(n4376), .B(P3_INSTQUEUE_REG_9__0__SCAN_IN), .Y(n4417));
  NAND3X1 g01431(.A(n4379), .B(n3994), .C(BUF2_REG_0__SCAN_IN), .Y(n4418));
  NAND4X1 g01432(.A(n3999), .B(n3994), .C(BUF2_REG_24__SCAN_IN), .D(n4381), .Y(n4419));
  AOI22X1 g01433(.A0(n4200), .A1(n4059), .B0(n4058), .B1(n4313), .Y(n4420));
  NAND4X1 g01434(.A(n4419), .B(n4418), .C(n4417), .D(n4420), .Y(P3_U2940));
  INVX1   g01435(.A(P3_INSTQUEUE_REG_8__7__SCAN_IN), .Y(n4422));
  INVX1   g01436(.A(n4195), .Y(n4423));
  NOR3X1  g01437(.A(n4957), .B(n4196), .C(n4423), .Y(n4424));
  NOR4X1  g01438(.A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n3516), .C(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .D(n3519), .Y(n4425));
  INVX1   g01439(.A(n4425), .Y(n4426));
  INVX1   g01440(.A(n4381), .Y(n4428));
  AOI21X1 g01441(.A0(n4428), .A1(n4426), .B0(n3989), .Y(n4429));
  NOR2X1  g01442(.A(n4429), .B(n4424), .Y(n4430));
  OAI21X1 g01443(.A0(n4269), .A1(n3509), .B0(n3994), .Y(n4432));
  NOR2X1  g01444(.A(n4432), .B(n4430), .Y(n4433));
  NOR4X1  g01445(.A(n4425), .B(n4074), .C(n3944), .D(n4381), .Y(n4434));
  OAI21X1 g01446(.A0(n4434), .A1(n3989), .B0(n4424), .Y(n4435));
  NOR3X1  g01447(.A(n4435), .B(n4007), .C(n3212), .Y(n4436));
  NOR4X1  g01448(.A(n4008), .B(n4007), .C(n3284), .D(n4426), .Y(n4437));
  OAI22X1 g01449(.A0(n4428), .A1(n4079), .B0(n4080), .B1(n4316), .Y(n4439));
  NOR3X1  g01450(.A(n4439), .B(n4437), .C(n4436), .Y(n4440));
  OAI21X1 g01451(.A0(n4433), .A1(n4422), .B0(n4440), .Y(P3_U2939));
  INVX1   g01452(.A(P3_INSTQUEUE_REG_8__6__SCAN_IN), .Y(n4442));
  NOR3X1  g01453(.A(n4435), .B(n4007), .C(n3209), .Y(n4443));
  NOR4X1  g01454(.A(n4008), .B(n4007), .C(n3281), .D(n4426), .Y(n4444));
  OAI22X1 g01455(.A0(n4428), .A1(n4088), .B0(n4089), .B1(n4316), .Y(n4445));
  NOR3X1  g01456(.A(n4445), .B(n4444), .C(n4443), .Y(n4446));
  OAI21X1 g01457(.A0(n4433), .A1(n4442), .B0(n4446), .Y(P3_U2938));
  INVX1   g01458(.A(P3_INSTQUEUE_REG_8__5__SCAN_IN), .Y(n4448));
  NOR3X1  g01459(.A(n4435), .B(n4007), .C(n3206), .Y(n4449));
  NOR4X1  g01460(.A(n4008), .B(n4007), .C(n3278), .D(n4426), .Y(n4450));
  OAI22X1 g01461(.A0(n4428), .A1(n4096), .B0(n4097), .B1(n4316), .Y(n4451));
  NOR3X1  g01462(.A(n4451), .B(n4450), .C(n4449), .Y(n4452));
  OAI21X1 g01463(.A0(n4433), .A1(n4448), .B0(n4452), .Y(P3_U2937));
  INVX1   g01464(.A(P3_INSTQUEUE_REG_8__4__SCAN_IN), .Y(n4454));
  NOR3X1  g01465(.A(n4435), .B(n4007), .C(n3203), .Y(n4455));
  NOR4X1  g01466(.A(n4008), .B(n4007), .C(n3275), .D(n4426), .Y(n4456));
  OAI22X1 g01467(.A0(n4428), .A1(n4104), .B0(n4105), .B1(n4316), .Y(n4457));
  NOR3X1  g01468(.A(n4457), .B(n4456), .C(n4455), .Y(n4458));
  OAI21X1 g01469(.A0(n4433), .A1(n4454), .B0(n4458), .Y(P3_U2936));
  INVX1   g01470(.A(P3_INSTQUEUE_REG_8__3__SCAN_IN), .Y(n4460));
  NOR3X1  g01471(.A(n4435), .B(n4007), .C(n3200), .Y(n4461));
  NOR4X1  g01472(.A(n4008), .B(n4007), .C(n3272), .D(n4426), .Y(n4462));
  OAI22X1 g01473(.A0(n4428), .A1(n4112), .B0(n4113), .B1(n4316), .Y(n4463));
  NOR3X1  g01474(.A(n4463), .B(n4462), .C(n4461), .Y(n4464));
  OAI21X1 g01475(.A0(n4433), .A1(n4460), .B0(n4464), .Y(P3_U2935));
  INVX1   g01476(.A(P3_INSTQUEUE_REG_8__2__SCAN_IN), .Y(n4466));
  NOR3X1  g01477(.A(n4435), .B(n4007), .C(n3197), .Y(n4467));
  NOR4X1  g01478(.A(n4008), .B(n4007), .C(n3269), .D(n4426), .Y(n4468));
  OAI22X1 g01479(.A0(n4428), .A1(n4120), .B0(n4121), .B1(n4316), .Y(n4469));
  NOR3X1  g01480(.A(n4469), .B(n4468), .C(n4467), .Y(n4470));
  OAI21X1 g01481(.A0(n4433), .A1(n4466), .B0(n4470), .Y(P3_U2934));
  INVX1   g01482(.A(P3_INSTQUEUE_REG_8__1__SCAN_IN), .Y(n4472));
  NOR3X1  g01483(.A(n4435), .B(n4007), .C(n3194), .Y(n4473));
  NOR4X1  g01484(.A(n4008), .B(n4007), .C(n3266), .D(n4426), .Y(n4474));
  OAI22X1 g01485(.A0(n4428), .A1(n4128), .B0(n4129), .B1(n4316), .Y(n4475));
  NOR3X1  g01486(.A(n4475), .B(n4474), .C(n4473), .Y(n4476));
  OAI21X1 g01487(.A0(n4433), .A1(n4472), .B0(n4476), .Y(P3_U2933));
  INVX1   g01488(.A(P3_INSTQUEUE_REG_8__0__SCAN_IN), .Y(n4478));
  NOR3X1  g01489(.A(n4435), .B(n4007), .C(n3190), .Y(n4479));
  NOR4X1  g01490(.A(n4008), .B(n4007), .C(n3263), .D(n4426), .Y(n4480));
  OAI22X1 g01491(.A0(n4428), .A1(n4136), .B0(n4137), .B1(n4316), .Y(n4481));
  NOR3X1  g01492(.A(n4481), .B(n4480), .C(n4479), .Y(n4482));
  OAI21X1 g01493(.A0(n4433), .A1(n4478), .B0(n4482), .Y(P3_U2932));
  NAND3X1 g01494(.A(n3518), .B(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C(n3513), .Y(n4485));
  OAI21X1 g01495(.A0(n4485), .A1(n3989), .B0(n4372), .Y(n4486));
  OAI21X1 g01496(.A0(n3995), .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B0(P3_STATE2_REG_3__SCAN_IN), .Y(n4487));
  NAND3X1 g01497(.A(n4487), .B(n4486), .C(n3994), .Y(n4488));
  NAND2X1 g01498(.A(n4488), .B(P3_INSTQUEUE_REG_7__7__SCAN_IN), .Y(n4489));
  NAND2X1 g01499(.A(n4485), .B(n3999), .Y(n4490));
  AOI21X1 g01500(.A0(n4490), .A1(n3988), .B0(n4372), .Y(n4491));
  NAND3X1 g01501(.A(n4491), .B(n3994), .C(BUF2_REG_7__SCAN_IN), .Y(n4492));
  NOR4X1  g01502(.A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n3516), .C(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .D(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Y(n4493));
  NAND4X1 g01503(.A(n3999), .B(n3994), .C(BUF2_REG_31__SCAN_IN), .D(n4493), .Y(n4494));
  AOI22X1 g01504(.A0(n4009), .A1(n4425), .B0(n4313), .B1(n4010), .Y(n4497));
  NAND4X1 g01505(.A(n4494), .B(n4492), .C(n4489), .D(n4497), .Y(P3_U2931));
  NAND2X1 g01506(.A(n4488), .B(P3_INSTQUEUE_REG_7__6__SCAN_IN), .Y(n4499));
  NAND3X1 g01507(.A(n4491), .B(n3994), .C(BUF2_REG_6__SCAN_IN), .Y(n4500));
  NAND4X1 g01508(.A(n3999), .B(n3994), .C(BUF2_REG_30__SCAN_IN), .D(n4493), .Y(n4501));
  AOI22X1 g01509(.A0(n4016), .A1(n4425), .B0(n4313), .B1(n4017), .Y(n4502));
  NAND4X1 g01510(.A(n4501), .B(n4500), .C(n4499), .D(n4502), .Y(P3_U2930));
  NAND2X1 g01511(.A(n4488), .B(P3_INSTQUEUE_REG_7__5__SCAN_IN), .Y(n4504));
  NAND3X1 g01512(.A(n4491), .B(n3994), .C(BUF2_REG_5__SCAN_IN), .Y(n4505));
  NAND4X1 g01513(.A(n3999), .B(n3994), .C(BUF2_REG_29__SCAN_IN), .D(n4493), .Y(n4506));
  AOI22X1 g01514(.A0(n4023), .A1(n4425), .B0(n4313), .B1(n4024), .Y(n4507));
  NAND4X1 g01515(.A(n4506), .B(n4505), .C(n4504), .D(n4507), .Y(P3_U2929));
  NAND2X1 g01516(.A(n4488), .B(P3_INSTQUEUE_REG_7__4__SCAN_IN), .Y(n4509));
  NAND3X1 g01517(.A(n4491), .B(n3994), .C(BUF2_REG_4__SCAN_IN), .Y(n4510));
  NAND4X1 g01518(.A(n3999), .B(n3994), .C(BUF2_REG_28__SCAN_IN), .D(n4493), .Y(n4511));
  AOI22X1 g01519(.A0(n4030), .A1(n4425), .B0(n4313), .B1(n4031), .Y(n4512));
  NAND4X1 g01520(.A(n4511), .B(n4510), .C(n4509), .D(n4512), .Y(P3_U2928));
  NAND2X1 g01521(.A(n4488), .B(P3_INSTQUEUE_REG_7__3__SCAN_IN), .Y(n4514));
  NAND3X1 g01522(.A(n4491), .B(n3994), .C(BUF2_REG_3__SCAN_IN), .Y(n4515));
  NAND4X1 g01523(.A(n3999), .B(n3994), .C(BUF2_REG_27__SCAN_IN), .D(n4493), .Y(n4516));
  AOI22X1 g01524(.A0(n4037), .A1(n4425), .B0(n4313), .B1(n4038), .Y(n4517));
  NAND4X1 g01525(.A(n4516), .B(n4515), .C(n4514), .D(n4517), .Y(P3_U2927));
  NAND2X1 g01526(.A(n4488), .B(P3_INSTQUEUE_REG_7__2__SCAN_IN), .Y(n4519));
  NAND3X1 g01527(.A(n4491), .B(n3994), .C(BUF2_REG_2__SCAN_IN), .Y(n4520));
  NAND4X1 g01528(.A(n3999), .B(n3994), .C(BUF2_REG_26__SCAN_IN), .D(n4493), .Y(n4521));
  AOI22X1 g01529(.A0(n4044), .A1(n4425), .B0(n4313), .B1(n4045), .Y(n4522));
  NAND4X1 g01530(.A(n4521), .B(n4520), .C(n4519), .D(n4522), .Y(P3_U2926));
  NAND2X1 g01531(.A(n4488), .B(P3_INSTQUEUE_REG_7__1__SCAN_IN), .Y(n4524));
  NAND3X1 g01532(.A(n4491), .B(n3994), .C(BUF2_REG_1__SCAN_IN), .Y(n4525));
  NAND4X1 g01533(.A(n3999), .B(n3994), .C(BUF2_REG_25__SCAN_IN), .D(n4493), .Y(n4526));
  AOI22X1 g01534(.A0(n4051), .A1(n4425), .B0(n4313), .B1(n4052), .Y(n4527));
  NAND4X1 g01535(.A(n4526), .B(n4525), .C(n4524), .D(n4527), .Y(P3_U2925));
  NAND2X1 g01536(.A(n4488), .B(P3_INSTQUEUE_REG_7__0__SCAN_IN), .Y(n4529));
  NAND3X1 g01537(.A(n4491), .B(n3994), .C(BUF2_REG_0__SCAN_IN), .Y(n4530));
  NAND4X1 g01538(.A(n3999), .B(n3994), .C(BUF2_REG_24__SCAN_IN), .D(n4493), .Y(n4531));
  AOI22X1 g01539(.A0(n4058), .A1(n4425), .B0(n4313), .B1(n4059), .Y(n4532));
  NAND4X1 g01540(.A(n4531), .B(n4530), .C(n4529), .D(n4532), .Y(P3_U2924));
  INVX1   g01541(.A(P3_INSTQUEUE_REG_6__7__SCAN_IN), .Y(n4534));
  NOR4X1  g01542(.A(n3518), .B(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .D(n3519), .Y(n4537));
  INVX1   g01543(.A(n4537), .Y(n4538));
  INVX1   g01544(.A(n4493), .Y(n4540));
  AOI21X1 g01545(.A0(n4540), .A1(n4538), .B0(n3989), .Y(n4541));
  NOR3X1  g01546(.A(n4541), .B(n4425), .C(n4381), .Y(n4542));
  OAI21X1 g01547(.A0(n4381), .A1(n3509), .B0(n3994), .Y(n4543));
  NOR2X1  g01548(.A(n4543), .B(n4542), .Y(n4544));
  NOR4X1  g01549(.A(n4537), .B(n4074), .C(n3944), .D(n4493), .Y(n4545));
  OAI22X1 g01550(.A0(n4425), .A1(n4381), .B0(n3989), .B1(n4545), .Y(n4546));
  NOR3X1  g01551(.A(n4546), .B(n4007), .C(n3212), .Y(n4547));
  NOR4X1  g01552(.A(n4008), .B(n4007), .C(n3284), .D(n4538), .Y(n4548));
  OAI22X1 g01553(.A0(n4428), .A1(n4080), .B0(n4079), .B1(n4540), .Y(n4550));
  NOR3X1  g01554(.A(n4550), .B(n4548), .C(n4547), .Y(n4551));
  OAI21X1 g01555(.A0(n4544), .A1(n4534), .B0(n4551), .Y(P3_U2923));
  INVX1   g01556(.A(P3_INSTQUEUE_REG_6__6__SCAN_IN), .Y(n4553));
  NOR3X1  g01557(.A(n4546), .B(n4007), .C(n3209), .Y(n4554));
  NOR4X1  g01558(.A(n4008), .B(n4007), .C(n3281), .D(n4538), .Y(n4555));
  OAI22X1 g01559(.A0(n4428), .A1(n4089), .B0(n4088), .B1(n4540), .Y(n4556));
  NOR3X1  g01560(.A(n4556), .B(n4555), .C(n4554), .Y(n4557));
  OAI21X1 g01561(.A0(n4544), .A1(n4553), .B0(n4557), .Y(P3_U2922));
  INVX1   g01562(.A(P3_INSTQUEUE_REG_6__5__SCAN_IN), .Y(n4559));
  NOR3X1  g01563(.A(n4546), .B(n4007), .C(n3206), .Y(n4560));
  NOR4X1  g01564(.A(n4008), .B(n4007), .C(n3278), .D(n4538), .Y(n4561));
  OAI22X1 g01565(.A0(n4428), .A1(n4097), .B0(n4096), .B1(n4540), .Y(n4562));
  NOR3X1  g01566(.A(n4562), .B(n4561), .C(n4560), .Y(n4563));
  OAI21X1 g01567(.A0(n4544), .A1(n4559), .B0(n4563), .Y(P3_U2921));
  INVX1   g01568(.A(P3_INSTQUEUE_REG_6__4__SCAN_IN), .Y(n4565));
  NOR3X1  g01569(.A(n4546), .B(n4007), .C(n3203), .Y(n4566));
  NOR4X1  g01570(.A(n4008), .B(n4007), .C(n3275), .D(n4538), .Y(n4567));
  OAI22X1 g01571(.A0(n4428), .A1(n4105), .B0(n4104), .B1(n4540), .Y(n4568));
  NOR3X1  g01572(.A(n4568), .B(n4567), .C(n4566), .Y(n4569));
  OAI21X1 g01573(.A0(n4544), .A1(n4565), .B0(n4569), .Y(P3_U2920));
  INVX1   g01574(.A(P3_INSTQUEUE_REG_6__3__SCAN_IN), .Y(n4571));
  NOR3X1  g01575(.A(n4546), .B(n4007), .C(n3200), .Y(n4572));
  NOR4X1  g01576(.A(n4008), .B(n4007), .C(n3272), .D(n4538), .Y(n4573));
  OAI22X1 g01577(.A0(n4428), .A1(n4113), .B0(n4112), .B1(n4540), .Y(n4574));
  NOR3X1  g01578(.A(n4574), .B(n4573), .C(n4572), .Y(n4575));
  OAI21X1 g01579(.A0(n4544), .A1(n4571), .B0(n4575), .Y(P3_U2919));
  INVX1   g01580(.A(P3_INSTQUEUE_REG_6__2__SCAN_IN), .Y(n4577));
  NOR3X1  g01581(.A(n4546), .B(n4007), .C(n3197), .Y(n4578));
  NOR4X1  g01582(.A(n4008), .B(n4007), .C(n3269), .D(n4538), .Y(n4579));
  OAI22X1 g01583(.A0(n4428), .A1(n4121), .B0(n4120), .B1(n4540), .Y(n4580));
  NOR3X1  g01584(.A(n4580), .B(n4579), .C(n4578), .Y(n4581));
  OAI21X1 g01585(.A0(n4544), .A1(n4577), .B0(n4581), .Y(P3_U2918));
  INVX1   g01586(.A(P3_INSTQUEUE_REG_6__1__SCAN_IN), .Y(n4583));
  NOR3X1  g01587(.A(n4546), .B(n4007), .C(n3194), .Y(n4584));
  NOR4X1  g01588(.A(n4008), .B(n4007), .C(n3266), .D(n4538), .Y(n4585));
  OAI22X1 g01589(.A0(n4428), .A1(n4129), .B0(n4128), .B1(n4540), .Y(n4586));
  NOR3X1  g01590(.A(n4586), .B(n4585), .C(n4584), .Y(n4587));
  OAI21X1 g01591(.A0(n4544), .A1(n4583), .B0(n4587), .Y(P3_U2917));
  INVX1   g01592(.A(P3_INSTQUEUE_REG_6__0__SCAN_IN), .Y(n4589));
  NOR3X1  g01593(.A(n4546), .B(n4007), .C(n3190), .Y(n4590));
  NOR4X1  g01594(.A(n4008), .B(n4007), .C(n3263), .D(n4538), .Y(n4591));
  OAI22X1 g01595(.A0(n4428), .A1(n4137), .B0(n4136), .B1(n4540), .Y(n4592));
  NOR3X1  g01596(.A(n4592), .B(n4591), .C(n4590), .Y(n4593));
  OAI21X1 g01597(.A0(n4544), .A1(n4589), .B0(n4593), .Y(P3_U2916));
  NAND3X1 g01598(.A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n3516), .C(n3513), .Y(n4596));
  OAI21X1 g01599(.A0(n4596), .A1(n3989), .B0(n4485), .Y(n4597));
  NAND2X1 g01600(.A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n3513), .Y(n4598));
  OAI21X1 g01601(.A0(n4598), .A1(n4144), .B0(P3_STATE2_REG_3__SCAN_IN), .Y(n4599));
  NAND3X1 g01602(.A(n4599), .B(n4597), .C(n3994), .Y(n4600));
  NAND2X1 g01603(.A(n4600), .B(P3_INSTQUEUE_REG_5__7__SCAN_IN), .Y(n4601));
  NAND2X1 g01604(.A(n4596), .B(n3999), .Y(n4602));
  AOI21X1 g01605(.A0(n4602), .A1(n3988), .B0(n4485), .Y(n4603));
  NAND3X1 g01606(.A(n4603), .B(n3994), .C(BUF2_REG_7__SCAN_IN), .Y(n4604));
  NOR4X1  g01607(.A(n3518), .B(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .D(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Y(n4605));
  NAND4X1 g01608(.A(n3999), .B(n3994), .C(BUF2_REG_31__SCAN_IN), .D(n4605), .Y(n4606));
  AOI22X1 g01609(.A0(n4425), .A1(n4010), .B0(n4009), .B1(n4537), .Y(n4609));
  NAND4X1 g01610(.A(n4606), .B(n4604), .C(n4601), .D(n4609), .Y(P3_U2915));
  NAND2X1 g01611(.A(n4600), .B(P3_INSTQUEUE_REG_5__6__SCAN_IN), .Y(n4611));
  NAND3X1 g01612(.A(n4603), .B(n3994), .C(BUF2_REG_6__SCAN_IN), .Y(n4612));
  NAND4X1 g01613(.A(n3999), .B(n3994), .C(BUF2_REG_30__SCAN_IN), .D(n4605), .Y(n4613));
  AOI22X1 g01614(.A0(n4425), .A1(n4017), .B0(n4016), .B1(n4537), .Y(n4614));
  NAND4X1 g01615(.A(n4613), .B(n4612), .C(n4611), .D(n4614), .Y(P3_U2914));
  NAND2X1 g01616(.A(n4600), .B(P3_INSTQUEUE_REG_5__5__SCAN_IN), .Y(n4616));
  NAND3X1 g01617(.A(n4603), .B(n3994), .C(BUF2_REG_5__SCAN_IN), .Y(n4617));
  NAND4X1 g01618(.A(n3999), .B(n3994), .C(BUF2_REG_29__SCAN_IN), .D(n4605), .Y(n4618));
  AOI22X1 g01619(.A0(n4425), .A1(n4024), .B0(n4023), .B1(n4537), .Y(n4619));
  NAND4X1 g01620(.A(n4618), .B(n4617), .C(n4616), .D(n4619), .Y(P3_U2913));
  NAND2X1 g01621(.A(n4600), .B(P3_INSTQUEUE_REG_5__4__SCAN_IN), .Y(n4621));
  NAND3X1 g01622(.A(n4603), .B(n3994), .C(BUF2_REG_4__SCAN_IN), .Y(n4622));
  NAND4X1 g01623(.A(n3999), .B(n3994), .C(BUF2_REG_28__SCAN_IN), .D(n4605), .Y(n4623));
  AOI22X1 g01624(.A0(n4425), .A1(n4031), .B0(n4030), .B1(n4537), .Y(n4624));
  NAND4X1 g01625(.A(n4623), .B(n4622), .C(n4621), .D(n4624), .Y(P3_U2912));
  NAND2X1 g01626(.A(n4600), .B(P3_INSTQUEUE_REG_5__3__SCAN_IN), .Y(n4626));
  NAND3X1 g01627(.A(n4603), .B(n3994), .C(BUF2_REG_3__SCAN_IN), .Y(n4627));
  NAND4X1 g01628(.A(n3999), .B(n3994), .C(BUF2_REG_27__SCAN_IN), .D(n4605), .Y(n4628));
  AOI22X1 g01629(.A0(n4425), .A1(n4038), .B0(n4037), .B1(n4537), .Y(n4629));
  NAND4X1 g01630(.A(n4628), .B(n4627), .C(n4626), .D(n4629), .Y(P3_U2911));
  NAND2X1 g01631(.A(n4600), .B(P3_INSTQUEUE_REG_5__2__SCAN_IN), .Y(n4631));
  NAND3X1 g01632(.A(n4603), .B(n3994), .C(BUF2_REG_2__SCAN_IN), .Y(n4632));
  NAND4X1 g01633(.A(n3999), .B(n3994), .C(BUF2_REG_26__SCAN_IN), .D(n4605), .Y(n4633));
  AOI22X1 g01634(.A0(n4425), .A1(n4045), .B0(n4044), .B1(n4537), .Y(n4634));
  NAND4X1 g01635(.A(n4633), .B(n4632), .C(n4631), .D(n4634), .Y(P3_U2910));
  NAND2X1 g01636(.A(n4600), .B(P3_INSTQUEUE_REG_5__1__SCAN_IN), .Y(n4636));
  NAND3X1 g01637(.A(n4603), .B(n3994), .C(BUF2_REG_1__SCAN_IN), .Y(n4637));
  NAND4X1 g01638(.A(n3999), .B(n3994), .C(BUF2_REG_25__SCAN_IN), .D(n4605), .Y(n4638));
  AOI22X1 g01639(.A0(n4425), .A1(n4052), .B0(n4051), .B1(n4537), .Y(n4639));
  NAND4X1 g01640(.A(n4638), .B(n4637), .C(n4636), .D(n4639), .Y(P3_U2909));
  NAND2X1 g01641(.A(n4600), .B(P3_INSTQUEUE_REG_5__0__SCAN_IN), .Y(n4641));
  NAND3X1 g01642(.A(n4603), .B(n3994), .C(BUF2_REG_0__SCAN_IN), .Y(n4642));
  NAND4X1 g01643(.A(n3999), .B(n3994), .C(BUF2_REG_24__SCAN_IN), .D(n4605), .Y(n4643));
  AOI22X1 g01644(.A0(n4425), .A1(n4059), .B0(n4058), .B1(n4537), .Y(n4644));
  NAND4X1 g01645(.A(n4643), .B(n4642), .C(n4641), .D(n4644), .Y(P3_U2908));
  NAND3X1 g01646(.A(n4197), .B(n4196), .C(n4423), .Y(n4646));
  NOR4X1  g01647(.A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .D(n3519), .Y(n4648));
  OAI21X1 g01648(.A0(n4648), .A1(n4605), .B0(n3988), .Y(n4649));
  NAND2X1 g01649(.A(n4649), .B(n4646), .Y(n4650));
  NAND2X1 g01650(.A(n4540), .B(P3_STATE2_REG_3__SCAN_IN), .Y(n4653));
  NAND3X1 g01651(.A(n4653), .B(n4650), .C(n3994), .Y(n4654));
  NAND2X1 g01652(.A(n4654), .B(P3_INSTQUEUE_REG_4__7__SCAN_IN), .Y(n4655));
  NAND4X1 g01653(.A(n3999), .B(n3994), .C(BUF2_REG_31__SCAN_IN), .D(n4648), .Y(n4656));
  NAND2X1 g01654(.A(n4493), .B(n4010), .Y(n4657));
  NOR2X1  g01655(.A(n4007), .B(n3212), .Y(n4658));
  INVX1   g01656(.A(n4196), .Y(n4659));
  NOR2X1  g01657(.A(P3_STATE2_REG_2__SCAN_IN), .B(n3509), .Y(n4660));
  NOR4X1  g01658(.A(n4957), .B(n4659), .C(n4195), .D(n4660), .Y(n4661));
  AOI22X1 g01659(.A0(n4605), .A1(n4009), .B0(n4658), .B1(n4661), .Y(n4662));
  NAND4X1 g01660(.A(n4657), .B(n4656), .C(n4655), .D(n4662), .Y(P3_U2907));
  NAND2X1 g01661(.A(n4654), .B(P3_INSTQUEUE_REG_4__6__SCAN_IN), .Y(n4664));
  NAND4X1 g01662(.A(n3999), .B(n3994), .C(BUF2_REG_30__SCAN_IN), .D(n4648), .Y(n4665));
  NAND2X1 g01663(.A(n4493), .B(n4017), .Y(n4666));
  NOR2X1  g01664(.A(n4007), .B(n3209), .Y(n4667));
  AOI22X1 g01665(.A0(n4605), .A1(n4016), .B0(n4667), .B1(n4661), .Y(n4668));
  NAND4X1 g01666(.A(n4666), .B(n4665), .C(n4664), .D(n4668), .Y(P3_U2906));
  NAND2X1 g01667(.A(n4654), .B(P3_INSTQUEUE_REG_4__5__SCAN_IN), .Y(n4670));
  NAND4X1 g01668(.A(n3999), .B(n3994), .C(BUF2_REG_29__SCAN_IN), .D(n4648), .Y(n4671));
  NAND2X1 g01669(.A(n4493), .B(n4024), .Y(n4672));
  NOR2X1  g01670(.A(n4007), .B(n3206), .Y(n4673));
  AOI22X1 g01671(.A0(n4605), .A1(n4023), .B0(n4673), .B1(n4661), .Y(n4674));
  NAND4X1 g01672(.A(n4672), .B(n4671), .C(n4670), .D(n4674), .Y(P3_U2905));
  NAND2X1 g01673(.A(n4654), .B(P3_INSTQUEUE_REG_4__4__SCAN_IN), .Y(n4676));
  NAND4X1 g01674(.A(n3999), .B(n3994), .C(BUF2_REG_28__SCAN_IN), .D(n4648), .Y(n4677));
  NAND2X1 g01675(.A(n4493), .B(n4031), .Y(n4678));
  NOR2X1  g01676(.A(n4007), .B(n3203), .Y(n4679));
  AOI22X1 g01677(.A0(n4605), .A1(n4030), .B0(n4679), .B1(n4661), .Y(n4680));
  NAND4X1 g01678(.A(n4678), .B(n4677), .C(n4676), .D(n4680), .Y(P3_U2904));
  NAND2X1 g01679(.A(n4654), .B(P3_INSTQUEUE_REG_4__3__SCAN_IN), .Y(n4682));
  NAND4X1 g01680(.A(n3999), .B(n3994), .C(BUF2_REG_27__SCAN_IN), .D(n4648), .Y(n4683));
  NAND2X1 g01681(.A(n4493), .B(n4038), .Y(n4684));
  NOR2X1  g01682(.A(n4007), .B(n3200), .Y(n4685));
  AOI22X1 g01683(.A0(n4605), .A1(n4037), .B0(n4685), .B1(n4661), .Y(n4686));
  NAND4X1 g01684(.A(n4684), .B(n4683), .C(n4682), .D(n4686), .Y(P3_U2903));
  NAND2X1 g01685(.A(n4654), .B(P3_INSTQUEUE_REG_4__2__SCAN_IN), .Y(n4688));
  NAND4X1 g01686(.A(n3999), .B(n3994), .C(BUF2_REG_26__SCAN_IN), .D(n4648), .Y(n4689));
  NAND2X1 g01687(.A(n4493), .B(n4045), .Y(n4690));
  NOR2X1  g01688(.A(n4007), .B(n3197), .Y(n4691));
  AOI22X1 g01689(.A0(n4605), .A1(n4044), .B0(n4691), .B1(n4661), .Y(n4692));
  NAND4X1 g01690(.A(n4690), .B(n4689), .C(n4688), .D(n4692), .Y(P3_U2902));
  NAND2X1 g01691(.A(n4654), .B(P3_INSTQUEUE_REG_4__1__SCAN_IN), .Y(n4694));
  NAND4X1 g01692(.A(n3999), .B(n3994), .C(BUF2_REG_25__SCAN_IN), .D(n4648), .Y(n4695));
  NAND2X1 g01693(.A(n4493), .B(n4052), .Y(n4696));
  NOR2X1  g01694(.A(n4007), .B(n3194), .Y(n4697));
  AOI22X1 g01695(.A0(n4605), .A1(n4051), .B0(n4697), .B1(n4661), .Y(n4698));
  NAND4X1 g01696(.A(n4696), .B(n4695), .C(n4694), .D(n4698), .Y(P3_U2901));
  NAND2X1 g01697(.A(n4654), .B(P3_INSTQUEUE_REG_4__0__SCAN_IN), .Y(n4700));
  NAND4X1 g01698(.A(n3999), .B(n3994), .C(BUF2_REG_24__SCAN_IN), .D(n4648), .Y(n4701));
  NAND2X1 g01699(.A(n4493), .B(n4059), .Y(n4702));
  NOR2X1  g01700(.A(n4007), .B(n3190), .Y(n4703));
  AOI22X1 g01701(.A0(n4605), .A1(n4058), .B0(n4703), .B1(n4661), .Y(n4704));
  NAND4X1 g01702(.A(n4702), .B(n4701), .C(n4700), .D(n4704), .Y(P3_U2900));
  NOR4X1  g01703(.A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .D(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Y(n4708));
  OAI21X1 g01704(.A0(n4708), .A1(n4648), .B0(n3988), .Y(n4709));
  NAND2X1 g01705(.A(n4709), .B(n4596), .Y(n4710));
  NAND2X1 g01706(.A(n3516), .B(n3513), .Y(n4711));
  OAI21X1 g01707(.A0(n4711), .A1(n4194), .B0(P3_STATE2_REG_3__SCAN_IN), .Y(n4712));
  NAND3X1 g01708(.A(n4712), .B(n4710), .C(n3994), .Y(n4713));
  NAND2X1 g01709(.A(n4713), .B(P3_INSTQUEUE_REG_3__7__SCAN_IN), .Y(n4714));
  NAND4X1 g01710(.A(n3999), .B(n3994), .C(BUF2_REG_31__SCAN_IN), .D(n4708), .Y(n4715));
  NAND2X1 g01711(.A(n4537), .B(n4010), .Y(n4717));
  NOR2X1  g01712(.A(n4596), .B(n4660), .Y(n4718));
  AOI22X1 g01713(.A0(n4648), .A1(n4009), .B0(n4658), .B1(n4718), .Y(n4719));
  NAND4X1 g01714(.A(n4717), .B(n4715), .C(n4714), .D(n4719), .Y(P3_U2899));
  NAND2X1 g01715(.A(n4713), .B(P3_INSTQUEUE_REG_3__6__SCAN_IN), .Y(n4721));
  NAND4X1 g01716(.A(n3999), .B(n3994), .C(BUF2_REG_30__SCAN_IN), .D(n4708), .Y(n4722));
  NAND2X1 g01717(.A(n4537), .B(n4017), .Y(n4723));
  AOI22X1 g01718(.A0(n4648), .A1(n4016), .B0(n4667), .B1(n4718), .Y(n4724));
  NAND4X1 g01719(.A(n4723), .B(n4722), .C(n4721), .D(n4724), .Y(P3_U2898));
  NAND2X1 g01720(.A(n4713), .B(P3_INSTQUEUE_REG_3__5__SCAN_IN), .Y(n4726));
  NAND4X1 g01721(.A(n3999), .B(n3994), .C(BUF2_REG_29__SCAN_IN), .D(n4708), .Y(n4727));
  NAND2X1 g01722(.A(n4537), .B(n4024), .Y(n4728));
  AOI22X1 g01723(.A0(n4648), .A1(n4023), .B0(n4673), .B1(n4718), .Y(n4729));
  NAND4X1 g01724(.A(n4728), .B(n4727), .C(n4726), .D(n4729), .Y(P3_U2897));
  NAND2X1 g01725(.A(n4713), .B(P3_INSTQUEUE_REG_3__4__SCAN_IN), .Y(n4731));
  NAND4X1 g01726(.A(n3999), .B(n3994), .C(BUF2_REG_28__SCAN_IN), .D(n4708), .Y(n4732));
  NAND2X1 g01727(.A(n4537), .B(n4031), .Y(n4733));
  AOI22X1 g01728(.A0(n4648), .A1(n4030), .B0(n4679), .B1(n4718), .Y(n4734));
  NAND4X1 g01729(.A(n4733), .B(n4732), .C(n4731), .D(n4734), .Y(P3_U2896));
  NAND2X1 g01730(.A(n4713), .B(P3_INSTQUEUE_REG_3__3__SCAN_IN), .Y(n4736));
  NAND4X1 g01731(.A(n3999), .B(n3994), .C(BUF2_REG_27__SCAN_IN), .D(n4708), .Y(n4737));
  NAND2X1 g01732(.A(n4537), .B(n4038), .Y(n4738));
  AOI22X1 g01733(.A0(n4648), .A1(n4037), .B0(n4685), .B1(n4718), .Y(n4739));
  NAND4X1 g01734(.A(n4738), .B(n4737), .C(n4736), .D(n4739), .Y(P3_U2895));
  NAND2X1 g01735(.A(n4713), .B(P3_INSTQUEUE_REG_3__2__SCAN_IN), .Y(n4741));
  NAND4X1 g01736(.A(n3999), .B(n3994), .C(BUF2_REG_26__SCAN_IN), .D(n4708), .Y(n4742));
  NAND2X1 g01737(.A(n4537), .B(n4045), .Y(n4743));
  AOI22X1 g01738(.A0(n4648), .A1(n4044), .B0(n4691), .B1(n4718), .Y(n4744));
  NAND4X1 g01739(.A(n4743), .B(n4742), .C(n4741), .D(n4744), .Y(P3_U2894));
  NAND2X1 g01740(.A(n4713), .B(P3_INSTQUEUE_REG_3__1__SCAN_IN), .Y(n4746));
  NAND4X1 g01741(.A(n3999), .B(n3994), .C(BUF2_REG_25__SCAN_IN), .D(n4708), .Y(n4747));
  NAND2X1 g01742(.A(n4537), .B(n4052), .Y(n4748));
  AOI22X1 g01743(.A0(n4648), .A1(n4051), .B0(n4697), .B1(n4718), .Y(n4749));
  NAND4X1 g01744(.A(n4748), .B(n4747), .C(n4746), .D(n4749), .Y(P3_U2893));
  NAND2X1 g01745(.A(n4713), .B(P3_INSTQUEUE_REG_3__0__SCAN_IN), .Y(n4751));
  NAND4X1 g01746(.A(n3999), .B(n3994), .C(BUF2_REG_24__SCAN_IN), .D(n4708), .Y(n4752));
  NAND2X1 g01747(.A(n4537), .B(n4059), .Y(n4753));
  AOI22X1 g01748(.A0(n4648), .A1(n4058), .B0(n4703), .B1(n4718), .Y(n4754));
  NAND4X1 g01749(.A(n4753), .B(n4752), .C(n4751), .D(n4754), .Y(P3_U2892));
  INVX1   g01750(.A(n4605), .Y(n4757));
  NAND4X1 g01751(.A(n3518), .B(n3516), .C(n3513), .D(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Y(n4758));
  OAI21X1 g01752(.A0(n4005), .A1(n4708), .B0(n3988), .Y(n4761));
  NAND3X1 g01753(.A(n4761), .B(n4758), .C(n4757), .Y(n4762));
  NAND2X1 g01754(.A(n4757), .B(P3_STATE2_REG_3__SCAN_IN), .Y(n4763));
  NAND3X1 g01755(.A(n4763), .B(n4762), .C(n3994), .Y(n4764));
  NAND2X1 g01756(.A(n4764), .B(P3_INSTQUEUE_REG_2__7__SCAN_IN), .Y(n4765));
  NAND4X1 g01757(.A(n3999), .B(n3994), .C(BUF2_REG_31__SCAN_IN), .D(n4005), .Y(n4766));
  NAND2X1 g01758(.A(n4605), .B(n4010), .Y(n4767));
  AOI21X1 g01759(.A0(n4758), .A1(n4757), .B0(n4660), .Y(n4768));
  AOI22X1 g01760(.A0(n4708), .A1(n4009), .B0(n4658), .B1(n4768), .Y(n4769));
  NAND4X1 g01761(.A(n4767), .B(n4766), .C(n4765), .D(n4769), .Y(P3_U2891));
  NAND2X1 g01762(.A(n4764), .B(P3_INSTQUEUE_REG_2__6__SCAN_IN), .Y(n4771));
  NAND4X1 g01763(.A(n3999), .B(n3994), .C(BUF2_REG_30__SCAN_IN), .D(n4005), .Y(n4772));
  NAND2X1 g01764(.A(n4605), .B(n4017), .Y(n4773));
  AOI22X1 g01765(.A0(n4708), .A1(n4016), .B0(n4667), .B1(n4768), .Y(n4774));
  NAND4X1 g01766(.A(n4773), .B(n4772), .C(n4771), .D(n4774), .Y(P3_U2890));
  NAND2X1 g01767(.A(n4764), .B(P3_INSTQUEUE_REG_2__5__SCAN_IN), .Y(n4776));
  NAND4X1 g01768(.A(n3999), .B(n3994), .C(BUF2_REG_29__SCAN_IN), .D(n4005), .Y(n4777));
  NAND2X1 g01769(.A(n4605), .B(n4024), .Y(n4778));
  AOI22X1 g01770(.A0(n4708), .A1(n4023), .B0(n4673), .B1(n4768), .Y(n4779));
  NAND4X1 g01771(.A(n4778), .B(n4777), .C(n4776), .D(n4779), .Y(P3_U2889));
  NAND2X1 g01772(.A(n4764), .B(P3_INSTQUEUE_REG_2__4__SCAN_IN), .Y(n4781));
  NAND4X1 g01773(.A(n3999), .B(n3994), .C(BUF2_REG_28__SCAN_IN), .D(n4005), .Y(n4782));
  NAND2X1 g01774(.A(n4605), .B(n4031), .Y(n4783));
  AOI22X1 g01775(.A0(n4708), .A1(n4030), .B0(n4679), .B1(n4768), .Y(n4784));
  NAND4X1 g01776(.A(n4783), .B(n4782), .C(n4781), .D(n4784), .Y(P3_U2888));
  NAND2X1 g01777(.A(n4764), .B(P3_INSTQUEUE_REG_2__3__SCAN_IN), .Y(n4786));
  NAND4X1 g01778(.A(n3999), .B(n3994), .C(BUF2_REG_27__SCAN_IN), .D(n4005), .Y(n4787));
  NAND2X1 g01779(.A(n4605), .B(n4038), .Y(n4788));
  AOI22X1 g01780(.A0(n4708), .A1(n4037), .B0(n4685), .B1(n4768), .Y(n4789));
  NAND4X1 g01781(.A(n4788), .B(n4787), .C(n4786), .D(n4789), .Y(P3_U2887));
  NAND2X1 g01782(.A(n4764), .B(P3_INSTQUEUE_REG_2__2__SCAN_IN), .Y(n4791));
  NAND4X1 g01783(.A(n3999), .B(n3994), .C(BUF2_REG_26__SCAN_IN), .D(n4005), .Y(n4792));
  NAND2X1 g01784(.A(n4605), .B(n4045), .Y(n4793));
  AOI22X1 g01785(.A0(n4708), .A1(n4044), .B0(n4691), .B1(n4768), .Y(n4794));
  NAND4X1 g01786(.A(n4793), .B(n4792), .C(n4791), .D(n4794), .Y(P3_U2886));
  NAND2X1 g01787(.A(n4764), .B(P3_INSTQUEUE_REG_2__1__SCAN_IN), .Y(n4796));
  NAND4X1 g01788(.A(n3999), .B(n3994), .C(BUF2_REG_25__SCAN_IN), .D(n4005), .Y(n4797));
  NAND2X1 g01789(.A(n4605), .B(n4052), .Y(n4798));
  AOI22X1 g01790(.A0(n4708), .A1(n4051), .B0(n4697), .B1(n4768), .Y(n4799));
  NAND4X1 g01791(.A(n4798), .B(n4797), .C(n4796), .D(n4799), .Y(P3_U2885));
  NAND2X1 g01792(.A(n4764), .B(P3_INSTQUEUE_REG_2__0__SCAN_IN), .Y(n4801));
  NAND4X1 g01793(.A(n3999), .B(n3994), .C(BUF2_REG_24__SCAN_IN), .D(n4005), .Y(n4802));
  NAND2X1 g01794(.A(n4605), .B(n4059), .Y(n4803));
  AOI22X1 g01795(.A0(n4708), .A1(n4058), .B0(n4703), .B1(n4768), .Y(n4804));
  NAND4X1 g01796(.A(n4803), .B(n4802), .C(n4801), .D(n4804), .Y(P3_U2884));
  NAND3X1 g01797(.A(n3518), .B(n3516), .C(n3513), .Y(n4806));
  OAI21X1 g01798(.A0(n4063), .A1(n4005), .B0(n3988), .Y(n4809));
  NAND2X1 g01799(.A(n4809), .B(n4806), .Y(n4810));
  OAI21X1 g01800(.A0(n4711), .A1(n4144), .B0(P3_STATE2_REG_3__SCAN_IN), .Y(n4811));
  NAND3X1 g01801(.A(n4811), .B(n4810), .C(n3994), .Y(n4812));
  NAND2X1 g01802(.A(n4812), .B(P3_INSTQUEUE_REG_1__7__SCAN_IN), .Y(n4813));
  NAND4X1 g01803(.A(n3999), .B(n3994), .C(BUF2_REG_31__SCAN_IN), .D(n4063), .Y(n4814));
  NAND2X1 g01804(.A(n4648), .B(n4010), .Y(n4816));
  NOR2X1  g01805(.A(n4806), .B(n4660), .Y(n4817));
  AOI22X1 g01806(.A0(n4005), .A1(n4009), .B0(n4658), .B1(n4817), .Y(n4818));
  NAND4X1 g01807(.A(n4816), .B(n4814), .C(n4813), .D(n4818), .Y(P3_U2883));
  NAND2X1 g01808(.A(n4812), .B(P3_INSTQUEUE_REG_1__6__SCAN_IN), .Y(n4820));
  NAND4X1 g01809(.A(n3999), .B(n3994), .C(BUF2_REG_30__SCAN_IN), .D(n4063), .Y(n4821));
  NAND2X1 g01810(.A(n4648), .B(n4017), .Y(n4822));
  AOI22X1 g01811(.A0(n4005), .A1(n4016), .B0(n4667), .B1(n4817), .Y(n4823));
  NAND4X1 g01812(.A(n4822), .B(n4821), .C(n4820), .D(n4823), .Y(P3_U2882));
  NAND2X1 g01813(.A(n4812), .B(P3_INSTQUEUE_REG_1__5__SCAN_IN), .Y(n4825));
  NAND4X1 g01814(.A(n3999), .B(n3994), .C(BUF2_REG_29__SCAN_IN), .D(n4063), .Y(n4826));
  NAND2X1 g01815(.A(n4648), .B(n4024), .Y(n4827));
  AOI22X1 g01816(.A0(n4005), .A1(n4023), .B0(n4673), .B1(n4817), .Y(n4828));
  NAND4X1 g01817(.A(n4827), .B(n4826), .C(n4825), .D(n4828), .Y(P3_U2881));
  NAND2X1 g01818(.A(n4812), .B(P3_INSTQUEUE_REG_1__4__SCAN_IN), .Y(n4830));
  NAND4X1 g01819(.A(n3999), .B(n3994), .C(BUF2_REG_28__SCAN_IN), .D(n4063), .Y(n4831));
  NAND2X1 g01820(.A(n4648), .B(n4031), .Y(n4832));
  AOI22X1 g01821(.A0(n4005), .A1(n4030), .B0(n4679), .B1(n4817), .Y(n4833));
  NAND4X1 g01822(.A(n4832), .B(n4831), .C(n4830), .D(n4833), .Y(P3_U2880));
  NAND2X1 g01823(.A(n4812), .B(P3_INSTQUEUE_REG_1__3__SCAN_IN), .Y(n4835));
  NAND4X1 g01824(.A(n3999), .B(n3994), .C(BUF2_REG_27__SCAN_IN), .D(n4063), .Y(n4836));
  NAND2X1 g01825(.A(n4648), .B(n4038), .Y(n4837));
  AOI22X1 g01826(.A0(n4005), .A1(n4037), .B0(n4685), .B1(n4817), .Y(n4838));
  NAND4X1 g01827(.A(n4837), .B(n4836), .C(n4835), .D(n4838), .Y(P3_U2879));
  NAND2X1 g01828(.A(n4812), .B(P3_INSTQUEUE_REG_1__2__SCAN_IN), .Y(n4840));
  NAND4X1 g01829(.A(n3999), .B(n3994), .C(BUF2_REG_26__SCAN_IN), .D(n4063), .Y(n4841));
  NAND2X1 g01830(.A(n4648), .B(n4045), .Y(n4842));
  AOI22X1 g01831(.A0(n4005), .A1(n4044), .B0(n4691), .B1(n4817), .Y(n4843));
  NAND4X1 g01832(.A(n4842), .B(n4841), .C(n4840), .D(n4843), .Y(P3_U2878));
  NAND2X1 g01833(.A(n4812), .B(P3_INSTQUEUE_REG_1__1__SCAN_IN), .Y(n4845));
  NAND4X1 g01834(.A(n3999), .B(n3994), .C(BUF2_REG_25__SCAN_IN), .D(n4063), .Y(n4846));
  NAND2X1 g01835(.A(n4648), .B(n4052), .Y(n4847));
  AOI22X1 g01836(.A0(n4005), .A1(n4051), .B0(n4697), .B1(n4817), .Y(n4848));
  NAND4X1 g01837(.A(n4847), .B(n4846), .C(n4845), .D(n4848), .Y(P3_U2877));
  NAND2X1 g01838(.A(n4812), .B(P3_INSTQUEUE_REG_1__0__SCAN_IN), .Y(n4850));
  NAND4X1 g01839(.A(n3999), .B(n3994), .C(BUF2_REG_24__SCAN_IN), .D(n4063), .Y(n4851));
  NAND2X1 g01840(.A(n4648), .B(n4059), .Y(n4852));
  AOI22X1 g01841(.A0(n4005), .A1(n4058), .B0(n4703), .B1(n4817), .Y(n4853));
  NAND4X1 g01842(.A(n4852), .B(n4851), .C(n4850), .D(n4853), .Y(P3_U2876));
  NAND3X1 g01843(.A(n4197), .B(n4196), .C(n4195), .Y(n4855));
  OAI21X1 g01844(.A0(n4006), .A1(n4063), .B0(n3988), .Y(n4858));
  NAND2X1 g01845(.A(n4858), .B(n4855), .Y(n4859));
  INVX1   g01846(.A(n4708), .Y(n4861));
  NAND2X1 g01847(.A(n4861), .B(P3_STATE2_REG_3__SCAN_IN), .Y(n4862));
  NAND3X1 g01848(.A(n4862), .B(n4859), .C(n3994), .Y(n4863));
  NAND2X1 g01849(.A(n4863), .B(P3_INSTQUEUE_REG_0__7__SCAN_IN), .Y(n4864));
  NAND4X1 g01850(.A(n3999), .B(n3994), .C(BUF2_REG_31__SCAN_IN), .D(n4006), .Y(n4865));
  NAND2X1 g01851(.A(n4708), .B(n4010), .Y(n4866));
  NOR2X1  g01852(.A(n4855), .B(n4660), .Y(n4867));
  AOI22X1 g01853(.A0(n4063), .A1(n4009), .B0(n4658), .B1(n4867), .Y(n4868));
  NAND4X1 g01854(.A(n4866), .B(n4865), .C(n4864), .D(n4868), .Y(P3_U2875));
  NAND2X1 g01855(.A(n4863), .B(P3_INSTQUEUE_REG_0__6__SCAN_IN), .Y(n4870));
  NAND4X1 g01856(.A(n3999), .B(n3994), .C(BUF2_REG_30__SCAN_IN), .D(n4006), .Y(n4871));
  NAND2X1 g01857(.A(n4708), .B(n4017), .Y(n4872));
  AOI22X1 g01858(.A0(n4063), .A1(n4016), .B0(n4667), .B1(n4867), .Y(n4873));
  NAND4X1 g01859(.A(n4872), .B(n4871), .C(n4870), .D(n4873), .Y(P3_U2874));
  NAND2X1 g01860(.A(n4863), .B(P3_INSTQUEUE_REG_0__5__SCAN_IN), .Y(n4875));
  NAND4X1 g01861(.A(n3999), .B(n3994), .C(BUF2_REG_29__SCAN_IN), .D(n4006), .Y(n4876));
  NAND2X1 g01862(.A(n4708), .B(n4024), .Y(n4877));
  AOI22X1 g01863(.A0(n4063), .A1(n4023), .B0(n4673), .B1(n4867), .Y(n4878));
  NAND4X1 g01864(.A(n4877), .B(n4876), .C(n4875), .D(n4878), .Y(P3_U2873));
  NAND2X1 g01865(.A(n4863), .B(P3_INSTQUEUE_REG_0__4__SCAN_IN), .Y(n4880));
  NAND4X1 g01866(.A(n3999), .B(n3994), .C(BUF2_REG_28__SCAN_IN), .D(n4006), .Y(n4881));
  NAND2X1 g01867(.A(n4708), .B(n4031), .Y(n4882));
  AOI22X1 g01868(.A0(n4063), .A1(n4030), .B0(n4679), .B1(n4867), .Y(n4883));
  NAND4X1 g01869(.A(n4882), .B(n4881), .C(n4880), .D(n4883), .Y(P3_U2872));
  NAND2X1 g01870(.A(n4863), .B(P3_INSTQUEUE_REG_0__3__SCAN_IN), .Y(n4885));
  NAND4X1 g01871(.A(n3999), .B(n3994), .C(BUF2_REG_27__SCAN_IN), .D(n4006), .Y(n4886));
  NAND2X1 g01872(.A(n4708), .B(n4038), .Y(n4887));
  AOI22X1 g01873(.A0(n4063), .A1(n4037), .B0(n4685), .B1(n4867), .Y(n4888));
  NAND4X1 g01874(.A(n4887), .B(n4886), .C(n4885), .D(n4888), .Y(P3_U2871));
  NAND2X1 g01875(.A(n4863), .B(P3_INSTQUEUE_REG_0__2__SCAN_IN), .Y(n4890));
  NAND4X1 g01876(.A(n3999), .B(n3994), .C(BUF2_REG_26__SCAN_IN), .D(n4006), .Y(n4891));
  NAND2X1 g01877(.A(n4708), .B(n4045), .Y(n4892));
  AOI22X1 g01878(.A0(n4063), .A1(n4044), .B0(n4691), .B1(n4867), .Y(n4893));
  NAND4X1 g01879(.A(n4892), .B(n4891), .C(n4890), .D(n4893), .Y(P3_U2870));
  NAND2X1 g01880(.A(n4863), .B(P3_INSTQUEUE_REG_0__1__SCAN_IN), .Y(n4895));
  NAND4X1 g01881(.A(n3999), .B(n3994), .C(BUF2_REG_25__SCAN_IN), .D(n4006), .Y(n4896));
  NAND2X1 g01882(.A(n4708), .B(n4052), .Y(n4897));
  AOI22X1 g01883(.A0(n4063), .A1(n4051), .B0(n4697), .B1(n4867), .Y(n4898));
  NAND4X1 g01884(.A(n4897), .B(n4896), .C(n4895), .D(n4898), .Y(P3_U2869));
  NAND2X1 g01885(.A(n4863), .B(P3_INSTQUEUE_REG_0__0__SCAN_IN), .Y(n4900));
  NAND4X1 g01886(.A(n3999), .B(n3994), .C(BUF2_REG_24__SCAN_IN), .D(n4006), .Y(n4901));
  NAND2X1 g01887(.A(n4708), .B(n4059), .Y(n4902));
  AOI22X1 g01888(.A0(n4063), .A1(n4058), .B0(n4703), .B1(n4867), .Y(n4903));
  NAND4X1 g01889(.A(n4902), .B(n4901), .C(n4900), .D(n4903), .Y(P3_U2868));
  INVX1   g01890(.A(n3955), .Y(n4905));
  NOR4X1  g01891(.A(n3510), .B(n3939), .C(n3511), .D(n3959), .Y(n4906));
  AOI21X1 g01892(.A0(n3510), .A1(P3_STATE2_REG_3__SCAN_IN), .B0(n4906), .Y(n4907));
  OAI21X1 g01893(.A0(n4905), .A1(n3752), .B0(n4907), .Y(n4908));
  INVX1   g01894(.A(n3949), .Y(n4909));
  NOR3X1  g01895(.A(n4909), .B(n3755), .C(n3753), .Y(n4910));
  NAND2X1 g01896(.A(n4910), .B(n4908), .Y(n4911));
  OAI21X1 g01897(.A0(n4908), .A1(n3531), .B0(n4911), .Y(P3_U3284));
  INVX1   g01898(.A(n3980), .Y(n4913));
  NOR2X1  g01899(.A(n3867), .B(n3571), .Y(n4914));
  OAI22X1 g01900(.A0(n4913), .A1(n4914), .B0(n4909), .B1(n3878), .Y(n4915));
  NAND2X1 g01901(.A(n4915), .B(n4908), .Y(n4916));
  OAI21X1 g01902(.A0(n4908), .A1(n3535), .B0(n4916), .Y(P3_U3285));
  INVX1   g01903(.A(n4908), .Y(n4918));
  NOR2X1  g01904(.A(n3974), .B(n3960), .Y(n4919));
  NAND2X1 g01905(.A(n4919), .B(P3_STATE2_REG_1__SCAN_IN), .Y(n4920));
  OAI21X1 g01906(.A0(n4913), .A1(n3824), .B0(n4920), .Y(n4921));
  AOI21X1 g01907(.A0(n3949), .A1(n3830), .B0(n4921), .Y(n4922));
  NAND2X1 g01908(.A(n4918), .B(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Y(n4923));
  OAI21X1 g01909(.A0(n4922), .A1(n4918), .B0(n4923), .Y(P3_U3288));
  INVX1   g01910(.A(n3960), .Y(n4925));
  NAND3X1 g01911(.A(n3974), .B(n4925), .C(P3_STATE2_REG_1__SCAN_IN), .Y(n4926));
  OAI21X1 g01912(.A0(n4913), .A1(n3839), .B0(n4926), .Y(n4927));
  AOI21X1 g01913(.A0(n3949), .A1(n3842), .B0(n4927), .Y(n4928));
  NAND2X1 g01914(.A(n4918), .B(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Y(n4929));
  OAI21X1 g01915(.A0(n4928), .A1(n4918), .B0(n4929), .Y(P3_U3289));
  OAI22X1 g01916(.A0(n4925), .A1(n3939), .B0(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(n4913), .Y(n4931));
  AOI21X1 g01917(.A0(n3949), .A1(n3848), .B0(n4931), .Y(n4932));
  NAND2X1 g01918(.A(n4918), .B(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n4933));
  OAI21X1 g01919(.A0(n4932), .A1(n4918), .B0(n4933), .Y(P3_U3290));
  NAND3X1 g01920(.A(n3976), .B(n3940), .C(P3_STATE2_REG_0__SCAN_IN), .Y(n4935));
  INVX1   g01921(.A(n4935), .Y(n4936));
  NOR4X1  g01922(.A(n4906), .B(n3994), .C(n3512), .D(n4936), .Y(P3_U2867));
  NOR3X1  g01923(.A(n4936), .B(n4906), .C(n3994), .Y(n4938));
  AOI21X1 g01924(.A0(n3995), .A1(P3_STATE2_REG_3__SCAN_IN), .B0(n4938), .Y(n4939));
  XOR2X1  g01925(.A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .Y(n4940));
  NAND3X1 g01926(.A(n3519), .B(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .Y(n4942));
  AOI21X1 g01927(.A0(n4942), .A1(n4659), .B0(n4381), .Y(n4943));
  AOI21X1 g01928(.A0(n4073), .A1(n3944), .B0(n3949), .Y(n4944));
  NAND2X1 g01929(.A(n4313), .B(P3_STATE2_REG_3__SCAN_IN), .Y(n4945));
  OAI21X1 g01930(.A0(n4944), .A1(n4943), .B0(n4945), .Y(n4946));
  AOI21X1 g01931(.A0(n4940), .A1(n3999), .B0(n4946), .Y(n4947));
  OAI22X1 g01932(.A0(n4939), .A1(n3513), .B0(n4938), .B1(n4947), .Y(P3_U2866));
  XOR2X1  g01933(.A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n3516), .Y(n4952));
  OAI22X1 g01934(.A0(n4952), .A1(n4944), .B0(n4262), .B1(n3509), .Y(n4953));
  AOI21X1 g01935(.A0(n3516), .A1(n3999), .B0(n4953), .Y(n4954));
  AOI21X1 g01936(.A0(n4194), .A1(P3_STATE2_REG_3__SCAN_IN), .B0(n4938), .Y(n4955));
  OAI22X1 g01937(.A0(n4954), .A1(n4938), .B0(n3516), .B1(n4955), .Y(P3_U2865));
  XOR2X1  g01938(.A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Y(n4957));
  OAI22X1 g01939(.A0(n4957), .A1(n4008), .B0(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(n3509), .Y(n4958));
  XOR2X1  g01940(.A(n4197), .B(n3519), .Y(n4959));
  NAND4X1 g01941(.A(P3_STATEBS16_REG_SCAN_IN), .B(n3519), .C(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .D(n4073), .Y(n4960));
  OAI21X1 g01942(.A0(n4944), .A1(n4959), .B0(n4960), .Y(n4961));
  AOI21X1 g01943(.A0(n4958), .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B0(n4961), .Y(n4962));
  AOI21X1 g01944(.A0(n3519), .A1(P3_STATE2_REG_3__SCAN_IN), .B0(n4938), .Y(n4963));
  OAI22X1 g01945(.A0(n4962), .A1(n4938), .B0(n3518), .B1(n4963), .Y(P3_U2864));
  NOR3X1  g01946(.A(n4938), .B(n4073), .C(n3949), .Y(n4965));
  AOI21X1 g01947(.A0(n3519), .A1(P3_STATE2_REG_3__SCAN_IN), .B0(n3977), .Y(n4966));
  OAI22X1 g01948(.A0(n4965), .A1(n3519), .B0(n4938), .B1(n4966), .Y(P3_U2863));
  NOR4X1  g01949(.A(P3_STATE2_REG_1__SCAN_IN), .B(P3_STATE2_REG_2__SCAN_IN), .C(P3_STATE2_REG_3__SCAN_IN), .D(P3_STATE2_REG_0__SCAN_IN), .Y(n4968));
  INVX1   g01950(.A(n4968), .Y(n4969));
  NOR4X1  g01951(.A(n3715), .B(n3714), .C(n3407), .D(n3726), .Y(n4970));
  AOI22X1 g01952(.A0(n3893), .A1(n3709), .B0(n3705), .B1(n4970), .Y(n4971));
  NAND3X1 g01953(.A(n3705), .B(n3650), .C(n3408), .Y(n4972));
  OAI21X1 g01954(.A0(n3891), .A1(n3708), .B0(n4972), .Y(n4973));
  AOI22X1 g01955(.A0(n3698), .A1(n3893), .B0(n3682), .B1(n4973), .Y(n4974));
  OAI21X1 g01956(.A0(n4971), .A1(n3682), .B0(n4974), .Y(n4975));
  INVX1   g01957(.A(n3744), .Y(n4976));
  AOI22X1 g01958(.A0(n3747), .A1(n3667), .B0(n3705), .B1(n3909), .Y(n4977));
  NOR4X1  g01959(.A(n3634), .B(n3547), .C(n3529), .D(n3698), .Y(n4978));
  AOI21X1 g01960(.A0(n3905), .A1(n3705), .B0(n4978), .Y(n4979));
  NAND3X1 g01961(.A(n4979), .B(n4977), .C(n4976), .Y(n4980));
  AOI21X1 g01962(.A0(n4975), .A1(n3583), .B0(n4980), .Y(n4981));
  OAI21X1 g01963(.A0(n4981), .A1(n4905), .B0(n4969), .Y(n4982));
  INVX1   g01964(.A(n4982), .Y(n4983));
  NOR2X1  g01965(.A(n4983), .B(n3511), .Y(n4984));
  INVX1   g01966(.A(n4984), .Y(n4985));
  AOI22X1 g01967(.A0(n3577), .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B0(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(n3550), .Y(n4988));
  AOI22X1 g01968(.A0(n3574), .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B0(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3562), .Y(n4991));
  AOI22X1 g01969(.A0(n3555), .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B0(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3575), .Y(n4994));
  AOI22X1 g01970(.A0(n3572), .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B0(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3568), .Y(n4997));
  NAND4X1 g01971(.A(n4994), .B(n4991), .C(n4988), .D(n4997), .Y(n4998));
  AOI22X1 g01972(.A0(n3565), .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B0(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3563), .Y(n5001));
  AOI22X1 g01973(.A0(n3578), .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B0(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3569), .Y(n5004));
  AOI22X1 g01974(.A0(n3571), .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B0(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3560), .Y(n5007));
  AOI22X1 g01975(.A0(n3566), .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B0(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3557), .Y(n5010));
  NAND4X1 g01976(.A(n5007), .B(n5004), .C(n5001), .D(n5010), .Y(n5011));
  NOR2X1  g01977(.A(n5011), .B(n4998), .Y(n5012));
  XOR2X1  g01978(.A(n5012), .B(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .Y(n5013));
  INVX1   g01979(.A(n5013), .Y(n5014));
  AOI22X1 g01980(.A0(n3577), .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B0(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3550), .Y(n5015));
  AOI22X1 g01981(.A0(n3574), .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B0(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3562), .Y(n5016));
  AOI22X1 g01982(.A0(n3555), .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B0(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3575), .Y(n5017));
  AOI22X1 g01983(.A0(n3572), .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B0(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3568), .Y(n5018));
  NAND4X1 g01984(.A(n5017), .B(n5016), .C(n5015), .D(n5018), .Y(n5019));
  AOI22X1 g01985(.A0(n3565), .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B0(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3563), .Y(n5020));
  AOI22X1 g01986(.A0(n3578), .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B0(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3569), .Y(n5021));
  AOI22X1 g01987(.A0(n3571), .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B0(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3560), .Y(n5022));
  AOI22X1 g01988(.A0(n3566), .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B0(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3557), .Y(n5023));
  NAND4X1 g01989(.A(n5022), .B(n5021), .C(n5020), .D(n5023), .Y(n5024));
  NOR2X1  g01990(.A(n5024), .B(n5019), .Y(n5025));
  NOR4X1  g01991(.A(n3719), .B(n3894), .C(n3618), .D(n5025), .Y(n5026));
  AOI22X1 g01992(.A0(n5014), .A1(n5026), .B0(n3858), .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .Y(n5027));
  AOI22X1 g01993(.A0(n3921), .A1(n5013), .B0(n3860), .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .Y(n5029));
  NOR3X1  g01994(.A(n3791), .B(n3667), .C(n3706), .Y(n5030));
  INVX1   g01995(.A(n5030), .Y(n5031));
  NOR3X1  g01996(.A(n3728), .B(n3894), .C(n3618), .Y(n5032));
  INVX1   g01997(.A(n5032), .Y(n5033));
  AOI21X1 g01998(.A0(n5033), .A1(n5031), .B0(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .Y(n5034));
  NOR3X1  g01999(.A(n3791), .B(n3789), .C(n3714), .Y(n5035));
  INVX1   g02000(.A(n5035), .Y(n5036));
  NAND4X1 g02001(.A(n3711), .B(n3584), .C(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .D(n3727), .Y(n5037));
  OAI21X1 g02002(.A0(n5036), .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B0(n5037), .Y(n5038));
  INVX1   g02003(.A(n5025), .Y(n5039));
  NOR4X1  g02004(.A(n3719), .B(n3894), .C(n3618), .D(n5039), .Y(n5040));
  INVX1   g02005(.A(n5040), .Y(n5041));
  NOR2X1  g02006(.A(n5041), .B(n5013), .Y(n5042));
  INVX1   g02007(.A(n3805), .Y(n5043));
  NOR3X1  g02008(.A(n3793), .B(n3789), .C(n3731), .Y(n5044));
  NOR3X1  g02009(.A(n3793), .B(n3789), .C(n3701), .Y(n5045));
  OAI21X1 g02010(.A0(n5045), .A1(n5044), .B0(n3960), .Y(n5046));
  OAI21X1 g02011(.A0(n5043), .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B0(n5046), .Y(n5047));
  NOR4X1  g02012(.A(n5042), .B(n5038), .C(n5034), .D(n5047), .Y(n5048));
  OAI21X1 g02013(.A0(n3732), .A1(n3720), .B0(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .Y(n5049));
  OAI21X1 g02014(.A0(n3924), .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B0(n5049), .Y(n5050));
  AOI21X1 g02015(.A0(n3835), .A1(n3797), .B0(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .Y(n5051));
  NAND4X1 g02016(.A(n3700), .B(n3584), .C(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .D(n3711), .Y(n5052));
  OAI21X1 g02017(.A0(n3925), .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B0(n5052), .Y(n5053));
  NOR3X1  g02018(.A(n5053), .B(n5051), .C(n5050), .Y(n5054));
  NAND4X1 g02019(.A(n5048), .B(n5029), .C(n5027), .D(n5054), .Y(n5055));
  AOI21X1 g02020(.A0(n3787), .A1(n3960), .B0(n5055), .Y(n5056));
  AOI22X1 g02021(.A0(n4983), .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B0(P3_REIP_REG_0__SCAN_IN), .B1(n4968), .Y(n5058));
  OAI21X1 g02022(.A0(n5056), .A1(n4985), .B0(n5058), .Y(P3_U2862));
  NAND2X1 g02023(.A(n3973), .B(n3787), .Y(n5061));
  AOI22X1 g02024(.A0(n3577), .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B0(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(n3550), .Y(n5062));
  AOI22X1 g02025(.A0(n3574), .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B0(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3562), .Y(n5063));
  AOI22X1 g02026(.A0(n3555), .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B0(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3575), .Y(n5064));
  AOI22X1 g02027(.A0(n3572), .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B0(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3568), .Y(n5065));
  NAND4X1 g02028(.A(n5064), .B(n5063), .C(n5062), .D(n5065), .Y(n5066));
  AOI22X1 g02029(.A0(n3565), .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B0(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3563), .Y(n5067));
  AOI22X1 g02030(.A0(n3578), .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B0(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3569), .Y(n5068));
  AOI22X1 g02031(.A0(n3571), .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B0(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3560), .Y(n5069));
  AOI22X1 g02032(.A0(n3566), .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B0(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3557), .Y(n5070));
  NAND4X1 g02033(.A(n5069), .B(n5068), .C(n5067), .D(n5070), .Y(n5071));
  NOR2X1  g02034(.A(n5071), .B(n5066), .Y(n5072));
  NOR2X1  g02035(.A(n5012), .B(n3960), .Y(n5073));
  XOR2X1  g02036(.A(n5073), .B(n3967), .Y(n5074));
  NOR4X1  g02037(.A(n5066), .B(n5012), .C(n3960), .D(n5071), .Y(n5075));
  INVX1   g02038(.A(n5072), .Y(n5076));
  NOR3X1  g02039(.A(n5076), .B(n5073), .C(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .Y(n5077));
  AOI21X1 g02040(.A0(n5075), .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B0(n5077), .Y(n5078));
  OAI21X1 g02041(.A0(n5074), .A1(n5072), .B0(n5078), .Y(n5079));
  OAI21X1 g02042(.A0(n5040), .A1(n5026), .B0(n5079), .Y(n5080));
  XOR2X1  g02043(.A(n5076), .B(n5012), .Y(n5081));
  INVX1   g02044(.A(n5081), .Y(n5082));
  NOR3X1  g02045(.A(n5011), .B(n4998), .C(n3960), .Y(n5083));
  XOR2X1  g02046(.A(n5083), .B(n3967), .Y(n5084));
  NOR4X1  g02047(.A(n5011), .B(n4998), .C(n3960), .D(n5072), .Y(n5085));
  NOR3X1  g02048(.A(n5081), .B(n5083), .C(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .Y(n5086));
  AOI21X1 g02049(.A0(n5085), .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B0(n5086), .Y(n5087));
  OAI21X1 g02050(.A0(n5084), .A1(n5082), .B0(n5087), .Y(n5088));
  NAND3X1 g02051(.A(n5088), .B(n3799), .C(n3730), .Y(n5089));
  NAND2X1 g02052(.A(n3860), .B(n3967), .Y(n5090));
  NAND2X1 g02053(.A(n3858), .B(n3967), .Y(n5091));
  NAND4X1 g02054(.A(n3792), .B(n3788), .C(n3730), .D(n3973), .Y(n5092));
  OAI21X1 g02055(.A0(n5045), .A1(n3805), .B0(n3973), .Y(n5093));
  NAND4X1 g02056(.A(n5092), .B(n5091), .C(n5090), .D(n5093), .Y(n5094));
  OAI21X1 g02057(.A0(n3834), .A1(n3798), .B0(n3973), .Y(n5095));
  OAI21X1 g02058(.A0(n3917), .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B0(n5095), .Y(n5096));
  OAI21X1 g02059(.A0(n3745), .A1(n3702), .B0(n3973), .Y(n5097));
  OAI21X1 g02060(.A0(n5035), .A1(n5030), .B0(n3973), .Y(n5098));
  AOI22X1 g02061(.A0(n3973), .A1(n5032), .B0(n3713), .B1(n3967), .Y(n5099));
  OAI21X1 g02062(.A0(n3732), .A1(n3720), .B0(n3967), .Y(n5100));
  NAND4X1 g02063(.A(n5099), .B(n5098), .C(n5097), .D(n5100), .Y(n5101));
  NOR3X1  g02064(.A(n5101), .B(n5096), .C(n5094), .Y(n5102));
  NAND4X1 g02065(.A(n5089), .B(n5080), .C(n5061), .D(n5102), .Y(n5103));
  AOI22X1 g02066(.A0(n4984), .A1(n5103), .B0(n4983), .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .Y(n5104));
  OAI21X1 g02067(.A0(n4969), .A1(n3399), .B0(n5104), .Y(P3_U2861));
  OAI21X1 g02068(.A0(n5082), .A1(n5083), .B0(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .Y(n5106));
  INVX1   g02069(.A(n5106), .Y(n5107));
  NOR2X1  g02070(.A(n5107), .B(n5085), .Y(n5108));
  INVX1   g02071(.A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .Y(n5109));
  AOI22X1 g02072(.A0(n3577), .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B0(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3550), .Y(n5110));
  AOI22X1 g02073(.A0(n3574), .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B0(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3562), .Y(n5111));
  AOI22X1 g02074(.A0(n3555), .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B0(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3575), .Y(n5112));
  AOI22X1 g02075(.A0(n3572), .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B0(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3568), .Y(n5113));
  NAND4X1 g02076(.A(n5112), .B(n5111), .C(n5110), .D(n5113), .Y(n5114));
  AOI22X1 g02077(.A0(n3565), .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B0(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3563), .Y(n5115));
  AOI22X1 g02078(.A0(n3578), .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B0(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3569), .Y(n5116));
  AOI22X1 g02079(.A0(n3571), .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B0(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3560), .Y(n5117));
  AOI22X1 g02080(.A0(n3566), .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B0(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3557), .Y(n5118));
  NAND4X1 g02081(.A(n5117), .B(n5116), .C(n5115), .D(n5118), .Y(n5119));
  NOR2X1  g02082(.A(n5119), .B(n5114), .Y(n5120));
  INVX1   g02083(.A(n5120), .Y(n5121));
  NOR2X1  g02084(.A(n5072), .B(n5012), .Y(n5122));
  XOR2X1  g02085(.A(n5122), .B(n5121), .Y(n5123));
  XOR2X1  g02086(.A(n5123), .B(n5109), .Y(n5124));
  NAND2X1 g02087(.A(n5108), .B(n5124), .Y(n5125));
  OAI21X1 g02088(.A0(n5124), .A1(n5108), .B0(n5125), .Y(n5127));
  NAND2X1 g02089(.A(n5127), .B(n3921), .Y(n5128));
  NAND2X1 g02090(.A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .Y(n5129));
  XOR2X1  g02091(.A(n5129), .B(n5109), .Y(n5130));
  NAND2X1 g02092(.A(n5130), .B(n3787), .Y(n5131));
  XOR2X1  g02093(.A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n3967), .Y(n5132));
  INVX1   g02094(.A(n5132), .Y(n5133));
  NAND2X1 g02095(.A(n5133), .B(n3858), .Y(n5134));
  NAND2X1 g02096(.A(n5133), .B(n3860), .Y(n5135));
  NAND4X1 g02097(.A(n3803), .B(n3759), .C(n3718), .D(n5130), .Y(n5136));
  OAI21X1 g02098(.A0(n5045), .A1(n5044), .B0(n5130), .Y(n5137));
  NAND4X1 g02099(.A(n5136), .B(n5135), .C(n5134), .D(n5137), .Y(n5138));
  OAI21X1 g02100(.A0(n3732), .A1(n3720), .B0(n5133), .Y(n5140));
  OAI21X1 g02101(.A0(n5130), .A1(n3924), .B0(n5140), .Y(n5141));
  OAI21X1 g02102(.A0(n5030), .A1(n3798), .B0(n5130), .Y(n5142));
  INVX1   g02103(.A(n5130), .Y(n5143));
  AOI22X1 g02104(.A0(n5133), .A1(n3713), .B0(n3745), .B1(n5143), .Y(n5144));
  AOI22X1 g02105(.A0(n5130), .A1(n3834), .B0(n3729), .B1(n5133), .Y(n5145));
  OAI21X1 g02106(.A0(n5035), .A1(n5032), .B0(n5130), .Y(n5146));
  NAND4X1 g02107(.A(n5145), .B(n5144), .C(n5142), .D(n5146), .Y(n5147));
  NOR3X1  g02108(.A(n5147), .B(n5141), .C(n5138), .Y(n5148));
  XOR2X1  g02109(.A(n5120), .B(n5076), .Y(n5149));
  INVX1   g02110(.A(n5075), .Y(n5151));
  OAI21X1 g02111(.A0(n5072), .A1(n5073), .B0(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .Y(n5152));
  NAND2X1 g02112(.A(n5152), .B(n5151), .Y(n5153));
  NOR2X1  g02113(.A(n5149), .B(n5109), .Y(n5156));
  XOR2X1  g02114(.A(n5149), .B(n5109), .Y(n5159));
  XOR2X1  g02115(.A(n5153), .B(n5159), .Y(n5162));
  AOI22X1 g02116(.A0(n5162), .A1(n5026), .B0(n5040), .B1(n5162), .Y(n5163));
  NAND4X1 g02117(.A(n5148), .B(n5131), .C(n5128), .D(n5163), .Y(n5164));
  AOI22X1 g02118(.A0(n4984), .A1(n5164), .B0(n4983), .B1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .Y(n5165));
  OAI21X1 g02119(.A0(n4969), .A1(n3396), .B0(n5165), .Y(P3_U2860));
  AOI22X1 g02120(.A0(n5149), .A1(n5109), .B0(n5151), .B1(n5152), .Y(n5167));
  NOR2X1  g02121(.A(n5167), .B(n5156), .Y(n5168));
  INVX1   g02122(.A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .Y(n5169));
  AOI22X1 g02123(.A0(n3577), .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B0(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3550), .Y(n5170));
  AOI22X1 g02124(.A0(n3574), .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B0(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3562), .Y(n5171));
  AOI22X1 g02125(.A0(n3555), .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B0(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3575), .Y(n5172));
  AOI22X1 g02126(.A0(n3572), .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B0(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3568), .Y(n5173));
  NAND4X1 g02127(.A(n5172), .B(n5171), .C(n5170), .D(n5173), .Y(n5174));
  AOI22X1 g02128(.A0(n3565), .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B0(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3563), .Y(n5175));
  AOI22X1 g02129(.A0(n3578), .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B0(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3569), .Y(n5176));
  AOI22X1 g02130(.A0(n3571), .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B0(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3560), .Y(n5177));
  AOI22X1 g02131(.A0(n3566), .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B0(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3557), .Y(n5178));
  NAND4X1 g02132(.A(n5177), .B(n5176), .C(n5175), .D(n5178), .Y(n5179));
  NOR2X1  g02133(.A(n5179), .B(n5174), .Y(n5180));
  NOR2X1  g02134(.A(n5120), .B(n5072), .Y(n5181));
  XOR2X1  g02135(.A(n5181), .B(n5180), .Y(n5182));
  AOI21X1 g02136(.A0(n5182), .A1(n5169), .B0(n5168), .Y(n5183));
  NOR2X1  g02137(.A(n5182), .B(n5169), .Y(n5184));
  INVX1   g02138(.A(n5184), .Y(n5185));
  XOR2X1  g02139(.A(n5182), .B(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .Y(n5186));
  AOI22X1 g02140(.A0(n5185), .A1(n5183), .B0(n5168), .B1(n5186), .Y(n5187));
  NAND2X1 g02141(.A(n5187), .B(n5040), .Y(n5188));
  NOR2X1  g02142(.A(n5123), .B(n5109), .Y(n5189));
  INVX1   g02143(.A(n5189), .Y(n5190));
  NOR2X1  g02144(.A(n5122), .B(n5121), .Y(n5191));
  XOR2X1  g02145(.A(n5180), .B(n5191), .Y(n5192));
  INVX1   g02146(.A(n5123), .Y(n5193));
  OAI22X1 g02147(.A0(n5193), .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B0(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(n5192), .Y(n5194));
  AOI21X1 g02148(.A0(n5192), .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B0(n5194), .Y(n5195));
  INVX1   g02149(.A(n5195), .Y(n5196));
  AOI21X1 g02150(.A0(n5190), .A1(n5108), .B0(n5196), .Y(n5197));
  OAI22X1 g02151(.A0(n5193), .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B0(n5085), .B1(n5107), .Y(n5198));
  INVX1   g02152(.A(n5192), .Y(n5199));
  AOI21X1 g02153(.A0(n5192), .A1(n5169), .B0(n5189), .Y(n5200));
  INVX1   g02154(.A(n5200), .Y(n5201));
  AOI21X1 g02155(.A0(n5199), .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B0(n5201), .Y(n5202));
  AOI21X1 g02156(.A0(n5202), .A1(n5198), .B0(n5197), .Y(n5203));
  NAND2X1 g02157(.A(n5203), .B(n3921), .Y(n5204));
  INVX1   g02158(.A(n5180), .Y(n5207));
  NAND2X1 g02159(.A(n5187), .B(n5026), .Y(n5213));
  NOR2X1  g02160(.A(n5129), .B(n5109), .Y(n5214));
  XOR2X1  g02161(.A(n5214), .B(n5169), .Y(n5215));
  INVX1   g02162(.A(n5215), .Y(n5216));
  NAND2X1 g02163(.A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .Y(n5217));
  XOR2X1  g02164(.A(n5217), .B(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .Y(n5218));
  NOR4X1  g02165(.A(n3760), .B(n3707), .C(n3600), .D(n5218), .Y(n5219));
  NOR4X1  g02166(.A(n3760), .B(n3634), .C(n3600), .D(n5218), .Y(n5220));
  OAI21X1 g02167(.A0(n5045), .A1(n5044), .B0(n5216), .Y(n5221));
  OAI21X1 g02168(.A0(n5215), .A1(n5043), .B0(n5221), .Y(n5222));
  NOR3X1  g02169(.A(n5222), .B(n5220), .C(n5219), .Y(n5223));
  AOI21X1 g02170(.A0(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B0(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .Y(n5224));
  XOR2X1  g02171(.A(n5224), .B(n5169), .Y(n5225));
  AOI21X1 g02172(.A0(n3918), .A1(n3920), .B0(n5218), .Y(n5226));
  AOI21X1 g02173(.A0(n5225), .A1(n3702), .B0(n5226), .Y(n5227));
  OAI21X1 g02174(.A0(n3834), .A1(n3798), .B0(n5216), .Y(n5228));
  AOI22X1 g02175(.A0(n5216), .A1(n5032), .B0(n3745), .B1(n5225), .Y(n5229));
  NAND2X1 g02176(.A(n5229), .B(n5228), .Y(n5230));
  OAI22X1 g02177(.A0(n5215), .A1(n5036), .B0(n3753), .B1(n5218), .Y(n5231));
  OAI22X1 g02178(.A0(n5215), .A1(n5031), .B0(n3917), .B1(n5218), .Y(n5232));
  NOR3X1  g02179(.A(n5232), .B(n5231), .C(n5230), .Y(n5233));
  NAND3X1 g02180(.A(n5233), .B(n5227), .C(n5223), .Y(n5234));
  AOI21X1 g02181(.A0(n5216), .A1(n3787), .B0(n5234), .Y(n5235));
  NAND4X1 g02182(.A(n5213), .B(n5204), .C(n5188), .D(n5235), .Y(n5236));
  AOI22X1 g02183(.A0(n4984), .A1(n5236), .B0(n4983), .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .Y(n5237));
  OAI21X1 g02184(.A0(n4969), .A1(n3393), .B0(n5237), .Y(P3_U2859));
  NOR2X1  g02185(.A(n5184), .B(n5183), .Y(n5239));
  NOR3X1  g02186(.A(n5180), .B(n5120), .C(n5072), .Y(n5240));
  AOI22X1 g02187(.A0(n3577), .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B0(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(n3550), .Y(n5241));
  AOI22X1 g02188(.A0(n3574), .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B0(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3562), .Y(n5242));
  AOI22X1 g02189(.A0(n3555), .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B0(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3575), .Y(n5243));
  AOI22X1 g02190(.A0(n3572), .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B0(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3568), .Y(n5244));
  NAND4X1 g02191(.A(n5243), .B(n5242), .C(n5241), .D(n5244), .Y(n5245));
  AOI22X1 g02192(.A0(n3565), .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B0(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3563), .Y(n5246));
  AOI22X1 g02193(.A0(n3578), .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B0(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3569), .Y(n5247));
  AOI22X1 g02194(.A0(n3571), .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B0(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3560), .Y(n5248));
  AOI22X1 g02195(.A0(n3566), .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B0(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3557), .Y(n5249));
  NAND4X1 g02196(.A(n5248), .B(n5247), .C(n5246), .D(n5249), .Y(n5250));
  NOR2X1  g02197(.A(n5250), .B(n5245), .Y(n5251));
  XOR2X1  g02198(.A(n5251), .B(n5240), .Y(n5252));
  XOR2X1  g02199(.A(n5252), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .Y(n5253));
  AOI21X1 g02200(.A0(n5252), .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B0(n5184), .Y(n5254));
  OAI21X1 g02201(.A0(n5252), .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B0(n5254), .Y(n5255));
  OAI22X1 g02202(.A0(n5253), .A1(n5239), .B0(n5183), .B1(n5255), .Y(n5256));
  NOR2X1  g02203(.A(n5256), .B(n5041), .Y(n5257));
  AOI21X1 g02204(.A0(n5199), .A1(n5190), .B0(n5169), .Y(n5258));
  AOI21X1 g02205(.A0(n5192), .A1(n5189), .B0(n5258), .Y(n5259));
  OAI21X1 g02206(.A0(n5194), .A1(n5108), .B0(n5259), .Y(n5260));
  NOR2X1  g02207(.A(n5180), .B(n5191), .Y(n5261));
  XOR2X1  g02208(.A(n5251), .B(n5261), .Y(n5262));
  XOR2X1  g02209(.A(n5262), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .Y(n5263));
  NOR2X1  g02210(.A(n5260), .B(n5263), .Y(n5264));
  AOI21X1 g02211(.A0(n5263), .A1(n5260), .B0(n5264), .Y(n5266));
  NOR2X1  g02212(.A(n5266), .B(n3922), .Y(n5267));
  INVX1   g02213(.A(n5026), .Y(n5268));
  AOI22X1 g02214(.A0(n5149), .A1(n5109), .B0(n5169), .B1(n5182), .Y(n5271));
  OAI21X1 g02215(.A0(n5156), .A1(n5153), .B0(n5271), .Y(n5272));
  INVX1   g02216(.A(n5251), .Y(n5275));
  XOR2X1  g02217(.A(n5275), .B(n5240), .Y(n5276));
  NOR2X1  g02218(.A(n5256), .B(n5268), .Y(n5281));
  NAND4X1 g02219(.A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .D(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .Y(n5282));
  XOR2X1  g02220(.A(n5282), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .Y(n5283));
  NAND3X1 g02221(.A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .C(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .Y(n5284));
  XOR2X1  g02222(.A(n5284), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .Y(n5285));
  INVX1   g02223(.A(n5285), .Y(n5286));
  NAND2X1 g02224(.A(n5286), .B(n3858), .Y(n5287));
  NAND2X1 g02225(.A(n5286), .B(n3860), .Y(n5288));
  INVX1   g02226(.A(n5283), .Y(n5289));
  NAND4X1 g02227(.A(n3803), .B(n3759), .C(n3718), .D(n5289), .Y(n5290));
  OAI21X1 g02228(.A0(n5045), .A1(n5044), .B0(n5289), .Y(n5291));
  NAND4X1 g02229(.A(n5290), .B(n5288), .C(n5287), .D(n5291), .Y(n5292));
  INVX1   g02230(.A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .Y(n5293));
  NOR2X1  g02231(.A(n5224), .B(n5169), .Y(n5294));
  XOR2X1  g02232(.A(n5294), .B(n5293), .Y(n5295));
  OAI21X1 g02233(.A0(n3732), .A1(n3720), .B0(n5286), .Y(n5296));
  OAI21X1 g02234(.A0(n5295), .A1(n3924), .B0(n5296), .Y(n5297));
  OAI21X1 g02235(.A0(n5030), .A1(n3798), .B0(n5289), .Y(n5298));
  INVX1   g02236(.A(n5295), .Y(n5299));
  AOI22X1 g02237(.A0(n5286), .A1(n3713), .B0(n3745), .B1(n5299), .Y(n5300));
  AOI22X1 g02238(.A0(n5289), .A1(n3834), .B0(n3729), .B1(n5286), .Y(n5301));
  OAI21X1 g02239(.A0(n5035), .A1(n5032), .B0(n5289), .Y(n5302));
  NAND4X1 g02240(.A(n5301), .B(n5300), .C(n5298), .D(n5302), .Y(n5303));
  NOR3X1  g02241(.A(n5303), .B(n5297), .C(n5292), .Y(n5304));
  OAI21X1 g02242(.A0(n5283), .A1(n3786), .B0(n5304), .Y(n5305));
  NOR4X1  g02243(.A(n5281), .B(n5267), .C(n5257), .D(n5305), .Y(n5306));
  AOI22X1 g02244(.A0(n4983), .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B0(P3_REIP_REG_4__SCAN_IN), .B1(n4968), .Y(n5307));
  OAI21X1 g02245(.A0(n5306), .A1(n4985), .B0(n5307), .Y(P3_U2858));
  NOR2X1  g02246(.A(n5262), .B(n5293), .Y(n5309));
  AOI22X1 g02247(.A0(n3577), .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B0(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3550), .Y(n5310));
  AOI22X1 g02248(.A0(n3574), .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B0(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3562), .Y(n5311));
  AOI22X1 g02249(.A0(n3555), .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B0(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3575), .Y(n5312));
  AOI22X1 g02250(.A0(n3572), .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B0(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3568), .Y(n5313));
  NAND4X1 g02251(.A(n5312), .B(n5311), .C(n5310), .D(n5313), .Y(n5314));
  AOI22X1 g02252(.A0(n3565), .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B0(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3563), .Y(n5315));
  AOI22X1 g02253(.A0(n3578), .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B0(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3569), .Y(n5316));
  AOI22X1 g02254(.A0(n3571), .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B0(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3560), .Y(n5317));
  AOI22X1 g02255(.A0(n3566), .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B0(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3557), .Y(n5318));
  NAND4X1 g02256(.A(n5317), .B(n5316), .C(n5315), .D(n5318), .Y(n5319));
  NOR2X1  g02257(.A(n5319), .B(n5314), .Y(n5320));
  NOR3X1  g02258(.A(n5251), .B(n5180), .C(n5191), .Y(n5321));
  XOR2X1  g02259(.A(n5321), .B(n5320), .Y(n5322));
  INVX1   g02260(.A(n5322), .Y(n5323));
  INVX1   g02261(.A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .Y(n5324));
  AOI22X1 g02262(.A0(n5262), .A1(n5293), .B0(n5324), .B1(n5322), .Y(n5325));
  INVX1   g02263(.A(n5325), .Y(n5326));
  AOI21X1 g02264(.A0(n5323), .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B0(n5326), .Y(n5327));
  OAI21X1 g02265(.A0(n5309), .A1(n5260), .B0(n5327), .Y(n5328));
  INVX1   g02266(.A(n5328), .Y(n5329));
  INVX1   g02267(.A(n5262), .Y(n5330));
  NOR2X1  g02268(.A(n5330), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .Y(n5331));
  INVX1   g02269(.A(n5331), .Y(n5332));
  AOI21X1 g02270(.A0(n5323), .A1(n5324), .B0(n5309), .Y(n5333));
  OAI21X1 g02271(.A0(n5323), .A1(n5324), .B0(n5333), .Y(n5334));
  AOI21X1 g02272(.A0(n5332), .A1(n5260), .B0(n5334), .Y(n5335));
  NOR3X1  g02273(.A(n5335), .B(n5329), .C(n3922), .Y(n5336));
  NOR2X1  g02274(.A(n5252), .B(n5293), .Y(n5337));
  AOI22X1 g02275(.A0(n5182), .A1(n5169), .B0(n5293), .B1(n5252), .Y(n5338));
  INVX1   g02276(.A(n5338), .Y(n5339));
  NOR2X1  g02277(.A(n5339), .B(n5168), .Y(n5340));
  NOR3X1  g02278(.A(n5349), .B(n5340), .C(n5337), .Y(n5342));
  NOR4X1  g02279(.A(n5180), .B(n5120), .C(n5072), .D(n5251), .Y(n5343));
  XOR2X1  g02280(.A(n5320), .B(n5343), .Y(n5344));
  XOR2X1  g02281(.A(n5344), .B(n5324), .Y(n5345));
  XOR2X1  g02282(.A(n5345), .B(n5342), .Y(n5346));
  NOR2X1  g02283(.A(n5346), .B(n5041), .Y(n5347));
  NOR2X1  g02284(.A(n5276), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .Y(n5348));
  NOR3X1  g02285(.A(n5348), .B(n5182), .C(n5169), .Y(n5349));
  AOI21X1 g02286(.A0(n5276), .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B0(n5349), .Y(n5350));
  OAI21X1 g02287(.A0(n5348), .A1(n5272), .B0(n5350), .Y(n5351));
  INVX1   g02288(.A(n5343), .Y(n5352));
  NOR2X1  g02289(.A(n5320), .B(n5251), .Y(n5353));
  AOI22X1 g02290(.A0(n5320), .A1(n5352), .B0(n5240), .B1(n5353), .Y(n5354));
  NOR2X1  g02291(.A(n5346), .B(n5268), .Y(n5357));
  NOR2X1  g02292(.A(n5282), .B(n5293), .Y(n5358));
  XOR2X1  g02293(.A(n5358), .B(n5324), .Y(n5359));
  NAND4X1 g02294(.A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .C(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .D(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .Y(n5360));
  XOR2X1  g02295(.A(n5360), .B(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .Y(n5361));
  INVX1   g02296(.A(n5361), .Y(n5362));
  NAND2X1 g02297(.A(n5362), .B(n3860), .Y(n5363));
  NAND2X1 g02298(.A(n5362), .B(n3858), .Y(n5364));
  NAND4X1 g02299(.A(n3803), .B(n3759), .C(n3718), .D(n5368), .Y(n5366));
  XOR2X1  g02300(.A(n5358), .B(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .Y(n5368));
  AOI22X1 g02301(.A0(n5368), .A1(n5044), .B0(n5045), .B1(n5368), .Y(n5369));
  NAND4X1 g02302(.A(n5366), .B(n5364), .C(n5363), .D(n5369), .Y(n5370));
  OAI21X1 g02303(.A0(n3732), .A1(n3713), .B0(n5362), .Y(n5371));
  OAI21X1 g02304(.A0(n5361), .A1(n3920), .B0(n5371), .Y(n5372));
  NOR3X1  g02305(.A(n5224), .B(n5293), .C(n5169), .Y(n5373));
  XOR2X1  g02306(.A(n5373), .B(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .Y(n5374));
  AOI22X1 g02307(.A0(n5368), .A1(n5032), .B0(n3745), .B1(n5374), .Y(n5375));
  AOI22X1 g02308(.A0(n5368), .A1(n5035), .B0(n3702), .B1(n5374), .Y(n5376));
  AOI22X1 g02309(.A0(n5368), .A1(n3834), .B0(n3729), .B1(n5362), .Y(n5377));
  OAI21X1 g02310(.A0(n5030), .A1(n3798), .B0(n5368), .Y(n5378));
  NAND4X1 g02311(.A(n5377), .B(n5376), .C(n5375), .D(n5378), .Y(n5379));
  NOR3X1  g02312(.A(n5379), .B(n5372), .C(n5370), .Y(n5380));
  OAI21X1 g02313(.A0(n5359), .A1(n3786), .B0(n5380), .Y(n5381));
  NOR4X1  g02314(.A(n5357), .B(n5347), .C(n5336), .D(n5381), .Y(n5382));
  AOI22X1 g02315(.A0(n4983), .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B0(P3_REIP_REG_5__SCAN_IN), .B1(n4968), .Y(n5383));
  OAI21X1 g02316(.A0(n5382), .A1(n4985), .B0(n5383), .Y(P3_U2857));
  AOI22X1 g02317(.A0(n3577), .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B0(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3550), .Y(n5389));
  AOI22X1 g02318(.A0(n3574), .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B0(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3562), .Y(n5390));
  AOI22X1 g02319(.A0(n3555), .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B0(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3575), .Y(n5391));
  AOI22X1 g02320(.A0(n3572), .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B0(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3568), .Y(n5392));
  NAND4X1 g02321(.A(n5391), .B(n5390), .C(n5389), .D(n5392), .Y(n5393));
  AOI22X1 g02322(.A0(n3565), .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B0(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3563), .Y(n5394));
  AOI22X1 g02323(.A0(n3578), .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B0(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3569), .Y(n5395));
  AOI22X1 g02324(.A0(n3571), .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B0(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3560), .Y(n5396));
  AOI22X1 g02325(.A0(n3566), .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B0(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3557), .Y(n5397));
  NAND4X1 g02326(.A(n5396), .B(n5395), .C(n5394), .D(n5397), .Y(n5398));
  NOR2X1  g02327(.A(n5398), .B(n5393), .Y(n5399));
  NOR2X1  g02328(.A(n5320), .B(n5352), .Y(n5400));
  XOR2X1  g02329(.A(n5400), .B(n5399), .Y(n5401));
  NOR2X1  g02330(.A(n5416), .B(n5041), .Y(n5404));
  NOR2X1  g02331(.A(n5354), .B(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .Y(n5405));
  INVX1   g02332(.A(n5405), .Y(n5406));
  NAND2X1 g02333(.A(n5354), .B(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .Y(n5407));
  INVX1   g02334(.A(n5407), .Y(n5408));
  AOI21X1 g02335(.A0(n5406), .A1(n5351), .B0(n5408), .Y(n5409));
  INVX1   g02336(.A(n5409), .Y(n5410));
  INVX1   g02337(.A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .Y(n5411));
  INVX1   g02338(.A(n5320), .Y(n5412));
  NAND3X1 g02339(.A(n5412), .B(n5275), .C(n5240), .Y(n5413));
  XOR2X1  g02340(.A(n5399), .B(n5413), .Y(n5414));
  XOR2X1  g02341(.A(n5414), .B(n5411), .Y(n5415));
  XOR2X1  g02342(.A(n5415), .B(n5410), .Y(n5416));
  NOR2X1  g02343(.A(n5416), .B(n5268), .Y(n5417));
  INVX1   g02344(.A(n5260), .Y(n5418));
  NOR3X1  g02345(.A(n5322), .B(n5262), .C(n5293), .Y(n5419));
  OAI21X1 g02346(.A0(n5262), .A1(n5293), .B0(n5322), .Y(n5420));
  AOI21X1 g02347(.A0(n5420), .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .B0(n5419), .Y(n5421));
  OAI21X1 g02348(.A0(n5326), .A1(n5418), .B0(n5421), .Y(n5422));
  NOR4X1  g02349(.A(n5251), .B(n5180), .C(n5191), .D(n5320), .Y(n5423));
  XOR2X1  g02350(.A(n5423), .B(n5399), .Y(n5424));
  XOR2X1  g02351(.A(n5424), .B(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .Y(n5425));
  XOR2X1  g02352(.A(n5425), .B(n5422), .Y(n5426));
  NOR2X1  g02353(.A(n5426), .B(n3922), .Y(n5427));
  NOR3X1  g02354(.A(n5282), .B(n5324), .C(n5293), .Y(n5428));
  XOR2X1  g02355(.A(n5428), .B(n5411), .Y(n5429));
  NOR2X1  g02356(.A(n5360), .B(n5324), .Y(n5430));
  XOR2X1  g02357(.A(n5430), .B(n5411), .Y(n5431));
  INVX1   g02358(.A(n5431), .Y(n5432));
  NAND2X1 g02359(.A(n5432), .B(n3860), .Y(n5433));
  NAND2X1 g02360(.A(n5432), .B(n3858), .Y(n5434));
  INVX1   g02361(.A(n5429), .Y(n5435));
  NAND4X1 g02362(.A(n3803), .B(n3759), .C(n3718), .D(n5435), .Y(n5436));
  AOI22X1 g02363(.A0(n5435), .A1(n5044), .B0(n5045), .B1(n5435), .Y(n5439));
  NAND4X1 g02364(.A(n5436), .B(n5434), .C(n5433), .D(n5439), .Y(n5440));
  OAI21X1 g02365(.A0(n3732), .A1(n3713), .B0(n5432), .Y(n5441));
  OAI21X1 g02366(.A0(n5431), .A1(n3920), .B0(n5441), .Y(n5442));
  NOR4X1  g02367(.A(n5324), .B(n5293), .C(n5169), .D(n5224), .Y(n5443));
  XOR2X1  g02368(.A(n5443), .B(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .Y(n5444));
  AOI22X1 g02369(.A0(n5435), .A1(n5032), .B0(n3745), .B1(n5444), .Y(n5445));
  AOI22X1 g02370(.A0(n5435), .A1(n5035), .B0(n3702), .B1(n5444), .Y(n5446));
  AOI22X1 g02371(.A0(n5435), .A1(n3834), .B0(n3729), .B1(n5432), .Y(n5447));
  OAI21X1 g02372(.A0(n5030), .A1(n3798), .B0(n5435), .Y(n5448));
  NAND4X1 g02373(.A(n5447), .B(n5446), .C(n5445), .D(n5448), .Y(n5449));
  NOR3X1  g02374(.A(n5449), .B(n5442), .C(n5440), .Y(n5450));
  OAI21X1 g02375(.A0(n5429), .A1(n3786), .B0(n5450), .Y(n5451));
  NOR4X1  g02376(.A(n5427), .B(n5417), .C(n5404), .D(n5451), .Y(n5452));
  AOI22X1 g02377(.A0(n4983), .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B0(P3_REIP_REG_6__SCAN_IN), .B1(n4968), .Y(n5453));
  OAI21X1 g02378(.A0(n5452), .A1(n4985), .B0(n5453), .Y(P3_U2856));
  NOR2X1  g02379(.A(n5401), .B(n5411), .Y(n5455));
  NOR3X1  g02380(.A(n5399), .B(n5320), .C(n5352), .Y(n5459));
  XOR2X1  g02381(.A(n5459), .B(n5025), .Y(n5460));
  XOR2X1  g02382(.A(n5460), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Y(n5461));
  NOR2X1  g02383(.A(n5474), .B(n5041), .Y(n5463));
  AOI21X1 g02384(.A0(n5401), .A1(n5411), .B0(n5409), .Y(n5466));
  NOR2X1  g02385(.A(n5466), .B(n5455), .Y(n5467));
  INVX1   g02386(.A(n5467), .Y(n5468));
  NOR2X1  g02387(.A(n5399), .B(n5025), .Y(n5470));
  INVX1   g02388(.A(n5470), .Y(n5471));
  XOR2X1  g02389(.A(n5461), .B(n5468), .Y(n5474));
  NOR2X1  g02390(.A(n5474), .B(n5268), .Y(n5475));
  NAND2X1 g02391(.A(n5424), .B(n5411), .Y(n5476));
  NAND2X1 g02392(.A(n5476), .B(n5422), .Y(n5477));
  OAI21X1 g02393(.A0(n5424), .A1(n5411), .B0(n5477), .Y(n5478));
  INVX1   g02394(.A(n5423), .Y(n5479));
  NOR2X1  g02395(.A(n5479), .B(n5399), .Y(n5480));
  XOR2X1  g02396(.A(n5480), .B(n5025), .Y(n5481));
  XOR2X1  g02397(.A(n5481), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Y(n5482));
  XOR2X1  g02398(.A(n5482), .B(n5478), .Y(n5483));
  INVX1   g02399(.A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Y(n5484));
  NOR4X1  g02400(.A(n5411), .B(n5324), .C(n5293), .D(n5282), .Y(n5485));
  XOR2X1  g02401(.A(n5485), .B(n5484), .Y(n5486));
  NOR2X1  g02402(.A(n5486), .B(n3786), .Y(n5487));
  NOR3X1  g02403(.A(n5360), .B(n5411), .C(n5324), .Y(n5488));
  XOR2X1  g02404(.A(n5488), .B(n5484), .Y(n5489));
  INVX1   g02405(.A(n5489), .Y(n5490));
  NAND2X1 g02406(.A(n5490), .B(n3860), .Y(n5491));
  NAND2X1 g02407(.A(n5490), .B(n3858), .Y(n5492));
  INVX1   g02408(.A(n5486), .Y(n5493));
  NAND4X1 g02409(.A(n3803), .B(n3759), .C(n3718), .D(n5493), .Y(n5494));
  AOI22X1 g02410(.A0(n5493), .A1(n5044), .B0(n5045), .B1(n5493), .Y(n5498));
  NAND4X1 g02411(.A(n5494), .B(n5492), .C(n5491), .D(n5498), .Y(n5499));
  OAI21X1 g02412(.A0(n3732), .A1(n3713), .B0(n5490), .Y(n5500));
  OAI21X1 g02413(.A0(n5489), .A1(n3920), .B0(n5500), .Y(n5501));
  NAND2X1 g02414(.A(n5443), .B(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .Y(n5502));
  XOR2X1  g02415(.A(n5502), .B(n5484), .Y(n5503));
  AOI22X1 g02416(.A0(n5493), .A1(n5032), .B0(n3745), .B1(n5503), .Y(n5504));
  AOI22X1 g02417(.A0(n5493), .A1(n5035), .B0(n3702), .B1(n5503), .Y(n5505));
  AOI22X1 g02418(.A0(n5493), .A1(n3834), .B0(n3729), .B1(n5490), .Y(n5506));
  OAI21X1 g02419(.A0(n5030), .A1(n3798), .B0(n5493), .Y(n5507));
  NAND4X1 g02420(.A(n5506), .B(n5505), .C(n5504), .D(n5507), .Y(n5508));
  NOR4X1  g02421(.A(n5501), .B(n5499), .C(n5487), .D(n5508), .Y(n5509));
  OAI21X1 g02422(.A0(n5483), .A1(n3922), .B0(n5509), .Y(n5510));
  NOR3X1  g02423(.A(n5510), .B(n5475), .C(n5463), .Y(n5511));
  AOI22X1 g02424(.A0(n4983), .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B0(P3_REIP_REG_7__SCAN_IN), .B1(n4968), .Y(n5512));
  OAI21X1 g02425(.A0(n5511), .A1(n4985), .B0(n5512), .Y(P3_U2855));
  INVX1   g02426(.A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .Y(n5517));
  NOR3X1  g02427(.A(n5471), .B(n5320), .C(n5352), .Y(n5518));
  XOR2X1  g02428(.A(n5518), .B(n5517), .Y(n5519));
  XOR2X1  g02429(.A(n5519), .B(n5571), .Y(n5520));
  NOR2X1  g02430(.A(n5520), .B(n5041), .Y(n5521));
  INVX1   g02431(.A(n5481), .Y(n5522));
  OAI21X1 g02432(.A0(n5522), .A1(n5478), .B0(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Y(n5523));
  INVX1   g02433(.A(n5523), .Y(n5524));
  AOI21X1 g02434(.A0(n5522), .A1(n5478), .B0(n5524), .Y(n5525));
  NOR2X1  g02435(.A(n5471), .B(n5479), .Y(n5526));
  XOR2X1  g02436(.A(n5526), .B(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .Y(n5527));
  XOR2X1  g02437(.A(n5527), .B(n5525), .Y(n5528));
  NOR2X1  g02438(.A(n5528), .B(n3922), .Y(n5529));
  AOI21X1 g02439(.A0(n5460), .A1(n5484), .B0(n5467), .Y(n5530));
  NOR2X1  g02440(.A(n5460), .B(n5484), .Y(n5531));
  NOR2X1  g02441(.A(n5531), .B(n5530), .Y(n5532));
  XOR2X1  g02442(.A(n5519), .B(n5532), .Y(n5535));
  NAND2X1 g02443(.A(n5485), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Y(n5536));
  XOR2X1  g02444(.A(n5536), .B(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .Y(n5537));
  NOR2X1  g02445(.A(n5537), .B(n3786), .Y(n5538));
  NOR4X1  g02446(.A(n5484), .B(n5411), .C(n5324), .D(n5360), .Y(n5539));
  XOR2X1  g02447(.A(n5539), .B(n5517), .Y(n5540));
  INVX1   g02448(.A(n5540), .Y(n5541));
  NAND2X1 g02449(.A(n5541), .B(n3860), .Y(n5542));
  NAND2X1 g02450(.A(n5541), .B(n3858), .Y(n5543));
  NAND4X1 g02451(.A(n3803), .B(n3759), .C(n3718), .D(n5547), .Y(n5545));
  XOR2X1  g02452(.A(n5536), .B(n5517), .Y(n5547));
  AOI22X1 g02453(.A0(n5547), .A1(n5044), .B0(n5045), .B1(n5547), .Y(n5548));
  NAND4X1 g02454(.A(n5545), .B(n5543), .C(n5542), .D(n5548), .Y(n5549));
  OAI21X1 g02455(.A0(n3732), .A1(n3713), .B0(n5541), .Y(n5550));
  OAI21X1 g02456(.A0(n5540), .A1(n3920), .B0(n5550), .Y(n5551));
  NAND3X1 g02457(.A(n5443), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .C(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .Y(n5552));
  XOR2X1  g02458(.A(n5552), .B(n5517), .Y(n5553));
  AOI22X1 g02459(.A0(n5547), .A1(n5032), .B0(n3745), .B1(n5553), .Y(n5554));
  AOI22X1 g02460(.A0(n5547), .A1(n5035), .B0(n3702), .B1(n5553), .Y(n5555));
  AOI22X1 g02461(.A0(n5547), .A1(n3834), .B0(n3729), .B1(n5541), .Y(n5556));
  OAI21X1 g02462(.A0(n5030), .A1(n3798), .B0(n5547), .Y(n5557));
  NAND4X1 g02463(.A(n5556), .B(n5555), .C(n5554), .D(n5557), .Y(n5558));
  NOR4X1  g02464(.A(n5551), .B(n5549), .C(n5538), .D(n5558), .Y(n5559));
  OAI21X1 g02465(.A0(n5535), .A1(n5268), .B0(n5559), .Y(n5560));
  NOR3X1  g02466(.A(n5560), .B(n5529), .C(n5521), .Y(n5561));
  AOI22X1 g02467(.A0(n4983), .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B0(P3_REIP_REG_8__SCAN_IN), .B1(n4968), .Y(n5562));
  OAI21X1 g02468(.A0(n5561), .A1(n4985), .B0(n5562), .Y(P3_U2854));
  INVX1   g02469(.A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .Y(n5564));
  NOR4X1  g02470(.A(n5320), .B(n5352), .C(n5517), .D(n5471), .Y(n5565));
  NOR2X1  g02471(.A(n5518), .B(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .Y(n5566));
  INVX1   g02472(.A(n5566), .Y(n5567));
  AOI21X1 g02473(.A0(n5567), .A1(n5571), .B0(n5565), .Y(n5568));
  XOR2X1  g02474(.A(n5568), .B(n5564), .Y(n5569));
  INVX1   g02475(.A(n5518), .Y(n5570));
  INVX1   g02476(.A(n5532), .Y(n5571));
  OAI21X1 g02477(.A0(n5571), .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B0(n5570), .Y(n5572));
  OAI21X1 g02478(.A0(n5532), .A1(n5517), .B0(n5572), .Y(n5573));
  XOR2X1  g02479(.A(n5518), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .Y(n5574));
  NAND2X1 g02480(.A(n5574), .B(n5573), .Y(n5576));
  OAI21X1 g02481(.A0(n5574), .A1(n5573), .B0(n5576), .Y(n5577));
  NAND2X1 g02482(.A(n5577), .B(n5026), .Y(n5578));
  AOI21X1 g02483(.A0(n5470), .A1(n5423), .B0(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .Y(n5579));
  NOR2X1  g02484(.A(n5579), .B(n5525), .Y(n5580));
  AOI21X1 g02485(.A0(n5526), .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B0(n5580), .Y(n5581));
  XOR2X1  g02486(.A(n5581), .B(n5564), .Y(n5582));
  NAND2X1 g02487(.A(n5582), .B(n3921), .Y(n5583));
  NAND3X1 g02488(.A(n5485), .B(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .C(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Y(n5584));
  XOR2X1  g02489(.A(n5584), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .Y(n5585));
  NOR2X1  g02490(.A(n5585), .B(n3786), .Y(n5586));
  NAND2X1 g02491(.A(n5539), .B(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .Y(n5587));
  XOR2X1  g02492(.A(n5587), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .Y(n5588));
  NOR4X1  g02493(.A(n3760), .B(n3707), .C(n3600), .D(n5588), .Y(n5589));
  NOR4X1  g02494(.A(n3760), .B(n3634), .C(n3600), .D(n5588), .Y(n5590));
  NOR4X1  g02495(.A(n3804), .B(n3802), .C(n3719), .D(n5585), .Y(n5591));
  INVX1   g02496(.A(n5044), .Y(n5592));
  INVX1   g02497(.A(n5045), .Y(n5593));
  OAI22X1 g02498(.A0(n5585), .A1(n5592), .B0(n5593), .B1(n5585), .Y(n5596));
  NOR4X1  g02499(.A(n5591), .B(n5590), .C(n5589), .D(n5596), .Y(n5597));
  NOR4X1  g02500(.A(n3719), .B(n3717), .C(n3618), .D(n5588), .Y(n5598));
  AOI21X1 g02501(.A0(n3918), .A1(n3753), .B0(n5588), .Y(n5599));
  NOR2X1  g02502(.A(n5599), .B(n5598), .Y(n5600));
  NAND4X1 g02503(.A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .C(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .D(n5443), .Y(n5601));
  XOR2X1  g02504(.A(n5601), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .Y(n5602));
  OAI22X1 g02505(.A0(n5585), .A1(n5033), .B0(n3925), .B1(n5602), .Y(n5603));
  OAI22X1 g02506(.A0(n5585), .A1(n5036), .B0(n3924), .B1(n5602), .Y(n5604));
  AOI21X1 g02507(.A0(n3835), .A1(n3797), .B0(n5585), .Y(n5605));
  OAI22X1 g02508(.A0(n5585), .A1(n5031), .B0(n3917), .B1(n5588), .Y(n5606));
  NOR4X1  g02509(.A(n5605), .B(n5604), .C(n5603), .D(n5606), .Y(n5607));
  NAND3X1 g02510(.A(n5607), .B(n5600), .C(n5597), .Y(n5608));
  NOR2X1  g02511(.A(n5608), .B(n5586), .Y(n5609));
  NAND3X1 g02512(.A(n5609), .B(n5583), .C(n5578), .Y(n5610));
  AOI21X1 g02513(.A0(n5569), .A1(n5040), .B0(n5610), .Y(n5611));
  AOI22X1 g02514(.A0(n4983), .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B0(P3_REIP_REG_9__SCAN_IN), .B1(n4968), .Y(n5612));
  OAI21X1 g02515(.A0(n5611), .A1(n4985), .B0(n5612), .Y(P3_U2853));
  INVX1   g02516(.A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .Y(n5614));
  OAI21X1 g02517(.A0(n5568), .A1(n5564), .B0(n5614), .Y(n5615));
  NOR3X1  g02518(.A(n5568), .B(n5614), .C(n5564), .Y(n5616));
  INVX1   g02519(.A(n5616), .Y(n5617));
  NAND2X1 g02520(.A(n5617), .B(n5615), .Y(n5618));
  NOR2X1  g02521(.A(n5618), .B(n5041), .Y(n5619));
  OAI21X1 g02522(.A0(n5570), .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B0(n5573), .Y(n5620));
  OAI21X1 g02523(.A0(n5518), .A1(n5564), .B0(n5620), .Y(n5621));
  XOR2X1  g02524(.A(n5518), .B(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .Y(n5622));
  NOR2X1  g02525(.A(n5622), .B(n5621), .Y(n5623));
  AOI21X1 g02526(.A0(n5622), .A1(n5621), .B0(n5623), .Y(n5625));
  NOR2X1  g02527(.A(n5625), .B(n5268), .Y(n5626));
  OAI21X1 g02528(.A0(n5581), .A1(n5564), .B0(n5614), .Y(n5627));
  NOR3X1  g02529(.A(n5581), .B(n5614), .C(n5564), .Y(n5628));
  INVX1   g02530(.A(n5628), .Y(n5629));
  NAND2X1 g02531(.A(n5629), .B(n5627), .Y(n5630));
  NAND4X1 g02532(.A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .C(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .D(n5485), .Y(n5631));
  XOR2X1  g02533(.A(n5631), .B(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .Y(n5632));
  NOR2X1  g02534(.A(n5632), .B(n3786), .Y(n5633));
  NAND3X1 g02535(.A(n5539), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .Y(n5634));
  XOR2X1  g02536(.A(n5634), .B(n5614), .Y(n5635));
  NAND2X1 g02537(.A(n5635), .B(n3858), .Y(n5636));
  NAND2X1 g02538(.A(n5635), .B(n3860), .Y(n5637));
  INVX1   g02539(.A(n5632), .Y(n5638));
  NAND4X1 g02540(.A(n3803), .B(n3759), .C(n3718), .D(n5638), .Y(n5639));
  AOI22X1 g02541(.A0(n5638), .A1(n5044), .B0(n5045), .B1(n5638), .Y(n5642));
  NAND4X1 g02542(.A(n5639), .B(n5637), .C(n5636), .D(n5642), .Y(n5643));
  NOR2X1  g02543(.A(n5601), .B(n5564), .Y(n5644));
  XOR2X1  g02544(.A(n5644), .B(n5614), .Y(n5645));
  INVX1   g02545(.A(n5645), .Y(n5646));
  AOI22X1 g02546(.A0(n5638), .A1(n5032), .B0(n3745), .B1(n5646), .Y(n5647));
  OAI21X1 g02547(.A0(n5632), .A1(n5036), .B0(n5647), .Y(n5648));
  OAI21X1 g02548(.A0(n3732), .A1(n3713), .B0(n5635), .Y(n5649));
  AOI22X1 g02549(.A0(n5635), .A1(n3720), .B0(n3702), .B1(n5646), .Y(n5650));
  AOI22X1 g02550(.A0(n5638), .A1(n3834), .B0(n3729), .B1(n5635), .Y(n5651));
  OAI21X1 g02551(.A0(n5030), .A1(n3798), .B0(n5638), .Y(n5652));
  NAND4X1 g02552(.A(n5651), .B(n5650), .C(n5649), .D(n5652), .Y(n5653));
  NOR4X1  g02553(.A(n5648), .B(n5643), .C(n5633), .D(n5653), .Y(n5654));
  OAI21X1 g02554(.A0(n5630), .A1(n3922), .B0(n5654), .Y(n5655));
  NOR3X1  g02555(.A(n5655), .B(n5626), .C(n5619), .Y(n5656));
  AOI22X1 g02556(.A0(n4983), .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B0(P3_REIP_REG_10__SCAN_IN), .B1(n4968), .Y(n5657));
  OAI21X1 g02557(.A0(n5656), .A1(n4985), .B0(n5657), .Y(P3_U2852));
  OAI21X1 g02558(.A0(n5614), .A1(n5564), .B0(n5518), .Y(n5659));
  OAI22X1 g02559(.A0(n5413), .A1(n5471), .B0(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .Y(n5660));
  INVX1   g02560(.A(n5660), .Y(n5661));
  AOI21X1 g02561(.A0(n5659), .A1(n5573), .B0(n5661), .Y(n5662));
  XOR2X1  g02562(.A(n5518), .B(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .Y(n5663));
  XOR2X1  g02563(.A(n5663), .B(n5662), .Y(n5664));
  INVX1   g02564(.A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .Y(n5665));
  XOR2X1  g02565(.A(n5616), .B(n5665), .Y(n5666));
  XOR2X1  g02566(.A(n5628), .B(n5665), .Y(n5667));
  NOR2X1  g02567(.A(n5667), .B(n3922), .Y(n5668));
  NOR2X1  g02568(.A(n5631), .B(n5614), .Y(n5669));
  XOR2X1  g02569(.A(n5669), .B(n5665), .Y(n5670));
  NAND4X1 g02570(.A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .D(n5539), .Y(n5671));
  XOR2X1  g02571(.A(n5671), .B(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .Y(n5672));
  INVX1   g02572(.A(n5672), .Y(n5673));
  NAND2X1 g02573(.A(n5673), .B(n3858), .Y(n5674));
  NAND2X1 g02574(.A(n5673), .B(n3860), .Y(n5675));
  INVX1   g02575(.A(n5670), .Y(n5676));
  AOI22X1 g02576(.A0(n5676), .A1(n3834), .B0(n5045), .B1(n5676), .Y(n5679));
  NAND3X1 g02577(.A(n5679), .B(n5675), .C(n5674), .Y(n5680));
  AOI21X1 g02578(.A0(n3918), .A1(n3753), .B0(n5672), .Y(n5681));
  NOR3X1  g02579(.A(n5601), .B(n5614), .C(n5564), .Y(n5682));
  XOR2X1  g02580(.A(n5682), .B(n5665), .Y(n5683));
  OAI22X1 g02581(.A0(n5672), .A1(n3920), .B0(n3924), .B1(n5683), .Y(n5684));
  OAI21X1 g02582(.A0(n5035), .A1(n3798), .B0(n5676), .Y(n5685));
  INVX1   g02583(.A(n5683), .Y(n5686));
  AOI22X1 g02584(.A0(n5676), .A1(n3805), .B0(n3745), .B1(n5686), .Y(n5687));
  OAI21X1 g02585(.A0(n5044), .A1(n5030), .B0(n5676), .Y(n5688));
  AOI22X1 g02586(.A0(n5676), .A1(n5032), .B0(n3729), .B1(n5673), .Y(n5689));
  NAND4X1 g02587(.A(n5688), .B(n5687), .C(n5685), .D(n5689), .Y(n5690));
  NOR4X1  g02588(.A(n5684), .B(n5681), .C(n5680), .D(n5690), .Y(n5691));
  OAI21X1 g02589(.A0(n5670), .A1(n3786), .B0(n5691), .Y(n5692));
  NOR2X1  g02590(.A(n5692), .B(n5668), .Y(n5693));
  OAI21X1 g02591(.A0(n5666), .A1(n5041), .B0(n5693), .Y(n5694));
  AOI21X1 g02592(.A0(n5664), .A1(n5026), .B0(n5694), .Y(n5695));
  AOI22X1 g02593(.A0(n4983), .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B0(P3_REIP_REG_11__SCAN_IN), .B1(n4968), .Y(n5696));
  OAI21X1 g02594(.A0(n5695), .A1(n4985), .B0(n5696), .Y(P3_U2851));
  AOI21X1 g02595(.A0(n5616), .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B0(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Y(n5698));
  INVX1   g02596(.A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Y(n5699));
  NOR3X1  g02597(.A(n5617), .B(n5699), .C(n5665), .Y(n5700));
  NOR3X1  g02598(.A(n5700), .B(n5698), .C(n5041), .Y(n5701));
  OAI21X1 g02599(.A0(n5570), .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B0(n5659), .Y(n5702));
  INVX1   g02600(.A(n5702), .Y(n5703));
  AOI21X1 g02601(.A0(n5570), .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B0(n5661), .Y(n5704));
  INVX1   g02602(.A(n5704), .Y(n5705));
  AOI21X1 g02603(.A0(n5703), .A1(n5573), .B0(n5705), .Y(n5706));
  INVX1   g02604(.A(n5706), .Y(n5707));
  XOR2X1  g02605(.A(n5518), .B(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Y(n5708));
  NOR2X1  g02606(.A(n5707), .B(n5708), .Y(n5709));
  AOI21X1 g02607(.A0(n5708), .A1(n5707), .B0(n5709), .Y(n5711));
  NOR2X1  g02608(.A(n5711), .B(n5268), .Y(n5712));
  AOI21X1 g02609(.A0(n5628), .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B0(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Y(n5713));
  NOR3X1  g02610(.A(n5629), .B(n5699), .C(n5665), .Y(n5714));
  NOR3X1  g02611(.A(n5714), .B(n5713), .C(n3922), .Y(n5715));
  NOR3X1  g02612(.A(n5631), .B(n5665), .C(n5614), .Y(n5716));
  XOR2X1  g02613(.A(n5716), .B(n5699), .Y(n5717));
  NOR2X1  g02614(.A(n5671), .B(n5665), .Y(n5718));
  XOR2X1  g02615(.A(n5718), .B(n5699), .Y(n5719));
  INVX1   g02616(.A(n5719), .Y(n5720));
  OAI21X1 g02617(.A0(n3732), .A1(n3720), .B0(n5720), .Y(n5721));
  OAI21X1 g02618(.A0(n5719), .A1(n3753), .B0(n5721), .Y(n5722));
  INVX1   g02619(.A(n5717), .Y(n5723));
  NAND4X1 g02620(.A(n3803), .B(n3759), .C(n3700), .D(n5723), .Y(n5724));
  AOI22X1 g02621(.A0(n5720), .A1(n3729), .B0(n5045), .B1(n5723), .Y(n5727));
  OAI21X1 g02622(.A0(n5032), .A1(n5030), .B0(n5723), .Y(n5728));
  NAND3X1 g02623(.A(n5728), .B(n5727), .C(n5724), .Y(n5729));
  NOR4X1  g02624(.A(n5665), .B(n5614), .C(n5564), .D(n5601), .Y(n5730));
  XOR2X1  g02625(.A(n5730), .B(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Y(n5731));
  AOI22X1 g02626(.A0(n5720), .A1(n3860), .B0(n3702), .B1(n5731), .Y(n5732));
  AOI22X1 g02627(.A0(n5723), .A1(n3798), .B0(n3745), .B1(n5731), .Y(n5733));
  OAI21X1 g02628(.A0(n5035), .A1(n3805), .B0(n5723), .Y(n5734));
  AOI22X1 g02629(.A0(n5723), .A1(n5044), .B0(n3858), .B1(n5720), .Y(n5735));
  NAND4X1 g02630(.A(n5734), .B(n5733), .C(n5732), .D(n5735), .Y(n5736));
  NOR3X1  g02631(.A(n5736), .B(n5729), .C(n5722), .Y(n5737));
  OAI21X1 g02632(.A0(n5717), .A1(n3786), .B0(n5737), .Y(n5738));
  NOR4X1  g02633(.A(n5715), .B(n5712), .C(n5701), .D(n5738), .Y(n5739));
  AOI22X1 g02634(.A0(n4983), .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B0(P3_REIP_REG_12__SCAN_IN), .B1(n4968), .Y(n5740));
  OAI21X1 g02635(.A0(n5739), .A1(n4985), .B0(n5740), .Y(P3_U2850));
  NOR2X1  g02636(.A(n5518), .B(n5699), .Y(n5742));
  INVX1   g02637(.A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .Y(n5743));
  NOR2X1  g02638(.A(n5518), .B(n5743), .Y(n5744));
  AOI21X1 g02639(.A0(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B0(n5570), .Y(n5745));
  NOR2X1  g02640(.A(n5745), .B(n5744), .Y(n5746));
  OAI21X1 g02641(.A0(n5742), .A1(n5707), .B0(n5746), .Y(n5747));
  AOI21X1 g02642(.A0(n5518), .A1(n5699), .B0(n5706), .Y(n5748));
  OAI22X1 g02643(.A0(n5413), .A1(n5471), .B0(n5743), .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Y(n5749));
  OAI21X1 g02644(.A0(n5570), .A1(n5743), .B0(n5749), .Y(n5750));
  OAI21X1 g02645(.A0(n5750), .A1(n5748), .B0(n5747), .Y(n5751));
  INVX1   g02646(.A(n5751), .Y(n5752));
  XOR2X1  g02647(.A(n5700), .B(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .Y(n5753));
  NAND2X1 g02648(.A(n5753), .B(n5040), .Y(n5754));
  XOR2X1  g02649(.A(n5714), .B(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .Y(n5755));
  NAND2X1 g02650(.A(n5755), .B(n3921), .Y(n5756));
  NOR3X1  g02651(.A(n5671), .B(n5699), .C(n5665), .Y(n5757));
  XOR2X1  g02652(.A(n5757), .B(n5743), .Y(n5758));
  INVX1   g02653(.A(n5758), .Y(n5759));
  OAI21X1 g02654(.A0(n3732), .A1(n3720), .B0(n5759), .Y(n5760));
  OAI21X1 g02655(.A0(n5758), .A1(n3917), .B0(n5760), .Y(n5761));
  OAI22X1 g02656(.A0(n5758), .A1(n3753), .B0(n5593), .B1(n5767), .Y(n5764));
  AOI21X1 g02657(.A0(n3861), .A1(n3859), .B0(n5758), .Y(n5765));
  NOR4X1  g02658(.A(n5699), .B(n5665), .C(n5614), .D(n5631), .Y(n5766));
  XOR2X1  g02659(.A(n5766), .B(n5743), .Y(n5767));
  AOI21X1 g02660(.A0(n3835), .A1(n5043), .B0(n5767), .Y(n5768));
  NOR4X1  g02661(.A(n5765), .B(n5764), .C(n5761), .D(n5768), .Y(n5769));
  NOR2X1  g02662(.A(n5767), .B(n3786), .Y(n5770));
  NAND2X1 g02663(.A(n5730), .B(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Y(n5771));
  XOR2X1  g02664(.A(n5771), .B(n5743), .Y(n5772));
  OAI21X1 g02665(.A0(n3745), .A1(n3702), .B0(n5772), .Y(n5773));
  OAI21X1 g02666(.A0(n5767), .A1(n3797), .B0(n5773), .Y(n5774));
  AOI21X1 g02667(.A0(n5036), .A1(n5033), .B0(n5767), .Y(n5775));
  AOI21X1 g02668(.A0(n5592), .A1(n5031), .B0(n5767), .Y(n5776));
  NOR4X1  g02669(.A(n5775), .B(n5774), .C(n5770), .D(n5776), .Y(n5777));
  NAND4X1 g02670(.A(n5769), .B(n5756), .C(n5754), .D(n5777), .Y(n5778));
  AOI21X1 g02671(.A0(n5752), .A1(n5026), .B0(n5778), .Y(n5779));
  AOI22X1 g02672(.A0(n4983), .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B0(P3_REIP_REG_13__SCAN_IN), .B1(n4968), .Y(n5780));
  OAI21X1 g02673(.A0(n5779), .A1(n4985), .B0(n5780), .Y(P3_U2849));
  INVX1   g02674(.A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .Y(n5782));
  NOR4X1  g02675(.A(n5743), .B(n5699), .C(n5665), .D(n5617), .Y(n5783));
  XOR2X1  g02676(.A(n5783), .B(n5782), .Y(n5784));
  NOR2X1  g02677(.A(n5784), .B(n5041), .Y(n5785));
  NOR4X1  g02678(.A(n5743), .B(n5699), .C(n5665), .D(n5629), .Y(n5786));
  XOR2X1  g02679(.A(n5786), .B(n5782), .Y(n5787));
  INVX1   g02680(.A(n5573), .Y(n5788));
  NOR3X1  g02681(.A(n5745), .B(n5702), .C(n5788), .Y(n5789));
  NOR4X1  g02682(.A(n5744), .B(n5742), .C(n5705), .D(n5789), .Y(n5790));
  XOR2X1  g02683(.A(n5518), .B(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .Y(n5791));
  XOR2X1  g02684(.A(n5791), .B(n5790), .Y(n5792));
  NOR4X1  g02685(.A(n5743), .B(n5699), .C(n5665), .D(n5671), .Y(n5793));
  XOR2X1  g02686(.A(n5793), .B(n5782), .Y(n5794));
  OAI22X1 g02687(.A0(n5794), .A1(n3917), .B0(n5593), .B1(n5800), .Y(n5797));
  AOI21X1 g02688(.A0(n3918), .A1(n3920), .B0(n5794), .Y(n5798));
  NAND2X1 g02689(.A(n5766), .B(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .Y(n5799));
  XOR2X1  g02690(.A(n5799), .B(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .Y(n5800));
  AOI21X1 g02691(.A0(n5036), .A1(n5033), .B0(n5800), .Y(n5801));
  NOR4X1  g02692(.A(n3712), .B(n3701), .C(n3583), .D(n5794), .Y(n5802));
  AOI21X1 g02693(.A0(n3861), .A1(n3859), .B0(n5794), .Y(n5803));
  NOR2X1  g02694(.A(n5803), .B(n5802), .Y(n5804));
  OAI21X1 g02695(.A0(n5800), .A1(n3786), .B0(n5804), .Y(n5805));
  NOR4X1  g02696(.A(n5801), .B(n5798), .C(n5797), .D(n5805), .Y(n5806));
  NAND3X1 g02697(.A(n5730), .B(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Y(n5807));
  XOR2X1  g02698(.A(n5807), .B(n5782), .Y(n5808));
  OAI21X1 g02699(.A0(n3745), .A1(n3702), .B0(n5808), .Y(n5809));
  OAI21X1 g02700(.A0(n5800), .A1(n3797), .B0(n5809), .Y(n5810));
  AOI21X1 g02701(.A0(n5592), .A1(n5031), .B0(n5800), .Y(n5811));
  AOI21X1 g02702(.A0(n3835), .A1(n5043), .B0(n5800), .Y(n5812));
  NOR3X1  g02703(.A(n5812), .B(n5811), .C(n5810), .Y(n5813));
  NAND2X1 g02704(.A(n5813), .B(n5806), .Y(n5814));
  AOI21X1 g02705(.A0(n5792), .A1(n5026), .B0(n5814), .Y(n5815));
  OAI21X1 g02706(.A0(n5787), .A1(n3922), .B0(n5815), .Y(n5816));
  OAI21X1 g02707(.A0(n5816), .A1(n5785), .B0(n4984), .Y(n5817));
  AOI22X1 g02708(.A0(n4983), .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B0(P3_REIP_REG_14__SCAN_IN), .B1(n4968), .Y(n5818));
  NAND2X1 g02709(.A(n5818), .B(n5817), .Y(P3_U2848));
  AOI21X1 g02710(.A0(n5783), .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B0(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .Y(n5820));
  NAND4X1 g02711(.A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .D(n5700), .Y(n5821));
  INVX1   g02712(.A(n5821), .Y(n5822));
  NOR3X1  g02713(.A(n5822), .B(n5820), .C(n5041), .Y(n5823));
  AOI21X1 g02714(.A0(n5518), .A1(n5782), .B0(n5790), .Y(n5824));
  AOI21X1 g02715(.A0(n5570), .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B0(n5824), .Y(n5825));
  INVX1   g02716(.A(n5825), .Y(n5826));
  XOR2X1  g02717(.A(n5518), .B(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .Y(n5827));
  XOR2X1  g02718(.A(n5827), .B(n5826), .Y(n5828));
  NOR2X1  g02719(.A(n5828), .B(n5268), .Y(n5829));
  AOI21X1 g02720(.A0(n5786), .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B0(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .Y(n5830));
  NAND4X1 g02721(.A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .D(n5714), .Y(n5831));
  INVX1   g02722(.A(n5831), .Y(n5832));
  NOR3X1  g02723(.A(n5832), .B(n5830), .C(n3922), .Y(n5833));
  NAND2X1 g02724(.A(n5793), .B(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .Y(n5834));
  XOR2X1  g02725(.A(n5834), .B(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .Y(n5835));
  INVX1   g02726(.A(n5835), .Y(n5836));
  OAI21X1 g02727(.A0(n3860), .A1(n3858), .B0(n5836), .Y(n5837));
  OAI21X1 g02728(.A0(n5835), .A1(n3753), .B0(n5837), .Y(n5838));
  INVX1   g02729(.A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .Y(n5839));
  OAI22X1 g02730(.A0(n5835), .A1(n3917), .B0(n5593), .B1(n5845), .Y(n5842));
  AOI21X1 g02731(.A0(n3918), .A1(n3920), .B0(n5835), .Y(n5843));
  NAND3X1 g02732(.A(n5766), .B(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .Y(n5844));
  XOR2X1  g02733(.A(n5844), .B(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .Y(n5845));
  AOI21X1 g02734(.A0(n5031), .A1(n3786), .B0(n5845), .Y(n5846));
  NOR4X1  g02735(.A(n5843), .B(n5842), .C(n5838), .D(n5846), .Y(n5847));
  NAND4X1 g02736(.A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .D(n5730), .Y(n5848));
  XOR2X1  g02737(.A(n5848), .B(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .Y(n5849));
  AOI21X1 g02738(.A0(n3925), .A1(n3924), .B0(n5849), .Y(n5850));
  AOI21X1 g02739(.A0(n5036), .A1(n3797), .B0(n5845), .Y(n5851));
  AOI21X1 g02740(.A0(n5592), .A1(n5033), .B0(n5845), .Y(n5852));
  AOI21X1 g02741(.A0(n3835), .A1(n5043), .B0(n5845), .Y(n5853));
  NOR4X1  g02742(.A(n5852), .B(n5851), .C(n5850), .D(n5853), .Y(n5854));
  NAND2X1 g02743(.A(n5854), .B(n5847), .Y(n5855));
  NOR4X1  g02744(.A(n5833), .B(n5829), .C(n5823), .D(n5855), .Y(n5856));
  AOI22X1 g02745(.A0(n4983), .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B0(P3_REIP_REG_15__SCAN_IN), .B1(n4968), .Y(n5857));
  OAI21X1 g02746(.A0(n5856), .A1(n4985), .B0(n5857), .Y(P3_U2847));
  NOR2X1  g02747(.A(n5518), .B(n5839), .Y(n5859));
  AOI21X1 g02748(.A0(n5518), .A1(n5839), .B0(n5825), .Y(n5860));
  NOR2X1  g02749(.A(n5860), .B(n5859), .Y(n5861));
  INVX1   g02750(.A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .Y(n5862));
  XOR2X1  g02751(.A(n5518), .B(n5862), .Y(n5863));
  XOR2X1  g02752(.A(n5863), .B(n5861), .Y(n5864));
  NOR2X1  g02753(.A(n5864), .B(n5268), .Y(n5865));
  XOR2X1  g02754(.A(n5821), .B(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .Y(n5866));
  NOR2X1  g02755(.A(n5866), .B(n5041), .Y(n5867));
  XOR2X1  g02756(.A(n5831), .B(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .Y(n5868));
  NOR2X1  g02757(.A(n5868), .B(n3922), .Y(n5869));
  NAND3X1 g02758(.A(n5793), .B(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .C(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .Y(n5870));
  XOR2X1  g02759(.A(n5870), .B(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .Y(n5871));
  INVX1   g02760(.A(n5871), .Y(n5872));
  OAI21X1 g02761(.A0(n3860), .A1(n3729), .B0(n5872), .Y(n5873));
  OAI21X1 g02762(.A0(n5871), .A1(n3918), .B0(n5873), .Y(n5874));
  OAI22X1 g02763(.A0(n5871), .A1(n3753), .B0(n5593), .B1(n5882), .Y(n5877));
  AOI21X1 g02764(.A0(n3859), .A1(n3920), .B0(n5871), .Y(n5878));
  NOR2X1  g02765(.A(n5848), .B(n5839), .Y(n5879));
  XOR2X1  g02766(.A(n5879), .B(n5862), .Y(n5880));
  NAND4X1 g02767(.A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .D(n5766), .Y(n5881));
  XOR2X1  g02768(.A(n5881), .B(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .Y(n5882));
  OAI22X1 g02769(.A0(n5880), .A1(n3924), .B0(n5043), .B1(n5882), .Y(n5883));
  NOR4X1  g02770(.A(n5878), .B(n5877), .C(n5874), .D(n5883), .Y(n5884));
  OAI22X1 g02771(.A0(n5880), .A1(n3925), .B0(n5033), .B1(n5882), .Y(n5885));
  AOI21X1 g02772(.A0(n5036), .A1(n3797), .B0(n5882), .Y(n5886));
  AOI21X1 g02773(.A0(n5031), .A1(n3835), .B0(n5882), .Y(n5887));
  AOI21X1 g02774(.A0(n5592), .A1(n3786), .B0(n5882), .Y(n5888));
  NOR4X1  g02775(.A(n5887), .B(n5886), .C(n5885), .D(n5888), .Y(n5889));
  NAND2X1 g02776(.A(n5889), .B(n5884), .Y(n5890));
  NOR4X1  g02777(.A(n5869), .B(n5867), .C(n5865), .D(n5890), .Y(n5891));
  AOI22X1 g02778(.A0(n4983), .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B0(P3_REIP_REG_16__SCAN_IN), .B1(n4968), .Y(n5892));
  OAI21X1 g02779(.A0(n5891), .A1(n4985), .B0(n5892), .Y(P3_U2846));
  INVX1   g02780(.A(n5861), .Y(n5894));
  INVX1   g02781(.A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .Y(n5895));
  NOR2X1  g02782(.A(n5895), .B(n5862), .Y(n5896));
  AOI21X1 g02783(.A0(n5896), .A1(n5894), .B0(n5570), .Y(n5897));
  NOR3X1  g02784(.A(n5860), .B(n5859), .C(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .Y(n5898));
  NOR2X1  g02785(.A(n5518), .B(n5895), .Y(n5899));
  NOR3X1  g02786(.A(n5899), .B(n5898), .C(n5897), .Y(n5900));
  AOI21X1 g02787(.A0(n5898), .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B0(n5518), .Y(n5901));
  INVX1   g02788(.A(n5901), .Y(n5902));
  AOI22X1 g02789(.A0(n5518), .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B0(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B1(n5894), .Y(n5903));
  AOI21X1 g02790(.A0(n5903), .A1(n5902), .B0(n5900), .Y(n5904));
  AOI21X1 g02791(.A0(n5822), .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B0(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .Y(n5905));
  INVX1   g02792(.A(n5896), .Y(n5906));
  NOR2X1  g02793(.A(n5906), .B(n5821), .Y(n5907));
  NOR2X1  g02794(.A(n5907), .B(n5905), .Y(n5908));
  NAND2X1 g02795(.A(n5908), .B(n5040), .Y(n5909));
  AOI21X1 g02796(.A0(n5832), .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B0(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .Y(n5910));
  NOR2X1  g02797(.A(n5906), .B(n5831), .Y(n5911));
  NOR3X1  g02798(.A(n5911), .B(n5910), .C(n3922), .Y(n5912));
  NAND4X1 g02799(.A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .C(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .D(n5793), .Y(n5913));
  XOR2X1  g02800(.A(n5913), .B(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .Y(n5914));
  INVX1   g02801(.A(n5914), .Y(n5915));
  AOI21X1 g02802(.A0(n3859), .A1(n3753), .B0(n5914), .Y(n5916));
  AOI21X1 g02803(.A0(n5915), .A1(n3732), .B0(n5916), .Y(n5917));
  AOI22X1 g02804(.A0(n5915), .A1(n3860), .B0(n5045), .B1(n5928), .Y(n5921));
  OAI21X1 g02805(.A0(n3729), .A1(n3720), .B0(n5915), .Y(n5922));
  NOR3X1  g02806(.A(n5848), .B(n5862), .C(n5839), .Y(n5923));
  XOR2X1  g02807(.A(n5923), .B(n5895), .Y(n5924));
  INVX1   g02808(.A(n5924), .Y(n5925));
  NOR2X1  g02809(.A(n5881), .B(n5862), .Y(n5926));
  XOR2X1  g02810(.A(n5926), .B(n5895), .Y(n5927));
  INVX1   g02811(.A(n5927), .Y(n5928));
  AOI22X1 g02812(.A0(n5925), .A1(n3745), .B0(n3805), .B1(n5928), .Y(n5929));
  NAND4X1 g02813(.A(n5922), .B(n5921), .C(n5917), .D(n5929), .Y(n5930));
  OAI21X1 g02814(.A0(n3834), .A1(n3787), .B0(n5928), .Y(n5931));
  AOI22X1 g02815(.A0(n5925), .A1(n3702), .B0(n5044), .B1(n5928), .Y(n5932));
  OAI21X1 g02816(.A0(n5035), .A1(n3798), .B0(n5928), .Y(n5933));
  OAI21X1 g02817(.A0(n5032), .A1(n5030), .B0(n5928), .Y(n5934));
  NAND4X1 g02818(.A(n5933), .B(n5932), .C(n5931), .D(n5934), .Y(n5935));
  NOR3X1  g02819(.A(n5935), .B(n5930), .C(n5912), .Y(n5936));
  NAND2X1 g02820(.A(n5936), .B(n5909), .Y(n5937));
  AOI21X1 g02821(.A0(n5904), .A1(n5026), .B0(n5937), .Y(n5938));
  AOI22X1 g02822(.A0(n4983), .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B0(P3_REIP_REG_17__SCAN_IN), .B1(n4968), .Y(n5939));
  OAI21X1 g02823(.A0(n5938), .A1(n4985), .B0(n5939), .Y(P3_U2845));
  AOI21X1 g02824(.A0(n5898), .A1(n5895), .B0(n5518), .Y(n5941));
  AOI21X1 g02825(.A0(n5896), .A1(n5894), .B0(n5941), .Y(n5942));
  INVX1   g02826(.A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .Y(n5943));
  XOR2X1  g02827(.A(n5518), .B(n5943), .Y(n5944));
  XOR2X1  g02828(.A(n5944), .B(n5942), .Y(n5945));
  NOR2X1  g02829(.A(n5945), .B(n5268), .Y(n5946));
  XOR2X1  g02830(.A(n5907), .B(n5943), .Y(n5947));
  NOR2X1  g02831(.A(n5947), .B(n5041), .Y(n5948));
  XOR2X1  g02832(.A(n5911), .B(n5943), .Y(n5949));
  NOR2X1  g02833(.A(n5913), .B(n5895), .Y(n5950));
  XOR2X1  g02834(.A(n5950), .B(n5943), .Y(n5951));
  INVX1   g02835(.A(n5951), .Y(n5952));
  AOI21X1 g02836(.A0(n3861), .A1(n3917), .B0(n5951), .Y(n5953));
  AOI21X1 g02837(.A0(n5952), .A1(n3732), .B0(n5953), .Y(n5954));
  AOI22X1 g02838(.A0(n5952), .A1(n3713), .B0(n5045), .B1(n5963), .Y(n5957));
  OAI21X1 g02839(.A0(n3858), .A1(n3720), .B0(n5952), .Y(n5958));
  NOR4X1  g02840(.A(n5895), .B(n5862), .C(n5839), .D(n5848), .Y(n5959));
  XOR2X1  g02841(.A(n5959), .B(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .Y(n5960));
  NOR3X1  g02842(.A(n5881), .B(n5895), .C(n5862), .Y(n5961));
  XOR2X1  g02843(.A(n5961), .B(n5943), .Y(n5962));
  INVX1   g02844(.A(n5962), .Y(n5963));
  AOI22X1 g02845(.A0(n5960), .A1(n3702), .B0(n3805), .B1(n5963), .Y(n5964));
  NAND4X1 g02846(.A(n5958), .B(n5957), .C(n5954), .D(n5964), .Y(n5965));
  AOI22X1 g02847(.A0(n5960), .A1(n3745), .B0(n5032), .B1(n5963), .Y(n5966));
  OAI21X1 g02848(.A0(n5035), .A1(n3798), .B0(n5963), .Y(n5967));
  NAND2X1 g02849(.A(n5967), .B(n5966), .Y(n5968));
  AOI21X1 g02850(.A0(n5031), .A1(n3835), .B0(n5962), .Y(n5969));
  AOI21X1 g02851(.A0(n5592), .A1(n3786), .B0(n5962), .Y(n5970));
  NOR4X1  g02852(.A(n5969), .B(n5968), .C(n5965), .D(n5970), .Y(n5971));
  OAI21X1 g02853(.A0(n5949), .A1(n3922), .B0(n5971), .Y(n5972));
  NOR3X1  g02854(.A(n5972), .B(n5948), .C(n5946), .Y(n5973));
  AOI22X1 g02855(.A0(n4983), .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B0(P3_REIP_REG_18__SCAN_IN), .B1(n4968), .Y(n5974));
  OAI21X1 g02856(.A0(n5973), .A1(n4985), .B0(n5974), .Y(P3_U2844));
  INVX1   g02857(.A(n5942), .Y(n5976));
  OAI21X1 g02858(.A0(n5570), .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B0(n5976), .Y(n5977));
  OAI21X1 g02859(.A0(n5518), .A1(n5943), .B0(n5977), .Y(n5978));
  XOR2X1  g02860(.A(n5518), .B(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .Y(n5979));
  NOR2X1  g02861(.A(n5978), .B(n5979), .Y(n5980));
  INVX1   g02862(.A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .Y(n5981));
  AOI21X1 g02863(.A0(n5979), .A1(n5978), .B0(n5980), .Y(n5984));
  NOR2X1  g02864(.A(n5984), .B(n5268), .Y(n5985));
  AOI21X1 g02865(.A0(n5907), .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B0(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .Y(n5986));
  NOR4X1  g02866(.A(n5821), .B(n5981), .C(n5943), .D(n5906), .Y(n5987));
  NOR3X1  g02867(.A(n5987), .B(n5986), .C(n5041), .Y(n5988));
  NOR3X1  g02868(.A(n5906), .B(n5831), .C(n5943), .Y(n5989));
  NOR4X1  g02869(.A(n5831), .B(n5981), .C(n5943), .D(n5906), .Y(n5990));
  INVX1   g02870(.A(n5990), .Y(n5991));
  OAI21X1 g02871(.A0(n5989), .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B0(n5991), .Y(n5992));
  NOR2X1  g02872(.A(n5992), .B(n3922), .Y(n5993));
  NOR3X1  g02873(.A(n5913), .B(n5943), .C(n5895), .Y(n5994));
  XOR2X1  g02874(.A(n5994), .B(n5981), .Y(n5995));
  INVX1   g02875(.A(n5995), .Y(n5996));
  OAI21X1 g02876(.A0(n3858), .A1(n3713), .B0(n5996), .Y(n5997));
  OAI21X1 g02877(.A0(n5995), .A1(n3918), .B0(n5997), .Y(n5998));
  OAI22X1 g02878(.A0(n5995), .A1(n3861), .B0(n5593), .B1(n6007), .Y(n6002));
  AOI21X1 g02879(.A0(n3917), .A1(n3920), .B0(n5995), .Y(n6003));
  NAND2X1 g02880(.A(n5959), .B(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .Y(n6004));
  XOR2X1  g02881(.A(n6004), .B(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .Y(n6005));
  NOR4X1  g02882(.A(n5943), .B(n5895), .C(n5862), .D(n5881), .Y(n6006));
  XOR2X1  g02883(.A(n6006), .B(n5981), .Y(n6007));
  OAI22X1 g02884(.A0(n6005), .A1(n3925), .B0(n5043), .B1(n6007), .Y(n6008));
  NOR4X1  g02885(.A(n6003), .B(n6002), .C(n5998), .D(n6008), .Y(n6009));
  AOI21X1 g02886(.A0(n3835), .A1(n3786), .B0(n6007), .Y(n6010));
  OAI22X1 g02887(.A0(n6005), .A1(n3924), .B0(n5592), .B1(n6007), .Y(n6011));
  AOI21X1 g02888(.A0(n5036), .A1(n3797), .B0(n6007), .Y(n6012));
  AOI21X1 g02889(.A0(n5033), .A1(n5031), .B0(n6007), .Y(n6013));
  NOR4X1  g02890(.A(n6012), .B(n6011), .C(n6010), .D(n6013), .Y(n6014));
  NAND2X1 g02891(.A(n6014), .B(n6009), .Y(n6015));
  NOR4X1  g02892(.A(n5993), .B(n5988), .C(n5985), .D(n6015), .Y(n6016));
  AOI22X1 g02893(.A0(n4983), .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B0(P3_REIP_REG_19__SCAN_IN), .B1(n4968), .Y(n6017));
  OAI21X1 g02894(.A0(n6016), .A1(n4985), .B0(n6017), .Y(P3_U2843));
  NOR2X1  g02895(.A(n5518), .B(n5981), .Y(n6019));
  INVX1   g02896(.A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .Y(n6020));
  NOR2X1  g02897(.A(n6020), .B(n5981), .Y(n6021));
  INVX1   g02898(.A(n6021), .Y(n6022));
  NOR2X1  g02899(.A(n5518), .B(n6020), .Y(n6023));
  AOI21X1 g02900(.A0(n6022), .A1(n5518), .B0(n6023), .Y(n6024));
  OAI21X1 g02901(.A0(n6019), .A1(n5978), .B0(n6024), .Y(n6025));
  NOR3X1  g02902(.A(n5978), .B(n6020), .C(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .Y(n6026));
  AOI22X1 g02903(.A0(n5518), .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B0(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B1(n5978), .Y(n6027));
  OAI21X1 g02904(.A0(n6026), .A1(n5518), .B0(n6027), .Y(n6028));
  NAND2X1 g02905(.A(n6028), .B(n6025), .Y(n6029));
  XOR2X1  g02906(.A(n5987), .B(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .Y(n6030));
  XOR2X1  g02907(.A(n5990), .B(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .Y(n6031));
  NAND2X1 g02908(.A(n6031), .B(n3921), .Y(n6032));
  NOR4X1  g02909(.A(n5981), .B(n5943), .C(n5895), .D(n5913), .Y(n6033));
  XOR2X1  g02910(.A(n6033), .B(n6020), .Y(n6034));
  INVX1   g02911(.A(n6034), .Y(n6035));
  OAI21X1 g02912(.A0(n3860), .A1(n3858), .B0(n6035), .Y(n6036));
  OAI21X1 g02913(.A0(n6034), .A1(n3917), .B0(n6036), .Y(n6037));
  OAI22X1 g02914(.A0(n6034), .A1(n3753), .B0(n5593), .B1(n6045), .Y(n6040));
  AOI21X1 g02915(.A0(n3918), .A1(n3920), .B0(n6034), .Y(n6041));
  NAND3X1 g02916(.A(n5959), .B(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .Y(n6042));
  XOR2X1  g02917(.A(n6042), .B(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .Y(n6043));
  NAND2X1 g02918(.A(n6006), .B(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .Y(n6044));
  XOR2X1  g02919(.A(n6044), .B(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .Y(n6045));
  OAI22X1 g02920(.A0(n6043), .A1(n3925), .B0(n5592), .B1(n6045), .Y(n6046));
  NOR4X1  g02921(.A(n6041), .B(n6040), .C(n6037), .D(n6046), .Y(n6047));
  AOI21X1 g02922(.A0(n5033), .A1(n5031), .B0(n6045), .Y(n6048));
  AOI21X1 g02923(.A0(n5036), .A1(n3797), .B0(n6045), .Y(n6049));
  AOI21X1 g02924(.A0(n5043), .A1(n3786), .B0(n6045), .Y(n6050));
  OAI22X1 g02925(.A0(n6043), .A1(n3924), .B0(n3835), .B1(n6045), .Y(n6051));
  NOR4X1  g02926(.A(n6050), .B(n6049), .C(n6048), .D(n6051), .Y(n6052));
  NAND3X1 g02927(.A(n6052), .B(n6047), .C(n6032), .Y(n6053));
  AOI21X1 g02928(.A0(n6030), .A1(n5040), .B0(n6053), .Y(n6054));
  OAI21X1 g02929(.A0(n6029), .A1(n5268), .B0(n6054), .Y(n6055));
  NAND2X1 g02930(.A(n6055), .B(n4984), .Y(n6056));
  AOI22X1 g02931(.A0(n4983), .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B0(P3_REIP_REG_20__SCAN_IN), .B1(n4968), .Y(n6057));
  NAND2X1 g02932(.A(n6057), .B(n6056), .Y(P3_U2842));
  OAI21X1 g02933(.A0(n5978), .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B0(n5570), .Y(n6059));
  AOI21X1 g02934(.A0(n6021), .A1(n5978), .B0(n6023), .Y(n6060));
  NAND2X1 g02935(.A(n6060), .B(n6059), .Y(n6061));
  XOR2X1  g02936(.A(n5518), .B(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .Y(n6062));
  XOR2X1  g02937(.A(n6062), .B(n6061), .Y(n6063));
  NOR2X1  g02938(.A(n6063), .B(n5268), .Y(n6064));
  INVX1   g02939(.A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .Y(n6065));
  NAND2X1 g02940(.A(n5987), .B(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .Y(n6066));
  XOR2X1  g02941(.A(n6066), .B(n6065), .Y(n6067));
  NAND2X1 g02942(.A(n6067), .B(n5040), .Y(n6068));
  OAI21X1 g02943(.A0(n5991), .A1(n6020), .B0(n6065), .Y(n6069));
  NOR3X1  g02944(.A(n5991), .B(n6065), .C(n6020), .Y(n6070));
  INVX1   g02945(.A(n6070), .Y(n6071));
  NAND3X1 g02946(.A(n6071), .B(n6069), .C(n3921), .Y(n6072));
  NAND2X1 g02947(.A(n6033), .B(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .Y(n6073));
  XOR2X1  g02948(.A(n6073), .B(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .Y(n6074));
  INVX1   g02949(.A(n6074), .Y(n6075));
  OAI21X1 g02950(.A0(n3860), .A1(n3858), .B0(n6075), .Y(n6076));
  OAI21X1 g02951(.A0(n6074), .A1(n3753), .B0(n6076), .Y(n6077));
  OAI22X1 g02952(.A0(n6074), .A1(n3917), .B0(n5593), .B1(n6083), .Y(n6080));
  AOI21X1 g02953(.A0(n3918), .A1(n3920), .B0(n6074), .Y(n6081));
  NAND3X1 g02954(.A(n6006), .B(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .C(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .Y(n6082));
  XOR2X1  g02955(.A(n6082), .B(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .Y(n6083));
  AOI21X1 g02956(.A0(n5592), .A1(n5043), .B0(n6083), .Y(n6084));
  NOR4X1  g02957(.A(n6081), .B(n6080), .C(n6077), .D(n6084), .Y(n6085));
  NAND4X1 g02958(.A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .C(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .D(n5959), .Y(n6086));
  XOR2X1  g02959(.A(n6086), .B(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .Y(n6087));
  AOI21X1 g02960(.A0(n3925), .A1(n3924), .B0(n6087), .Y(n6088));
  AOI21X1 g02961(.A0(n3835), .A1(n3786), .B0(n6083), .Y(n6089));
  AOI21X1 g02962(.A0(n5036), .A1(n3797), .B0(n6083), .Y(n6090));
  AOI21X1 g02963(.A0(n5033), .A1(n5031), .B0(n6083), .Y(n6091));
  NOR4X1  g02964(.A(n6090), .B(n6089), .C(n6088), .D(n6091), .Y(n6092));
  NAND4X1 g02965(.A(n6085), .B(n6072), .C(n6068), .D(n6092), .Y(n6093));
  OAI21X1 g02966(.A0(n6093), .A1(n6064), .B0(n4984), .Y(n6094));
  AOI22X1 g02967(.A0(n4983), .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B0(P3_REIP_REG_21__SCAN_IN), .B1(n4968), .Y(n6095));
  NAND2X1 g02968(.A(n6095), .B(n6094), .Y(P3_U2841));
  NOR3X1  g02969(.A(n6065), .B(n6020), .C(n5981), .Y(n6097));
  AOI21X1 g02970(.A0(n6097), .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B0(n5570), .Y(n6098));
  NOR2X1  g02971(.A(n6098), .B(n5942), .Y(n6099));
  NOR2X1  g02972(.A(n5518), .B(n6065), .Y(n6100));
  AOI21X1 g02973(.A0(n5981), .A1(n5943), .B0(n5518), .Y(n6101));
  NOR3X1  g02974(.A(n6101), .B(n6100), .C(n6023), .Y(n6102));
  INVX1   g02975(.A(n6102), .Y(n6103));
  NOR2X1  g02976(.A(n6103), .B(n6099), .Y(n6104));
  XOR2X1  g02977(.A(n5518), .B(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .Y(n6105));
  XOR2X1  g02978(.A(n6105), .B(n6104), .Y(n6106));
  INVX1   g02979(.A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .Y(n6107));
  NOR2X1  g02980(.A(n6066), .B(n6065), .Y(n6108));
  XOR2X1  g02981(.A(n6108), .B(n6107), .Y(n6109));
  XOR2X1  g02982(.A(n6070), .B(n6107), .Y(n6110));
  NOR2X1  g02983(.A(n6110), .B(n3922), .Y(n6111));
  NAND3X1 g02984(.A(n6033), .B(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .C(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .Y(n6112));
  XOR2X1  g02985(.A(n6112), .B(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .Y(n6113));
  INVX1   g02986(.A(n6113), .Y(n6114));
  OAI21X1 g02987(.A0(n3860), .A1(n3713), .B0(n6114), .Y(n6115));
  OAI21X1 g02988(.A0(n6113), .A1(n3859), .B0(n6115), .Y(n6116));
  OAI22X1 g02989(.A0(n6113), .A1(n3917), .B0(n5593), .B1(n6122), .Y(n6119));
  AOI21X1 g02990(.A0(n3918), .A1(n3920), .B0(n6113), .Y(n6120));
  NAND4X1 g02991(.A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .C(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .D(n6006), .Y(n6121));
  XOR2X1  g02992(.A(n6121), .B(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .Y(n6122));
  AOI21X1 g02993(.A0(n5592), .A1(n3786), .B0(n6122), .Y(n6123));
  NOR4X1  g02994(.A(n6120), .B(n6119), .C(n6116), .D(n6123), .Y(n6124));
  NOR2X1  g02995(.A(n6086), .B(n6065), .Y(n6125));
  XOR2X1  g02996(.A(n6125), .B(n6107), .Y(n6126));
  AOI21X1 g02997(.A0(n3925), .A1(n3924), .B0(n6126), .Y(n6127));
  AOI21X1 g02998(.A0(n5033), .A1(n5031), .B0(n6122), .Y(n6128));
  AOI21X1 g02999(.A0(n3835), .A1(n3797), .B0(n6122), .Y(n6129));
  AOI21X1 g03000(.A0(n5036), .A1(n5043), .B0(n6122), .Y(n6130));
  NOR4X1  g03001(.A(n6129), .B(n6128), .C(n6127), .D(n6130), .Y(n6131));
  NAND2X1 g03002(.A(n6131), .B(n6124), .Y(n6132));
  NOR2X1  g03003(.A(n6132), .B(n6111), .Y(n6133));
  OAI21X1 g03004(.A0(n6109), .A1(n5041), .B0(n6133), .Y(n6134));
  AOI21X1 g03005(.A0(n6106), .A1(n5026), .B0(n6134), .Y(n6135));
  AOI22X1 g03006(.A0(n4983), .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B0(P3_REIP_REG_22__SCAN_IN), .B1(n4968), .Y(n6136));
  OAI21X1 g03007(.A0(n6135), .A1(n4985), .B0(n6136), .Y(P3_U2840));
  AOI21X1 g03008(.A0(n5518), .A1(n6107), .B0(n6098), .Y(n6138));
  AOI21X1 g03009(.A0(n5570), .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B0(n6103), .Y(n6139));
  INVX1   g03010(.A(n6139), .Y(n6140));
  AOI21X1 g03011(.A0(n6138), .A1(n5976), .B0(n6140), .Y(n6141));
  XOR2X1  g03012(.A(n5518), .B(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .Y(n6142));
  XOR2X1  g03013(.A(n6142), .B(n6141), .Y(n6143));
  INVX1   g03014(.A(n6143), .Y(n6144));
  NOR2X1  g03015(.A(n6144), .B(n5268), .Y(n6145));
  NOR3X1  g03016(.A(n6066), .B(n6107), .C(n6065), .Y(n6146));
  INVX1   g03017(.A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .Y(n6147));
  NOR4X1  g03018(.A(n6147), .B(n6107), .C(n6065), .D(n6066), .Y(n6148));
  INVX1   g03019(.A(n6148), .Y(n6149));
  OAI21X1 g03020(.A0(n6146), .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B0(n6149), .Y(n6150));
  NOR2X1  g03021(.A(n6150), .B(n5041), .Y(n6151));
  OAI21X1 g03022(.A0(n6071), .A1(n6107), .B0(n6147), .Y(n6152));
  NOR3X1  g03023(.A(n6071), .B(n6147), .C(n6107), .Y(n6153));
  INVX1   g03024(.A(n6153), .Y(n6154));
  NAND3X1 g03025(.A(n6154), .B(n6152), .C(n3921), .Y(n6155));
  NAND4X1 g03026(.A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .C(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .D(n6033), .Y(n6156));
  XOR2X1  g03027(.A(n6156), .B(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .Y(n6157));
  INVX1   g03028(.A(n6157), .Y(n6158));
  OAI21X1 g03029(.A0(n3860), .A1(n3713), .B0(n6158), .Y(n6159));
  OAI21X1 g03030(.A0(n6157), .A1(n3859), .B0(n6159), .Y(n6160));
  OAI22X1 g03031(.A0(n6157), .A1(n3917), .B0(n5593), .B1(n6166), .Y(n6163));
  AOI21X1 g03032(.A0(n3918), .A1(n3920), .B0(n6157), .Y(n6164));
  NOR2X1  g03033(.A(n6121), .B(n6107), .Y(n6165));
  XOR2X1  g03034(.A(n6165), .B(n6147), .Y(n6166));
  AOI21X1 g03035(.A0(n5592), .A1(n3786), .B0(n6166), .Y(n6167));
  NOR4X1  g03036(.A(n6164), .B(n6163), .C(n6160), .D(n6167), .Y(n6168));
  NOR3X1  g03037(.A(n6086), .B(n6107), .C(n6065), .Y(n6169));
  XOR2X1  g03038(.A(n6169), .B(n6147), .Y(n6170));
  AOI21X1 g03039(.A0(n3925), .A1(n3924), .B0(n6170), .Y(n6171));
  AOI21X1 g03040(.A0(n5033), .A1(n5031), .B0(n6166), .Y(n6172));
  AOI21X1 g03041(.A0(n3835), .A1(n3797), .B0(n6166), .Y(n6173));
  AOI21X1 g03042(.A0(n5036), .A1(n5043), .B0(n6166), .Y(n6174));
  NOR4X1  g03043(.A(n6173), .B(n6172), .C(n6171), .D(n6174), .Y(n6175));
  NAND3X1 g03044(.A(n6175), .B(n6168), .C(n6155), .Y(n6176));
  NOR3X1  g03045(.A(n6176), .B(n6151), .C(n6145), .Y(n6177));
  AOI22X1 g03046(.A0(n4983), .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B0(P3_REIP_REG_23__SCAN_IN), .B1(n4968), .Y(n6178));
  OAI21X1 g03047(.A0(n6177), .A1(n4985), .B0(n6178), .Y(P3_U2839));
  OAI21X1 g03048(.A0(n5570), .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B0(n6138), .Y(n6180));
  NOR2X1  g03049(.A(n6180), .B(n5942), .Y(n6181));
  AOI21X1 g03050(.A0(n5570), .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B0(n6140), .Y(n6182));
  INVX1   g03051(.A(n6182), .Y(n6183));
  NOR2X1  g03052(.A(n6183), .B(n6181), .Y(n6184));
  XOR2X1  g03053(.A(n5518), .B(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .Y(n6185));
  XOR2X1  g03054(.A(n6185), .B(n6184), .Y(n6186));
  XOR2X1  g03055(.A(n6148), .B(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .Y(n6187));
  NAND2X1 g03056(.A(n6187), .B(n5040), .Y(n6188));
  INVX1   g03057(.A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .Y(n6189));
  XOR2X1  g03058(.A(n6153), .B(n6189), .Y(n6190));
  INVX1   g03059(.A(n6190), .Y(n6191));
  NAND2X1 g03060(.A(n6191), .B(n3921), .Y(n6192));
  NOR2X1  g03061(.A(n6156), .B(n6147), .Y(n6193));
  XOR2X1  g03062(.A(n6193), .B(n6189), .Y(n6194));
  INVX1   g03063(.A(n6194), .Y(n6195));
  OAI21X1 g03064(.A0(n3729), .A1(n3713), .B0(n6195), .Y(n6196));
  OAI21X1 g03065(.A0(n6194), .A1(n3861), .B0(n6196), .Y(n6197));
  OAI22X1 g03066(.A0(n6194), .A1(n3859), .B0(n5593), .B1(n6203), .Y(n6200));
  AOI21X1 g03067(.A0(n3918), .A1(n3920), .B0(n6194), .Y(n6201));
  NOR3X1  g03068(.A(n6121), .B(n6147), .C(n6107), .Y(n6202));
  XOR2X1  g03069(.A(n6202), .B(n6189), .Y(n6203));
  AOI21X1 g03070(.A0(n5592), .A1(n3797), .B0(n6203), .Y(n6204));
  NOR4X1  g03071(.A(n6201), .B(n6200), .C(n6197), .D(n6204), .Y(n6205));
  NOR4X1  g03072(.A(n6147), .B(n6107), .C(n6065), .D(n6086), .Y(n6206));
  XOR2X1  g03073(.A(n6206), .B(n6189), .Y(n6207));
  OAI22X1 g03074(.A0(n6203), .A1(n5031), .B0(n3925), .B1(n6207), .Y(n6208));
  OAI22X1 g03075(.A0(n6203), .A1(n5036), .B0(n3924), .B1(n6207), .Y(n6209));
  AOI21X1 g03076(.A0(n3835), .A1(n3786), .B0(n6203), .Y(n6210));
  AOI21X1 g03077(.A0(n5033), .A1(n5043), .B0(n6203), .Y(n6211));
  NOR4X1  g03078(.A(n6210), .B(n6209), .C(n6208), .D(n6211), .Y(n6212));
  NAND4X1 g03079(.A(n6205), .B(n6192), .C(n6188), .D(n6212), .Y(n6213));
  AOI21X1 g03080(.A0(n6186), .A1(n5026), .B0(n6213), .Y(n6214));
  AOI22X1 g03081(.A0(n4983), .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B0(P3_REIP_REG_24__SCAN_IN), .B1(n4968), .Y(n6215));
  OAI21X1 g03082(.A0(n6214), .A1(n4985), .B0(n6215), .Y(P3_U2838));
  XOR2X1  g03083(.A(n5518), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Y(n6217));
  AOI21X1 g03084(.A0(n5518), .A1(n6189), .B0(n6180), .Y(n6218));
  AOI21X1 g03085(.A0(n5570), .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B0(n6183), .Y(n6219));
  INVX1   g03086(.A(n6219), .Y(n6220));
  AOI21X1 g03087(.A0(n6218), .A1(n5976), .B0(n6220), .Y(n6221));
  INVX1   g03088(.A(n6221), .Y(n6222));
  NOR3X1  g03089(.A(n5471), .B(n5413), .C(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Y(n6223));
  INVX1   g03090(.A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Y(n6224));
  NOR2X1  g03091(.A(n5518), .B(n6224), .Y(n6225));
  OAI21X1 g03092(.A0(n6225), .A1(n6223), .B0(n6222), .Y(n6226));
  OAI21X1 g03093(.A0(n6222), .A1(n6217), .B0(n6226), .Y(n6227));
  AOI21X1 g03094(.A0(n6148), .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B0(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Y(n6228));
  NOR3X1  g03095(.A(n6149), .B(n6224), .C(n6189), .Y(n6229));
  NOR2X1  g03096(.A(n6229), .B(n6228), .Y(n6230));
  NAND2X1 g03097(.A(n6230), .B(n5040), .Y(n6231));
  AOI21X1 g03098(.A0(n6153), .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B0(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Y(n6232));
  NOR3X1  g03099(.A(n6154), .B(n6224), .C(n6189), .Y(n6233));
  NOR2X1  g03100(.A(n6233), .B(n6232), .Y(n6234));
  NAND2X1 g03101(.A(n6234), .B(n3921), .Y(n6235));
  NOR3X1  g03102(.A(n6156), .B(n6189), .C(n6147), .Y(n6236));
  XOR2X1  g03103(.A(n6236), .B(n6224), .Y(n6237));
  INVX1   g03104(.A(n6237), .Y(n6238));
  OAI21X1 g03105(.A0(n3729), .A1(n3713), .B0(n6238), .Y(n6239));
  OAI21X1 g03106(.A0(n6237), .A1(n3861), .B0(n6239), .Y(n6240));
  OAI22X1 g03107(.A0(n6237), .A1(n3859), .B0(n5593), .B1(n6246), .Y(n6243));
  AOI21X1 g03108(.A0(n3918), .A1(n3920), .B0(n6237), .Y(n6244));
  NOR4X1  g03109(.A(n6189), .B(n6147), .C(n6107), .D(n6121), .Y(n6245));
  XOR2X1  g03110(.A(n6245), .B(n6224), .Y(n6246));
  AOI21X1 g03111(.A0(n5592), .A1(n3835), .B0(n6246), .Y(n6247));
  NOR4X1  g03112(.A(n6244), .B(n6243), .C(n6240), .D(n6247), .Y(n6248));
  NAND2X1 g03113(.A(n6206), .B(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .Y(n6249));
  XOR2X1  g03114(.A(n6249), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Y(n6250));
  OAI22X1 g03115(.A0(n6246), .A1(n5031), .B0(n3925), .B1(n6250), .Y(n6251));
  OAI22X1 g03116(.A0(n6246), .A1(n5036), .B0(n3924), .B1(n6250), .Y(n6252));
  AOI21X1 g03117(.A0(n5043), .A1(n3786), .B0(n6246), .Y(n6253));
  AOI21X1 g03118(.A0(n5033), .A1(n3797), .B0(n6246), .Y(n6254));
  NOR4X1  g03119(.A(n6253), .B(n6252), .C(n6251), .D(n6254), .Y(n6255));
  NAND4X1 g03120(.A(n6248), .B(n6235), .C(n6231), .D(n6255), .Y(n6256));
  AOI21X1 g03121(.A0(n6227), .A1(n5026), .B0(n6256), .Y(n6257));
  AOI22X1 g03122(.A0(n4983), .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B0(P3_REIP_REG_25__SCAN_IN), .B1(n4968), .Y(n6258));
  OAI21X1 g03123(.A0(n6257), .A1(n4985), .B0(n6258), .Y(P3_U2837));
  INVX1   g03124(.A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .Y(n6260));
  NOR2X1  g03125(.A(n5518), .B(n6260), .Y(n6261));
  AOI21X1 g03126(.A0(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B0(n5570), .Y(n6262));
  NOR2X1  g03127(.A(n6262), .B(n6261), .Y(n6263));
  OAI21X1 g03128(.A0(n6225), .A1(n6222), .B0(n6263), .Y(n6264));
  NOR2X1  g03129(.A(n6223), .B(n6221), .Y(n6265));
  OAI22X1 g03130(.A0(n5413), .A1(n5471), .B0(n6260), .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Y(n6266));
  OAI21X1 g03131(.A0(n5570), .A1(n6260), .B0(n6266), .Y(n6267));
  OAI21X1 g03132(.A0(n6267), .A1(n6265), .B0(n6264), .Y(n6268));
  NOR2X1  g03133(.A(n6268), .B(n5268), .Y(n6269));
  XOR2X1  g03134(.A(n6229), .B(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .Y(n6270));
  NAND2X1 g03135(.A(n6270), .B(n5040), .Y(n6271));
  XOR2X1  g03136(.A(n6233), .B(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .Y(n6272));
  NAND2X1 g03137(.A(n6272), .B(n3921), .Y(n6273));
  NOR4X1  g03138(.A(n6224), .B(n6189), .C(n6147), .D(n6156), .Y(n6274));
  XOR2X1  g03139(.A(n6274), .B(n6260), .Y(n6275));
  INVX1   g03140(.A(n6275), .Y(n6276));
  OAI21X1 g03141(.A0(n3729), .A1(n3713), .B0(n6276), .Y(n6277));
  OAI21X1 g03142(.A0(n6275), .A1(n3861), .B0(n6277), .Y(n6278));
  OAI22X1 g03143(.A0(n6275), .A1(n3859), .B0(n5593), .B1(n6284), .Y(n6281));
  AOI21X1 g03144(.A0(n3918), .A1(n3920), .B0(n6275), .Y(n6282));
  NAND2X1 g03145(.A(n6245), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Y(n6283));
  XOR2X1  g03146(.A(n6283), .B(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .Y(n6284));
  AOI21X1 g03147(.A0(n5592), .A1(n3835), .B0(n6284), .Y(n6285));
  NOR4X1  g03148(.A(n6282), .B(n6281), .C(n6278), .D(n6285), .Y(n6286));
  NAND3X1 g03149(.A(n6206), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .C(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .Y(n6287));
  XOR2X1  g03150(.A(n6287), .B(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .Y(n6288));
  OAI22X1 g03151(.A0(n6284), .A1(n5031), .B0(n3925), .B1(n6288), .Y(n6289));
  OAI22X1 g03152(.A0(n6284), .A1(n5036), .B0(n3924), .B1(n6288), .Y(n6290));
  AOI21X1 g03153(.A0(n5043), .A1(n3786), .B0(n6284), .Y(n6291));
  AOI21X1 g03154(.A0(n5033), .A1(n3797), .B0(n6284), .Y(n6292));
  NOR4X1  g03155(.A(n6291), .B(n6290), .C(n6289), .D(n6292), .Y(n6293));
  NAND4X1 g03156(.A(n6286), .B(n6273), .C(n6271), .D(n6293), .Y(n6294));
  OAI21X1 g03157(.A0(n6294), .A1(n6269), .B0(n4984), .Y(n6295));
  AOI22X1 g03158(.A0(n4983), .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B0(P3_REIP_REG_26__SCAN_IN), .B1(n4968), .Y(n6296));
  NAND2X1 g03159(.A(n6296), .B(n6295), .Y(P3_U2836));
  NOR2X1  g03160(.A(n6262), .B(n6221), .Y(n6298));
  NOR3X1  g03161(.A(n6298), .B(n6261), .C(n6225), .Y(n6299));
  INVX1   g03162(.A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .Y(n6300));
  XOR2X1  g03163(.A(n5518), .B(n6300), .Y(n6301));
  XOR2X1  g03164(.A(n6301), .B(n6299), .Y(n6302));
  NOR2X1  g03165(.A(n6302), .B(n5268), .Y(n6303));
  NOR4X1  g03166(.A(n6260), .B(n6224), .C(n6189), .D(n6149), .Y(n6304));
  XOR2X1  g03167(.A(n6304), .B(n6300), .Y(n6305));
  NOR2X1  g03168(.A(n6305), .B(n5041), .Y(n6306));
  NOR4X1  g03169(.A(n6260), .B(n6224), .C(n6189), .D(n6154), .Y(n6307));
  XOR2X1  g03170(.A(n6307), .B(n6300), .Y(n6308));
  NOR2X1  g03171(.A(n6308), .B(n3922), .Y(n6309));
  NAND2X1 g03172(.A(n6274), .B(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .Y(n6310));
  XOR2X1  g03173(.A(n6310), .B(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .Y(n6311));
  INVX1   g03174(.A(n6311), .Y(n6312));
  OAI21X1 g03175(.A0(n3729), .A1(n3713), .B0(n6312), .Y(n6313));
  OAI21X1 g03176(.A0(n6311), .A1(n3861), .B0(n6313), .Y(n6314));
  OAI22X1 g03177(.A0(n6311), .A1(n3859), .B0(n5593), .B1(n6320), .Y(n6317));
  AOI21X1 g03178(.A0(n3918), .A1(n3920), .B0(n6311), .Y(n6318));
  NAND3X1 g03179(.A(n6245), .B(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .C(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Y(n6319));
  XOR2X1  g03180(.A(n6319), .B(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .Y(n6320));
  AOI21X1 g03181(.A0(n5592), .A1(n3835), .B0(n6320), .Y(n6321));
  NOR4X1  g03182(.A(n6318), .B(n6317), .C(n6314), .D(n6321), .Y(n6322));
  NAND4X1 g03183(.A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .C(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .D(n6206), .Y(n6323));
  XOR2X1  g03184(.A(n6323), .B(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .Y(n6324));
  OAI22X1 g03185(.A0(n6320), .A1(n5031), .B0(n3925), .B1(n6324), .Y(n6325));
  OAI22X1 g03186(.A0(n6320), .A1(n5036), .B0(n3924), .B1(n6324), .Y(n6326));
  AOI21X1 g03187(.A0(n5043), .A1(n3786), .B0(n6320), .Y(n6327));
  AOI21X1 g03188(.A0(n5033), .A1(n3797), .B0(n6320), .Y(n6328));
  NOR4X1  g03189(.A(n6327), .B(n6326), .C(n6325), .D(n6328), .Y(n6329));
  NAND2X1 g03190(.A(n6329), .B(n6322), .Y(n6330));
  NOR4X1  g03191(.A(n6309), .B(n6306), .C(n6303), .D(n6330), .Y(n6331));
  AOI22X1 g03192(.A0(n4983), .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B0(P3_REIP_REG_27__SCAN_IN), .B1(n4968), .Y(n6332));
  OAI21X1 g03193(.A0(n6331), .A1(n4985), .B0(n6332), .Y(P3_U2835));
  NAND2X1 g03194(.A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .Y(n6334));
  NOR2X1  g03195(.A(n6334), .B(n6299), .Y(n6335));
  NOR2X1  g03196(.A(n6335), .B(n5570), .Y(n6336));
  INVX1   g03197(.A(n6336), .Y(n6337));
  NOR4X1  g03198(.A(n6261), .B(n6225), .C(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .D(n6298), .Y(n6338));
  AOI21X1 g03199(.A0(n5570), .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B0(n6338), .Y(n6339));
  AOI21X1 g03200(.A0(n6338), .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B0(n5518), .Y(n6340));
  NOR2X1  g03201(.A(n6299), .B(n6300), .Y(n6341));
  INVX1   g03202(.A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .Y(n6342));
  NOR3X1  g03203(.A(n5471), .B(n5413), .C(n6342), .Y(n6343));
  NOR3X1  g03204(.A(n6343), .B(n6341), .C(n6340), .Y(n6344));
  AOI21X1 g03205(.A0(n6339), .A1(n6337), .B0(n6344), .Y(n6345));
  INVX1   g03206(.A(n6304), .Y(n6346));
  NOR2X1  g03207(.A(n6346), .B(n6300), .Y(n6347));
  OAI22X1 g03208(.A0(n6334), .A1(n6346), .B0(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B1(n6347), .Y(n6348));
  AOI21X1 g03209(.A0(n6307), .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B0(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .Y(n6349));
  INVX1   g03210(.A(n6307), .Y(n6350));
  NOR2X1  g03211(.A(n6334), .B(n6350), .Y(n6351));
  NOR3X1  g03212(.A(n6351), .B(n6349), .C(n3922), .Y(n6352));
  NAND3X1 g03213(.A(n6274), .B(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .C(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .Y(n6353));
  XOR2X1  g03214(.A(n6353), .B(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .Y(n6354));
  INVX1   g03215(.A(n6354), .Y(n6355));
  OAI21X1 g03216(.A0(n3729), .A1(n3713), .B0(n6355), .Y(n6356));
  OAI21X1 g03217(.A0(n6354), .A1(n3861), .B0(n6356), .Y(n6357));
  OAI22X1 g03218(.A0(n6354), .A1(n3859), .B0(n5593), .B1(n6363), .Y(n6360));
  AOI21X1 g03219(.A0(n3918), .A1(n3920), .B0(n6354), .Y(n6361));
  NAND4X1 g03220(.A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .C(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .D(n6245), .Y(n6362));
  XOR2X1  g03221(.A(n6362), .B(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .Y(n6363));
  AOI21X1 g03222(.A0(n5592), .A1(n3835), .B0(n6363), .Y(n6364));
  NOR4X1  g03223(.A(n6361), .B(n6360), .C(n6357), .D(n6364), .Y(n6365));
  NOR2X1  g03224(.A(n6323), .B(n6300), .Y(n6366));
  XOR2X1  g03225(.A(n6366), .B(n6342), .Y(n6367));
  OAI22X1 g03226(.A0(n6363), .A1(n5031), .B0(n3925), .B1(n6367), .Y(n6368));
  OAI22X1 g03227(.A0(n6363), .A1(n5036), .B0(n3924), .B1(n6367), .Y(n6369));
  AOI21X1 g03228(.A0(n5043), .A1(n3786), .B0(n6363), .Y(n6370));
  AOI21X1 g03229(.A0(n5033), .A1(n3797), .B0(n6363), .Y(n6371));
  NOR4X1  g03230(.A(n6370), .B(n6369), .C(n6368), .D(n6371), .Y(n6372));
  NAND2X1 g03231(.A(n6372), .B(n6365), .Y(n6373));
  NOR2X1  g03232(.A(n6373), .B(n6352), .Y(n6374));
  OAI21X1 g03233(.A0(n6348), .A1(n5041), .B0(n6374), .Y(n6375));
  AOI21X1 g03234(.A0(n6345), .A1(n5026), .B0(n6375), .Y(n6376));
  AOI22X1 g03235(.A0(n4983), .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B0(P3_REIP_REG_28__SCAN_IN), .B1(n4968), .Y(n6377));
  OAI21X1 g03236(.A0(n6376), .A1(n4985), .B0(n6377), .Y(P3_U2834));
  NOR2X1  g03237(.A(n6338), .B(n5518), .Y(n6379));
  OAI22X1 g03238(.A0(n6299), .A1(n6334), .B0(n5518), .B1(n6342), .Y(n6380));
  NOR2X1  g03239(.A(n6380), .B(n6379), .Y(n6381));
  INVX1   g03240(.A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .Y(n6382));
  XOR2X1  g03241(.A(n5518), .B(n6382), .Y(n6383));
  XOR2X1  g03242(.A(n6383), .B(n6381), .Y(n6384));
  NOR2X1  g03243(.A(n6384), .B(n5268), .Y(n6385));
  NAND3X1 g03244(.A(n6304), .B(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .C(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .Y(n6386));
  XOR2X1  g03245(.A(n6386), .B(n6382), .Y(n6387));
  NAND2X1 g03246(.A(n6387), .B(n5040), .Y(n6388));
  XOR2X1  g03247(.A(n6351), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .Y(n6389));
  NAND2X1 g03248(.A(n6389), .B(n3921), .Y(n6390));
  NAND4X1 g03249(.A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .C(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .D(n6274), .Y(n6391));
  XOR2X1  g03250(.A(n6391), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .Y(n6392));
  INVX1   g03251(.A(n6392), .Y(n6393));
  OAI21X1 g03252(.A0(n3729), .A1(n3713), .B0(n6393), .Y(n6394));
  OAI21X1 g03253(.A0(n6392), .A1(n3861), .B0(n6394), .Y(n6395));
  OAI22X1 g03254(.A0(n6392), .A1(n3859), .B0(n5593), .B1(n6401), .Y(n6398));
  AOI21X1 g03255(.A0(n3918), .A1(n3920), .B0(n6392), .Y(n6399));
  NOR2X1  g03256(.A(n6362), .B(n6342), .Y(n6400));
  XOR2X1  g03257(.A(n6400), .B(n6382), .Y(n6401));
  AOI21X1 g03258(.A0(n5592), .A1(n3835), .B0(n6401), .Y(n6402));
  NOR4X1  g03259(.A(n6399), .B(n6398), .C(n6395), .D(n6402), .Y(n6403));
  NOR3X1  g03260(.A(n6323), .B(n6342), .C(n6300), .Y(n6404));
  XOR2X1  g03261(.A(n6404), .B(n6382), .Y(n6405));
  OAI22X1 g03262(.A0(n6401), .A1(n5031), .B0(n3925), .B1(n6405), .Y(n6406));
  OAI22X1 g03263(.A0(n6401), .A1(n5036), .B0(n3924), .B1(n6405), .Y(n6407));
  AOI21X1 g03264(.A0(n5043), .A1(n3786), .B0(n6401), .Y(n6408));
  AOI21X1 g03265(.A0(n5033), .A1(n3797), .B0(n6401), .Y(n6409));
  NOR4X1  g03266(.A(n6408), .B(n6407), .C(n6406), .D(n6409), .Y(n6410));
  NAND4X1 g03267(.A(n6403), .B(n6390), .C(n6388), .D(n6410), .Y(n6411));
  OAI21X1 g03268(.A0(n6411), .A1(n6385), .B0(n4984), .Y(n6412));
  AOI22X1 g03269(.A0(n4983), .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B0(P3_REIP_REG_29__SCAN_IN), .B1(n4968), .Y(n6413));
  NAND2X1 g03270(.A(n6413), .B(n6412), .Y(P3_U2833));
  XOR2X1  g03271(.A(n5518), .B(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .Y(n6415));
  INVX1   g03272(.A(n6415), .Y(n6416));
  NOR2X1  g03273(.A(n6381), .B(n6382), .Y(n6417));
  NOR2X1  g03274(.A(n5518), .B(n6382), .Y(n6418));
  NOR2X1  g03275(.A(n6381), .B(n5518), .Y(n6419));
  NOR3X1  g03276(.A(n6419), .B(n6418), .C(n6417), .Y(n6420));
  XOR2X1  g03277(.A(n6420), .B(n6416), .Y(n6421));
  NOR2X1  g03278(.A(n6421), .B(n5268), .Y(n6422));
  NAND4X1 g03279(.A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .C(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .D(n6304), .Y(n6423));
  XOR2X1  g03280(.A(n6423), .B(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .Y(n6424));
  NOR2X1  g03281(.A(n6424), .B(n5041), .Y(n6425));
  INVX1   g03282(.A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .Y(n6426));
  NOR3X1  g03283(.A(n6334), .B(n6350), .C(n6382), .Y(n6427));
  XOR2X1  g03284(.A(n6427), .B(n6426), .Y(n6428));
  NOR2X1  g03285(.A(n6428), .B(n3922), .Y(n6429));
  NOR2X1  g03286(.A(n6391), .B(n6382), .Y(n6430));
  XOR2X1  g03287(.A(n6430), .B(n6426), .Y(n6431));
  INVX1   g03288(.A(n6431), .Y(n6432));
  OAI21X1 g03289(.A0(n3729), .A1(n3713), .B0(n6432), .Y(n6433));
  OAI21X1 g03290(.A0(n6431), .A1(n3861), .B0(n6433), .Y(n6434));
  OAI22X1 g03291(.A0(n6431), .A1(n3859), .B0(n5593), .B1(n6440), .Y(n6437));
  AOI21X1 g03292(.A0(n3918), .A1(n3920), .B0(n6431), .Y(n6438));
  NOR3X1  g03293(.A(n6362), .B(n6382), .C(n6342), .Y(n6439));
  XOR2X1  g03294(.A(n6439), .B(n6426), .Y(n6440));
  AOI21X1 g03295(.A0(n5592), .A1(n3835), .B0(n6440), .Y(n6441));
  NOR4X1  g03296(.A(n6438), .B(n6437), .C(n6434), .D(n6441), .Y(n6442));
  NOR4X1  g03297(.A(n6382), .B(n6342), .C(n6300), .D(n6323), .Y(n6443));
  XOR2X1  g03298(.A(n6443), .B(n6426), .Y(n6444));
  OAI22X1 g03299(.A0(n6440), .A1(n5031), .B0(n3925), .B1(n6444), .Y(n6445));
  OAI22X1 g03300(.A0(n6440), .A1(n5036), .B0(n3924), .B1(n6444), .Y(n6446));
  AOI21X1 g03301(.A0(n5043), .A1(n3786), .B0(n6440), .Y(n6447));
  AOI21X1 g03302(.A0(n5033), .A1(n3797), .B0(n6440), .Y(n6448));
  NOR4X1  g03303(.A(n6447), .B(n6446), .C(n6445), .D(n6448), .Y(n6449));
  NAND2X1 g03304(.A(n6449), .B(n6442), .Y(n6450));
  NOR4X1  g03305(.A(n6429), .B(n6425), .C(n6422), .D(n6450), .Y(n6451));
  AOI22X1 g03306(.A0(n4983), .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B0(P3_REIP_REG_30__SCAN_IN), .B1(n4968), .Y(n6452));
  OAI21X1 g03307(.A0(n6451), .A1(n4985), .B0(n6452), .Y(P3_U2832));
  NOR2X1  g03308(.A(n3961), .B(n6426), .Y(n6454));
  INVX1   g03309(.A(n6454), .Y(n6455));
  OAI21X1 g03310(.A0(n6455), .A1(n6420), .B0(n5518), .Y(n6456));
  AOI22X1 g03311(.A0(n5570), .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B0(n6426), .B1(n6420), .Y(n6457));
  NOR2X1  g03312(.A(n6420), .B(n6426), .Y(n6458));
  INVX1   g03313(.A(n6458), .Y(n6459));
  NOR3X1  g03314(.A(n6418), .B(n3961), .C(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .Y(n6460));
  AOI21X1 g03315(.A0(n6460), .A1(n6381), .B0(n5518), .Y(n6461));
  AOI21X1 g03316(.A0(n5518), .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B0(n6461), .Y(n6462));
  AOI22X1 g03317(.A0(n6459), .A1(n6462), .B0(n6457), .B1(n6456), .Y(n6463));
  NAND2X1 g03318(.A(n6463), .B(n5026), .Y(n6464));
  NOR2X1  g03319(.A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n6426), .Y(n6465));
  INVX1   g03320(.A(n6465), .Y(n6466));
  OAI21X1 g03321(.A0(n6423), .A1(n6426), .B0(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .Y(n6467));
  OAI21X1 g03322(.A0(n6466), .A1(n6423), .B0(n6467), .Y(n6468));
  AOI21X1 g03323(.A0(n6427), .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B0(n3961), .Y(n6469));
  AOI21X1 g03324(.A0(n6465), .A1(n6427), .B0(n6469), .Y(n6470));
  NOR3X1  g03325(.A(n6391), .B(n6426), .C(n6382), .Y(n6471));
  XOR2X1  g03326(.A(n6471), .B(n3961), .Y(n6472));
  INVX1   g03327(.A(n6472), .Y(n6473));
  OAI21X1 g03328(.A0(n3858), .A1(n3732), .B0(n6473), .Y(n6474));
  OAI21X1 g03329(.A0(n6472), .A1(n3753), .B0(n6474), .Y(n6475));
  NAND2X1 g03330(.A(n6473), .B(n3729), .Y(n6476));
  INVX1   g03331(.A(P3_REIP_REG_31__SCAN_IN), .Y(n6477));
  NOR2X1  g03332(.A(n4969), .B(n6477), .Y(n6478));
  OAI22X1 g03333(.A0(n5593), .A1(n6485), .B0(n4982), .B1(n3961), .Y(n6481));
  NOR2X1  g03334(.A(n6481), .B(n6478), .Y(n6482));
  OAI21X1 g03335(.A0(n3860), .A1(n3720), .B0(n6473), .Y(n6483));
  NOR4X1  g03336(.A(n6426), .B(n6382), .C(n6342), .D(n6362), .Y(n6484));
  XOR2X1  g03337(.A(n6484), .B(n3961), .Y(n6485));
  INVX1   g03338(.A(n6485), .Y(n6486));
  OAI21X1 g03339(.A0(n5044), .A1(n3787), .B0(n6486), .Y(n6487));
  NAND4X1 g03340(.A(n6483), .B(n6482), .C(n6476), .D(n6487), .Y(n6488));
  OAI21X1 g03341(.A0(n5035), .A1(n3798), .B0(n6486), .Y(n6489));
  NAND2X1 g03342(.A(n6443), .B(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .Y(n6490));
  XOR2X1  g03343(.A(n6490), .B(n3961), .Y(n6491));
  AOI22X1 g03344(.A0(n6486), .A1(n5032), .B0(n3702), .B1(n6491), .Y(n6492));
  OAI21X1 g03345(.A0(n3834), .A1(n3805), .B0(n6486), .Y(n6493));
  AOI22X1 g03346(.A0(n6486), .A1(n5030), .B0(n3745), .B1(n6491), .Y(n6494));
  NAND4X1 g03347(.A(n6493), .B(n6492), .C(n6489), .D(n6494), .Y(n6495));
  NOR3X1  g03348(.A(n6495), .B(n6488), .C(n6475), .Y(n6496));
  OAI21X1 g03349(.A0(n6470), .A1(n3922), .B0(n6496), .Y(n6497));
  AOI21X1 g03350(.A0(n6468), .A1(n5040), .B0(n6497), .Y(n6498));
  NOR2X1  g03351(.A(n4982), .B(n3961), .Y(n6499));
  NOR3X1  g03352(.A(n6499), .B(n6478), .C(n4984), .Y(n6500));
  AOI21X1 g03353(.A0(n6498), .A1(n6464), .B0(n6500), .Y(P3_U2831));
  NOR2X1  g03354(.A(n4073), .B(n3949), .Y(n6502));
  AOI22X1 g03355(.A0(n3914), .A1(n3890), .B0(n3893), .B1(n3921), .Y(n6503));
  OAI22X1 g03356(.A0(n6502), .A1(P3_STATE2_REG_0__SCAN_IN), .B0(n4905), .B1(n6503), .Y(n6504));
  INVX1   g03357(.A(n6504), .Y(n6505));
  AOI22X1 g03358(.A0(n6505), .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B0(P3_REIP_REG_0__SCAN_IN), .B1(n4968), .Y(n6507));
  NOR4X1  g03359(.A(P3_STATE2_REG_1__SCAN_IN), .B(n3511), .C(P3_STATE2_REG_3__SCAN_IN), .D(P3_STATE2_REG_0__SCAN_IN), .Y(n6508));
  NOR3X1  g03360(.A(n6505), .B(n3682), .C(n3510), .Y(n6509));
  AOI22X1 g03361(.A0(n6508), .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B0(n5013), .B1(n6509), .Y(n6510));
  NOR3X1  g03362(.A(n6505), .B(P3_STATEBS16_REG_SCAN_IN), .C(n3939), .Y(n6511));
  NOR4X1  g03363(.A(n5025), .B(n3681), .C(n3510), .D(n6505), .Y(n6512));
  AOI22X1 g03364(.A0(n6511), .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B0(n5014), .B1(n6512), .Y(n6513));
  NOR3X1  g03365(.A(n6505), .B(n3944), .C(n3939), .Y(n6514));
  NOR4X1  g03366(.A(n5039), .B(n3681), .C(n3510), .D(n6505), .Y(n6515));
  AOI22X1 g03367(.A0(n6514), .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B0(n5014), .B1(n6515), .Y(n6516));
  NAND4X1 g03368(.A(n6513), .B(n6510), .C(n6507), .D(n6516), .Y(P3_U2830));
  AOI22X1 g03369(.A0(n6505), .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B0(P3_REIP_REG_1__SCAN_IN), .B1(n4968), .Y(n6518));
  INVX1   g03370(.A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .Y(n6519));
  AOI22X1 g03371(.A0(n6508), .A1(n6519), .B0(n5088), .B1(n6509), .Y(n6520));
  AOI22X1 g03372(.A0(n6511), .A1(n6519), .B0(n5079), .B1(n6512), .Y(n6521));
  AOI22X1 g03373(.A0(n6514), .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B0(n5079), .B1(n6515), .Y(n6522));
  NAND4X1 g03374(.A(n6521), .B(n6520), .C(n6518), .D(n6522), .Y(P3_U2829));
  AOI22X1 g03375(.A0(n6505), .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B0(n5127), .B1(n6509), .Y(n6524));
  XOR2X1  g03376(.A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .Y(n6525));
  AOI22X1 g03377(.A0(n6508), .A1(n6525), .B0(n4968), .B1(P3_REIP_REG_2__SCAN_IN), .Y(n6526));
  AOI22X1 g03378(.A0(n6512), .A1(n5162), .B0(n6511), .B1(n6525), .Y(n6527));
  INVX1   g03379(.A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .Y(n6528));
  AOI22X1 g03380(.A0(n6514), .A1(n6528), .B0(n5162), .B1(n6515), .Y(n6529));
  NAND4X1 g03381(.A(n6527), .B(n6526), .C(n6524), .D(n6529), .Y(P3_U2828));
  XOR2X1  g03382(.A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .Y(n6531));
  NAND4X1 g03383(.A(n6504), .B(P3_STATEBS16_REG_SCAN_IN), .C(P3_STATE2_REG_1__SCAN_IN), .D(n6531), .Y(n6532));
  NAND2X1 g03384(.A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .Y(n6533));
  XOR2X1  g03385(.A(n6533), .B(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .Y(n6534));
  INVX1   g03386(.A(n6534), .Y(n6535));
  AOI22X1 g03387(.A0(n6512), .A1(n5187), .B0(n6511), .B1(n6535), .Y(n6536));
  NAND2X1 g03388(.A(n6515), .B(n5187), .Y(n6537));
  AOI22X1 g03389(.A0(n6508), .A1(n6535), .B0(n6505), .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .Y(n6539));
  OAI21X1 g03390(.A0(n4969), .A1(n3393), .B0(n6539), .Y(n6540));
  AOI21X1 g03391(.A0(n6509), .A1(n5203), .B0(n6540), .Y(n6541));
  NAND4X1 g03392(.A(n6537), .B(n6536), .C(n6532), .D(n6541), .Y(P3_U2827));
  INVX1   g03393(.A(n6512), .Y(n6543));
  NOR2X1  g03394(.A(n6543), .B(n5256), .Y(n6544));
  NAND3X1 g03395(.A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .C(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .Y(n6545));
  XOR2X1  g03396(.A(n6545), .B(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .Y(n6546));
  INVX1   g03397(.A(n6546), .Y(n6547));
  AOI22X1 g03398(.A0(n6508), .A1(n6547), .B0(n6505), .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .Y(n6548));
  OAI21X1 g03399(.A0(n4969), .A1(n3390), .B0(n6548), .Y(n6549));
  INVX1   g03400(.A(n6511), .Y(n6550));
  INVX1   g03401(.A(n6514), .Y(n6551));
  NAND2X1 g03402(.A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .Y(n6552));
  XOR2X1  g03403(.A(n6552), .B(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .Y(n6553));
  OAI22X1 g03404(.A0(n6546), .A1(n6550), .B0(n6551), .B1(n6553), .Y(n6554));
  NOR3X1  g03405(.A(n6554), .B(n6549), .C(n6544), .Y(n6555));
  INVX1   g03406(.A(n5256), .Y(n6556));
  NOR4X1  g03407(.A(n5266), .B(n3682), .C(n3510), .D(n6505), .Y(n6557));
  AOI21X1 g03408(.A0(n6515), .A1(n6556), .B0(n6557), .Y(n6558));
  NAND2X1 g03409(.A(n6558), .B(n6555), .Y(P3_U2826));
  NOR2X1  g03410(.A(n5335), .B(n5329), .Y(n6560));
  NAND2X1 g03411(.A(n6509), .B(n6560), .Y(n6561));
  NOR2X1  g03412(.A(n6543), .B(n5346), .Y(n6562));
  INVX1   g03413(.A(n6515), .Y(n6563));
  NOR2X1  g03414(.A(n6563), .B(n5346), .Y(n6564));
  NAND4X1 g03415(.A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .C(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .D(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .Y(n6565));
  XOR2X1  g03416(.A(n6565), .B(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .Y(n6566));
  INVX1   g03417(.A(n6566), .Y(n6567));
  AOI22X1 g03418(.A0(n6508), .A1(n6567), .B0(n6505), .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .Y(n6568));
  OAI21X1 g03419(.A0(n4969), .A1(n3387), .B0(n6568), .Y(n6569));
  NAND3X1 g03420(.A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .C(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .Y(n6570));
  XOR2X1  g03421(.A(n6570), .B(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .Y(n6571));
  OAI22X1 g03422(.A0(n6566), .A1(n6550), .B0(n6551), .B1(n6571), .Y(n6572));
  NOR4X1  g03423(.A(n6569), .B(n6564), .C(n6562), .D(n6572), .Y(n6573));
  NAND2X1 g03424(.A(n6573), .B(n6561), .Y(P3_U2825));
  NOR2X1  g03425(.A(n6543), .B(n5416), .Y(n6575));
  NOR4X1  g03426(.A(n5426), .B(n3682), .C(n3510), .D(n6505), .Y(n6576));
  INVX1   g03427(.A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .Y(n6577));
  INVX1   g03428(.A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .Y(n6578));
  NOR2X1  g03429(.A(n6565), .B(n6578), .Y(n6579));
  XOR2X1  g03430(.A(n6579), .B(n6577), .Y(n6580));
  INVX1   g03431(.A(n6580), .Y(n6581));
  AOI22X1 g03432(.A0(n6508), .A1(n6581), .B0(n6505), .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .Y(n6582));
  OAI21X1 g03433(.A0(n4969), .A1(n3384), .B0(n6582), .Y(n6583));
  NAND4X1 g03434(.A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .C(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .D(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .Y(n6584));
  XOR2X1  g03435(.A(n6584), .B(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .Y(n6585));
  OAI22X1 g03436(.A0(n6580), .A1(n6550), .B0(n6551), .B1(n6585), .Y(n6586));
  NOR4X1  g03437(.A(n6583), .B(n6576), .C(n6575), .D(n6586), .Y(n6587));
  OAI21X1 g03438(.A0(n6563), .A1(n5416), .B0(n6587), .Y(P3_U2824));
  NOR2X1  g03439(.A(n6543), .B(n5474), .Y(n6589));
  INVX1   g03440(.A(n6509), .Y(n6590));
  NOR2X1  g03441(.A(n6590), .B(n5483), .Y(n6591));
  INVX1   g03442(.A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .Y(n6592));
  NOR3X1  g03443(.A(n6565), .B(n6577), .C(n6578), .Y(n6593));
  XOR2X1  g03444(.A(n6593), .B(n6592), .Y(n6594));
  INVX1   g03445(.A(n6594), .Y(n6595));
  AOI22X1 g03446(.A0(n6508), .A1(n6595), .B0(n6505), .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .Y(n6596));
  OAI21X1 g03447(.A0(n4969), .A1(n3381), .B0(n6596), .Y(n6597));
  NOR2X1  g03448(.A(n6584), .B(n6577), .Y(n6598));
  XOR2X1  g03449(.A(n6598), .B(n6592), .Y(n6599));
  OAI22X1 g03450(.A0(n6594), .A1(n6550), .B0(n6551), .B1(n6599), .Y(n6600));
  NOR4X1  g03451(.A(n6597), .B(n6591), .C(n6589), .D(n6600), .Y(n6601));
  OAI21X1 g03452(.A0(n6563), .A1(n5474), .B0(n6601), .Y(P3_U2823));
  NOR2X1  g03453(.A(n6590), .B(n5528), .Y(n6603));
  NOR2X1  g03454(.A(n6543), .B(n5535), .Y(n6604));
  INVX1   g03455(.A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .Y(n6605));
  NOR4X1  g03456(.A(n6592), .B(n6577), .C(n6578), .D(n6565), .Y(n6606));
  XOR2X1  g03457(.A(n6606), .B(n6605), .Y(n6607));
  INVX1   g03458(.A(n6607), .Y(n6608));
  AOI22X1 g03459(.A0(n6508), .A1(n6608), .B0(n6505), .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .Y(n6609));
  OAI21X1 g03460(.A0(n4969), .A1(n3378), .B0(n6609), .Y(n6610));
  NOR3X1  g03461(.A(n6584), .B(n6592), .C(n6577), .Y(n6611));
  XOR2X1  g03462(.A(n6611), .B(n6605), .Y(n6612));
  OAI22X1 g03463(.A0(n6607), .A1(n6550), .B0(n6551), .B1(n6612), .Y(n6613));
  NOR4X1  g03464(.A(n6610), .B(n6604), .C(n6603), .D(n6613), .Y(n6614));
  OAI21X1 g03465(.A0(n6563), .A1(n5520), .B0(n6614), .Y(P3_U2822));
  NAND2X1 g03466(.A(n6515), .B(n5569), .Y(n6616));
  NAND2X1 g03467(.A(n6512), .B(n5577), .Y(n6617));
  NAND2X1 g03468(.A(n6509), .B(n5582), .Y(n6618));
  NAND2X1 g03469(.A(n6606), .B(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .Y(n6619));
  XOR2X1  g03470(.A(n6619), .B(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .Y(n6620));
  INVX1   g03471(.A(n6620), .Y(n6621));
  AOI22X1 g03472(.A0(n6508), .A1(n6621), .B0(n6505), .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .Y(n6622));
  OAI21X1 g03473(.A0(n4969), .A1(n3375), .B0(n6622), .Y(n6623));
  INVX1   g03474(.A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .Y(n6624));
  NOR4X1  g03475(.A(n6605), .B(n6592), .C(n6577), .D(n6584), .Y(n6625));
  XOR2X1  g03476(.A(n6625), .B(n6624), .Y(n6626));
  OAI22X1 g03477(.A0(n6620), .A1(n6550), .B0(n6551), .B1(n6626), .Y(n6627));
  NOR2X1  g03478(.A(n6627), .B(n6623), .Y(n6628));
  NAND4X1 g03479(.A(n6618), .B(n6617), .C(n6616), .D(n6628), .Y(P3_U2821));
  NOR2X1  g03480(.A(n6563), .B(n5618), .Y(n6630));
  NOR2X1  g03481(.A(n6590), .B(n5630), .Y(n6631));
  NAND3X1 g03482(.A(n6606), .B(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .C(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .Y(n6632));
  XOR2X1  g03483(.A(n6632), .B(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .Y(n6633));
  INVX1   g03484(.A(n6633), .Y(n6634));
  AOI22X1 g03485(.A0(n6508), .A1(n6634), .B0(n6505), .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .Y(n6635));
  OAI21X1 g03486(.A0(n4969), .A1(n3372), .B0(n6635), .Y(n6636));
  NAND2X1 g03487(.A(n6625), .B(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .Y(n6637));
  XOR2X1  g03488(.A(n6637), .B(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .Y(n6638));
  OAI22X1 g03489(.A0(n6633), .A1(n6550), .B0(n6551), .B1(n6638), .Y(n6639));
  NOR4X1  g03490(.A(n6636), .B(n6631), .C(n6630), .D(n6639), .Y(n6640));
  OAI21X1 g03491(.A0(n6543), .A1(n5625), .B0(n6640), .Y(P3_U2820));
  NAND2X1 g03492(.A(n6512), .B(n5664), .Y(n6642));
  NOR2X1  g03493(.A(n6563), .B(n5666), .Y(n6643));
  NOR2X1  g03494(.A(n6590), .B(n5667), .Y(n6644));
  NAND4X1 g03495(.A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .C(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .D(n6606), .Y(n6645));
  XOR2X1  g03496(.A(n6645), .B(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .Y(n6646));
  INVX1   g03497(.A(n6646), .Y(n6647));
  AOI22X1 g03498(.A0(n6508), .A1(n6647), .B0(n6505), .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .Y(n6648));
  OAI21X1 g03499(.A0(n4969), .A1(n3369), .B0(n6648), .Y(n6649));
  NAND3X1 g03500(.A(n6625), .B(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .C(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .Y(n6650));
  XOR2X1  g03501(.A(n6650), .B(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .Y(n6651));
  OAI22X1 g03502(.A0(n6646), .A1(n6550), .B0(n6551), .B1(n6651), .Y(n6652));
  NOR4X1  g03503(.A(n6649), .B(n6644), .C(n6643), .D(n6652), .Y(n6653));
  NAND2X1 g03504(.A(n6653), .B(n6642), .Y(P3_U2819));
  NOR2X1  g03505(.A(n5700), .B(n5698), .Y(n6655));
  NAND2X1 g03506(.A(n6515), .B(n6655), .Y(n6656));
  NOR2X1  g03507(.A(n6543), .B(n5711), .Y(n6657));
  NOR3X1  g03508(.A(n6590), .B(n5714), .C(n5713), .Y(n6658));
  INVX1   g03509(.A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .Y(n6659));
  INVX1   g03510(.A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .Y(n6660));
  NOR2X1  g03511(.A(n6645), .B(n6660), .Y(n6661));
  XOR2X1  g03512(.A(n6661), .B(n6659), .Y(n6662));
  INVX1   g03513(.A(n6662), .Y(n6663));
  AOI22X1 g03514(.A0(n6508), .A1(n6663), .B0(n6505), .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .Y(n6664));
  OAI21X1 g03515(.A0(n4969), .A1(n3366), .B0(n6664), .Y(n6665));
  NAND4X1 g03516(.A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .C(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .D(n6625), .Y(n6666));
  XOR2X1  g03517(.A(n6666), .B(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .Y(n6667));
  OAI22X1 g03518(.A0(n6662), .A1(n6550), .B0(n6551), .B1(n6667), .Y(n6668));
  NOR4X1  g03519(.A(n6665), .B(n6658), .C(n6657), .D(n6668), .Y(n6669));
  NAND2X1 g03520(.A(n6669), .B(n6656), .Y(P3_U2818));
  NAND2X1 g03521(.A(n6515), .B(n5753), .Y(n6671));
  NAND2X1 g03522(.A(n6512), .B(n5752), .Y(n6672));
  NAND2X1 g03523(.A(n6509), .B(n5755), .Y(n6673));
  INVX1   g03524(.A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .Y(n6674));
  NOR3X1  g03525(.A(n6645), .B(n6659), .C(n6660), .Y(n6675));
  XOR2X1  g03526(.A(n6675), .B(n6674), .Y(n6676));
  INVX1   g03527(.A(n6676), .Y(n6677));
  AOI22X1 g03528(.A0(n6508), .A1(n6677), .B0(n6505), .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .Y(n6678));
  OAI21X1 g03529(.A0(n4969), .A1(n3363), .B0(n6678), .Y(n6679));
  NOR2X1  g03530(.A(n6666), .B(n6659), .Y(n6680));
  XOR2X1  g03531(.A(n6680), .B(n6674), .Y(n6681));
  OAI22X1 g03532(.A0(n6676), .A1(n6550), .B0(n6551), .B1(n6681), .Y(n6682));
  NOR2X1  g03533(.A(n6682), .B(n6679), .Y(n6683));
  NAND4X1 g03534(.A(n6673), .B(n6672), .C(n6671), .D(n6683), .Y(P3_U2817));
  NOR2X1  g03535(.A(n6590), .B(n5787), .Y(n6685));
  NAND2X1 g03536(.A(n6512), .B(n5792), .Y(n6686));
  INVX1   g03537(.A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .Y(n6687));
  INVX1   g03538(.A(n6508), .Y(n6688));
  NOR4X1  g03539(.A(n6674), .B(n6659), .C(n6660), .D(n6645), .Y(n6689));
  XOR2X1  g03540(.A(n6689), .B(n6687), .Y(n6690));
  OAI22X1 g03541(.A0(n6688), .A1(n6690), .B0(n6504), .B1(n6687), .Y(n6691));
  AOI21X1 g03542(.A0(n4968), .A1(P3_REIP_REG_14__SCAN_IN), .B0(n6691), .Y(n6692));
  INVX1   g03543(.A(n6690), .Y(n6693));
  NOR3X1  g03544(.A(n6666), .B(n6674), .C(n6659), .Y(n6694));
  XOR2X1  g03545(.A(n6694), .B(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .Y(n6695));
  AOI22X1 g03546(.A0(n6693), .A1(n6511), .B0(n6514), .B1(n6695), .Y(n6696));
  NAND3X1 g03547(.A(n6696), .B(n6692), .C(n6686), .Y(n6697));
  NOR2X1  g03548(.A(n6697), .B(n6685), .Y(n6698));
  OAI21X1 g03549(.A0(n6563), .A1(n5784), .B0(n6698), .Y(P3_U2816));
  INVX1   g03550(.A(n5820), .Y(n6700));
  NAND3X1 g03551(.A(n6515), .B(n5821), .C(n6700), .Y(n6701));
  NOR2X1  g03552(.A(n6543), .B(n5828), .Y(n6702));
  NOR3X1  g03553(.A(n6590), .B(n5832), .C(n5830), .Y(n6703));
  NAND2X1 g03554(.A(n6689), .B(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .Y(n6704));
  XOR2X1  g03555(.A(n6704), .B(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .Y(n6705));
  INVX1   g03556(.A(n6705), .Y(n6706));
  AOI22X1 g03557(.A0(n6508), .A1(n6706), .B0(n6505), .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .Y(n6707));
  OAI21X1 g03558(.A0(n4969), .A1(n3357), .B0(n6707), .Y(n6708));
  INVX1   g03559(.A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .Y(n6709));
  NOR4X1  g03560(.A(n6687), .B(n6674), .C(n6659), .D(n6666), .Y(n6710));
  XOR2X1  g03561(.A(n6710), .B(n6709), .Y(n6711));
  OAI22X1 g03562(.A0(n6705), .A1(n6550), .B0(n6551), .B1(n6711), .Y(n6712));
  NOR4X1  g03563(.A(n6708), .B(n6703), .C(n6702), .D(n6712), .Y(n6713));
  NAND2X1 g03564(.A(n6713), .B(n6701), .Y(P3_U2815));
  NOR2X1  g03565(.A(n6563), .B(n5866), .Y(n6715));
  NOR2X1  g03566(.A(n6590), .B(n5868), .Y(n6716));
  NAND3X1 g03567(.A(n6689), .B(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .Y(n6717));
  XOR2X1  g03568(.A(n6717), .B(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .Y(n6718));
  INVX1   g03569(.A(n6718), .Y(n6719));
  AOI22X1 g03570(.A0(n6508), .A1(n6719), .B0(n6505), .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .Y(n6720));
  OAI21X1 g03571(.A0(n4969), .A1(n3354), .B0(n6720), .Y(n6721));
  NAND2X1 g03572(.A(n6710), .B(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .Y(n6722));
  XOR2X1  g03573(.A(n6722), .B(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .Y(n6723));
  OAI22X1 g03574(.A0(n6718), .A1(n6550), .B0(n6551), .B1(n6723), .Y(n6724));
  NOR4X1  g03575(.A(n6721), .B(n6716), .C(n6715), .D(n6724), .Y(n6725));
  OAI21X1 g03576(.A0(n6543), .A1(n5864), .B0(n6725), .Y(P3_U2814));
  NAND2X1 g03577(.A(n6512), .B(n5904), .Y(n6727));
  NOR3X1  g03578(.A(n6563), .B(n5907), .C(n5905), .Y(n6728));
  NOR3X1  g03579(.A(n6590), .B(n5911), .C(n5910), .Y(n6729));
  INVX1   g03580(.A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .Y(n6730));
  NAND4X1 g03581(.A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .D(n6689), .Y(n6731));
  XOR2X1  g03582(.A(n6731), .B(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .Y(n6732));
  OAI22X1 g03583(.A0(n6688), .A1(n6732), .B0(n6504), .B1(n6730), .Y(n6733));
  AOI21X1 g03584(.A0(n4968), .A1(P3_REIP_REG_17__SCAN_IN), .B0(n6733), .Y(n6734));
  INVX1   g03585(.A(n6732), .Y(n6735));
  NAND3X1 g03586(.A(n6710), .B(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .C(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .Y(n6736));
  XOR2X1  g03587(.A(n6736), .B(n6730), .Y(n6737));
  AOI22X1 g03588(.A0(n6735), .A1(n6511), .B0(n6514), .B1(n6737), .Y(n6738));
  NAND2X1 g03589(.A(n6738), .B(n6734), .Y(n6739));
  NOR3X1  g03590(.A(n6739), .B(n6729), .C(n6728), .Y(n6740));
  NAND2X1 g03591(.A(n6740), .B(n6727), .Y(P3_U2813));
  NOR2X1  g03592(.A(n6563), .B(n5947), .Y(n6742));
  NOR2X1  g03593(.A(n6590), .B(n5949), .Y(n6743));
  INVX1   g03594(.A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .Y(n6744));
  NOR2X1  g03595(.A(n6731), .B(n6730), .Y(n6745));
  XOR2X1  g03596(.A(n6745), .B(n6744), .Y(n6746));
  OAI22X1 g03597(.A0(n6688), .A1(n6746), .B0(n6504), .B1(n6744), .Y(n6747));
  AOI21X1 g03598(.A0(n4968), .A1(P3_REIP_REG_18__SCAN_IN), .B0(n6747), .Y(n6748));
  INVX1   g03599(.A(n6746), .Y(n6749));
  NAND4X1 g03600(.A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .C(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .D(n6710), .Y(n6750));
  XOR2X1  g03601(.A(n6750), .B(n6744), .Y(n6751));
  AOI22X1 g03602(.A0(n6749), .A1(n6511), .B0(n6514), .B1(n6751), .Y(n6752));
  NAND2X1 g03603(.A(n6752), .B(n6748), .Y(n6753));
  NOR3X1  g03604(.A(n6753), .B(n6743), .C(n6742), .Y(n6754));
  OAI21X1 g03605(.A0(n6543), .A1(n5945), .B0(n6754), .Y(P3_U2812));
  NOR3X1  g03606(.A(n6563), .B(n5987), .C(n5986), .Y(n6756));
  NOR2X1  g03607(.A(n6590), .B(n5992), .Y(n6757));
  INVX1   g03608(.A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .Y(n6758));
  NOR3X1  g03609(.A(n6731), .B(n6744), .C(n6730), .Y(n6759));
  XOR2X1  g03610(.A(n6759), .B(n6758), .Y(n6760));
  AOI22X1 g03611(.A0(n6505), .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B0(P3_REIP_REG_19__SCAN_IN), .B1(n4968), .Y(n6761));
  OAI21X1 g03612(.A0(n6760), .A1(n6688), .B0(n6761), .Y(n6762));
  NOR2X1  g03613(.A(n6750), .B(n6744), .Y(n6763));
  XOR2X1  g03614(.A(n6763), .B(n6758), .Y(n6764));
  OAI22X1 g03615(.A0(n6760), .A1(n6550), .B0(n6551), .B1(n6764), .Y(n6765));
  NOR4X1  g03616(.A(n6762), .B(n6757), .C(n6756), .D(n6765), .Y(n6766));
  OAI21X1 g03617(.A0(n6543), .A1(n5984), .B0(n6766), .Y(P3_U2811));
  NAND2X1 g03618(.A(n6509), .B(n6031), .Y(n6768));
  INVX1   g03619(.A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .Y(n6769));
  NOR4X1  g03620(.A(n6758), .B(n6744), .C(n6730), .D(n6731), .Y(n6770));
  XOR2X1  g03621(.A(n6770), .B(n6769), .Y(n6771));
  NOR4X1  g03622(.A(n6505), .B(P3_STATEBS16_REG_SCAN_IN), .C(n3939), .D(n6771), .Y(n6772));
  NOR2X1  g03623(.A(n6771), .B(n6688), .Y(n6773));
  NOR3X1  g03624(.A(n6750), .B(n6758), .C(n6744), .Y(n6774));
  XOR2X1  g03625(.A(n6774), .B(n6769), .Y(n6775));
  NOR4X1  g03626(.A(n6505), .B(n3944), .C(n3939), .D(n6775), .Y(n6776));
  OAI22X1 g03627(.A0(n6504), .A1(n6769), .B0(n3342), .B1(n4969), .Y(n6777));
  NOR4X1  g03628(.A(n6776), .B(n6773), .C(n6772), .D(n6777), .Y(n6778));
  NAND2X1 g03629(.A(n6778), .B(n6768), .Y(n6779));
  AOI21X1 g03630(.A0(n6515), .A1(n6030), .B0(n6779), .Y(n6780));
  OAI21X1 g03631(.A0(n6543), .A1(n6029), .B0(n6780), .Y(P3_U2810));
  NAND3X1 g03632(.A(n6509), .B(n6071), .C(n6069), .Y(n6782));
  NAND2X1 g03633(.A(n6770), .B(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .Y(n6783));
  XOR2X1  g03634(.A(n6783), .B(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .Y(n6784));
  NOR4X1  g03635(.A(n6505), .B(P3_STATEBS16_REG_SCAN_IN), .C(n3939), .D(n6784), .Y(n6785));
  NOR2X1  g03636(.A(n6784), .B(n6688), .Y(n6786));
  INVX1   g03637(.A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .Y(n6787));
  NOR4X1  g03638(.A(n6769), .B(n6758), .C(n6744), .D(n6750), .Y(n6788));
  XOR2X1  g03639(.A(n6788), .B(n6787), .Y(n6789));
  NOR4X1  g03640(.A(n6505), .B(n3944), .C(n3939), .D(n6789), .Y(n6790));
  OAI22X1 g03641(.A0(n6504), .A1(n6787), .B0(n3339), .B1(n4969), .Y(n6791));
  NOR4X1  g03642(.A(n6790), .B(n6786), .C(n6785), .D(n6791), .Y(n6792));
  NAND2X1 g03643(.A(n6792), .B(n6782), .Y(n6793));
  AOI21X1 g03644(.A0(n6515), .A1(n6067), .B0(n6793), .Y(n6794));
  OAI21X1 g03645(.A0(n6543), .A1(n6063), .B0(n6794), .Y(P3_U2809));
  NAND2X1 g03646(.A(n6512), .B(n6106), .Y(n6796));
  NOR2X1  g03647(.A(n6563), .B(n6109), .Y(n6797));
  NAND3X1 g03648(.A(n6770), .B(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .Y(n6798));
  XOR2X1  g03649(.A(n6798), .B(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .Y(n6799));
  NOR4X1  g03650(.A(n6505), .B(P3_STATEBS16_REG_SCAN_IN), .C(n3939), .D(n6799), .Y(n6800));
  NOR2X1  g03651(.A(n6799), .B(n6688), .Y(n6801));
  NAND2X1 g03652(.A(n6788), .B(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .Y(n6802));
  XOR2X1  g03653(.A(n6802), .B(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .Y(n6803));
  AOI22X1 g03654(.A0(n6505), .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B0(P3_REIP_REG_22__SCAN_IN), .B1(n4968), .Y(n6804));
  OAI21X1 g03655(.A0(n6803), .A1(n6551), .B0(n6804), .Y(n6805));
  NOR3X1  g03656(.A(n6805), .B(n6801), .C(n6800), .Y(n6806));
  OAI21X1 g03657(.A0(n6590), .A1(n6110), .B0(n6806), .Y(n6807));
  NOR2X1  g03658(.A(n6807), .B(n6797), .Y(n6808));
  NAND2X1 g03659(.A(n6808), .B(n6796), .Y(P3_U2808));
  NAND2X1 g03660(.A(n6512), .B(n6143), .Y(n6810));
  INVX1   g03661(.A(n6150), .Y(n6811));
  NAND2X1 g03662(.A(n6515), .B(n6811), .Y(n6812));
  NAND3X1 g03663(.A(n6509), .B(n6154), .C(n6152), .Y(n6813));
  NAND4X1 g03664(.A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .D(n6770), .Y(n6814));
  XOR2X1  g03665(.A(n6814), .B(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .Y(n6815));
  NOR4X1  g03666(.A(n6505), .B(P3_STATEBS16_REG_SCAN_IN), .C(n3939), .D(n6815), .Y(n6816));
  NOR2X1  g03667(.A(n6815), .B(n6688), .Y(n6817));
  NAND3X1 g03668(.A(n6788), .B(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .C(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .Y(n6818));
  XOR2X1  g03669(.A(n6818), .B(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .Y(n6819));
  NOR4X1  g03670(.A(n6505), .B(n3944), .C(n3939), .D(n6819), .Y(n6820));
  INVX1   g03671(.A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .Y(n6821));
  OAI22X1 g03672(.A0(n6504), .A1(n6821), .B0(n3333), .B1(n4969), .Y(n6822));
  NOR4X1  g03673(.A(n6820), .B(n6817), .C(n6816), .D(n6822), .Y(n6823));
  NAND4X1 g03674(.A(n6813), .B(n6812), .C(n6810), .D(n6823), .Y(P3_U2807));
  NAND2X1 g03675(.A(n6512), .B(n6186), .Y(n6825));
  INVX1   g03676(.A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .Y(n6826));
  NOR2X1  g03677(.A(n6814), .B(n6821), .Y(n6827));
  XOR2X1  g03678(.A(n6827), .B(n6826), .Y(n6828));
  NOR4X1  g03679(.A(n6505), .B(P3_STATEBS16_REG_SCAN_IN), .C(n3939), .D(n6828), .Y(n6829));
  NOR2X1  g03680(.A(n6828), .B(n6688), .Y(n6830));
  NAND4X1 g03681(.A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .C(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .D(n6788), .Y(n6831));
  XOR2X1  g03682(.A(n6831), .B(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .Y(n6832));
  NOR4X1  g03683(.A(n6505), .B(n3944), .C(n3939), .D(n6832), .Y(n6833));
  OAI22X1 g03684(.A0(n6504), .A1(n6826), .B0(n3330), .B1(n4969), .Y(n6834));
  NOR4X1  g03685(.A(n6833), .B(n6830), .C(n6829), .D(n6834), .Y(n6835));
  OAI21X1 g03686(.A0(n6590), .A1(n6190), .B0(n6835), .Y(n6836));
  AOI21X1 g03687(.A0(n6515), .A1(n6187), .B0(n6836), .Y(n6837));
  NAND2X1 g03688(.A(n6837), .B(n6825), .Y(P3_U2806));
  NAND2X1 g03689(.A(n6512), .B(n6227), .Y(n6839));
  NAND2X1 g03690(.A(n6515), .B(n6230), .Y(n6840));
  INVX1   g03691(.A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .Y(n6841));
  NOR3X1  g03692(.A(n6814), .B(n6826), .C(n6821), .Y(n6842));
  XOR2X1  g03693(.A(n6842), .B(n6841), .Y(n6843));
  INVX1   g03694(.A(n6843), .Y(n6844));
  NOR2X1  g03695(.A(n6831), .B(n6826), .Y(n6845));
  XOR2X1  g03696(.A(n6845), .B(n6841), .Y(n6846));
  AOI22X1 g03697(.A0(n6505), .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B0(P3_REIP_REG_25__SCAN_IN), .B1(n4968), .Y(n6847));
  OAI21X1 g03698(.A0(n6846), .A1(n6551), .B0(n6847), .Y(n6848));
  AOI21X1 g03699(.A0(n6844), .A1(n6508), .B0(n6848), .Y(n6849));
  OAI21X1 g03700(.A0(n6843), .A1(n6550), .B0(n6849), .Y(n6850));
  AOI21X1 g03701(.A0(n6509), .A1(n6234), .B0(n6850), .Y(n6851));
  NAND3X1 g03702(.A(n6851), .B(n6840), .C(n6839), .Y(P3_U2805));
  NAND2X1 g03703(.A(n6509), .B(n6272), .Y(n6853));
  INVX1   g03704(.A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .Y(n6854));
  NOR4X1  g03705(.A(n6841), .B(n6826), .C(n6821), .D(n6814), .Y(n6855));
  XOR2X1  g03706(.A(n6855), .B(n6854), .Y(n6856));
  NOR2X1  g03707(.A(n6856), .B(n6688), .Y(n6857));
  NOR4X1  g03708(.A(n6505), .B(P3_STATEBS16_REG_SCAN_IN), .C(n3939), .D(n6856), .Y(n6858));
  NOR3X1  g03709(.A(n6831), .B(n6841), .C(n6826), .Y(n6859));
  XOR2X1  g03710(.A(n6859), .B(n6854), .Y(n6860));
  NOR4X1  g03711(.A(n6505), .B(n3944), .C(n3939), .D(n6860), .Y(n6861));
  OAI22X1 g03712(.A0(n6504), .A1(n6854), .B0(n3324), .B1(n4969), .Y(n6862));
  NOR4X1  g03713(.A(n6861), .B(n6858), .C(n6857), .D(n6862), .Y(n6863));
  NAND2X1 g03714(.A(n6863), .B(n6853), .Y(n6864));
  AOI21X1 g03715(.A0(n6515), .A1(n6270), .B0(n6864), .Y(n6865));
  OAI21X1 g03716(.A0(n6543), .A1(n6268), .B0(n6865), .Y(P3_U2804));
  NOR2X1  g03717(.A(n6563), .B(n6305), .Y(n6867));
  NAND2X1 g03718(.A(n6855), .B(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .Y(n6868));
  XOR2X1  g03719(.A(n6868), .B(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .Y(n6869));
  NOR2X1  g03720(.A(n6869), .B(n6688), .Y(n6870));
  NOR4X1  g03721(.A(n6505), .B(P3_STATEBS16_REG_SCAN_IN), .C(n3939), .D(n6869), .Y(n6871));
  INVX1   g03722(.A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .Y(n6872));
  NOR4X1  g03723(.A(n6854), .B(n6841), .C(n6826), .D(n6831), .Y(n6873));
  XOR2X1  g03724(.A(n6873), .B(n6872), .Y(n6874));
  NOR4X1  g03725(.A(n6505), .B(n3944), .C(n3939), .D(n6874), .Y(n6875));
  OAI22X1 g03726(.A0(n6504), .A1(n6872), .B0(n3321), .B1(n4969), .Y(n6876));
  NOR4X1  g03727(.A(n6875), .B(n6871), .C(n6870), .D(n6876), .Y(n6877));
  OAI21X1 g03728(.A0(n6590), .A1(n6308), .B0(n6877), .Y(n6878));
  NOR2X1  g03729(.A(n6878), .B(n6867), .Y(n6879));
  OAI21X1 g03730(.A0(n6543), .A1(n6302), .B0(n6879), .Y(P3_U2803));
  NAND2X1 g03731(.A(n6512), .B(n6345), .Y(n6881));
  NOR2X1  g03732(.A(n6563), .B(n6348), .Y(n6882));
  NOR3X1  g03733(.A(n6590), .B(n6351), .C(n6349), .Y(n6883));
  NAND3X1 g03734(.A(n6855), .B(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .Y(n6884));
  XOR2X1  g03735(.A(n6884), .B(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .Y(n6885));
  NOR2X1  g03736(.A(n6885), .B(n6688), .Y(n6886));
  NAND2X1 g03737(.A(n6873), .B(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .Y(n6887));
  XOR2X1  g03738(.A(n6887), .B(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .Y(n6888));
  AOI22X1 g03739(.A0(n6505), .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B0(P3_REIP_REG_28__SCAN_IN), .B1(n4968), .Y(n6889));
  OAI21X1 g03740(.A0(n6888), .A1(n6551), .B0(n6889), .Y(n6890));
  NOR2X1  g03741(.A(n6890), .B(n6886), .Y(n6891));
  OAI21X1 g03742(.A0(n6885), .A1(n6550), .B0(n6891), .Y(n6892));
  NOR3X1  g03743(.A(n6892), .B(n6883), .C(n6882), .Y(n6893));
  NAND2X1 g03744(.A(n6893), .B(n6881), .Y(P3_U2802));
  NAND2X1 g03745(.A(n6509), .B(n6389), .Y(n6895));
  NAND4X1 g03746(.A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .D(n6855), .Y(n6896));
  XOR2X1  g03747(.A(n6896), .B(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .Y(n6897));
  NOR4X1  g03748(.A(n6505), .B(P3_STATEBS16_REG_SCAN_IN), .C(n3939), .D(n6897), .Y(n6898));
  NOR2X1  g03749(.A(n6897), .B(n6688), .Y(n6899));
  NAND3X1 g03750(.A(n6873), .B(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .Y(n6900));
  XOR2X1  g03751(.A(n6900), .B(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .Y(n6901));
  NOR4X1  g03752(.A(n6505), .B(n3944), .C(n3939), .D(n6901), .Y(n6902));
  INVX1   g03753(.A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .Y(n6903));
  OAI22X1 g03754(.A0(n6504), .A1(n6903), .B0(n3315), .B1(n4969), .Y(n6904));
  NOR4X1  g03755(.A(n6902), .B(n6899), .C(n6898), .D(n6904), .Y(n6905));
  NAND2X1 g03756(.A(n6905), .B(n6895), .Y(n6906));
  AOI21X1 g03757(.A0(n6515), .A1(n6387), .B0(n6906), .Y(n6907));
  OAI21X1 g03758(.A0(n6543), .A1(n6384), .B0(n6907), .Y(P3_U2801));
  NOR2X1  g03759(.A(n6563), .B(n6424), .Y(n6909));
  NOR2X1  g03760(.A(n6590), .B(n6428), .Y(n6910));
  INVX1   g03761(.A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .Y(n6911));
  NOR2X1  g03762(.A(n6896), .B(n6903), .Y(n6912));
  XOR2X1  g03763(.A(n6912), .B(n6911), .Y(n6913));
  NOR4X1  g03764(.A(n6505), .B(P3_STATEBS16_REG_SCAN_IN), .C(n3939), .D(n6913), .Y(n6914));
  NAND4X1 g03765(.A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .D(n6873), .Y(n6915));
  XOR2X1  g03766(.A(n6915), .B(n6911), .Y(n6916));
  OAI22X1 g03767(.A0(n6504), .A1(n6911), .B0(n3310), .B1(n4969), .Y(n6917));
  AOI21X1 g03768(.A0(n6916), .A1(n6514), .B0(n6917), .Y(n6918));
  OAI21X1 g03769(.A0(n6913), .A1(n6688), .B0(n6918), .Y(n6919));
  NOR4X1  g03770(.A(n6914), .B(n6910), .C(n6909), .D(n6919), .Y(n6920));
  OAI21X1 g03771(.A0(n6543), .A1(n6421), .B0(n6920), .Y(P3_U2800));
  NAND2X1 g03772(.A(n6512), .B(n6463), .Y(n6922));
  INVX1   g03773(.A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .Y(n6923));
  NOR3X1  g03774(.A(n6896), .B(n6911), .C(n6903), .Y(n6924));
  XOR2X1  g03775(.A(n6924), .B(n6923), .Y(n6925));
  NOR4X1  g03776(.A(n6505), .B(P3_STATEBS16_REG_SCAN_IN), .C(n3939), .D(n6925), .Y(n6926));
  NOR2X1  g03777(.A(n6925), .B(n6688), .Y(n6927));
  NOR2X1  g03778(.A(n6915), .B(n6911), .Y(n6928));
  XOR2X1  g03779(.A(n6928), .B(n6923), .Y(n6929));
  NOR4X1  g03780(.A(n6505), .B(n3944), .C(n3939), .D(n6929), .Y(n6930));
  OAI22X1 g03781(.A0(n6504), .A1(n6923), .B0(n6477), .B1(n4969), .Y(n6931));
  NOR4X1  g03782(.A(n6930), .B(n6927), .C(n6926), .D(n6931), .Y(n6932));
  OAI21X1 g03783(.A0(n6590), .A1(n6470), .B0(n6932), .Y(n6933));
  AOI21X1 g03784(.A0(n6515), .A1(n6468), .B0(n6933), .Y(n6934));
  NAND2X1 g03785(.A(n6934), .B(n6922), .Y(P3_U2799));
  NOR3X1  g03786(.A(n3918), .B(n3704), .C(n3529), .Y(n6936));
  NOR4X1  g03787(.A(n3704), .B(n3529), .C(n3407), .D(n3920), .Y(n6937));
  OAI21X1 g03788(.A0(n6937), .A1(n6936), .B0(n3955), .Y(n6938));
  INVX1   g03789(.A(n6938), .Y(n6939));
  NAND2X1 g03790(.A(n6939), .B(n3682), .Y(n6940));
  NOR2X1  g03791(.A(n6938), .B(n3682), .Y(n6941));
  AOI22X1 g03792(.A0(n6938), .A1(P3_LWORD_REG_15__SCAN_IN), .B0(P3_EAX_REG_15__SCAN_IN), .B1(n6941), .Y(n6942));
  OAI21X1 g03793(.A0(n6940), .A1(n3236), .B0(n6942), .Y(P3_U2798));
  AOI22X1 g03794(.A0(n6938), .A1(P3_LWORD_REG_14__SCAN_IN), .B0(P3_EAX_REG_14__SCAN_IN), .B1(n6941), .Y(n6944));
  OAI21X1 g03795(.A0(n6940), .A1(n3233), .B0(n6944), .Y(P3_U2797));
  AOI22X1 g03796(.A0(n6938), .A1(P3_LWORD_REG_13__SCAN_IN), .B0(P3_EAX_REG_13__SCAN_IN), .B1(n6941), .Y(n6946));
  OAI21X1 g03797(.A0(n6940), .A1(n3230), .B0(n6946), .Y(P3_U2796));
  AOI22X1 g03798(.A0(n6938), .A1(P3_LWORD_REG_12__SCAN_IN), .B0(P3_EAX_REG_12__SCAN_IN), .B1(n6941), .Y(n6948));
  OAI21X1 g03799(.A0(n6940), .A1(n3227), .B0(n6948), .Y(P3_U2795));
  AOI22X1 g03800(.A0(n6938), .A1(P3_LWORD_REG_11__SCAN_IN), .B0(P3_EAX_REG_11__SCAN_IN), .B1(n6941), .Y(n6950));
  OAI21X1 g03801(.A0(n6940), .A1(n3224), .B0(n6950), .Y(P3_U2794));
  AOI22X1 g03802(.A0(n6938), .A1(P3_LWORD_REG_10__SCAN_IN), .B0(P3_EAX_REG_10__SCAN_IN), .B1(n6941), .Y(n6952));
  OAI21X1 g03803(.A0(n6940), .A1(n3221), .B0(n6952), .Y(P3_U2793));
  AOI22X1 g03804(.A0(n6938), .A1(P3_LWORD_REG_9__SCAN_IN), .B0(P3_EAX_REG_9__SCAN_IN), .B1(n6941), .Y(n6954));
  OAI21X1 g03805(.A0(n6940), .A1(n3218), .B0(n6954), .Y(P3_U2792));
  AOI22X1 g03806(.A0(n6938), .A1(P3_LWORD_REG_8__SCAN_IN), .B0(P3_EAX_REG_8__SCAN_IN), .B1(n6941), .Y(n6956));
  OAI21X1 g03807(.A0(n6940), .A1(n3215), .B0(n6956), .Y(P3_U2791));
  AOI22X1 g03808(.A0(n6938), .A1(P3_LWORD_REG_7__SCAN_IN), .B0(P3_EAX_REG_7__SCAN_IN), .B1(n6941), .Y(n6958));
  OAI21X1 g03809(.A0(n6940), .A1(n3212), .B0(n6958), .Y(P3_U2790));
  AOI22X1 g03810(.A0(n6938), .A1(P3_LWORD_REG_6__SCAN_IN), .B0(P3_EAX_REG_6__SCAN_IN), .B1(n6941), .Y(n6960));
  OAI21X1 g03811(.A0(n6940), .A1(n3209), .B0(n6960), .Y(P3_U2789));
  AOI22X1 g03812(.A0(n6938), .A1(P3_LWORD_REG_5__SCAN_IN), .B0(P3_EAX_REG_5__SCAN_IN), .B1(n6941), .Y(n6962));
  OAI21X1 g03813(.A0(n6940), .A1(n3206), .B0(n6962), .Y(P3_U2788));
  AOI22X1 g03814(.A0(n6938), .A1(P3_LWORD_REG_4__SCAN_IN), .B0(P3_EAX_REG_4__SCAN_IN), .B1(n6941), .Y(n6964));
  OAI21X1 g03815(.A0(n6940), .A1(n3203), .B0(n6964), .Y(P3_U2787));
  AOI22X1 g03816(.A0(n6938), .A1(P3_LWORD_REG_3__SCAN_IN), .B0(P3_EAX_REG_3__SCAN_IN), .B1(n6941), .Y(n6966));
  OAI21X1 g03817(.A0(n6940), .A1(n3200), .B0(n6966), .Y(P3_U2786));
  AOI22X1 g03818(.A0(n6938), .A1(P3_LWORD_REG_2__SCAN_IN), .B0(P3_EAX_REG_2__SCAN_IN), .B1(n6941), .Y(n6968));
  OAI21X1 g03819(.A0(n6940), .A1(n3197), .B0(n6968), .Y(P3_U2785));
  AOI22X1 g03820(.A0(n6938), .A1(P3_LWORD_REG_1__SCAN_IN), .B0(P3_EAX_REG_1__SCAN_IN), .B1(n6941), .Y(n6970));
  OAI21X1 g03821(.A0(n6940), .A1(n3194), .B0(n6970), .Y(P3_U2784));
  AOI22X1 g03822(.A0(n6938), .A1(P3_LWORD_REG_0__SCAN_IN), .B0(P3_EAX_REG_0__SCAN_IN), .B1(n6941), .Y(n6972));
  OAI21X1 g03823(.A0(n6940), .A1(n3190), .B0(n6972), .Y(P3_U2783));
  AOI22X1 g03824(.A0(n6938), .A1(P3_UWORD_REG_14__SCAN_IN), .B0(P3_EAX_REG_30__SCAN_IN), .B1(n6941), .Y(n6974));
  OAI21X1 g03825(.A0(n6940), .A1(n3233), .B0(n6974), .Y(P3_U2782));
  AOI22X1 g03826(.A0(n6938), .A1(P3_UWORD_REG_13__SCAN_IN), .B0(P3_EAX_REG_29__SCAN_IN), .B1(n6941), .Y(n6976));
  OAI21X1 g03827(.A0(n6940), .A1(n3230), .B0(n6976), .Y(P3_U2781));
  AOI22X1 g03828(.A0(n6938), .A1(P3_UWORD_REG_12__SCAN_IN), .B0(P3_EAX_REG_28__SCAN_IN), .B1(n6941), .Y(n6978));
  OAI21X1 g03829(.A0(n6940), .A1(n3227), .B0(n6978), .Y(P3_U2780));
  AOI22X1 g03830(.A0(n6938), .A1(P3_UWORD_REG_11__SCAN_IN), .B0(P3_EAX_REG_27__SCAN_IN), .B1(n6941), .Y(n6980));
  OAI21X1 g03831(.A0(n6940), .A1(n3224), .B0(n6980), .Y(P3_U2779));
  AOI22X1 g03832(.A0(n6938), .A1(P3_UWORD_REG_10__SCAN_IN), .B0(P3_EAX_REG_26__SCAN_IN), .B1(n6941), .Y(n6982));
  OAI21X1 g03833(.A0(n6940), .A1(n3221), .B0(n6982), .Y(P3_U2778));
  AOI22X1 g03834(.A0(n6938), .A1(P3_UWORD_REG_9__SCAN_IN), .B0(P3_EAX_REG_25__SCAN_IN), .B1(n6941), .Y(n6984));
  OAI21X1 g03835(.A0(n6940), .A1(n3218), .B0(n6984), .Y(P3_U2777));
  AOI22X1 g03836(.A0(n6938), .A1(P3_UWORD_REG_8__SCAN_IN), .B0(P3_EAX_REG_24__SCAN_IN), .B1(n6941), .Y(n6986));
  OAI21X1 g03837(.A0(n6940), .A1(n3215), .B0(n6986), .Y(P3_U2776));
  AOI22X1 g03838(.A0(n6938), .A1(P3_UWORD_REG_7__SCAN_IN), .B0(P3_EAX_REG_23__SCAN_IN), .B1(n6941), .Y(n6988));
  OAI21X1 g03839(.A0(n6940), .A1(n3212), .B0(n6988), .Y(P3_U2775));
  AOI22X1 g03840(.A0(n6938), .A1(P3_UWORD_REG_6__SCAN_IN), .B0(P3_EAX_REG_22__SCAN_IN), .B1(n6941), .Y(n6990));
  OAI21X1 g03841(.A0(n6940), .A1(n3209), .B0(n6990), .Y(P3_U2774));
  AOI22X1 g03842(.A0(n6938), .A1(P3_UWORD_REG_5__SCAN_IN), .B0(P3_EAX_REG_21__SCAN_IN), .B1(n6941), .Y(n6992));
  OAI21X1 g03843(.A0(n6940), .A1(n3206), .B0(n6992), .Y(P3_U2773));
  AOI22X1 g03844(.A0(n6938), .A1(P3_UWORD_REG_4__SCAN_IN), .B0(P3_EAX_REG_20__SCAN_IN), .B1(n6941), .Y(n6994));
  OAI21X1 g03845(.A0(n6940), .A1(n3203), .B0(n6994), .Y(P3_U2772));
  AOI22X1 g03846(.A0(n6938), .A1(P3_UWORD_REG_3__SCAN_IN), .B0(P3_EAX_REG_19__SCAN_IN), .B1(n6941), .Y(n6996));
  OAI21X1 g03847(.A0(n6940), .A1(n3200), .B0(n6996), .Y(P3_U2771));
  AOI22X1 g03848(.A0(n6938), .A1(P3_UWORD_REG_2__SCAN_IN), .B0(P3_EAX_REG_18__SCAN_IN), .B1(n6941), .Y(n6998));
  OAI21X1 g03849(.A0(n6940), .A1(n3197), .B0(n6998), .Y(P3_U2770));
  AOI22X1 g03850(.A0(n6938), .A1(P3_UWORD_REG_1__SCAN_IN), .B0(P3_EAX_REG_17__SCAN_IN), .B1(n6941), .Y(n7000));
  OAI21X1 g03851(.A0(n6940), .A1(n3194), .B0(n7000), .Y(P3_U2769));
  AOI22X1 g03852(.A0(n6938), .A1(P3_UWORD_REG_0__SCAN_IN), .B0(P3_EAX_REG_16__SCAN_IN), .B1(n6941), .Y(n7002));
  OAI21X1 g03853(.A0(n6940), .A1(n3190), .B0(n7002), .Y(P3_U2768));
  INVX1   g03854(.A(P3_EAX_REG_0__SCAN_IN), .Y(n7004));
  NAND2X1 g03855(.A(n3955), .B(n3725), .Y(n7005));
  OAI22X1 g03856(.A0(n3733), .A1(n7005), .B0(n3958), .B1(P3_STATE2_REG_0__SCAN_IN), .Y(n7006));
  INVX1   g03857(.A(n7006), .Y(n7007));
  NOR2X1  g03858(.A(n7007), .B(n3510), .Y(n7008));
  INVX1   g03859(.A(n7008), .Y(n7009));
  NOR3X1  g03860(.A(P3_STATE2_REG_0__SCAN_IN), .B(n3939), .C(n3511), .Y(n7010));
  AOI22X1 g03861(.A0(n7007), .A1(P3_DATAO_REG_0__SCAN_IN), .B0(P3_LWORD_REG_0__SCAN_IN), .B1(n7010), .Y(n7011));
  OAI21X1 g03862(.A0(n7009), .A1(n7004), .B0(n7011), .Y(P3_U2767));
  NAND3X1 g03863(.A(n7006), .B(P3_EAX_REG_1__SCAN_IN), .C(P3_STATE2_REG_0__SCAN_IN), .Y(n7013));
  AOI22X1 g03864(.A0(n7007), .A1(P3_DATAO_REG_1__SCAN_IN), .B0(P3_LWORD_REG_1__SCAN_IN), .B1(n7010), .Y(n7014));
  NAND2X1 g03865(.A(n7014), .B(n7013), .Y(P3_U2766));
  INVX1   g03866(.A(P3_EAX_REG_2__SCAN_IN), .Y(n7016));
  AOI22X1 g03867(.A0(n7007), .A1(P3_DATAO_REG_2__SCAN_IN), .B0(P3_LWORD_REG_2__SCAN_IN), .B1(n7010), .Y(n7017));
  OAI21X1 g03868(.A0(n7009), .A1(n7016), .B0(n7017), .Y(P3_U2765));
  INVX1   g03869(.A(P3_EAX_REG_3__SCAN_IN), .Y(n7019));
  AOI22X1 g03870(.A0(n7007), .A1(P3_DATAO_REG_3__SCAN_IN), .B0(P3_LWORD_REG_3__SCAN_IN), .B1(n7010), .Y(n7020));
  OAI21X1 g03871(.A0(n7009), .A1(n7019), .B0(n7020), .Y(P3_U2764));
  INVX1   g03872(.A(P3_EAX_REG_4__SCAN_IN), .Y(n7022));
  AOI22X1 g03873(.A0(n7007), .A1(P3_DATAO_REG_4__SCAN_IN), .B0(P3_LWORD_REG_4__SCAN_IN), .B1(n7010), .Y(n7023));
  OAI21X1 g03874(.A0(n7009), .A1(n7022), .B0(n7023), .Y(P3_U2763));
  INVX1   g03875(.A(P3_EAX_REG_5__SCAN_IN), .Y(n7025));
  AOI22X1 g03876(.A0(n7007), .A1(P3_DATAO_REG_5__SCAN_IN), .B0(P3_LWORD_REG_5__SCAN_IN), .B1(n7010), .Y(n7026));
  OAI21X1 g03877(.A0(n7009), .A1(n7025), .B0(n7026), .Y(P3_U2762));
  INVX1   g03878(.A(P3_EAX_REG_6__SCAN_IN), .Y(n7028));
  AOI22X1 g03879(.A0(n7007), .A1(P3_DATAO_REG_6__SCAN_IN), .B0(P3_LWORD_REG_6__SCAN_IN), .B1(n7010), .Y(n7029));
  OAI21X1 g03880(.A0(n7009), .A1(n7028), .B0(n7029), .Y(P3_U2761));
  NAND3X1 g03881(.A(n7006), .B(P3_EAX_REG_7__SCAN_IN), .C(P3_STATE2_REG_0__SCAN_IN), .Y(n7031));
  AOI22X1 g03882(.A0(n7007), .A1(P3_DATAO_REG_7__SCAN_IN), .B0(P3_LWORD_REG_7__SCAN_IN), .B1(n7010), .Y(n7032));
  NAND2X1 g03883(.A(n7032), .B(n7031), .Y(P3_U2760));
  INVX1   g03884(.A(P3_EAX_REG_8__SCAN_IN), .Y(n7034));
  AOI22X1 g03885(.A0(n7007), .A1(P3_DATAO_REG_8__SCAN_IN), .B0(P3_LWORD_REG_8__SCAN_IN), .B1(n7010), .Y(n7035));
  OAI21X1 g03886(.A0(n7009), .A1(n7034), .B0(n7035), .Y(P3_U2759));
  INVX1   g03887(.A(P3_EAX_REG_9__SCAN_IN), .Y(n7037));
  AOI22X1 g03888(.A0(n7007), .A1(P3_DATAO_REG_9__SCAN_IN), .B0(P3_LWORD_REG_9__SCAN_IN), .B1(n7010), .Y(n7038));
  OAI21X1 g03889(.A0(n7009), .A1(n7037), .B0(n7038), .Y(P3_U2758));
  INVX1   g03890(.A(P3_EAX_REG_10__SCAN_IN), .Y(n7040));
  AOI22X1 g03891(.A0(n7007), .A1(P3_DATAO_REG_10__SCAN_IN), .B0(P3_LWORD_REG_10__SCAN_IN), .B1(n7010), .Y(n7041));
  OAI21X1 g03892(.A0(n7009), .A1(n7040), .B0(n7041), .Y(P3_U2757));
  INVX1   g03893(.A(P3_EAX_REG_11__SCAN_IN), .Y(n7043));
  AOI22X1 g03894(.A0(n7007), .A1(P3_DATAO_REG_11__SCAN_IN), .B0(P3_LWORD_REG_11__SCAN_IN), .B1(n7010), .Y(n7044));
  OAI21X1 g03895(.A0(n7009), .A1(n7043), .B0(n7044), .Y(P3_U2756));
  NAND3X1 g03896(.A(n7006), .B(P3_EAX_REG_12__SCAN_IN), .C(P3_STATE2_REG_0__SCAN_IN), .Y(n7046));
  AOI22X1 g03897(.A0(n7007), .A1(P3_DATAO_REG_12__SCAN_IN), .B0(P3_LWORD_REG_12__SCAN_IN), .B1(n7010), .Y(n7047));
  NAND2X1 g03898(.A(n7047), .B(n7046), .Y(P3_U2755));
  INVX1   g03899(.A(P3_EAX_REG_13__SCAN_IN), .Y(n7049));
  AOI22X1 g03900(.A0(n7007), .A1(P3_DATAO_REG_13__SCAN_IN), .B0(P3_LWORD_REG_13__SCAN_IN), .B1(n7010), .Y(n7050));
  OAI21X1 g03901(.A0(n7009), .A1(n7049), .B0(n7050), .Y(P3_U2754));
  INVX1   g03902(.A(P3_EAX_REG_14__SCAN_IN), .Y(n7052));
  AOI22X1 g03903(.A0(n7007), .A1(P3_DATAO_REG_14__SCAN_IN), .B0(P3_LWORD_REG_14__SCAN_IN), .B1(n7010), .Y(n7053));
  OAI21X1 g03904(.A0(n7009), .A1(n7052), .B0(n7053), .Y(P3_U2753));
  INVX1   g03905(.A(P3_EAX_REG_15__SCAN_IN), .Y(n7055));
  AOI22X1 g03906(.A0(n7007), .A1(P3_DATAO_REG_15__SCAN_IN), .B0(P3_LWORD_REG_15__SCAN_IN), .B1(n7010), .Y(n7056));
  OAI21X1 g03907(.A0(n7009), .A1(n7055), .B0(n7056), .Y(P3_U2752));
  INVX1   g03908(.A(P3_EAX_REG_16__SCAN_IN), .Y(n7058));
  NAND3X1 g03909(.A(n7006), .B(n3699), .C(P3_STATE2_REG_0__SCAN_IN), .Y(n7059));
  AOI22X1 g03910(.A0(n7007), .A1(P3_DATAO_REG_16__SCAN_IN), .B0(P3_UWORD_REG_0__SCAN_IN), .B1(n7010), .Y(n7060));
  OAI21X1 g03911(.A0(n7059), .A1(n7058), .B0(n7060), .Y(P3_U2751));
  NAND4X1 g03912(.A(n3699), .B(P3_EAX_REG_17__SCAN_IN), .C(P3_STATE2_REG_0__SCAN_IN), .D(n7006), .Y(n7062));
  AOI22X1 g03913(.A0(n7007), .A1(P3_DATAO_REG_17__SCAN_IN), .B0(P3_UWORD_REG_1__SCAN_IN), .B1(n7010), .Y(n7063));
  NAND2X1 g03914(.A(n7063), .B(n7062), .Y(P3_U2750));
  INVX1   g03915(.A(P3_EAX_REG_18__SCAN_IN), .Y(n7065));
  AOI22X1 g03916(.A0(n7007), .A1(P3_DATAO_REG_18__SCAN_IN), .B0(P3_UWORD_REG_2__SCAN_IN), .B1(n7010), .Y(n7066));
  OAI21X1 g03917(.A0(n7059), .A1(n7065), .B0(n7066), .Y(P3_U2749));
  INVX1   g03918(.A(P3_EAX_REG_19__SCAN_IN), .Y(n7068));
  AOI22X1 g03919(.A0(n7007), .A1(P3_DATAO_REG_19__SCAN_IN), .B0(P3_UWORD_REG_3__SCAN_IN), .B1(n7010), .Y(n7069));
  OAI21X1 g03920(.A0(n7059), .A1(n7068), .B0(n7069), .Y(P3_U2748));
  INVX1   g03921(.A(P3_EAX_REG_20__SCAN_IN), .Y(n7071));
  AOI22X1 g03922(.A0(n7007), .A1(P3_DATAO_REG_20__SCAN_IN), .B0(P3_UWORD_REG_4__SCAN_IN), .B1(n7010), .Y(n7072));
  OAI21X1 g03923(.A0(n7059), .A1(n7071), .B0(n7072), .Y(P3_U2747));
  INVX1   g03924(.A(P3_EAX_REG_21__SCAN_IN), .Y(n7074));
  AOI22X1 g03925(.A0(n7007), .A1(P3_DATAO_REG_21__SCAN_IN), .B0(P3_UWORD_REG_5__SCAN_IN), .B1(n7010), .Y(n7075));
  OAI21X1 g03926(.A0(n7059), .A1(n7074), .B0(n7075), .Y(P3_U2746));
  NAND4X1 g03927(.A(n3699), .B(P3_EAX_REG_22__SCAN_IN), .C(P3_STATE2_REG_0__SCAN_IN), .D(n7006), .Y(n7077));
  AOI22X1 g03928(.A0(n7007), .A1(P3_DATAO_REG_22__SCAN_IN), .B0(P3_UWORD_REG_6__SCAN_IN), .B1(n7010), .Y(n7078));
  NAND2X1 g03929(.A(n7078), .B(n7077), .Y(P3_U2745));
  INVX1   g03930(.A(P3_EAX_REG_23__SCAN_IN), .Y(n7080));
  AOI22X1 g03931(.A0(n7007), .A1(P3_DATAO_REG_23__SCAN_IN), .B0(P3_UWORD_REG_7__SCAN_IN), .B1(n7010), .Y(n7081));
  OAI21X1 g03932(.A0(n7059), .A1(n7080), .B0(n7081), .Y(P3_U2744));
  INVX1   g03933(.A(P3_EAX_REG_24__SCAN_IN), .Y(n7083));
  AOI22X1 g03934(.A0(n7007), .A1(P3_DATAO_REG_24__SCAN_IN), .B0(P3_UWORD_REG_8__SCAN_IN), .B1(n7010), .Y(n7084));
  OAI21X1 g03935(.A0(n7059), .A1(n7083), .B0(n7084), .Y(P3_U2743));
  INVX1   g03936(.A(P3_EAX_REG_25__SCAN_IN), .Y(n7086));
  AOI22X1 g03937(.A0(n7007), .A1(P3_DATAO_REG_25__SCAN_IN), .B0(P3_UWORD_REG_9__SCAN_IN), .B1(n7010), .Y(n7087));
  OAI21X1 g03938(.A0(n7059), .A1(n7086), .B0(n7087), .Y(P3_U2742));
  NAND4X1 g03939(.A(n3699), .B(P3_EAX_REG_26__SCAN_IN), .C(P3_STATE2_REG_0__SCAN_IN), .D(n7006), .Y(n7089));
  AOI22X1 g03940(.A0(n7007), .A1(P3_DATAO_REG_26__SCAN_IN), .B0(P3_UWORD_REG_10__SCAN_IN), .B1(n7010), .Y(n7090));
  NAND2X1 g03941(.A(n7090), .B(n7089), .Y(P3_U2741));
  INVX1   g03942(.A(P3_EAX_REG_27__SCAN_IN), .Y(n7092));
  AOI22X1 g03943(.A0(n7007), .A1(P3_DATAO_REG_27__SCAN_IN), .B0(P3_UWORD_REG_11__SCAN_IN), .B1(n7010), .Y(n7093));
  OAI21X1 g03944(.A0(n7059), .A1(n7092), .B0(n7093), .Y(P3_U2740));
  INVX1   g03945(.A(P3_EAX_REG_28__SCAN_IN), .Y(n7095));
  AOI22X1 g03946(.A0(n7007), .A1(P3_DATAO_REG_28__SCAN_IN), .B0(P3_UWORD_REG_12__SCAN_IN), .B1(n7010), .Y(n7096));
  OAI21X1 g03947(.A0(n7059), .A1(n7095), .B0(n7096), .Y(P3_U2739));
  INVX1   g03948(.A(P3_EAX_REG_29__SCAN_IN), .Y(n7098));
  AOI22X1 g03949(.A0(n7007), .A1(P3_DATAO_REG_29__SCAN_IN), .B0(P3_UWORD_REG_13__SCAN_IN), .B1(n7010), .Y(n7099));
  OAI21X1 g03950(.A0(n7059), .A1(n7098), .B0(n7099), .Y(P3_U2738));
  INVX1   g03951(.A(P3_EAX_REG_30__SCAN_IN), .Y(n7101));
  AOI22X1 g03952(.A0(n7007), .A1(P3_DATAO_REG_30__SCAN_IN), .B0(P3_UWORD_REG_14__SCAN_IN), .B1(n7010), .Y(n7102));
  OAI21X1 g03953(.A0(n7059), .A1(n7101), .B0(n7102), .Y(P3_U2737));
  NOR2X1  g03954(.A(n7006), .B(n2964), .Y(P3_U2736));
  AOI21X1 g03955(.A0(n3835), .A1(n3723), .B0(n4905), .Y(n7105));
  NAND4X1 g03956(.A(n3667), .B(n3774), .C(BUF2_REG_0__SCAN_IN), .D(n7105), .Y(n7106));
  INVX1   g03957(.A(n7105), .Y(n7107));
  NOR2X1  g03958(.A(n7107), .B(n3667), .Y(n7108));
  OAI21X1 g03959(.A0(n5011), .A1(n4998), .B0(n7108), .Y(n7109));
  NOR2X1  g03960(.A(n7105), .B(n7004), .Y(n7110));
  NOR2X1  g03961(.A(n7107), .B(n3774), .Y(n7111));
  AOI21X1 g03962(.A0(n7111), .A1(n7004), .B0(n7110), .Y(n7112));
  NAND3X1 g03963(.A(n7112), .B(n7109), .C(n7106), .Y(P3_U2735));
  NAND4X1 g03964(.A(n3667), .B(n3774), .C(BUF2_REG_1__SCAN_IN), .D(n7105), .Y(n7114));
  NAND3X1 g03965(.A(n7105), .B(n5076), .C(n3666), .Y(n7115));
  XOR2X1  g03966(.A(P3_EAX_REG_1__SCAN_IN), .B(P3_EAX_REG_0__SCAN_IN), .Y(n7116));
  AOI22X1 g03967(.A0(n7111), .A1(n7116), .B0(n7107), .B1(P3_EAX_REG_1__SCAN_IN), .Y(n7117));
  NAND3X1 g03968(.A(n7117), .B(n7115), .C(n7114), .Y(P3_U2734));
  NAND4X1 g03969(.A(n3667), .B(n3774), .C(BUF2_REG_2__SCAN_IN), .D(n7105), .Y(n7119));
  NAND3X1 g03970(.A(n7105), .B(n5121), .C(n3666), .Y(n7120));
  NAND2X1 g03971(.A(P3_EAX_REG_1__SCAN_IN), .B(P3_EAX_REG_0__SCAN_IN), .Y(n7121));
  XOR2X1  g03972(.A(n7121), .B(n7016), .Y(n7122));
  AOI22X1 g03973(.A0(n7111), .A1(n7122), .B0(n7107), .B1(P3_EAX_REG_2__SCAN_IN), .Y(n7123));
  NAND3X1 g03974(.A(n7123), .B(n7120), .C(n7119), .Y(P3_U2733));
  NAND4X1 g03975(.A(n3667), .B(n3774), .C(BUF2_REG_3__SCAN_IN), .D(n7105), .Y(n7125));
  NAND3X1 g03976(.A(n7105), .B(n5207), .C(n3666), .Y(n7126));
  NOR2X1  g03977(.A(n7121), .B(n7016), .Y(n7127));
  XOR2X1  g03978(.A(n7127), .B(P3_EAX_REG_3__SCAN_IN), .Y(n7128));
  AOI22X1 g03979(.A0(n7111), .A1(n7128), .B0(n7107), .B1(P3_EAX_REG_3__SCAN_IN), .Y(n7129));
  NAND3X1 g03980(.A(n7129), .B(n7126), .C(n7125), .Y(P3_U2732));
  NAND4X1 g03981(.A(n3667), .B(n3774), .C(BUF2_REG_4__SCAN_IN), .D(n7105), .Y(n7131));
  NAND3X1 g03982(.A(n7105), .B(n5275), .C(n3666), .Y(n7132));
  NAND4X1 g03983(.A(P3_EAX_REG_2__SCAN_IN), .B(P3_EAX_REG_1__SCAN_IN), .C(P3_EAX_REG_0__SCAN_IN), .D(P3_EAX_REG_3__SCAN_IN), .Y(n7133));
  XOR2X1  g03984(.A(n7133), .B(n7022), .Y(n7134));
  AOI22X1 g03985(.A0(n7111), .A1(n7134), .B0(n7107), .B1(P3_EAX_REG_4__SCAN_IN), .Y(n7135));
  NAND3X1 g03986(.A(n7135), .B(n7132), .C(n7131), .Y(P3_U2731));
  NAND4X1 g03987(.A(n3667), .B(n3774), .C(BUF2_REG_5__SCAN_IN), .D(n7105), .Y(n7137));
  NAND3X1 g03988(.A(n7105), .B(n5412), .C(n3666), .Y(n7138));
  NOR4X1  g03989(.A(n7022), .B(n7019), .C(n7016), .D(n7121), .Y(n7139));
  XOR2X1  g03990(.A(n7139), .B(P3_EAX_REG_5__SCAN_IN), .Y(n7140));
  AOI22X1 g03991(.A0(n7111), .A1(n7140), .B0(n7107), .B1(P3_EAX_REG_5__SCAN_IN), .Y(n7141));
  NAND3X1 g03992(.A(n7141), .B(n7138), .C(n7137), .Y(P3_U2730));
  NAND4X1 g03993(.A(n3667), .B(n3774), .C(BUF2_REG_6__SCAN_IN), .D(n7105), .Y(n7143));
  OAI21X1 g03994(.A0(n5398), .A1(n5393), .B0(n7108), .Y(n7144));
  NAND2X1 g03995(.A(n7139), .B(P3_EAX_REG_5__SCAN_IN), .Y(n7145));
  XOR2X1  g03996(.A(n7145), .B(n7028), .Y(n7146));
  AOI22X1 g03997(.A0(n7111), .A1(n7146), .B0(n7107), .B1(P3_EAX_REG_6__SCAN_IN), .Y(n7147));
  NAND3X1 g03998(.A(n7147), .B(n7144), .C(n7143), .Y(P3_U2729));
  NAND4X1 g03999(.A(n3667), .B(n3774), .C(BUF2_REG_7__SCAN_IN), .D(n7105), .Y(n7149));
  NAND3X1 g04000(.A(n7105), .B(n5039), .C(n3666), .Y(n7150));
  INVX1   g04001(.A(n7139), .Y(n7151));
  NOR3X1  g04002(.A(n7151), .B(n7028), .C(n7025), .Y(n7152));
  XOR2X1  g04003(.A(n7152), .B(P3_EAX_REG_7__SCAN_IN), .Y(n7153));
  AOI22X1 g04004(.A0(n7111), .A1(n7153), .B0(n7107), .B1(P3_EAX_REG_7__SCAN_IN), .Y(n7154));
  NAND3X1 g04005(.A(n7154), .B(n7150), .C(n7149), .Y(P3_U2728));
  NAND4X1 g04006(.A(n3667), .B(n3774), .C(BUF2_REG_8__SCAN_IN), .D(n7105), .Y(n7156));
  INVX1   g04007(.A(P3_INSTQUEUE_REG_15__0__SCAN_IN), .Y(n7157));
  NAND4X1 g04008(.A(n3517), .B(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .D(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n7158));
  NAND4X1 g04009(.A(n3517), .B(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .D(n3541), .Y(n7159));
  OAI22X1 g04010(.A0(n7158), .A1(n7157), .B0(n4133), .B1(n7159), .Y(n7160));
  INVX1   g04011(.A(P3_INSTQUEUE_REG_13__0__SCAN_IN), .Y(n7161));
  NAND4X1 g04012(.A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n3515), .C(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .D(n3541), .Y(n7162));
  NAND4X1 g04013(.A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n3515), .C(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .D(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n7163));
  OAI22X1 g04014(.A0(n7162), .A1(n4253), .B0(n7161), .B1(n7163), .Y(n7164));
  INVX1   g04015(.A(P3_INSTQUEUE_REG_11__0__SCAN_IN), .Y(n7165));
  NAND4X1 g04016(.A(n3517), .B(n3515), .C(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .D(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n7166));
  NAND4X1 g04017(.A(n3517), .B(n3515), .C(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .D(n3541), .Y(n7167));
  OAI22X1 g04018(.A0(n7166), .A1(n7165), .B0(n4365), .B1(n7167), .Y(n7168));
  NAND4X1 g04019(.A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(n3535), .D(n3541), .Y(n7169));
  NAND4X1 g04020(.A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(n3535), .D(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n7170));
  OAI22X1 g04021(.A0(n7169), .A1(n4478), .B0(n3685), .B1(n7170), .Y(n7171));
  NOR4X1  g04022(.A(n7168), .B(n7164), .C(n7160), .D(n7171), .Y(n7172));
  INVX1   g04023(.A(P3_INSTQUEUE_REG_2__0__SCAN_IN), .Y(n7173));
  NAND4X1 g04024(.A(n3517), .B(n3515), .C(n3535), .D(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n7174));
  OAI22X1 g04025(.A0(n7174), .A1(n3686), .B0(n7173), .B1(n3551), .Y(n7176));
  INVX1   g04026(.A(P3_INSTQUEUE_REG_1__0__SCAN_IN), .Y(n7177));
  NAND4X1 g04027(.A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .D(n3541), .Y(n7178));
  NAND4X1 g04028(.A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .D(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n7179));
  OAI22X1 g04029(.A0(n7178), .A1(n3683), .B0(n7177), .B1(n7179), .Y(n7180));
  INVX1   g04030(.A(P3_INSTQUEUE_REG_7__0__SCAN_IN), .Y(n7181));
  NAND4X1 g04031(.A(n3517), .B(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(n3535), .D(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n7182));
  NAND4X1 g04032(.A(n3517), .B(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(n3535), .D(n3541), .Y(n7183));
  OAI22X1 g04033(.A0(n7182), .A1(n7181), .B0(n4589), .B1(n7183), .Y(n7184));
  INVX1   g04034(.A(P3_INSTQUEUE_REG_5__0__SCAN_IN), .Y(n7185));
  INVX1   g04035(.A(P3_INSTQUEUE_REG_4__0__SCAN_IN), .Y(n7186));
  NAND4X1 g04036(.A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n3515), .C(n3535), .D(n3541), .Y(n7187));
  NAND4X1 g04037(.A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n3515), .C(n3535), .D(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n7188));
  OAI22X1 g04038(.A0(n7187), .A1(n7186), .B0(n7185), .B1(n7188), .Y(n7189));
  NOR4X1  g04039(.A(n7184), .B(n7180), .C(n7176), .D(n7189), .Y(n7190));
  NAND2X1 g04040(.A(n7190), .B(n7172), .Y(n7191));
  NAND3X1 g04041(.A(n7191), .B(n7105), .C(n3666), .Y(n7192));
  NAND4X1 g04042(.A(P3_EAX_REG_7__SCAN_IN), .B(P3_EAX_REG_6__SCAN_IN), .C(P3_EAX_REG_5__SCAN_IN), .D(n7139), .Y(n7193));
  XOR2X1  g04043(.A(n7193), .B(n7034), .Y(n7194));
  AOI22X1 g04044(.A0(n7111), .A1(n7194), .B0(n7107), .B1(P3_EAX_REG_8__SCAN_IN), .Y(n7195));
  NAND3X1 g04045(.A(n7195), .B(n7192), .C(n7156), .Y(P3_U2727));
  NAND4X1 g04046(.A(n3667), .B(n3774), .C(BUF2_REG_9__SCAN_IN), .D(n7105), .Y(n7197));
  INVX1   g04047(.A(P3_INSTQUEUE_REG_15__1__SCAN_IN), .Y(n7198));
  OAI22X1 g04048(.A0(n7158), .A1(n7198), .B0(n4125), .B1(n7159), .Y(n7199));
  INVX1   g04049(.A(P3_INSTQUEUE_REG_13__1__SCAN_IN), .Y(n7200));
  OAI22X1 g04050(.A0(n7162), .A1(n4247), .B0(n7200), .B1(n7163), .Y(n7201));
  INVX1   g04051(.A(P3_INSTQUEUE_REG_11__1__SCAN_IN), .Y(n7202));
  OAI22X1 g04052(.A0(n7166), .A1(n7202), .B0(n4359), .B1(n7167), .Y(n7203));
  INVX1   g04053(.A(P3_INSTQUEUE_REG_9__1__SCAN_IN), .Y(n7204));
  OAI22X1 g04054(.A0(n7169), .A1(n4472), .B0(n7204), .B1(n7170), .Y(n7205));
  NOR4X1  g04055(.A(n7203), .B(n7201), .C(n7199), .D(n7205), .Y(n7206));
  INVX1   g04056(.A(P3_INSTQUEUE_REG_3__1__SCAN_IN), .Y(n7207));
  INVX1   g04057(.A(P3_INSTQUEUE_REG_2__1__SCAN_IN), .Y(n7208));
  OAI22X1 g04058(.A0(n7174), .A1(n7207), .B0(n7208), .B1(n3551), .Y(n7209));
  INVX1   g04059(.A(P3_INSTQUEUE_REG_1__1__SCAN_IN), .Y(n7210));
  OAI22X1 g04060(.A0(n7178), .A1(n3668), .B0(n7210), .B1(n7179), .Y(n7211));
  INVX1   g04061(.A(P3_INSTQUEUE_REG_7__1__SCAN_IN), .Y(n7212));
  OAI22X1 g04062(.A0(n7182), .A1(n7212), .B0(n4583), .B1(n7183), .Y(n7213));
  INVX1   g04063(.A(P3_INSTQUEUE_REG_5__1__SCAN_IN), .Y(n7214));
  INVX1   g04064(.A(P3_INSTQUEUE_REG_4__1__SCAN_IN), .Y(n7215));
  OAI22X1 g04065(.A0(n7187), .A1(n7215), .B0(n7214), .B1(n7188), .Y(n7216));
  NOR4X1  g04066(.A(n7213), .B(n7211), .C(n7209), .D(n7216), .Y(n7217));
  NAND2X1 g04067(.A(n7217), .B(n7206), .Y(n7218));
  NAND3X1 g04068(.A(n7218), .B(n7105), .C(n3666), .Y(n7219));
  NAND3X1 g04069(.A(n7152), .B(P3_EAX_REG_8__SCAN_IN), .C(P3_EAX_REG_7__SCAN_IN), .Y(n7220));
  XOR2X1  g04070(.A(n7220), .B(n7037), .Y(n7221));
  AOI22X1 g04071(.A0(n7111), .A1(n7221), .B0(n7107), .B1(P3_EAX_REG_9__SCAN_IN), .Y(n7222));
  NAND3X1 g04072(.A(n7222), .B(n7219), .C(n7197), .Y(P3_U2726));
  NAND4X1 g04073(.A(n3667), .B(n3774), .C(BUF2_REG_10__SCAN_IN), .D(n7105), .Y(n7224));
  INVX1   g04074(.A(P3_INSTQUEUE_REG_15__2__SCAN_IN), .Y(n7225));
  OAI22X1 g04075(.A0(n7158), .A1(n7225), .B0(n4117), .B1(n7159), .Y(n7226));
  INVX1   g04076(.A(P3_INSTQUEUE_REG_13__2__SCAN_IN), .Y(n7227));
  OAI22X1 g04077(.A0(n7162), .A1(n4241), .B0(n7227), .B1(n7163), .Y(n7228));
  INVX1   g04078(.A(P3_INSTQUEUE_REG_11__2__SCAN_IN), .Y(n7229));
  OAI22X1 g04079(.A0(n7166), .A1(n7229), .B0(n4353), .B1(n7167), .Y(n7230));
  OAI22X1 g04080(.A0(n7169), .A1(n4466), .B0(n3553), .B1(n7170), .Y(n7231));
  NOR4X1  g04081(.A(n7230), .B(n7228), .C(n7226), .D(n7231), .Y(n7232));
  INVX1   g04082(.A(P3_INSTQUEUE_REG_2__2__SCAN_IN), .Y(n7233));
  OAI22X1 g04083(.A0(n7174), .A1(n3554), .B0(n7233), .B1(n3551), .Y(n7234));
  INVX1   g04084(.A(P3_INSTQUEUE_REG_1__2__SCAN_IN), .Y(n7235));
  OAI22X1 g04085(.A0(n7178), .A1(n3549), .B0(n7235), .B1(n7179), .Y(n7236));
  INVX1   g04086(.A(P3_INSTQUEUE_REG_7__2__SCAN_IN), .Y(n7237));
  OAI22X1 g04087(.A0(n7182), .A1(n7237), .B0(n4577), .B1(n7183), .Y(n7238));
  INVX1   g04088(.A(P3_INSTQUEUE_REG_5__2__SCAN_IN), .Y(n7239));
  INVX1   g04089(.A(P3_INSTQUEUE_REG_4__2__SCAN_IN), .Y(n7240));
  OAI22X1 g04090(.A0(n7187), .A1(n7240), .B0(n7239), .B1(n7188), .Y(n7241));
  NOR4X1  g04091(.A(n7238), .B(n7236), .C(n7234), .D(n7241), .Y(n7242));
  NAND2X1 g04092(.A(n7242), .B(n7232), .Y(n7243));
  NAND3X1 g04093(.A(n7243), .B(n7105), .C(n3666), .Y(n7244));
  NAND4X1 g04094(.A(P3_EAX_REG_9__SCAN_IN), .B(P3_EAX_REG_8__SCAN_IN), .C(P3_EAX_REG_7__SCAN_IN), .D(n7152), .Y(n7245));
  XOR2X1  g04095(.A(n7245), .B(n7040), .Y(n7246));
  AOI22X1 g04096(.A0(n7111), .A1(n7246), .B0(n7107), .B1(P3_EAX_REG_10__SCAN_IN), .Y(n7247));
  NAND3X1 g04097(.A(n7247), .B(n7244), .C(n7224), .Y(P3_U2725));
  NAND4X1 g04098(.A(n3667), .B(n3774), .C(BUF2_REG_11__SCAN_IN), .D(n7105), .Y(n7249));
  INVX1   g04099(.A(P3_INSTQUEUE_REG_15__3__SCAN_IN), .Y(n7250));
  OAI22X1 g04100(.A0(n7158), .A1(n7250), .B0(n4109), .B1(n7159), .Y(n7251));
  INVX1   g04101(.A(P3_INSTQUEUE_REG_13__3__SCAN_IN), .Y(n7252));
  OAI22X1 g04102(.A0(n7162), .A1(n4235), .B0(n7252), .B1(n7163), .Y(n7253));
  INVX1   g04103(.A(P3_INSTQUEUE_REG_11__3__SCAN_IN), .Y(n7254));
  OAI22X1 g04104(.A0(n7166), .A1(n7254), .B0(n4347), .B1(n7167), .Y(n7255));
  OAI22X1 g04105(.A0(n7169), .A1(n4460), .B0(n3603), .B1(n7170), .Y(n7256));
  NOR4X1  g04106(.A(n7255), .B(n7253), .C(n7251), .D(n7256), .Y(n7257));
  INVX1   g04107(.A(P3_INSTQUEUE_REG_2__3__SCAN_IN), .Y(n7258));
  OAI22X1 g04108(.A0(n7174), .A1(n3604), .B0(n7258), .B1(n3551), .Y(n7259));
  INVX1   g04109(.A(P3_INSTQUEUE_REG_1__3__SCAN_IN), .Y(n7260));
  OAI22X1 g04110(.A0(n7178), .A1(n3601), .B0(n7260), .B1(n7179), .Y(n7261));
  INVX1   g04111(.A(P3_INSTQUEUE_REG_7__3__SCAN_IN), .Y(n7262));
  OAI22X1 g04112(.A0(n7182), .A1(n7262), .B0(n4571), .B1(n7183), .Y(n7263));
  INVX1   g04113(.A(P3_INSTQUEUE_REG_5__3__SCAN_IN), .Y(n7264));
  INVX1   g04114(.A(P3_INSTQUEUE_REG_4__3__SCAN_IN), .Y(n7265));
  OAI22X1 g04115(.A0(n7187), .A1(n7265), .B0(n7264), .B1(n7188), .Y(n7266));
  NOR4X1  g04116(.A(n7263), .B(n7261), .C(n7259), .D(n7266), .Y(n7267));
  NAND2X1 g04117(.A(n7267), .B(n7257), .Y(n7268));
  NAND3X1 g04118(.A(n7268), .B(n7105), .C(n3666), .Y(n7269));
  NOR3X1  g04119(.A(n7220), .B(n7040), .C(n7037), .Y(n7270));
  XOR2X1  g04120(.A(n7270), .B(P3_EAX_REG_11__SCAN_IN), .Y(n7271));
  AOI22X1 g04121(.A0(n7111), .A1(n7271), .B0(n7107), .B1(P3_EAX_REG_11__SCAN_IN), .Y(n7272));
  NAND3X1 g04122(.A(n7272), .B(n7269), .C(n7249), .Y(P3_U2724));
  NAND4X1 g04123(.A(n3667), .B(n3774), .C(BUF2_REG_12__SCAN_IN), .D(n7105), .Y(n7274));
  INVX1   g04124(.A(P3_INSTQUEUE_REG_15__4__SCAN_IN), .Y(n7275));
  OAI22X1 g04125(.A0(n7158), .A1(n7275), .B0(n4101), .B1(n7159), .Y(n7276));
  INVX1   g04126(.A(P3_INSTQUEUE_REG_13__4__SCAN_IN), .Y(n7277));
  OAI22X1 g04127(.A0(n7162), .A1(n4229), .B0(n7277), .B1(n7163), .Y(n7278));
  INVX1   g04128(.A(P3_INSTQUEUE_REG_11__4__SCAN_IN), .Y(n7279));
  OAI22X1 g04129(.A0(n7166), .A1(n7279), .B0(n4341), .B1(n7167), .Y(n7280));
  OAI22X1 g04130(.A0(n7169), .A1(n4454), .B0(n3621), .B1(n7170), .Y(n7281));
  NOR4X1  g04131(.A(n7280), .B(n7278), .C(n7276), .D(n7281), .Y(n7282));
  INVX1   g04132(.A(P3_INSTQUEUE_REG_2__4__SCAN_IN), .Y(n7283));
  OAI22X1 g04133(.A0(n7174), .A1(n3622), .B0(n7283), .B1(n3551), .Y(n7284));
  INVX1   g04134(.A(P3_INSTQUEUE_REG_1__4__SCAN_IN), .Y(n7285));
  OAI22X1 g04135(.A0(n7178), .A1(n3619), .B0(n7285), .B1(n7179), .Y(n7286));
  INVX1   g04136(.A(P3_INSTQUEUE_REG_7__4__SCAN_IN), .Y(n7287));
  OAI22X1 g04137(.A0(n7182), .A1(n7287), .B0(n4565), .B1(n7183), .Y(n7288));
  INVX1   g04138(.A(P3_INSTQUEUE_REG_5__4__SCAN_IN), .Y(n7289));
  INVX1   g04139(.A(P3_INSTQUEUE_REG_4__4__SCAN_IN), .Y(n7290));
  OAI22X1 g04140(.A0(n7187), .A1(n7290), .B0(n7289), .B1(n7188), .Y(n7291));
  NOR4X1  g04141(.A(n7288), .B(n7286), .C(n7284), .D(n7291), .Y(n7292));
  NAND2X1 g04142(.A(n7292), .B(n7282), .Y(n7293));
  NAND3X1 g04143(.A(n7293), .B(n7105), .C(n3666), .Y(n7294));
  NOR4X1  g04144(.A(n7043), .B(n7040), .C(n7037), .D(n7220), .Y(n7295));
  XOR2X1  g04145(.A(n7295), .B(P3_EAX_REG_12__SCAN_IN), .Y(n7296));
  AOI22X1 g04146(.A0(n7111), .A1(n7296), .B0(n7107), .B1(P3_EAX_REG_12__SCAN_IN), .Y(n7297));
  NAND3X1 g04147(.A(n7297), .B(n7294), .C(n7274), .Y(P3_U2723));
  NAND4X1 g04148(.A(n3667), .B(n3774), .C(BUF2_REG_13__SCAN_IN), .D(n7105), .Y(n7299));
  INVX1   g04149(.A(P3_INSTQUEUE_REG_15__5__SCAN_IN), .Y(n7300));
  OAI22X1 g04150(.A0(n7158), .A1(n7300), .B0(n4093), .B1(n7159), .Y(n7301));
  INVX1   g04151(.A(P3_INSTQUEUE_REG_13__5__SCAN_IN), .Y(n7302));
  OAI22X1 g04152(.A0(n7162), .A1(n4223), .B0(n7302), .B1(n7163), .Y(n7303));
  INVX1   g04153(.A(P3_INSTQUEUE_REG_11__5__SCAN_IN), .Y(n7304));
  OAI22X1 g04154(.A0(n7166), .A1(n7304), .B0(n4335), .B1(n7167), .Y(n7305));
  OAI22X1 g04155(.A0(n7169), .A1(n4448), .B0(n3637), .B1(n7170), .Y(n7306));
  NOR4X1  g04156(.A(n7305), .B(n7303), .C(n7301), .D(n7306), .Y(n7307));
  INVX1   g04157(.A(P3_INSTQUEUE_REG_2__5__SCAN_IN), .Y(n7308));
  OAI22X1 g04158(.A0(n7174), .A1(n3638), .B0(n7308), .B1(n3551), .Y(n7309));
  INVX1   g04159(.A(P3_INSTQUEUE_REG_1__5__SCAN_IN), .Y(n7310));
  OAI22X1 g04160(.A0(n7178), .A1(n3635), .B0(n7310), .B1(n7179), .Y(n7311));
  INVX1   g04161(.A(P3_INSTQUEUE_REG_7__5__SCAN_IN), .Y(n7312));
  OAI22X1 g04162(.A0(n7182), .A1(n7312), .B0(n4559), .B1(n7183), .Y(n7313));
  INVX1   g04163(.A(P3_INSTQUEUE_REG_5__5__SCAN_IN), .Y(n7314));
  INVX1   g04164(.A(P3_INSTQUEUE_REG_4__5__SCAN_IN), .Y(n7315));
  OAI22X1 g04165(.A0(n7187), .A1(n7315), .B0(n7314), .B1(n7188), .Y(n7316));
  NOR4X1  g04166(.A(n7313), .B(n7311), .C(n7309), .D(n7316), .Y(n7317));
  NAND2X1 g04167(.A(n7317), .B(n7307), .Y(n7318));
  NAND3X1 g04168(.A(n7318), .B(n7105), .C(n3666), .Y(n7319));
  NAND3X1 g04169(.A(n7270), .B(P3_EAX_REG_12__SCAN_IN), .C(P3_EAX_REG_11__SCAN_IN), .Y(n7320));
  XOR2X1  g04170(.A(n7320), .B(n7049), .Y(n7321));
  AOI22X1 g04171(.A0(n7111), .A1(n7321), .B0(n7107), .B1(P3_EAX_REG_13__SCAN_IN), .Y(n7322));
  NAND3X1 g04172(.A(n7322), .B(n7319), .C(n7299), .Y(P3_U2722));
  NAND4X1 g04173(.A(n3667), .B(n3774), .C(BUF2_REG_14__SCAN_IN), .D(n7105), .Y(n7324));
  INVX1   g04174(.A(P3_INSTQUEUE_REG_15__6__SCAN_IN), .Y(n7325));
  OAI22X1 g04175(.A0(n7158), .A1(n7325), .B0(n4085), .B1(n7159), .Y(n7326));
  INVX1   g04176(.A(P3_INSTQUEUE_REG_13__6__SCAN_IN), .Y(n7327));
  OAI22X1 g04177(.A0(n7162), .A1(n4217), .B0(n7327), .B1(n7163), .Y(n7328));
  INVX1   g04178(.A(P3_INSTQUEUE_REG_11__6__SCAN_IN), .Y(n7329));
  OAI22X1 g04179(.A0(n7166), .A1(n7329), .B0(n4329), .B1(n7167), .Y(n7330));
  OAI22X1 g04180(.A0(n7169), .A1(n4442), .B0(n3653), .B1(n7170), .Y(n7331));
  NOR4X1  g04181(.A(n7330), .B(n7328), .C(n7326), .D(n7331), .Y(n7332));
  INVX1   g04182(.A(P3_INSTQUEUE_REG_2__6__SCAN_IN), .Y(n7333));
  OAI22X1 g04183(.A0(n7174), .A1(n3654), .B0(n7333), .B1(n3551), .Y(n7334));
  INVX1   g04184(.A(P3_INSTQUEUE_REG_1__6__SCAN_IN), .Y(n7335));
  OAI22X1 g04185(.A0(n7178), .A1(n3651), .B0(n7335), .B1(n7179), .Y(n7336));
  INVX1   g04186(.A(P3_INSTQUEUE_REG_7__6__SCAN_IN), .Y(n7337));
  OAI22X1 g04187(.A0(n7182), .A1(n7337), .B0(n4553), .B1(n7183), .Y(n7338));
  INVX1   g04188(.A(P3_INSTQUEUE_REG_5__6__SCAN_IN), .Y(n7339));
  INVX1   g04189(.A(P3_INSTQUEUE_REG_4__6__SCAN_IN), .Y(n7340));
  OAI22X1 g04190(.A0(n7187), .A1(n7340), .B0(n7339), .B1(n7188), .Y(n7341));
  NOR4X1  g04191(.A(n7338), .B(n7336), .C(n7334), .D(n7341), .Y(n7342));
  NAND2X1 g04192(.A(n7342), .B(n7332), .Y(n7343));
  NAND3X1 g04193(.A(n7343), .B(n7105), .C(n3666), .Y(n7344));
  NAND4X1 g04194(.A(P3_EAX_REG_13__SCAN_IN), .B(P3_EAX_REG_12__SCAN_IN), .C(P3_EAX_REG_11__SCAN_IN), .D(n7270), .Y(n7345));
  XOR2X1  g04195(.A(n7345), .B(n7052), .Y(n7346));
  AOI22X1 g04196(.A0(n7111), .A1(n7346), .B0(n7107), .B1(P3_EAX_REG_14__SCAN_IN), .Y(n7347));
  NAND3X1 g04197(.A(n7347), .B(n7344), .C(n7324), .Y(P3_U2721));
  NAND4X1 g04198(.A(n3667), .B(n3774), .C(BUF2_REG_15__SCAN_IN), .D(n7105), .Y(n7349));
  INVX1   g04199(.A(P3_INSTQUEUE_REG_15__7__SCAN_IN), .Y(n7350));
  OAI22X1 g04200(.A0(n7158), .A1(n7350), .B0(n4062), .B1(n7159), .Y(n7351));
  INVX1   g04201(.A(P3_INSTQUEUE_REG_13__7__SCAN_IN), .Y(n7352));
  OAI22X1 g04202(.A0(n7162), .A1(n4193), .B0(n7352), .B1(n7163), .Y(n7353));
  INVX1   g04203(.A(P3_INSTQUEUE_REG_11__7__SCAN_IN), .Y(n7354));
  OAI22X1 g04204(.A0(n7166), .A1(n7354), .B0(n4310), .B1(n7167), .Y(n7355));
  OAI22X1 g04205(.A0(n7169), .A1(n4422), .B0(n3587), .B1(n7170), .Y(n7356));
  NOR4X1  g04206(.A(n7355), .B(n7353), .C(n7351), .D(n7356), .Y(n7357));
  INVX1   g04207(.A(P3_INSTQUEUE_REG_2__7__SCAN_IN), .Y(n7358));
  OAI22X1 g04208(.A0(n7174), .A1(n3588), .B0(n7358), .B1(n3551), .Y(n7359));
  INVX1   g04209(.A(P3_INSTQUEUE_REG_1__7__SCAN_IN), .Y(n7360));
  OAI22X1 g04210(.A0(n7178), .A1(n3585), .B0(n7360), .B1(n7179), .Y(n7361));
  INVX1   g04211(.A(P3_INSTQUEUE_REG_7__7__SCAN_IN), .Y(n7362));
  OAI22X1 g04212(.A0(n7182), .A1(n7362), .B0(n4534), .B1(n7183), .Y(n7363));
  INVX1   g04213(.A(P3_INSTQUEUE_REG_5__7__SCAN_IN), .Y(n7364));
  INVX1   g04214(.A(P3_INSTQUEUE_REG_4__7__SCAN_IN), .Y(n7365));
  OAI22X1 g04215(.A0(n7187), .A1(n7365), .B0(n7364), .B1(n7188), .Y(n7366));
  NOR4X1  g04216(.A(n7363), .B(n7361), .C(n7359), .D(n7366), .Y(n7367));
  NAND2X1 g04217(.A(n7367), .B(n7357), .Y(n7368));
  NAND3X1 g04218(.A(n7368), .B(n7105), .C(n3666), .Y(n7369));
  NOR3X1  g04219(.A(n7320), .B(n7052), .C(n7049), .Y(n7370));
  XOR2X1  g04220(.A(n7370), .B(P3_EAX_REG_15__SCAN_IN), .Y(n7371));
  AOI22X1 g04221(.A0(n7111), .A1(n7371), .B0(n7107), .B1(P3_EAX_REG_15__SCAN_IN), .Y(n7372));
  NAND3X1 g04222(.A(n7372), .B(n7369), .C(n7349), .Y(P3_U2720));
  OAI22X1 g04223(.A0(n7183), .A1(n7181), .B0(n4589), .B1(n7188), .Y(n7378));
  OAI22X1 g04224(.A0(n7174), .A1(n7186), .B0(n7185), .B1(n7187), .Y(n7383));
  OAI22X1 g04225(.A0(n3551), .A1(n3686), .B0(n7173), .B1(n7179), .Y(n7388));
  OAI22X1 g04226(.A0(n7158), .A1(n3683), .B0(n7177), .B1(n7178), .Y(n7393));
  NOR4X1  g04227(.A(n7388), .B(n7383), .C(n7378), .D(n7393), .Y(n7394));
  OAI22X1 g04228(.A0(n7167), .A1(n7165), .B0(n4365), .B1(n7170), .Y(n7399));
  OAI22X1 g04229(.A0(n7182), .A1(n4478), .B0(n3685), .B1(n7169), .Y(n7404));
  OAI22X1 g04230(.A0(n7159), .A1(n7157), .B0(n4133), .B1(n7163), .Y(n7409));
  OAI22X1 g04231(.A0(n7166), .A1(n4253), .B0(n7161), .B1(n7162), .Y(n7414));
  NOR4X1  g04232(.A(n7409), .B(n7404), .C(n7399), .D(n7414), .Y(n7415));
  NAND2X1 g04233(.A(n7415), .B(n7394), .Y(n7416));
  NAND3X1 g04234(.A(n7416), .B(n7105), .C(n3666), .Y(n7417));
  NOR4X1  g04235(.A(n7055), .B(n7052), .C(n7049), .D(n7320), .Y(n7418));
  XOR2X1  g04236(.A(n7418), .B(P3_EAX_REG_16__SCAN_IN), .Y(n7419));
  AOI22X1 g04237(.A0(n7111), .A1(n7419), .B0(n7107), .B1(P3_EAX_REG_16__SCAN_IN), .Y(n7420));
  NOR3X1  g04238(.A(n7107), .B(n3708), .C(n3600), .Y(n7421));
  NOR3X1  g04239(.A(n7107), .B(n3714), .C(n3600), .Y(n7422));
  AOI22X1 g04240(.A0(n7421), .A1(BUF2_REG_16__SCAN_IN), .B0(BUF2_REG_0__SCAN_IN), .B1(n7422), .Y(n7423));
  NAND3X1 g04241(.A(n7423), .B(n7420), .C(n7417), .Y(P3_U2719));
  OAI22X1 g04242(.A0(n7183), .A1(n7212), .B0(n4583), .B1(n7188), .Y(n7425));
  OAI22X1 g04243(.A0(n7174), .A1(n7215), .B0(n7214), .B1(n7187), .Y(n7426));
  OAI22X1 g04244(.A0(n3551), .A1(n7207), .B0(n7208), .B1(n7179), .Y(n7427));
  OAI22X1 g04245(.A0(n7158), .A1(n3668), .B0(n7210), .B1(n7178), .Y(n7428));
  NOR4X1  g04246(.A(n7427), .B(n7426), .C(n7425), .D(n7428), .Y(n7429));
  OAI22X1 g04247(.A0(n7167), .A1(n7202), .B0(n4359), .B1(n7170), .Y(n7430));
  OAI22X1 g04248(.A0(n7182), .A1(n4472), .B0(n7204), .B1(n7169), .Y(n7431));
  OAI22X1 g04249(.A0(n7159), .A1(n7198), .B0(n4125), .B1(n7163), .Y(n7432));
  OAI22X1 g04250(.A0(n7166), .A1(n4247), .B0(n7200), .B1(n7162), .Y(n7433));
  NOR4X1  g04251(.A(n7432), .B(n7431), .C(n7430), .D(n7433), .Y(n7434));
  NAND2X1 g04252(.A(n7434), .B(n7429), .Y(n7435));
  NAND3X1 g04253(.A(n7435), .B(n7105), .C(n3666), .Y(n7436));
  NAND2X1 g04254(.A(P3_EAX_REG_16__SCAN_IN), .B(P3_EAX_REG_15__SCAN_IN), .Y(n7437));
  NOR4X1  g04255(.A(n7320), .B(n7052), .C(n7049), .D(n7437), .Y(n7438));
  XOR2X1  g04256(.A(n7438), .B(P3_EAX_REG_17__SCAN_IN), .Y(n7439));
  AOI22X1 g04257(.A0(n7111), .A1(n7439), .B0(n7107), .B1(P3_EAX_REG_17__SCAN_IN), .Y(n7440));
  AOI22X1 g04258(.A0(n7421), .A1(BUF2_REG_17__SCAN_IN), .B0(BUF2_REG_1__SCAN_IN), .B1(n7422), .Y(n7441));
  NAND3X1 g04259(.A(n7441), .B(n7440), .C(n7436), .Y(P3_U2718));
  OAI22X1 g04260(.A0(n7183), .A1(n7237), .B0(n4577), .B1(n7188), .Y(n7443));
  OAI22X1 g04261(.A0(n7174), .A1(n7240), .B0(n7239), .B1(n7187), .Y(n7444));
  OAI22X1 g04262(.A0(n3551), .A1(n3554), .B0(n7233), .B1(n7179), .Y(n7445));
  OAI22X1 g04263(.A0(n7158), .A1(n3549), .B0(n7235), .B1(n7178), .Y(n7446));
  NOR4X1  g04264(.A(n7445), .B(n7444), .C(n7443), .D(n7446), .Y(n7447));
  OAI22X1 g04265(.A0(n7167), .A1(n7229), .B0(n4353), .B1(n7170), .Y(n7448));
  OAI22X1 g04266(.A0(n7182), .A1(n4466), .B0(n3553), .B1(n7169), .Y(n7449));
  OAI22X1 g04267(.A0(n7159), .A1(n7225), .B0(n4117), .B1(n7163), .Y(n7450));
  OAI22X1 g04268(.A0(n7166), .A1(n4241), .B0(n7227), .B1(n7162), .Y(n7451));
  NOR4X1  g04269(.A(n7450), .B(n7449), .C(n7448), .D(n7451), .Y(n7452));
  NAND2X1 g04270(.A(n7452), .B(n7447), .Y(n7453));
  NAND3X1 g04271(.A(n7453), .B(n7105), .C(n3666), .Y(n7454));
  NAND2X1 g04272(.A(n7438), .B(P3_EAX_REG_17__SCAN_IN), .Y(n7455));
  XOR2X1  g04273(.A(n7455), .B(n7065), .Y(n7456));
  AOI22X1 g04274(.A0(n7111), .A1(n7456), .B0(n7107), .B1(P3_EAX_REG_18__SCAN_IN), .Y(n7457));
  AOI22X1 g04275(.A0(n7421), .A1(BUF2_REG_18__SCAN_IN), .B0(BUF2_REG_2__SCAN_IN), .B1(n7422), .Y(n7458));
  NAND3X1 g04276(.A(n7458), .B(n7457), .C(n7454), .Y(P3_U2717));
  OAI22X1 g04277(.A0(n7183), .A1(n7262), .B0(n4571), .B1(n7188), .Y(n7460));
  OAI22X1 g04278(.A0(n7174), .A1(n7265), .B0(n7264), .B1(n7187), .Y(n7461));
  OAI22X1 g04279(.A0(n3551), .A1(n3604), .B0(n7258), .B1(n7179), .Y(n7462));
  OAI22X1 g04280(.A0(n7158), .A1(n3601), .B0(n7260), .B1(n7178), .Y(n7463));
  NOR4X1  g04281(.A(n7462), .B(n7461), .C(n7460), .D(n7463), .Y(n7464));
  OAI22X1 g04282(.A0(n7167), .A1(n7254), .B0(n4347), .B1(n7170), .Y(n7465));
  OAI22X1 g04283(.A0(n7182), .A1(n4460), .B0(n3603), .B1(n7169), .Y(n7466));
  OAI22X1 g04284(.A0(n7159), .A1(n7250), .B0(n4109), .B1(n7163), .Y(n7467));
  OAI22X1 g04285(.A0(n7166), .A1(n4235), .B0(n7252), .B1(n7162), .Y(n7468));
  NOR4X1  g04286(.A(n7467), .B(n7466), .C(n7465), .D(n7468), .Y(n7469));
  NAND2X1 g04287(.A(n7469), .B(n7464), .Y(n7470));
  NAND3X1 g04288(.A(n7470), .B(n7105), .C(n3666), .Y(n7471));
  NAND3X1 g04289(.A(n7438), .B(P3_EAX_REG_18__SCAN_IN), .C(P3_EAX_REG_17__SCAN_IN), .Y(n7472));
  XOR2X1  g04290(.A(n7472), .B(n7068), .Y(n7473));
  AOI22X1 g04291(.A0(n7111), .A1(n7473), .B0(n7107), .B1(P3_EAX_REG_19__SCAN_IN), .Y(n7474));
  AOI22X1 g04292(.A0(n7421), .A1(BUF2_REG_19__SCAN_IN), .B0(BUF2_REG_3__SCAN_IN), .B1(n7422), .Y(n7475));
  NAND3X1 g04293(.A(n7475), .B(n7474), .C(n7471), .Y(P3_U2716));
  OAI22X1 g04294(.A0(n7183), .A1(n7287), .B0(n4565), .B1(n7188), .Y(n7477));
  OAI22X1 g04295(.A0(n7174), .A1(n7290), .B0(n7289), .B1(n7187), .Y(n7478));
  OAI22X1 g04296(.A0(n3551), .A1(n3622), .B0(n7283), .B1(n7179), .Y(n7479));
  OAI22X1 g04297(.A0(n7158), .A1(n3619), .B0(n7285), .B1(n7178), .Y(n7480));
  NOR4X1  g04298(.A(n7479), .B(n7478), .C(n7477), .D(n7480), .Y(n7481));
  OAI22X1 g04299(.A0(n7167), .A1(n7279), .B0(n4341), .B1(n7170), .Y(n7482));
  OAI22X1 g04300(.A0(n7182), .A1(n4454), .B0(n3621), .B1(n7169), .Y(n7483));
  OAI22X1 g04301(.A0(n7159), .A1(n7275), .B0(n4101), .B1(n7163), .Y(n7484));
  OAI22X1 g04302(.A0(n7166), .A1(n4229), .B0(n7277), .B1(n7162), .Y(n7485));
  NOR4X1  g04303(.A(n7484), .B(n7483), .C(n7482), .D(n7485), .Y(n7486));
  NAND2X1 g04304(.A(n7486), .B(n7481), .Y(n7487));
  NAND3X1 g04305(.A(n7487), .B(n7105), .C(n3666), .Y(n7488));
  NAND4X1 g04306(.A(P3_EAX_REG_19__SCAN_IN), .B(P3_EAX_REG_18__SCAN_IN), .C(P3_EAX_REG_17__SCAN_IN), .D(n7438), .Y(n7489));
  XOR2X1  g04307(.A(n7489), .B(n7071), .Y(n7490));
  AOI22X1 g04308(.A0(n7111), .A1(n7490), .B0(n7107), .B1(P3_EAX_REG_20__SCAN_IN), .Y(n7491));
  AOI22X1 g04309(.A0(n7421), .A1(BUF2_REG_20__SCAN_IN), .B0(BUF2_REG_4__SCAN_IN), .B1(n7422), .Y(n7492));
  NAND3X1 g04310(.A(n7492), .B(n7491), .C(n7488), .Y(P3_U2715));
  OAI22X1 g04311(.A0(n7183), .A1(n7312), .B0(n4559), .B1(n7188), .Y(n7494));
  OAI22X1 g04312(.A0(n7174), .A1(n7315), .B0(n7314), .B1(n7187), .Y(n7495));
  OAI22X1 g04313(.A0(n3551), .A1(n3638), .B0(n7308), .B1(n7179), .Y(n7496));
  OAI22X1 g04314(.A0(n7158), .A1(n3635), .B0(n7310), .B1(n7178), .Y(n7497));
  NOR4X1  g04315(.A(n7496), .B(n7495), .C(n7494), .D(n7497), .Y(n7498));
  OAI22X1 g04316(.A0(n7167), .A1(n7304), .B0(n4335), .B1(n7170), .Y(n7499));
  OAI22X1 g04317(.A0(n7182), .A1(n4448), .B0(n3637), .B1(n7169), .Y(n7500));
  OAI22X1 g04318(.A0(n7159), .A1(n7300), .B0(n4093), .B1(n7163), .Y(n7501));
  OAI22X1 g04319(.A0(n7166), .A1(n4223), .B0(n7302), .B1(n7162), .Y(n7502));
  NOR4X1  g04320(.A(n7501), .B(n7500), .C(n7499), .D(n7502), .Y(n7503));
  NAND2X1 g04321(.A(n7503), .B(n7498), .Y(n7504));
  NAND3X1 g04322(.A(n7504), .B(n7105), .C(n3666), .Y(n7505));
  NOR3X1  g04323(.A(n7472), .B(n7071), .C(n7068), .Y(n7506));
  XOR2X1  g04324(.A(n7506), .B(P3_EAX_REG_21__SCAN_IN), .Y(n7507));
  AOI22X1 g04325(.A0(n7111), .A1(n7507), .B0(n7107), .B1(P3_EAX_REG_21__SCAN_IN), .Y(n7508));
  AOI22X1 g04326(.A0(n7421), .A1(BUF2_REG_21__SCAN_IN), .B0(BUF2_REG_5__SCAN_IN), .B1(n7422), .Y(n7509));
  NAND3X1 g04327(.A(n7509), .B(n7508), .C(n7505), .Y(P3_U2714));
  OAI22X1 g04328(.A0(n7183), .A1(n7337), .B0(n4553), .B1(n7188), .Y(n7511));
  OAI22X1 g04329(.A0(n7174), .A1(n7340), .B0(n7339), .B1(n7187), .Y(n7512));
  OAI22X1 g04330(.A0(n3551), .A1(n3654), .B0(n7333), .B1(n7179), .Y(n7513));
  OAI22X1 g04331(.A0(n7158), .A1(n3651), .B0(n7335), .B1(n7178), .Y(n7514));
  NOR4X1  g04332(.A(n7513), .B(n7512), .C(n7511), .D(n7514), .Y(n7515));
  OAI22X1 g04333(.A0(n7167), .A1(n7329), .B0(n4329), .B1(n7170), .Y(n7516));
  OAI22X1 g04334(.A0(n7182), .A1(n4442), .B0(n3653), .B1(n7169), .Y(n7517));
  OAI22X1 g04335(.A0(n7159), .A1(n7325), .B0(n4085), .B1(n7163), .Y(n7518));
  OAI22X1 g04336(.A0(n7166), .A1(n4217), .B0(n7327), .B1(n7162), .Y(n7519));
  NOR4X1  g04337(.A(n7518), .B(n7517), .C(n7516), .D(n7519), .Y(n7520));
  NAND2X1 g04338(.A(n7520), .B(n7515), .Y(n7521));
  NAND3X1 g04339(.A(n7521), .B(n7105), .C(n3666), .Y(n7522));
  NOR4X1  g04340(.A(n7074), .B(n7071), .C(n7068), .D(n7472), .Y(n7523));
  XOR2X1  g04341(.A(n7523), .B(P3_EAX_REG_22__SCAN_IN), .Y(n7524));
  AOI22X1 g04342(.A0(n7111), .A1(n7524), .B0(n7107), .B1(P3_EAX_REG_22__SCAN_IN), .Y(n7525));
  AOI22X1 g04343(.A0(n7421), .A1(BUF2_REG_22__SCAN_IN), .B0(BUF2_REG_6__SCAN_IN), .B1(n7422), .Y(n7526));
  NAND3X1 g04344(.A(n7526), .B(n7525), .C(n7522), .Y(P3_U2713));
  AOI22X1 g04345(.A0(n3571), .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B0(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3572), .Y(n7530));
  AOI22X1 g04346(.A0(n3575), .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B0(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3568), .Y(n7533));
  NAND2X1 g04347(.A(n7533), .B(n7530), .Y(n7534));
  AOI22X1 g04348(.A0(n3563), .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B0(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3578), .Y(n7537));
  AOI22X1 g04349(.A0(n3569), .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B0(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3577), .Y(n7540));
  NAND2X1 g04350(.A(n7540), .B(n7537), .Y(n7541));
  AOI22X1 g04351(.A0(n3565), .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B0(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3574), .Y(n7544));
  AOI22X1 g04352(.A0(n3562), .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B0(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3555), .Y(n7547));
  AOI22X1 g04353(.A0(n3566), .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B0(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3550), .Y(n7550));
  AOI22X1 g04354(.A0(n3560), .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B0(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3557), .Y(n7553));
  NAND4X1 g04355(.A(n7550), .B(n7547), .C(n7544), .D(n7553), .Y(n7554));
  NOR3X1  g04356(.A(n7554), .B(n7541), .C(n7534), .Y(n7555));
  AOI22X1 g04357(.A0(n3575), .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B0(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3555), .Y(n7556));
  AOI22X1 g04358(.A0(n3562), .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B0(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3574), .Y(n7557));
  AOI22X1 g04359(.A0(n3550), .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B0(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3577), .Y(n7558));
  AOI22X1 g04360(.A0(n3569), .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B0(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3578), .Y(n7559));
  NAND4X1 g04361(.A(n7558), .B(n7557), .C(n7556), .D(n7559), .Y(n7560));
  AOI22X1 g04362(.A0(n3560), .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B0(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3571), .Y(n7561));
  AOI22X1 g04363(.A0(n3568), .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B0(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3572), .Y(n7562));
  AOI22X1 g04364(.A0(n3563), .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B0(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3565), .Y(n7563));
  AOI22X1 g04365(.A0(n3557), .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B0(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3566), .Y(n7564));
  NAND4X1 g04366(.A(n7563), .B(n7562), .C(n7561), .D(n7564), .Y(n7565));
  NOR2X1  g04367(.A(n7565), .B(n7560), .Y(n7566));
  XOR2X1  g04368(.A(n7566), .B(n7555), .Y(n7567));
  NAND3X1 g04369(.A(n7567), .B(n7105), .C(n3666), .Y(n7568));
  NAND3X1 g04370(.A(n7506), .B(P3_EAX_REG_22__SCAN_IN), .C(P3_EAX_REG_21__SCAN_IN), .Y(n7569));
  XOR2X1  g04371(.A(n7569), .B(n7080), .Y(n7570));
  AOI22X1 g04372(.A0(n7111), .A1(n7570), .B0(n7107), .B1(P3_EAX_REG_23__SCAN_IN), .Y(n7571));
  AOI22X1 g04373(.A0(n7421), .A1(BUF2_REG_23__SCAN_IN), .B0(BUF2_REG_7__SCAN_IN), .B1(n7422), .Y(n7572));
  NAND3X1 g04374(.A(n7572), .B(n7571), .C(n7568), .Y(P3_U2712));
  NOR2X1  g04375(.A(n7566), .B(n7555), .Y(n7574));
  AOI22X1 g04376(.A0(n3571), .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B0(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3572), .Y(n7575));
  AOI22X1 g04377(.A0(n3575), .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B0(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3568), .Y(n7576));
  NAND2X1 g04378(.A(n7576), .B(n7575), .Y(n7577));
  AOI22X1 g04379(.A0(n3563), .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B0(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3578), .Y(n7578));
  INVX1   g04380(.A(n7578), .Y(n7579));
  AOI22X1 g04381(.A0(n3569), .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B0(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3577), .Y(n7580));
  INVX1   g04382(.A(n7580), .Y(n7581));
  AOI22X1 g04383(.A0(n3565), .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B0(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3574), .Y(n7582));
  AOI22X1 g04384(.A0(n3562), .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B0(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3555), .Y(n7583));
  AOI22X1 g04385(.A0(n3566), .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B0(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3550), .Y(n7584));
  AOI22X1 g04386(.A0(n3560), .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B0(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3557), .Y(n7585));
  NAND4X1 g04387(.A(n7584), .B(n7583), .C(n7582), .D(n7585), .Y(n7586));
  NOR4X1  g04388(.A(n7581), .B(n7579), .C(n7577), .D(n7586), .Y(n7587));
  INVX1   g04389(.A(n7587), .Y(n7588));
  XOR2X1  g04390(.A(n7588), .B(n7574), .Y(n7589));
  NAND3X1 g04391(.A(n7589), .B(n7105), .C(n3666), .Y(n7590));
  NAND4X1 g04392(.A(P3_EAX_REG_23__SCAN_IN), .B(P3_EAX_REG_22__SCAN_IN), .C(P3_EAX_REG_21__SCAN_IN), .D(n7506), .Y(n7591));
  XOR2X1  g04393(.A(n7591), .B(n7083), .Y(n7592));
  AOI22X1 g04394(.A0(n7111), .A1(n7592), .B0(n7107), .B1(P3_EAX_REG_24__SCAN_IN), .Y(n7593));
  AOI22X1 g04395(.A0(n7421), .A1(BUF2_REG_24__SCAN_IN), .B0(BUF2_REG_8__SCAN_IN), .B1(n7422), .Y(n7594));
  NAND3X1 g04396(.A(n7594), .B(n7593), .C(n7590), .Y(P3_U2711));
  NOR3X1  g04397(.A(n7587), .B(n7566), .C(n7555), .Y(n7596));
  AOI22X1 g04398(.A0(n3571), .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B0(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3572), .Y(n7597));
  AOI22X1 g04399(.A0(n3575), .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B0(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3568), .Y(n7598));
  NAND2X1 g04400(.A(n7598), .B(n7597), .Y(n7599));
  AOI22X1 g04401(.A0(n3563), .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B0(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3578), .Y(n7600));
  INVX1   g04402(.A(n7600), .Y(n7601));
  AOI22X1 g04403(.A0(n3569), .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B0(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3577), .Y(n7602));
  INVX1   g04404(.A(n7602), .Y(n7603));
  AOI22X1 g04405(.A0(n3565), .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B0(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3574), .Y(n7604));
  AOI22X1 g04406(.A0(n3562), .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B0(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3555), .Y(n7605));
  AOI22X1 g04407(.A0(n3566), .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B0(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3550), .Y(n7606));
  AOI22X1 g04408(.A0(n3560), .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B0(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3557), .Y(n7607));
  NAND4X1 g04409(.A(n7606), .B(n7605), .C(n7604), .D(n7607), .Y(n7608));
  NOR4X1  g04410(.A(n7603), .B(n7601), .C(n7599), .D(n7608), .Y(n7609));
  INVX1   g04411(.A(n7609), .Y(n7610));
  XOR2X1  g04412(.A(n7610), .B(n7596), .Y(n7611));
  NAND3X1 g04413(.A(n7611), .B(n7105), .C(n3666), .Y(n7612));
  NOR3X1  g04414(.A(n7569), .B(n7083), .C(n7080), .Y(n7613));
  XOR2X1  g04415(.A(n7613), .B(P3_EAX_REG_25__SCAN_IN), .Y(n7614));
  AOI22X1 g04416(.A0(n7111), .A1(n7614), .B0(n7107), .B1(P3_EAX_REG_25__SCAN_IN), .Y(n7615));
  AOI22X1 g04417(.A0(n7421), .A1(BUF2_REG_25__SCAN_IN), .B0(BUF2_REG_9__SCAN_IN), .B1(n7422), .Y(n7616));
  NAND3X1 g04418(.A(n7616), .B(n7615), .C(n7612), .Y(P3_U2710));
  NOR4X1  g04419(.A(n7587), .B(n7566), .C(n7555), .D(n7609), .Y(n7618));
  AOI22X1 g04420(.A0(n3571), .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B0(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3572), .Y(n7619));
  AOI22X1 g04421(.A0(n3575), .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B0(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3568), .Y(n7620));
  NAND2X1 g04422(.A(n7620), .B(n7619), .Y(n7621));
  AOI22X1 g04423(.A0(n3563), .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B0(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3578), .Y(n7622));
  AOI22X1 g04424(.A0(n3569), .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B0(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3577), .Y(n7623));
  NAND2X1 g04425(.A(n7623), .B(n7622), .Y(n7624));
  AOI22X1 g04426(.A0(n3565), .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B0(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3574), .Y(n7625));
  AOI22X1 g04427(.A0(n3562), .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B0(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3555), .Y(n7626));
  AOI22X1 g04428(.A0(n3566), .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B0(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3550), .Y(n7627));
  AOI22X1 g04429(.A0(n3560), .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B0(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3557), .Y(n7628));
  NAND4X1 g04430(.A(n7627), .B(n7626), .C(n7625), .D(n7628), .Y(n7629));
  NOR3X1  g04431(.A(n7629), .B(n7624), .C(n7621), .Y(n7630));
  INVX1   g04432(.A(n7630), .Y(n7631));
  XOR2X1  g04433(.A(n7631), .B(n7618), .Y(n7632));
  NAND3X1 g04434(.A(n7632), .B(n7105), .C(n3666), .Y(n7633));
  NOR4X1  g04435(.A(n7086), .B(n7083), .C(n7080), .D(n7569), .Y(n7634));
  XOR2X1  g04436(.A(n7634), .B(P3_EAX_REG_26__SCAN_IN), .Y(n7635));
  AOI22X1 g04437(.A0(n7111), .A1(n7635), .B0(n7107), .B1(P3_EAX_REG_26__SCAN_IN), .Y(n7636));
  AOI22X1 g04438(.A0(n7421), .A1(BUF2_REG_26__SCAN_IN), .B0(BUF2_REG_10__SCAN_IN), .B1(n7422), .Y(n7637));
  NAND3X1 g04439(.A(n7637), .B(n7636), .C(n7633), .Y(P3_U2709));
  NAND2X1 g04440(.A(n7631), .B(n7618), .Y(n7639));
  AOI22X1 g04441(.A0(n3571), .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B0(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3572), .Y(n7640));
  AOI22X1 g04442(.A0(n3575), .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B0(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3568), .Y(n7641));
  NAND2X1 g04443(.A(n7641), .B(n7640), .Y(n7642));
  AOI22X1 g04444(.A0(n3563), .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B0(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3578), .Y(n7643));
  INVX1   g04445(.A(n7643), .Y(n7644));
  AOI22X1 g04446(.A0(n3569), .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B0(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3577), .Y(n7645));
  INVX1   g04447(.A(n7645), .Y(n7646));
  AOI22X1 g04448(.A0(n3565), .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B0(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3574), .Y(n7647));
  AOI22X1 g04449(.A0(n3562), .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B0(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3555), .Y(n7648));
  AOI22X1 g04450(.A0(n3566), .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B0(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3550), .Y(n7649));
  AOI22X1 g04451(.A0(n3560), .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B0(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3557), .Y(n7650));
  NAND4X1 g04452(.A(n7649), .B(n7648), .C(n7647), .D(n7650), .Y(n7651));
  NOR4X1  g04453(.A(n7646), .B(n7644), .C(n7642), .D(n7651), .Y(n7652));
  XOR2X1  g04454(.A(n7652), .B(n7639), .Y(n7653));
  NAND3X1 g04455(.A(n7653), .B(n7105), .C(n3666), .Y(n7654));
  NAND3X1 g04456(.A(n7613), .B(P3_EAX_REG_26__SCAN_IN), .C(P3_EAX_REG_25__SCAN_IN), .Y(n7655));
  XOR2X1  g04457(.A(n7655), .B(n7092), .Y(n7656));
  AOI22X1 g04458(.A0(n7111), .A1(n7656), .B0(n7107), .B1(P3_EAX_REG_27__SCAN_IN), .Y(n7657));
  AOI22X1 g04459(.A0(n7421), .A1(BUF2_REG_27__SCAN_IN), .B0(BUF2_REG_11__SCAN_IN), .B1(n7422), .Y(n7658));
  NAND3X1 g04460(.A(n7658), .B(n7657), .C(n7654), .Y(P3_U2708));
  INVX1   g04461(.A(n7652), .Y(n7660));
  NAND3X1 g04462(.A(n7660), .B(n7631), .C(n7618), .Y(n7661));
  AOI22X1 g04463(.A0(n3571), .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B0(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3572), .Y(n7662));
  AOI22X1 g04464(.A0(n3575), .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B0(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3568), .Y(n7663));
  NAND2X1 g04465(.A(n7663), .B(n7662), .Y(n7664));
  OAI22X1 g04466(.A0(n7159), .A1(n3635), .B0(n7308), .B1(n7178), .Y(n7667));
  OAI22X1 g04467(.A0(n7158), .A1(n7310), .B0(n3638), .B1(n7179), .Y(n7670));
  AOI22X1 g04468(.A0(n3565), .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B0(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3574), .Y(n7671));
  AOI22X1 g04469(.A0(n3562), .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B0(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3555), .Y(n7672));
  AOI22X1 g04470(.A0(n3566), .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B0(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3550), .Y(n7673));
  AOI22X1 g04471(.A0(n3560), .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B0(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3557), .Y(n7674));
  NAND4X1 g04472(.A(n7673), .B(n7672), .C(n7671), .D(n7674), .Y(n7675));
  NOR4X1  g04473(.A(n7670), .B(n7667), .C(n7664), .D(n7675), .Y(n7676));
  XOR2X1  g04474(.A(n7676), .B(n7661), .Y(n7677));
  NAND3X1 g04475(.A(n7677), .B(n7105), .C(n3666), .Y(n7678));
  NAND4X1 g04476(.A(P3_EAX_REG_27__SCAN_IN), .B(P3_EAX_REG_26__SCAN_IN), .C(P3_EAX_REG_25__SCAN_IN), .D(n7613), .Y(n7679));
  XOR2X1  g04477(.A(n7679), .B(n7095), .Y(n7680));
  AOI22X1 g04478(.A0(n7111), .A1(n7680), .B0(n7107), .B1(P3_EAX_REG_28__SCAN_IN), .Y(n7681));
  AOI22X1 g04479(.A0(n7421), .A1(BUF2_REG_28__SCAN_IN), .B0(BUF2_REG_12__SCAN_IN), .B1(n7422), .Y(n7682));
  NAND3X1 g04480(.A(n7682), .B(n7681), .C(n7678), .Y(P3_U2707));
  NOR2X1  g04481(.A(n7676), .B(n7661), .Y(n7684));
  AOI22X1 g04482(.A0(n3571), .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B0(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3572), .Y(n7685));
  AOI22X1 g04483(.A0(n3575), .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B0(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3568), .Y(n7686));
  OAI22X1 g04484(.A0(n7159), .A1(n3651), .B0(n7333), .B1(n7178), .Y(n7687));
  OAI22X1 g04485(.A0(n7158), .A1(n7335), .B0(n3654), .B1(n7179), .Y(n7688));
  AOI22X1 g04486(.A0(n3565), .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B0(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3574), .Y(n7689));
  AOI22X1 g04487(.A0(n3562), .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B0(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3555), .Y(n7690));
  AOI22X1 g04488(.A0(n3566), .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B0(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3550), .Y(n7691));
  AOI22X1 g04489(.A0(n3560), .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B0(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3557), .Y(n7692));
  NAND4X1 g04490(.A(n7691), .B(n7690), .C(n7689), .D(n7692), .Y(n7693));
  NOR3X1  g04491(.A(n7693), .B(n7688), .C(n7687), .Y(n7694));
  NAND3X1 g04492(.A(n7694), .B(n7686), .C(n7685), .Y(n7695));
  XOR2X1  g04493(.A(n7695), .B(n7684), .Y(n7696));
  NAND3X1 g04494(.A(n7696), .B(n7105), .C(n3666), .Y(n7697));
  NAND2X1 g04495(.A(P3_EAX_REG_28__SCAN_IN), .B(P3_EAX_REG_27__SCAN_IN), .Y(n7698));
  NOR2X1  g04496(.A(n7698), .B(n7655), .Y(n7699));
  XOR2X1  g04497(.A(n7699), .B(P3_EAX_REG_29__SCAN_IN), .Y(n7700));
  AOI22X1 g04498(.A0(n7111), .A1(n7700), .B0(n7107), .B1(P3_EAX_REG_29__SCAN_IN), .Y(n7701));
  AOI22X1 g04499(.A0(n7421), .A1(BUF2_REG_29__SCAN_IN), .B0(BUF2_REG_13__SCAN_IN), .B1(n7422), .Y(n7702));
  NAND3X1 g04500(.A(n7702), .B(n7701), .C(n7697), .Y(P3_U2706));
  NAND2X1 g04501(.A(n7695), .B(n7684), .Y(n7704));
  AOI22X1 g04502(.A0(n3571), .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B0(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3572), .Y(n7705));
  AOI22X1 g04503(.A0(n3575), .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B0(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3568), .Y(n7706));
  NAND2X1 g04504(.A(n7706), .B(n7705), .Y(n7707));
  OAI22X1 g04505(.A0(n7159), .A1(n3585), .B0(n7358), .B1(n7178), .Y(n7708));
  OAI22X1 g04506(.A0(n7158), .A1(n7360), .B0(n3588), .B1(n7179), .Y(n7709));
  AOI22X1 g04507(.A0(n3565), .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B0(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3574), .Y(n7710));
  AOI22X1 g04508(.A0(n3562), .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B0(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3555), .Y(n7711));
  AOI22X1 g04509(.A0(n3566), .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B0(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3550), .Y(n7712));
  AOI22X1 g04510(.A0(n3560), .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B0(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3557), .Y(n7713));
  NAND4X1 g04511(.A(n7712), .B(n7711), .C(n7710), .D(n7713), .Y(n7714));
  NOR4X1  g04512(.A(n7709), .B(n7708), .C(n7707), .D(n7714), .Y(n7715));
  XOR2X1  g04513(.A(n7715), .B(n7704), .Y(n7716));
  NAND3X1 g04514(.A(n7716), .B(n7105), .C(n3666), .Y(n7717));
  NOR3X1  g04515(.A(n7698), .B(n7655), .C(n7098), .Y(n7718));
  XOR2X1  g04516(.A(n7718), .B(P3_EAX_REG_30__SCAN_IN), .Y(n7719));
  AOI22X1 g04517(.A0(n7111), .A1(n7719), .B0(n7107), .B1(P3_EAX_REG_30__SCAN_IN), .Y(n7720));
  AOI22X1 g04518(.A0(n7421), .A1(BUF2_REG_30__SCAN_IN), .B0(BUF2_REG_14__SCAN_IN), .B1(n7422), .Y(n7721));
  NAND3X1 g04519(.A(n7721), .B(n7720), .C(n7717), .Y(P3_U2705));
  NAND4X1 g04520(.A(n3715), .B(n3774), .C(BUF2_REG_31__SCAN_IN), .D(n7105), .Y(n7723));
  NOR4X1  g04521(.A(n7655), .B(n7101), .C(n7098), .D(n7698), .Y(n7724));
  XOR2X1  g04522(.A(n7724), .B(P3_EAX_REG_31__SCAN_IN), .Y(n7725));
  AOI22X1 g04523(.A0(n7111), .A1(n7725), .B0(n7107), .B1(P3_EAX_REG_31__SCAN_IN), .Y(n7726));
  NAND2X1 g04524(.A(n7726), .B(n7723), .Y(P3_U2704));
  AOI21X1 g04525(.A0(n5043), .A1(n3746), .B0(n4905), .Y(n7728));
  INVX1   g04526(.A(n7728), .Y(n7729));
  NOR2X1  g04527(.A(n7729), .B(n3774), .Y(n7730));
  INVX1   g04528(.A(n7730), .Y(n7731));
  NOR2X1  g04529(.A(n7729), .B(n3600), .Y(n7732));
  AOI22X1 g04530(.A0(n7729), .A1(P3_EBX_REG_0__SCAN_IN), .B0(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(n7732), .Y(n7733));
  OAI21X1 g04531(.A0(n7731), .A1(P3_EBX_REG_0__SCAN_IN), .B0(n7733), .Y(P3_U2703));
  INVX1   g04532(.A(P3_EBX_REG_0__SCAN_IN), .Y(n7735));
  XOR2X1  g04533(.A(P3_EBX_REG_1__SCAN_IN), .B(n7735), .Y(n7736));
  AOI22X1 g04534(.A0(n7729), .A1(P3_EBX_REG_1__SCAN_IN), .B0(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(n7732), .Y(n7737));
  OAI21X1 g04535(.A0(n7736), .A1(n7731), .B0(n7737), .Y(P3_U2702));
  NAND2X1 g04536(.A(P3_EBX_REG_1__SCAN_IN), .B(P3_EBX_REG_0__SCAN_IN), .Y(n7739));
  XOR2X1  g04537(.A(n7739), .B(P3_EBX_REG_2__SCAN_IN), .Y(n7740));
  AOI22X1 g04538(.A0(n7729), .A1(P3_EBX_REG_2__SCAN_IN), .B0(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(n7732), .Y(n7741));
  OAI21X1 g04539(.A0(n7740), .A1(n7731), .B0(n7741), .Y(P3_U2701));
  INVX1   g04540(.A(P3_EBX_REG_3__SCAN_IN), .Y(n7743));
  INVX1   g04541(.A(P3_EBX_REG_2__SCAN_IN), .Y(n7744));
  NOR2X1  g04542(.A(n7739), .B(n7744), .Y(n7745));
  XOR2X1  g04543(.A(n7745), .B(n7743), .Y(n7746));
  AOI22X1 g04544(.A0(n7729), .A1(P3_EBX_REG_3__SCAN_IN), .B0(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(n7732), .Y(n7747));
  OAI21X1 g04545(.A0(n7746), .A1(n7731), .B0(n7747), .Y(P3_U2700));
  NAND4X1 g04546(.A(P3_EBX_REG_2__SCAN_IN), .B(P3_EBX_REG_1__SCAN_IN), .C(P3_EBX_REG_0__SCAN_IN), .D(P3_EBX_REG_3__SCAN_IN), .Y(n7749));
  XOR2X1  g04547(.A(n7749), .B(P3_EBX_REG_4__SCAN_IN), .Y(n7750));
  AOI22X1 g04548(.A0(n7729), .A1(P3_EBX_REG_4__SCAN_IN), .B0(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(n7732), .Y(n7751));
  OAI21X1 g04549(.A0(n7750), .A1(n7731), .B0(n7751), .Y(P3_U2699));
  INVX1   g04550(.A(P3_EBX_REG_5__SCAN_IN), .Y(n7753));
  INVX1   g04551(.A(P3_EBX_REG_4__SCAN_IN), .Y(n7754));
  NOR4X1  g04552(.A(n7754), .B(n7743), .C(n7744), .D(n7739), .Y(n7755));
  XOR2X1  g04553(.A(n7755), .B(n7753), .Y(n7756));
  AOI22X1 g04554(.A0(n7729), .A1(P3_EBX_REG_5__SCAN_IN), .B0(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(n7732), .Y(n7757));
  OAI21X1 g04555(.A0(n7756), .A1(n7731), .B0(n7757), .Y(P3_U2698));
  NAND2X1 g04556(.A(n7755), .B(P3_EBX_REG_5__SCAN_IN), .Y(n7759));
  XOR2X1  g04557(.A(n7759), .B(P3_EBX_REG_6__SCAN_IN), .Y(n7760));
  AOI22X1 g04558(.A0(n7729), .A1(P3_EBX_REG_6__SCAN_IN), .B0(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(n7732), .Y(n7761));
  OAI21X1 g04559(.A0(n7760), .A1(n7731), .B0(n7761), .Y(P3_U2697));
  NAND2X1 g04560(.A(P3_EBX_REG_4__SCAN_IN), .B(P3_EBX_REG_3__SCAN_IN), .Y(n7763));
  NAND2X1 g04561(.A(P3_EBX_REG_6__SCAN_IN), .B(P3_EBX_REG_5__SCAN_IN), .Y(n7764));
  NOR4X1  g04562(.A(n7763), .B(n7739), .C(n7744), .D(n7764), .Y(n7765));
  XOR2X1  g04563(.A(n7765), .B(P3_EBX_REG_7__SCAN_IN), .Y(n7766));
  NAND3X1 g04564(.A(n7766), .B(n7728), .C(n3600), .Y(n7767));
  AOI22X1 g04565(.A0(n7729), .A1(P3_EBX_REG_7__SCAN_IN), .B0(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(n7732), .Y(n7768));
  NAND2X1 g04566(.A(n7768), .B(n7767), .Y(P3_U2696));
  NAND2X1 g04567(.A(n7765), .B(P3_EBX_REG_7__SCAN_IN), .Y(n7770));
  XOR2X1  g04568(.A(n7770), .B(P3_EBX_REG_8__SCAN_IN), .Y(n7771));
  AOI22X1 g04569(.A0(n7729), .A1(P3_EBX_REG_8__SCAN_IN), .B0(n7191), .B1(n7732), .Y(n7772));
  OAI21X1 g04570(.A0(n7771), .A1(n7731), .B0(n7772), .Y(P3_U2695));
  NAND3X1 g04571(.A(n7765), .B(P3_EBX_REG_8__SCAN_IN), .C(P3_EBX_REG_7__SCAN_IN), .Y(n7774));
  XOR2X1  g04572(.A(n7774), .B(P3_EBX_REG_9__SCAN_IN), .Y(n7775));
  AOI22X1 g04573(.A0(n7729), .A1(P3_EBX_REG_9__SCAN_IN), .B0(n7218), .B1(n7732), .Y(n7776));
  OAI21X1 g04574(.A0(n7775), .A1(n7731), .B0(n7776), .Y(P3_U2694));
  NAND3X1 g04575(.A(n7728), .B(n7243), .C(n3774), .Y(n7778));
  INVX1   g04576(.A(P3_EBX_REG_10__SCAN_IN), .Y(n7779));
  NAND4X1 g04577(.A(P3_EBX_REG_9__SCAN_IN), .B(P3_EBX_REG_8__SCAN_IN), .C(P3_EBX_REG_7__SCAN_IN), .D(n7765), .Y(n7780));
  XOR2X1  g04578(.A(n7780), .B(n7779), .Y(n7781));
  AOI22X1 g04579(.A0(n7730), .A1(n7781), .B0(n7729), .B1(P3_EBX_REG_10__SCAN_IN), .Y(n7782));
  NAND2X1 g04580(.A(n7782), .B(n7778), .Y(P3_U2693));
  NAND3X1 g04581(.A(n7728), .B(n7268), .C(n3774), .Y(n7784));
  INVX1   g04582(.A(P3_EBX_REG_9__SCAN_IN), .Y(n7785));
  NOR3X1  g04583(.A(n7774), .B(n7779), .C(n7785), .Y(n7786));
  XOR2X1  g04584(.A(n7786), .B(P3_EBX_REG_11__SCAN_IN), .Y(n7787));
  AOI22X1 g04585(.A0(n7730), .A1(n7787), .B0(n7729), .B1(P3_EBX_REG_11__SCAN_IN), .Y(n7788));
  NAND2X1 g04586(.A(n7788), .B(n7784), .Y(P3_U2692));
  NAND3X1 g04587(.A(n7728), .B(n7293), .C(n3774), .Y(n7790));
  INVX1   g04588(.A(P3_EBX_REG_11__SCAN_IN), .Y(n7791));
  NOR4X1  g04589(.A(n7791), .B(n7779), .C(n7785), .D(n7774), .Y(n7792));
  XOR2X1  g04590(.A(n7792), .B(P3_EBX_REG_12__SCAN_IN), .Y(n7793));
  AOI22X1 g04591(.A0(n7730), .A1(n7793), .B0(n7729), .B1(P3_EBX_REG_12__SCAN_IN), .Y(n7794));
  NAND2X1 g04592(.A(n7794), .B(n7790), .Y(P3_U2691));
  NAND3X1 g04593(.A(n7728), .B(n7318), .C(n3774), .Y(n7796));
  INVX1   g04594(.A(P3_EBX_REG_13__SCAN_IN), .Y(n7797));
  NAND3X1 g04595(.A(n7786), .B(P3_EBX_REG_12__SCAN_IN), .C(P3_EBX_REG_11__SCAN_IN), .Y(n7798));
  XOR2X1  g04596(.A(n7798), .B(n7797), .Y(n7799));
  AOI22X1 g04597(.A0(n7730), .A1(n7799), .B0(n7729), .B1(P3_EBX_REG_13__SCAN_IN), .Y(n7800));
  NAND2X1 g04598(.A(n7800), .B(n7796), .Y(P3_U2690));
  NAND3X1 g04599(.A(n7728), .B(n7343), .C(n3774), .Y(n7802));
  INVX1   g04600(.A(P3_EBX_REG_14__SCAN_IN), .Y(n7803));
  NAND4X1 g04601(.A(P3_EBX_REG_13__SCAN_IN), .B(P3_EBX_REG_12__SCAN_IN), .C(P3_EBX_REG_11__SCAN_IN), .D(n7786), .Y(n7804));
  XOR2X1  g04602(.A(n7804), .B(n7803), .Y(n7805));
  AOI22X1 g04603(.A0(n7730), .A1(n7805), .B0(n7729), .B1(P3_EBX_REG_14__SCAN_IN), .Y(n7806));
  NAND2X1 g04604(.A(n7806), .B(n7802), .Y(P3_U2689));
  NAND3X1 g04605(.A(n7728), .B(n7368), .C(n3774), .Y(n7808));
  NOR3X1  g04606(.A(n7798), .B(n7803), .C(n7797), .Y(n7809));
  XOR2X1  g04607(.A(n7809), .B(P3_EBX_REG_15__SCAN_IN), .Y(n7810));
  AOI22X1 g04608(.A0(n7730), .A1(n7810), .B0(n7729), .B1(P3_EBX_REG_15__SCAN_IN), .Y(n7811));
  NAND2X1 g04609(.A(n7811), .B(n7808), .Y(P3_U2688));
  NAND3X1 g04610(.A(n7728), .B(n7416), .C(n3774), .Y(n7813));
  INVX1   g04611(.A(P3_EBX_REG_15__SCAN_IN), .Y(n7814));
  NOR4X1  g04612(.A(n7814), .B(n7803), .C(n7797), .D(n7798), .Y(n7815));
  XOR2X1  g04613(.A(n7815), .B(P3_EBX_REG_16__SCAN_IN), .Y(n7816));
  AOI22X1 g04614(.A0(n7730), .A1(n7816), .B0(n7729), .B1(P3_EBX_REG_16__SCAN_IN), .Y(n7817));
  NAND2X1 g04615(.A(n7817), .B(n7813), .Y(P3_U2687));
  NAND3X1 g04616(.A(n7728), .B(n7435), .C(n3774), .Y(n7819));
  NAND2X1 g04617(.A(P3_EBX_REG_16__SCAN_IN), .B(P3_EBX_REG_15__SCAN_IN), .Y(n7820));
  NOR4X1  g04618(.A(n7798), .B(n7803), .C(n7797), .D(n7820), .Y(n7821));
  XOR2X1  g04619(.A(n7821), .B(P3_EBX_REG_17__SCAN_IN), .Y(n7822));
  AOI22X1 g04620(.A0(n7730), .A1(n7822), .B0(n7729), .B1(P3_EBX_REG_17__SCAN_IN), .Y(n7823));
  NAND2X1 g04621(.A(n7823), .B(n7819), .Y(P3_U2686));
  NAND3X1 g04622(.A(n7728), .B(n7453), .C(n3774), .Y(n7825));
  INVX1   g04623(.A(P3_EBX_REG_17__SCAN_IN), .Y(n7826));
  NAND2X1 g04624(.A(P3_EBX_REG_14__SCAN_IN), .B(P3_EBX_REG_13__SCAN_IN), .Y(n7827));
  NOR4X1  g04625(.A(n7827), .B(n7798), .C(n7826), .D(n7820), .Y(n7828));
  XOR2X1  g04626(.A(n7828), .B(P3_EBX_REG_18__SCAN_IN), .Y(n7829));
  AOI22X1 g04627(.A0(n7730), .A1(n7829), .B0(n7729), .B1(P3_EBX_REG_18__SCAN_IN), .Y(n7830));
  NAND2X1 g04628(.A(n7830), .B(n7825), .Y(P3_U2685));
  NAND3X1 g04629(.A(n7728), .B(n7470), .C(n3774), .Y(n7832));
  INVX1   g04630(.A(P3_EBX_REG_19__SCAN_IN), .Y(n7833));
  NAND3X1 g04631(.A(n7821), .B(P3_EBX_REG_18__SCAN_IN), .C(P3_EBX_REG_17__SCAN_IN), .Y(n7834));
  XOR2X1  g04632(.A(n7834), .B(n7833), .Y(n7835));
  AOI22X1 g04633(.A0(n7730), .A1(n7835), .B0(n7729), .B1(P3_EBX_REG_19__SCAN_IN), .Y(n7836));
  NAND2X1 g04634(.A(n7836), .B(n7832), .Y(P3_U2684));
  NAND3X1 g04635(.A(n7728), .B(n7487), .C(n3774), .Y(n7838));
  INVX1   g04636(.A(P3_EBX_REG_20__SCAN_IN), .Y(n7839));
  NAND4X1 g04637(.A(P3_EBX_REG_19__SCAN_IN), .B(P3_EBX_REG_18__SCAN_IN), .C(P3_EBX_REG_17__SCAN_IN), .D(n7821), .Y(n7840));
  XOR2X1  g04638(.A(n7840), .B(n7839), .Y(n7841));
  AOI22X1 g04639(.A0(n7730), .A1(n7841), .B0(n7729), .B1(P3_EBX_REG_20__SCAN_IN), .Y(n7842));
  NAND2X1 g04640(.A(n7842), .B(n7838), .Y(P3_U2683));
  NAND3X1 g04641(.A(n7728), .B(n7504), .C(n3774), .Y(n7844));
  NOR3X1  g04642(.A(n7834), .B(n7839), .C(n7833), .Y(n7845));
  XOR2X1  g04643(.A(n7845), .B(P3_EBX_REG_21__SCAN_IN), .Y(n7846));
  AOI22X1 g04644(.A0(n7730), .A1(n7846), .B0(n7729), .B1(P3_EBX_REG_21__SCAN_IN), .Y(n7847));
  NAND2X1 g04645(.A(n7847), .B(n7844), .Y(P3_U2682));
  NAND3X1 g04646(.A(n7728), .B(n7521), .C(n3774), .Y(n7849));
  INVX1   g04647(.A(P3_EBX_REG_21__SCAN_IN), .Y(n7850));
  NOR4X1  g04648(.A(n7850), .B(n7839), .C(n7833), .D(n7834), .Y(n7851));
  XOR2X1  g04649(.A(n7851), .B(P3_EBX_REG_22__SCAN_IN), .Y(n7852));
  AOI22X1 g04650(.A0(n7730), .A1(n7852), .B0(n7729), .B1(P3_EBX_REG_22__SCAN_IN), .Y(n7853));
  NAND2X1 g04651(.A(n7853), .B(n7849), .Y(P3_U2681));
  NAND3X1 g04652(.A(n7728), .B(n7567), .C(n3774), .Y(n7855));
  INVX1   g04653(.A(P3_EBX_REG_23__SCAN_IN), .Y(n7856));
  NAND3X1 g04654(.A(n7845), .B(P3_EBX_REG_22__SCAN_IN), .C(P3_EBX_REG_21__SCAN_IN), .Y(n7857));
  XOR2X1  g04655(.A(n7857), .B(n7856), .Y(n7858));
  AOI22X1 g04656(.A0(n7730), .A1(n7858), .B0(n7729), .B1(P3_EBX_REG_23__SCAN_IN), .Y(n7859));
  NAND2X1 g04657(.A(n7859), .B(n7855), .Y(P3_U2680));
  NAND3X1 g04658(.A(n7728), .B(n7589), .C(n3774), .Y(n7861));
  INVX1   g04659(.A(P3_EBX_REG_24__SCAN_IN), .Y(n7862));
  NAND4X1 g04660(.A(P3_EBX_REG_23__SCAN_IN), .B(P3_EBX_REG_22__SCAN_IN), .C(P3_EBX_REG_21__SCAN_IN), .D(n7845), .Y(n7863));
  XOR2X1  g04661(.A(n7863), .B(n7862), .Y(n7864));
  AOI22X1 g04662(.A0(n7730), .A1(n7864), .B0(n7729), .B1(P3_EBX_REG_24__SCAN_IN), .Y(n7865));
  NAND2X1 g04663(.A(n7865), .B(n7861), .Y(P3_U2679));
  NAND3X1 g04664(.A(n7728), .B(n7611), .C(n3774), .Y(n7867));
  NOR3X1  g04665(.A(n7857), .B(n7862), .C(n7856), .Y(n7868));
  XOR2X1  g04666(.A(n7868), .B(P3_EBX_REG_25__SCAN_IN), .Y(n7869));
  AOI22X1 g04667(.A0(n7730), .A1(n7869), .B0(n7729), .B1(P3_EBX_REG_25__SCAN_IN), .Y(n7870));
  NAND2X1 g04668(.A(n7870), .B(n7867), .Y(P3_U2678));
  NAND3X1 g04669(.A(n7728), .B(n7632), .C(n3774), .Y(n7872));
  INVX1   g04670(.A(P3_EBX_REG_25__SCAN_IN), .Y(n7873));
  NOR4X1  g04671(.A(n7873), .B(n7862), .C(n7856), .D(n7857), .Y(n7874));
  XOR2X1  g04672(.A(n7874), .B(P3_EBX_REG_26__SCAN_IN), .Y(n7875));
  AOI22X1 g04673(.A0(n7730), .A1(n7875), .B0(n7729), .B1(P3_EBX_REG_26__SCAN_IN), .Y(n7876));
  NAND2X1 g04674(.A(n7876), .B(n7872), .Y(P3_U2677));
  NAND3X1 g04675(.A(n7728), .B(n7653), .C(n3774), .Y(n7878));
  INVX1   g04676(.A(P3_EBX_REG_27__SCAN_IN), .Y(n7879));
  NAND3X1 g04677(.A(n7868), .B(P3_EBX_REG_26__SCAN_IN), .C(P3_EBX_REG_25__SCAN_IN), .Y(n7880));
  XOR2X1  g04678(.A(n7880), .B(n7879), .Y(n7881));
  AOI22X1 g04679(.A0(n7730), .A1(n7881), .B0(n7729), .B1(P3_EBX_REG_27__SCAN_IN), .Y(n7882));
  NAND2X1 g04680(.A(n7882), .B(n7878), .Y(P3_U2676));
  NAND3X1 g04681(.A(n7728), .B(n7677), .C(n3774), .Y(n7884));
  INVX1   g04682(.A(P3_EBX_REG_28__SCAN_IN), .Y(n7885));
  NAND4X1 g04683(.A(P3_EBX_REG_27__SCAN_IN), .B(P3_EBX_REG_26__SCAN_IN), .C(P3_EBX_REG_25__SCAN_IN), .D(n7868), .Y(n7886));
  XOR2X1  g04684(.A(n7886), .B(n7885), .Y(n7887));
  AOI22X1 g04685(.A0(n7730), .A1(n7887), .B0(n7729), .B1(P3_EBX_REG_28__SCAN_IN), .Y(n7888));
  NAND2X1 g04686(.A(n7888), .B(n7884), .Y(P3_U2675));
  NAND3X1 g04687(.A(n7728), .B(n7696), .C(n3774), .Y(n7890));
  NOR3X1  g04688(.A(n7880), .B(n7885), .C(n7879), .Y(n7891));
  XOR2X1  g04689(.A(n7891), .B(P3_EBX_REG_29__SCAN_IN), .Y(n7892));
  AOI22X1 g04690(.A0(n7730), .A1(n7892), .B0(n7729), .B1(P3_EBX_REG_29__SCAN_IN), .Y(n7893));
  NAND2X1 g04691(.A(n7893), .B(n7890), .Y(P3_U2674));
  NAND3X1 g04692(.A(n7728), .B(n7716), .C(n3774), .Y(n7895));
  INVX1   g04693(.A(P3_EBX_REG_29__SCAN_IN), .Y(n7896));
  NOR4X1  g04694(.A(n7896), .B(n7885), .C(n7879), .D(n7880), .Y(n7897));
  XOR2X1  g04695(.A(n7897), .B(P3_EBX_REG_30__SCAN_IN), .Y(n7898));
  AOI22X1 g04696(.A0(n7730), .A1(n7898), .B0(n7729), .B1(P3_EBX_REG_30__SCAN_IN), .Y(n7899));
  NAND2X1 g04697(.A(n7899), .B(n7895), .Y(P3_U2673));
  INVX1   g04698(.A(P3_EBX_REG_31__SCAN_IN), .Y(n7901));
  NAND2X1 g04699(.A(n7897), .B(P3_EBX_REG_30__SCAN_IN), .Y(n7902));
  XOR2X1  g04700(.A(n7902), .B(P3_EBX_REG_31__SCAN_IN), .Y(n7903));
  OAI22X1 g04701(.A0(n7731), .A1(n7903), .B0(n7728), .B1(n7901), .Y(P3_U2672));
  INVX1   g04702(.A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .Y(n7905));
  INVX1   g04703(.A(n6925), .Y(n7906));
  AOI21X1 g04704(.A0(n3733), .A1(n3721), .B0(n4905), .Y(n7907));
  NOR4X1  g04705(.A(n4968), .B(n3984), .C(n3954), .D(n7907), .Y(n7908));
  NOR3X1  g04706(.A(n7908), .B(n7906), .C(n3939), .Y(n7909));
  INVX1   g04707(.A(n7909), .Y(n7910));
  NOR3X1  g04708(.A(n7908), .B(n6925), .C(n3939), .Y(n7911));
  NAND3X1 g04709(.A(n7907), .B(n3932), .C(n3718), .Y(n7913));
  OAI21X1 g04710(.A0(n3932), .A1(n3726), .B0(n6941), .Y(n7915));
  OAI21X1 g04711(.A0(n7913), .A1(P3_EBX_REG_31__SCAN_IN), .B0(n7915), .Y(n7916));
  INVX1   g04712(.A(n7916), .Y(n7917));
  INVX1   g04713(.A(P3_REIP_REG_0__SCAN_IN), .Y(n7918));
  NOR4X1  g04714(.A(n3932), .B(n3719), .C(n3511), .D(n7908), .Y(n7919));
  INVX1   g04715(.A(n7919), .Y(n7920));
  NOR2X1  g04716(.A(n7920), .B(n7918), .Y(n7921));
  NOR3X1  g04717(.A(n7908), .B(n3728), .C(n3511), .Y(n7922));
  INVX1   g04718(.A(n7922), .Y(n7923));
  NOR3X1  g04719(.A(n7908), .B(n3701), .C(n3511), .Y(n7924));
  INVX1   g04720(.A(n7908), .Y(n7925));
  NOR2X1  g04721(.A(n7908), .B(n3509), .Y(n7926));
  INVX1   g04722(.A(n7926), .Y(n7927));
  OAI22X1 g04723(.A0(n7925), .A1(n7918), .B0(n7905), .B1(n7927), .Y(n7928));
  AOI21X1 g04724(.A0(n7924), .A1(n3541), .B0(n7928), .Y(n7929));
  OAI21X1 g04725(.A0(n7923), .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B0(n7929), .Y(n7930));
  NAND3X1 g04726(.A(n6941), .B(n3931), .C(n3725), .Y(n7931));
  NOR2X1  g04727(.A(n7913), .B(n7901), .Y(n7932));
  INVX1   g04728(.A(n7932), .Y(n7933));
  OAI22X1 g04729(.A0(n7931), .A1(n7918), .B0(n7735), .B1(n7933), .Y(n7934));
  NOR3X1  g04730(.A(n7934), .B(n7930), .C(n7921), .Y(n7935));
  OAI21X1 g04731(.A0(n7917), .A1(n7735), .B0(n7935), .Y(n7936));
  AOI21X1 g04732(.A0(n7911), .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B0(n7936), .Y(n7937));
  OAI21X1 g04733(.A0(n7910), .A1(n7905), .B0(n7937), .Y(P3_U2671));
  NAND2X1 g04734(.A(n7909), .B(n6519), .Y(n7939));
  XOR2X1  g04735(.A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B(n7905), .Y(n7940));
  NAND2X1 g04736(.A(n7940), .B(n7911), .Y(n7941));
  NAND2X1 g04737(.A(n7916), .B(P3_EBX_REG_1__SCAN_IN), .Y(n7942));
  NAND2X1 g04738(.A(n7919), .B(n3399), .Y(n7943));
  NOR2X1  g04739(.A(n3541), .B(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Y(n7944));
  OAI21X1 g04740(.A0(n3833), .A1(n7944), .B0(n7922), .Y(n7945));
  OAI21X1 g04741(.A0(n3833), .A1(n7944), .B0(n7924), .Y(n7946));
  AOI22X1 g04742(.A0(n7908), .A1(P3_REIP_REG_1__SCAN_IN), .B0(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n7926), .Y(n7947));
  NAND4X1 g04743(.A(n7946), .B(n7945), .C(n7943), .D(n7947), .Y(n7948));
  OAI22X1 g04744(.A0(n7931), .A1(P3_REIP_REG_1__SCAN_IN), .B0(n7736), .B1(n7933), .Y(n7949));
  NOR2X1  g04745(.A(n7949), .B(n7948), .Y(n7950));
  NAND4X1 g04746(.A(n7942), .B(n7941), .C(n7939), .D(n7950), .Y(P3_U2670));
  NAND2X1 g04747(.A(n7909), .B(n6525), .Y(n7952));
  NAND2X1 g04748(.A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B(n7905), .Y(n7953));
  XOR2X1  g04749(.A(n7953), .B(n6525), .Y(n7954));
  NAND2X1 g04750(.A(n7954), .B(n7911), .Y(n7955));
  NOR2X1  g04751(.A(n7917), .B(n7744), .Y(n7956));
  XOR2X1  g04752(.A(P3_REIP_REG_2__SCAN_IN), .B(n3399), .Y(n7957));
  NOR2X1  g04753(.A(n7957), .B(n7920), .Y(n7958));
  OAI22X1 g04754(.A0(n7925), .A1(n3396), .B0(n6528), .B1(n7927), .Y(n7959));
  AOI21X1 g04755(.A0(n7924), .A1(n3825), .B0(n7959), .Y(n7960));
  OAI21X1 g04756(.A0(n7923), .A1(n3824), .B0(n7960), .Y(n7961));
  NOR2X1  g04757(.A(P3_EBX_REG_1__SCAN_IN), .B(P3_EBX_REG_0__SCAN_IN), .Y(n7962));
  XOR2X1  g04758(.A(n7962), .B(P3_EBX_REG_2__SCAN_IN), .Y(n7963));
  OAI22X1 g04759(.A0(n7957), .A1(n7931), .B0(n7933), .B1(n7963), .Y(n7964));
  NOR4X1  g04760(.A(n7961), .B(n7958), .C(n7956), .D(n7964), .Y(n7965));
  NAND3X1 g04761(.A(n7965), .B(n7955), .C(n7952), .Y(P3_U2669));
  NAND2X1 g04762(.A(n7909), .B(n6535), .Y(n7967));
  NOR3X1  g04763(.A(n6528), .B(n6519), .C(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .Y(n7968));
  XOR2X1  g04764(.A(n7968), .B(n6534), .Y(n7969));
  NAND2X1 g04765(.A(n7969), .B(n7911), .Y(n7970));
  NOR2X1  g04766(.A(n7917), .B(n7743), .Y(n7971));
  NAND2X1 g04767(.A(P3_REIP_REG_2__SCAN_IN), .B(P3_REIP_REG_1__SCAN_IN), .Y(n7972));
  XOR2X1  g04768(.A(n7972), .B(P3_REIP_REG_3__SCAN_IN), .Y(n7973));
  NOR2X1  g04769(.A(n7973), .B(n7920), .Y(n7974));
  XOR2X1  g04770(.A(n3866), .B(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n7975));
  NAND2X1 g04771(.A(n7975), .B(n7922), .Y(n7976));
  NAND2X1 g04772(.A(n7975), .B(n7924), .Y(n7977));
  AOI22X1 g04773(.A0(n7908), .A1(P3_REIP_REG_3__SCAN_IN), .B0(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(n7926), .Y(n7978));
  NAND3X1 g04774(.A(n7978), .B(n7977), .C(n7976), .Y(n7979));
  NOR3X1  g04775(.A(P3_EBX_REG_2__SCAN_IN), .B(P3_EBX_REG_1__SCAN_IN), .C(P3_EBX_REG_0__SCAN_IN), .Y(n7980));
  XOR2X1  g04776(.A(n7980), .B(P3_EBX_REG_3__SCAN_IN), .Y(n7981));
  OAI22X1 g04777(.A0(n7973), .A1(n7931), .B0(n7933), .B1(n7981), .Y(n7982));
  NOR4X1  g04778(.A(n7979), .B(n7974), .C(n7971), .D(n7982), .Y(n7983));
  NAND3X1 g04779(.A(n7983), .B(n7970), .C(n7967), .Y(P3_U2668));
  INVX1   g04780(.A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .Y(n7985));
  NOR4X1  g04781(.A(n6528), .B(n6519), .C(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .D(n7985), .Y(n7986));
  XOR2X1  g04782(.A(n7986), .B(n6547), .Y(n7987));
  NOR4X1  g04783(.A(n7908), .B(n6925), .C(n3939), .D(n7987), .Y(n7988));
  NOR2X1  g04784(.A(n7917), .B(n7754), .Y(n7989));
  NAND3X1 g04785(.A(P3_REIP_REG_3__SCAN_IN), .B(P3_REIP_REG_2__SCAN_IN), .C(P3_REIP_REG_1__SCAN_IN), .Y(n7990));
  XOR2X1  g04786(.A(n7990), .B(P3_REIP_REG_4__SCAN_IN), .Y(n7991));
  XOR2X1  g04787(.A(n7179), .B(n3531), .Y(n7993));
  NAND2X1 g04788(.A(n7993), .B(n7922), .Y(n7994));
  NAND2X1 g04789(.A(n7926), .B(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .Y(n7995));
  NOR3X1  g04790(.A(P3_STATE2_REG_1__SCAN_IN), .B(P3_STATE2_REG_2__SCAN_IN), .C(P3_STATE2_REG_3__SCAN_IN), .Y(n7996));
  INVX1   g04791(.A(n7996), .Y(n7997));
  AOI21X1 g04792(.A0(n7908), .A1(P3_REIP_REG_4__SCAN_IN), .B0(n4968), .Y(n7999));
  NAND3X1 g04793(.A(n7999), .B(n7995), .C(n7994), .Y(n8000));
  AOI21X1 g04794(.A0(n7993), .A1(n7924), .B0(n8000), .Y(n8001));
  OAI21X1 g04795(.A0(n7991), .A1(n7920), .B0(n8001), .Y(n8002));
  NOR4X1  g04796(.A(P3_EBX_REG_2__SCAN_IN), .B(P3_EBX_REG_1__SCAN_IN), .C(P3_EBX_REG_0__SCAN_IN), .D(P3_EBX_REG_3__SCAN_IN), .Y(n8003));
  NAND3X1 g04797(.A(n7980), .B(n7754), .C(n7743), .Y(n8004));
  OAI21X1 g04798(.A0(n8003), .A1(n7754), .B0(n8004), .Y(n8005));
  OAI22X1 g04799(.A0(n7991), .A1(n7931), .B0(n7933), .B1(n8005), .Y(n8006));
  NOR4X1  g04800(.A(n8002), .B(n7989), .C(n7988), .D(n8006), .Y(n8007));
  OAI21X1 g04801(.A0(n7910), .A1(n6546), .B0(n8007), .Y(P3_U2667));
  NAND2X1 g04802(.A(n7986), .B(n6546), .Y(n8009));
  XOR2X1  g04803(.A(n8009), .B(n6566), .Y(n8010));
  NOR4X1  g04804(.A(n7908), .B(n6925), .C(n3939), .D(n8010), .Y(n8011));
  NOR2X1  g04805(.A(n7917), .B(n7753), .Y(n8012));
  NAND4X1 g04806(.A(P3_REIP_REG_3__SCAN_IN), .B(P3_REIP_REG_2__SCAN_IN), .C(P3_REIP_REG_1__SCAN_IN), .D(P3_REIP_REG_4__SCAN_IN), .Y(n8013));
  XOR2X1  g04807(.A(n8013), .B(P3_REIP_REG_5__SCAN_IN), .Y(n8014));
  INVX1   g04808(.A(n8014), .Y(n8015));
  NAND2X1 g04809(.A(n8015), .B(n7919), .Y(n8016));
  NAND4X1 g04810(.A(n3866), .B(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .D(n7924), .Y(n8017));
  NAND4X1 g04811(.A(n3866), .B(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .D(n7922), .Y(n8018));
  NAND2X1 g04812(.A(n7908), .B(P3_REIP_REG_5__SCAN_IN), .Y(n8019));
  OAI21X1 g04813(.A0(n7908), .A1(n7997), .B0(n8019), .Y(n8020));
  AOI21X1 g04814(.A0(n7926), .A1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B0(n8020), .Y(n8021));
  NAND4X1 g04815(.A(n8018), .B(n8017), .C(n8016), .D(n8021), .Y(n8022));
  XOR2X1  g04816(.A(n8004), .B(n7753), .Y(n8023));
  OAI22X1 g04817(.A0(n8014), .A1(n7931), .B0(n7933), .B1(n8023), .Y(n8024));
  NOR4X1  g04818(.A(n8022), .B(n8012), .C(n8011), .D(n8024), .Y(n8025));
  OAI21X1 g04819(.A0(n7910), .A1(n6566), .B0(n8025), .Y(P3_U2666));
  OAI21X1 g04820(.A0(n8009), .A1(n6567), .B0(n6581), .Y(n8027));
  NOR3X1  g04821(.A(n8009), .B(n6581), .C(n6567), .Y(n8028));
  INVX1   g04822(.A(n8028), .Y(n8029));
  NAND3X1 g04823(.A(n8029), .B(n8027), .C(n7911), .Y(n8030));
  NAND2X1 g04824(.A(n7909), .B(n6581), .Y(n8031));
  NAND2X1 g04825(.A(n7916), .B(P3_EBX_REG_6__SCAN_IN), .Y(n8032));
  OAI21X1 g04826(.A0(n8004), .A1(P3_EBX_REG_5__SCAN_IN), .B0(P3_EBX_REG_6__SCAN_IN), .Y(n8033));
  NOR3X1  g04827(.A(n8004), .B(P3_EBX_REG_6__SCAN_IN), .C(P3_EBX_REG_5__SCAN_IN), .Y(n8034));
  INVX1   g04828(.A(n8034), .Y(n8035));
  NAND2X1 g04829(.A(n8035), .B(n8033), .Y(n8036));
  NOR3X1  g04830(.A(n8036), .B(n7913), .C(n7901), .Y(n8037));
  NOR2X1  g04831(.A(n8013), .B(n3387), .Y(n8038));
  XOR2X1  g04832(.A(n8038), .B(n3384), .Y(n8039));
  NOR2X1  g04833(.A(n8039), .B(n7931), .Y(n8040));
  NOR2X1  g04834(.A(n8039), .B(n7920), .Y(n8041));
  AOI21X1 g04835(.A0(n7908), .A1(P3_REIP_REG_6__SCAN_IN), .B0(n4968), .Y(n8042));
  OAI21X1 g04836(.A0(n7927), .A1(n6577), .B0(n8042), .Y(n8043));
  NOR4X1  g04837(.A(n8041), .B(n8040), .C(n8037), .D(n8043), .Y(n8044));
  NAND4X1 g04838(.A(n8032), .B(n8031), .C(n8030), .D(n8044), .Y(P3_U2665));
  XOR2X1  g04839(.A(n8028), .B(n6594), .Y(n8046));
  NAND2X1 g04840(.A(n8046), .B(n7911), .Y(n8047));
  NAND2X1 g04841(.A(n7909), .B(n6595), .Y(n8048));
  NAND2X1 g04842(.A(n7916), .B(P3_EBX_REG_7__SCAN_IN), .Y(n8049));
  XOR2X1  g04843(.A(n8034), .B(P3_EBX_REG_7__SCAN_IN), .Y(n8050));
  NOR3X1  g04844(.A(n8050), .B(n7913), .C(n7901), .Y(n8051));
  NOR3X1  g04845(.A(n8013), .B(n3384), .C(n3387), .Y(n8052));
  XOR2X1  g04846(.A(n8052), .B(n3381), .Y(n8053));
  NOR2X1  g04847(.A(n8053), .B(n7931), .Y(n8054));
  NOR2X1  g04848(.A(n8053), .B(n7920), .Y(n8055));
  AOI21X1 g04849(.A0(n7908), .A1(P3_REIP_REG_7__SCAN_IN), .B0(n4968), .Y(n8056));
  OAI21X1 g04850(.A0(n7927), .A1(n6592), .B0(n8056), .Y(n8057));
  NOR4X1  g04851(.A(n8055), .B(n8054), .C(n8051), .D(n8057), .Y(n8058));
  NAND4X1 g04852(.A(n8049), .B(n8048), .C(n8047), .D(n8058), .Y(P3_U2664));
  NOR4X1  g04853(.A(n6595), .B(n6581), .C(n6567), .D(n8009), .Y(n8060));
  XOR2X1  g04854(.A(n8060), .B(n6607), .Y(n8061));
  NAND2X1 g04855(.A(n8061), .B(n7911), .Y(n8062));
  NAND2X1 g04856(.A(n7909), .B(n6608), .Y(n8063));
  NAND2X1 g04857(.A(n7916), .B(P3_EBX_REG_8__SCAN_IN), .Y(n8064));
  OAI21X1 g04858(.A0(n8035), .A1(P3_EBX_REG_7__SCAN_IN), .B0(P3_EBX_REG_8__SCAN_IN), .Y(n8065));
  NOR3X1  g04859(.A(n8035), .B(P3_EBX_REG_8__SCAN_IN), .C(P3_EBX_REG_7__SCAN_IN), .Y(n8066));
  INVX1   g04860(.A(n8066), .Y(n8067));
  NAND2X1 g04861(.A(n8067), .B(n8065), .Y(n8068));
  NOR3X1  g04862(.A(n8068), .B(n7913), .C(n7901), .Y(n8069));
  NOR4X1  g04863(.A(n3381), .B(n3384), .C(n3387), .D(n8013), .Y(n8070));
  XOR2X1  g04864(.A(n8070), .B(n3378), .Y(n8071));
  NOR2X1  g04865(.A(n8071), .B(n7931), .Y(n8072));
  NOR2X1  g04866(.A(n8071), .B(n7920), .Y(n8073));
  AOI21X1 g04867(.A0(n7908), .A1(P3_REIP_REG_8__SCAN_IN), .B0(n4968), .Y(n8074));
  OAI21X1 g04868(.A0(n7927), .A1(n6605), .B0(n8074), .Y(n8075));
  NOR4X1  g04869(.A(n8073), .B(n8072), .C(n8069), .D(n8075), .Y(n8076));
  NAND4X1 g04870(.A(n8064), .B(n8063), .C(n8062), .D(n8076), .Y(P3_U2663));
  NOR4X1  g04871(.A(n6621), .B(n6608), .C(n6595), .D(n8029), .Y(n8078));
  AOI21X1 g04872(.A0(n8060), .A1(n6607), .B0(n6620), .Y(n8079));
  NOR2X1  g04873(.A(n8079), .B(n8078), .Y(n8080));
  NAND2X1 g04874(.A(n8080), .B(n7911), .Y(n8081));
  NAND2X1 g04875(.A(n7909), .B(n6621), .Y(n8082));
  NAND2X1 g04876(.A(n7916), .B(P3_EBX_REG_9__SCAN_IN), .Y(n8083));
  XOR2X1  g04877(.A(n8066), .B(P3_EBX_REG_9__SCAN_IN), .Y(n8084));
  NOR3X1  g04878(.A(n8084), .B(n7913), .C(n7901), .Y(n8085));
  NAND2X1 g04879(.A(n8070), .B(P3_REIP_REG_8__SCAN_IN), .Y(n8086));
  XOR2X1  g04880(.A(n8086), .B(P3_REIP_REG_9__SCAN_IN), .Y(n8087));
  NOR2X1  g04881(.A(n8087), .B(n7931), .Y(n8088));
  NOR2X1  g04882(.A(n8087), .B(n7920), .Y(n8089));
  AOI21X1 g04883(.A0(n7908), .A1(P3_REIP_REG_9__SCAN_IN), .B0(n4968), .Y(n8090));
  OAI21X1 g04884(.A0(n7927), .A1(n6624), .B0(n8090), .Y(n8091));
  NOR4X1  g04885(.A(n8089), .B(n8088), .C(n8085), .D(n8091), .Y(n8092));
  NAND4X1 g04886(.A(n8083), .B(n8082), .C(n8081), .D(n8092), .Y(P3_U2662));
  XOR2X1  g04887(.A(n8078), .B(n6633), .Y(n8094));
  NAND2X1 g04888(.A(n8094), .B(n7911), .Y(n8095));
  NAND2X1 g04889(.A(n7909), .B(n6634), .Y(n8096));
  NAND2X1 g04890(.A(n7916), .B(P3_EBX_REG_10__SCAN_IN), .Y(n8097));
  AOI21X1 g04891(.A0(n8066), .A1(n7785), .B0(n7779), .Y(n8098));
  NOR3X1  g04892(.A(n8067), .B(P3_EBX_REG_10__SCAN_IN), .C(P3_EBX_REG_9__SCAN_IN), .Y(n8099));
  NOR4X1  g04893(.A(n8098), .B(n7913), .C(n7901), .D(n8099), .Y(n8100));
  NAND3X1 g04894(.A(n8070), .B(P3_REIP_REG_9__SCAN_IN), .C(P3_REIP_REG_8__SCAN_IN), .Y(n8101));
  XOR2X1  g04895(.A(n8101), .B(P3_REIP_REG_10__SCAN_IN), .Y(n8102));
  NOR2X1  g04896(.A(n8102), .B(n7931), .Y(n8103));
  NOR2X1  g04897(.A(n8102), .B(n7920), .Y(n8104));
  NAND2X1 g04898(.A(n7926), .B(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .Y(n8105));
  AOI21X1 g04899(.A0(n7908), .A1(P3_REIP_REG_10__SCAN_IN), .B0(n4968), .Y(n8106));
  NAND2X1 g04900(.A(n8106), .B(n8105), .Y(n8107));
  NOR4X1  g04901(.A(n8104), .B(n8103), .C(n8100), .D(n8107), .Y(n8108));
  NAND4X1 g04902(.A(n8097), .B(n8096), .C(n8095), .D(n8108), .Y(P3_U2661));
  NAND4X1 g04903(.A(n6633), .B(n6620), .C(n6607), .D(n8060), .Y(n8110));
  XOR2X1  g04904(.A(n8110), .B(n6647), .Y(n8111));
  NAND2X1 g04905(.A(n8111), .B(n7911), .Y(n8112));
  NAND2X1 g04906(.A(n7909), .B(n6647), .Y(n8113));
  NAND2X1 g04907(.A(n7916), .B(P3_EBX_REG_11__SCAN_IN), .Y(n8114));
  XOR2X1  g04908(.A(n8099), .B(P3_EBX_REG_11__SCAN_IN), .Y(n8115));
  NOR3X1  g04909(.A(n8115), .B(n7913), .C(n7901), .Y(n8116));
  NAND4X1 g04910(.A(P3_REIP_REG_10__SCAN_IN), .B(P3_REIP_REG_9__SCAN_IN), .C(P3_REIP_REG_8__SCAN_IN), .D(n8070), .Y(n8117));
  XOR2X1  g04911(.A(n8117), .B(P3_REIP_REG_11__SCAN_IN), .Y(n8118));
  NOR2X1  g04912(.A(n8118), .B(n7931), .Y(n8119));
  NOR2X1  g04913(.A(n8118), .B(n7920), .Y(n8120));
  AOI21X1 g04914(.A0(n7908), .A1(P3_REIP_REG_11__SCAN_IN), .B0(n4968), .Y(n8121));
  OAI21X1 g04915(.A0(n7927), .A1(n6660), .B0(n8121), .Y(n8122));
  NOR4X1  g04916(.A(n8120), .B(n8119), .C(n8116), .D(n8122), .Y(n8123));
  NAND4X1 g04917(.A(n8114), .B(n8113), .C(n8112), .D(n8123), .Y(P3_U2660));
  OAI21X1 g04918(.A0(n8110), .A1(n6647), .B0(n6663), .Y(n8125));
  NOR3X1  g04919(.A(n8110), .B(n6663), .C(n6647), .Y(n8126));
  INVX1   g04920(.A(n8126), .Y(n8127));
  NAND3X1 g04921(.A(n8127), .B(n8125), .C(n7911), .Y(n8128));
  NAND2X1 g04922(.A(n7909), .B(n6663), .Y(n8129));
  NAND2X1 g04923(.A(n7916), .B(P3_EBX_REG_12__SCAN_IN), .Y(n8130));
  INVX1   g04924(.A(P3_EBX_REG_12__SCAN_IN), .Y(n8131));
  AOI21X1 g04925(.A0(n8099), .A1(n7791), .B0(n8131), .Y(n8132));
  NAND3X1 g04926(.A(n8099), .B(n8131), .C(n7791), .Y(n8133));
  INVX1   g04927(.A(n8133), .Y(n8134));
  NOR4X1  g04928(.A(n8132), .B(n7913), .C(n7901), .D(n8134), .Y(n8135));
  NOR2X1  g04929(.A(n8117), .B(n3369), .Y(n8136));
  XOR2X1  g04930(.A(n8136), .B(n3366), .Y(n8137));
  NOR2X1  g04931(.A(n8137), .B(n7931), .Y(n8138));
  NOR2X1  g04932(.A(n8137), .B(n7920), .Y(n8139));
  AOI21X1 g04933(.A0(n7908), .A1(P3_REIP_REG_12__SCAN_IN), .B0(n4968), .Y(n8140));
  OAI21X1 g04934(.A0(n7927), .A1(n6659), .B0(n8140), .Y(n8141));
  NOR4X1  g04935(.A(n8139), .B(n8138), .C(n8135), .D(n8141), .Y(n8142));
  NAND4X1 g04936(.A(n8130), .B(n8129), .C(n8128), .D(n8142), .Y(P3_U2659));
  XOR2X1  g04937(.A(n8126), .B(n6676), .Y(n8144));
  NAND2X1 g04938(.A(n8144), .B(n7911), .Y(n8145));
  NAND2X1 g04939(.A(n7909), .B(n6677), .Y(n8146));
  NAND2X1 g04940(.A(n7916), .B(P3_EBX_REG_13__SCAN_IN), .Y(n8147));
  XOR2X1  g04941(.A(n8133), .B(n7797), .Y(n8148));
  NOR3X1  g04942(.A(n8148), .B(n7913), .C(n7901), .Y(n8149));
  NOR3X1  g04943(.A(n8117), .B(n3366), .C(n3369), .Y(n8150));
  XOR2X1  g04944(.A(n8150), .B(n3363), .Y(n8151));
  NOR2X1  g04945(.A(n8151), .B(n7931), .Y(n8152));
  NOR2X1  g04946(.A(n8151), .B(n7920), .Y(n8153));
  AOI21X1 g04947(.A0(n7908), .A1(P3_REIP_REG_13__SCAN_IN), .B0(n4968), .Y(n8154));
  OAI21X1 g04948(.A0(n7927), .A1(n6674), .B0(n8154), .Y(n8155));
  NOR4X1  g04949(.A(n8153), .B(n8152), .C(n8149), .D(n8155), .Y(n8156));
  NAND4X1 g04950(.A(n8147), .B(n8146), .C(n8145), .D(n8156), .Y(P3_U2658));
  NOR4X1  g04951(.A(n6677), .B(n6663), .C(n6647), .D(n8110), .Y(n8158));
  XOR2X1  g04952(.A(n8158), .B(n6690), .Y(n8159));
  NAND2X1 g04953(.A(n8159), .B(n7911), .Y(n8160));
  NAND2X1 g04954(.A(n7909), .B(n6693), .Y(n8161));
  NAND2X1 g04955(.A(n7916), .B(P3_EBX_REG_14__SCAN_IN), .Y(n8162));
  AOI21X1 g04956(.A0(n8134), .A1(n7797), .B0(n7803), .Y(n8163));
  NOR3X1  g04957(.A(n8133), .B(P3_EBX_REG_14__SCAN_IN), .C(P3_EBX_REG_13__SCAN_IN), .Y(n8164));
  NOR4X1  g04958(.A(n8163), .B(n7913), .C(n7901), .D(n8164), .Y(n8165));
  NOR4X1  g04959(.A(n3363), .B(n3366), .C(n3369), .D(n8117), .Y(n8166));
  XOR2X1  g04960(.A(n8166), .B(n3360), .Y(n8167));
  NOR2X1  g04961(.A(n8167), .B(n7931), .Y(n8168));
  NOR2X1  g04962(.A(n8167), .B(n7920), .Y(n8169));
  AOI21X1 g04963(.A0(n7908), .A1(P3_REIP_REG_14__SCAN_IN), .B0(n4968), .Y(n8170));
  OAI21X1 g04964(.A0(n7927), .A1(n6687), .B0(n8170), .Y(n8171));
  NOR4X1  g04965(.A(n8169), .B(n8168), .C(n8165), .D(n8171), .Y(n8172));
  NAND4X1 g04966(.A(n8162), .B(n8161), .C(n8160), .D(n8172), .Y(P3_U2657));
  NOR4X1  g04967(.A(n6706), .B(n6693), .C(n6677), .D(n8127), .Y(n8174));
  AOI21X1 g04968(.A0(n8158), .A1(n6690), .B0(n6705), .Y(n8175));
  NOR2X1  g04969(.A(n8175), .B(n8174), .Y(n8176));
  NAND2X1 g04970(.A(n8176), .B(n7911), .Y(n8177));
  NAND2X1 g04971(.A(n7909), .B(n6706), .Y(n8178));
  NAND2X1 g04972(.A(n7916), .B(P3_EBX_REG_15__SCAN_IN), .Y(n8179));
  XOR2X1  g04973(.A(n8164), .B(P3_EBX_REG_15__SCAN_IN), .Y(n8180));
  NOR3X1  g04974(.A(n8180), .B(n7913), .C(n7901), .Y(n8181));
  NAND2X1 g04975(.A(n8166), .B(P3_REIP_REG_14__SCAN_IN), .Y(n8182));
  XOR2X1  g04976(.A(n8182), .B(P3_REIP_REG_15__SCAN_IN), .Y(n8183));
  NOR2X1  g04977(.A(n8183), .B(n7931), .Y(n8184));
  NOR2X1  g04978(.A(n8183), .B(n7920), .Y(n8185));
  AOI21X1 g04979(.A0(n7908), .A1(P3_REIP_REG_15__SCAN_IN), .B0(n4968), .Y(n8186));
  OAI21X1 g04980(.A0(n7927), .A1(n6709), .B0(n8186), .Y(n8187));
  NOR4X1  g04981(.A(n8185), .B(n8184), .C(n8181), .D(n8187), .Y(n8188));
  NAND4X1 g04982(.A(n8179), .B(n8178), .C(n8177), .D(n8188), .Y(P3_U2656));
  XOR2X1  g04983(.A(n8174), .B(n6718), .Y(n8190));
  NAND2X1 g04984(.A(n8190), .B(n7911), .Y(n8191));
  NAND2X1 g04985(.A(n7909), .B(n6719), .Y(n8192));
  NAND2X1 g04986(.A(n7916), .B(P3_EBX_REG_16__SCAN_IN), .Y(n8193));
  INVX1   g04987(.A(P3_EBX_REG_16__SCAN_IN), .Y(n8194));
  NOR4X1  g04988(.A(P3_EBX_REG_15__SCAN_IN), .B(P3_EBX_REG_14__SCAN_IN), .C(P3_EBX_REG_13__SCAN_IN), .D(n8133), .Y(n8195));
  NAND3X1 g04989(.A(n8164), .B(n8194), .C(n7814), .Y(n8196));
  OAI21X1 g04990(.A0(n8195), .A1(n8194), .B0(n8196), .Y(n8197));
  NOR3X1  g04991(.A(n8197), .B(n7913), .C(n7901), .Y(n8198));
  NAND3X1 g04992(.A(n8166), .B(P3_REIP_REG_15__SCAN_IN), .C(P3_REIP_REG_14__SCAN_IN), .Y(n8199));
  XOR2X1  g04993(.A(n8199), .B(P3_REIP_REG_16__SCAN_IN), .Y(n8200));
  NOR2X1  g04994(.A(n8200), .B(n7931), .Y(n8201));
  NOR2X1  g04995(.A(n8200), .B(n7920), .Y(n8202));
  NAND2X1 g04996(.A(n7926), .B(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .Y(n8203));
  AOI21X1 g04997(.A0(n7908), .A1(P3_REIP_REG_16__SCAN_IN), .B0(n4968), .Y(n8204));
  NAND2X1 g04998(.A(n8204), .B(n8203), .Y(n8205));
  NOR4X1  g04999(.A(n8202), .B(n8201), .C(n8198), .D(n8205), .Y(n8206));
  NAND4X1 g05000(.A(n8193), .B(n8192), .C(n8191), .D(n8206), .Y(P3_U2655));
  NAND4X1 g05001(.A(n6718), .B(n6705), .C(n6690), .D(n8158), .Y(n8208));
  XOR2X1  g05002(.A(n8208), .B(n6735), .Y(n8209));
  NAND2X1 g05003(.A(n8209), .B(n7911), .Y(n8210));
  NAND2X1 g05004(.A(n7909), .B(n6735), .Y(n8211));
  NAND2X1 g05005(.A(n7916), .B(P3_EBX_REG_17__SCAN_IN), .Y(n8212));
  XOR2X1  g05006(.A(n8196), .B(n7826), .Y(n8213));
  NOR3X1  g05007(.A(n8213), .B(n7913), .C(n7901), .Y(n8214));
  NAND4X1 g05008(.A(P3_REIP_REG_16__SCAN_IN), .B(P3_REIP_REG_15__SCAN_IN), .C(P3_REIP_REG_14__SCAN_IN), .D(n8166), .Y(n8215));
  XOR2X1  g05009(.A(n8215), .B(P3_REIP_REG_17__SCAN_IN), .Y(n8216));
  NOR2X1  g05010(.A(n8216), .B(n7931), .Y(n8217));
  NOR2X1  g05011(.A(n8216), .B(n7920), .Y(n8218));
  AOI21X1 g05012(.A0(n7908), .A1(P3_REIP_REG_17__SCAN_IN), .B0(n4968), .Y(n8219));
  OAI21X1 g05013(.A0(n7927), .A1(n6730), .B0(n8219), .Y(n8220));
  NOR4X1  g05014(.A(n8218), .B(n8217), .C(n8214), .D(n8220), .Y(n8221));
  NAND4X1 g05015(.A(n8212), .B(n8211), .C(n8210), .D(n8221), .Y(P3_U2654));
  OAI21X1 g05016(.A0(n8208), .A1(n6735), .B0(n6749), .Y(n8223));
  NOR3X1  g05017(.A(n8208), .B(n6749), .C(n6735), .Y(n8224));
  INVX1   g05018(.A(n8224), .Y(n8225));
  NAND3X1 g05019(.A(n8225), .B(n8223), .C(n7911), .Y(n8226));
  NAND2X1 g05020(.A(n7909), .B(n6749), .Y(n8227));
  NAND2X1 g05021(.A(n7916), .B(P3_EBX_REG_18__SCAN_IN), .Y(n8228));
  OAI21X1 g05022(.A0(n8196), .A1(P3_EBX_REG_17__SCAN_IN), .B0(P3_EBX_REG_18__SCAN_IN), .Y(n8229));
  NOR3X1  g05023(.A(n8196), .B(P3_EBX_REG_18__SCAN_IN), .C(P3_EBX_REG_17__SCAN_IN), .Y(n8230));
  INVX1   g05024(.A(n8230), .Y(n8231));
  NAND2X1 g05025(.A(n8231), .B(n8229), .Y(n8232));
  NOR3X1  g05026(.A(n8232), .B(n7913), .C(n7901), .Y(n8233));
  NOR2X1  g05027(.A(n8215), .B(n3351), .Y(n8234));
  XOR2X1  g05028(.A(n8234), .B(n3348), .Y(n8235));
  NOR2X1  g05029(.A(n8235), .B(n7931), .Y(n8236));
  NOR2X1  g05030(.A(n8235), .B(n7920), .Y(n8237));
  AOI21X1 g05031(.A0(n7908), .A1(P3_REIP_REG_18__SCAN_IN), .B0(n4968), .Y(n8238));
  OAI21X1 g05032(.A0(n7927), .A1(n6744), .B0(n8238), .Y(n8239));
  NOR4X1  g05033(.A(n8237), .B(n8236), .C(n8233), .D(n8239), .Y(n8240));
  NAND4X1 g05034(.A(n8228), .B(n8227), .C(n8226), .D(n8240), .Y(P3_U2653));
  XOR2X1  g05035(.A(n8224), .B(n6760), .Y(n8242));
  NAND2X1 g05036(.A(n8242), .B(n7911), .Y(n8243));
  INVX1   g05037(.A(n6760), .Y(n8244));
  NAND2X1 g05038(.A(n7909), .B(n8244), .Y(n8245));
  NAND2X1 g05039(.A(n7916), .B(P3_EBX_REG_19__SCAN_IN), .Y(n8246));
  XOR2X1  g05040(.A(n8230), .B(P3_EBX_REG_19__SCAN_IN), .Y(n8247));
  NOR3X1  g05041(.A(n8247), .B(n7913), .C(n7901), .Y(n8248));
  NOR3X1  g05042(.A(n8215), .B(n3348), .C(n3351), .Y(n8249));
  XOR2X1  g05043(.A(n8249), .B(n3345), .Y(n8250));
  NOR2X1  g05044(.A(n8250), .B(n7931), .Y(n8251));
  NOR2X1  g05045(.A(n8250), .B(n7920), .Y(n8252));
  AOI21X1 g05046(.A0(n7908), .A1(P3_REIP_REG_19__SCAN_IN), .B0(n4968), .Y(n8253));
  OAI21X1 g05047(.A0(n7927), .A1(n6758), .B0(n8253), .Y(n8254));
  NOR4X1  g05048(.A(n8252), .B(n8251), .C(n8248), .D(n8254), .Y(n8255));
  NAND4X1 g05049(.A(n8246), .B(n8245), .C(n8243), .D(n8255), .Y(P3_U2652));
  NOR4X1  g05050(.A(n8244), .B(n6749), .C(n6735), .D(n8208), .Y(n8257));
  XOR2X1  g05051(.A(n8257), .B(n6771), .Y(n8258));
  NAND2X1 g05052(.A(n8258), .B(n7911), .Y(n8259));
  INVX1   g05053(.A(n6771), .Y(n8260));
  NAND2X1 g05054(.A(n7909), .B(n8260), .Y(n8261));
  NAND2X1 g05055(.A(n7916), .B(P3_EBX_REG_20__SCAN_IN), .Y(n8262));
  NOR4X1  g05056(.A(n3345), .B(n3348), .C(n3351), .D(n8215), .Y(n8263));
  XOR2X1  g05057(.A(n8263), .B(n3342), .Y(n8264));
  NOR2X1  g05058(.A(n8264), .B(n7931), .Y(n8265));
  AOI21X1 g05059(.A0(n8230), .A1(n7833), .B0(n7839), .Y(n8266));
  NOR3X1  g05060(.A(n8231), .B(P3_EBX_REG_20__SCAN_IN), .C(P3_EBX_REG_19__SCAN_IN), .Y(n8267));
  NOR4X1  g05061(.A(n8266), .B(n7913), .C(n7901), .D(n8267), .Y(n8268));
  AOI22X1 g05062(.A0(n7908), .A1(P3_REIP_REG_20__SCAN_IN), .B0(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B1(n7926), .Y(n8269));
  OAI21X1 g05063(.A0(n8264), .A1(n7920), .B0(n8269), .Y(n8270));
  NOR3X1  g05064(.A(n8270), .B(n8268), .C(n8265), .Y(n8271));
  NAND4X1 g05065(.A(n8262), .B(n8261), .C(n8259), .D(n8271), .Y(P3_U2651));
  INVX1   g05066(.A(n6784), .Y(n8273));
  NOR4X1  g05067(.A(n8273), .B(n8260), .C(n8244), .D(n8225), .Y(n8274));
  AOI21X1 g05068(.A0(n8257), .A1(n6771), .B0(n6784), .Y(n8275));
  NOR2X1  g05069(.A(n8275), .B(n8274), .Y(n8276));
  NAND2X1 g05070(.A(n8276), .B(n7911), .Y(n8277));
  NAND2X1 g05071(.A(n7909), .B(n8273), .Y(n8278));
  NAND2X1 g05072(.A(n7916), .B(P3_EBX_REG_21__SCAN_IN), .Y(n8279));
  NAND2X1 g05073(.A(n8263), .B(P3_REIP_REG_20__SCAN_IN), .Y(n8280));
  XOR2X1  g05074(.A(n8280), .B(P3_REIP_REG_21__SCAN_IN), .Y(n8281));
  NOR2X1  g05075(.A(n8281), .B(n7931), .Y(n8282));
  XOR2X1  g05076(.A(n8267), .B(P3_EBX_REG_21__SCAN_IN), .Y(n8283));
  NOR3X1  g05077(.A(n8283), .B(n7913), .C(n7901), .Y(n8284));
  AOI22X1 g05078(.A0(n7908), .A1(P3_REIP_REG_21__SCAN_IN), .B0(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B1(n7926), .Y(n8285));
  OAI21X1 g05079(.A0(n8281), .A1(n7920), .B0(n8285), .Y(n8286));
  NOR3X1  g05080(.A(n8286), .B(n8284), .C(n8282), .Y(n8287));
  NAND4X1 g05081(.A(n8279), .B(n8278), .C(n8277), .D(n8287), .Y(P3_U2650));
  XOR2X1  g05082(.A(n8274), .B(n6799), .Y(n8289));
  NAND2X1 g05083(.A(n8289), .B(n7911), .Y(n8290));
  INVX1   g05084(.A(n6799), .Y(n8291));
  NAND2X1 g05085(.A(n7909), .B(n8291), .Y(n8292));
  NAND2X1 g05086(.A(n7916), .B(P3_EBX_REG_22__SCAN_IN), .Y(n8293));
  NAND3X1 g05087(.A(n8263), .B(P3_REIP_REG_21__SCAN_IN), .C(P3_REIP_REG_20__SCAN_IN), .Y(n8294));
  XOR2X1  g05088(.A(n8294), .B(P3_REIP_REG_22__SCAN_IN), .Y(n8295));
  AOI22X1 g05089(.A0(n7908), .A1(P3_REIP_REG_22__SCAN_IN), .B0(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(n7926), .Y(n8296));
  OAI21X1 g05090(.A0(n8295), .A1(n7920), .B0(n8296), .Y(n8297));
  INVX1   g05091(.A(n8267), .Y(n8298));
  OAI21X1 g05092(.A0(n8298), .A1(P3_EBX_REG_21__SCAN_IN), .B0(P3_EBX_REG_22__SCAN_IN), .Y(n8299));
  NOR3X1  g05093(.A(n8298), .B(P3_EBX_REG_22__SCAN_IN), .C(P3_EBX_REG_21__SCAN_IN), .Y(n8300));
  INVX1   g05094(.A(n8300), .Y(n8301));
  NAND3X1 g05095(.A(n8301), .B(n8299), .C(n7932), .Y(n8302));
  OAI21X1 g05096(.A0(n8295), .A1(n7931), .B0(n8302), .Y(n8303));
  NOR2X1  g05097(.A(n8303), .B(n8297), .Y(n8304));
  NAND4X1 g05098(.A(n8293), .B(n8292), .C(n8290), .D(n8304), .Y(P3_U2649));
  INVX1   g05099(.A(n6815), .Y(n8306));
  NAND4X1 g05100(.A(n6799), .B(n6784), .C(n6771), .D(n8257), .Y(n8307));
  XOR2X1  g05101(.A(n8307), .B(n8306), .Y(n8308));
  NAND2X1 g05102(.A(n8308), .B(n7911), .Y(n8309));
  NAND2X1 g05103(.A(n7909), .B(n8306), .Y(n8310));
  NAND2X1 g05104(.A(n7916), .B(P3_EBX_REG_23__SCAN_IN), .Y(n8311));
  NAND4X1 g05105(.A(P3_REIP_REG_22__SCAN_IN), .B(P3_REIP_REG_21__SCAN_IN), .C(P3_REIP_REG_20__SCAN_IN), .D(n8263), .Y(n8312));
  XOR2X1  g05106(.A(n8312), .B(P3_REIP_REG_23__SCAN_IN), .Y(n8313));
  NOR2X1  g05107(.A(n8313), .B(n7931), .Y(n8314));
  NOR2X1  g05108(.A(n8313), .B(n7920), .Y(n8315));
  XOR2X1  g05109(.A(n8300), .B(P3_EBX_REG_23__SCAN_IN), .Y(n8316));
  NOR3X1  g05110(.A(n8316), .B(n7913), .C(n7901), .Y(n8317));
  OAI22X1 g05111(.A0(n7925), .A1(n3333), .B0(n6821), .B1(n7927), .Y(n8318));
  NOR4X1  g05112(.A(n8317), .B(n8315), .C(n8314), .D(n8318), .Y(n8319));
  NAND4X1 g05113(.A(n8311), .B(n8310), .C(n8309), .D(n8319), .Y(P3_U2648));
  INVX1   g05114(.A(n6828), .Y(n8321));
  NAND2X1 g05115(.A(n7909), .B(n8321), .Y(n8322));
  OAI21X1 g05116(.A0(n8307), .A1(n8306), .B0(n8321), .Y(n8323));
  NOR3X1  g05117(.A(n8307), .B(n8321), .C(n8306), .Y(n8324));
  INVX1   g05118(.A(n8324), .Y(n8325));
  NAND3X1 g05119(.A(n8325), .B(n8323), .C(n7911), .Y(n8326));
  NAND2X1 g05120(.A(n7916), .B(P3_EBX_REG_24__SCAN_IN), .Y(n8327));
  OAI21X1 g05121(.A0(n8301), .A1(P3_EBX_REG_23__SCAN_IN), .B0(P3_EBX_REG_24__SCAN_IN), .Y(n8328));
  NOR3X1  g05122(.A(n8301), .B(P3_EBX_REG_24__SCAN_IN), .C(P3_EBX_REG_23__SCAN_IN), .Y(n8329));
  INVX1   g05123(.A(n8329), .Y(n8330));
  NAND3X1 g05124(.A(n8330), .B(n8328), .C(n7932), .Y(n8331));
  AOI22X1 g05125(.A0(n7908), .A1(P3_REIP_REG_24__SCAN_IN), .B0(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B1(n7926), .Y(n8332));
  NAND3X1 g05126(.A(n8332), .B(n8331), .C(n8327), .Y(n8333));
  NOR2X1  g05127(.A(n8312), .B(n3333), .Y(n8334));
  XOR2X1  g05128(.A(n8334), .B(n3330), .Y(n8335));
  AOI21X1 g05129(.A0(n7931), .A1(n7920), .B0(n8335), .Y(n8336));
  NOR2X1  g05130(.A(n8336), .B(n8333), .Y(n8337));
  NAND3X1 g05131(.A(n8337), .B(n8326), .C(n8322), .Y(P3_U2647));
  XOR2X1  g05132(.A(n8324), .B(n6843), .Y(n8339));
  NOR3X1  g05133(.A(n8312), .B(n3330), .C(n3333), .Y(n8340));
  XOR2X1  g05134(.A(n8340), .B(P3_REIP_REG_25__SCAN_IN), .Y(n8341));
  NAND2X1 g05135(.A(n8341), .B(n7919), .Y(n8342));
  NAND4X1 g05136(.A(n6941), .B(n3931), .C(n3725), .D(n8341), .Y(n8343));
  NAND2X1 g05137(.A(n7916), .B(P3_EBX_REG_25__SCAN_IN), .Y(n8344));
  XOR2X1  g05138(.A(n8329), .B(n7873), .Y(n8345));
  OAI22X1 g05139(.A0(n7925), .A1(n3327), .B0(n6841), .B1(n7927), .Y(n8346));
  AOI21X1 g05140(.A0(n8345), .A1(n7932), .B0(n8346), .Y(n8347));
  NAND4X1 g05141(.A(n8344), .B(n8343), .C(n8342), .D(n8347), .Y(n8348));
  AOI21X1 g05142(.A0(n8339), .A1(n7911), .B0(n8348), .Y(n8349));
  OAI21X1 g05143(.A0(n7910), .A1(n6843), .B0(n8349), .Y(P3_U2646));
  INVX1   g05144(.A(n6856), .Y(n8351));
  NOR4X1  g05145(.A(n6844), .B(n8321), .C(n8306), .D(n8307), .Y(n8352));
  XOR2X1  g05146(.A(n8352), .B(n8351), .Y(n8353));
  NOR4X1  g05147(.A(n7908), .B(n6925), .C(n3939), .D(n8353), .Y(n8354));
  NOR4X1  g05148(.A(n3327), .B(n3330), .C(n3333), .D(n8312), .Y(n8355));
  XOR2X1  g05149(.A(n8355), .B(n3324), .Y(n8356));
  NOR2X1  g05150(.A(n8356), .B(n7920), .Y(n8357));
  NOR2X1  g05151(.A(n8356), .B(n7931), .Y(n8358));
  NAND2X1 g05152(.A(n7916), .B(P3_EBX_REG_26__SCAN_IN), .Y(n8359));
  NAND4X1 g05153(.A(n7873), .B(n7862), .C(n7856), .D(n8300), .Y(n8360));
  NOR3X1  g05154(.A(n8330), .B(P3_EBX_REG_26__SCAN_IN), .C(P3_EBX_REG_25__SCAN_IN), .Y(n8361));
  AOI21X1 g05155(.A0(n8360), .A1(P3_EBX_REG_26__SCAN_IN), .B0(n8361), .Y(n8362));
  OAI22X1 g05156(.A0(n7925), .A1(n3324), .B0(n6854), .B1(n7927), .Y(n8363));
  AOI21X1 g05157(.A0(n8362), .A1(n7932), .B0(n8363), .Y(n8364));
  NAND2X1 g05158(.A(n8364), .B(n8359), .Y(n8365));
  NOR4X1  g05159(.A(n8358), .B(n8357), .C(n8354), .D(n8365), .Y(n8366));
  OAI21X1 g05160(.A0(n7910), .A1(n6856), .B0(n8366), .Y(P3_U2645));
  INVX1   g05161(.A(n6869), .Y(n8368));
  NOR4X1  g05162(.A(n8368), .B(n8351), .C(n6844), .D(n8325), .Y(n8369));
  AOI21X1 g05163(.A0(n8352), .A1(n6856), .B0(n6869), .Y(n8370));
  NOR2X1  g05164(.A(n8370), .B(n8369), .Y(n8371));
  NAND2X1 g05165(.A(n8355), .B(P3_REIP_REG_26__SCAN_IN), .Y(n8372));
  XOR2X1  g05166(.A(n8372), .B(n3321), .Y(n8373));
  NAND2X1 g05167(.A(n8373), .B(n7919), .Y(n8374));
  NAND4X1 g05168(.A(n6941), .B(n3931), .C(n3725), .D(n8373), .Y(n8375));
  NAND2X1 g05169(.A(n7916), .B(P3_EBX_REG_27__SCAN_IN), .Y(n8376));
  XOR2X1  g05170(.A(n8361), .B(n7879), .Y(n8377));
  OAI22X1 g05171(.A0(n7925), .A1(n3321), .B0(n6872), .B1(n7927), .Y(n8378));
  AOI21X1 g05172(.A0(n8377), .A1(n7932), .B0(n8378), .Y(n8379));
  NAND4X1 g05173(.A(n8376), .B(n8375), .C(n8374), .D(n8379), .Y(n8380));
  AOI21X1 g05174(.A0(n8371), .A1(n7911), .B0(n8380), .Y(n8381));
  OAI21X1 g05175(.A0(n7910), .A1(n6869), .B0(n8381), .Y(P3_U2644));
  XOR2X1  g05176(.A(n8369), .B(n6885), .Y(n8383));
  NAND3X1 g05177(.A(n8355), .B(P3_REIP_REG_27__SCAN_IN), .C(P3_REIP_REG_26__SCAN_IN), .Y(n8384));
  XOR2X1  g05178(.A(n8384), .B(P3_REIP_REG_28__SCAN_IN), .Y(n8385));
  NOR2X1  g05179(.A(n8385), .B(n7931), .Y(n8386));
  NOR2X1  g05180(.A(n7917), .B(n7885), .Y(n8387));
  NOR4X1  g05181(.A(P3_EBX_REG_27__SCAN_IN), .B(P3_EBX_REG_26__SCAN_IN), .C(P3_EBX_REG_25__SCAN_IN), .D(n8330), .Y(n8388));
  NAND3X1 g05182(.A(n8361), .B(n7885), .C(n7879), .Y(n8389));
  OAI21X1 g05183(.A0(n8388), .A1(n7885), .B0(n8389), .Y(n8390));
  AOI22X1 g05184(.A0(n7908), .A1(P3_REIP_REG_28__SCAN_IN), .B0(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B1(n7926), .Y(n8391));
  OAI21X1 g05185(.A0(n8390), .A1(n7933), .B0(n8391), .Y(n8392));
  NOR3X1  g05186(.A(n8392), .B(n8387), .C(n8386), .Y(n8393));
  OAI21X1 g05187(.A0(n8385), .A1(n7920), .B0(n8393), .Y(n8394));
  AOI21X1 g05188(.A0(n8383), .A1(n7911), .B0(n8394), .Y(n8395));
  OAI21X1 g05189(.A0(n7910), .A1(n6885), .B0(n8395), .Y(P3_U2643));
  INVX1   g05190(.A(n6897), .Y(n8397));
  NAND4X1 g05191(.A(n6885), .B(n6869), .C(n6856), .D(n8352), .Y(n8398));
  XOR2X1  g05192(.A(n8398), .B(n8397), .Y(n8399));
  NAND4X1 g05193(.A(P3_REIP_REG_28__SCAN_IN), .B(P3_REIP_REG_27__SCAN_IN), .C(P3_REIP_REG_26__SCAN_IN), .D(n8355), .Y(n8400));
  XOR2X1  g05194(.A(n8400), .B(n3315), .Y(n8401));
  NAND2X1 g05195(.A(n8401), .B(n7919), .Y(n8402));
  NAND4X1 g05196(.A(n6941), .B(n3931), .C(n3725), .D(n8401), .Y(n8403));
  NAND2X1 g05197(.A(n7916), .B(P3_EBX_REG_29__SCAN_IN), .Y(n8404));
  XOR2X1  g05198(.A(n8389), .B(P3_EBX_REG_29__SCAN_IN), .Y(n8405));
  OAI22X1 g05199(.A0(n7925), .A1(n3315), .B0(n6903), .B1(n7927), .Y(n8406));
  AOI21X1 g05200(.A0(n8405), .A1(n7932), .B0(n8406), .Y(n8407));
  NAND4X1 g05201(.A(n8404), .B(n8403), .C(n8402), .D(n8407), .Y(n8408));
  AOI21X1 g05202(.A0(n8399), .A1(n7911), .B0(n8408), .Y(n8409));
  OAI21X1 g05203(.A0(n7910), .A1(n6897), .B0(n8409), .Y(P3_U2642));
  NOR2X1  g05204(.A(n8398), .B(n8397), .Y(n8411));
  XOR2X1  g05205(.A(n8411), .B(n6913), .Y(n8412));
  NOR2X1  g05206(.A(n8400), .B(n3315), .Y(n8413));
  XOR2X1  g05207(.A(n8413), .B(P3_REIP_REG_30__SCAN_IN), .Y(n8414));
  NAND2X1 g05208(.A(n8414), .B(n7919), .Y(n8415));
  NAND4X1 g05209(.A(n6941), .B(n3931), .C(n3725), .D(n8414), .Y(n8416));
  NAND2X1 g05210(.A(n7916), .B(P3_EBX_REG_30__SCAN_IN), .Y(n8417));
  INVX1   g05211(.A(P3_EBX_REG_30__SCAN_IN), .Y(n8418));
  NOR2X1  g05212(.A(n8389), .B(P3_EBX_REG_29__SCAN_IN), .Y(n8419));
  XOR2X1  g05213(.A(n8419), .B(n8418), .Y(n8420));
  OAI22X1 g05214(.A0(n7925), .A1(n3310), .B0(n6911), .B1(n7927), .Y(n8421));
  AOI21X1 g05215(.A0(n8420), .A1(n7932), .B0(n8421), .Y(n8422));
  NAND4X1 g05216(.A(n8417), .B(n8416), .C(n8415), .D(n8422), .Y(n8423));
  AOI21X1 g05217(.A0(n8412), .A1(n7911), .B0(n8423), .Y(n8424));
  OAI21X1 g05218(.A0(n7910), .A1(n6913), .B0(n8424), .Y(P3_U2641));
  NOR3X1  g05219(.A(n8400), .B(n3310), .C(n3315), .Y(n8426));
  XOR2X1  g05220(.A(n8426), .B(n6477), .Y(n8427));
  NOR2X1  g05221(.A(n8427), .B(n7931), .Y(n8428));
  NOR2X1  g05222(.A(n8427), .B(n7920), .Y(n8429));
  NOR2X1  g05223(.A(n7917), .B(n7901), .Y(n8430));
  NOR3X1  g05224(.A(n8389), .B(P3_EBX_REG_30__SCAN_IN), .C(P3_EBX_REG_29__SCAN_IN), .Y(n8431));
  XOR2X1  g05225(.A(n8431), .B(P3_EBX_REG_31__SCAN_IN), .Y(n8432));
  AOI22X1 g05226(.A0(n7908), .A1(P3_REIP_REG_31__SCAN_IN), .B0(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B1(n7926), .Y(n8433));
  OAI21X1 g05227(.A0(n8432), .A1(n7933), .B0(n8433), .Y(n8434));
  NOR4X1  g05228(.A(n8430), .B(n8429), .C(n8428), .D(n8434), .Y(n8435));
  NAND2X1 g05229(.A(n8411), .B(n6913), .Y(n8436));
  XOR2X1  g05230(.A(n8436), .B(n7906), .Y(n8437));
  AOI21X1 g05231(.A0(n7909), .A1(n7906), .B0(n8437), .Y(n8438));
  NAND3X1 g05232(.A(n7925), .B(n7906), .C(P3_STATE2_REG_1__SCAN_IN), .Y(n8439));
  OAI21X1 g05233(.A0(n8439), .A1(n8438), .B0(n8435), .Y(P3_U2640));
  NOR4X1  g05234(.A(P3_DATAWIDTH_REG_15__SCAN_IN), .B(P3_DATAWIDTH_REG_14__SCAN_IN), .C(P3_DATAWIDTH_REG_13__SCAN_IN), .D(P3_DATAWIDTH_REG_16__SCAN_IN), .Y(n8441));
  NOR4X1  g05235(.A(P3_DATAWIDTH_REG_12__SCAN_IN), .B(P3_DATAWIDTH_REG_11__SCAN_IN), .C(P3_DATAWIDTH_REG_10__SCAN_IN), .D(P3_DATAWIDTH_REG_26__SCAN_IN), .Y(n8442));
  NOR4X1  g05236(.A(P3_DATAWIDTH_REG_7__SCAN_IN), .B(P3_DATAWIDTH_REG_6__SCAN_IN), .C(P3_DATAWIDTH_REG_5__SCAN_IN), .D(P3_DATAWIDTH_REG_8__SCAN_IN), .Y(n8443));
  NOR4X1  g05237(.A(P3_DATAWIDTH_REG_4__SCAN_IN), .B(P3_DATAWIDTH_REG_3__SCAN_IN), .C(P3_DATAWIDTH_REG_2__SCAN_IN), .D(P3_DATAWIDTH_REG_17__SCAN_IN), .Y(n8444));
  NAND4X1 g05238(.A(n8443), .B(n8442), .C(n8441), .D(n8444), .Y(n8445));
  NOR4X1  g05239(.A(P3_DATAWIDTH_REG_22__SCAN_IN), .B(P3_DATAWIDTH_REG_21__SCAN_IN), .C(P3_DATAWIDTH_REG_20__SCAN_IN), .D(P3_DATAWIDTH_REG_23__SCAN_IN), .Y(n8446));
  INVX1   g05240(.A(P3_DATAWIDTH_REG_0__SCAN_IN), .Y(n8447));
  NOR2X1  g05241(.A(n3445), .B(n8447), .Y(n8448));
  NOR3X1  g05242(.A(n8448), .B(P3_DATAWIDTH_REG_19__SCAN_IN), .C(P3_DATAWIDTH_REG_18__SCAN_IN), .Y(n8449));
  NOR4X1  g05243(.A(P3_DATAWIDTH_REG_29__SCAN_IN), .B(P3_DATAWIDTH_REG_28__SCAN_IN), .C(P3_DATAWIDTH_REG_27__SCAN_IN), .D(P3_DATAWIDTH_REG_30__SCAN_IN), .Y(n8450));
  NOR4X1  g05244(.A(P3_DATAWIDTH_REG_25__SCAN_IN), .B(P3_DATAWIDTH_REG_24__SCAN_IN), .C(P3_DATAWIDTH_REG_9__SCAN_IN), .D(P3_DATAWIDTH_REG_31__SCAN_IN), .Y(n8451));
  NAND4X1 g05245(.A(n8450), .B(n8449), .C(n8446), .D(n8451), .Y(n8452));
  NOR2X1  g05246(.A(n8452), .B(n8445), .Y(n8453));
  NAND3X1 g05247(.A(n8453), .B(n3399), .C(n3445), .Y(n8454));
  NOR2X1  g05248(.A(P3_DATAWIDTH_REG_1__SCAN_IN), .B(P3_DATAWIDTH_REG_0__SCAN_IN), .Y(n8455));
  NAND3X1 g05249(.A(n8455), .B(n8453), .C(n7918), .Y(n8456));
  OAI21X1 g05250(.A0(n8452), .A1(n8445), .B0(P3_BYTEENABLE_REG_3__SCAN_IN), .Y(n8457));
  NAND3X1 g05251(.A(n8457), .B(n8456), .C(n8454), .Y(P3_U2639));
  NAND2X1 g05252(.A(P3_REIP_REG_1__SCAN_IN), .B(P3_REIP_REG_0__SCAN_IN), .Y(n8459));
  AOI21X1 g05253(.A0(n7918), .A1(P3_DATAWIDTH_REG_0__SCAN_IN), .B0(n8455), .Y(n8460));
  OAI21X1 g05254(.A0(n8460), .A1(P3_REIP_REG_1__SCAN_IN), .B0(n8459), .Y(n8461));
  NAND2X1 g05255(.A(n8461), .B(n8453), .Y(n8462));
  OAI21X1 g05256(.A0(n8453), .A1(n3299), .B0(n8462), .Y(P3_U3292));
  NAND2X1 g05257(.A(n8453), .B(P3_REIP_REG_1__SCAN_IN), .Y(n8464));
  OAI21X1 g05258(.A0(n8452), .A1(n8445), .B0(P3_BYTEENABLE_REG_1__SCAN_IN), .Y(n8465));
  NAND3X1 g05259(.A(n8465), .B(n8464), .C(n8456), .Y(P3_U2638));
  OAI21X1 g05260(.A0(P3_REIP_REG_1__SCAN_IN), .A1(P3_REIP_REG_0__SCAN_IN), .B0(n8453), .Y(n8467));
  OAI21X1 g05261(.A0(n8453), .A1(n3307), .B0(n8467), .Y(P3_U3293));
  OAI21X1 g05262(.A0(P3_STATE_REG_0__SCAN_IN), .A1(n3296), .B0(P3_W_R_N_REG_SCAN_IN), .Y(n8469));
  OAI21X1 g05263(.A0(n3301), .A1(P3_READREQUEST_REG_SCAN_IN), .B0(n8469), .Y(P3_U3294));
  NAND2X1 g05264(.A(n3955), .B(n3897), .Y(n8471));
  NOR2X1  g05265(.A(n4905), .B(n3912), .Y(n8472));
  OAI21X1 g05266(.A0(n8472), .A1(n3959), .B0(n8471), .Y(P3_U2637));
  INVX1   g05267(.A(n8472), .Y(n8474));
  OAI21X1 g05268(.A0(n4905), .A1(n3912), .B0(P3_MORE_REG_SCAN_IN), .Y(n8475));
  OAI21X1 g05269(.A0(n8474), .A1(n3927), .B0(n8475), .Y(P3_U3295));
  AOI22X1 g05270(.A0(n3416), .A1(n3294), .B0(P3_STATEBS16_REG_SCAN_IN), .B1(n3442), .Y(n8477));
  OAI21X1 g05271(.A0(n3442), .A1(n3439), .B0(n8477), .Y(P3_U2636));
  INVX1   g05272(.A(n7907), .Y(n8479));
  OAI21X1 g05273(.A0(n3958), .A1(n3407), .B0(n4909), .Y(n8480));
  AOI21X1 g05274(.A0(n8480), .A1(n3510), .B0(n4073), .Y(n8481));
  NAND2X1 g05275(.A(n8481), .B(n8479), .Y(n8482));
  OAI21X1 g05276(.A0(n3730), .A1(n3727), .B0(n3726), .Y(n8483));
  OAI21X1 g05277(.A0(n3404), .A1(n3403), .B0(P3_STATE2_REG_2__SCAN_IN), .Y(n8484));
  AOI21X1 g05278(.A0(n3730), .A1(n3944), .B0(n8484), .Y(n8485));
  AOI21X1 g05279(.A0(n8485), .A1(n8483), .B0(n3510), .Y(n8486));
  OAI21X1 g05280(.A0(n8486), .A1(n3979), .B0(n8482), .Y(n8487));
  OAI21X1 g05281(.A0(n8482), .A1(n3409), .B0(n8487), .Y(P3_U3296));
  OAI21X1 g05282(.A0(P3_STATE_REG_0__SCAN_IN), .A1(n3296), .B0(P3_D_C_N_REG_SCAN_IN), .Y(n8489));
  INVX1   g05283(.A(P3_CODEFETCH_REG_SCAN_IN), .Y(n8490));
  AOI22X1 g05284(.A0(n3300), .A1(n8490), .B0(n3294), .B1(n3416), .Y(n8491));
  NAND2X1 g05285(.A(n8491), .B(n8489), .Y(P3_U2635));
  NAND3X1 g05286(.A(P3_MEMORYFETCH_REG_SCAN_IN), .B(n3294), .C(P3_STATE_REG_1__SCAN_IN), .Y(n8493));
  OAI21X1 g05287(.A0(n3300), .A1(n3290), .B0(n8493), .Y(P3_U3297));
  OAI22X1 g05288(.A0(n7997), .A1(n3510), .B0(n8490), .B1(n7907), .Y(P3_U2634));
  NAND2X1 g05289(.A(P3_ADS_N_REG_SCAN_IN), .B(P3_STATE_REG_0__SCAN_IN), .Y(n8497));
  NAND2X1 g05290(.A(n8497), .B(n3442), .Y(P3_U2633));
  NAND2X1 g05291(.A(n3813), .B(P3_STATE2_REG_2__SCAN_IN), .Y(n8499));
  OAI21X1 g05292(.A0(n7907), .A1(n7996), .B0(n8499), .Y(n8500));
  NAND3X1 g05293(.A(n8479), .B(n7997), .C(P3_READREQUEST_REG_SCAN_IN), .Y(n8501));
  NAND2X1 g05294(.A(n8501), .B(n8500), .Y(P3_U3298));
  OAI22X1 g05295(.A0(n7996), .A1(n7907), .B0(n3699), .B1(n3511), .Y(n8503));
  NAND3X1 g05296(.A(n8479), .B(n7997), .C(P3_MEMORYFETCH_REG_SCAN_IN), .Y(n8504));
  NAND2X1 g05297(.A(n8504), .B(n8503), .Y(P3_U3299));
  INVX1   g05298(.A(P2_STATE_REG_0__SCAN_IN), .Y(n8506));
  NAND3X1 g05299(.A(P2_BYTEENABLE_REG_3__SCAN_IN), .B(n8506), .C(P2_STATE_REG_1__SCAN_IN), .Y(n8507));
  INVX1   g05300(.A(P2_STATE_REG_1__SCAN_IN), .Y(n8508));
  OAI21X1 g05301(.A0(P2_STATE_REG_0__SCAN_IN), .A1(n8508), .B0(P2_BE_N_REG_3__SCAN_IN), .Y(n8509));
  NAND2X1 g05302(.A(n8509), .B(n8507), .Y(P2_U3585));
  INVX1   g05303(.A(P2_BYTEENABLE_REG_2__SCAN_IN), .Y(n8511));
  NOR2X1  g05304(.A(P2_STATE_REG_0__SCAN_IN), .B(n8508), .Y(n8512));
  INVX1   g05305(.A(n8512), .Y(n8513));
  OAI21X1 g05306(.A0(P2_STATE_REG_0__SCAN_IN), .A1(n8508), .B0(P2_BE_N_REG_2__SCAN_IN), .Y(n8514));
  OAI21X1 g05307(.A0(n8513), .A1(n8511), .B0(n8514), .Y(P2_U3586));
  NAND3X1 g05308(.A(P2_BYTEENABLE_REG_1__SCAN_IN), .B(n8506), .C(P2_STATE_REG_1__SCAN_IN), .Y(n8516));
  OAI21X1 g05309(.A0(P2_STATE_REG_0__SCAN_IN), .A1(n8508), .B0(P2_BE_N_REG_1__SCAN_IN), .Y(n8517));
  NAND2X1 g05310(.A(n8517), .B(n8516), .Y(P2_U3587));
  NAND3X1 g05311(.A(P2_BYTEENABLE_REG_0__SCAN_IN), .B(n8506), .C(P2_STATE_REG_1__SCAN_IN), .Y(n8519));
  OAI21X1 g05312(.A0(P2_STATE_REG_0__SCAN_IN), .A1(n8508), .B0(P2_BE_N_REG_0__SCAN_IN), .Y(n8520));
  NAND2X1 g05313(.A(n8520), .B(n8519), .Y(P2_U3588));
  INVX1   g05314(.A(P2_REIP_REG_30__SCAN_IN), .Y(n8522));
  NAND3X1 g05315(.A(n8506), .B(P2_STATE_REG_1__SCAN_IN), .C(P2_STATE_REG_2__SCAN_IN), .Y(n8523));
  NOR3X1  g05316(.A(P2_STATE_REG_0__SCAN_IN), .B(n8508), .C(P2_STATE_REG_2__SCAN_IN), .Y(n8524));
  AOI22X1 g05317(.A0(n8513), .A1(P2_ADDRESS_REG_29__SCAN_IN), .B0(P2_REIP_REG_31__SCAN_IN), .B1(n8524), .Y(n8525));
  OAI21X1 g05318(.A0(n8523), .A1(n8522), .B0(n8525), .Y(P2_U3241));
  INVX1   g05319(.A(P2_REIP_REG_29__SCAN_IN), .Y(n8527));
  AOI22X1 g05320(.A0(n8513), .A1(P2_ADDRESS_REG_28__SCAN_IN), .B0(P2_REIP_REG_30__SCAN_IN), .B1(n8524), .Y(n8528));
  OAI21X1 g05321(.A0(n8523), .A1(n8527), .B0(n8528), .Y(P2_U3240));
  INVX1   g05322(.A(P2_REIP_REG_28__SCAN_IN), .Y(n8530));
  AOI22X1 g05323(.A0(n8513), .A1(P2_ADDRESS_REG_27__SCAN_IN), .B0(P2_REIP_REG_29__SCAN_IN), .B1(n8524), .Y(n8531));
  OAI21X1 g05324(.A0(n8523), .A1(n8530), .B0(n8531), .Y(P2_U3239));
  INVX1   g05325(.A(P2_REIP_REG_27__SCAN_IN), .Y(n8533));
  AOI22X1 g05326(.A0(n8513), .A1(P2_ADDRESS_REG_26__SCAN_IN), .B0(P2_REIP_REG_28__SCAN_IN), .B1(n8524), .Y(n8534));
  OAI21X1 g05327(.A0(n8523), .A1(n8533), .B0(n8534), .Y(P2_U3238));
  INVX1   g05328(.A(P2_REIP_REG_26__SCAN_IN), .Y(n8536));
  AOI22X1 g05329(.A0(n8513), .A1(P2_ADDRESS_REG_25__SCAN_IN), .B0(P2_REIP_REG_27__SCAN_IN), .B1(n8524), .Y(n8537));
  OAI21X1 g05330(.A0(n8523), .A1(n8536), .B0(n8537), .Y(P2_U3237));
  INVX1   g05331(.A(P2_REIP_REG_25__SCAN_IN), .Y(n8539));
  AOI22X1 g05332(.A0(n8513), .A1(P2_ADDRESS_REG_24__SCAN_IN), .B0(P2_REIP_REG_26__SCAN_IN), .B1(n8524), .Y(n8540));
  OAI21X1 g05333(.A0(n8523), .A1(n8539), .B0(n8540), .Y(P2_U3236));
  INVX1   g05334(.A(P2_REIP_REG_24__SCAN_IN), .Y(n8542));
  AOI22X1 g05335(.A0(n8513), .A1(P2_ADDRESS_REG_23__SCAN_IN), .B0(P2_REIP_REG_25__SCAN_IN), .B1(n8524), .Y(n8543));
  OAI21X1 g05336(.A0(n8523), .A1(n8542), .B0(n8543), .Y(P2_U3235));
  INVX1   g05337(.A(P2_REIP_REG_23__SCAN_IN), .Y(n8545));
  AOI22X1 g05338(.A0(n8513), .A1(P2_ADDRESS_REG_22__SCAN_IN), .B0(P2_REIP_REG_24__SCAN_IN), .B1(n8524), .Y(n8546));
  OAI21X1 g05339(.A0(n8523), .A1(n8545), .B0(n8546), .Y(P2_U3234));
  INVX1   g05340(.A(P2_REIP_REG_22__SCAN_IN), .Y(n8548));
  AOI22X1 g05341(.A0(n8513), .A1(P2_ADDRESS_REG_21__SCAN_IN), .B0(P2_REIP_REG_23__SCAN_IN), .B1(n8524), .Y(n8549));
  OAI21X1 g05342(.A0(n8523), .A1(n8548), .B0(n8549), .Y(P2_U3233));
  INVX1   g05343(.A(P2_REIP_REG_21__SCAN_IN), .Y(n8551));
  AOI22X1 g05344(.A0(n8513), .A1(P2_ADDRESS_REG_20__SCAN_IN), .B0(P2_REIP_REG_22__SCAN_IN), .B1(n8524), .Y(n8552));
  OAI21X1 g05345(.A0(n8523), .A1(n8551), .B0(n8552), .Y(P2_U3232));
  INVX1   g05346(.A(P2_REIP_REG_20__SCAN_IN), .Y(n8554));
  AOI22X1 g05347(.A0(n8513), .A1(P2_ADDRESS_REG_19__SCAN_IN), .B0(P2_REIP_REG_21__SCAN_IN), .B1(n8524), .Y(n8555));
  OAI21X1 g05348(.A0(n8523), .A1(n8554), .B0(n8555), .Y(P2_U3231));
  INVX1   g05349(.A(P2_REIP_REG_19__SCAN_IN), .Y(n8557));
  AOI22X1 g05350(.A0(n8513), .A1(P2_ADDRESS_REG_18__SCAN_IN), .B0(P2_REIP_REG_20__SCAN_IN), .B1(n8524), .Y(n8558));
  OAI21X1 g05351(.A0(n8523), .A1(n8557), .B0(n8558), .Y(P2_U3230));
  INVX1   g05352(.A(P2_REIP_REG_18__SCAN_IN), .Y(n8560));
  AOI22X1 g05353(.A0(n8513), .A1(P2_ADDRESS_REG_17__SCAN_IN), .B0(P2_REIP_REG_19__SCAN_IN), .B1(n8524), .Y(n8561));
  OAI21X1 g05354(.A0(n8523), .A1(n8560), .B0(n8561), .Y(P2_U3229));
  INVX1   g05355(.A(P2_REIP_REG_17__SCAN_IN), .Y(n8563));
  AOI22X1 g05356(.A0(n8513), .A1(P2_ADDRESS_REG_16__SCAN_IN), .B0(P2_REIP_REG_18__SCAN_IN), .B1(n8524), .Y(n8564));
  OAI21X1 g05357(.A0(n8523), .A1(n8563), .B0(n8564), .Y(P2_U3228));
  INVX1   g05358(.A(P2_REIP_REG_16__SCAN_IN), .Y(n8566));
  AOI22X1 g05359(.A0(n8513), .A1(P2_ADDRESS_REG_15__SCAN_IN), .B0(P2_REIP_REG_17__SCAN_IN), .B1(n8524), .Y(n8567));
  OAI21X1 g05360(.A0(n8523), .A1(n8566), .B0(n8567), .Y(P2_U3227));
  INVX1   g05361(.A(P2_REIP_REG_15__SCAN_IN), .Y(n8569));
  AOI22X1 g05362(.A0(n8513), .A1(P2_ADDRESS_REG_14__SCAN_IN), .B0(P2_REIP_REG_16__SCAN_IN), .B1(n8524), .Y(n8570));
  OAI21X1 g05363(.A0(n8523), .A1(n8569), .B0(n8570), .Y(P2_U3226));
  INVX1   g05364(.A(P2_REIP_REG_14__SCAN_IN), .Y(n8572));
  AOI22X1 g05365(.A0(n8513), .A1(P2_ADDRESS_REG_13__SCAN_IN), .B0(P2_REIP_REG_15__SCAN_IN), .B1(n8524), .Y(n8573));
  OAI21X1 g05366(.A0(n8523), .A1(n8572), .B0(n8573), .Y(P2_U3225));
  INVX1   g05367(.A(P2_REIP_REG_13__SCAN_IN), .Y(n8575));
  AOI22X1 g05368(.A0(n8513), .A1(P2_ADDRESS_REG_12__SCAN_IN), .B0(P2_REIP_REG_14__SCAN_IN), .B1(n8524), .Y(n8576));
  OAI21X1 g05369(.A0(n8523), .A1(n8575), .B0(n8576), .Y(P2_U3224));
  INVX1   g05370(.A(P2_REIP_REG_12__SCAN_IN), .Y(n8578));
  AOI22X1 g05371(.A0(n8513), .A1(P2_ADDRESS_REG_11__SCAN_IN), .B0(P2_REIP_REG_13__SCAN_IN), .B1(n8524), .Y(n8579));
  OAI21X1 g05372(.A0(n8523), .A1(n8578), .B0(n8579), .Y(P2_U3223));
  INVX1   g05373(.A(P2_REIP_REG_11__SCAN_IN), .Y(n8581));
  AOI22X1 g05374(.A0(n8513), .A1(P2_ADDRESS_REG_10__SCAN_IN), .B0(P2_REIP_REG_12__SCAN_IN), .B1(n8524), .Y(n8582));
  OAI21X1 g05375(.A0(n8523), .A1(n8581), .B0(n8582), .Y(P2_U3222));
  NAND4X1 g05376(.A(n8506), .B(P2_STATE_REG_1__SCAN_IN), .C(P2_STATE_REG_2__SCAN_IN), .D(P2_REIP_REG_10__SCAN_IN), .Y(n8584));
  AOI22X1 g05377(.A0(n8513), .A1(P2_ADDRESS_REG_9__SCAN_IN), .B0(P2_REIP_REG_11__SCAN_IN), .B1(n8524), .Y(n8585));
  NAND2X1 g05378(.A(n8585), .B(n8584), .Y(P2_U3221));
  INVX1   g05379(.A(P2_REIP_REG_9__SCAN_IN), .Y(n8587));
  AOI22X1 g05380(.A0(n8513), .A1(P2_ADDRESS_REG_8__SCAN_IN), .B0(P2_REIP_REG_10__SCAN_IN), .B1(n8524), .Y(n8588));
  OAI21X1 g05381(.A0(n8523), .A1(n8587), .B0(n8588), .Y(P2_U3220));
  NAND4X1 g05382(.A(n8506), .B(P2_STATE_REG_1__SCAN_IN), .C(P2_STATE_REG_2__SCAN_IN), .D(P2_REIP_REG_8__SCAN_IN), .Y(n8590));
  AOI22X1 g05383(.A0(n8513), .A1(P2_ADDRESS_REG_7__SCAN_IN), .B0(P2_REIP_REG_9__SCAN_IN), .B1(n8524), .Y(n8591));
  NAND2X1 g05384(.A(n8591), .B(n8590), .Y(P2_U3219));
  INVX1   g05385(.A(P2_REIP_REG_7__SCAN_IN), .Y(n8593));
  AOI22X1 g05386(.A0(n8513), .A1(P2_ADDRESS_REG_6__SCAN_IN), .B0(P2_REIP_REG_8__SCAN_IN), .B1(n8524), .Y(n8594));
  OAI21X1 g05387(.A0(n8523), .A1(n8593), .B0(n8594), .Y(P2_U3218));
  NAND4X1 g05388(.A(n8506), .B(P2_STATE_REG_1__SCAN_IN), .C(P2_STATE_REG_2__SCAN_IN), .D(P2_REIP_REG_6__SCAN_IN), .Y(n8596));
  AOI22X1 g05389(.A0(n8513), .A1(P2_ADDRESS_REG_5__SCAN_IN), .B0(P2_REIP_REG_7__SCAN_IN), .B1(n8524), .Y(n8597));
  NAND2X1 g05390(.A(n8597), .B(n8596), .Y(P2_U3217));
  INVX1   g05391(.A(P2_REIP_REG_5__SCAN_IN), .Y(n8599));
  AOI22X1 g05392(.A0(n8513), .A1(P2_ADDRESS_REG_4__SCAN_IN), .B0(P2_REIP_REG_6__SCAN_IN), .B1(n8524), .Y(n8600));
  OAI21X1 g05393(.A0(n8523), .A1(n8599), .B0(n8600), .Y(P2_U3216));
  INVX1   g05394(.A(P2_REIP_REG_4__SCAN_IN), .Y(n8602));
  AOI22X1 g05395(.A0(n8513), .A1(P2_ADDRESS_REG_3__SCAN_IN), .B0(P2_REIP_REG_5__SCAN_IN), .B1(n8524), .Y(n8603));
  OAI21X1 g05396(.A0(n8523), .A1(n8602), .B0(n8603), .Y(P2_U3215));
  NAND4X1 g05397(.A(n8506), .B(P2_STATE_REG_1__SCAN_IN), .C(P2_STATE_REG_2__SCAN_IN), .D(P2_REIP_REG_3__SCAN_IN), .Y(n8605));
  AOI22X1 g05398(.A0(n8513), .A1(P2_ADDRESS_REG_2__SCAN_IN), .B0(P2_REIP_REG_4__SCAN_IN), .B1(n8524), .Y(n8606));
  NAND2X1 g05399(.A(n8606), .B(n8605), .Y(P2_U3214));
  INVX1   g05400(.A(P2_REIP_REG_2__SCAN_IN), .Y(n8608));
  AOI22X1 g05401(.A0(n8513), .A1(P2_ADDRESS_REG_1__SCAN_IN), .B0(P2_REIP_REG_3__SCAN_IN), .B1(n8524), .Y(n8609));
  OAI21X1 g05402(.A0(n8523), .A1(n8608), .B0(n8609), .Y(P2_U3213));
  INVX1   g05403(.A(P2_REIP_REG_1__SCAN_IN), .Y(n8611));
  AOI22X1 g05404(.A0(n8513), .A1(P2_ADDRESS_REG_0__SCAN_IN), .B0(P2_REIP_REG_2__SCAN_IN), .B1(n8524), .Y(n8612));
  OAI21X1 g05405(.A0(n8523), .A1(n8611), .B0(n8612), .Y(P2_U3212));
  INVX1   g05406(.A(P2_STATE_REG_2__SCAN_IN), .Y(n8614));
  INVX1   g05407(.A(READY12_REG_SCAN_IN), .Y(n8615));
  INVX1   g05408(.A(READY21_REG_SCAN_IN), .Y(n8616));
  NOR2X1  g05409(.A(P2_REQUESTPENDING_REG_SCAN_IN), .B(HOLD), .Y(n8617));
  OAI21X1 g05410(.A0(n8616), .A1(n8615), .B0(n8617), .Y(n8618));
  NOR2X1  g05411(.A(n8616), .B(n8615), .Y(n8619));
  INVX1   g05412(.A(n8619), .Y(n8620));
  INVX1   g05413(.A(P2_REQUESTPENDING_REG_SCAN_IN), .Y(n8621));
  NOR2X1  g05414(.A(n8621), .B(HOLD), .Y(n8622));
  AOI21X1 g05415(.A0(n8622), .A1(n8620), .B0(n8508), .Y(n8623));
  NAND2X1 g05416(.A(P2_STATE_REG_0__SCAN_IN), .B(HOLD), .Y(n8624));
  OAI21X1 g05417(.A0(P2_STATE_REG_0__SCAN_IN), .A1(NA), .B0(n8624), .Y(n8625));
  AOI21X1 g05418(.A0(n8623), .A1(n8618), .B0(n8625), .Y(n8626));
  NAND3X1 g05419(.A(P2_STATE_REG_1__SCAN_IN), .B(READY21_REG_SCAN_IN), .C(READY12_REG_SCAN_IN), .Y(n8627));
  NOR2X1  g05420(.A(P2_STATE_REG_1__SCAN_IN), .B(P2_STATE_REG_2__SCAN_IN), .Y(n8628));
  NAND3X1 g05421(.A(n8628), .B(n8621), .C(HOLD), .Y(n8629));
  OAI21X1 g05422(.A0(n8627), .A1(n8617), .B0(n8629), .Y(n8630));
  NOR3X1  g05423(.A(n8508), .B(P2_STATE_REG_2__SCAN_IN), .C(n3419), .Y(n8631));
  NOR2X1  g05424(.A(n8631), .B(n8506), .Y(n8632));
  AOI22X1 g05425(.A0(n8630), .A1(n8632), .B0(n8512), .B1(P2_STATE_REG_2__SCAN_IN), .Y(n8633));
  OAI21X1 g05426(.A0(n8626), .A1(n8614), .B0(n8633), .Y(P2_U3211));
  NOR3X1  g05427(.A(n8621), .B(n8506), .C(HOLD), .Y(n8635));
  NAND3X1 g05428(.A(P2_REQUESTPENDING_REG_SCAN_IN), .B(P2_STATE_REG_0__SCAN_IN), .C(n8614), .Y(n8636));
  OAI21X1 g05429(.A0(P2_STATE_REG_0__SCAN_IN), .A1(n8614), .B0(n8636), .Y(n8637));
  OAI21X1 g05430(.A0(n8637), .A1(n8635), .B0(n8508), .Y(n8638));
  AOI21X1 g05431(.A0(READY21_REG_SCAN_IN), .A1(READY12_REG_SCAN_IN), .B0(n3428), .Y(n8639));
  OAI21X1 g05432(.A0(n8639), .A1(n8506), .B0(P2_STATE_REG_2__SCAN_IN), .Y(n8640));
  NAND3X1 g05433(.A(n8640), .B(n8618), .C(P2_STATE_REG_1__SCAN_IN), .Y(n8641));
  OAI21X1 g05434(.A0(n8619), .A1(n8614), .B0(n8512), .Y(n8642));
  NAND3X1 g05435(.A(n8642), .B(n8641), .C(n8638), .Y(P2_U3210));
  NAND2X1 g05436(.A(P2_REQUESTPENDING_REG_SCAN_IN), .B(P2_STATE_REG_0__SCAN_IN), .Y(n8644));
  OAI21X1 g05437(.A0(n8644), .A1(n8623), .B0(n8614), .Y(n8645));
  OAI22X1 g05438(.A0(P2_STATE_REG_0__SCAN_IN), .A1(n3419), .B0(n8614), .B1(n8622), .Y(n8646));
  NOR3X1  g05439(.A(n8622), .B(n8506), .C(n8614), .Y(n8647));
  AOI21X1 g05440(.A0(n8646), .A1(n8508), .B0(n8647), .Y(n8648));
  NAND2X1 g05441(.A(n8648), .B(n8645), .Y(P2_U3209));
  OAI21X1 g05442(.A0(P2_STATE_REG_1__SCAN_IN), .A1(P2_STATE_REG_2__SCAN_IN), .B0(n3439), .Y(n8650));
  NOR3X1  g05443(.A(n8506), .B(n8508), .C(P2_STATE_REG_2__SCAN_IN), .Y(n8651));
  AOI21X1 g05444(.A0(n8506), .A1(n8508), .B0(n8651), .Y(n8652));
  NAND2X1 g05445(.A(n8652), .B(P2_DATAWIDTH_REG_0__SCAN_IN), .Y(n8653));
  OAI21X1 g05446(.A0(n8652), .A1(n8650), .B0(n8653), .Y(P2_U3591));
  INVX1   g05447(.A(P2_DATAWIDTH_REG_1__SCAN_IN), .Y(n8655));
  INVX1   g05448(.A(n8652), .Y(n8656));
  NAND2X1 g05449(.A(n8656), .B(n8650), .Y(n8657));
  OAI21X1 g05450(.A0(n8656), .A1(n8655), .B0(n8657), .Y(P2_U3592));
  INVX1   g05451(.A(P2_DATAWIDTH_REG_2__SCAN_IN), .Y(n8659));
  NOR2X1  g05452(.A(n8656), .B(n8659), .Y(P2_U3208));
  INVX1   g05453(.A(P2_DATAWIDTH_REG_3__SCAN_IN), .Y(n8661));
  NOR2X1  g05454(.A(n8656), .B(n8661), .Y(P2_U3207));
  INVX1   g05455(.A(P2_DATAWIDTH_REG_4__SCAN_IN), .Y(n8663));
  NOR2X1  g05456(.A(n8656), .B(n8663), .Y(P2_U3206));
  INVX1   g05457(.A(P2_DATAWIDTH_REG_5__SCAN_IN), .Y(n8665));
  NOR2X1  g05458(.A(n8656), .B(n8665), .Y(P2_U3205));
  INVX1   g05459(.A(P2_DATAWIDTH_REG_6__SCAN_IN), .Y(n8667));
  NOR2X1  g05460(.A(n8656), .B(n8667), .Y(P2_U3204));
  INVX1   g05461(.A(P2_DATAWIDTH_REG_7__SCAN_IN), .Y(n8669));
  NOR2X1  g05462(.A(n8656), .B(n8669), .Y(P2_U3203));
  INVX1   g05463(.A(P2_DATAWIDTH_REG_8__SCAN_IN), .Y(n8671));
  NOR2X1  g05464(.A(n8656), .B(n8671), .Y(P2_U3202));
  INVX1   g05465(.A(P2_DATAWIDTH_REG_9__SCAN_IN), .Y(n8673));
  NOR2X1  g05466(.A(n8656), .B(n8673), .Y(P2_U3201));
  INVX1   g05467(.A(P2_DATAWIDTH_REG_10__SCAN_IN), .Y(n8675));
  NOR2X1  g05468(.A(n8656), .B(n8675), .Y(P2_U3200));
  INVX1   g05469(.A(P2_DATAWIDTH_REG_11__SCAN_IN), .Y(n8677));
  NOR2X1  g05470(.A(n8656), .B(n8677), .Y(P2_U3199));
  INVX1   g05471(.A(P2_DATAWIDTH_REG_12__SCAN_IN), .Y(n8679));
  NOR2X1  g05472(.A(n8656), .B(n8679), .Y(P2_U3198));
  INVX1   g05473(.A(P2_DATAWIDTH_REG_13__SCAN_IN), .Y(n8681));
  NOR2X1  g05474(.A(n8656), .B(n8681), .Y(P2_U3197));
  INVX1   g05475(.A(P2_DATAWIDTH_REG_14__SCAN_IN), .Y(n8683));
  NOR2X1  g05476(.A(n8656), .B(n8683), .Y(P2_U3196));
  INVX1   g05477(.A(P2_DATAWIDTH_REG_15__SCAN_IN), .Y(n8685));
  NOR2X1  g05478(.A(n8656), .B(n8685), .Y(P2_U3195));
  INVX1   g05479(.A(P2_DATAWIDTH_REG_16__SCAN_IN), .Y(n8687));
  NOR2X1  g05480(.A(n8656), .B(n8687), .Y(P2_U3194));
  INVX1   g05481(.A(P2_DATAWIDTH_REG_17__SCAN_IN), .Y(n8689));
  NOR2X1  g05482(.A(n8656), .B(n8689), .Y(P2_U3193));
  INVX1   g05483(.A(P2_DATAWIDTH_REG_18__SCAN_IN), .Y(n8691));
  NOR2X1  g05484(.A(n8656), .B(n8691), .Y(P2_U3192));
  INVX1   g05485(.A(P2_DATAWIDTH_REG_19__SCAN_IN), .Y(n8693));
  NOR2X1  g05486(.A(n8656), .B(n8693), .Y(P2_U3191));
  INVX1   g05487(.A(P2_DATAWIDTH_REG_20__SCAN_IN), .Y(n8695));
  NOR2X1  g05488(.A(n8656), .B(n8695), .Y(P2_U3190));
  INVX1   g05489(.A(P2_DATAWIDTH_REG_21__SCAN_IN), .Y(n8697));
  NOR2X1  g05490(.A(n8656), .B(n8697), .Y(P2_U3189));
  INVX1   g05491(.A(P2_DATAWIDTH_REG_22__SCAN_IN), .Y(n8699));
  NOR2X1  g05492(.A(n8656), .B(n8699), .Y(P2_U3188));
  INVX1   g05493(.A(P2_DATAWIDTH_REG_23__SCAN_IN), .Y(n8701));
  NOR2X1  g05494(.A(n8656), .B(n8701), .Y(P2_U3187));
  INVX1   g05495(.A(P2_DATAWIDTH_REG_24__SCAN_IN), .Y(n8703));
  NOR2X1  g05496(.A(n8656), .B(n8703), .Y(P2_U3186));
  INVX1   g05497(.A(P2_DATAWIDTH_REG_25__SCAN_IN), .Y(n8705));
  NOR2X1  g05498(.A(n8656), .B(n8705), .Y(P2_U3185));
  INVX1   g05499(.A(P2_DATAWIDTH_REG_26__SCAN_IN), .Y(n8707));
  NOR2X1  g05500(.A(n8656), .B(n8707), .Y(P2_U3184));
  INVX1   g05501(.A(P2_DATAWIDTH_REG_27__SCAN_IN), .Y(n8709));
  NOR2X1  g05502(.A(n8656), .B(n8709), .Y(P2_U3183));
  INVX1   g05503(.A(P2_DATAWIDTH_REG_28__SCAN_IN), .Y(n8711));
  NOR2X1  g05504(.A(n8656), .B(n8711), .Y(P2_U3182));
  INVX1   g05505(.A(P2_DATAWIDTH_REG_29__SCAN_IN), .Y(n8713));
  NOR2X1  g05506(.A(n8656), .B(n8713), .Y(P2_U3181));
  INVX1   g05507(.A(P2_DATAWIDTH_REG_30__SCAN_IN), .Y(n8715));
  NOR2X1  g05508(.A(n8656), .B(n8715), .Y(P2_U3180));
  INVX1   g05509(.A(P2_DATAWIDTH_REG_31__SCAN_IN), .Y(n8717));
  NOR2X1  g05510(.A(n8656), .B(n8717), .Y(P2_U3179));
  INVX1   g05511(.A(P2_STATE2_REG_3__SCAN_IN), .Y(n8719));
  INVX1   g05512(.A(P2_STATE2_REG_0__SCAN_IN), .Y(n8720));
  INVX1   g05513(.A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n8721));
  NAND3X1 g05514(.A(n8721), .B(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Y(n8722));
  NOR2X1  g05515(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_6__4__SCAN_IN), .Y(n8723));
  INVX1   g05516(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n8724));
  NOR2X1  g05517(.A(n8724), .B(P2_INSTQUEUE_REG_14__4__SCAN_IN), .Y(n8725));
  NOR3X1  g05518(.A(n8725), .B(n8723), .C(n8722), .Y(n8726));
  INVX1   g05519(.A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Y(n8727));
  NAND3X1 g05520(.A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C(n8727), .Y(n8728));
  NOR2X1  g05521(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_3__4__SCAN_IN), .Y(n8729));
  NOR2X1  g05522(.A(n8724), .B(P2_INSTQUEUE_REG_11__4__SCAN_IN), .Y(n8730));
  NOR3X1  g05523(.A(n8730), .B(n8729), .C(n8728), .Y(n8731));
  INVX1   g05524(.A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Y(n8732));
  NAND3X1 g05525(.A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(n8732), .C(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Y(n8733));
  NOR2X1  g05526(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_5__4__SCAN_IN), .Y(n8734));
  NOR2X1  g05527(.A(n8724), .B(P2_INSTQUEUE_REG_13__4__SCAN_IN), .Y(n8735));
  NOR3X1  g05528(.A(n8735), .B(n8734), .C(n8733), .Y(n8736));
  NAND3X1 g05529(.A(n8721), .B(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C(n8727), .Y(n8737));
  NOR2X1  g05530(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_2__4__SCAN_IN), .Y(n8738));
  NOR2X1  g05531(.A(n8724), .B(P2_INSTQUEUE_REG_10__4__SCAN_IN), .Y(n8739));
  NOR3X1  g05532(.A(n8739), .B(n8738), .C(n8737), .Y(n8740));
  NOR4X1  g05533(.A(n8736), .B(n8731), .C(n8726), .D(n8740), .Y(n8741));
  NAND3X1 g05534(.A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Y(n8742));
  NOR2X1  g05535(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_7__4__SCAN_IN), .Y(n8743));
  NOR2X1  g05536(.A(n8724), .B(P2_INSTQUEUE_REG_15__4__SCAN_IN), .Y(n8744));
  NOR3X1  g05537(.A(n8744), .B(n8743), .C(n8742), .Y(n8745));
  NAND3X1 g05538(.A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(n8732), .C(n8727), .Y(n8746));
  NOR2X1  g05539(.A(n8724), .B(P2_INSTQUEUE_REG_9__4__SCAN_IN), .Y(n8747));
  NOR2X1  g05540(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_1__4__SCAN_IN), .Y(n8748));
  NOR3X1  g05541(.A(n8748), .B(n8747), .C(n8746), .Y(n8749));
  NAND3X1 g05542(.A(n8721), .B(n8732), .C(n8727), .Y(n8750));
  NOR2X1  g05543(.A(n8724), .B(P2_INSTQUEUE_REG_8__4__SCAN_IN), .Y(n8751));
  NOR2X1  g05544(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_0__4__SCAN_IN), .Y(n8752));
  NOR3X1  g05545(.A(n8752), .B(n8751), .C(n8750), .Y(n8753));
  NAND3X1 g05546(.A(n8721), .B(n8732), .C(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Y(n8754));
  NOR2X1  g05547(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_4__4__SCAN_IN), .Y(n8755));
  NOR2X1  g05548(.A(n8724), .B(P2_INSTQUEUE_REG_12__4__SCAN_IN), .Y(n8756));
  NOR3X1  g05549(.A(n8756), .B(n8755), .C(n8754), .Y(n8757));
  NOR4X1  g05550(.A(n8753), .B(n8749), .C(n8745), .D(n8757), .Y(n8758));
  NOR3X1  g05551(.A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(n8732), .C(n8727), .Y(n8759));
  NOR3X1  g05552(.A(n8721), .B(n8732), .C(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Y(n8760));
  INVX1   g05553(.A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .Y(n8761));
  NOR2X1  g05554(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_6__6__SCAN_IN), .Y(n8762));
  AOI21X1 g05555(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8761), .B0(n8762), .Y(n8763));
  INVX1   g05556(.A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .Y(n8764));
  NOR2X1  g05557(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_3__6__SCAN_IN), .Y(n8765));
  AOI21X1 g05558(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8764), .B0(n8765), .Y(n8766));
  AOI22X1 g05559(.A0(n8763), .A1(n8759), .B0(n8760), .B1(n8766), .Y(n8767));
  NOR3X1  g05560(.A(n8721), .B(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C(n8727), .Y(n8768));
  NOR3X1  g05561(.A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(n8732), .C(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Y(n8769));
  INVX1   g05562(.A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .Y(n8770));
  NOR2X1  g05563(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_5__6__SCAN_IN), .Y(n8771));
  AOI21X1 g05564(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8770), .B0(n8771), .Y(n8772));
  INVX1   g05565(.A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .Y(n8773));
  NOR2X1  g05566(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_2__6__SCAN_IN), .Y(n8774));
  AOI21X1 g05567(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8773), .B0(n8774), .Y(n8775));
  AOI22X1 g05568(.A0(n8772), .A1(n8768), .B0(n8769), .B1(n8775), .Y(n8776));
  NAND2X1 g05569(.A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Y(n8777));
  NOR2X1  g05570(.A(n8777), .B(n8721), .Y(n8778));
  NOR3X1  g05571(.A(n8721), .B(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Y(n8779));
  INVX1   g05572(.A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .Y(n8780));
  NOR2X1  g05573(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_7__6__SCAN_IN), .Y(n8781));
  AOI21X1 g05574(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8780), .B0(n8781), .Y(n8782));
  INVX1   g05575(.A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .Y(n8783));
  NOR2X1  g05576(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_1__6__SCAN_IN), .Y(n8784));
  AOI21X1 g05577(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8783), .B0(n8784), .Y(n8785));
  AOI22X1 g05578(.A0(n8782), .A1(n8778), .B0(n8779), .B1(n8785), .Y(n8786));
  NOR3X1  g05579(.A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Y(n8787));
  NOR3X1  g05580(.A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C(n8727), .Y(n8788));
  INVX1   g05581(.A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .Y(n8789));
  NOR2X1  g05582(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_0__6__SCAN_IN), .Y(n8790));
  AOI21X1 g05583(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8789), .B0(n8790), .Y(n8791));
  INVX1   g05584(.A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .Y(n8792));
  NOR2X1  g05585(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_4__6__SCAN_IN), .Y(n8793));
  AOI21X1 g05586(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8792), .B0(n8793), .Y(n8794));
  AOI22X1 g05587(.A0(n8791), .A1(n8787), .B0(n8788), .B1(n8794), .Y(n8795));
  NAND4X1 g05588(.A(n8786), .B(n8776), .C(n8767), .D(n8795), .Y(n8796));
  INVX1   g05589(.A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .Y(n8797));
  NOR2X1  g05590(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_6__5__SCAN_IN), .Y(n8798));
  AOI21X1 g05591(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8797), .B0(n8798), .Y(n8799));
  INVX1   g05592(.A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .Y(n8800));
  NOR2X1  g05593(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_3__5__SCAN_IN), .Y(n8801));
  AOI21X1 g05594(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8800), .B0(n8801), .Y(n8802));
  AOI22X1 g05595(.A0(n8799), .A1(n8759), .B0(n8760), .B1(n8802), .Y(n8803));
  INVX1   g05596(.A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .Y(n8804));
  NOR2X1  g05597(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_5__5__SCAN_IN), .Y(n8805));
  AOI21X1 g05598(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8804), .B0(n8805), .Y(n8806));
  INVX1   g05599(.A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .Y(n8807));
  NOR2X1  g05600(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_2__5__SCAN_IN), .Y(n8808));
  AOI21X1 g05601(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8807), .B0(n8808), .Y(n8809));
  AOI22X1 g05602(.A0(n8806), .A1(n8768), .B0(n8769), .B1(n8809), .Y(n8810));
  INVX1   g05603(.A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .Y(n8811));
  NOR2X1  g05604(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_7__5__SCAN_IN), .Y(n8812));
  AOI21X1 g05605(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8811), .B0(n8812), .Y(n8813));
  INVX1   g05606(.A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .Y(n8814));
  NOR2X1  g05607(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_1__5__SCAN_IN), .Y(n8815));
  AOI21X1 g05608(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8814), .B0(n8815), .Y(n8816));
  AOI22X1 g05609(.A0(n8813), .A1(n8778), .B0(n8779), .B1(n8816), .Y(n8817));
  INVX1   g05610(.A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .Y(n8818));
  NOR2X1  g05611(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .Y(n8819));
  AOI21X1 g05612(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8818), .B0(n8819), .Y(n8820));
  INVX1   g05613(.A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .Y(n8821));
  NOR2X1  g05614(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_4__5__SCAN_IN), .Y(n8822));
  AOI21X1 g05615(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8821), .B0(n8822), .Y(n8823));
  AOI22X1 g05616(.A0(n8820), .A1(n8787), .B0(n8788), .B1(n8823), .Y(n8824));
  NAND4X1 g05617(.A(n8817), .B(n8810), .C(n8803), .D(n8824), .Y(n8825));
  NAND4X1 g05618(.A(n8796), .B(n8758), .C(n8741), .D(n8825), .Y(n8826));
  INVX1   g05619(.A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .Y(n8827));
  NOR2X1  g05620(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_6__2__SCAN_IN), .Y(n8828));
  AOI21X1 g05621(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8827), .B0(n8828), .Y(n8829));
  INVX1   g05622(.A(P2_INSTQUEUE_REG_11__2__SCAN_IN), .Y(n8830));
  NOR2X1  g05623(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_3__2__SCAN_IN), .Y(n8831));
  AOI21X1 g05624(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8830), .B0(n8831), .Y(n8832));
  AOI22X1 g05625(.A0(n8829), .A1(n8759), .B0(n8760), .B1(n8832), .Y(n8833));
  INVX1   g05626(.A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .Y(n8834));
  NOR2X1  g05627(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_5__2__SCAN_IN), .Y(n8835));
  AOI21X1 g05628(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8834), .B0(n8835), .Y(n8836));
  INVX1   g05629(.A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .Y(n8837));
  NOR2X1  g05630(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_2__2__SCAN_IN), .Y(n8838));
  AOI21X1 g05631(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8837), .B0(n8838), .Y(n8839));
  AOI22X1 g05632(.A0(n8836), .A1(n8768), .B0(n8769), .B1(n8839), .Y(n8840));
  INVX1   g05633(.A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .Y(n8841));
  NOR2X1  g05634(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_7__2__SCAN_IN), .Y(n8842));
  AOI21X1 g05635(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8841), .B0(n8842), .Y(n8843));
  INVX1   g05636(.A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .Y(n8844));
  NOR2X1  g05637(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_1__2__SCAN_IN), .Y(n8845));
  AOI21X1 g05638(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8844), .B0(n8845), .Y(n8846));
  AOI22X1 g05639(.A0(n8843), .A1(n8778), .B0(n8779), .B1(n8846), .Y(n8847));
  INVX1   g05640(.A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .Y(n8848));
  NOR2X1  g05641(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_0__2__SCAN_IN), .Y(n8849));
  AOI21X1 g05642(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8848), .B0(n8849), .Y(n8850));
  INVX1   g05643(.A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .Y(n8851));
  NOR2X1  g05644(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_4__2__SCAN_IN), .Y(n8852));
  AOI21X1 g05645(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8851), .B0(n8852), .Y(n8853));
  AOI22X1 g05646(.A0(n8850), .A1(n8787), .B0(n8788), .B1(n8853), .Y(n8854));
  NAND4X1 g05647(.A(n8847), .B(n8840), .C(n8833), .D(n8854), .Y(n8855));
  INVX1   g05648(.A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .Y(n8856));
  NOR2X1  g05649(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_6__7__SCAN_IN), .Y(n8857));
  AOI21X1 g05650(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8856), .B0(n8857), .Y(n8858));
  INVX1   g05651(.A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .Y(n8859));
  NOR2X1  g05652(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_3__7__SCAN_IN), .Y(n8860));
  AOI21X1 g05653(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8859), .B0(n8860), .Y(n8861));
  AOI22X1 g05654(.A0(n8858), .A1(n8759), .B0(n8760), .B1(n8861), .Y(n8862));
  INVX1   g05655(.A(P2_INSTQUEUE_REG_13__7__SCAN_IN), .Y(n8863));
  NOR2X1  g05656(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_5__7__SCAN_IN), .Y(n8864));
  AOI21X1 g05657(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8863), .B0(n8864), .Y(n8865));
  INVX1   g05658(.A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .Y(n8866));
  NOR2X1  g05659(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_2__7__SCAN_IN), .Y(n8867));
  AOI21X1 g05660(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8866), .B0(n8867), .Y(n8868));
  AOI22X1 g05661(.A0(n8865), .A1(n8768), .B0(n8769), .B1(n8868), .Y(n8869));
  INVX1   g05662(.A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .Y(n8870));
  NOR2X1  g05663(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_7__7__SCAN_IN), .Y(n8871));
  AOI21X1 g05664(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8870), .B0(n8871), .Y(n8872));
  INVX1   g05665(.A(P2_INSTQUEUE_REG_9__7__SCAN_IN), .Y(n8873));
  NOR2X1  g05666(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_1__7__SCAN_IN), .Y(n8874));
  AOI21X1 g05667(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8873), .B0(n8874), .Y(n8875));
  AOI22X1 g05668(.A0(n8872), .A1(n8778), .B0(n8779), .B1(n8875), .Y(n8876));
  INVX1   g05669(.A(P2_INSTQUEUE_REG_8__7__SCAN_IN), .Y(n8877));
  NOR2X1  g05670(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .Y(n8878));
  AOI21X1 g05671(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8877), .B0(n8878), .Y(n8879));
  INVX1   g05672(.A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .Y(n8880));
  NOR2X1  g05673(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_4__7__SCAN_IN), .Y(n8881));
  AOI21X1 g05674(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8880), .B0(n8881), .Y(n8882));
  AOI22X1 g05675(.A0(n8879), .A1(n8787), .B0(n8788), .B1(n8882), .Y(n8883));
  NAND4X1 g05676(.A(n8876), .B(n8869), .C(n8862), .D(n8883), .Y(n8884));
  INVX1   g05677(.A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .Y(n8885));
  NOR2X1  g05678(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_6__3__SCAN_IN), .Y(n8886));
  AOI21X1 g05679(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8885), .B0(n8886), .Y(n8887));
  INVX1   g05680(.A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .Y(n8888));
  NOR2X1  g05681(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_3__3__SCAN_IN), .Y(n8889));
  AOI21X1 g05682(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8888), .B0(n8889), .Y(n8890));
  AOI22X1 g05683(.A0(n8887), .A1(n8759), .B0(n8760), .B1(n8890), .Y(n8891));
  INVX1   g05684(.A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .Y(n8892));
  NOR2X1  g05685(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_5__3__SCAN_IN), .Y(n8893));
  AOI21X1 g05686(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8892), .B0(n8893), .Y(n8894));
  INVX1   g05687(.A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .Y(n8895));
  NOR2X1  g05688(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_2__3__SCAN_IN), .Y(n8896));
  AOI21X1 g05689(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8895), .B0(n8896), .Y(n8897));
  AOI22X1 g05690(.A0(n8894), .A1(n8768), .B0(n8769), .B1(n8897), .Y(n8898));
  INVX1   g05691(.A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .Y(n8899));
  NOR2X1  g05692(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_7__3__SCAN_IN), .Y(n8900));
  AOI21X1 g05693(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8899), .B0(n8900), .Y(n8901));
  INVX1   g05694(.A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .Y(n8902));
  NOR2X1  g05695(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_1__3__SCAN_IN), .Y(n8903));
  AOI21X1 g05696(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8902), .B0(n8903), .Y(n8904));
  AOI22X1 g05697(.A0(n8901), .A1(n8778), .B0(n8779), .B1(n8904), .Y(n8905));
  INVX1   g05698(.A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .Y(n8906));
  NOR2X1  g05699(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_0__3__SCAN_IN), .Y(n8907));
  AOI21X1 g05700(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8906), .B0(n8907), .Y(n8908));
  INVX1   g05701(.A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .Y(n8909));
  NOR2X1  g05702(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_4__3__SCAN_IN), .Y(n8910));
  AOI21X1 g05703(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8909), .B0(n8910), .Y(n8911));
  AOI22X1 g05704(.A0(n8908), .A1(n8787), .B0(n8788), .B1(n8911), .Y(n8912));
  NAND4X1 g05705(.A(n8905), .B(n8898), .C(n8891), .D(n8912), .Y(n8913));
  NAND2X1 g05706(.A(n8913), .B(n8884), .Y(n8914));
  NOR3X1  g05707(.A(n8914), .B(n8855), .C(n8826), .Y(n8915));
  INVX1   g05708(.A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .Y(n8916));
  NOR2X1  g05709(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_6__0__SCAN_IN), .Y(n8917));
  AOI21X1 g05710(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8916), .B0(n8917), .Y(n8918));
  INVX1   g05711(.A(P2_INSTQUEUE_REG_11__0__SCAN_IN), .Y(n8919));
  NOR2X1  g05712(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_3__0__SCAN_IN), .Y(n8920));
  AOI21X1 g05713(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8919), .B0(n8920), .Y(n8921));
  AOI22X1 g05714(.A0(n8918), .A1(n8759), .B0(n8760), .B1(n8921), .Y(n8922));
  INVX1   g05715(.A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .Y(n8923));
  NOR2X1  g05716(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_5__0__SCAN_IN), .Y(n8924));
  AOI21X1 g05717(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8923), .B0(n8924), .Y(n8925));
  INVX1   g05718(.A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .Y(n8926));
  NOR2X1  g05719(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_2__0__SCAN_IN), .Y(n8927));
  AOI21X1 g05720(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8926), .B0(n8927), .Y(n8928));
  AOI22X1 g05721(.A0(n8925), .A1(n8768), .B0(n8769), .B1(n8928), .Y(n8929));
  NAND2X1 g05722(.A(n8929), .B(n8922), .Y(n8930));
  INVX1   g05723(.A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .Y(n8931));
  NOR2X1  g05724(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_7__0__SCAN_IN), .Y(n8932));
  AOI21X1 g05725(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8931), .B0(n8932), .Y(n8933));
  INVX1   g05726(.A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .Y(n8934));
  NOR2X1  g05727(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_1__0__SCAN_IN), .Y(n8935));
  AOI21X1 g05728(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8934), .B0(n8935), .Y(n8936));
  AOI22X1 g05729(.A0(n8933), .A1(n8778), .B0(n8779), .B1(n8936), .Y(n8937));
  INVX1   g05730(.A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .Y(n8938));
  NOR2X1  g05731(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_0__0__SCAN_IN), .Y(n8939));
  AOI21X1 g05732(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8938), .B0(n8939), .Y(n8940));
  INVX1   g05733(.A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .Y(n8941));
  NOR2X1  g05734(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_4__0__SCAN_IN), .Y(n8942));
  AOI21X1 g05735(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8941), .B0(n8942), .Y(n8943));
  AOI22X1 g05736(.A0(n8940), .A1(n8787), .B0(n8788), .B1(n8943), .Y(n8944));
  NAND2X1 g05737(.A(n8944), .B(n8937), .Y(n8945));
  NOR2X1  g05738(.A(n8945), .B(n8930), .Y(n8946));
  INVX1   g05739(.A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .Y(n8947));
  NOR2X1  g05740(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_6__1__SCAN_IN), .Y(n8948));
  AOI21X1 g05741(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8947), .B0(n8948), .Y(n8949));
  INVX1   g05742(.A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .Y(n8950));
  NOR2X1  g05743(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_3__1__SCAN_IN), .Y(n8951));
  AOI21X1 g05744(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8950), .B0(n8951), .Y(n8952));
  AOI22X1 g05745(.A0(n8949), .A1(n8759), .B0(n8760), .B1(n8952), .Y(n8953));
  INVX1   g05746(.A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .Y(n8954));
  NOR2X1  g05747(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_5__1__SCAN_IN), .Y(n8955));
  AOI21X1 g05748(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8954), .B0(n8955), .Y(n8956));
  INVX1   g05749(.A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .Y(n8957));
  NOR2X1  g05750(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_2__1__SCAN_IN), .Y(n8958));
  AOI21X1 g05751(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8957), .B0(n8958), .Y(n8959));
  AOI22X1 g05752(.A0(n8956), .A1(n8768), .B0(n8769), .B1(n8959), .Y(n8960));
  INVX1   g05753(.A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .Y(n8961));
  NOR2X1  g05754(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_7__1__SCAN_IN), .Y(n8962));
  AOI21X1 g05755(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8961), .B0(n8962), .Y(n8963));
  INVX1   g05756(.A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .Y(n8964));
  NOR2X1  g05757(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_1__1__SCAN_IN), .Y(n8965));
  AOI21X1 g05758(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8964), .B0(n8965), .Y(n8966));
  AOI22X1 g05759(.A0(n8963), .A1(n8778), .B0(n8779), .B1(n8966), .Y(n8967));
  INVX1   g05760(.A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .Y(n8968));
  NOR2X1  g05761(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_0__1__SCAN_IN), .Y(n8969));
  AOI21X1 g05762(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8968), .B0(n8969), .Y(n8970));
  INVX1   g05763(.A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .Y(n8971));
  NOR2X1  g05764(.A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P2_INSTQUEUE_REG_4__1__SCAN_IN), .Y(n8972));
  AOI21X1 g05765(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n8971), .B0(n8972), .Y(n8973));
  AOI22X1 g05766(.A0(n8970), .A1(n8787), .B0(n8788), .B1(n8973), .Y(n8974));
  NAND4X1 g05767(.A(n8967), .B(n8960), .C(n8953), .D(n8974), .Y(n8975));
  NOR2X1  g05768(.A(n8975), .B(n8946), .Y(n8976));
  INVX1   g05769(.A(n8976), .Y(n8977));
  NAND4X1 g05770(.A(n8937), .B(n8929), .C(n8922), .D(n8944), .Y(n8978));
  NAND2X1 g05771(.A(n8975), .B(n8978), .Y(n8979));
  NOR4X1  g05772(.A(n8732), .B(n8727), .C(n8724), .D(n8721), .Y(n8980));
  NOR4X1  g05773(.A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .D(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n8981));
  AOI22X1 g05774(.A0(n8980), .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B0(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(n8981), .Y(n8982));
  NOR4X1  g05775(.A(n8732), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .D(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n8983));
  NOR4X1  g05776(.A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .D(n8721), .Y(n8984));
  AOI22X1 g05777(.A0(n8983), .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B0(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(n8984), .Y(n8985));
  NOR4X1  g05778(.A(n8732), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .D(n8721), .Y(n8986));
  NOR4X1  g05779(.A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n8727), .C(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .D(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n8987));
  AOI22X1 g05780(.A0(n8986), .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B0(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(n8987), .Y(n8988));
  NOR4X1  g05781(.A(n8732), .B(n8727), .C(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .D(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n8989));
  NOR4X1  g05782(.A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n8727), .C(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .D(n8721), .Y(n8990));
  AOI22X1 g05783(.A0(n8989), .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B0(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(n8990), .Y(n8991));
  NAND4X1 g05784(.A(n8988), .B(n8985), .C(n8982), .D(n8991), .Y(n8992));
  NOR4X1  g05785(.A(n8732), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(n8724), .D(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n8993));
  NOR4X1  g05786(.A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(n8724), .D(n8721), .Y(n8994));
  AOI22X1 g05787(.A0(n8993), .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B0(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(n8994), .Y(n8995));
  NOR4X1  g05788(.A(n8732), .B(n8727), .C(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .D(n8721), .Y(n8996));
  NOR4X1  g05789(.A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(n8724), .D(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n8997));
  AOI22X1 g05790(.A0(n8996), .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B0(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(n8997), .Y(n8998));
  NOR4X1  g05791(.A(n8732), .B(n8727), .C(n8724), .D(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n8999));
  NOR4X1  g05792(.A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n8727), .C(n8724), .D(n8721), .Y(n9000));
  AOI22X1 g05793(.A0(n8999), .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B0(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(n9000), .Y(n9001));
  NOR4X1  g05794(.A(n8732), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(n8724), .D(n8721), .Y(n9002));
  NOR4X1  g05795(.A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n8727), .C(n8724), .D(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n9003));
  AOI22X1 g05796(.A0(n9002), .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B0(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(n9003), .Y(n9004));
  NAND4X1 g05797(.A(n9001), .B(n8998), .C(n8995), .D(n9004), .Y(n9005));
  NOR3X1  g05798(.A(n9005), .B(n8992), .C(n8979), .Y(n9006));
  INVX1   g05799(.A(n8979), .Y(n9007));
  AOI22X1 g05800(.A0(n8980), .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B0(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(n8981), .Y(n9008));
  AOI22X1 g05801(.A0(n8983), .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B0(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(n8984), .Y(n9009));
  AOI22X1 g05802(.A0(n8986), .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B0(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(n8987), .Y(n9010));
  AOI22X1 g05803(.A0(n8989), .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B0(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(n8990), .Y(n9011));
  NAND4X1 g05804(.A(n9010), .B(n9009), .C(n9008), .D(n9011), .Y(n9012));
  AOI22X1 g05805(.A0(n8993), .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B0(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(n8994), .Y(n9013));
  AOI22X1 g05806(.A0(n8996), .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B0(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(n8997), .Y(n9014));
  AOI22X1 g05807(.A0(n8999), .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B0(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(n9000), .Y(n9015));
  AOI22X1 g05808(.A0(n9002), .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B0(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(n9003), .Y(n9016));
  NAND4X1 g05809(.A(n9015), .B(n9014), .C(n9013), .D(n9016), .Y(n9017));
  NOR2X1  g05810(.A(n9017), .B(n9012), .Y(n9018));
  INVX1   g05811(.A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .Y(n9019));
  NAND2X1 g05812(.A(n8960), .B(n8953), .Y(n9020));
  NAND2X1 g05813(.A(n8974), .B(n8967), .Y(n9021));
  NOR2X1  g05814(.A(n9021), .B(n9020), .Y(n9022));
  AOI22X1 g05815(.A0(n8980), .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B0(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(n8981), .Y(n9024));
  AOI22X1 g05816(.A0(n8983), .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B0(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(n8984), .Y(n9025));
  AOI22X1 g05817(.A0(n8986), .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B0(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(n8987), .Y(n9026));
  AOI22X1 g05818(.A0(n8989), .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B0(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(n8990), .Y(n9027));
  NAND4X1 g05819(.A(n9026), .B(n9025), .C(n9024), .D(n9027), .Y(n9028));
  AOI22X1 g05820(.A0(n8993), .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B0(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(n8994), .Y(n9029));
  AOI22X1 g05821(.A0(n8996), .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B0(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(n8997), .Y(n9030));
  AOI22X1 g05822(.A0(n8999), .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B0(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(n9000), .Y(n9031));
  AOI22X1 g05823(.A0(n9002), .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B0(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(n9003), .Y(n9032));
  NAND4X1 g05824(.A(n9031), .B(n9030), .C(n9029), .D(n9032), .Y(n9033));
  NOR2X1  g05825(.A(n9033), .B(n9028), .Y(n9034));
  NOR4X1  g05826(.A(n9007), .B(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C(n9019), .D(n9007), .Y(n9035));
  AOI22X1 g05827(.A0(n8980), .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B0(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(n8981), .Y(n9036));
  AOI22X1 g05828(.A0(n8983), .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B0(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(n8984), .Y(n9037));
  AOI22X1 g05829(.A0(n8986), .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B0(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(n8987), .Y(n9038));
  AOI22X1 g05830(.A0(n8989), .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B0(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(n8990), .Y(n9039));
  NAND4X1 g05831(.A(n9038), .B(n9037), .C(n9036), .D(n9039), .Y(n9040));
  AOI22X1 g05832(.A0(n8993), .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B0(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(n8994), .Y(n9041));
  AOI22X1 g05833(.A0(n8996), .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B0(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(n8997), .Y(n9042));
  AOI22X1 g05834(.A0(n8999), .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B0(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(n9000), .Y(n9043));
  AOI22X1 g05835(.A0(n9002), .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B0(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(n9003), .Y(n9044));
  NAND4X1 g05836(.A(n9043), .B(n9042), .C(n9041), .D(n9044), .Y(n9045));
  NOR2X1  g05837(.A(n9045), .B(n9040), .Y(n9046));
  NOR4X1  g05838(.A(n9007), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C(n8724), .D(n9007), .Y(n9047));
  AOI21X1 g05839(.A0(n8975), .A1(n8978), .B0(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .Y(n9048));
  INVX1   g05840(.A(n9048), .Y(n9049));
  INVX1   g05841(.A(n9046), .Y(n9051));
  AOI22X1 g05842(.A0(n8979), .A1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B0(n9007), .B1(n9051), .Y(n9052));
  AOI21X1 g05843(.A0(n8975), .A1(n8978), .B0(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .Y(n9053));
  INVX1   g05844(.A(n9053), .Y(n9054));
  AOI22X1 g05845(.A0(n8980), .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B0(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(n8981), .Y(n9055));
  AOI22X1 g05846(.A0(n8983), .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B0(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(n8984), .Y(n9056));
  AOI22X1 g05847(.A0(n8986), .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B0(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(n8987), .Y(n9057));
  AOI22X1 g05848(.A0(n8989), .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B0(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(n8990), .Y(n9058));
  NAND4X1 g05849(.A(n9057), .B(n9056), .C(n9055), .D(n9058), .Y(n9059));
  AOI22X1 g05850(.A0(n8993), .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B0(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(n8994), .Y(n9060));
  AOI22X1 g05851(.A0(n8996), .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B0(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(n8997), .Y(n9061));
  AOI22X1 g05852(.A0(n8999), .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B0(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(n9000), .Y(n9062));
  AOI22X1 g05853(.A0(n9002), .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B0(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(n9003), .Y(n9063));
  NAND4X1 g05854(.A(n9062), .B(n9061), .C(n9060), .D(n9063), .Y(n9064));
  NOR2X1  g05855(.A(n9064), .B(n9059), .Y(n9065));
  INVX1   g05856(.A(n9065), .Y(n9066));
  AOI22X1 g05857(.A0(n8979), .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B0(n9007), .B1(n9066), .Y(n9067));
  AOI22X1 g05858(.A0(n9054), .A1(n9067), .B0(n9052), .B1(n9049), .Y(n9068));
  NOR3X1  g05859(.A(n9068), .B(n9047), .C(n9035), .Y(n9069));
  INVX1   g05860(.A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .Y(n9070));
  INVX1   g05861(.A(n8980), .Y(n9071));
  NAND2X1 g05862(.A(n8981), .B(P2_INSTQUEUE_REG_1__1__SCAN_IN), .Y(n9072));
  OAI21X1 g05863(.A0(n9071), .A1(n9070), .B0(n9072), .Y(n9073));
  INVX1   g05864(.A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .Y(n9074));
  INVX1   g05865(.A(n8983), .Y(n9075));
  NAND2X1 g05866(.A(n8984), .B(P2_INSTQUEUE_REG_2__1__SCAN_IN), .Y(n9076));
  OAI21X1 g05867(.A0(n9075), .A1(n9074), .B0(n9076), .Y(n9077));
  NOR2X1  g05868(.A(n9077), .B(n9073), .Y(n9078));
  AOI22X1 g05869(.A0(n8986), .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B0(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(n8987), .Y(n9079));
  AOI22X1 g05870(.A0(n8989), .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B0(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(n8990), .Y(n9080));
  INVX1   g05871(.A(n8993), .Y(n9081));
  INVX1   g05872(.A(n8994), .Y(n9082));
  OAI22X1 g05873(.A0(n9081), .A1(n8950), .B0(n8957), .B1(n9082), .Y(n9083));
  INVX1   g05874(.A(n8996), .Y(n9084));
  INVX1   g05875(.A(n8997), .Y(n9085));
  OAI22X1 g05876(.A0(n9084), .A1(n8968), .B0(n8964), .B1(n9085), .Y(n9086));
  INVX1   g05877(.A(n8999), .Y(n9087));
  INVX1   g05878(.A(n9000), .Y(n9088));
  OAI22X1 g05879(.A0(n9087), .A1(n8961), .B0(n8947), .B1(n9088), .Y(n9089));
  INVX1   g05880(.A(n9002), .Y(n9090));
  INVX1   g05881(.A(n9003), .Y(n9091));
  OAI22X1 g05882(.A0(n9090), .A1(n8971), .B0(n8954), .B1(n9091), .Y(n9092));
  NOR4X1  g05883(.A(n9089), .B(n9086), .C(n9083), .D(n9092), .Y(n9093));
  NAND4X1 g05884(.A(n9080), .B(n9079), .C(n9078), .D(n9093), .Y(n9094));
  AOI22X1 g05885(.A0(n8979), .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B0(n9007), .B1(n9094), .Y(n9095));
  AOI21X1 g05886(.A0(n8975), .A1(n8978), .B0(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Y(n9096));
  INVX1   g05887(.A(n9096), .Y(n9097));
  NOR2X1  g05888(.A(n9097), .B(n9095), .Y(n9098));
  INVX1   g05889(.A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .Y(n9099));
  NAND2X1 g05890(.A(n8981), .B(P2_INSTQUEUE_REG_1__0__SCAN_IN), .Y(n9100));
  OAI21X1 g05891(.A0(n9071), .A1(n9099), .B0(n9100), .Y(n9101));
  INVX1   g05892(.A(P2_INSTQUEUE_REG_3__0__SCAN_IN), .Y(n9102));
  NAND2X1 g05893(.A(n8984), .B(P2_INSTQUEUE_REG_2__0__SCAN_IN), .Y(n9103));
  OAI21X1 g05894(.A0(n9075), .A1(n9102), .B0(n9103), .Y(n9104));
  NOR2X1  g05895(.A(n9104), .B(n9101), .Y(n9105));
  NAND2X1 g05896(.A(n8986), .B(P2_INSTQUEUE_REG_4__0__SCAN_IN), .Y(n9106));
  NAND2X1 g05897(.A(n8987), .B(P2_INSTQUEUE_REG_5__0__SCAN_IN), .Y(n9107));
  NAND2X1 g05898(.A(n9107), .B(n9106), .Y(n9108));
  NAND2X1 g05899(.A(n8989), .B(P2_INSTQUEUE_REG_7__0__SCAN_IN), .Y(n9109));
  NAND2X1 g05900(.A(n8990), .B(P2_INSTQUEUE_REG_6__0__SCAN_IN), .Y(n9110));
  NAND2X1 g05901(.A(n9110), .B(n9109), .Y(n9111));
  NOR2X1  g05902(.A(n9111), .B(n9108), .Y(n9112));
  OAI22X1 g05903(.A0(n9081), .A1(n8919), .B0(n8926), .B1(n9082), .Y(n9113));
  OAI22X1 g05904(.A0(n9084), .A1(n8938), .B0(n8934), .B1(n9085), .Y(n9114));
  NOR2X1  g05905(.A(n9114), .B(n9113), .Y(n9115));
  OAI22X1 g05906(.A0(n9087), .A1(n8931), .B0(n8916), .B1(n9088), .Y(n9116));
  OAI22X1 g05907(.A0(n9090), .A1(n8941), .B0(n8923), .B1(n9091), .Y(n9117));
  NOR2X1  g05908(.A(n9117), .B(n9116), .Y(n9118));
  NAND4X1 g05909(.A(n9115), .B(n9112), .C(n9105), .D(n9118), .Y(n9119));
  INVX1   g05910(.A(n9119), .Y(n9120));
  NOR4X1  g05911(.A(n9007), .B(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .C(n8721), .D(n9007), .Y(n9121));
  NOR2X1  g05912(.A(n9121), .B(n9098), .Y(n9122));
  AOI21X1 g05913(.A0(n9097), .A1(n9095), .B0(n9122), .Y(n9123));
  NOR2X1  g05914(.A(n9034), .B(n8979), .Y(n9124));
  AOI21X1 g05915(.A0(n8979), .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B0(n9124), .Y(n9125));
  AOI21X1 g05916(.A0(n8975), .A1(n8978), .B0(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .Y(n9126));
  INVX1   g05917(.A(n9126), .Y(n9127));
  NOR4X1  g05918(.A(n9007), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C(n8727), .D(n9007), .Y(n9128));
  NOR2X1  g05919(.A(n9128), .B(n9047), .Y(n9129));
  OAI21X1 g05920(.A0(n9127), .A1(n9125), .B0(n9129), .Y(n9130));
  NAND2X1 g05921(.A(n9127), .B(n9125), .Y(n9131));
  OAI21X1 g05922(.A0(n9130), .A1(n9123), .B0(n9131), .Y(n9132));
  NOR2X1  g05923(.A(n9132), .B(n9069), .Y(n9133));
  INVX1   g05924(.A(n9133), .Y(n9134));
  XOR2X1  g05925(.A(n9134), .B(n9006), .Y(n9137));
  INVX1   g05926(.A(n9137), .Y(n9138));
  NOR3X1  g05927(.A(n9017), .B(n9012), .C(n8979), .Y(n9139));
  XOR2X1  g05928(.A(n9139), .B(n9134), .Y(n9140));
  INVX1   g05929(.A(n9140), .Y(n9141));
  XOR2X1  g05930(.A(n9052), .B(n9049), .Y(n9142));
  INVX1   g05931(.A(n9142), .Y(n9143));
  NOR2X1  g05932(.A(n9128), .B(n9123), .Y(n9144));
  AOI21X1 g05933(.A0(n9067), .A1(n9054), .B0(n9144), .Y(n9145));
  XOR2X1  g05934(.A(n9145), .B(n9143), .Y(n9146));
  XOR2X1  g05935(.A(n9067), .B(n9054), .Y(n9147));
  XOR2X1  g05936(.A(n9147), .B(n9123), .Y(n9148));
  XOR2X1  g05937(.A(n9097), .B(n9095), .Y(n9149));
  XOR2X1  g05938(.A(n9149), .B(n9121), .Y(n9150));
  AOI22X1 g05939(.A0(n8979), .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B0(n9007), .B1(n9119), .Y(n9151));
  AOI21X1 g05940(.A0(n8975), .A1(n8978), .B0(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Y(n9152));
  XOR2X1  g05941(.A(n9152), .B(n9151), .Y(n9153));
  INVX1   g05942(.A(n9153), .Y(n9154));
  AOI21X1 g05943(.A0(n9154), .A1(n9150), .B0(n9148), .Y(n9155));
  XOR2X1  g05944(.A(n9127), .B(n9125), .Y(n9156));
  INVX1   g05945(.A(n9129), .Y(n9157));
  OAI22X1 g05946(.A0(n9123), .A1(n9157), .B0(n9068), .B1(n9047), .Y(n9158));
  XOR2X1  g05947(.A(n9158), .B(n9156), .Y(n9159));
  NOR4X1  g05948(.A(n9155), .B(n9146), .C(n9141), .D(n9159), .Y(n9160));
  NOR2X1  g05949(.A(n9160), .B(n9138), .Y(n9161));
  INVX1   g05950(.A(P2_FLUSH_REG_SCAN_IN), .Y(n9162));
  INVX1   g05951(.A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .Y(n9163));
  NOR2X1  g05952(.A(n9163), .B(n8720), .Y(n9164));
  INVX1   g05953(.A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .Y(n9165));
  INVX1   g05954(.A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .Y(n9166));
  INVX1   g05955(.A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .Y(n9167));
  INVX1   g05956(.A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .Y(n9168));
  INVX1   g05957(.A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .Y(n9169));
  INVX1   g05958(.A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .Y(n9170));
  INVX1   g05959(.A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .Y(n9171));
  INVX1   g05960(.A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .Y(n9172));
  INVX1   g05961(.A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .Y(n9173));
  INVX1   g05962(.A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .Y(n9174));
  INVX1   g05963(.A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .Y(n9175));
  INVX1   g05964(.A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .Y(n9176));
  INVX1   g05965(.A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .Y(n9177));
  INVX1   g05966(.A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .Y(n9178));
  INVX1   g05967(.A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .Y(n9179));
  NAND4X1 g05968(.A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .C(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .D(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .Y(n9180));
  NOR4X1  g05969(.A(n9179), .B(n9178), .C(n9177), .D(n9180), .Y(n9181));
  NAND4X1 g05970(.A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .C(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .D(n9181), .Y(n9182));
  NOR4X1  g05971(.A(n9176), .B(n9175), .C(n9174), .D(n9182), .Y(n9183));
  NAND4X1 g05972(.A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .C(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .D(n9183), .Y(n9184));
  NOR4X1  g05973(.A(n9173), .B(n9172), .C(n9171), .D(n9184), .Y(n9185));
  NAND4X1 g05974(.A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .C(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .D(n9185), .Y(n9186));
  NOR4X1  g05975(.A(n9170), .B(n9169), .C(n9168), .D(n9186), .Y(n9187));
  NAND4X1 g05976(.A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .B(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .C(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .D(n9187), .Y(n9188));
  NOR3X1  g05977(.A(n9188), .B(n9167), .C(n9166), .Y(n9189));
  XOR2X1  g05978(.A(n9189), .B(n9165), .Y(n9190));
  INVX1   g05979(.A(n9190), .Y(n9191));
  AOI21X1 g05980(.A0(n9191), .A1(n8720), .B0(n9164), .Y(n9192));
  INVX1   g05981(.A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .Y(n9193));
  NOR2X1  g05982(.A(n9193), .B(P2_STATE2_REG_0__SCAN_IN), .Y(n9194));
  AOI21X1 g05983(.A0(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A1(P2_STATE2_REG_0__SCAN_IN), .B0(n9194), .Y(n9195));
  NOR2X1  g05984(.A(n9195), .B(n9192), .Y(n9196));
  AOI21X1 g05985(.A0(n9192), .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B0(n9196), .Y(n9197));
  NOR2X1  g05986(.A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B(P2_STATE2_REG_0__SCAN_IN), .Y(n9198));
  AOI21X1 g05987(.A0(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A1(P2_STATE2_REG_0__SCAN_IN), .B0(n9198), .Y(n9199));
  INVX1   g05988(.A(n9199), .Y(n9200));
  XOR2X1  g05989(.A(n9200), .B(n9195), .Y(n9201));
  NOR2X1  g05990(.A(n9201), .B(n9192), .Y(n9202));
  AOI21X1 g05991(.A0(n9192), .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B0(n9202), .Y(n9203));
  NOR3X1  g05992(.A(n9203), .B(n9197), .C(n9162), .Y(n9204));
  INVX1   g05993(.A(P2_STATE2_REG_1__SCAN_IN), .Y(n9205));
  AOI21X1 g05994(.A0(n9162), .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B0(n9205), .Y(n9206));
  INVX1   g05995(.A(n9206), .Y(n9207));
  INVX1   g05996(.A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Y(n9208));
  INVX1   g05997(.A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Y(n9209));
  AOI21X1 g05998(.A0(n9209), .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B0(n9208), .Y(n9210));
  NAND3X1 g05999(.A(n9209), .B(n9208), .C(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n9211));
  AOI21X1 g06000(.A0(n9211), .A1(n8732), .B0(n9210), .Y(n9212));
  XOR2X1  g06001(.A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n8727), .Y(n9213));
  XOR2X1  g06002(.A(n9213), .B(n9212), .Y(n9214));
  OAI22X1 g06003(.A0(n9207), .A1(n9204), .B0(P2_STATE2_REG_1__SCAN_IN), .B1(n9214), .Y(n9215));
  INVX1   g06004(.A(n9197), .Y(n9216));
  AOI21X1 g06005(.A0(n9162), .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B0(n9205), .Y(n9217));
  OAI21X1 g06006(.A0(n9216), .A1(n9162), .B0(n9217), .Y(n9218));
  NOR3X1  g06007(.A(P2_FLUSH_REG_SCAN_IN), .B(n9019), .C(n9205), .Y(n9219));
  NOR2X1  g06008(.A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B(n9019), .Y(n9220));
  INVX1   g06009(.A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .Y(n9221));
  NOR2X1  g06010(.A(n9221), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n9222));
  INVX1   g06011(.A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .Y(n9223));
  AOI21X1 g06012(.A0(n9223), .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B0(n9212), .Y(n9224));
  AOI21X1 g06013(.A0(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A1(n8727), .B0(n9224), .Y(n9225));
  AOI21X1 g06014(.A0(n9221), .A1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B0(n9225), .Y(n9226));
  INVX1   g06015(.A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .Y(n9227));
  NOR2X1  g06016(.A(n9227), .B(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .Y(n9228));
  NOR3X1  g06017(.A(n9228), .B(n9226), .C(n9222), .Y(n9229));
  NOR2X1  g06018(.A(n9229), .B(n9220), .Y(n9230));
  NOR2X1  g06019(.A(n9230), .B(P2_STATE2_REG_1__SCAN_IN), .Y(n9231));
  NOR2X1  g06020(.A(n9231), .B(n9219), .Y(n9232));
  NOR2X1  g06021(.A(n9226), .B(n9222), .Y(n9233));
  XOR2X1  g06022(.A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B(n9019), .Y(n9234));
  XOR2X1  g06023(.A(n9234), .B(n9233), .Y(n9235));
  INVX1   g06024(.A(n9235), .Y(n9236));
  AOI21X1 g06025(.A0(n9236), .A1(n9205), .B0(n9219), .Y(n9237));
  AOI21X1 g06026(.A0(n9162), .A1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B0(n9205), .Y(n9238));
  XOR2X1  g06027(.A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n8724), .Y(n9239));
  XOR2X1  g06028(.A(n9239), .B(n9225), .Y(n9240));
  NOR2X1  g06029(.A(n9240), .B(P2_STATE2_REG_1__SCAN_IN), .Y(n9241));
  NOR2X1  g06030(.A(n9241), .B(n9238), .Y(n9242));
  INVX1   g06031(.A(n9242), .Y(n9243));
  XOR2X1  g06032(.A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n8721), .Y(n9244));
  INVX1   g06033(.A(n9244), .Y(n9245));
  AOI21X1 g06034(.A0(n9245), .A1(n9205), .B0(n9243), .Y(n9246));
  NAND4X1 g06035(.A(n9237), .B(n9232), .C(n9218), .D(n9246), .Y(n9247));
  NOR2X1  g06036(.A(n9247), .B(n9215), .Y(n9248));
  NAND2X1 g06037(.A(n9203), .B(n9216), .Y(n9249));
  AOI21X1 g06038(.A0(n9162), .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B0(n9205), .Y(n9250));
  OAI21X1 g06039(.A0(n9249), .A1(n9162), .B0(n9250), .Y(n9251));
  NOR2X1  g06040(.A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n8721), .Y(n9252));
  XOR2X1  g06041(.A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n8732), .Y(n9253));
  XOR2X1  g06042(.A(n9253), .B(n9252), .Y(n9254));
  INVX1   g06043(.A(n9254), .Y(n9255));
  AOI21X1 g06044(.A0(n9255), .A1(n9205), .B0(n9243), .Y(n9256));
  NAND4X1 g06045(.A(n9251), .B(n9237), .C(n9232), .D(n9256), .Y(n9257));
  OAI21X1 g06046(.A0(n9257), .A1(n9215), .B0(n9232), .Y(n9258));
  NOR2X1  g06047(.A(n9258), .B(n9248), .Y(n9259));
  OAI22X1 g06048(.A0(n9161), .A1(n8977), .B0(n8979), .B1(n9259), .Y(n9260));
  NAND2X1 g06049(.A(n9260), .B(n8915), .Y(n9261));
  NAND2X1 g06050(.A(n8978), .B(P2_STATE2_REG_0__SCAN_IN), .Y(n9262));
  NOR2X1  g06051(.A(n9262), .B(n9230), .Y(n9263));
  OAI21X1 g06052(.A0(n9022), .A1(n8946), .B0(P2_STATE2_REG_0__SCAN_IN), .Y(n9264));
  NOR3X1  g06053(.A(n9264), .B(n9263), .C(n9140), .Y(n9265));
  INVX1   g06054(.A(n9264), .Y(n9266));
  AOI21X1 g06055(.A0(n9266), .A1(n9146), .B0(n8720), .Y(n9267));
  OAI22X1 g06056(.A0(n9240), .A1(n9262), .B0(n8724), .B1(P2_STATE2_REG_0__SCAN_IN), .Y(n9268));
  INVX1   g06057(.A(n9150), .Y(n9269));
  AOI21X1 g06058(.A0(n9266), .A1(n9269), .B0(n8720), .Y(n9270));
  NOR3X1  g06059(.A(n9022), .B(n8978), .C(n8720), .Y(n9271));
  AOI21X1 g06060(.A0(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A1(n8720), .B0(n9271), .Y(n9272));
  OAI21X1 g06061(.A0(n9262), .A1(n9254), .B0(n9272), .Y(n9273));
  NOR2X1  g06062(.A(n8978), .B(n8720), .Y(n9274));
  NOR2X1  g06063(.A(n9262), .B(n9022), .Y(n9275));
  NAND3X1 g06064(.A(n9275), .B(n9274), .C(n9154), .Y(n9276));
  NOR2X1  g06065(.A(n8946), .B(n8720), .Y(n9277));
  NAND2X1 g06066(.A(n9022), .B(P2_STATE2_REG_0__SCAN_IN), .Y(n9278));
  OAI21X1 g06067(.A0(n8721), .A1(P2_STATE2_REG_0__SCAN_IN), .B0(n9278), .Y(n9279));
  AOI21X1 g06068(.A0(n9277), .A1(n9245), .B0(n9279), .Y(n9280));
  AOI21X1 g06069(.A0(n9274), .A1(n9154), .B0(n9275), .Y(n9281));
  OAI21X1 g06070(.A0(n9281), .A1(n9280), .B0(n9276), .Y(n9282));
  AOI21X1 g06071(.A0(n9273), .A1(n9270), .B0(n9282), .Y(n9283));
  NOR2X1  g06072(.A(n8975), .B(n8720), .Y(n9284));
  AOI21X1 g06073(.A0(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A1(n8720), .B0(n9284), .Y(n9285));
  OAI21X1 g06074(.A0(n9262), .A1(n9214), .B0(n9285), .Y(n9286));
  INVX1   g06075(.A(n9148), .Y(n9287));
  NOR3X1  g06076(.A(n9287), .B(n8978), .C(n8720), .Y(n9288));
  OAI22X1 g06077(.A0(n9286), .A1(n9288), .B0(n9273), .B1(n9270), .Y(n9289));
  NAND3X1 g06078(.A(n9286), .B(n9274), .C(n9148), .Y(n9290));
  OAI21X1 g06079(.A0(n9289), .A1(n9283), .B0(n9290), .Y(n9291));
  AOI21X1 g06080(.A0(n9268), .A1(n9267), .B0(n9291), .Y(n9292));
  AOI22X1 g06081(.A0(n9236), .A1(n9277), .B0(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B1(n8720), .Y(n9293));
  NAND3X1 g06082(.A(n9293), .B(n9266), .C(n9159), .Y(n9294));
  OAI21X1 g06083(.A0(n9268), .A1(n9267), .B0(n9294), .Y(n9295));
  NOR2X1  g06084(.A(n9295), .B(n9292), .Y(n9296));
  INVX1   g06085(.A(n9263), .Y(n9297));
  NOR2X1  g06086(.A(n9264), .B(n9140), .Y(n9298));
  NOR2X1  g06087(.A(n9298), .B(n9297), .Y(n9299));
  AOI21X1 g06088(.A0(n9266), .A1(n9159), .B0(n9293), .Y(n9300));
  NOR3X1  g06089(.A(n9300), .B(n9299), .C(n9296), .Y(n9301));
  XOR2X1  g06090(.A(n9298), .B(n9297), .Y(n9303));
  OAI21X1 g06091(.A0(n9301), .A1(n9265), .B0(n9303), .Y(n9304));
  NOR4X1  g06092(.A(n9263), .B(n9137), .C(P2_STATE2_REG_0__SCAN_IN), .D(n9264), .Y(n9305));
  NOR2X1  g06093(.A(n9299), .B(n9305), .Y(n9307));
  NAND2X1 g06094(.A(n9307), .B(n9304), .Y(n9308));
  NOR2X1  g06095(.A(n9022), .B(n8978), .Y(n9309));
  NOR2X1  g06096(.A(n8975), .B(n8978), .Y(n9310));
  INVX1   g06097(.A(n9310), .Y(n9311));
  AOI21X1 g06098(.A0(n8758), .A1(n8741), .B0(n8855), .Y(n9312));
  INVX1   g06099(.A(n9312), .Y(n9313));
  NOR2X1  g06100(.A(n8724), .B(P2_INSTQUEUE_REG_14__6__SCAN_IN), .Y(n9314));
  NOR3X1  g06101(.A(n9314), .B(n8762), .C(n8722), .Y(n9315));
  NOR2X1  g06102(.A(n8724), .B(P2_INSTQUEUE_REG_11__6__SCAN_IN), .Y(n9316));
  NOR3X1  g06103(.A(n9316), .B(n8765), .C(n8728), .Y(n9317));
  NOR2X1  g06104(.A(n8724), .B(P2_INSTQUEUE_REG_13__6__SCAN_IN), .Y(n9318));
  NOR3X1  g06105(.A(n9318), .B(n8771), .C(n8733), .Y(n9319));
  NOR2X1  g06106(.A(n8724), .B(P2_INSTQUEUE_REG_10__6__SCAN_IN), .Y(n9320));
  NOR3X1  g06107(.A(n9320), .B(n8774), .C(n8737), .Y(n9321));
  NOR4X1  g06108(.A(n9319), .B(n9317), .C(n9315), .D(n9321), .Y(n9322));
  NOR2X1  g06109(.A(n8724), .B(P2_INSTQUEUE_REG_15__6__SCAN_IN), .Y(n9323));
  NOR3X1  g06110(.A(n9323), .B(n8781), .C(n8742), .Y(n9324));
  NOR2X1  g06111(.A(n8724), .B(P2_INSTQUEUE_REG_9__6__SCAN_IN), .Y(n9325));
  NOR3X1  g06112(.A(n8784), .B(n9325), .C(n8746), .Y(n9326));
  NOR2X1  g06113(.A(n8724), .B(P2_INSTQUEUE_REG_8__6__SCAN_IN), .Y(n9327));
  NOR3X1  g06114(.A(n8790), .B(n9327), .C(n8750), .Y(n9328));
  NOR2X1  g06115(.A(n8724), .B(P2_INSTQUEUE_REG_12__6__SCAN_IN), .Y(n9329));
  NOR3X1  g06116(.A(n9329), .B(n8793), .C(n8754), .Y(n9330));
  NOR4X1  g06117(.A(n9328), .B(n9326), .C(n9324), .D(n9330), .Y(n9331));
  NAND3X1 g06118(.A(n8825), .B(n9331), .C(n9322), .Y(n9332));
  NOR4X1  g06119(.A(n9313), .B(n9311), .C(n8914), .D(n9332), .Y(n9333));
  NAND2X1 g06120(.A(n8840), .B(n8833), .Y(n9334));
  NAND2X1 g06121(.A(n8854), .B(n8847), .Y(n9335));
  NOR2X1  g06122(.A(n9335), .B(n9334), .Y(n9336));
  NAND2X1 g06123(.A(n8869), .B(n8862), .Y(n9337));
  NAND2X1 g06124(.A(n8883), .B(n8876), .Y(n9338));
  NOR2X1  g06125(.A(n9338), .B(n9337), .Y(n9339));
  NOR4X1  g06126(.A(n9339), .B(n9336), .C(n8826), .D(n8913), .Y(n9340));
  AOI21X1 g06127(.A0(n9340), .A1(n9309), .B0(n9333), .Y(n9341));
  NOR2X1  g06128(.A(n9341), .B(n9308), .Y(n9342));
  INVX1   g06129(.A(n9342), .Y(n9343));
  NOR3X1  g06130(.A(n9214), .B(n8975), .C(n8946), .Y(n9347));
  AOI21X1 g06131(.A0(n9255), .A1(n8977), .B0(n9347), .Y(n9348));
  AOI21X1 g06132(.A0(n9022), .A1(n8978), .B0(n9214), .Y(n9349));
  AOI21X1 g06133(.A0(n9255), .A1(n8976), .B0(n9349), .Y(n9350));
  NAND3X1 g06134(.A(n9240), .B(n9350), .C(n9348), .Y(n9354));
  AOI21X1 g06135(.A0(n9236), .A1(n8977), .B0(n9354), .Y(n9355));
  OAI21X1 g06136(.A0(n9235), .A1(n8977), .B0(n9355), .Y(n9356));
  NAND2X1 g06137(.A(n9356), .B(n9230), .Y(n9357));
  INVX1   g06138(.A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .Y(n9358));
  AOI21X1 g06139(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n9358), .B0(n8723), .Y(n9359));
  INVX1   g06140(.A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .Y(n9360));
  AOI21X1 g06141(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n9360), .B0(n8729), .Y(n9361));
  AOI22X1 g06142(.A0(n8760), .A1(n9361), .B0(n9359), .B1(n8759), .Y(n9362));
  INVX1   g06143(.A(P2_INSTQUEUE_REG_13__4__SCAN_IN), .Y(n9363));
  AOI21X1 g06144(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n9363), .B0(n8734), .Y(n9364));
  INVX1   g06145(.A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .Y(n9365));
  AOI21X1 g06146(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n9365), .B0(n8738), .Y(n9366));
  AOI22X1 g06147(.A0(n8769), .A1(n9366), .B0(n9364), .B1(n8768), .Y(n9367));
  INVX1   g06148(.A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .Y(n9368));
  AOI21X1 g06149(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n9368), .B0(n8743), .Y(n9369));
  INVX1   g06150(.A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .Y(n9370));
  AOI21X1 g06151(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n9370), .B0(n8748), .Y(n9371));
  AOI22X1 g06152(.A0(n8779), .A1(n9371), .B0(n9369), .B1(n8778), .Y(n9372));
  INVX1   g06153(.A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .Y(n9373));
  AOI21X1 g06154(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n9373), .B0(n8752), .Y(n9374));
  INVX1   g06155(.A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .Y(n9375));
  AOI21X1 g06156(.A0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n9375), .B0(n8755), .Y(n9376));
  AOI22X1 g06157(.A0(n8788), .A1(n9376), .B0(n9374), .B1(n8787), .Y(n9377));
  NAND4X1 g06158(.A(n9372), .B(n9367), .C(n9362), .D(n9377), .Y(n9378));
  NOR2X1  g06159(.A(n8724), .B(P2_INSTQUEUE_REG_14__5__SCAN_IN), .Y(n9379));
  NOR3X1  g06160(.A(n9379), .B(n8798), .C(n8722), .Y(n9380));
  NOR2X1  g06161(.A(n8724), .B(P2_INSTQUEUE_REG_11__5__SCAN_IN), .Y(n9381));
  NOR3X1  g06162(.A(n9381), .B(n8801), .C(n8728), .Y(n9382));
  NOR2X1  g06163(.A(n8724), .B(P2_INSTQUEUE_REG_13__5__SCAN_IN), .Y(n9383));
  NOR3X1  g06164(.A(n9383), .B(n8805), .C(n8733), .Y(n9384));
  NOR2X1  g06165(.A(n8724), .B(P2_INSTQUEUE_REG_10__5__SCAN_IN), .Y(n9385));
  NOR3X1  g06166(.A(n9385), .B(n8808), .C(n8737), .Y(n9386));
  NOR4X1  g06167(.A(n9384), .B(n9382), .C(n9380), .D(n9386), .Y(n9387));
  NOR2X1  g06168(.A(n8724), .B(P2_INSTQUEUE_REG_15__5__SCAN_IN), .Y(n9388));
  NOR3X1  g06169(.A(n9388), .B(n8812), .C(n8742), .Y(n9389));
  NOR2X1  g06170(.A(n8724), .B(P2_INSTQUEUE_REG_9__5__SCAN_IN), .Y(n9390));
  NOR3X1  g06171(.A(n8815), .B(n9390), .C(n8746), .Y(n9391));
  NOR2X1  g06172(.A(n8724), .B(P2_INSTQUEUE_REG_8__5__SCAN_IN), .Y(n9392));
  NOR3X1  g06173(.A(n8819), .B(n9392), .C(n8750), .Y(n9393));
  NOR2X1  g06174(.A(n8724), .B(P2_INSTQUEUE_REG_12__5__SCAN_IN), .Y(n9394));
  NOR3X1  g06175(.A(n9394), .B(n8822), .C(n8754), .Y(n9395));
  NOR4X1  g06176(.A(n9393), .B(n9391), .C(n9389), .D(n9395), .Y(n9396));
  NAND4X1 g06177(.A(n8884), .B(n9396), .C(n9387), .D(n8913), .Y(n9397));
  NOR4X1  g06178(.A(n8855), .B(n8796), .C(n9378), .D(n9397), .Y(n9398));
  AOI22X1 g06179(.A0(n9340), .A1(n9310), .B0(n8978), .B1(n9398), .Y(n9399));
  INVX1   g06180(.A(n9399), .Y(n9400));
  NOR4X1  g06181(.A(n9313), .B(n8979), .C(n8914), .D(n9332), .Y(n9401));
  AOI22X1 g06182(.A0(n9400), .A1(n9357), .B0(n9308), .B1(n9401), .Y(n9402));
  NAND3X1 g06183(.A(n9402), .B(n9343), .C(n9261), .Y(n9403));
  INVX1   g06184(.A(n8915), .Y(n9404));
  NOR3X1  g06185(.A(n9160), .B(n9138), .C(n8977), .Y(n9405));
  AOI21X1 g06186(.A0(n9259), .A1(n9007), .B0(n9405), .Y(n9406));
  NOR2X1  g06187(.A(n9406), .B(n9404), .Y(n9407));
  INVX1   g06188(.A(n9407), .Y(n9408));
  AOI22X1 g06189(.A0(n9340), .A1(n9310), .B0(n9007), .B1(n9398), .Y(n9409));
  NOR3X1  g06190(.A(n9409), .B(n9357), .C(n8619), .Y(n9410));
  AOI21X1 g06191(.A0(n9333), .A1(n9308), .B0(n9410), .Y(n9411));
  INVX1   g06192(.A(n9401), .Y(n9412));
  NOR2X1  g06193(.A(n9412), .B(n9308), .Y(n9413));
  INVX1   g06194(.A(n9413), .Y(n9414));
  INVX1   g06195(.A(n9309), .Y(n9415));
  INVX1   g06196(.A(n9340), .Y(n9416));
  XOR2X1  g06197(.A(P2_STATE_REG_1__SCAN_IN), .B(n8614), .Y(n9417));
  NOR3X1  g06198(.A(n9417), .B(n8619), .C(P2_STATE_REG_0__SCAN_IN), .Y(n9418));
  INVX1   g06199(.A(n9418), .Y(n9419));
  NOR3X1  g06200(.A(n9419), .B(n9416), .C(n9415), .Y(n9420));
  NAND4X1 g06201(.A(n9398), .B(n9356), .C(n9230), .D(n9418), .Y(n9421));
  NOR3X1  g06202(.A(n8913), .B(n9339), .C(n8826), .Y(n9422));
  AOI21X1 g06203(.A0(n9422), .A1(n8946), .B0(n9336), .Y(n9423));
  NOR2X1  g06204(.A(n8978), .B(n9378), .Y(n9424));
  NOR3X1  g06205(.A(n9424), .B(n9309), .C(n8914), .Y(n9425));
  NAND3X1 g06206(.A(n9396), .B(n9387), .C(n8796), .Y(n9426));
  NAND3X1 g06207(.A(n9426), .B(n9332), .C(n8884), .Y(n9427));
  OAI21X1 g06208(.A0(n9332), .A1(n9378), .B0(n9426), .Y(n9428));
  AOI21X1 g06209(.A0(n9427), .A1(n8976), .B0(n9428), .Y(n9429));
  OAI21X1 g06210(.A0(n9425), .A1(n8855), .B0(n9429), .Y(n9430));
  NAND2X1 g06211(.A(n9367), .B(n9362), .Y(n9431));
  NAND2X1 g06212(.A(n9377), .B(n9372), .Y(n9432));
  NOR2X1  g06213(.A(n9432), .B(n9431), .Y(n9433));
  AOI21X1 g06214(.A0(n9396), .A1(n9387), .B0(n8796), .Y(n9434));
  NOR3X1  g06215(.A(n9434), .B(n8855), .C(n9433), .Y(n9435));
  NOR3X1  g06216(.A(n9435), .B(n9430), .C(n9423), .Y(n9436));
  NAND2X1 g06217(.A(n9436), .B(n9421), .Y(n9437));
  AOI21X1 g06218(.A0(n9420), .A1(n9308), .B0(n9437), .Y(n9438));
  NAND3X1 g06219(.A(n9438), .B(n9414), .C(n9411), .Y(n9439));
  NAND2X1 g06220(.A(n8898), .B(n8891), .Y(n9440));
  NAND2X1 g06221(.A(n8912), .B(n8905), .Y(n9441));
  NOR2X1  g06222(.A(n9441), .B(n9440), .Y(n9442));
  NAND2X1 g06223(.A(n9434), .B(n9433), .Y(n9443));
  NAND2X1 g06224(.A(n9332), .B(n9378), .Y(n9444));
  NAND4X1 g06225(.A(n9443), .B(n9426), .C(n8884), .D(n9444), .Y(n9445));
  NAND2X1 g06226(.A(n9445), .B(n8975), .Y(n9446));
  AOI21X1 g06227(.A0(n9427), .A1(n8976), .B0(n8855), .Y(n9447));
  AOI21X1 g06228(.A0(n9447), .A1(n9446), .B0(n9442), .Y(n9448));
  NAND4X1 g06229(.A(n8825), .B(n8796), .C(n9433), .D(n8884), .Y(n9449));
  NOR3X1  g06230(.A(n8855), .B(n8796), .C(n9378), .Y(n9450));
  AOI21X1 g06231(.A0(n8758), .A1(n8741), .B0(n8884), .Y(n9451));
  NOR2X1  g06232(.A(n9451), .B(n9450), .Y(n9452));
  AOI22X1 g06233(.A0(n9387), .A1(n9396), .B0(n9331), .B1(n9322), .Y(n9453));
  AOI22X1 g06234(.A0(n8913), .A1(n9332), .B0(n9336), .B1(n9453), .Y(n9454));
  NAND2X1 g06235(.A(n9454), .B(n9452), .Y(n9455));
  AOI21X1 g06236(.A0(n9449), .A1(n8855), .B0(n9455), .Y(n9456));
  NOR2X1  g06237(.A(n8913), .B(n8855), .Y(n9457));
  XOR2X1  g06238(.A(n9022), .B(n8978), .Y(n9458));
  NOR3X1  g06239(.A(n9426), .B(n8884), .C(n9378), .Y(n9459));
  NOR2X1  g06240(.A(n9434), .B(n8975), .Y(n9460));
  OAI21X1 g06241(.A0(n9460), .A1(n9459), .B0(n9458), .Y(n9461));
  AOI21X1 g06242(.A0(n9331), .A1(n9322), .B0(n8825), .Y(n9462));
  NOR2X1  g06243(.A(n8884), .B(n9378), .Y(n9463));
  NAND4X1 g06244(.A(n9457), .B(n9462), .C(n9310), .D(n9463), .Y(n9464));
  OAI21X1 g06245(.A0(n9309), .A1(n8976), .B0(n9378), .Y(n9465));
  NAND2X1 g06246(.A(n8810), .B(n8803), .Y(n9466));
  NAND2X1 g06247(.A(n8824), .B(n8817), .Y(n9467));
  NOR2X1  g06248(.A(n9467), .B(n9466), .Y(n9468));
  OAI21X1 g06249(.A0(n9339), .A1(n9468), .B0(n9309), .Y(n9469));
  INVX1   g06250(.A(n8796), .Y(n9470));
  OAI21X1 g06251(.A0(n8978), .A1(n9470), .B0(n8855), .Y(n9471));
  NAND4X1 g06252(.A(n9469), .B(n9465), .C(n9464), .D(n9471), .Y(n9472));
  AOI21X1 g06253(.A0(n9461), .A1(n9457), .B0(n9472), .Y(n9473));
  OAI21X1 g06254(.A0(n9456), .A1(n9311), .B0(n9473), .Y(n9474));
  NOR3X1  g06255(.A(n9474), .B(n9448), .C(n8915), .Y(n9475));
  INVX1   g06256(.A(n9417), .Y(n9476));
  NAND4X1 g06257(.A(n9398), .B(n8976), .C(P2_STATE2_REG_0__SCAN_IN), .D(n9476), .Y(n9477));
  NAND3X1 g06258(.A(n9422), .B(n9274), .C(n8855), .Y(n9478));
  NOR3X1  g06259(.A(n8975), .B(n8796), .C(n8720), .Y(n9479));
  NOR4X1  g06260(.A(n9339), .B(n8855), .C(n8825), .D(n8913), .Y(n9480));
  NAND4X1 g06261(.A(n9479), .B(n8946), .C(n9378), .D(n9480), .Y(n9481));
  NAND4X1 g06262(.A(n9284), .B(n8946), .C(n8796), .D(n9480), .Y(n9482));
  NAND4X1 g06263(.A(n9481), .B(n9478), .C(n9477), .D(n9482), .Y(n9483));
  INVX1   g06264(.A(P2_EBX_REG_1__SCAN_IN), .Y(n9484));
  NAND4X1 g06265(.A(n9457), .B(n9007), .C(P2_STATE2_REG_0__SCAN_IN), .D(n9459), .Y(n9485));
  NAND3X1 g06266(.A(n8975), .B(n8978), .C(P2_STATE2_REG_0__SCAN_IN), .Y(n9486));
  NAND4X1 g06267(.A(n8913), .B(n8884), .C(n9468), .D(n9450), .Y(n9487));
  NOR2X1  g06268(.A(n9487), .B(n9486), .Y(n9488));
  AOI22X1 g06269(.A0(P2_REIP_REG_1__SCAN_IN), .A1(n9488), .B0(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(P2_STATE2_REG_1__SCAN_IN), .Y(n9489));
  OAI21X1 g06270(.A0(n9485), .A1(n9484), .B0(n9489), .Y(n9490));
  AOI21X1 g06271(.A0(n9483), .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B0(n9490), .Y(n9491));
  NAND2X1 g06272(.A(n9479), .B(n8946), .Y(n9492));
  OAI22X1 g06273(.A0(n9464), .A1(n8720), .B0(n9468), .B1(n9492), .Y(n9493));
  NOR2X1  g06274(.A(n9332), .B(n9378), .Y(n9494));
  NOR2X1  g06275(.A(n9434), .B(n9433), .Y(n9495));
  NOR4X1  g06276(.A(n9494), .B(n9462), .C(n9339), .D(n9495), .Y(n9496));
  NAND3X1 g06277(.A(n8913), .B(n8758), .C(n8741), .Y(n9497));
  NOR2X1  g06278(.A(n9262), .B(n8975), .Y(n9498));
  OAI21X1 g06279(.A0(n9497), .A1(n9427), .B0(n9498), .Y(n9499));
  NAND4X1 g06280(.A(n8978), .B(n8913), .C(P2_STATE2_REG_0__SCAN_IN), .D(n8975), .Y(n9500));
  OAI21X1 g06281(.A0(n9500), .A1(n9496), .B0(n9499), .Y(n9501));
  NAND2X1 g06282(.A(n9463), .B(n9462), .Y(n9502));
  NAND3X1 g06283(.A(n9502), .B(n9275), .C(n9442), .Y(n9503));
  NOR4X1  g06284(.A(n8914), .B(n8855), .C(n8826), .D(n9262), .Y(n9504));
  NOR2X1  g06285(.A(n9262), .B(n9336), .Y(n9505));
  NOR3X1  g06286(.A(n9505), .B(n9504), .C(n9271), .Y(n9506));
  NAND2X1 g06287(.A(n9506), .B(n9503), .Y(n9507));
  NAND4X1 g06288(.A(n8825), .B(n8758), .C(n8741), .D(n8884), .Y(n9508));
  OAI21X1 g06289(.A0(n9508), .A1(n9434), .B0(n8855), .Y(n9509));
  NAND2X1 g06290(.A(n8825), .B(n8796), .Y(n9510));
  OAI22X1 g06291(.A0(n9442), .A1(n9434), .B0(n8855), .B1(n9510), .Y(n9511));
  NOR3X1  g06292(.A(n9511), .B(n9451), .C(n9450), .Y(n9512));
  NAND2X1 g06293(.A(n9284), .B(n8946), .Y(n9513));
  AOI21X1 g06294(.A0(n9512), .A1(n9509), .B0(n9513), .Y(n9514));
  NOR4X1  g06295(.A(n9507), .B(n9501), .C(n9493), .D(n9514), .Y(n9515));
  NAND2X1 g06296(.A(n9442), .B(n8884), .Y(n9516));
  NAND2X1 g06297(.A(n9274), .B(n8855), .Y(n9517));
  NOR3X1  g06298(.A(n9517), .B(n9516), .C(n8826), .Y(n9518));
  NAND3X1 g06299(.A(n9457), .B(n8884), .C(n9468), .Y(n9519));
  NOR4X1  g06300(.A(n9278), .B(n8978), .C(n9470), .D(n9519), .Y(n9520));
  NAND3X1 g06301(.A(n9476), .B(n8978), .C(P2_STATE2_REG_0__SCAN_IN), .Y(n9521));
  NOR2X1  g06302(.A(P2_STATE2_REG_0__SCAN_IN), .B(P2_STATE2_REG_1__SCAN_IN), .Y(n9522));
  INVX1   g06303(.A(n9522), .Y(n9523));
  OAI22X1 g06304(.A0(n9521), .A1(n9487), .B0(n9208), .B1(n9523), .Y(n9524));
  NOR4X1  g06305(.A(n9488), .B(n9520), .C(n9518), .D(n9524), .Y(n9525));
  OAI21X1 g06306(.A0(n9515), .A1(n8732), .B0(n9525), .Y(n9526));
  OAI21X1 g06307(.A0(n9459), .A1(n8913), .B0(n8978), .Y(n9527));
  AOI21X1 g06308(.A0(n9445), .A1(n8913), .B0(n9527), .Y(n9528));
  NAND2X1 g06309(.A(n9332), .B(n9022), .Y(n9529));
  OAI21X1 g06310(.A0(n9529), .A1(n9459), .B0(P2_STATE2_REG_0__SCAN_IN), .Y(n9530));
  NOR2X1  g06311(.A(n9530), .B(n9528), .Y(n9531));
  INVX1   g06312(.A(P2_EBX_REG_0__SCAN_IN), .Y(n9532));
  NAND3X1 g06313(.A(n9463), .B(n9457), .C(n9462), .Y(n9533));
  NOR4X1  g06314(.A(n8979), .B(n9532), .C(n8720), .D(n9533), .Y(n9534));
  OAI21X1 g06315(.A0(n9193), .A1(n9205), .B0(n9523), .Y(n9535));
  NOR3X1  g06316(.A(n9535), .B(n9505), .C(n9504), .Y(n9536));
  NAND2X1 g06317(.A(n9536), .B(n9499), .Y(n9537));
  INVX1   g06318(.A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .Y(n9538));
  NAND4X1 g06319(.A(n9022), .B(n8978), .C(P2_STATE2_REG_0__SCAN_IN), .D(n9476), .Y(n9539));
  NOR2X1  g06320(.A(n9539), .B(n9487), .Y(n9540));
  NOR3X1  g06321(.A(n9519), .B(n9492), .C(n9433), .Y(n9541));
  NOR4X1  g06322(.A(n9541), .B(n9518), .C(n9540), .D(n9520), .Y(n9542));
  AOI22X1 g06323(.A0(n9284), .A1(n8946), .B0(P2_REIP_REG_0__SCAN_IN), .B1(n9488), .Y(n9543));
  OAI22X1 g06324(.A0(n9542), .A1(n9538), .B0(n9456), .B1(n9543), .Y(n9544));
  NOR4X1  g06325(.A(n9537), .B(n9534), .C(n9531), .D(n9544), .Y(n9545));
  OAI22X1 g06326(.A0(n9533), .A1(n9486), .B0(n9209), .B1(n9523), .Y(n9546));
  INVX1   g06327(.A(n9500), .Y(n9547));
  AOI21X1 g06328(.A0(n9547), .A1(n9445), .B0(n9546), .Y(n9548));
  NAND2X1 g06329(.A(n9548), .B(n9499), .Y(n9549));
  NOR3X1  g06330(.A(n9459), .B(n9486), .C(n8913), .Y(n9550));
  NOR4X1  g06331(.A(n9504), .B(n9550), .C(n9271), .D(n9505), .Y(n9551));
  NAND3X1 g06332(.A(n9454), .B(n9452), .C(n9509), .Y(n9552));
  NAND3X1 g06333(.A(n9552), .B(n9284), .C(n8946), .Y(n9553));
  NOR2X1  g06334(.A(n9464), .B(n8720), .Y(n9554));
  NOR2X1  g06335(.A(n9492), .B(n9468), .Y(n9555));
  NOR3X1  g06336(.A(n9555), .B(n9554), .C(n9541), .Y(n9556));
  NAND3X1 g06337(.A(n9556), .B(n9553), .C(n9551), .Y(n9557));
  NAND2X1 g06338(.A(n9481), .B(n8721), .Y(n9558));
  OAI22X1 g06339(.A0(n9557), .A1(n9549), .B0(n9546), .B1(n9558), .Y(n9559));
  NOR2X1  g06340(.A(n9559), .B(n9545), .Y(n9560));
  XOR2X1  g06341(.A(n9560), .B(n9526), .Y(n9561));
  NOR2X1  g06342(.A(n9555), .B(n9554), .Y(n9562));
  NOR4X1  g06343(.A(n9462), .B(n9434), .C(n9339), .D(n9497), .Y(n9563));
  NOR3X1  g06344(.A(n9563), .B(n9262), .C(n8975), .Y(n9564));
  AOI21X1 g06345(.A0(n9547), .A1(n9445), .B0(n9564), .Y(n9565));
  NAND4X1 g06346(.A(n9551), .B(n9565), .C(n9562), .D(n9553), .Y(n9566));
  NAND2X1 g06347(.A(n9398), .B(n9275), .Y(n9567));
  INVX1   g06348(.A(n9521), .Y(n9568));
  AOI22X1 g06349(.A0(n9568), .A1(n9398), .B0(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(n9522), .Y(n9569));
  NAND4X1 g06350(.A(n9567), .B(n9482), .C(n9478), .D(n9569), .Y(n9570));
  AOI21X1 g06351(.A0(n9566), .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B0(n9570), .Y(n9571));
  INVX1   g06352(.A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .Y(n9572));
  NOR3X1  g06353(.A(n9533), .B(n8979), .C(n8720), .Y(n9573));
  INVX1   g06354(.A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .Y(n9574));
  OAI22X1 g06355(.A0(n8611), .A1(n9567), .B0(n9574), .B1(n9205), .Y(n9575));
  AOI21X1 g06356(.A0(n9573), .A1(P2_EBX_REG_1__SCAN_IN), .B0(n9575), .Y(n9576));
  OAI21X1 g06357(.A0(n9542), .A1(n9572), .B0(n9576), .Y(n9577));
  NOR2X1  g06358(.A(n9496), .B(n9442), .Y(n9578));
  AOI21X1 g06359(.A0(n9460), .A1(n9502), .B0(n8720), .Y(n9579));
  OAI21X1 g06360(.A0(n9527), .A1(n9578), .B0(n9579), .Y(n9580));
  NOR2X1  g06361(.A(n9537), .B(n9534), .Y(n9581));
  INVX1   g06362(.A(P2_REIP_REG_0__SCAN_IN), .Y(n9582));
  OAI21X1 g06363(.A0(n9567), .A1(n9582), .B0(n9513), .Y(n9583));
  AOI22X1 g06364(.A0(n9483), .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B0(n9552), .B1(n9583), .Y(n9584));
  NAND3X1 g06365(.A(n9584), .B(n9581), .C(n9580), .Y(n9585));
  NOR2X1  g06366(.A(n9500), .B(n9496), .Y(n9586));
  NOR3X1  g06367(.A(n9546), .B(n9586), .C(n9564), .Y(n9587));
  OAI21X1 g06368(.A0(n9492), .A1(n9468), .B0(n9481), .Y(n9588));
  NOR4X1  g06369(.A(n9514), .B(n9507), .C(n9554), .D(n9588), .Y(n9589));
  NOR3X1  g06370(.A(n9546), .B(n9541), .C(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n9590));
  AOI21X1 g06371(.A0(n9589), .A1(n9587), .B0(n9590), .Y(n9591));
  NAND3X1 g06372(.A(n9591), .B(n9585), .C(n9577), .Y(n9592));
  NAND2X1 g06373(.A(n9571), .B(n9577), .Y(n9593));
  OAI22X1 g06374(.A0(n9592), .A1(n9571), .B0(n9560), .B1(n9593), .Y(n9594));
  AOI21X1 g06375(.A0(n9561), .A1(n9491), .B0(n9594), .Y(n9595));
  NOR2X1  g06376(.A(n9487), .B(n8946), .Y(n9596));
  NOR4X1  g06377(.A(n8978), .B(n9336), .C(n8826), .D(n9516), .Y(n9597));
  NOR3X1  g06378(.A(n9519), .B(n9311), .C(n9470), .Y(n9598));
  NOR3X1  g06379(.A(n9598), .B(n9597), .C(n9596), .Y(n9599));
  INVX1   g06380(.A(n9599), .Y(n9600));
  XOR2X1  g06381(.A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(n8732), .Y(n9601));
  NAND4X1 g06382(.A(n8884), .B(n9470), .C(n9378), .D(n9310), .Y(n9602));
  OAI21X1 g06383(.A0(n9502), .A1(n8979), .B0(n9602), .Y(n9603));
  NOR2X1  g06384(.A(n8913), .B(n8825), .Y(n9604));
  XOR2X1  g06385(.A(n8975), .B(n8978), .Y(n9605));
  NOR4X1  g06386(.A(n9442), .B(n9339), .C(n9433), .D(n9332), .Y(n9607));
  AOI22X1 g06387(.A0(n9458), .A1(n9607), .B0(n9604), .B1(n9603), .Y(n9608));
  NOR3X1  g06388(.A(n9608), .B(n9601), .C(n8855), .Y(n9609));
  AOI21X1 g06389(.A0(n9600), .A1(n8732), .B0(n9609), .Y(n9610));
  OAI21X1 g06390(.A0(n9595), .A1(n9475), .B0(n9610), .Y(n9611));
  NAND2X1 g06391(.A(n9611), .B(n9439), .Y(n9612));
  OAI21X1 g06392(.A0(n9439), .A1(n8732), .B0(n9612), .Y(n9613));
  XOR2X1  g06393(.A(n9559), .B(n9585), .Y(n9614));
  NOR3X1  g06394(.A(n9608), .B(n8855), .C(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n9615));
  AOI21X1 g06395(.A0(n9600), .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B0(n9615), .Y(n9616));
  OAI21X1 g06396(.A0(n9614), .A1(n9475), .B0(n9616), .Y(n9617));
  AOI21X1 g06397(.A0(n9617), .A1(n9439), .B0(n9209), .Y(n9618));
  OAI21X1 g06398(.A0(n9439), .A1(n8721), .B0(n9618), .Y(n9619));
  AOI21X1 g06399(.A0(n9613), .A1(n9208), .B0(n9619), .Y(n9620));
  INVX1   g06400(.A(n9439), .Y(n9621));
  NOR3X1  g06401(.A(n9559), .B(n9545), .C(n9491), .Y(n9622));
  OAI21X1 g06402(.A0(n9559), .A1(n9545), .B0(n9491), .Y(n9623));
  AOI21X1 g06403(.A0(n9623), .A1(n9526), .B0(n9622), .Y(n9624));
  NAND2X1 g06404(.A(n9573), .B(P2_EBX_REG_2__SCAN_IN), .Y(n9625));
  AOI22X1 g06405(.A0(P2_REIP_REG_2__SCAN_IN), .A1(n9488), .B0(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(P2_STATE2_REG_1__SCAN_IN), .Y(n9626));
  NAND2X1 g06406(.A(n9626), .B(n9625), .Y(n9627));
  AOI21X1 g06407(.A0(n9483), .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B0(n9627), .Y(n9628));
  AOI21X1 g06408(.A0(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A1(n8720), .B0(P2_STATE2_REG_1__SCAN_IN), .Y(n9629));
  INVX1   g06409(.A(n9629), .Y(n9630));
  AOI21X1 g06410(.A0(n9566), .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B0(n9630), .Y(n9631));
  XOR2X1  g06411(.A(n9631), .B(n9628), .Y(n9632));
  XOR2X1  g06412(.A(n9632), .B(n9624), .Y(n9633));
  NOR2X1  g06413(.A(n9633), .B(n9475), .Y(n9634));
  XOR2X1  g06414(.A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n8727), .Y(n9635));
  NOR2X1  g06415(.A(n9635), .B(n9599), .Y(n9636));
  OAI21X1 g06416(.A0(n8721), .A1(n8732), .B0(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Y(n9637));
  NAND2X1 g06417(.A(n9637), .B(n8728), .Y(n9638));
  NOR2X1  g06418(.A(n9533), .B(n8979), .Y(n9639));
  NOR4X1  g06419(.A(n9311), .B(n8796), .C(n9433), .D(n9519), .Y(n9640));
  OAI21X1 g06420(.A0(n9640), .A1(n9639), .B0(n9638), .Y(n9641));
  NOR2X1  g06421(.A(n9401), .B(n9333), .Y(n9642));
  OAI21X1 g06422(.A0(n9642), .A1(n9638), .B0(n9641), .Y(n9643));
  NOR3X1  g06423(.A(n9643), .B(n9636), .C(n9634), .Y(n9644));
  NOR2X1  g06424(.A(n9644), .B(n9621), .Y(n9645));
  AOI21X1 g06425(.A0(n9621), .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B0(n9645), .Y(n9646));
  NAND2X1 g06426(.A(n9646), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .Y(n9647));
  OAI21X1 g06427(.A0(n9613), .A1(n9208), .B0(n9647), .Y(n9648));
  NOR2X1  g06428(.A(n9648), .B(n9620), .Y(n9649));
  NAND2X1 g06429(.A(n9483), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .Y(n9650));
  NAND3X1 g06430(.A(n9626), .B(n9625), .C(n9650), .Y(n9651));
  OAI21X1 g06431(.A0(n9515), .A1(n8727), .B0(n9629), .Y(n9652));
  NAND2X1 g06432(.A(n9652), .B(n9651), .Y(n9653));
  NOR2X1  g06433(.A(n9652), .B(n9651), .Y(n9654));
  OAI21X1 g06434(.A0(n9654), .A1(n9624), .B0(n9653), .Y(n9655));
  AOI22X1 g06435(.A0(n9566), .A1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B0(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B1(n9522), .Y(n9656));
  INVX1   g06436(.A(n9656), .Y(n9657));
  INVX1   g06437(.A(P2_EBX_REG_3__SCAN_IN), .Y(n9658));
  AOI22X1 g06438(.A0(P2_REIP_REG_3__SCAN_IN), .A1(n9488), .B0(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(P2_STATE2_REG_1__SCAN_IN), .Y(n9659));
  OAI21X1 g06439(.A0(n9485), .A1(n9658), .B0(n9659), .Y(n9660));
  AOI21X1 g06440(.A0(n9483), .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B0(n9660), .Y(n9661));
  XOR2X1  g06441(.A(n9661), .B(n9657), .Y(n9662));
  XOR2X1  g06442(.A(n9662), .B(n9655), .Y(n9663));
  XOR2X1  g06443(.A(n8777), .B(n8724), .Y(n9664));
  XOR2X1  g06444(.A(n8742), .B(n8724), .Y(n9665));
  OAI21X1 g06445(.A0(n9640), .A1(n9639), .B0(n9665), .Y(n9666));
  AOI21X1 g06446(.A0(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B0(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Y(n9667));
  XOR2X1  g06447(.A(n9667), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n9668));
  OAI21X1 g06448(.A0(n9668), .A1(n9642), .B0(n9666), .Y(n9669));
  AOI21X1 g06449(.A0(n9664), .A1(n9600), .B0(n9669), .Y(n9670));
  OAI21X1 g06450(.A0(n9663), .A1(n9475), .B0(n9670), .Y(n9671));
  NOR2X1  g06451(.A(n9439), .B(n8724), .Y(n9672));
  AOI21X1 g06452(.A0(n9671), .A1(n9439), .B0(n9672), .Y(n9673));
  OAI22X1 g06453(.A0(n9646), .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B0(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B1(n9673), .Y(n9674));
  NOR4X1  g06454(.A(n9311), .B(n9336), .C(n8826), .D(n9516), .Y(n9675));
  INVX1   g06455(.A(n9675), .Y(n9676));
  NOR2X1  g06456(.A(n8777), .B(n8724), .Y(n9677));
  NAND3X1 g06457(.A(n9022), .B(n8855), .C(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .Y(n9678));
  XOR2X1  g06458(.A(n9678), .B(n9677), .Y(n9679));
  NOR3X1  g06459(.A(n9679), .B(n9621), .C(n9676), .Y(n9680));
  AOI21X1 g06460(.A0(n9621), .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B0(n9680), .Y(n9681));
  AOI22X1 g06461(.A0(n9673), .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B0(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B1(n9681), .Y(n9682));
  OAI21X1 g06462(.A0(n9674), .A1(n9649), .B0(n9682), .Y(n9683));
  NOR2X1  g06463(.A(n9673), .B(n9646), .Y(n9684));
  NOR2X1  g06464(.A(n9681), .B(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .Y(n9685));
  INVX1   g06465(.A(n9357), .Y(n9687));
  OAI22X1 g06466(.A0(n9419), .A1(n9458), .B0(n8619), .B1(n9605), .Y(n9693));
  NOR2X1  g06467(.A(n9693), .B(n13918), .Y(n9694));
  OAI21X1 g06468(.A0(P2_MORE_REG_SCAN_IN), .A1(P2_FLUSH_REG_SCAN_IN), .B0(n9694), .Y(n9695));
  NAND2X1 g06469(.A(n9695), .B(n9681), .Y(n9696));
  NOR3X1  g06470(.A(n9696), .B(n9685), .C(n9684), .Y(n9697));
  NAND3X1 g06471(.A(n9697), .B(n9683), .C(n9408), .Y(n9698));
  NOR3X1  g06472(.A(n9698), .B(n9403), .C(P2_STATE2_REG_1__SCAN_IN), .Y(n9699));
  INVX1   g06473(.A(P2_STATE2_REG_2__SCAN_IN), .Y(n9700));
  AOI21X1 g06474(.A0(READY21_REG_SCAN_IN), .A1(READY12_REG_SCAN_IN), .B0(P2_STATEBS16_REG_SCAN_IN), .Y(n9701));
  INVX1   g06475(.A(n9701), .Y(n9702));
  NOR4X1  g06476(.A(n9539), .B(n9487), .C(P2_STATE_REG_0__SCAN_IN), .D(n9702), .Y(n9703));
  AOI21X1 g06477(.A0(READY21_REG_SCAN_IN), .A1(READY12_REG_SCAN_IN), .B0(P2_STATE2_REG_0__SCAN_IN), .Y(n9704));
  NOR4X1  g06478(.A(n9703), .B(n9522), .C(n9700), .D(n9704), .Y(n9705));
  AOI21X1 g06479(.A0(n9705), .A1(n9699), .B0(n8720), .Y(n9706));
  NOR2X1  g06480(.A(n9698), .B(n9403), .Y(n9707));
  NAND3X1 g06481(.A(P2_STATE2_REG_0__SCAN_IN), .B(P2_STATE2_REG_1__SCAN_IN), .C(P2_STATE2_REG_2__SCAN_IN), .Y(n9708));
  OAI21X1 g06482(.A0(n9706), .A1(n8719), .B0(n9708), .Y(P2_U3593));
  INVX1   g06483(.A(P2_STATEBS16_REG_SCAN_IN), .Y(n9710));
  NOR2X1  g06484(.A(n8720), .B(P2_STATE2_REG_2__SCAN_IN), .Y(n9711));
  OAI21X1 g06485(.A0(n8616), .A1(n8615), .B0(n9711), .Y(n9712));
  OAI21X1 g06486(.A0(n9710), .A1(P2_STATE2_REG_0__SCAN_IN), .B0(n9712), .Y(n9713));
  NOR2X1  g06487(.A(P2_STATE2_REG_1__SCAN_IN), .B(n9700), .Y(n9714));
  AOI21X1 g06488(.A0(n9713), .A1(P2_STATE2_REG_1__SCAN_IN), .B0(n9714), .Y(n9715));
  OAI21X1 g06489(.A0(n9706), .A1(n9700), .B0(n9715), .Y(P2_U3178));
  NOR2X1  g06490(.A(P2_STATE2_REG_1__SCAN_IN), .B(P2_STATE2_REG_3__SCAN_IN), .Y(n9717));
  NAND3X1 g06491(.A(n9717), .B(n9706), .C(n8620), .Y(n9718));
  OAI21X1 g06492(.A0(n9699), .A1(n8720), .B0(n9705), .Y(n9719));
  INVX1   g06493(.A(n9719), .Y(n9720));
  NOR4X1  g06494(.A(P2_STATE2_REG_2__SCAN_IN), .B(n8616), .C(n8615), .D(n8720), .Y(n9721));
  OAI21X1 g06495(.A0(n9721), .A1(n9720), .B0(P2_STATE2_REG_1__SCAN_IN), .Y(n9722));
  NOR4X1  g06496(.A(P2_STATE2_REG_0__SCAN_IN), .B(n9205), .C(P2_STATE2_REG_2__SCAN_IN), .D(P2_STATEBS16_REG_SCAN_IN), .Y(n9723));
  NOR3X1  g06497(.A(n8720), .B(P2_STATE2_REG_1__SCAN_IN), .C(n9700), .Y(n9724));
  AOI21X1 g06498(.A0(n9724), .A1(n9719), .B0(n9723), .Y(n9725));
  NAND3X1 g06499(.A(n9725), .B(n9722), .C(n9718), .Y(P2_U3177));
  NOR4X1  g06500(.A(n9248), .B(n9205), .C(n9700), .D(n9258), .Y(n9727));
  OAI21X1 g06501(.A0(n9727), .A1(n9720), .B0(P2_STATE2_REG_0__SCAN_IN), .Y(n9728));
  NOR2X1  g06502(.A(P2_STATE2_REG_1__SCAN_IN), .B(P2_STATE2_REG_2__SCAN_IN), .Y(n9729));
  AOI21X1 g06503(.A0(n9307), .A1(n9304), .B0(n8719), .Y(n9730));
  AOI21X1 g06504(.A0(n9730), .A1(n9729), .B0(P2_STATE2_REG_0__SCAN_IN), .Y(n9731));
  INVX1   g06505(.A(n9724), .Y(n9732));
  NOR4X1  g06506(.A(P2_STATE2_REG_1__SCAN_IN), .B(P2_STATE2_REG_2__SCAN_IN), .C(n8719), .D(n8720), .Y(n9733));
  NOR2X1  g06507(.A(n9733), .B(n9721), .Y(n9734));
  OAI21X1 g06508(.A0(n9732), .A1(n9707), .B0(n9734), .Y(n9735));
  AOI21X1 g06509(.A0(n9731), .A1(n9719), .B0(n9735), .Y(n9736));
  NAND2X1 g06510(.A(n9736), .B(n9728), .Y(P2_U3176));
  INVX1   g06511(.A(n9730), .Y(n9738));
  XOR2X1  g06512(.A(P2_STATE2_REG_1__SCAN_IN), .B(n9700), .Y(n9739));
  AOI21X1 g06513(.A0(n9739), .A1(n9738), .B0(P2_STATE2_REG_0__SCAN_IN), .Y(n9740));
  INVX1   g06514(.A(BUF1_REG_7__SCAN_IN), .Y(n9741));
  NOR2X1  g06515(.A(n3086), .B(n9741), .Y(n9742));
  AOI21X1 g06516(.A0(n3086), .A1(BUF2_REG_7__SCAN_IN), .B0(n9742), .Y(n9743));
  INVX1   g06517(.A(n9743), .Y(n9744));
  NAND2X1 g06518(.A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Y(n9745));
  NOR3X1  g06519(.A(n9745), .B(n9223), .C(n9221), .Y(n9746));
  XOR2X1  g06520(.A(n9560), .B(n9571), .Y(n9747));
  NAND2X1 g06521(.A(n9591), .B(n9585), .Y(n9748));
  NOR2X1  g06522(.A(n9526), .B(n9491), .Y(n9749));
  AOI22X1 g06523(.A0(n9622), .A1(n9526), .B0(n9748), .B1(n9749), .Y(n9750));
  OAI21X1 g06524(.A0(n9747), .A1(n9577), .B0(n9750), .Y(n9751));
  XOR2X1  g06525(.A(n9559), .B(n9545), .Y(n9752));
  NAND2X1 g06526(.A(n9752), .B(n9751), .Y(n9753));
  NOR3X1  g06527(.A(n9753), .B(n9663), .C(n9633), .Y(n9754));
  OAI21X1 g06528(.A0(n9754), .A1(n9746), .B0(P2_STATE2_REG_2__SCAN_IN), .Y(n9755));
  NAND3X1 g06529(.A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .Y(n9756));
  NOR3X1  g06530(.A(P2_STATEBS16_REG_SCAN_IN), .B(P2_STATE2_REG_2__SCAN_IN), .C(P2_STATE2_REG_3__SCAN_IN), .Y(n9757));
  NOR3X1  g06531(.A(n9710), .B(P2_STATE2_REG_2__SCAN_IN), .C(P2_STATE2_REG_3__SCAN_IN), .Y(n9758));
  INVX1   g06532(.A(n9758), .Y(n9759));
  NAND4X1 g06533(.A(n9331), .B(n9322), .C(P2_STATE2_REG_0__SCAN_IN), .D(n8975), .Y(n9760));
  NOR2X1  g06534(.A(n9760), .B(n9099), .Y(n9761));
  NAND3X1 g06535(.A(P2_STATE2_REG_0__SCAN_IN), .B(P2_STATE2_REG_2__SCAN_IN), .C(n8719), .Y(n9762));
  NOR3X1  g06536(.A(n9762), .B(n9761), .C(n8796), .Y(n9763));
  INVX1   g06537(.A(n9763), .Y(n9764));
  NOR2X1  g06538(.A(P2_STATE2_REG_0__SCAN_IN), .B(n9700), .Y(n9765));
  NOR2X1  g06539(.A(P2_STATE2_REG_2__SCAN_IN), .B(P2_STATE2_REG_3__SCAN_IN), .Y(n9766));
  INVX1   g06540(.A(n9766), .Y(n9767));
  AOI21X1 g06541(.A0(n8796), .A1(P2_STATE2_REG_0__SCAN_IN), .B0(P2_STATE2_REG_3__SCAN_IN), .Y(n9768));
  OAI22X1 g06542(.A0(n9767), .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B0(n8721), .B1(n9768), .Y(n9769));
  AOI21X1 g06543(.A0(n9765), .A1(n9752), .B0(n9769), .Y(n9770));
  XOR2X1  g06544(.A(n9770), .B(n9764), .Y(n9771));
  INVX1   g06545(.A(n9771), .Y(n9772));
  NOR2X1  g06546(.A(n9760), .B(n9070), .Y(n9773));
  INVX1   g06547(.A(n9765), .Y(n9774));
  INVX1   g06548(.A(n9769), .Y(n9775));
  OAI21X1 g06549(.A0(n9774), .A1(n9614), .B0(n9775), .Y(n9776));
  XOR2X1  g06550(.A(n9770), .B(n9773), .Y(n9778));
  XOR2X1  g06551(.A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n9208), .Y(n9779));
  INVX1   g06552(.A(n9779), .Y(n9780));
  INVX1   g06553(.A(n9768), .Y(n9781));
  AOI22X1 g06554(.A0(n9766), .A1(n9780), .B0(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(n9781), .Y(n9782));
  OAI21X1 g06555(.A0(n9774), .A1(n9595), .B0(n9782), .Y(n9783));
  XOR2X1  g06556(.A(n9783), .B(n9778), .Y(n9784));
  INVX1   g06557(.A(n9760), .Y(n9785));
  XOR2X1  g06558(.A(n9745), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .Y(n9786));
  INVX1   g06559(.A(n9786), .Y(n9787));
  AOI22X1 g06560(.A0(n9766), .A1(n9787), .B0(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(n9781), .Y(n9788));
  OAI21X1 g06561(.A0(n9774), .A1(n9633), .B0(n9788), .Y(n9789));
  AOI21X1 g06562(.A0(n9785), .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B0(n9789), .Y(n9790));
  INVX1   g06563(.A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .Y(n9791));
  AOI21X1 g06564(.A0(n9591), .A1(n9585), .B0(n9577), .Y(n9792));
  OAI21X1 g06565(.A0(n9792), .A1(n9571), .B0(n9592), .Y(n9793));
  XOR2X1  g06566(.A(n9632), .B(n9793), .Y(n9794));
  INVX1   g06567(.A(n9788), .Y(n9795));
  AOI21X1 g06568(.A0(n9765), .A1(n9794), .B0(n9795), .Y(n9796));
  NOR3X1  g06569(.A(n9796), .B(n9760), .C(n9791), .Y(n9797));
  OAI22X1 g06570(.A0(n9763), .A1(n9770), .B0(n9760), .B1(n9070), .Y(n9798));
  NOR4X1  g06571(.A(n9763), .B(n9760), .C(n9070), .D(n9770), .Y(n9799));
  OAI21X1 g06572(.A0(n9799), .A1(n9783), .B0(n9798), .Y(n9800));
  NOR3X1  g06573(.A(n9800), .B(n9797), .C(n9790), .Y(n9801));
  AOI21X1 g06574(.A0(n9785), .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B0(n9796), .Y(n9802));
  NOR3X1  g06575(.A(n9789), .B(n9760), .C(n9791), .Y(n9803));
  INVX1   g06576(.A(n9782), .Y(n9804));
  AOI21X1 g06577(.A0(n9765), .A1(n9751), .B0(n9804), .Y(n9805));
  AOI21X1 g06578(.A0(n9776), .A1(n9764), .B0(n9773), .Y(n9806));
  NAND3X1 g06579(.A(n9773), .B(n9776), .C(n9764), .Y(n9807));
  OAI21X1 g06580(.A0(n9806), .A1(n9805), .B0(n9807), .Y(n9808));
  NOR3X1  g06581(.A(n9808), .B(n9803), .C(n9802), .Y(n9809));
  NOR2X1  g06582(.A(n9809), .B(n9801), .Y(n9810));
  INVX1   g06583(.A(n9810), .Y(n9811));
  NAND3X1 g06584(.A(n9789), .B(n9785), .C(P2_INSTQUEUE_REG_0__2__SCAN_IN), .Y(n9812));
  OAI21X1 g06585(.A0(n9800), .A1(n9790), .B0(n9812), .Y(n9813));
  XOR2X1  g06586(.A(n9661), .B(n9656), .Y(n9814));
  XOR2X1  g06587(.A(n9814), .B(n9655), .Y(n9815));
  AOI21X1 g06588(.A0(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B0(n9221), .Y(n9816));
  NOR3X1  g06589(.A(n9745), .B(n9223), .C(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .Y(n9817));
  NOR2X1  g06590(.A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n9221), .Y(n9818));
  NOR3X1  g06591(.A(n9818), .B(n9817), .C(n9816), .Y(n9819));
  INVX1   g06592(.A(n9819), .Y(n9820));
  AOI22X1 g06593(.A0(n9766), .A1(n9820), .B0(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(n9781), .Y(n9821));
  INVX1   g06594(.A(n9821), .Y(n9822));
  AOI21X1 g06595(.A0(n9765), .A1(n9815), .B0(n9822), .Y(n9823));
  INVX1   g06596(.A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .Y(n9824));
  NOR2X1  g06597(.A(n9760), .B(n9824), .Y(n9825));
  XOR2X1  g06598(.A(n9825), .B(n9823), .Y(n9826));
  XOR2X1  g06599(.A(n9826), .B(n9813), .Y(n9827));
  NOR4X1  g06600(.A(n9811), .B(n9784), .C(n9772), .D(n9827), .Y(n9828));
  NOR2X1  g06601(.A(n9784), .B(n9771), .Y(n9829));
  INVX1   g06602(.A(n9829), .Y(n9830));
  NOR4X1  g06603(.A(n9809), .B(n9801), .C(n9830), .D(n9827), .Y(n9831));
  NOR3X1  g06604(.A(n9831), .B(n9828), .C(n9759), .Y(n9832));
  NOR2X1  g06605(.A(n9832), .B(n9757), .Y(n9833));
  OAI21X1 g06606(.A0(n9833), .A1(n9756), .B0(n9755), .Y(n9834));
  NAND3X1 g06607(.A(n9834), .B(n9744), .C(n9740), .Y(n9835));
  INVX1   g06608(.A(n9740), .Y(n9836));
  NOR4X1  g06609(.A(n9828), .B(n9759), .C(n9836), .D(n9831), .Y(n9837));
  OAI21X1 g06610(.A0(n9837), .A1(n9757), .B0(n9756), .Y(n9838));
  INVX1   g06611(.A(n9746), .Y(n9839));
  NOR3X1  g06612(.A(n9754), .B(n9746), .C(n9700), .Y(n9840));
  AOI21X1 g06613(.A0(n9839), .A1(P2_STATE2_REG_3__SCAN_IN), .B0(n9840), .Y(n9841));
  NAND3X1 g06614(.A(n9841), .B(n9838), .C(n9740), .Y(n9842));
  NAND2X1 g06615(.A(n9842), .B(P2_INSTQUEUE_REG_15__7__SCAN_IN), .Y(n9843));
  INVX1   g06616(.A(BUF1_REG_31__SCAN_IN), .Y(n9844));
  NOR2X1  g06617(.A(n3086), .B(n9844), .Y(n9845));
  AOI21X1 g06618(.A0(n3086), .A1(BUF2_REG_31__SCAN_IN), .B0(n9845), .Y(n9846));
  NOR3X1  g06619(.A(n9846), .B(n9759), .C(n9836), .Y(n9847));
  INVX1   g06620(.A(n9831), .Y(n9848));
  INVX1   g06621(.A(BUF1_REG_23__SCAN_IN), .Y(n9849));
  NOR2X1  g06622(.A(n3086), .B(n9849), .Y(n9850));
  AOI21X1 g06623(.A0(n3086), .A1(BUF2_REG_23__SCAN_IN), .B0(n9850), .Y(n9851));
  INVX1   g06624(.A(n9851), .Y(n9852));
  NAND3X1 g06625(.A(n9852), .B(n9758), .C(n9740), .Y(n9853));
  NAND3X1 g06626(.A(n9740), .B(n8884), .C(P2_STATE2_REG_3__SCAN_IN), .Y(n9854));
  OAI22X1 g06627(.A0(n9853), .A1(n9848), .B0(n9839), .B1(n9854), .Y(n9855));
  AOI21X1 g06628(.A0(n9847), .A1(n9828), .B0(n9855), .Y(n9856));
  NAND3X1 g06629(.A(n9856), .B(n9843), .C(n9835), .Y(P2_U3175));
  INVX1   g06630(.A(BUF1_REG_6__SCAN_IN), .Y(n9858));
  NOR2X1  g06631(.A(n3086), .B(n9858), .Y(n9859));
  AOI21X1 g06632(.A0(n3086), .A1(BUF2_REG_6__SCAN_IN), .B0(n9859), .Y(n9860));
  INVX1   g06633(.A(n9860), .Y(n9861));
  NAND3X1 g06634(.A(n9861), .B(n9834), .C(n9740), .Y(n9862));
  NAND2X1 g06635(.A(n9842), .B(P2_INSTQUEUE_REG_15__6__SCAN_IN), .Y(n9863));
  INVX1   g06636(.A(BUF1_REG_30__SCAN_IN), .Y(n9864));
  NOR2X1  g06637(.A(n3086), .B(n9864), .Y(n9865));
  AOI21X1 g06638(.A0(n3086), .A1(BUF2_REG_30__SCAN_IN), .B0(n9865), .Y(n9866));
  NOR3X1  g06639(.A(n9866), .B(n9759), .C(n9836), .Y(n9867));
  INVX1   g06640(.A(BUF1_REG_22__SCAN_IN), .Y(n9868));
  NOR2X1  g06641(.A(n3086), .B(n9868), .Y(n9869));
  AOI21X1 g06642(.A0(n3086), .A1(BUF2_REG_22__SCAN_IN), .B0(n9869), .Y(n9870));
  INVX1   g06643(.A(n9870), .Y(n9871));
  NAND3X1 g06644(.A(n9871), .B(n9758), .C(n9740), .Y(n9872));
  NAND3X1 g06645(.A(n9740), .B(n8796), .C(P2_STATE2_REG_3__SCAN_IN), .Y(n9873));
  OAI22X1 g06646(.A0(n9872), .A1(n9848), .B0(n9839), .B1(n9873), .Y(n9874));
  AOI21X1 g06647(.A0(n9867), .A1(n9828), .B0(n9874), .Y(n9875));
  NAND3X1 g06648(.A(n9875), .B(n9863), .C(n9862), .Y(P2_U3174));
  INVX1   g06649(.A(BUF1_REG_5__SCAN_IN), .Y(n9877));
  NOR2X1  g06650(.A(n3086), .B(n9877), .Y(n9878));
  AOI21X1 g06651(.A0(n3086), .A1(BUF2_REG_5__SCAN_IN), .B0(n9878), .Y(n9879));
  INVX1   g06652(.A(n9879), .Y(n9880));
  NAND3X1 g06653(.A(n9880), .B(n9834), .C(n9740), .Y(n9881));
  NAND2X1 g06654(.A(n9842), .B(P2_INSTQUEUE_REG_15__5__SCAN_IN), .Y(n9882));
  INVX1   g06655(.A(BUF1_REG_29__SCAN_IN), .Y(n9883));
  NOR2X1  g06656(.A(n3086), .B(n9883), .Y(n9884));
  AOI21X1 g06657(.A0(n3086), .A1(BUF2_REG_29__SCAN_IN), .B0(n9884), .Y(n9885));
  NOR3X1  g06658(.A(n9885), .B(n9759), .C(n9836), .Y(n9886));
  INVX1   g06659(.A(BUF1_REG_21__SCAN_IN), .Y(n9887));
  NOR2X1  g06660(.A(n3086), .B(n9887), .Y(n9888));
  AOI21X1 g06661(.A0(n3086), .A1(BUF2_REG_21__SCAN_IN), .B0(n9888), .Y(n9889));
  INVX1   g06662(.A(n9889), .Y(n9890));
  NAND3X1 g06663(.A(n9890), .B(n9758), .C(n9740), .Y(n9891));
  NAND3X1 g06664(.A(n9740), .B(n8825), .C(P2_STATE2_REG_3__SCAN_IN), .Y(n9892));
  OAI22X1 g06665(.A0(n9891), .A1(n9848), .B0(n9839), .B1(n9892), .Y(n9893));
  AOI21X1 g06666(.A0(n9886), .A1(n9828), .B0(n9893), .Y(n9894));
  NAND3X1 g06667(.A(n9894), .B(n9882), .C(n9881), .Y(P2_U3173));
  INVX1   g06668(.A(BUF1_REG_4__SCAN_IN), .Y(n9896));
  NOR2X1  g06669(.A(n3086), .B(n9896), .Y(n9897));
  AOI21X1 g06670(.A0(n3086), .A1(BUF2_REG_4__SCAN_IN), .B0(n9897), .Y(n9898));
  INVX1   g06671(.A(n9898), .Y(n9899));
  NAND3X1 g06672(.A(n9899), .B(n9834), .C(n9740), .Y(n9900));
  NAND2X1 g06673(.A(n9842), .B(P2_INSTQUEUE_REG_15__4__SCAN_IN), .Y(n9901));
  INVX1   g06674(.A(BUF1_REG_28__SCAN_IN), .Y(n9902));
  NOR2X1  g06675(.A(n3086), .B(n9902), .Y(n9903));
  AOI21X1 g06676(.A0(n3086), .A1(BUF2_REG_28__SCAN_IN), .B0(n9903), .Y(n9904));
  NOR3X1  g06677(.A(n9904), .B(n9759), .C(n9836), .Y(n9905));
  INVX1   g06678(.A(BUF1_REG_20__SCAN_IN), .Y(n9906));
  NOR2X1  g06679(.A(n3086), .B(n9906), .Y(n9907));
  AOI21X1 g06680(.A0(n3086), .A1(BUF2_REG_20__SCAN_IN), .B0(n9907), .Y(n9908));
  INVX1   g06681(.A(n9908), .Y(n9909));
  NAND3X1 g06682(.A(n9909), .B(n9758), .C(n9740), .Y(n9910));
  NAND3X1 g06683(.A(n9740), .B(n9378), .C(P2_STATE2_REG_3__SCAN_IN), .Y(n9911));
  OAI22X1 g06684(.A0(n9910), .A1(n9848), .B0(n9839), .B1(n9911), .Y(n9912));
  AOI21X1 g06685(.A0(n9905), .A1(n9828), .B0(n9912), .Y(n9913));
  NAND3X1 g06686(.A(n9913), .B(n9901), .C(n9900), .Y(P2_U3172));
  INVX1   g06687(.A(BUF1_REG_3__SCAN_IN), .Y(n9915));
  NOR2X1  g06688(.A(n3086), .B(n9915), .Y(n9916));
  AOI21X1 g06689(.A0(n3086), .A1(BUF2_REG_3__SCAN_IN), .B0(n9916), .Y(n9917));
  INVX1   g06690(.A(n9917), .Y(n9918));
  NAND3X1 g06691(.A(n9918), .B(n9834), .C(n9740), .Y(n9919));
  NAND2X1 g06692(.A(n9842), .B(P2_INSTQUEUE_REG_15__3__SCAN_IN), .Y(n9920));
  INVX1   g06693(.A(BUF1_REG_27__SCAN_IN), .Y(n9921));
  NOR2X1  g06694(.A(n3086), .B(n9921), .Y(n9922));
  AOI21X1 g06695(.A0(n3086), .A1(BUF2_REG_27__SCAN_IN), .B0(n9922), .Y(n9923));
  NOR3X1  g06696(.A(n9923), .B(n9759), .C(n9836), .Y(n9924));
  INVX1   g06697(.A(BUF1_REG_19__SCAN_IN), .Y(n9925));
  NOR2X1  g06698(.A(n3086), .B(n9925), .Y(n9926));
  AOI21X1 g06699(.A0(n3086), .A1(BUF2_REG_19__SCAN_IN), .B0(n9926), .Y(n9927));
  INVX1   g06700(.A(n9927), .Y(n9928));
  NAND3X1 g06701(.A(n9928), .B(n9758), .C(n9740), .Y(n9929));
  NAND3X1 g06702(.A(n9740), .B(n8913), .C(P2_STATE2_REG_3__SCAN_IN), .Y(n9930));
  OAI22X1 g06703(.A0(n9929), .A1(n9848), .B0(n9839), .B1(n9930), .Y(n9931));
  AOI21X1 g06704(.A0(n9924), .A1(n9828), .B0(n9931), .Y(n9932));
  NAND3X1 g06705(.A(n9932), .B(n9920), .C(n9919), .Y(P2_U3171));
  INVX1   g06706(.A(BUF1_REG_2__SCAN_IN), .Y(n9934));
  NOR2X1  g06707(.A(n3086), .B(n9934), .Y(n9935));
  AOI21X1 g06708(.A0(n3086), .A1(BUF2_REG_2__SCAN_IN), .B0(n9935), .Y(n9936));
  INVX1   g06709(.A(n9936), .Y(n9937));
  NAND3X1 g06710(.A(n9937), .B(n9834), .C(n9740), .Y(n9938));
  NAND2X1 g06711(.A(n9842), .B(P2_INSTQUEUE_REG_15__2__SCAN_IN), .Y(n9939));
  INVX1   g06712(.A(BUF1_REG_26__SCAN_IN), .Y(n9940));
  NOR2X1  g06713(.A(n3086), .B(n9940), .Y(n9941));
  AOI21X1 g06714(.A0(n3086), .A1(BUF2_REG_26__SCAN_IN), .B0(n9941), .Y(n9942));
  NOR3X1  g06715(.A(n9942), .B(n9759), .C(n9836), .Y(n9943));
  INVX1   g06716(.A(BUF1_REG_18__SCAN_IN), .Y(n9944));
  NOR2X1  g06717(.A(n3086), .B(n9944), .Y(n9945));
  AOI21X1 g06718(.A0(n3086), .A1(BUF2_REG_18__SCAN_IN), .B0(n9945), .Y(n9946));
  INVX1   g06719(.A(n9946), .Y(n9947));
  NAND3X1 g06720(.A(n9947), .B(n9758), .C(n9740), .Y(n9948));
  NAND3X1 g06721(.A(n9740), .B(n8855), .C(P2_STATE2_REG_3__SCAN_IN), .Y(n9949));
  OAI22X1 g06722(.A0(n9948), .A1(n9848), .B0(n9839), .B1(n9949), .Y(n9950));
  AOI21X1 g06723(.A0(n9943), .A1(n9828), .B0(n9950), .Y(n9951));
  NAND3X1 g06724(.A(n9951), .B(n9939), .C(n9938), .Y(P2_U3170));
  INVX1   g06725(.A(BUF1_REG_1__SCAN_IN), .Y(n9953));
  NOR2X1  g06726(.A(n3086), .B(n9953), .Y(n9954));
  AOI21X1 g06727(.A0(n3086), .A1(BUF2_REG_1__SCAN_IN), .B0(n9954), .Y(n9955));
  INVX1   g06728(.A(n9955), .Y(n9956));
  NAND3X1 g06729(.A(n9956), .B(n9834), .C(n9740), .Y(n9957));
  NAND2X1 g06730(.A(n9842), .B(P2_INSTQUEUE_REG_15__1__SCAN_IN), .Y(n9958));
  INVX1   g06731(.A(BUF1_REG_25__SCAN_IN), .Y(n9959));
  NOR2X1  g06732(.A(n3086), .B(n9959), .Y(n9960));
  AOI21X1 g06733(.A0(n3086), .A1(BUF2_REG_25__SCAN_IN), .B0(n9960), .Y(n9961));
  NOR3X1  g06734(.A(n9961), .B(n9759), .C(n9836), .Y(n9962));
  INVX1   g06735(.A(BUF1_REG_17__SCAN_IN), .Y(n9963));
  NOR2X1  g06736(.A(n3086), .B(n9963), .Y(n9964));
  AOI21X1 g06737(.A0(n3086), .A1(BUF2_REG_17__SCAN_IN), .B0(n9964), .Y(n9965));
  INVX1   g06738(.A(n9965), .Y(n9966));
  NAND3X1 g06739(.A(n9966), .B(n9758), .C(n9740), .Y(n9967));
  NAND3X1 g06740(.A(n9740), .B(n8975), .C(P2_STATE2_REG_3__SCAN_IN), .Y(n9968));
  OAI22X1 g06741(.A0(n9967), .A1(n9848), .B0(n9839), .B1(n9968), .Y(n9969));
  AOI21X1 g06742(.A0(n9962), .A1(n9828), .B0(n9969), .Y(n9970));
  NAND3X1 g06743(.A(n9970), .B(n9958), .C(n9957), .Y(P2_U3169));
  INVX1   g06744(.A(BUF1_REG_0__SCAN_IN), .Y(n9972));
  NOR2X1  g06745(.A(n3086), .B(n9972), .Y(n9973));
  AOI21X1 g06746(.A0(n3086), .A1(BUF2_REG_0__SCAN_IN), .B0(n9973), .Y(n9974));
  INVX1   g06747(.A(n9974), .Y(n9975));
  NAND3X1 g06748(.A(n9975), .B(n9834), .C(n9740), .Y(n9976));
  NAND2X1 g06749(.A(n9842), .B(P2_INSTQUEUE_REG_15__0__SCAN_IN), .Y(n9977));
  INVX1   g06750(.A(BUF1_REG_24__SCAN_IN), .Y(n9978));
  NOR2X1  g06751(.A(n3086), .B(n9978), .Y(n9979));
  AOI21X1 g06752(.A0(n3086), .A1(BUF2_REG_24__SCAN_IN), .B0(n9979), .Y(n9980));
  NOR3X1  g06753(.A(n9980), .B(n9759), .C(n9836), .Y(n9981));
  INVX1   g06754(.A(BUF1_REG_16__SCAN_IN), .Y(n9982));
  NOR2X1  g06755(.A(n3086), .B(n9982), .Y(n9983));
  AOI21X1 g06756(.A0(n3086), .A1(BUF2_REG_16__SCAN_IN), .B0(n9983), .Y(n9984));
  INVX1   g06757(.A(n9984), .Y(n9985));
  NAND3X1 g06758(.A(n9985), .B(n9758), .C(n9740), .Y(n9986));
  NAND3X1 g06759(.A(n9740), .B(n8978), .C(P2_STATE2_REG_3__SCAN_IN), .Y(n9987));
  OAI22X1 g06760(.A0(n9986), .A1(n9848), .B0(n9839), .B1(n9987), .Y(n9988));
  AOI21X1 g06761(.A0(n9981), .A1(n9828), .B0(n9988), .Y(n9989));
  NAND3X1 g06762(.A(n9989), .B(n9977), .C(n9976), .Y(P2_U3168));
  NOR4X1  g06763(.A(n9208), .B(n9223), .C(n9221), .D(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Y(n9991));
  NAND2X1 g06764(.A(n9614), .B(n9751), .Y(n9992));
  NOR3X1  g06765(.A(n9992), .B(n9663), .C(n9633), .Y(n9993));
  OAI21X1 g06766(.A0(n9993), .A1(n9991), .B0(P2_STATE2_REG_2__SCAN_IN), .Y(n9994));
  NOR3X1  g06767(.A(n9779), .B(n9819), .C(n9786), .Y(n9995));
  XOR2X1  g06768(.A(n9805), .B(n9778), .Y(n9996));
  NOR4X1  g06769(.A(n9811), .B(n9996), .C(n9771), .D(n9827), .Y(n9997));
  NOR3X1  g06770(.A(n9828), .B(n9997), .C(n9759), .Y(n9999));
  OAI21X1 g06771(.A0(n9999), .A1(n9757), .B0(n9995), .Y(n10000));
  NAND2X1 g06772(.A(n10000), .B(n9994), .Y(n10001));
  NAND3X1 g06773(.A(n10001), .B(n9744), .C(n9740), .Y(n10002));
  NOR2X1  g06774(.A(n9819), .B(n9786), .Y(n10003));
  INVX1   g06775(.A(n10003), .Y(n10004));
  NOR4X1  g06776(.A(n9997), .B(n9759), .C(n9836), .D(n9828), .Y(n10005));
  OAI22X1 g06777(.A0(n9757), .A1(n10005), .B0(n9779), .B1(n10004), .Y(n10006));
  INVX1   g06778(.A(n9991), .Y(n10007));
  NOR3X1  g06779(.A(n9993), .B(n9991), .C(n9700), .Y(n10008));
  AOI21X1 g06780(.A0(n10007), .A1(P2_STATE2_REG_3__SCAN_IN), .B0(n10008), .Y(n10009));
  NAND3X1 g06781(.A(n10009), .B(n10006), .C(n9740), .Y(n10010));
  NAND2X1 g06782(.A(n10010), .B(P2_INSTQUEUE_REG_14__7__SCAN_IN), .Y(n10011));
  INVX1   g06783(.A(n9828), .Y(n10012));
  OAI22X1 g06784(.A0(n10007), .A1(n9854), .B0(n9853), .B1(n10012), .Y(n10013));
  AOI21X1 g06785(.A0(n9997), .A1(n9847), .B0(n10013), .Y(n10014));
  NAND3X1 g06786(.A(n10014), .B(n10011), .C(n10002), .Y(P2_U3167));
  NAND3X1 g06787(.A(n10001), .B(n9861), .C(n9740), .Y(n10016));
  NAND2X1 g06788(.A(n10010), .B(P2_INSTQUEUE_REG_14__6__SCAN_IN), .Y(n10017));
  OAI22X1 g06789(.A0(n10007), .A1(n9873), .B0(n9872), .B1(n10012), .Y(n10018));
  AOI21X1 g06790(.A0(n9997), .A1(n9867), .B0(n10018), .Y(n10019));
  NAND3X1 g06791(.A(n10019), .B(n10017), .C(n10016), .Y(P2_U3166));
  NAND3X1 g06792(.A(n10001), .B(n9880), .C(n9740), .Y(n10021));
  NAND2X1 g06793(.A(n10010), .B(P2_INSTQUEUE_REG_14__5__SCAN_IN), .Y(n10022));
  OAI22X1 g06794(.A0(n10007), .A1(n9892), .B0(n9891), .B1(n10012), .Y(n10023));
  AOI21X1 g06795(.A0(n9997), .A1(n9886), .B0(n10023), .Y(n10024));
  NAND3X1 g06796(.A(n10024), .B(n10022), .C(n10021), .Y(P2_U3165));
  NAND3X1 g06797(.A(n10001), .B(n9899), .C(n9740), .Y(n10026));
  NAND2X1 g06798(.A(n10010), .B(P2_INSTQUEUE_REG_14__4__SCAN_IN), .Y(n10027));
  OAI22X1 g06799(.A0(n10007), .A1(n9911), .B0(n9910), .B1(n10012), .Y(n10028));
  AOI21X1 g06800(.A0(n9997), .A1(n9905), .B0(n10028), .Y(n10029));
  NAND3X1 g06801(.A(n10029), .B(n10027), .C(n10026), .Y(P2_U3164));
  NAND3X1 g06802(.A(n10001), .B(n9918), .C(n9740), .Y(n10031));
  NAND2X1 g06803(.A(n10010), .B(P2_INSTQUEUE_REG_14__3__SCAN_IN), .Y(n10032));
  OAI22X1 g06804(.A0(n10007), .A1(n9930), .B0(n9929), .B1(n10012), .Y(n10033));
  AOI21X1 g06805(.A0(n9997), .A1(n9924), .B0(n10033), .Y(n10034));
  NAND3X1 g06806(.A(n10034), .B(n10032), .C(n10031), .Y(P2_U3163));
  NAND3X1 g06807(.A(n10001), .B(n9937), .C(n9740), .Y(n10036));
  NAND2X1 g06808(.A(n10010), .B(P2_INSTQUEUE_REG_14__2__SCAN_IN), .Y(n10037));
  OAI22X1 g06809(.A0(n10007), .A1(n9949), .B0(n9948), .B1(n10012), .Y(n10038));
  AOI21X1 g06810(.A0(n9997), .A1(n9943), .B0(n10038), .Y(n10039));
  NAND3X1 g06811(.A(n10039), .B(n10037), .C(n10036), .Y(P2_U3162));
  NAND3X1 g06812(.A(n10001), .B(n9956), .C(n9740), .Y(n10041));
  NAND2X1 g06813(.A(n10010), .B(P2_INSTQUEUE_REG_14__1__SCAN_IN), .Y(n10042));
  OAI22X1 g06814(.A0(n10007), .A1(n9968), .B0(n9967), .B1(n10012), .Y(n10043));
  AOI21X1 g06815(.A0(n9997), .A1(n9962), .B0(n10043), .Y(n10044));
  NAND3X1 g06816(.A(n10044), .B(n10042), .C(n10041), .Y(P2_U3161));
  NAND3X1 g06817(.A(n10001), .B(n9975), .C(n9740), .Y(n10046));
  NAND2X1 g06818(.A(n10010), .B(P2_INSTQUEUE_REG_14__0__SCAN_IN), .Y(n10047));
  OAI22X1 g06819(.A0(n10007), .A1(n9987), .B0(n9986), .B1(n10012), .Y(n10048));
  AOI21X1 g06820(.A0(n9997), .A1(n9981), .B0(n10048), .Y(n10049));
  NAND3X1 g06821(.A(n10049), .B(n10047), .C(n10046), .Y(P2_U3160));
  NOR4X1  g06822(.A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n9223), .C(n9221), .D(n9209), .Y(n10051));
  NAND2X1 g06823(.A(n9752), .B(n9595), .Y(n10052));
  NOR3X1  g06824(.A(n10052), .B(n9663), .C(n9633), .Y(n10053));
  OAI21X1 g06825(.A0(n10053), .A1(n10051), .B0(P2_STATE2_REG_2__SCAN_IN), .Y(n10054));
  NAND3X1 g06826(.A(n9208), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .Y(n10055));
  NOR4X1  g06827(.A(n9811), .B(n9996), .C(n9772), .D(n9827), .Y(n10056));
  NOR3X1  g06828(.A(n9997), .B(n10056), .C(n9759), .Y(n10058));
  NOR2X1  g06829(.A(n10058), .B(n9757), .Y(n10059));
  OAI21X1 g06830(.A0(n10059), .A1(n10055), .B0(n10054), .Y(n10060));
  NAND3X1 g06831(.A(n10060), .B(n9744), .C(n9740), .Y(n10061));
  NOR4X1  g06832(.A(n10056), .B(n9759), .C(n9836), .D(n9997), .Y(n10062));
  OAI21X1 g06833(.A0(n10062), .A1(n9757), .B0(n10055), .Y(n10063));
  INVX1   g06834(.A(n10051), .Y(n10064));
  NOR3X1  g06835(.A(n10053), .B(n10051), .C(n9700), .Y(n10065));
  AOI21X1 g06836(.A0(n10064), .A1(P2_STATE2_REG_3__SCAN_IN), .B0(n10065), .Y(n10066));
  NAND3X1 g06837(.A(n10066), .B(n10063), .C(n9740), .Y(n10067));
  NAND2X1 g06838(.A(n10067), .B(P2_INSTQUEUE_REG_13__7__SCAN_IN), .Y(n10068));
  INVX1   g06839(.A(n9997), .Y(n10069));
  OAI22X1 g06840(.A0(n10064), .A1(n9854), .B0(n9853), .B1(n10069), .Y(n10070));
  AOI21X1 g06841(.A0(n10056), .A1(n9847), .B0(n10070), .Y(n10071));
  NAND3X1 g06842(.A(n10071), .B(n10068), .C(n10061), .Y(P2_U3159));
  NAND3X1 g06843(.A(n10060), .B(n9861), .C(n9740), .Y(n10073));
  NAND2X1 g06844(.A(n10067), .B(P2_INSTQUEUE_REG_13__6__SCAN_IN), .Y(n10074));
  OAI22X1 g06845(.A0(n10064), .A1(n9873), .B0(n9872), .B1(n10069), .Y(n10075));
  AOI21X1 g06846(.A0(n10056), .A1(n9867), .B0(n10075), .Y(n10076));
  NAND3X1 g06847(.A(n10076), .B(n10074), .C(n10073), .Y(P2_U3158));
  NAND3X1 g06848(.A(n10060), .B(n9880), .C(n9740), .Y(n10078));
  NAND2X1 g06849(.A(n10067), .B(P2_INSTQUEUE_REG_13__5__SCAN_IN), .Y(n10079));
  OAI22X1 g06850(.A0(n10064), .A1(n9892), .B0(n9891), .B1(n10069), .Y(n10080));
  AOI21X1 g06851(.A0(n10056), .A1(n9886), .B0(n10080), .Y(n10081));
  NAND3X1 g06852(.A(n10081), .B(n10079), .C(n10078), .Y(P2_U3157));
  NAND3X1 g06853(.A(n10060), .B(n9899), .C(n9740), .Y(n10083));
  NAND2X1 g06854(.A(n10067), .B(P2_INSTQUEUE_REG_13__4__SCAN_IN), .Y(n10084));
  OAI22X1 g06855(.A0(n10064), .A1(n9911), .B0(n9910), .B1(n10069), .Y(n10085));
  AOI21X1 g06856(.A0(n10056), .A1(n9905), .B0(n10085), .Y(n10086));
  NAND3X1 g06857(.A(n10086), .B(n10084), .C(n10083), .Y(P2_U3156));
  NAND3X1 g06858(.A(n10060), .B(n9918), .C(n9740), .Y(n10088));
  NAND2X1 g06859(.A(n10067), .B(P2_INSTQUEUE_REG_13__3__SCAN_IN), .Y(n10089));
  OAI22X1 g06860(.A0(n10064), .A1(n9930), .B0(n9929), .B1(n10069), .Y(n10090));
  AOI21X1 g06861(.A0(n10056), .A1(n9924), .B0(n10090), .Y(n10091));
  NAND3X1 g06862(.A(n10091), .B(n10089), .C(n10088), .Y(P2_U3155));
  NAND3X1 g06863(.A(n10060), .B(n9937), .C(n9740), .Y(n10093));
  NAND2X1 g06864(.A(n10067), .B(P2_INSTQUEUE_REG_13__2__SCAN_IN), .Y(n10094));
  OAI22X1 g06865(.A0(n10064), .A1(n9949), .B0(n9948), .B1(n10069), .Y(n10095));
  AOI21X1 g06866(.A0(n10056), .A1(n9943), .B0(n10095), .Y(n10096));
  NAND3X1 g06867(.A(n10096), .B(n10094), .C(n10093), .Y(P2_U3154));
  NAND3X1 g06868(.A(n10060), .B(n9956), .C(n9740), .Y(n10098));
  NAND2X1 g06869(.A(n10067), .B(P2_INSTQUEUE_REG_13__1__SCAN_IN), .Y(n10099));
  OAI22X1 g06870(.A0(n10064), .A1(n9968), .B0(n9967), .B1(n10069), .Y(n10100));
  AOI21X1 g06871(.A0(n10056), .A1(n9962), .B0(n10100), .Y(n10101));
  NAND3X1 g06872(.A(n10101), .B(n10099), .C(n10098), .Y(P2_U3153));
  NAND3X1 g06873(.A(n10060), .B(n9975), .C(n9740), .Y(n10103));
  NAND2X1 g06874(.A(n10067), .B(P2_INSTQUEUE_REG_13__0__SCAN_IN), .Y(n10104));
  OAI22X1 g06875(.A0(n10064), .A1(n9987), .B0(n9986), .B1(n10069), .Y(n10105));
  AOI21X1 g06876(.A0(n10056), .A1(n9981), .B0(n10105), .Y(n10106));
  NAND3X1 g06877(.A(n10106), .B(n10104), .C(n10103), .Y(P2_U3152));
  NOR4X1  g06878(.A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n9223), .C(n9221), .D(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Y(n10108));
  NAND2X1 g06879(.A(n9614), .B(n9595), .Y(n10109));
  NOR3X1  g06880(.A(n10109), .B(n9663), .C(n9633), .Y(n10110));
  OAI21X1 g06881(.A0(n10110), .A1(n10108), .B0(P2_STATE2_REG_2__SCAN_IN), .Y(n10111));
  NOR3X1  g06882(.A(n9780), .B(n9819), .C(n9786), .Y(n10112));
  NOR4X1  g06883(.A(n9810), .B(n9784), .C(n9771), .D(n9827), .Y(n10113));
  NOR3X1  g06884(.A(n10056), .B(n10113), .C(n9759), .Y(n10115));
  OAI21X1 g06885(.A0(n10115), .A1(n9757), .B0(n10112), .Y(n10116));
  NAND2X1 g06886(.A(n10116), .B(n10111), .Y(n10117));
  NAND3X1 g06887(.A(n10117), .B(n9744), .C(n9740), .Y(n10118));
  NOR4X1  g06888(.A(n10113), .B(n9759), .C(n9836), .D(n10056), .Y(n10119));
  OAI22X1 g06889(.A0(n9757), .A1(n10119), .B0(n9780), .B1(n10004), .Y(n10120));
  INVX1   g06890(.A(n10108), .Y(n10121));
  NOR3X1  g06891(.A(n10110), .B(n10108), .C(n9700), .Y(n10122));
  AOI21X1 g06892(.A0(n10121), .A1(P2_STATE2_REG_3__SCAN_IN), .B0(n10122), .Y(n10123));
  NAND3X1 g06893(.A(n10123), .B(n10120), .C(n9740), .Y(n10124));
  NAND2X1 g06894(.A(n10124), .B(P2_INSTQUEUE_REG_12__7__SCAN_IN), .Y(n10125));
  INVX1   g06895(.A(n10056), .Y(n10126));
  OAI22X1 g06896(.A0(n10121), .A1(n9854), .B0(n9853), .B1(n10126), .Y(n10127));
  AOI21X1 g06897(.A0(n10113), .A1(n9847), .B0(n10127), .Y(n10128));
  NAND3X1 g06898(.A(n10128), .B(n10125), .C(n10118), .Y(P2_U3151));
  NAND3X1 g06899(.A(n10117), .B(n9861), .C(n9740), .Y(n10130));
  NAND2X1 g06900(.A(n10124), .B(P2_INSTQUEUE_REG_12__6__SCAN_IN), .Y(n10131));
  OAI22X1 g06901(.A0(n10121), .A1(n9873), .B0(n9872), .B1(n10126), .Y(n10132));
  AOI21X1 g06902(.A0(n10113), .A1(n9867), .B0(n10132), .Y(n10133));
  NAND3X1 g06903(.A(n10133), .B(n10131), .C(n10130), .Y(P2_U3150));
  NAND3X1 g06904(.A(n10117), .B(n9880), .C(n9740), .Y(n10135));
  NAND2X1 g06905(.A(n10124), .B(P2_INSTQUEUE_REG_12__5__SCAN_IN), .Y(n10136));
  OAI22X1 g06906(.A0(n10121), .A1(n9892), .B0(n9891), .B1(n10126), .Y(n10137));
  AOI21X1 g06907(.A0(n10113), .A1(n9886), .B0(n10137), .Y(n10138));
  NAND3X1 g06908(.A(n10138), .B(n10136), .C(n10135), .Y(P2_U3149));
  NAND3X1 g06909(.A(n10117), .B(n9899), .C(n9740), .Y(n10140));
  NAND2X1 g06910(.A(n10124), .B(P2_INSTQUEUE_REG_12__4__SCAN_IN), .Y(n10141));
  OAI22X1 g06911(.A0(n10121), .A1(n9911), .B0(n9910), .B1(n10126), .Y(n10142));
  AOI21X1 g06912(.A0(n10113), .A1(n9905), .B0(n10142), .Y(n10143));
  NAND3X1 g06913(.A(n10143), .B(n10141), .C(n10140), .Y(P2_U3148));
  NAND3X1 g06914(.A(n10117), .B(n9918), .C(n9740), .Y(n10145));
  NAND2X1 g06915(.A(n10124), .B(P2_INSTQUEUE_REG_12__3__SCAN_IN), .Y(n10146));
  OAI22X1 g06916(.A0(n10121), .A1(n9930), .B0(n9929), .B1(n10126), .Y(n10147));
  AOI21X1 g06917(.A0(n10113), .A1(n9924), .B0(n10147), .Y(n10148));
  NAND3X1 g06918(.A(n10148), .B(n10146), .C(n10145), .Y(P2_U3147));
  NAND3X1 g06919(.A(n10117), .B(n9937), .C(n9740), .Y(n10150));
  NAND2X1 g06920(.A(n10124), .B(P2_INSTQUEUE_REG_12__2__SCAN_IN), .Y(n10151));
  OAI22X1 g06921(.A0(n10121), .A1(n9949), .B0(n9948), .B1(n10126), .Y(n10152));
  AOI21X1 g06922(.A0(n10113), .A1(n9943), .B0(n10152), .Y(n10153));
  NAND3X1 g06923(.A(n10153), .B(n10151), .C(n10150), .Y(P2_U3146));
  NAND3X1 g06924(.A(n10117), .B(n9956), .C(n9740), .Y(n10155));
  NAND2X1 g06925(.A(n10124), .B(P2_INSTQUEUE_REG_12__1__SCAN_IN), .Y(n10156));
  OAI22X1 g06926(.A0(n10121), .A1(n9968), .B0(n9967), .B1(n10126), .Y(n10157));
  AOI21X1 g06927(.A0(n10113), .A1(n9962), .B0(n10157), .Y(n10158));
  NAND3X1 g06928(.A(n10158), .B(n10156), .C(n10155), .Y(P2_U3145));
  NAND3X1 g06929(.A(n10117), .B(n9975), .C(n9740), .Y(n10160));
  NAND2X1 g06930(.A(n10124), .B(P2_INSTQUEUE_REG_12__0__SCAN_IN), .Y(n10161));
  OAI22X1 g06931(.A0(n10121), .A1(n9987), .B0(n9986), .B1(n10126), .Y(n10162));
  AOI21X1 g06932(.A0(n10113), .A1(n9981), .B0(n10162), .Y(n10163));
  NAND3X1 g06933(.A(n10163), .B(n10161), .C(n10160), .Y(P2_U3144));
  NOR3X1  g06934(.A(n9745), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C(n9221), .Y(n10165));
  NOR2X1  g06935(.A(n9614), .B(n9595), .Y(n10166));
  NAND3X1 g06936(.A(n10166), .B(n9815), .C(n9633), .Y(n10167));
  INVX1   g06937(.A(n10167), .Y(n10168));
  OAI21X1 g06938(.A0(n10168), .A1(n10165), .B0(P2_STATE2_REG_2__SCAN_IN), .Y(n10169));
  NAND3X1 g06939(.A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n9223), .C(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .Y(n10170));
  NOR4X1  g06940(.A(n9810), .B(n9784), .C(n9772), .D(n9827), .Y(n10171));
  NOR3X1  g06941(.A(n10113), .B(n10171), .C(n9759), .Y(n10173));
  NOR2X1  g06942(.A(n10173), .B(n9757), .Y(n10174));
  OAI21X1 g06943(.A0(n10174), .A1(n10170), .B0(n10169), .Y(n10175));
  NAND3X1 g06944(.A(n10175), .B(n9744), .C(n9740), .Y(n10176));
  NOR4X1  g06945(.A(n10171), .B(n9759), .C(n9836), .D(n10113), .Y(n10177));
  OAI21X1 g06946(.A0(n10177), .A1(n9757), .B0(n10170), .Y(n10178));
  INVX1   g06947(.A(n10165), .Y(n10179));
  NOR3X1  g06948(.A(n10168), .B(n10165), .C(n9700), .Y(n10180));
  AOI21X1 g06949(.A0(n10179), .A1(P2_STATE2_REG_3__SCAN_IN), .B0(n10180), .Y(n10181));
  NAND3X1 g06950(.A(n10181), .B(n10178), .C(n9740), .Y(n10182));
  NAND2X1 g06951(.A(n10182), .B(P2_INSTQUEUE_REG_11__7__SCAN_IN), .Y(n10183));
  INVX1   g06952(.A(n10113), .Y(n10184));
  OAI22X1 g06953(.A0(n10179), .A1(n9854), .B0(n9853), .B1(n10184), .Y(n10185));
  AOI21X1 g06954(.A0(n10171), .A1(n9847), .B0(n10185), .Y(n10186));
  NAND3X1 g06955(.A(n10186), .B(n10183), .C(n10176), .Y(P2_U3143));
  NAND3X1 g06956(.A(n10175), .B(n9861), .C(n9740), .Y(n10188));
  NAND2X1 g06957(.A(n10182), .B(P2_INSTQUEUE_REG_11__6__SCAN_IN), .Y(n10189));
  OAI22X1 g06958(.A0(n10179), .A1(n9873), .B0(n9872), .B1(n10184), .Y(n10190));
  AOI21X1 g06959(.A0(n10171), .A1(n9867), .B0(n10190), .Y(n10191));
  NAND3X1 g06960(.A(n10191), .B(n10189), .C(n10188), .Y(P2_U3142));
  NAND3X1 g06961(.A(n10175), .B(n9880), .C(n9740), .Y(n10193));
  NAND2X1 g06962(.A(n10182), .B(P2_INSTQUEUE_REG_11__5__SCAN_IN), .Y(n10194));
  OAI22X1 g06963(.A0(n10179), .A1(n9892), .B0(n9891), .B1(n10184), .Y(n10195));
  AOI21X1 g06964(.A0(n10171), .A1(n9886), .B0(n10195), .Y(n10196));
  NAND3X1 g06965(.A(n10196), .B(n10194), .C(n10193), .Y(P2_U3141));
  NAND3X1 g06966(.A(n10175), .B(n9899), .C(n9740), .Y(n10198));
  NAND2X1 g06967(.A(n10182), .B(P2_INSTQUEUE_REG_11__4__SCAN_IN), .Y(n10199));
  OAI22X1 g06968(.A0(n10179), .A1(n9911), .B0(n9910), .B1(n10184), .Y(n10200));
  AOI21X1 g06969(.A0(n10171), .A1(n9905), .B0(n10200), .Y(n10201));
  NAND3X1 g06970(.A(n10201), .B(n10199), .C(n10198), .Y(P2_U3140));
  NAND3X1 g06971(.A(n10175), .B(n9918), .C(n9740), .Y(n10203));
  NAND2X1 g06972(.A(n10182), .B(P2_INSTQUEUE_REG_11__3__SCAN_IN), .Y(n10204));
  OAI22X1 g06973(.A0(n10179), .A1(n9930), .B0(n9929), .B1(n10184), .Y(n10205));
  AOI21X1 g06974(.A0(n10171), .A1(n9924), .B0(n10205), .Y(n10206));
  NAND3X1 g06975(.A(n10206), .B(n10204), .C(n10203), .Y(P2_U3139));
  NAND3X1 g06976(.A(n10175), .B(n9937), .C(n9740), .Y(n10208));
  NAND2X1 g06977(.A(n10182), .B(P2_INSTQUEUE_REG_11__2__SCAN_IN), .Y(n10209));
  OAI22X1 g06978(.A0(n10179), .A1(n9949), .B0(n9948), .B1(n10184), .Y(n10210));
  AOI21X1 g06979(.A0(n10171), .A1(n9943), .B0(n10210), .Y(n10211));
  NAND3X1 g06980(.A(n10211), .B(n10209), .C(n10208), .Y(P2_U3138));
  NAND3X1 g06981(.A(n10175), .B(n9956), .C(n9740), .Y(n10213));
  NAND2X1 g06982(.A(n10182), .B(P2_INSTQUEUE_REG_11__1__SCAN_IN), .Y(n10214));
  OAI22X1 g06983(.A0(n10179), .A1(n9968), .B0(n9967), .B1(n10184), .Y(n10215));
  AOI21X1 g06984(.A0(n10171), .A1(n9962), .B0(n10215), .Y(n10216));
  NAND3X1 g06985(.A(n10216), .B(n10214), .C(n10213), .Y(P2_U3137));
  NAND3X1 g06986(.A(n10175), .B(n9975), .C(n9740), .Y(n10218));
  NAND2X1 g06987(.A(n10182), .B(P2_INSTQUEUE_REG_11__0__SCAN_IN), .Y(n10219));
  OAI22X1 g06988(.A0(n10179), .A1(n9987), .B0(n9986), .B1(n10184), .Y(n10220));
  AOI21X1 g06989(.A0(n10171), .A1(n9981), .B0(n10220), .Y(n10221));
  NAND3X1 g06990(.A(n10221), .B(n10219), .C(n10218), .Y(P2_U3136));
  NOR4X1  g06991(.A(n9208), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C(n9221), .D(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Y(n10223));
  NOR2X1  g06992(.A(n9752), .B(n9595), .Y(n10224));
  NAND3X1 g06993(.A(n10224), .B(n9815), .C(n9633), .Y(n10225));
  INVX1   g06994(.A(n10225), .Y(n10226));
  OAI21X1 g06995(.A0(n10226), .A1(n10223), .B0(P2_STATE2_REG_2__SCAN_IN), .Y(n10227));
  NOR3X1  g06996(.A(n9779), .B(n9819), .C(n9787), .Y(n10228));
  NOR4X1  g06997(.A(n9810), .B(n9996), .C(n9771), .D(n9827), .Y(n10229));
  NOR3X1  g06998(.A(n10171), .B(n10229), .C(n9759), .Y(n10231));
  OAI21X1 g06999(.A0(n10231), .A1(n9757), .B0(n10228), .Y(n10232));
  NAND2X1 g07000(.A(n10232), .B(n10227), .Y(n10233));
  NAND3X1 g07001(.A(n10233), .B(n9744), .C(n9740), .Y(n10234));
  NOR2X1  g07002(.A(n9819), .B(n9787), .Y(n10235));
  INVX1   g07003(.A(n10235), .Y(n10236));
  NOR4X1  g07004(.A(n10229), .B(n9759), .C(n9836), .D(n10171), .Y(n10237));
  OAI22X1 g07005(.A0(n10236), .A1(n9779), .B0(n9757), .B1(n10237), .Y(n10238));
  INVX1   g07006(.A(n10223), .Y(n10239));
  NOR3X1  g07007(.A(n10226), .B(n10223), .C(n9700), .Y(n10240));
  AOI21X1 g07008(.A0(n10239), .A1(P2_STATE2_REG_3__SCAN_IN), .B0(n10240), .Y(n10241));
  NAND3X1 g07009(.A(n10241), .B(n10238), .C(n9740), .Y(n10242));
  NAND2X1 g07010(.A(n10242), .B(P2_INSTQUEUE_REG_10__7__SCAN_IN), .Y(n10243));
  INVX1   g07011(.A(n10171), .Y(n10244));
  OAI22X1 g07012(.A0(n10239), .A1(n9854), .B0(n9853), .B1(n10244), .Y(n10245));
  AOI21X1 g07013(.A0(n10229), .A1(n9847), .B0(n10245), .Y(n10246));
  NAND3X1 g07014(.A(n10246), .B(n10243), .C(n10234), .Y(P2_U3135));
  NAND3X1 g07015(.A(n10233), .B(n9861), .C(n9740), .Y(n10248));
  NAND2X1 g07016(.A(n10242), .B(P2_INSTQUEUE_REG_10__6__SCAN_IN), .Y(n10249));
  OAI22X1 g07017(.A0(n10239), .A1(n9873), .B0(n9872), .B1(n10244), .Y(n10250));
  AOI21X1 g07018(.A0(n10229), .A1(n9867), .B0(n10250), .Y(n10251));
  NAND3X1 g07019(.A(n10251), .B(n10249), .C(n10248), .Y(P2_U3134));
  NAND3X1 g07020(.A(n10233), .B(n9880), .C(n9740), .Y(n10253));
  NAND2X1 g07021(.A(n10242), .B(P2_INSTQUEUE_REG_10__5__SCAN_IN), .Y(n10254));
  OAI22X1 g07022(.A0(n10239), .A1(n9892), .B0(n9891), .B1(n10244), .Y(n10255));
  AOI21X1 g07023(.A0(n10229), .A1(n9886), .B0(n10255), .Y(n10256));
  NAND3X1 g07024(.A(n10256), .B(n10254), .C(n10253), .Y(P2_U3133));
  NAND3X1 g07025(.A(n10233), .B(n9899), .C(n9740), .Y(n10258));
  NAND2X1 g07026(.A(n10242), .B(P2_INSTQUEUE_REG_10__4__SCAN_IN), .Y(n10259));
  OAI22X1 g07027(.A0(n10239), .A1(n9911), .B0(n9910), .B1(n10244), .Y(n10260));
  AOI21X1 g07028(.A0(n10229), .A1(n9905), .B0(n10260), .Y(n10261));
  NAND3X1 g07029(.A(n10261), .B(n10259), .C(n10258), .Y(P2_U3132));
  NAND3X1 g07030(.A(n10233), .B(n9918), .C(n9740), .Y(n10263));
  NAND2X1 g07031(.A(n10242), .B(P2_INSTQUEUE_REG_10__3__SCAN_IN), .Y(n10264));
  OAI22X1 g07032(.A0(n10239), .A1(n9930), .B0(n9929), .B1(n10244), .Y(n10265));
  AOI21X1 g07033(.A0(n10229), .A1(n9924), .B0(n10265), .Y(n10266));
  NAND3X1 g07034(.A(n10266), .B(n10264), .C(n10263), .Y(P2_U3131));
  NAND3X1 g07035(.A(n10233), .B(n9937), .C(n9740), .Y(n10268));
  NAND2X1 g07036(.A(n10242), .B(P2_INSTQUEUE_REG_10__2__SCAN_IN), .Y(n10269));
  OAI22X1 g07037(.A0(n10239), .A1(n9949), .B0(n9948), .B1(n10244), .Y(n10270));
  AOI21X1 g07038(.A0(n10229), .A1(n9943), .B0(n10270), .Y(n10271));
  NAND3X1 g07039(.A(n10271), .B(n10269), .C(n10268), .Y(P2_U3130));
  NAND3X1 g07040(.A(n10233), .B(n9956), .C(n9740), .Y(n10273));
  NAND2X1 g07041(.A(n10242), .B(P2_INSTQUEUE_REG_10__1__SCAN_IN), .Y(n10274));
  OAI22X1 g07042(.A0(n10239), .A1(n9968), .B0(n9967), .B1(n10244), .Y(n10275));
  AOI21X1 g07043(.A0(n10229), .A1(n9962), .B0(n10275), .Y(n10276));
  NAND3X1 g07044(.A(n10276), .B(n10274), .C(n10273), .Y(P2_U3129));
  NAND3X1 g07045(.A(n10233), .B(n9975), .C(n9740), .Y(n10278));
  NAND2X1 g07046(.A(n10242), .B(P2_INSTQUEUE_REG_10__0__SCAN_IN), .Y(n10279));
  OAI22X1 g07047(.A0(n10239), .A1(n9987), .B0(n9986), .B1(n10244), .Y(n10280));
  AOI21X1 g07048(.A0(n10229), .A1(n9981), .B0(n10280), .Y(n10281));
  NAND3X1 g07049(.A(n10281), .B(n10279), .C(n10278), .Y(P2_U3128));
  NOR4X1  g07050(.A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C(n9221), .D(n9209), .Y(n10283));
  NOR2X1  g07051(.A(n9614), .B(n9751), .Y(n10284));
  NAND3X1 g07052(.A(n10284), .B(n9815), .C(n9633), .Y(n10285));
  INVX1   g07053(.A(n10285), .Y(n10286));
  OAI21X1 g07054(.A0(n10286), .A1(n10283), .B0(P2_STATE2_REG_2__SCAN_IN), .Y(n10287));
  NAND3X1 g07055(.A(n9208), .B(n9223), .C(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .Y(n10288));
  NOR4X1  g07056(.A(n9810), .B(n9996), .C(n9772), .D(n9827), .Y(n10289));
  NOR3X1  g07057(.A(n10229), .B(n10289), .C(n9759), .Y(n10291));
  NOR2X1  g07058(.A(n10291), .B(n9757), .Y(n10292));
  OAI21X1 g07059(.A0(n10292), .A1(n10288), .B0(n10287), .Y(n10293));
  NAND3X1 g07060(.A(n10293), .B(n9744), .C(n9740), .Y(n10294));
  NOR4X1  g07061(.A(n10289), .B(n9759), .C(n9836), .D(n10229), .Y(n10295));
  OAI21X1 g07062(.A0(n10295), .A1(n9757), .B0(n10288), .Y(n10296));
  INVX1   g07063(.A(n10283), .Y(n10297));
  NOR3X1  g07064(.A(n10286), .B(n10283), .C(n9700), .Y(n10298));
  AOI21X1 g07065(.A0(n10297), .A1(P2_STATE2_REG_3__SCAN_IN), .B0(n10298), .Y(n10299));
  NAND3X1 g07066(.A(n10299), .B(n10296), .C(n9740), .Y(n10300));
  NAND2X1 g07067(.A(n10300), .B(P2_INSTQUEUE_REG_9__7__SCAN_IN), .Y(n10301));
  INVX1   g07068(.A(n10229), .Y(n10302));
  OAI22X1 g07069(.A0(n10297), .A1(n9854), .B0(n9853), .B1(n10302), .Y(n10303));
  AOI21X1 g07070(.A0(n10289), .A1(n9847), .B0(n10303), .Y(n10304));
  NAND3X1 g07071(.A(n10304), .B(n10301), .C(n10294), .Y(P2_U3127));
  NAND3X1 g07072(.A(n10293), .B(n9861), .C(n9740), .Y(n10306));
  NAND2X1 g07073(.A(n10300), .B(P2_INSTQUEUE_REG_9__6__SCAN_IN), .Y(n10307));
  OAI22X1 g07074(.A0(n10297), .A1(n9873), .B0(n9872), .B1(n10302), .Y(n10308));
  AOI21X1 g07075(.A0(n10289), .A1(n9867), .B0(n10308), .Y(n10309));
  NAND3X1 g07076(.A(n10309), .B(n10307), .C(n10306), .Y(P2_U3126));
  NAND3X1 g07077(.A(n10293), .B(n9880), .C(n9740), .Y(n10311));
  NAND2X1 g07078(.A(n10300), .B(P2_INSTQUEUE_REG_9__5__SCAN_IN), .Y(n10312));
  OAI22X1 g07079(.A0(n10297), .A1(n9892), .B0(n9891), .B1(n10302), .Y(n10313));
  AOI21X1 g07080(.A0(n10289), .A1(n9886), .B0(n10313), .Y(n10314));
  NAND3X1 g07081(.A(n10314), .B(n10312), .C(n10311), .Y(P2_U3125));
  NAND3X1 g07082(.A(n10293), .B(n9899), .C(n9740), .Y(n10316));
  NAND2X1 g07083(.A(n10300), .B(P2_INSTQUEUE_REG_9__4__SCAN_IN), .Y(n10317));
  OAI22X1 g07084(.A0(n10297), .A1(n9911), .B0(n9910), .B1(n10302), .Y(n10318));
  AOI21X1 g07085(.A0(n10289), .A1(n9905), .B0(n10318), .Y(n10319));
  NAND3X1 g07086(.A(n10319), .B(n10317), .C(n10316), .Y(P2_U3124));
  NAND3X1 g07087(.A(n10293), .B(n9918), .C(n9740), .Y(n10321));
  NAND2X1 g07088(.A(n10300), .B(P2_INSTQUEUE_REG_9__3__SCAN_IN), .Y(n10322));
  OAI22X1 g07089(.A0(n10297), .A1(n9930), .B0(n9929), .B1(n10302), .Y(n10323));
  AOI21X1 g07090(.A0(n10289), .A1(n9924), .B0(n10323), .Y(n10324));
  NAND3X1 g07091(.A(n10324), .B(n10322), .C(n10321), .Y(P2_U3123));
  NAND3X1 g07092(.A(n10293), .B(n9937), .C(n9740), .Y(n10326));
  NAND2X1 g07093(.A(n10300), .B(P2_INSTQUEUE_REG_9__2__SCAN_IN), .Y(n10327));
  OAI22X1 g07094(.A0(n10297), .A1(n9949), .B0(n9948), .B1(n10302), .Y(n10328));
  AOI21X1 g07095(.A0(n10289), .A1(n9943), .B0(n10328), .Y(n10329));
  NAND3X1 g07096(.A(n10329), .B(n10327), .C(n10326), .Y(P2_U3122));
  NAND3X1 g07097(.A(n10293), .B(n9956), .C(n9740), .Y(n10331));
  NAND2X1 g07098(.A(n10300), .B(P2_INSTQUEUE_REG_9__1__SCAN_IN), .Y(n10332));
  OAI22X1 g07099(.A0(n10297), .A1(n9968), .B0(n9967), .B1(n10302), .Y(n10333));
  AOI21X1 g07100(.A0(n10289), .A1(n9962), .B0(n10333), .Y(n10334));
  NAND3X1 g07101(.A(n10334), .B(n10332), .C(n10331), .Y(P2_U3121));
  NAND3X1 g07102(.A(n10293), .B(n9975), .C(n9740), .Y(n10336));
  NAND2X1 g07103(.A(n10300), .B(P2_INSTQUEUE_REG_9__0__SCAN_IN), .Y(n10337));
  OAI22X1 g07104(.A0(n10297), .A1(n9987), .B0(n9986), .B1(n10302), .Y(n10338));
  AOI21X1 g07105(.A0(n10289), .A1(n9981), .B0(n10338), .Y(n10339));
  NAND3X1 g07106(.A(n10339), .B(n10337), .C(n10336), .Y(P2_U3120));
  NOR4X1  g07107(.A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C(n9221), .D(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Y(n10341));
  NOR2X1  g07108(.A(n9752), .B(n9751), .Y(n10342));
  NAND3X1 g07109(.A(n10342), .B(n9815), .C(n9633), .Y(n10343));
  INVX1   g07110(.A(n10343), .Y(n10344));
  OAI21X1 g07111(.A0(n10344), .A1(n10341), .B0(P2_STATE2_REG_2__SCAN_IN), .Y(n10345));
  NOR3X1  g07112(.A(n9780), .B(n9819), .C(n9787), .Y(n10346));
  OAI21X1 g07113(.A0(n9760), .A1(n9791), .B0(n9796), .Y(n10347));
  AOI21X1 g07114(.A0(n9808), .A1(n10347), .B0(n9797), .Y(n10349));
  XOR2X1  g07115(.A(n9826), .B(n10349), .Y(n10350));
  NOR3X1  g07116(.A(n10289), .B(n10406), .C(n9759), .Y(n10353));
  OAI21X1 g07117(.A0(n10353), .A1(n9757), .B0(n10346), .Y(n10354));
  NAND2X1 g07118(.A(n10354), .B(n10345), .Y(n10355));
  NAND3X1 g07119(.A(n10355), .B(n9744), .C(n9740), .Y(n10356));
  NOR4X1  g07120(.A(n10406), .B(n9759), .C(n9836), .D(n10289), .Y(n10357));
  OAI22X1 g07121(.A0(n10236), .A1(n9780), .B0(n9757), .B1(n10357), .Y(n10358));
  INVX1   g07122(.A(n10341), .Y(n10359));
  NOR3X1  g07123(.A(n10344), .B(n10341), .C(n9700), .Y(n10360));
  AOI21X1 g07124(.A0(n10359), .A1(P2_STATE2_REG_3__SCAN_IN), .B0(n10360), .Y(n10361));
  NAND3X1 g07125(.A(n10361), .B(n10358), .C(n9740), .Y(n10362));
  NAND2X1 g07126(.A(n10362), .B(P2_INSTQUEUE_REG_8__7__SCAN_IN), .Y(n10363));
  INVX1   g07127(.A(n10289), .Y(n10364));
  OAI22X1 g07128(.A0(n10359), .A1(n9854), .B0(n9853), .B1(n10364), .Y(n10365));
  AOI21X1 g07129(.A0(n10406), .A1(n9847), .B0(n10365), .Y(n10366));
  NAND3X1 g07130(.A(n10366), .B(n10363), .C(n10356), .Y(P2_U3119));
  NAND3X1 g07131(.A(n10355), .B(n9861), .C(n9740), .Y(n10368));
  NAND2X1 g07132(.A(n10362), .B(P2_INSTQUEUE_REG_8__6__SCAN_IN), .Y(n10369));
  OAI22X1 g07133(.A0(n10359), .A1(n9873), .B0(n9872), .B1(n10364), .Y(n10370));
  AOI21X1 g07134(.A0(n10406), .A1(n9867), .B0(n10370), .Y(n10371));
  NAND3X1 g07135(.A(n10371), .B(n10369), .C(n10368), .Y(P2_U3118));
  NAND3X1 g07136(.A(n10355), .B(n9880), .C(n9740), .Y(n10373));
  NAND2X1 g07137(.A(n10362), .B(P2_INSTQUEUE_REG_8__5__SCAN_IN), .Y(n10374));
  OAI22X1 g07138(.A0(n10359), .A1(n9892), .B0(n9891), .B1(n10364), .Y(n10375));
  AOI21X1 g07139(.A0(n10406), .A1(n9886), .B0(n10375), .Y(n10376));
  NAND3X1 g07140(.A(n10376), .B(n10374), .C(n10373), .Y(P2_U3117));
  NAND3X1 g07141(.A(n10355), .B(n9899), .C(n9740), .Y(n10378));
  NAND2X1 g07142(.A(n10362), .B(P2_INSTQUEUE_REG_8__4__SCAN_IN), .Y(n10379));
  OAI22X1 g07143(.A0(n10359), .A1(n9911), .B0(n9910), .B1(n10364), .Y(n10380));
  AOI21X1 g07144(.A0(n10406), .A1(n9905), .B0(n10380), .Y(n10381));
  NAND3X1 g07145(.A(n10381), .B(n10379), .C(n10378), .Y(P2_U3116));
  NAND3X1 g07146(.A(n10355), .B(n9918), .C(n9740), .Y(n10383));
  NAND2X1 g07147(.A(n10362), .B(P2_INSTQUEUE_REG_8__3__SCAN_IN), .Y(n10384));
  OAI22X1 g07148(.A0(n10359), .A1(n9930), .B0(n9929), .B1(n10364), .Y(n10385));
  AOI21X1 g07149(.A0(n10406), .A1(n9924), .B0(n10385), .Y(n10386));
  NAND3X1 g07150(.A(n10386), .B(n10384), .C(n10383), .Y(P2_U3115));
  NAND3X1 g07151(.A(n10355), .B(n9937), .C(n9740), .Y(n10388));
  NAND2X1 g07152(.A(n10362), .B(P2_INSTQUEUE_REG_8__2__SCAN_IN), .Y(n10389));
  OAI22X1 g07153(.A0(n10359), .A1(n9949), .B0(n9948), .B1(n10364), .Y(n10390));
  AOI21X1 g07154(.A0(n10406), .A1(n9943), .B0(n10390), .Y(n10391));
  NAND3X1 g07155(.A(n10391), .B(n10389), .C(n10388), .Y(P2_U3114));
  NAND3X1 g07156(.A(n10355), .B(n9956), .C(n9740), .Y(n10393));
  NAND2X1 g07157(.A(n10362), .B(P2_INSTQUEUE_REG_8__1__SCAN_IN), .Y(n10394));
  OAI22X1 g07158(.A0(n10359), .A1(n9968), .B0(n9967), .B1(n10364), .Y(n10395));
  AOI21X1 g07159(.A0(n10406), .A1(n9962), .B0(n10395), .Y(n10396));
  NAND3X1 g07160(.A(n10396), .B(n10394), .C(n10393), .Y(P2_U3113));
  NAND3X1 g07161(.A(n10355), .B(n9975), .C(n9740), .Y(n10398));
  NAND2X1 g07162(.A(n10362), .B(P2_INSTQUEUE_REG_8__0__SCAN_IN), .Y(n10399));
  OAI22X1 g07163(.A0(n10359), .A1(n9987), .B0(n9986), .B1(n10364), .Y(n10400));
  AOI21X1 g07164(.A0(n10406), .A1(n9981), .B0(n10400), .Y(n10401));
  NAND3X1 g07165(.A(n10401), .B(n10399), .C(n10398), .Y(P2_U3112));
  NOR3X1  g07166(.A(n9753), .B(n9815), .C(n9633), .Y(n10403));
  OAI21X1 g07167(.A0(n10403), .A1(n9817), .B0(P2_STATE2_REG_2__SCAN_IN), .Y(n10404));
  NAND3X1 g07168(.A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C(n9221), .Y(n10405));
  NOR4X1  g07169(.A(n9809), .B(n9801), .C(n9830), .D(n10350), .Y(n10406));
  NOR4X1  g07170(.A(n9811), .B(n9784), .C(n9772), .D(n10350), .Y(n10407));
  NOR3X1  g07171(.A(n10407), .B(n10406), .C(n9759), .Y(n10408));
  NOR2X1  g07172(.A(n10408), .B(n9757), .Y(n10409));
  OAI21X1 g07173(.A0(n10409), .A1(n10405), .B0(n10404), .Y(n10410));
  NAND3X1 g07174(.A(n10410), .B(n9744), .C(n9740), .Y(n10411));
  NOR4X1  g07175(.A(n10406), .B(n9759), .C(n9836), .D(n10407), .Y(n10412));
  OAI21X1 g07176(.A0(n10412), .A1(n9757), .B0(n10405), .Y(n10413));
  INVX1   g07177(.A(n9817), .Y(n10414));
  NOR3X1  g07178(.A(n10403), .B(n9817), .C(n9700), .Y(n10415));
  AOI21X1 g07179(.A0(n10414), .A1(P2_STATE2_REG_3__SCAN_IN), .B0(n10415), .Y(n10416));
  NAND3X1 g07180(.A(n10416), .B(n10413), .C(n9740), .Y(n10417));
  NAND2X1 g07181(.A(n10417), .B(P2_INSTQUEUE_REG_7__7__SCAN_IN), .Y(n10418));
  INVX1   g07182(.A(n10406), .Y(n10419));
  OAI22X1 g07183(.A0(n9853), .A1(n10419), .B0(n10414), .B1(n9854), .Y(n10420));
  AOI21X1 g07184(.A0(n10407), .A1(n9847), .B0(n10420), .Y(n10421));
  NAND3X1 g07185(.A(n10421), .B(n10418), .C(n10411), .Y(P2_U3111));
  NAND3X1 g07186(.A(n10410), .B(n9861), .C(n9740), .Y(n10423));
  NAND2X1 g07187(.A(n10417), .B(P2_INSTQUEUE_REG_7__6__SCAN_IN), .Y(n10424));
  OAI22X1 g07188(.A0(n9872), .A1(n10419), .B0(n10414), .B1(n9873), .Y(n10425));
  AOI21X1 g07189(.A0(n10407), .A1(n9867), .B0(n10425), .Y(n10426));
  NAND3X1 g07190(.A(n10426), .B(n10424), .C(n10423), .Y(P2_U3110));
  NAND3X1 g07191(.A(n10410), .B(n9880), .C(n9740), .Y(n10428));
  NAND2X1 g07192(.A(n10417), .B(P2_INSTQUEUE_REG_7__5__SCAN_IN), .Y(n10429));
  OAI22X1 g07193(.A0(n9891), .A1(n10419), .B0(n10414), .B1(n9892), .Y(n10430));
  AOI21X1 g07194(.A0(n10407), .A1(n9886), .B0(n10430), .Y(n10431));
  NAND3X1 g07195(.A(n10431), .B(n10429), .C(n10428), .Y(P2_U3109));
  NAND3X1 g07196(.A(n10410), .B(n9899), .C(n9740), .Y(n10433));
  NAND2X1 g07197(.A(n10417), .B(P2_INSTQUEUE_REG_7__4__SCAN_IN), .Y(n10434));
  OAI22X1 g07198(.A0(n9910), .A1(n10419), .B0(n10414), .B1(n9911), .Y(n10435));
  AOI21X1 g07199(.A0(n10407), .A1(n9905), .B0(n10435), .Y(n10436));
  NAND3X1 g07200(.A(n10436), .B(n10434), .C(n10433), .Y(P2_U3108));
  NAND3X1 g07201(.A(n10410), .B(n9918), .C(n9740), .Y(n10438));
  NAND2X1 g07202(.A(n10417), .B(P2_INSTQUEUE_REG_7__3__SCAN_IN), .Y(n10439));
  OAI22X1 g07203(.A0(n9929), .A1(n10419), .B0(n10414), .B1(n9930), .Y(n10440));
  AOI21X1 g07204(.A0(n10407), .A1(n9924), .B0(n10440), .Y(n10441));
  NAND3X1 g07205(.A(n10441), .B(n10439), .C(n10438), .Y(P2_U3107));
  NAND3X1 g07206(.A(n10410), .B(n9937), .C(n9740), .Y(n10443));
  NAND2X1 g07207(.A(n10417), .B(P2_INSTQUEUE_REG_7__2__SCAN_IN), .Y(n10444));
  OAI22X1 g07208(.A0(n9948), .A1(n10419), .B0(n10414), .B1(n9949), .Y(n10445));
  AOI21X1 g07209(.A0(n10407), .A1(n9943), .B0(n10445), .Y(n10446));
  NAND3X1 g07210(.A(n10446), .B(n10444), .C(n10443), .Y(P2_U3106));
  NAND3X1 g07211(.A(n10410), .B(n9956), .C(n9740), .Y(n10448));
  NAND2X1 g07212(.A(n10417), .B(P2_INSTQUEUE_REG_7__1__SCAN_IN), .Y(n10449));
  OAI22X1 g07213(.A0(n9967), .A1(n10419), .B0(n10414), .B1(n9968), .Y(n10450));
  AOI21X1 g07214(.A0(n10407), .A1(n9962), .B0(n10450), .Y(n10451));
  NAND3X1 g07215(.A(n10451), .B(n10449), .C(n10448), .Y(P2_U3105));
  NAND3X1 g07216(.A(n10410), .B(n9975), .C(n9740), .Y(n10453));
  NAND2X1 g07217(.A(n10417), .B(P2_INSTQUEUE_REG_7__0__SCAN_IN), .Y(n10454));
  OAI22X1 g07218(.A0(n9986), .A1(n10419), .B0(n10414), .B1(n9987), .Y(n10455));
  AOI21X1 g07219(.A0(n10407), .A1(n9981), .B0(n10455), .Y(n10456));
  NAND3X1 g07220(.A(n10456), .B(n10454), .C(n10453), .Y(P2_U3104));
  NOR4X1  g07221(.A(n9208), .B(n9223), .C(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .D(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Y(n10458));
  NOR3X1  g07222(.A(n9992), .B(n9815), .C(n9633), .Y(n10459));
  OAI21X1 g07223(.A0(n10459), .A1(n10458), .B0(P2_STATE2_REG_2__SCAN_IN), .Y(n10460));
  NOR4X1  g07224(.A(n9817), .B(n9816), .C(n9786), .D(n9818), .Y(n10461));
  INVX1   g07225(.A(n10461), .Y(n10462));
  NOR2X1  g07226(.A(n10462), .B(n9779), .Y(n10463));
  NOR4X1  g07227(.A(n9811), .B(n9996), .C(n9771), .D(n10350), .Y(n10464));
  NOR3X1  g07228(.A(n10407), .B(n10464), .C(n9759), .Y(n10466));
  OAI21X1 g07229(.A0(n10466), .A1(n9757), .B0(n10463), .Y(n10467));
  NAND2X1 g07230(.A(n10467), .B(n10460), .Y(n10468));
  NAND3X1 g07231(.A(n10468), .B(n9744), .C(n9740), .Y(n10469));
  NOR4X1  g07232(.A(n10464), .B(n9759), .C(n9836), .D(n10407), .Y(n10470));
  OAI22X1 g07233(.A0(n10462), .A1(n9779), .B0(n9757), .B1(n10470), .Y(n10471));
  INVX1   g07234(.A(n10458), .Y(n10472));
  NOR3X1  g07235(.A(n10459), .B(n10458), .C(n9700), .Y(n10473));
  AOI21X1 g07236(.A0(n10472), .A1(P2_STATE2_REG_3__SCAN_IN), .B0(n10473), .Y(n10474));
  NAND3X1 g07237(.A(n10474), .B(n10471), .C(n9740), .Y(n10475));
  NAND2X1 g07238(.A(n10475), .B(P2_INSTQUEUE_REG_6__7__SCAN_IN), .Y(n10476));
  INVX1   g07239(.A(n10407), .Y(n10477));
  OAI22X1 g07240(.A0(n10472), .A1(n9854), .B0(n9853), .B1(n10477), .Y(n10478));
  AOI21X1 g07241(.A0(n10464), .A1(n9847), .B0(n10478), .Y(n10479));
  NAND3X1 g07242(.A(n10479), .B(n10476), .C(n10469), .Y(P2_U3103));
  NAND3X1 g07243(.A(n10468), .B(n9861), .C(n9740), .Y(n10481));
  NAND2X1 g07244(.A(n10475), .B(P2_INSTQUEUE_REG_6__6__SCAN_IN), .Y(n10482));
  OAI22X1 g07245(.A0(n10472), .A1(n9873), .B0(n9872), .B1(n10477), .Y(n10483));
  AOI21X1 g07246(.A0(n10464), .A1(n9867), .B0(n10483), .Y(n10484));
  NAND3X1 g07247(.A(n10484), .B(n10482), .C(n10481), .Y(P2_U3102));
  NAND3X1 g07248(.A(n10468), .B(n9880), .C(n9740), .Y(n10486));
  NAND2X1 g07249(.A(n10475), .B(P2_INSTQUEUE_REG_6__5__SCAN_IN), .Y(n10487));
  OAI22X1 g07250(.A0(n10472), .A1(n9892), .B0(n9891), .B1(n10477), .Y(n10488));
  AOI21X1 g07251(.A0(n10464), .A1(n9886), .B0(n10488), .Y(n10489));
  NAND3X1 g07252(.A(n10489), .B(n10487), .C(n10486), .Y(P2_U3101));
  NAND3X1 g07253(.A(n10468), .B(n9899), .C(n9740), .Y(n10491));
  NAND2X1 g07254(.A(n10475), .B(P2_INSTQUEUE_REG_6__4__SCAN_IN), .Y(n10492));
  OAI22X1 g07255(.A0(n10472), .A1(n9911), .B0(n9910), .B1(n10477), .Y(n10493));
  AOI21X1 g07256(.A0(n10464), .A1(n9905), .B0(n10493), .Y(n10494));
  NAND3X1 g07257(.A(n10494), .B(n10492), .C(n10491), .Y(P2_U3100));
  NAND3X1 g07258(.A(n10468), .B(n9918), .C(n9740), .Y(n10496));
  NAND2X1 g07259(.A(n10475), .B(P2_INSTQUEUE_REG_6__3__SCAN_IN), .Y(n10497));
  OAI22X1 g07260(.A0(n10472), .A1(n9930), .B0(n9929), .B1(n10477), .Y(n10498));
  AOI21X1 g07261(.A0(n10464), .A1(n9924), .B0(n10498), .Y(n10499));
  NAND3X1 g07262(.A(n10499), .B(n10497), .C(n10496), .Y(P2_U3099));
  NAND3X1 g07263(.A(n10468), .B(n9937), .C(n9740), .Y(n10501));
  NAND2X1 g07264(.A(n10475), .B(P2_INSTQUEUE_REG_6__2__SCAN_IN), .Y(n10502));
  OAI22X1 g07265(.A0(n10472), .A1(n9949), .B0(n9948), .B1(n10477), .Y(n10503));
  AOI21X1 g07266(.A0(n10464), .A1(n9943), .B0(n10503), .Y(n10504));
  NAND3X1 g07267(.A(n10504), .B(n10502), .C(n10501), .Y(P2_U3098));
  NAND3X1 g07268(.A(n10468), .B(n9956), .C(n9740), .Y(n10506));
  NAND2X1 g07269(.A(n10475), .B(P2_INSTQUEUE_REG_6__1__SCAN_IN), .Y(n10507));
  OAI22X1 g07270(.A0(n10472), .A1(n9968), .B0(n9967), .B1(n10477), .Y(n10508));
  AOI21X1 g07271(.A0(n10464), .A1(n9962), .B0(n10508), .Y(n10509));
  NAND3X1 g07272(.A(n10509), .B(n10507), .C(n10506), .Y(P2_U3097));
  NAND3X1 g07273(.A(n10468), .B(n9975), .C(n9740), .Y(n10511));
  NAND2X1 g07274(.A(n10475), .B(P2_INSTQUEUE_REG_6__0__SCAN_IN), .Y(n10512));
  OAI22X1 g07275(.A0(n10472), .A1(n9987), .B0(n9986), .B1(n10477), .Y(n10513));
  AOI21X1 g07276(.A0(n10464), .A1(n9981), .B0(n10513), .Y(n10514));
  NAND3X1 g07277(.A(n10514), .B(n10512), .C(n10511), .Y(P2_U3096));
  NOR4X1  g07278(.A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n9223), .C(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .D(n9209), .Y(n10516));
  NOR3X1  g07279(.A(n10052), .B(n9815), .C(n9633), .Y(n10517));
  OAI21X1 g07280(.A0(n10517), .A1(n10516), .B0(P2_STATE2_REG_2__SCAN_IN), .Y(n10518));
  NAND3X1 g07281(.A(n9208), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C(n9221), .Y(n10519));
  NOR4X1  g07282(.A(n9811), .B(n9996), .C(n9772), .D(n10350), .Y(n10520));
  NOR3X1  g07283(.A(n10464), .B(n10520), .C(n9759), .Y(n10522));
  NOR2X1  g07284(.A(n10522), .B(n9757), .Y(n10523));
  OAI21X1 g07285(.A0(n10523), .A1(n10519), .B0(n10518), .Y(n10524));
  NAND3X1 g07286(.A(n10524), .B(n9744), .C(n9740), .Y(n10525));
  NOR4X1  g07287(.A(n10520), .B(n9759), .C(n9836), .D(n10464), .Y(n10526));
  OAI21X1 g07288(.A0(n10526), .A1(n9757), .B0(n10519), .Y(n10527));
  INVX1   g07289(.A(n10516), .Y(n10528));
  NOR3X1  g07290(.A(n10517), .B(n10516), .C(n9700), .Y(n10529));
  AOI21X1 g07291(.A0(n10528), .A1(P2_STATE2_REG_3__SCAN_IN), .B0(n10529), .Y(n10530));
  NAND3X1 g07292(.A(n10530), .B(n10527), .C(n9740), .Y(n10531));
  NAND2X1 g07293(.A(n10531), .B(P2_INSTQUEUE_REG_5__7__SCAN_IN), .Y(n10532));
  INVX1   g07294(.A(n10464), .Y(n10533));
  OAI22X1 g07295(.A0(n10528), .A1(n9854), .B0(n9853), .B1(n10533), .Y(n10534));
  AOI21X1 g07296(.A0(n10520), .A1(n9847), .B0(n10534), .Y(n10535));
  NAND3X1 g07297(.A(n10535), .B(n10532), .C(n10525), .Y(P2_U3095));
  NAND3X1 g07298(.A(n10524), .B(n9861), .C(n9740), .Y(n10537));
  NAND2X1 g07299(.A(n10531), .B(P2_INSTQUEUE_REG_5__6__SCAN_IN), .Y(n10538));
  OAI22X1 g07300(.A0(n10528), .A1(n9873), .B0(n9872), .B1(n10533), .Y(n10539));
  AOI21X1 g07301(.A0(n10520), .A1(n9867), .B0(n10539), .Y(n10540));
  NAND3X1 g07302(.A(n10540), .B(n10538), .C(n10537), .Y(P2_U3094));
  NAND3X1 g07303(.A(n10524), .B(n9880), .C(n9740), .Y(n10542));
  NAND2X1 g07304(.A(n10531), .B(P2_INSTQUEUE_REG_5__5__SCAN_IN), .Y(n10543));
  OAI22X1 g07305(.A0(n10528), .A1(n9892), .B0(n9891), .B1(n10533), .Y(n10544));
  AOI21X1 g07306(.A0(n10520), .A1(n9886), .B0(n10544), .Y(n10545));
  NAND3X1 g07307(.A(n10545), .B(n10543), .C(n10542), .Y(P2_U3093));
  NAND3X1 g07308(.A(n10524), .B(n9899), .C(n9740), .Y(n10547));
  NAND2X1 g07309(.A(n10531), .B(P2_INSTQUEUE_REG_5__4__SCAN_IN), .Y(n10548));
  OAI22X1 g07310(.A0(n10528), .A1(n9911), .B0(n9910), .B1(n10533), .Y(n10549));
  AOI21X1 g07311(.A0(n10520), .A1(n9905), .B0(n10549), .Y(n10550));
  NAND3X1 g07312(.A(n10550), .B(n10548), .C(n10547), .Y(P2_U3092));
  NAND3X1 g07313(.A(n10524), .B(n9918), .C(n9740), .Y(n10552));
  NAND2X1 g07314(.A(n10531), .B(P2_INSTQUEUE_REG_5__3__SCAN_IN), .Y(n10553));
  OAI22X1 g07315(.A0(n10528), .A1(n9930), .B0(n9929), .B1(n10533), .Y(n10554));
  AOI21X1 g07316(.A0(n10520), .A1(n9924), .B0(n10554), .Y(n10555));
  NAND3X1 g07317(.A(n10555), .B(n10553), .C(n10552), .Y(P2_U3091));
  NAND3X1 g07318(.A(n10524), .B(n9937), .C(n9740), .Y(n10557));
  NAND2X1 g07319(.A(n10531), .B(P2_INSTQUEUE_REG_5__2__SCAN_IN), .Y(n10558));
  OAI22X1 g07320(.A0(n10528), .A1(n9949), .B0(n9948), .B1(n10533), .Y(n10559));
  AOI21X1 g07321(.A0(n10520), .A1(n9943), .B0(n10559), .Y(n10560));
  NAND3X1 g07322(.A(n10560), .B(n10558), .C(n10557), .Y(P2_U3090));
  NAND3X1 g07323(.A(n10524), .B(n9956), .C(n9740), .Y(n10562));
  NAND2X1 g07324(.A(n10531), .B(P2_INSTQUEUE_REG_5__1__SCAN_IN), .Y(n10563));
  OAI22X1 g07325(.A0(n10528), .A1(n9968), .B0(n9967), .B1(n10533), .Y(n10564));
  AOI21X1 g07326(.A0(n10520), .A1(n9962), .B0(n10564), .Y(n10565));
  NAND3X1 g07327(.A(n10565), .B(n10563), .C(n10562), .Y(P2_U3089));
  NAND3X1 g07328(.A(n10524), .B(n9975), .C(n9740), .Y(n10567));
  NAND2X1 g07329(.A(n10531), .B(P2_INSTQUEUE_REG_5__0__SCAN_IN), .Y(n10568));
  OAI22X1 g07330(.A0(n10528), .A1(n9987), .B0(n9986), .B1(n10533), .Y(n10569));
  AOI21X1 g07331(.A0(n10520), .A1(n9981), .B0(n10569), .Y(n10570));
  NAND3X1 g07332(.A(n10570), .B(n10568), .C(n10567), .Y(P2_U3088));
  NOR4X1  g07333(.A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n9223), .C(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .D(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Y(n10572));
  NOR3X1  g07334(.A(n10109), .B(n9815), .C(n9633), .Y(n10573));
  OAI21X1 g07335(.A0(n10573), .A1(n10572), .B0(P2_STATE2_REG_2__SCAN_IN), .Y(n10574));
  NOR2X1  g07336(.A(n10462), .B(n9780), .Y(n10575));
  NOR4X1  g07337(.A(n9810), .B(n9784), .C(n9771), .D(n10350), .Y(n10576));
  NOR3X1  g07338(.A(n10520), .B(n10576), .C(n9759), .Y(n10578));
  OAI21X1 g07339(.A0(n10578), .A1(n9757), .B0(n10575), .Y(n10579));
  NAND2X1 g07340(.A(n10579), .B(n10574), .Y(n10580));
  NAND3X1 g07341(.A(n10580), .B(n9744), .C(n9740), .Y(n10581));
  NOR4X1  g07342(.A(n10576), .B(n9759), .C(n9836), .D(n10520), .Y(n10582));
  OAI22X1 g07343(.A0(n10462), .A1(n9780), .B0(n9757), .B1(n10582), .Y(n10583));
  INVX1   g07344(.A(n10572), .Y(n10584));
  NOR3X1  g07345(.A(n10573), .B(n10572), .C(n9700), .Y(n10585));
  AOI21X1 g07346(.A0(n10584), .A1(P2_STATE2_REG_3__SCAN_IN), .B0(n10585), .Y(n10586));
  NAND3X1 g07347(.A(n10586), .B(n10583), .C(n9740), .Y(n10587));
  NAND2X1 g07348(.A(n10587), .B(P2_INSTQUEUE_REG_4__7__SCAN_IN), .Y(n10588));
  INVX1   g07349(.A(n10520), .Y(n10589));
  OAI22X1 g07350(.A0(n10584), .A1(n9854), .B0(n9853), .B1(n10589), .Y(n10590));
  AOI21X1 g07351(.A0(n10576), .A1(n9847), .B0(n10590), .Y(n10591));
  NAND3X1 g07352(.A(n10591), .B(n10588), .C(n10581), .Y(P2_U3087));
  NAND3X1 g07353(.A(n10580), .B(n9861), .C(n9740), .Y(n10593));
  NAND2X1 g07354(.A(n10587), .B(P2_INSTQUEUE_REG_4__6__SCAN_IN), .Y(n10594));
  OAI22X1 g07355(.A0(n10584), .A1(n9873), .B0(n9872), .B1(n10589), .Y(n10595));
  AOI21X1 g07356(.A0(n10576), .A1(n9867), .B0(n10595), .Y(n10596));
  NAND3X1 g07357(.A(n10596), .B(n10594), .C(n10593), .Y(P2_U3086));
  NAND3X1 g07358(.A(n10580), .B(n9880), .C(n9740), .Y(n10598));
  NAND2X1 g07359(.A(n10587), .B(P2_INSTQUEUE_REG_4__5__SCAN_IN), .Y(n10599));
  OAI22X1 g07360(.A0(n10584), .A1(n9892), .B0(n9891), .B1(n10589), .Y(n10600));
  AOI21X1 g07361(.A0(n10576), .A1(n9886), .B0(n10600), .Y(n10601));
  NAND3X1 g07362(.A(n10601), .B(n10599), .C(n10598), .Y(P2_U3085));
  NAND3X1 g07363(.A(n10580), .B(n9899), .C(n9740), .Y(n10603));
  NAND2X1 g07364(.A(n10587), .B(P2_INSTQUEUE_REG_4__4__SCAN_IN), .Y(n10604));
  OAI22X1 g07365(.A0(n10584), .A1(n9911), .B0(n9910), .B1(n10589), .Y(n10605));
  AOI21X1 g07366(.A0(n10576), .A1(n9905), .B0(n10605), .Y(n10606));
  NAND3X1 g07367(.A(n10606), .B(n10604), .C(n10603), .Y(P2_U3084));
  NAND3X1 g07368(.A(n10580), .B(n9918), .C(n9740), .Y(n10608));
  NAND2X1 g07369(.A(n10587), .B(P2_INSTQUEUE_REG_4__3__SCAN_IN), .Y(n10609));
  OAI22X1 g07370(.A0(n10584), .A1(n9930), .B0(n9929), .B1(n10589), .Y(n10610));
  AOI21X1 g07371(.A0(n10576), .A1(n9924), .B0(n10610), .Y(n10611));
  NAND3X1 g07372(.A(n10611), .B(n10609), .C(n10608), .Y(P2_U3083));
  NAND3X1 g07373(.A(n10580), .B(n9937), .C(n9740), .Y(n10613));
  NAND2X1 g07374(.A(n10587), .B(P2_INSTQUEUE_REG_4__2__SCAN_IN), .Y(n10614));
  OAI22X1 g07375(.A0(n10584), .A1(n9949), .B0(n9948), .B1(n10589), .Y(n10615));
  AOI21X1 g07376(.A0(n10576), .A1(n9943), .B0(n10615), .Y(n10616));
  NAND3X1 g07377(.A(n10616), .B(n10614), .C(n10613), .Y(P2_U3082));
  NAND3X1 g07378(.A(n10580), .B(n9956), .C(n9740), .Y(n10618));
  NAND2X1 g07379(.A(n10587), .B(P2_INSTQUEUE_REG_4__1__SCAN_IN), .Y(n10619));
  OAI22X1 g07380(.A0(n10584), .A1(n9968), .B0(n9967), .B1(n10589), .Y(n10620));
  AOI21X1 g07381(.A0(n10576), .A1(n9962), .B0(n10620), .Y(n10621));
  NAND3X1 g07382(.A(n10621), .B(n10619), .C(n10618), .Y(P2_U3081));
  NAND3X1 g07383(.A(n10580), .B(n9975), .C(n9740), .Y(n10623));
  NAND2X1 g07384(.A(n10587), .B(P2_INSTQUEUE_REG_4__0__SCAN_IN), .Y(n10624));
  OAI22X1 g07385(.A0(n10584), .A1(n9987), .B0(n9986), .B1(n10589), .Y(n10625));
  AOI21X1 g07386(.A0(n10576), .A1(n9981), .B0(n10625), .Y(n10626));
  NAND3X1 g07387(.A(n10626), .B(n10624), .C(n10623), .Y(P2_U3080));
  NOR3X1  g07388(.A(n9745), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .Y(n10628));
  NOR3X1  g07389(.A(n9753), .B(n9815), .C(n9794), .Y(n10629));
  OAI21X1 g07390(.A0(n10629), .A1(n10628), .B0(P2_STATE2_REG_2__SCAN_IN), .Y(n10630));
  NAND3X1 g07391(.A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n9223), .C(n9221), .Y(n10631));
  NOR4X1  g07392(.A(n9810), .B(n9784), .C(n9772), .D(n10350), .Y(n10632));
  NOR3X1  g07393(.A(n10576), .B(n10632), .C(n9759), .Y(n10634));
  NOR2X1  g07394(.A(n10634), .B(n9757), .Y(n10635));
  OAI21X1 g07395(.A0(n10635), .A1(n10631), .B0(n10630), .Y(n10636));
  NAND3X1 g07396(.A(n10636), .B(n9744), .C(n9740), .Y(n10637));
  NOR4X1  g07397(.A(n10632), .B(n9759), .C(n9836), .D(n10576), .Y(n10638));
  OAI21X1 g07398(.A0(n10638), .A1(n9757), .B0(n10631), .Y(n10639));
  INVX1   g07399(.A(n10628), .Y(n10640));
  NOR3X1  g07400(.A(n10629), .B(n10628), .C(n9700), .Y(n10641));
  AOI21X1 g07401(.A0(n10640), .A1(P2_STATE2_REG_3__SCAN_IN), .B0(n10641), .Y(n10642));
  NAND3X1 g07402(.A(n10642), .B(n10639), .C(n9740), .Y(n10643));
  NAND2X1 g07403(.A(n10643), .B(P2_INSTQUEUE_REG_3__7__SCAN_IN), .Y(n10644));
  INVX1   g07404(.A(n10576), .Y(n10645));
  OAI22X1 g07405(.A0(n10640), .A1(n9854), .B0(n9853), .B1(n10645), .Y(n10646));
  AOI21X1 g07406(.A0(n10632), .A1(n9847), .B0(n10646), .Y(n10647));
  NAND3X1 g07407(.A(n10647), .B(n10644), .C(n10637), .Y(P2_U3079));
  NAND3X1 g07408(.A(n10636), .B(n9861), .C(n9740), .Y(n10649));
  NAND2X1 g07409(.A(n10643), .B(P2_INSTQUEUE_REG_3__6__SCAN_IN), .Y(n10650));
  OAI22X1 g07410(.A0(n10640), .A1(n9873), .B0(n9872), .B1(n10645), .Y(n10651));
  AOI21X1 g07411(.A0(n10632), .A1(n9867), .B0(n10651), .Y(n10652));
  NAND3X1 g07412(.A(n10652), .B(n10650), .C(n10649), .Y(P2_U3078));
  NAND3X1 g07413(.A(n10636), .B(n9880), .C(n9740), .Y(n10654));
  NAND2X1 g07414(.A(n10643), .B(P2_INSTQUEUE_REG_3__5__SCAN_IN), .Y(n10655));
  OAI22X1 g07415(.A0(n10640), .A1(n9892), .B0(n9891), .B1(n10645), .Y(n10656));
  AOI21X1 g07416(.A0(n10632), .A1(n9886), .B0(n10656), .Y(n10657));
  NAND3X1 g07417(.A(n10657), .B(n10655), .C(n10654), .Y(P2_U3077));
  NAND3X1 g07418(.A(n10636), .B(n9899), .C(n9740), .Y(n10659));
  NAND2X1 g07419(.A(n10643), .B(P2_INSTQUEUE_REG_3__4__SCAN_IN), .Y(n10660));
  OAI22X1 g07420(.A0(n10640), .A1(n9911), .B0(n9910), .B1(n10645), .Y(n10661));
  AOI21X1 g07421(.A0(n10632), .A1(n9905), .B0(n10661), .Y(n10662));
  NAND3X1 g07422(.A(n10662), .B(n10660), .C(n10659), .Y(P2_U3076));
  NAND3X1 g07423(.A(n10636), .B(n9918), .C(n9740), .Y(n10664));
  NAND2X1 g07424(.A(n10643), .B(P2_INSTQUEUE_REG_3__3__SCAN_IN), .Y(n10665));
  OAI22X1 g07425(.A0(n10640), .A1(n9930), .B0(n9929), .B1(n10645), .Y(n10666));
  AOI21X1 g07426(.A0(n10632), .A1(n9924), .B0(n10666), .Y(n10667));
  NAND3X1 g07427(.A(n10667), .B(n10665), .C(n10664), .Y(P2_U3075));
  NAND3X1 g07428(.A(n10636), .B(n9937), .C(n9740), .Y(n10669));
  NAND2X1 g07429(.A(n10643), .B(P2_INSTQUEUE_REG_3__2__SCAN_IN), .Y(n10670));
  OAI22X1 g07430(.A0(n10640), .A1(n9949), .B0(n9948), .B1(n10645), .Y(n10671));
  AOI21X1 g07431(.A0(n10632), .A1(n9943), .B0(n10671), .Y(n10672));
  NAND3X1 g07432(.A(n10672), .B(n10670), .C(n10669), .Y(P2_U3074));
  NAND3X1 g07433(.A(n10636), .B(n9956), .C(n9740), .Y(n10674));
  NAND2X1 g07434(.A(n10643), .B(P2_INSTQUEUE_REG_3__1__SCAN_IN), .Y(n10675));
  OAI22X1 g07435(.A0(n10640), .A1(n9968), .B0(n9967), .B1(n10645), .Y(n10676));
  AOI21X1 g07436(.A0(n10632), .A1(n9962), .B0(n10676), .Y(n10677));
  NAND3X1 g07437(.A(n10677), .B(n10675), .C(n10674), .Y(P2_U3073));
  NAND3X1 g07438(.A(n10636), .B(n9975), .C(n9740), .Y(n10679));
  NAND2X1 g07439(.A(n10643), .B(P2_INSTQUEUE_REG_3__0__SCAN_IN), .Y(n10680));
  OAI22X1 g07440(.A0(n10640), .A1(n9987), .B0(n9986), .B1(n10645), .Y(n10681));
  AOI21X1 g07441(.A0(n10632), .A1(n9981), .B0(n10681), .Y(n10682));
  NAND3X1 g07442(.A(n10682), .B(n10680), .C(n10679), .Y(P2_U3072));
  NOR4X1  g07443(.A(n9208), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .D(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Y(n10684));
  NOR3X1  g07444(.A(n9992), .B(n9815), .C(n9794), .Y(n10685));
  OAI21X1 g07445(.A0(n10685), .A1(n10684), .B0(P2_STATE2_REG_2__SCAN_IN), .Y(n10686));
  NOR3X1  g07446(.A(n9779), .B(n9820), .C(n9787), .Y(n10687));
  NOR4X1  g07447(.A(n9810), .B(n9996), .C(n9771), .D(n10350), .Y(n10688));
  NOR3X1  g07448(.A(n10632), .B(n10688), .C(n9759), .Y(n10690));
  OAI21X1 g07449(.A0(n10690), .A1(n9757), .B0(n10687), .Y(n10691));
  NAND2X1 g07450(.A(n10691), .B(n10686), .Y(n10692));
  NAND3X1 g07451(.A(n10692), .B(n9744), .C(n9740), .Y(n10693));
  NOR4X1  g07452(.A(n9817), .B(n9816), .C(n9787), .D(n9818), .Y(n10694));
  INVX1   g07453(.A(n10694), .Y(n10695));
  NOR4X1  g07454(.A(n10688), .B(n9759), .C(n9836), .D(n10632), .Y(n10696));
  OAI22X1 g07455(.A0(n10695), .A1(n9779), .B0(n9757), .B1(n10696), .Y(n10697));
  INVX1   g07456(.A(n10684), .Y(n10698));
  NOR3X1  g07457(.A(n10685), .B(n10684), .C(n9700), .Y(n10699));
  AOI21X1 g07458(.A0(n10698), .A1(P2_STATE2_REG_3__SCAN_IN), .B0(n10699), .Y(n10700));
  NAND3X1 g07459(.A(n10700), .B(n10697), .C(n9740), .Y(n10701));
  NAND2X1 g07460(.A(n10701), .B(P2_INSTQUEUE_REG_2__7__SCAN_IN), .Y(n10702));
  INVX1   g07461(.A(n10632), .Y(n10703));
  OAI22X1 g07462(.A0(n10698), .A1(n9854), .B0(n9853), .B1(n10703), .Y(n10704));
  AOI21X1 g07463(.A0(n10688), .A1(n9847), .B0(n10704), .Y(n10705));
  NAND3X1 g07464(.A(n10705), .B(n10702), .C(n10693), .Y(P2_U3071));
  NAND3X1 g07465(.A(n10692), .B(n9861), .C(n9740), .Y(n10707));
  NAND2X1 g07466(.A(n10701), .B(P2_INSTQUEUE_REG_2__6__SCAN_IN), .Y(n10708));
  OAI22X1 g07467(.A0(n10698), .A1(n9873), .B0(n9872), .B1(n10703), .Y(n10709));
  AOI21X1 g07468(.A0(n10688), .A1(n9867), .B0(n10709), .Y(n10710));
  NAND3X1 g07469(.A(n10710), .B(n10708), .C(n10707), .Y(P2_U3070));
  NAND3X1 g07470(.A(n10692), .B(n9880), .C(n9740), .Y(n10712));
  NAND2X1 g07471(.A(n10701), .B(P2_INSTQUEUE_REG_2__5__SCAN_IN), .Y(n10713));
  OAI22X1 g07472(.A0(n10698), .A1(n9892), .B0(n9891), .B1(n10703), .Y(n10714));
  AOI21X1 g07473(.A0(n10688), .A1(n9886), .B0(n10714), .Y(n10715));
  NAND3X1 g07474(.A(n10715), .B(n10713), .C(n10712), .Y(P2_U3069));
  NAND3X1 g07475(.A(n10692), .B(n9899), .C(n9740), .Y(n10717));
  NAND2X1 g07476(.A(n10701), .B(P2_INSTQUEUE_REG_2__4__SCAN_IN), .Y(n10718));
  OAI22X1 g07477(.A0(n10698), .A1(n9911), .B0(n9910), .B1(n10703), .Y(n10719));
  AOI21X1 g07478(.A0(n10688), .A1(n9905), .B0(n10719), .Y(n10720));
  NAND3X1 g07479(.A(n10720), .B(n10718), .C(n10717), .Y(P2_U3068));
  NAND3X1 g07480(.A(n10692), .B(n9918), .C(n9740), .Y(n10722));
  NAND2X1 g07481(.A(n10701), .B(P2_INSTQUEUE_REG_2__3__SCAN_IN), .Y(n10723));
  OAI22X1 g07482(.A0(n10698), .A1(n9930), .B0(n9929), .B1(n10703), .Y(n10724));
  AOI21X1 g07483(.A0(n10688), .A1(n9924), .B0(n10724), .Y(n10725));
  NAND3X1 g07484(.A(n10725), .B(n10723), .C(n10722), .Y(P2_U3067));
  NAND3X1 g07485(.A(n10692), .B(n9937), .C(n9740), .Y(n10727));
  NAND2X1 g07486(.A(n10701), .B(P2_INSTQUEUE_REG_2__2__SCAN_IN), .Y(n10728));
  OAI22X1 g07487(.A0(n10698), .A1(n9949), .B0(n9948), .B1(n10703), .Y(n10729));
  AOI21X1 g07488(.A0(n10688), .A1(n9943), .B0(n10729), .Y(n10730));
  NAND3X1 g07489(.A(n10730), .B(n10728), .C(n10727), .Y(P2_U3066));
  NAND3X1 g07490(.A(n10692), .B(n9956), .C(n9740), .Y(n10732));
  NAND2X1 g07491(.A(n10701), .B(P2_INSTQUEUE_REG_2__1__SCAN_IN), .Y(n10733));
  OAI22X1 g07492(.A0(n10698), .A1(n9968), .B0(n9967), .B1(n10703), .Y(n10734));
  AOI21X1 g07493(.A0(n10688), .A1(n9962), .B0(n10734), .Y(n10735));
  NAND3X1 g07494(.A(n10735), .B(n10733), .C(n10732), .Y(P2_U3065));
  NAND3X1 g07495(.A(n10692), .B(n9975), .C(n9740), .Y(n10737));
  NAND2X1 g07496(.A(n10701), .B(P2_INSTQUEUE_REG_2__0__SCAN_IN), .Y(n10738));
  OAI22X1 g07497(.A0(n10698), .A1(n9987), .B0(n9986), .B1(n10703), .Y(n10739));
  AOI21X1 g07498(.A0(n10688), .A1(n9981), .B0(n10739), .Y(n10740));
  NAND3X1 g07499(.A(n10740), .B(n10738), .C(n10737), .Y(P2_U3064));
  NOR4X1  g07500(.A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .D(n9209), .Y(n10742));
  NOR3X1  g07501(.A(n10052), .B(n9815), .C(n9794), .Y(n10743));
  OAI21X1 g07502(.A0(n10743), .A1(n10742), .B0(P2_STATE2_REG_2__SCAN_IN), .Y(n10744));
  NAND3X1 g07503(.A(n9208), .B(n9223), .C(n9221), .Y(n10745));
  NOR4X1  g07504(.A(n9810), .B(n9996), .C(n9772), .D(n10350), .Y(n10746));
  NOR3X1  g07505(.A(n10688), .B(n10746), .C(n9759), .Y(n10748));
  NOR2X1  g07506(.A(n10748), .B(n9757), .Y(n10749));
  OAI21X1 g07507(.A0(n10749), .A1(n10745), .B0(n10744), .Y(n10750));
  NAND3X1 g07508(.A(n10750), .B(n9744), .C(n9740), .Y(n10751));
  NOR4X1  g07509(.A(n10746), .B(n9759), .C(n9836), .D(n10688), .Y(n10752));
  OAI21X1 g07510(.A0(n10752), .A1(n9757), .B0(n10745), .Y(n10753));
  INVX1   g07511(.A(n10742), .Y(n10754));
  NOR3X1  g07512(.A(n10743), .B(n10742), .C(n9700), .Y(n10755));
  AOI21X1 g07513(.A0(n10754), .A1(P2_STATE2_REG_3__SCAN_IN), .B0(n10755), .Y(n10756));
  NAND3X1 g07514(.A(n10756), .B(n10753), .C(n9740), .Y(n10757));
  NAND2X1 g07515(.A(n10757), .B(P2_INSTQUEUE_REG_1__7__SCAN_IN), .Y(n10758));
  INVX1   g07516(.A(n10688), .Y(n10759));
  OAI22X1 g07517(.A0(n10754), .A1(n9854), .B0(n9853), .B1(n10759), .Y(n10760));
  AOI21X1 g07518(.A0(n10746), .A1(n9847), .B0(n10760), .Y(n10761));
  NAND3X1 g07519(.A(n10761), .B(n10758), .C(n10751), .Y(P2_U3063));
  NAND3X1 g07520(.A(n10750), .B(n9861), .C(n9740), .Y(n10763));
  NAND2X1 g07521(.A(n10757), .B(P2_INSTQUEUE_REG_1__6__SCAN_IN), .Y(n10764));
  OAI22X1 g07522(.A0(n10754), .A1(n9873), .B0(n9872), .B1(n10759), .Y(n10765));
  AOI21X1 g07523(.A0(n10746), .A1(n9867), .B0(n10765), .Y(n10766));
  NAND3X1 g07524(.A(n10766), .B(n10764), .C(n10763), .Y(P2_U3062));
  NAND3X1 g07525(.A(n10750), .B(n9880), .C(n9740), .Y(n10768));
  NAND2X1 g07526(.A(n10757), .B(P2_INSTQUEUE_REG_1__5__SCAN_IN), .Y(n10769));
  OAI22X1 g07527(.A0(n10754), .A1(n9892), .B0(n9891), .B1(n10759), .Y(n10770));
  AOI21X1 g07528(.A0(n10746), .A1(n9886), .B0(n10770), .Y(n10771));
  NAND3X1 g07529(.A(n10771), .B(n10769), .C(n10768), .Y(P2_U3061));
  NAND3X1 g07530(.A(n10750), .B(n9899), .C(n9740), .Y(n10773));
  NAND2X1 g07531(.A(n10757), .B(P2_INSTQUEUE_REG_1__4__SCAN_IN), .Y(n10774));
  OAI22X1 g07532(.A0(n10754), .A1(n9911), .B0(n9910), .B1(n10759), .Y(n10775));
  AOI21X1 g07533(.A0(n10746), .A1(n9905), .B0(n10775), .Y(n10776));
  NAND3X1 g07534(.A(n10776), .B(n10774), .C(n10773), .Y(P2_U3060));
  NAND3X1 g07535(.A(n10750), .B(n9918), .C(n9740), .Y(n10778));
  NAND2X1 g07536(.A(n10757), .B(P2_INSTQUEUE_REG_1__3__SCAN_IN), .Y(n10779));
  OAI22X1 g07537(.A0(n10754), .A1(n9930), .B0(n9929), .B1(n10759), .Y(n10780));
  AOI21X1 g07538(.A0(n10746), .A1(n9924), .B0(n10780), .Y(n10781));
  NAND3X1 g07539(.A(n10781), .B(n10779), .C(n10778), .Y(P2_U3059));
  NAND3X1 g07540(.A(n10750), .B(n9937), .C(n9740), .Y(n10783));
  NAND2X1 g07541(.A(n10757), .B(P2_INSTQUEUE_REG_1__2__SCAN_IN), .Y(n10784));
  OAI22X1 g07542(.A0(n10754), .A1(n9949), .B0(n9948), .B1(n10759), .Y(n10785));
  AOI21X1 g07543(.A0(n10746), .A1(n9943), .B0(n10785), .Y(n10786));
  NAND3X1 g07544(.A(n10786), .B(n10784), .C(n10783), .Y(P2_U3058));
  NAND3X1 g07545(.A(n10750), .B(n9956), .C(n9740), .Y(n10788));
  NAND2X1 g07546(.A(n10757), .B(P2_INSTQUEUE_REG_1__1__SCAN_IN), .Y(n10789));
  OAI22X1 g07547(.A0(n10754), .A1(n9968), .B0(n9967), .B1(n10759), .Y(n10790));
  AOI21X1 g07548(.A0(n10746), .A1(n9962), .B0(n10790), .Y(n10791));
  NAND3X1 g07549(.A(n10791), .B(n10789), .C(n10788), .Y(P2_U3057));
  NAND3X1 g07550(.A(n10750), .B(n9975), .C(n9740), .Y(n10793));
  NAND2X1 g07551(.A(n10757), .B(P2_INSTQUEUE_REG_1__0__SCAN_IN), .Y(n10794));
  OAI22X1 g07552(.A0(n10754), .A1(n9987), .B0(n9986), .B1(n10759), .Y(n10795));
  AOI21X1 g07553(.A0(n10746), .A1(n9981), .B0(n10795), .Y(n10796));
  NAND3X1 g07554(.A(n10796), .B(n10794), .C(n10793), .Y(P2_U3056));
  NOR4X1  g07555(.A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .D(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Y(n10798));
  NOR3X1  g07556(.A(n10109), .B(n9815), .C(n9794), .Y(n10799));
  OAI21X1 g07557(.A0(n10799), .A1(n10798), .B0(P2_STATE2_REG_2__SCAN_IN), .Y(n10800));
  NOR3X1  g07558(.A(n9780), .B(n9820), .C(n9787), .Y(n10801));
  NOR3X1  g07559(.A(n10746), .B(n9831), .C(n9759), .Y(n10804));
  OAI21X1 g07560(.A0(n10804), .A1(n9757), .B0(n10801), .Y(n10805));
  NAND2X1 g07561(.A(n10805), .B(n10800), .Y(n10806));
  NAND3X1 g07562(.A(n10806), .B(n9744), .C(n9740), .Y(n10807));
  NOR4X1  g07563(.A(n9831), .B(n9759), .C(n9836), .D(n10746), .Y(n10808));
  OAI22X1 g07564(.A0(n10695), .A1(n9780), .B0(n9757), .B1(n10808), .Y(n10809));
  INVX1   g07565(.A(n10798), .Y(n10810));
  NOR3X1  g07566(.A(n10799), .B(n10798), .C(n9700), .Y(n10811));
  AOI21X1 g07567(.A0(n10810), .A1(P2_STATE2_REG_3__SCAN_IN), .B0(n10811), .Y(n10812));
  NAND3X1 g07568(.A(n10812), .B(n10809), .C(n9740), .Y(n10813));
  NAND2X1 g07569(.A(n10813), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .Y(n10814));
  INVX1   g07570(.A(n10746), .Y(n10815));
  OAI22X1 g07571(.A0(n10810), .A1(n9854), .B0(n9853), .B1(n10815), .Y(n10816));
  AOI21X1 g07572(.A0(n9831), .A1(n9847), .B0(n10816), .Y(n10817));
  NAND3X1 g07573(.A(n10817), .B(n10814), .C(n10807), .Y(P2_U3055));
  NAND3X1 g07574(.A(n10806), .B(n9861), .C(n9740), .Y(n10819));
  NAND2X1 g07575(.A(n10813), .B(P2_INSTQUEUE_REG_0__6__SCAN_IN), .Y(n10820));
  OAI22X1 g07576(.A0(n10810), .A1(n9873), .B0(n9872), .B1(n10815), .Y(n10821));
  AOI21X1 g07577(.A0(n9831), .A1(n9867), .B0(n10821), .Y(n10822));
  NAND3X1 g07578(.A(n10822), .B(n10820), .C(n10819), .Y(P2_U3054));
  NAND3X1 g07579(.A(n10806), .B(n9880), .C(n9740), .Y(n10824));
  NAND2X1 g07580(.A(n10813), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .Y(n10825));
  OAI22X1 g07581(.A0(n10810), .A1(n9892), .B0(n9891), .B1(n10815), .Y(n10826));
  AOI21X1 g07582(.A0(n9831), .A1(n9886), .B0(n10826), .Y(n10827));
  NAND3X1 g07583(.A(n10827), .B(n10825), .C(n10824), .Y(P2_U3053));
  NAND3X1 g07584(.A(n10806), .B(n9899), .C(n9740), .Y(n10829));
  NAND2X1 g07585(.A(n10813), .B(P2_INSTQUEUE_REG_0__4__SCAN_IN), .Y(n10830));
  OAI22X1 g07586(.A0(n10810), .A1(n9911), .B0(n9910), .B1(n10815), .Y(n10831));
  AOI21X1 g07587(.A0(n9831), .A1(n9905), .B0(n10831), .Y(n10832));
  NAND3X1 g07588(.A(n10832), .B(n10830), .C(n10829), .Y(P2_U3052));
  NAND3X1 g07589(.A(n10806), .B(n9918), .C(n9740), .Y(n10834));
  NAND2X1 g07590(.A(n10813), .B(P2_INSTQUEUE_REG_0__3__SCAN_IN), .Y(n10835));
  OAI22X1 g07591(.A0(n10810), .A1(n9930), .B0(n9929), .B1(n10815), .Y(n10836));
  AOI21X1 g07592(.A0(n9831), .A1(n9924), .B0(n10836), .Y(n10837));
  NAND3X1 g07593(.A(n10837), .B(n10835), .C(n10834), .Y(P2_U3051));
  NAND3X1 g07594(.A(n10806), .B(n9937), .C(n9740), .Y(n10839));
  NAND2X1 g07595(.A(n10813), .B(P2_INSTQUEUE_REG_0__2__SCAN_IN), .Y(n10840));
  OAI22X1 g07596(.A0(n10810), .A1(n9949), .B0(n9948), .B1(n10815), .Y(n10841));
  AOI21X1 g07597(.A0(n9831), .A1(n9943), .B0(n10841), .Y(n10842));
  NAND3X1 g07598(.A(n10842), .B(n10840), .C(n10839), .Y(P2_U3050));
  NAND3X1 g07599(.A(n10806), .B(n9956), .C(n9740), .Y(n10844));
  NAND2X1 g07600(.A(n10813), .B(P2_INSTQUEUE_REG_0__1__SCAN_IN), .Y(n10845));
  OAI22X1 g07601(.A0(n10810), .A1(n9968), .B0(n9967), .B1(n10815), .Y(n10846));
  AOI21X1 g07602(.A0(n9831), .A1(n9962), .B0(n10846), .Y(n10847));
  NAND3X1 g07603(.A(n10847), .B(n10845), .C(n10844), .Y(P2_U3049));
  NAND3X1 g07604(.A(n10806), .B(n9975), .C(n9740), .Y(n10849));
  NAND2X1 g07605(.A(n10813), .B(P2_INSTQUEUE_REG_0__0__SCAN_IN), .Y(n10850));
  OAI22X1 g07606(.A0(n10810), .A1(n9987), .B0(n9986), .B1(n10815), .Y(n10851));
  AOI21X1 g07607(.A0(n9831), .A1(n9981), .B0(n10851), .Y(n10852));
  NAND3X1 g07608(.A(n10852), .B(n10850), .C(n10849), .Y(P2_U3048));
  NOR4X1  g07609(.A(n8720), .B(n9205), .C(n9700), .D(n9162), .Y(n10854));
  AOI21X1 g07610(.A0(n8720), .A1(P2_STATE2_REG_3__SCAN_IN), .B0(n10854), .Y(n10855));
  OAI21X1 g07611(.A0(n9732), .A1(n9621), .B0(n10855), .Y(n10856));
  INVX1   g07612(.A(n9717), .Y(n10857));
  NOR4X1  g07613(.A(n9679), .B(n9416), .C(n9311), .D(n10857), .Y(n10858));
  NAND2X1 g07614(.A(n10858), .B(n10856), .Y(n10859));
  OAI21X1 g07615(.A0(n10856), .A1(n9019), .B0(n10859), .Y(P2_U3595));
  NAND2X1 g07616(.A(n9717), .B(n9671), .Y(n10861));
  OAI21X1 g07617(.A0(n9827), .A1(n9738), .B0(n10861), .Y(n10862));
  NAND2X1 g07618(.A(n10862), .B(n10856), .Y(n10863));
  OAI21X1 g07619(.A0(n10856), .A1(n8724), .B0(n10863), .Y(P2_U3596));
  NOR3X1  g07620(.A(n9203), .B(n9197), .C(n9205), .Y(n10865));
  OAI22X1 g07621(.A0(n9738), .A1(n9811), .B0(n10857), .B1(n9644), .Y(n10866));
  OAI21X1 g07622(.A0(n10866), .A1(n10865), .B0(n10856), .Y(n10867));
  OAI21X1 g07623(.A0(n10856), .A1(n8727), .B0(n10867), .Y(P2_U3599));
  AOI22X1 g07624(.A0(n9730), .A1(n9996), .B0(n9717), .B1(n9611), .Y(n10869));
  OAI21X1 g07625(.A0(n9249), .A1(n9205), .B0(n10869), .Y(n10870));
  NAND2X1 g07626(.A(n10870), .B(n10856), .Y(n10871));
  OAI21X1 g07627(.A0(n10856), .A1(n8732), .B0(n10871), .Y(P2_U3600));
  AOI22X1 g07628(.A0(n9730), .A1(n9772), .B0(n9717), .B1(n9617), .Y(n10873));
  OAI21X1 g07629(.A0(n9216), .A1(n9205), .B0(n10873), .Y(n10874));
  NAND2X1 g07630(.A(n10874), .B(n10856), .Y(n10875));
  OAI21X1 g07631(.A0(n10856), .A1(n8721), .B0(n10875), .Y(P2_U3601));
  NOR4X1  g07632(.A(n8720), .B(n9205), .C(n9700), .D(n9259), .Y(n10877));
  NOR4X1  g07633(.A(n10854), .B(n9740), .C(n9227), .D(n10877), .Y(P2_U3047));
  NOR3X1  g07634(.A(n10877), .B(n10854), .C(n9740), .Y(n10879));
  INVX1   g07635(.A(n10879), .Y(n10880));
  NAND2X1 g07636(.A(n9996), .B(n9771), .Y(n10882));
  XOR2X1  g07637(.A(n9810), .B(n9830), .Y(n10883));
  AOI21X1 g07638(.A0(n9810), .A1(n9829), .B0(n9827), .Y(n10884));
  OAI22X1 g07639(.A0(n10406), .A1(n10884), .B0(n10883), .B1(n10882), .Y(n10885));
  AOI21X1 g07640(.A0(n10885), .A1(n10477), .B0(n9759), .Y(n10886));
  NOR2X1  g07641(.A(n9757), .B(n9717), .Y(n10887));
  INVX1   g07642(.A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .Y(n10888));
  NOR3X1  g07643(.A(n9022), .B(n8825), .C(P2_STATE2_REG_3__SCAN_IN), .Y(n10889));
  NOR3X1  g07644(.A(n9332), .B(n9022), .C(P2_STATE2_REG_3__SCAN_IN), .Y(n10890));
  NOR4X1  g07645(.A(n9339), .B(n9470), .C(P2_STATE2_REG_3__SCAN_IN), .D(n9417), .Y(n10891));
  NOR3X1  g07646(.A(n10891), .B(n10890), .C(n10889), .Y(n10892));
  NOR3X1  g07647(.A(n9417), .B(n9339), .C(P2_STATE2_REG_3__SCAN_IN), .Y(n10893));
  NAND3X1 g07648(.A(n10893), .B(n9022), .C(n9468), .Y(n10894));
  INVX1   g07649(.A(n10894), .Y(n10895));
  NOR2X1  g07650(.A(n8884), .B(P2_STATE2_REG_3__SCAN_IN), .Y(n10896));
  AOI22X1 g07651(.A0(n10895), .A1(P2_REIP_REG_2__SCAN_IN), .B0(P2_EAX_REG_2__SCAN_IN), .B1(n10896), .Y(n10897));
  OAI21X1 g07652(.A0(n10892), .A1(n10888), .B0(n10897), .Y(n10898));
  NOR3X1  g07653(.A(n8975), .B(n9468), .C(P2_STATE2_REG_3__SCAN_IN), .Y(n10899));
  INVX1   g07654(.A(n10890), .Y(n10900));
  NAND2X1 g07655(.A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(P2_STATE2_REG_3__SCAN_IN), .Y(n10901));
  NAND2X1 g07656(.A(n10901), .B(n10900), .Y(n10902));
  AOI21X1 g07657(.A0(n10899), .A1(n9066), .B0(n10902), .Y(n10903));
  INVX1   g07658(.A(n10903), .Y(n10904));
  NAND2X1 g07659(.A(n10904), .B(n10898), .Y(n10905));
  NOR4X1  g07660(.A(n9434), .B(n9339), .C(P2_STATE2_REG_3__SCAN_IN), .D(n9417), .Y(n10906));
  NOR2X1  g07661(.A(n9208), .B(n8719), .Y(n10907));
  NOR3X1  g07662(.A(n10907), .B(n10906), .C(n10889), .Y(n10908));
  INVX1   g07663(.A(n10908), .Y(n10909));
  AOI21X1 g07664(.A0(n10899), .A1(n9094), .B0(n10909), .Y(n10910));
  NOR2X1  g07665(.A(n10892), .B(n9538), .Y(n10911));
  AOI21X1 g07666(.A0(n10896), .A1(P2_EAX_REG_0__SCAN_IN), .B0(P2_STATE2_REG_3__SCAN_IN), .Y(n10912));
  OAI21X1 g07667(.A0(n10894), .A1(n9582), .B0(n10912), .Y(n10913));
  NOR2X1  g07668(.A(n10913), .B(n10911), .Y(n10914));
  INVX1   g07669(.A(n10899), .Y(n10915));
  NOR2X1  g07670(.A(n10915), .B(n9120), .Y(n10916));
  NOR2X1  g07671(.A(n9209), .B(n8719), .Y(n10917));
  NOR4X1  g07672(.A(n10916), .B(n10896), .C(n10890), .D(n10917), .Y(n10918));
  NOR3X1  g07673(.A(n10918), .B(n10914), .C(n10910), .Y(n10919));
  NOR2X1  g07674(.A(n10918), .B(n10914), .Y(n10920));
  INVX1   g07675(.A(n10920), .Y(n10921));
  AOI22X1 g07676(.A0(n10895), .A1(P2_REIP_REG_1__SCAN_IN), .B0(P2_EAX_REG_1__SCAN_IN), .B1(n10896), .Y(n10922));
  OAI21X1 g07677(.A0(n10892), .A1(n9572), .B0(n10922), .Y(n10923));
  INVX1   g07678(.A(n10923), .Y(n10924));
  AOI21X1 g07679(.A0(n10921), .A1(n10910), .B0(n10924), .Y(n10925));
  OAI22X1 g07680(.A0(n10919), .A1(n10925), .B0(n10904), .B1(n10898), .Y(n10926));
  NAND2X1 g07681(.A(n10926), .B(n10905), .Y(n10927));
  AOI22X1 g07682(.A0(n9051), .A1(n10899), .B0(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B1(P2_STATE2_REG_3__SCAN_IN), .Y(n10928));
  INVX1   g07683(.A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .Y(n10929));
  AOI22X1 g07684(.A0(n10895), .A1(P2_REIP_REG_3__SCAN_IN), .B0(P2_EAX_REG_3__SCAN_IN), .B1(n10896), .Y(n10930));
  OAI21X1 g07685(.A0(n10892), .A1(n10929), .B0(n10930), .Y(n10931));
  XOR2X1  g07686(.A(n10931), .B(n10928), .Y(n10932));
  XOR2X1  g07687(.A(n10932), .B(n10927), .Y(n10933));
  OAI22X1 g07688(.A0(n10887), .A1(n9827), .B0(n8719), .B1(n10933), .Y(n10934));
  OAI21X1 g07689(.A0(n10934), .A1(n10886), .B0(n10880), .Y(n10935));
  OAI21X1 g07690(.A0(n10880), .A1(n9221), .B0(n10935), .Y(P2_U3602));
  XOR2X1  g07691(.A(n10883), .B(n10882), .Y(n10937));
  NOR2X1  g07692(.A(n10925), .B(n10919), .Y(n10938));
  XOR2X1  g07693(.A(n10903), .B(n10898), .Y(n10939));
  XOR2X1  g07694(.A(n10939), .B(n10938), .Y(n10940));
  INVX1   g07695(.A(n10940), .Y(n10941));
  OAI22X1 g07696(.A0(n10887), .A1(n9811), .B0(n8719), .B1(n10941), .Y(n10942));
  AOI21X1 g07697(.A0(n10937), .A1(n9758), .B0(n10942), .Y(n10943));
  NAND2X1 g07698(.A(n10879), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .Y(n10944));
  OAI21X1 g07699(.A0(n10943), .A1(n10879), .B0(n10944), .Y(P2_U3603));
  NAND2X1 g07700(.A(n9784), .B(n9772), .Y(n10946));
  NAND2X1 g07701(.A(n9784), .B(n9771), .Y(n10947));
  AOI21X1 g07702(.A0(n10947), .A1(n10946), .B0(n9759), .Y(n10948));
  INVX1   g07703(.A(n10910), .Y(n10949));
  XOR2X1  g07704(.A(n10923), .B(n10921), .Y(n10950));
  NOR3X1  g07705(.A(n10923), .B(n10920), .C(n10910), .Y(n10951));
  AOI21X1 g07706(.A0(n10923), .A1(n10919), .B0(n10951), .Y(n10952));
  OAI21X1 g07707(.A0(n10950), .A1(n10949), .B0(n10952), .Y(n10953));
  INVX1   g07708(.A(n10953), .Y(n10954));
  OAI22X1 g07709(.A0(n10887), .A1(n9784), .B0(n8719), .B1(n10954), .Y(n10955));
  OAI21X1 g07710(.A0(n10955), .A1(n10948), .B0(n10880), .Y(n10956));
  OAI21X1 g07711(.A0(n10880), .A1(n9208), .B0(n10956), .Y(P2_U3604));
  NOR2X1  g07712(.A(n9766), .B(n9717), .Y(n10958));
  XOR2X1  g07713(.A(n10918), .B(n10914), .Y(n10959));
  INVX1   g07714(.A(n10959), .Y(n10960));
  OAI22X1 g07715(.A0(n10958), .A1(n9771), .B0(n8719), .B1(n10960), .Y(n10961));
  OAI21X1 g07716(.A0(n10961), .A1(n9727), .B0(n10880), .Y(n10962));
  OAI21X1 g07717(.A0(n10880), .A1(n9209), .B0(n10962), .Y(P2_U3605));
  NOR2X1  g07718(.A(n9474), .B(n9448), .Y(n10964));
  NOR4X1  g07719(.A(P2_STATE2_REG_1__SCAN_IN), .B(P2_STATE2_REG_2__SCAN_IN), .C(P2_STATE2_REG_3__SCAN_IN), .D(P2_STATE2_REG_0__SCAN_IN), .Y(n10965));
  INVX1   g07720(.A(n10965), .Y(n10966));
  AOI21X1 g07721(.A0(n9259), .A1(n8975), .B0(n9405), .Y(n10967));
  NOR2X1  g07722(.A(n10967), .B(n9404), .Y(n10968));
  NOR3X1  g07723(.A(n9308), .B(n8946), .C(n9433), .Y(n10969));
  NAND3X1 g07724(.A(n9418), .B(n8975), .C(n8855), .Y(n10970));
  OAI21X1 g07725(.A0(n9313), .A1(n8975), .B0(n10970), .Y(n10971));
  NAND2X1 g07726(.A(n10971), .B(n9308), .Y(n10972));
  OAI21X1 g07727(.A0(n8975), .A1(n8855), .B0(n8620), .Y(n10973));
  AOI21X1 g07728(.A0(n9487), .A1(n8975), .B0(n10973), .Y(n10974));
  NAND3X1 g07729(.A(n10974), .B(n9356), .C(n9230), .Y(n10975));
  NAND4X1 g07730(.A(n10972), .B(n9436), .C(n9421), .D(n10975), .Y(n10976));
  NOR3X1  g07731(.A(n10976), .B(n10969), .C(n10968), .Y(n10977));
  OAI21X1 g07732(.A0(n10977), .A1(n9732), .B0(n10966), .Y(n10978));
  INVX1   g07733(.A(n10978), .Y(n10979));
  NOR2X1  g07734(.A(n10979), .B(n9700), .Y(n10980));
  INVX1   g07735(.A(n10980), .Y(n10981));
  AOI21X1 g07736(.A0(n9309), .A1(n8915), .B0(n9639), .Y(n10982));
  AOI21X1 g07737(.A0(n10982), .A1(n10964), .B0(n10981), .Y(n10983));
  NOR2X1  g07738(.A(n9416), .B(n9415), .Y(n10984));
  OAI21X1 g07739(.A0(n9487), .A1(n8979), .B0(n9412), .Y(n10985));
  OAI21X1 g07740(.A0(n10985), .A1(n10984), .B0(n10980), .Y(n10986));
  INVX1   g07741(.A(n9333), .Y(n10987));
  NOR3X1  g07742(.A(n10979), .B(n10987), .C(n9700), .Y(n10988));
  INVX1   g07743(.A(n10988), .Y(n10989));
  OAI22X1 g07744(.A0(n10986), .A1(n10960), .B0(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(n10989), .Y(n10990));
  AOI21X1 g07745(.A0(n10983), .A1(n9538), .B0(n10990), .Y(n10991));
  AOI22X1 g07746(.A0(n8980), .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B0(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(n8981), .Y(n10992));
  AOI22X1 g07747(.A0(n8983), .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B0(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(n8984), .Y(n10993));
  AOI22X1 g07748(.A0(n8986), .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B0(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(n8987), .Y(n10994));
  AOI22X1 g07749(.A0(n8989), .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B0(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(n8990), .Y(n10995));
  NAND4X1 g07750(.A(n10994), .B(n10993), .C(n10992), .D(n10995), .Y(n10996));
  AOI22X1 g07751(.A0(n8993), .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B0(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(n8994), .Y(n10997));
  AOI22X1 g07752(.A0(n8996), .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B0(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(n8997), .Y(n10998));
  AOI22X1 g07753(.A0(n8999), .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B0(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(n9000), .Y(n10999));
  AOI22X1 g07754(.A0(n9002), .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B0(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(n9003), .Y(n11000));
  NAND4X1 g07755(.A(n10999), .B(n10998), .C(n10997), .D(n11000), .Y(n11001));
  NOR2X1  g07756(.A(n11001), .B(n10996), .Y(n11002));
  NOR2X1  g07757(.A(n8825), .B(n9532), .Y(n11003));
  AOI21X1 g07758(.A0(n9153), .A1(n8825), .B0(n11003), .Y(n11004));
  XOR2X1  g07759(.A(n11004), .B(n8825), .Y(n11005));
  NOR2X1  g07760(.A(n11005), .B(n11002), .Y(n11006));
  INVX1   g07761(.A(n11002), .Y(n11007));
  NAND3X1 g07762(.A(n10166), .B(n9815), .C(n9794), .Y(n11008));
  NAND3X1 g07763(.A(n10224), .B(n9815), .C(n9794), .Y(n11009));
  OAI22X1 g07764(.A0(n11008), .A1(n8931), .B0(n8916), .B1(n11009), .Y(n11010));
  NAND3X1 g07765(.A(n10284), .B(n9815), .C(n9794), .Y(n11011));
  NAND3X1 g07766(.A(n10342), .B(n9815), .C(n9794), .Y(n11012));
  OAI22X1 g07767(.A0(n11011), .A1(n8923), .B0(n8941), .B1(n11012), .Y(n11013));
  NOR2X1  g07768(.A(n11013), .B(n11010), .Y(n11014));
  OAI22X1 g07769(.A0(n10167), .A1(n8919), .B0(n8926), .B1(n10225), .Y(n11015));
  OAI22X1 g07770(.A0(n10285), .A1(n8934), .B0(n8938), .B1(n10343), .Y(n11016));
  NOR2X1  g07771(.A(n11016), .B(n11015), .Y(n11017));
  NAND3X1 g07772(.A(n10166), .B(n9663), .C(n9633), .Y(n11018));
  NAND4X1 g07773(.A(n9663), .B(n9633), .C(P2_INSTQUEUE_REG_2__0__SCAN_IN), .D(n10224), .Y(n11019));
  OAI21X1 g07774(.A0(n11018), .A1(n9102), .B0(n11019), .Y(n11020));
  NAND3X1 g07775(.A(n10342), .B(n9663), .C(n9633), .Y(n11021));
  NAND4X1 g07776(.A(n9663), .B(n9633), .C(P2_INSTQUEUE_REG_1__0__SCAN_IN), .D(n10284), .Y(n11022));
  OAI21X1 g07777(.A0(n11021), .A1(n9099), .B0(n11022), .Y(n11023));
  AOI22X1 g07778(.A0(n10403), .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B0(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(n10459), .Y(n11024));
  AOI22X1 g07779(.A0(n10517), .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B0(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(n10573), .Y(n11025));
  NAND2X1 g07780(.A(n11025), .B(n11024), .Y(n11026));
  NOR3X1  g07781(.A(n11026), .B(n11023), .C(n11020), .Y(n11027));
  NAND3X1 g07782(.A(n11027), .B(n11017), .C(n11014), .Y(n11028));
  NOR2X1  g07783(.A(n9120), .B(n8975), .Y(n11029));
  AOI21X1 g07784(.A0(n11028), .A1(n8975), .B0(n11029), .Y(n11030));
  XOR2X1  g07785(.A(n11030), .B(n9022), .Y(n11031));
  NOR2X1  g07786(.A(n11031), .B(n11007), .Y(n11032));
  NOR2X1  g07787(.A(n11032), .B(n11006), .Y(n11033));
  XOR2X1  g07788(.A(n11033), .B(n9538), .Y(n11034));
  NOR4X1  g07789(.A(n8979), .B(n9404), .C(n9700), .D(n10979), .Y(n11035));
  NAND2X1 g07790(.A(n11035), .B(n11034), .Y(n11036));
  XOR2X1  g07791(.A(n11031), .B(n9538), .Y(n11037));
  NOR3X1  g07792(.A(n9487), .B(n8975), .C(n8946), .Y(n11039));
  NOR4X1  g07793(.A(n9640), .B(n9598), .C(n9675), .D(n11039), .Y(n11040));
  NOR3X1  g07794(.A(n11040), .B(n10979), .C(n9700), .Y(n11041));
  INVX1   g07795(.A(n11041), .Y(n11042));
  AOI22X1 g07796(.A0(n10979), .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B0(P2_REIP_REG_0__SCAN_IN), .B1(n10965), .Y(n11044));
  OAI21X1 g07797(.A0(n11042), .A1(n9614), .B0(n11044), .Y(n11045));
  AOI21X1 g07798(.A0(n12547), .A1(n11037), .B0(n11045), .Y(n11046));
  NAND3X1 g07799(.A(n11046), .B(n11036), .C(n10991), .Y(P2_U3046));
  XOR2X1  g07800(.A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n9538), .Y(n11048));
  INVX1   g07801(.A(n11048), .Y(n11049));
  OAI22X1 g07802(.A0(n10989), .A1(n11048), .B0(n10986), .B1(n10954), .Y(n11050));
  AOI21X1 g07803(.A0(n11049), .A1(n10983), .B0(n11050), .Y(n11051));
  OAI21X1 g07804(.A0(n11032), .A1(n11006), .B0(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .Y(n11052));
  NOR2X1  g07805(.A(n8825), .B(n9484), .Y(n11054));
  AOI21X1 g07806(.A0(n9269), .A1(n8825), .B0(n11054), .Y(n11055));
  XOR2X1  g07807(.A(n11055), .B(n11003), .Y(n11056));
  NOR2X1  g07808(.A(n11056), .B(n11002), .Y(n11057));
  AOI22X1 g07809(.A0(n9754), .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B0(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(n9993), .Y(n11058));
  AOI22X1 g07810(.A0(n10053), .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B0(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(n10110), .Y(n11059));
  NAND2X1 g07811(.A(n11059), .B(n11058), .Y(n11060));
  OAI22X1 g07812(.A0(n10167), .A1(n8950), .B0(n8957), .B1(n10225), .Y(n11061));
  OAI22X1 g07813(.A0(n10285), .A1(n8964), .B0(n8968), .B1(n10343), .Y(n11062));
  AOI22X1 g07814(.A0(n10629), .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B0(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(n10685), .Y(n11063));
  AOI22X1 g07815(.A0(n10743), .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B0(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(n10799), .Y(n11064));
  AOI22X1 g07816(.A0(n10403), .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B0(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(n10459), .Y(n11065));
  AOI22X1 g07817(.A0(n10517), .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B0(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(n10573), .Y(n11066));
  NAND4X1 g07818(.A(n11065), .B(n11064), .C(n11063), .D(n11066), .Y(n11067));
  NOR4X1  g07819(.A(n11062), .B(n11061), .C(n11060), .D(n11067), .Y(n11068));
  NAND2X1 g07820(.A(n9094), .B(n9022), .Y(n11069));
  OAI21X1 g07821(.A0(n11068), .A1(n9022), .B0(n11069), .Y(n11070));
  NOR2X1  g07822(.A(n9119), .B(n8975), .Y(n11071));
  NAND3X1 g07823(.A(n11070), .B(n11030), .C(n9022), .Y(n11072));
  OAI21X1 g07824(.A0(n11071), .A1(n11070), .B0(n11072), .Y(n11073));
  AOI21X1 g07825(.A0(n11073), .A1(n11002), .B0(n11057), .Y(n11074));
  NOR3X1  g07826(.A(n11074), .B(n11052), .C(n9572), .Y(n11075));
  INVX1   g07827(.A(n11074), .Y(n11076));
  XOR2X1  g07828(.A(n11052), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .Y(n11077));
  NAND3X1 g07829(.A(n11076), .B(n11052), .C(n9572), .Y(n11078));
  OAI21X1 g07830(.A0(n11077), .A1(n11076), .B0(n11078), .Y(n11079));
  OAI21X1 g07831(.A0(n11079), .A1(n11075), .B0(n11035), .Y(n11080));
  NOR2X1  g07832(.A(n11031), .B(n9538), .Y(n11081));
  NAND3X1 g07833(.A(n11081), .B(n11073), .C(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .Y(n11082));
  INVX1   g07834(.A(n11073), .Y(n11083));
  XOR2X1  g07835(.A(n11081), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .Y(n11084));
  NAND2X1 g07836(.A(n11084), .B(n11083), .Y(n11085));
  INVX1   g07837(.A(n11081), .Y(n11086));
  NAND3X1 g07838(.A(n11086), .B(n11073), .C(n9572), .Y(n11087));
  NAND3X1 g07839(.A(n11087), .B(n11085), .C(n11082), .Y(n11088));
  AOI22X1 g07840(.A0(n10979), .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B0(P2_REIP_REG_1__SCAN_IN), .B1(n10965), .Y(n11089));
  OAI21X1 g07841(.A0(n11042), .A1(n9595), .B0(n11089), .Y(n11090));
  AOI21X1 g07842(.A0(n11088), .A1(n12547), .B0(n11090), .Y(n11091));
  NAND3X1 g07843(.A(n11091), .B(n11080), .C(n11051), .Y(P2_U3045));
  NAND2X1 g07844(.A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .Y(n11093));
  XOR2X1  g07845(.A(n11093), .B(n10888), .Y(n11094));
  NAND2X1 g07846(.A(n11094), .B(n10983), .Y(n11095));
  INVX1   g07847(.A(n10986), .Y(n11096));
  XOR2X1  g07848(.A(n11093), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .Y(n11097));
  AOI22X1 g07849(.A0(n10988), .A1(n11097), .B0(n11096), .B1(n10940), .Y(n11098));
  NOR2X1  g07850(.A(n11074), .B(n11052), .Y(n11099));
  AOI21X1 g07851(.A0(n11074), .A1(n11052), .B0(n9572), .Y(n11100));
  NOR2X1  g07852(.A(n11100), .B(n11099), .Y(n11101));
  OAI21X1 g07853(.A0(n11004), .A1(n8825), .B0(n11055), .Y(n11102));
  INVX1   g07854(.A(n11102), .Y(n11103));
  NOR2X1  g07855(.A(n9148), .B(n9468), .Y(n11104));
  AOI21X1 g07856(.A0(n9468), .A1(P2_EBX_REG_2__SCAN_IN), .B0(n11104), .Y(n11105));
  XOR2X1  g07857(.A(n11105), .B(n11103), .Y(n11106));
  NAND2X1 g07858(.A(n11106), .B(n11007), .Y(n11107));
  NOR2X1  g07859(.A(n11068), .B(n9022), .Y(n11108));
  AOI21X1 g07860(.A0(n9094), .A1(n9022), .B0(n11108), .Y(n11109));
  AOI21X1 g07861(.A0(n11030), .A1(n9022), .B0(n11109), .Y(n11110));
  AOI22X1 g07862(.A0(n9754), .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B0(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(n9993), .Y(n11111));
  AOI22X1 g07863(.A0(n10053), .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B0(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(n10110), .Y(n11112));
  NAND2X1 g07864(.A(n11112), .B(n11111), .Y(n11113));
  OAI22X1 g07865(.A0(n10167), .A1(n8830), .B0(n8837), .B1(n10225), .Y(n11114));
  OAI22X1 g07866(.A0(n10285), .A1(n8844), .B0(n8848), .B1(n10343), .Y(n11115));
  AOI22X1 g07867(.A0(n10629), .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B0(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(n10685), .Y(n11116));
  AOI22X1 g07868(.A0(n10743), .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B0(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(n10799), .Y(n11117));
  AOI22X1 g07869(.A0(n10403), .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B0(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(n10459), .Y(n11118));
  AOI22X1 g07870(.A0(n10517), .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B0(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(n10573), .Y(n11119));
  NAND4X1 g07871(.A(n11118), .B(n11117), .C(n11116), .D(n11119), .Y(n11120));
  NOR4X1  g07872(.A(n11115), .B(n11114), .C(n11113), .D(n11120), .Y(n11121));
  OAI21X1 g07873(.A0(n9064), .A1(n9059), .B0(n9022), .Y(n11122));
  OAI21X1 g07874(.A0(n11121), .A1(n9022), .B0(n11122), .Y(n11123));
  XOR2X1  g07875(.A(n11123), .B(n8975), .Y(n11124));
  XOR2X1  g07876(.A(n11124), .B(n11110), .Y(n11125));
  OAI21X1 g07877(.A0(n11125), .A1(n11007), .B0(n11107), .Y(n11126));
  XOR2X1  g07878(.A(n11126), .B(n10888), .Y(n11127));
  XOR2X1  g07879(.A(n11127), .B(n11101), .Y(n11128));
  NAND2X1 g07880(.A(n11128), .B(n11035), .Y(n11129));
  OAI21X1 g07881(.A0(n11081), .A1(n11073), .B0(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .Y(n11130));
  OAI21X1 g07882(.A0(n11086), .A1(n11083), .B0(n11130), .Y(n11131));
  XOR2X1  g07883(.A(n11125), .B(n10888), .Y(n11132));
  XOR2X1  g07884(.A(n11132), .B(n11131), .Y(n11133));
  AOI22X1 g07885(.A0(n10979), .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B0(P2_REIP_REG_2__SCAN_IN), .B1(n10965), .Y(n11134));
  OAI21X1 g07886(.A0(n11042), .A1(n9633), .B0(n11134), .Y(n11135));
  AOI21X1 g07887(.A0(n11133), .A1(n12547), .B0(n11135), .Y(n11136));
  NAND4X1 g07888(.A(n11129), .B(n11098), .C(n11095), .D(n11136), .Y(P2_U3044));
  NAND3X1 g07889(.A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .Y(n11138));
  XOR2X1  g07890(.A(n11138), .B(n10929), .Y(n11139));
  NAND2X1 g07891(.A(n11139), .B(n10983), .Y(n11140));
  INVX1   g07892(.A(n10933), .Y(n11141));
  AOI21X1 g07893(.A0(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B0(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .Y(n11142));
  XOR2X1  g07894(.A(n11142), .B(n10929), .Y(n11143));
  AOI22X1 g07895(.A0(n10988), .A1(n11143), .B0(n11096), .B1(n11141), .Y(n11144));
  NAND2X1 g07896(.A(n11126), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .Y(n11145));
  OAI22X1 g07897(.A0(n11100), .A1(n11099), .B0(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B1(n11126), .Y(n11146));
  NAND2X1 g07898(.A(n11146), .B(n11145), .Y(n11147));
  NAND2X1 g07899(.A(n11105), .B(n11103), .Y(n11148));
  NOR2X1  g07900(.A(n8825), .B(n9658), .Y(n11149));
  AOI21X1 g07901(.A0(n9146), .A1(n8825), .B0(n11149), .Y(n11150));
  XOR2X1  g07902(.A(n11150), .B(n11148), .Y(n11151));
  NOR2X1  g07903(.A(n11151), .B(n11002), .Y(n11152));
  INVX1   g07904(.A(n11152), .Y(n11153));
  NOR2X1  g07905(.A(n9065), .B(n8975), .Y(n11154));
  NAND3X1 g07906(.A(n11122), .B(n11121), .C(n8975), .Y(n11155));
  AOI21X1 g07907(.A0(n11155), .A1(n11110), .B0(n11154), .Y(n11156));
  OAI22X1 g07908(.A0(n11008), .A1(n8899), .B0(n8885), .B1(n11009), .Y(n11157));
  OAI22X1 g07909(.A0(n11011), .A1(n8892), .B0(n8909), .B1(n11012), .Y(n11158));
  OAI22X1 g07910(.A0(n10167), .A1(n8888), .B0(n8895), .B1(n10225), .Y(n11159));
  OAI22X1 g07911(.A0(n10285), .A1(n8902), .B0(n8906), .B1(n10343), .Y(n11160));
  NOR4X1  g07912(.A(n11159), .B(n11158), .C(n11157), .D(n11160), .Y(n11161));
  INVX1   g07913(.A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .Y(n11162));
  NAND4X1 g07914(.A(n9663), .B(n9633), .C(P2_INSTQUEUE_REG_2__3__SCAN_IN), .D(n10224), .Y(n11163));
  OAI21X1 g07915(.A0(n11018), .A1(n11162), .B0(n11163), .Y(n11164));
  NAND4X1 g07916(.A(n9663), .B(n9633), .C(P2_INSTQUEUE_REG_1__3__SCAN_IN), .D(n10284), .Y(n11165));
  OAI21X1 g07917(.A0(n11021), .A1(n9824), .B0(n11165), .Y(n11166));
  NOR2X1  g07918(.A(n11166), .B(n11164), .Y(n11167));
  AOI22X1 g07919(.A0(n10403), .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B0(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(n10459), .Y(n11168));
  AOI22X1 g07920(.A0(n10517), .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B0(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(n10573), .Y(n11169));
  NAND4X1 g07921(.A(n11168), .B(n11167), .C(n11161), .D(n11169), .Y(n11170));
  NAND2X1 g07922(.A(n11170), .B(n8975), .Y(n11171));
  OAI21X1 g07923(.A0(n9045), .A1(n9040), .B0(n9022), .Y(n11172));
  NAND2X1 g07924(.A(n11172), .B(n11171), .Y(n11173));
  XOR2X1  g07925(.A(n11173), .B(n11156), .Y(n11174));
  OAI21X1 g07926(.A0(n11174), .A1(n11007), .B0(n11153), .Y(n11175));
  XOR2X1  g07927(.A(n11175), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .Y(n11176));
  XOR2X1  g07928(.A(n11176), .B(n11147), .Y(n11177));
  NAND2X1 g07929(.A(n11177), .B(n11035), .Y(n11178));
  NOR2X1  g07930(.A(n11125), .B(n10888), .Y(n11179));
  NAND2X1 g07931(.A(n11125), .B(n10888), .Y(n11180));
  AOI21X1 g07932(.A0(n11180), .A1(n11131), .B0(n11179), .Y(n11181));
  XOR2X1  g07933(.A(n11174), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .Y(n11182));
  XOR2X1  g07934(.A(n11182), .B(n11181), .Y(n11183));
  AOI22X1 g07935(.A0(n10979), .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B0(P2_REIP_REG_3__SCAN_IN), .B1(n10965), .Y(n11184));
  OAI21X1 g07936(.A0(n11042), .A1(n9663), .B0(n11184), .Y(n11185));
  AOI21X1 g07937(.A0(n11183), .A1(n12547), .B0(n11185), .Y(n11186));
  NAND4X1 g07938(.A(n11178), .B(n11144), .C(n11140), .D(n11186), .Y(P2_U3043));
  INVX1   g07939(.A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .Y(n11188));
  NAND4X1 g07940(.A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .D(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .Y(n11189));
  XOR2X1  g07941(.A(n11189), .B(n11188), .Y(n11190));
  NAND2X1 g07942(.A(n11190), .B(n10983), .Y(n11191));
  INVX1   g07943(.A(n10931), .Y(n11192));
  NOR2X1  g07944(.A(n11192), .B(n10928), .Y(n11193));
  AOI22X1 g07945(.A0(n10928), .A1(n11192), .B0(n10926), .B1(n10905), .Y(n11194));
  NOR2X1  g07946(.A(n11194), .B(n11193), .Y(n11195));
  NOR4X1  g07947(.A(n8975), .B(n9468), .C(P2_STATE2_REG_3__SCAN_IN), .D(n9034), .Y(n11196));
  INVX1   g07948(.A(n11196), .Y(n11197));
  AOI22X1 g07949(.A0(n10895), .A1(P2_REIP_REG_4__SCAN_IN), .B0(P2_EAX_REG_4__SCAN_IN), .B1(n10896), .Y(n11198));
  OAI21X1 g07950(.A0(n10892), .A1(n11188), .B0(n11198), .Y(n11199));
  XOR2X1  g07951(.A(n11199), .B(n11197), .Y(n11200));
  XOR2X1  g07952(.A(n11200), .B(n11195), .Y(n11201));
  NOR2X1  g07953(.A(n11142), .B(n10929), .Y(n11202));
  XOR2X1  g07954(.A(n11202), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .Y(n11203));
  AOI22X1 g07955(.A0(n11201), .A1(n11096), .B0(n10988), .B1(n11203), .Y(n11204));
  NOR2X1  g07956(.A(n11175), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .Y(n11205));
  NOR2X1  g07957(.A(n11205), .B(n11146), .Y(n11206));
  NOR2X1  g07958(.A(n9046), .B(n8975), .Y(n11207));
  AOI21X1 g07959(.A0(n11170), .A1(n8975), .B0(n11207), .Y(n11208));
  XOR2X1  g07960(.A(n11208), .B(n11156), .Y(n11209));
  AOI21X1 g07961(.A0(n11209), .A1(n11002), .B0(n11152), .Y(n11210));
  AOI21X1 g07962(.A0(n11210), .A1(n10929), .B0(n11145), .Y(n11211));
  NOR2X1  g07963(.A(n11210), .B(n10929), .Y(n11212));
  NOR3X1  g07964(.A(n11212), .B(n11211), .C(n11206), .Y(n11213));
  NAND3X1 g07965(.A(n11150), .B(n11105), .C(n11103), .Y(n11214));
  INVX1   g07966(.A(P2_EBX_REG_4__SCAN_IN), .Y(n11215));
  NOR2X1  g07967(.A(n8825), .B(n11215), .Y(n11216));
  AOI21X1 g07968(.A0(n9159), .A1(n8825), .B0(n11216), .Y(n11217));
  XOR2X1  g07969(.A(n11217), .B(n11214), .Y(n11218));
  NOR2X1  g07970(.A(n11218), .B(n11002), .Y(n11219));
  AOI21X1 g07971(.A0(n11172), .A1(n11171), .B0(n11156), .Y(n11220));
  AOI22X1 g07972(.A0(n9754), .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B0(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(n9993), .Y(n11221));
  AOI22X1 g07973(.A0(n10053), .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B0(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(n10110), .Y(n11222));
  AOI22X1 g07974(.A0(n10168), .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B0(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(n10226), .Y(n11223));
  AOI22X1 g07975(.A0(n10286), .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B0(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(n10344), .Y(n11224));
  NAND4X1 g07976(.A(n11223), .B(n11222), .C(n11221), .D(n11224), .Y(n11225));
  AOI22X1 g07977(.A0(n10629), .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B0(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(n10685), .Y(n11226));
  AOI22X1 g07978(.A0(n10743), .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B0(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(n10799), .Y(n11227));
  AOI22X1 g07979(.A0(n10403), .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B0(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(n10459), .Y(n11228));
  AOI22X1 g07980(.A0(n10517), .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B0(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(n10573), .Y(n11229));
  NAND4X1 g07981(.A(n11228), .B(n11227), .C(n11226), .D(n11229), .Y(n11230));
  OAI21X1 g07982(.A0(n11230), .A1(n11225), .B0(n8975), .Y(n11231));
  OAI21X1 g07983(.A0(n9034), .A1(n8975), .B0(n11231), .Y(n11232));
  XOR2X1  g07984(.A(n11232), .B(n11220), .Y(n11233));
  AOI21X1 g07985(.A0(n11233), .A1(n11002), .B0(n11219), .Y(n11234));
  XOR2X1  g07986(.A(n11234), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .Y(n11235));
  XOR2X1  g07987(.A(n11235), .B(n11213), .Y(n11236));
  NAND2X1 g07988(.A(n11236), .B(n11035), .Y(n11237));
  AOI21X1 g07989(.A0(n11174), .A1(n10929), .B0(n11181), .Y(n11238));
  AOI21X1 g07990(.A0(n11209), .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B0(n11238), .Y(n11239));
  XOR2X1  g07991(.A(n11233), .B(n11188), .Y(n11240));
  INVX1   g07992(.A(n11240), .Y(n11241));
  XOR2X1  g07993(.A(n11241), .B(n11239), .Y(n11242));
  NOR4X1  g07994(.A(n10981), .B(n8977), .C(n9404), .D(n11242), .Y(n11243));
  NOR2X1  g07995(.A(n9661), .B(n9656), .Y(n11244));
  NAND2X1 g07996(.A(n9661), .B(n9656), .Y(n11245));
  AOI21X1 g07997(.A0(n11245), .A1(n9655), .B0(n11244), .Y(n11246));
  AOI22X1 g07998(.A0(P2_REIP_REG_4__SCAN_IN), .A1(n9488), .B0(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(P2_STATE2_REG_1__SCAN_IN), .Y(n11247));
  OAI21X1 g07999(.A0(n9485), .A1(n11215), .B0(n11247), .Y(n11248));
  AOI21X1 g08000(.A0(n9483), .A1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B0(n11248), .Y(n11249));
  INVX1   g08001(.A(n11249), .Y(n11250));
  XOR2X1  g08002(.A(n11250), .B(n11246), .Y(n11251));
  AOI22X1 g08003(.A0(n10979), .A1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B0(P2_REIP_REG_4__SCAN_IN), .B1(n10965), .Y(n11252));
  OAI21X1 g08004(.A0(n11251), .A1(n11042), .B0(n11252), .Y(n11253));
  NOR2X1  g08005(.A(n11253), .B(n11243), .Y(n11254));
  NAND4X1 g08006(.A(n11237), .B(n11204), .C(n11191), .D(n11254), .Y(P2_U3042));
  NOR2X1  g08007(.A(n11189), .B(n11188), .Y(n11256));
  XOR2X1  g08008(.A(n11256), .B(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .Y(n11257));
  NAND2X1 g08009(.A(n11257), .B(n10983), .Y(n11258));
  INVX1   g08010(.A(n11199), .Y(n11259));
  OAI22X1 g08011(.A0(n11196), .A1(n11199), .B0(n11194), .B1(n11193), .Y(n11260));
  OAI21X1 g08012(.A0(n11259), .A1(n11197), .B0(n11260), .Y(n11261));
  NOR4X1  g08013(.A(n8975), .B(n9468), .C(P2_STATE2_REG_3__SCAN_IN), .D(n9018), .Y(n11262));
  INVX1   g08014(.A(n11262), .Y(n11263));
  INVX1   g08015(.A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .Y(n11264));
  AOI22X1 g08016(.A0(n10895), .A1(P2_REIP_REG_5__SCAN_IN), .B0(P2_EAX_REG_5__SCAN_IN), .B1(n10896), .Y(n11265));
  OAI21X1 g08017(.A0(n10892), .A1(n11264), .B0(n11265), .Y(n11266));
  XOR2X1  g08018(.A(n11266), .B(n11263), .Y(n11267));
  XOR2X1  g08019(.A(n11267), .B(n11261), .Y(n11268));
  INVX1   g08020(.A(n11268), .Y(n11269));
  NOR3X1  g08021(.A(n11142), .B(n11188), .C(n10929), .Y(n11270));
  XOR2X1  g08022(.A(n11270), .B(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .Y(n11271));
  AOI22X1 g08023(.A0(n11269), .A1(n11096), .B0(n10988), .B1(n11271), .Y(n11272));
  NOR2X1  g08024(.A(n11234), .B(n11188), .Y(n11273));
  AOI21X1 g08025(.A0(n11234), .A1(n11188), .B0(n11213), .Y(n11274));
  NOR2X1  g08026(.A(n11274), .B(n11273), .Y(n11275));
  NAND4X1 g08027(.A(n11150), .B(n11105), .C(n11103), .D(n11217), .Y(n11276));
  INVX1   g08028(.A(n11276), .Y(n11277));
  INVX1   g08029(.A(P2_EBX_REG_5__SCAN_IN), .Y(n11278));
  NOR2X1  g08030(.A(n8825), .B(n11278), .Y(n11279));
  AOI21X1 g08031(.A0(n9141), .A1(n8825), .B0(n11279), .Y(n11280));
  XOR2X1  g08032(.A(n11280), .B(n11277), .Y(n11281));
  INVX1   g08033(.A(n11281), .Y(n11282));
  NOR2X1  g08034(.A(n11282), .B(n11002), .Y(n11283));
  NAND2X1 g08035(.A(n11232), .B(n11220), .Y(n11284));
  AOI22X1 g08036(.A0(n9754), .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B0(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(n9993), .Y(n11285));
  AOI22X1 g08037(.A0(n10053), .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B0(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(n10110), .Y(n11286));
  AOI22X1 g08038(.A0(n10168), .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B0(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(n10226), .Y(n11287));
  AOI22X1 g08039(.A0(n10286), .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B0(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(n10344), .Y(n11288));
  NAND4X1 g08040(.A(n11287), .B(n11286), .C(n11285), .D(n11288), .Y(n11289));
  AOI22X1 g08041(.A0(n10629), .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B0(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(n10685), .Y(n11290));
  AOI22X1 g08042(.A0(n10743), .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B0(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(n10799), .Y(n11291));
  AOI22X1 g08043(.A0(n10403), .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B0(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(n10459), .Y(n11292));
  AOI22X1 g08044(.A0(n10517), .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B0(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(n10573), .Y(n11293));
  NAND4X1 g08045(.A(n11292), .B(n11291), .C(n11290), .D(n11293), .Y(n11294));
  NOR2X1  g08046(.A(n11294), .B(n11289), .Y(n11295));
  NOR2X1  g08047(.A(n9018), .B(n8975), .Y(n11296));
  INVX1   g08048(.A(n11296), .Y(n11297));
  OAI21X1 g08049(.A0(n11295), .A1(n9022), .B0(n11297), .Y(n11298));
  INVX1   g08050(.A(n11298), .Y(n11299));
  XOR2X1  g08051(.A(n11299), .B(n11284), .Y(n11300));
  AOI21X1 g08052(.A0(n11300), .A1(n11002), .B0(n11283), .Y(n11301));
  XOR2X1  g08053(.A(n11301), .B(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .Y(n11302));
  XOR2X1  g08054(.A(n11302), .B(n11275), .Y(n11303));
  NAND2X1 g08055(.A(n11303), .B(n11035), .Y(n11304));
  NOR2X1  g08056(.A(n11233), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .Y(n11305));
  NOR2X1  g08057(.A(n11305), .B(n11239), .Y(n11306));
  AOI21X1 g08058(.A0(n11233), .A1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B0(n11306), .Y(n11307));
  XOR2X1  g08059(.A(n11298), .B(n11284), .Y(n11308));
  XOR2X1  g08060(.A(n11308), .B(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .Y(n11309));
  XOR2X1  g08061(.A(n11309), .B(n11307), .Y(n11310));
  NOR2X1  g08062(.A(n11249), .B(n11246), .Y(n11311));
  AOI22X1 g08063(.A0(P2_REIP_REG_5__SCAN_IN), .A1(n9488), .B0(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(P2_STATE2_REG_1__SCAN_IN), .Y(n11312));
  OAI21X1 g08064(.A0(n9485), .A1(n11278), .B0(n11312), .Y(n11313));
  AOI21X1 g08065(.A0(n9483), .A1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B0(n11313), .Y(n11314));
  XOR2X1  g08066(.A(n11314), .B(n11311), .Y(n11315));
  AOI22X1 g08067(.A0(n10979), .A1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B0(P2_REIP_REG_5__SCAN_IN), .B1(n10965), .Y(n11316));
  OAI21X1 g08068(.A0(n11315), .A1(n11042), .B0(n11316), .Y(n11317));
  AOI21X1 g08069(.A0(n11310), .A1(n12547), .B0(n11317), .Y(n11318));
  NAND4X1 g08070(.A(n11304), .B(n11272), .C(n11258), .D(n11318), .Y(P2_U3041));
  NOR3X1  g08071(.A(n11189), .B(n11264), .C(n11188), .Y(n11320));
  XOR2X1  g08072(.A(n11320), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .Y(n11321));
  NAND2X1 g08073(.A(n11321), .B(n10983), .Y(n11322));
  INVX1   g08074(.A(n11266), .Y(n11323));
  NOR2X1  g08075(.A(n11323), .B(n11263), .Y(n11324));
  NOR2X1  g08076(.A(n11266), .B(n11262), .Y(n11325));
  INVX1   g08077(.A(n11325), .Y(n11326));
  AOI21X1 g08078(.A0(n11326), .A1(n11261), .B0(n11324), .Y(n11327));
  NOR2X1  g08079(.A(n9005), .B(n8992), .Y(n11328));
  NOR4X1  g08080(.A(n8975), .B(n9468), .C(P2_STATE2_REG_3__SCAN_IN), .D(n11328), .Y(n11329));
  INVX1   g08081(.A(n11329), .Y(n11330));
  INVX1   g08082(.A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .Y(n11331));
  AOI22X1 g08083(.A0(n10895), .A1(P2_REIP_REG_6__SCAN_IN), .B0(P2_EAX_REG_6__SCAN_IN), .B1(n10896), .Y(n11332));
  OAI21X1 g08084(.A0(n10892), .A1(n11331), .B0(n11332), .Y(n11333));
  XOR2X1  g08085(.A(n11333), .B(n11330), .Y(n11334));
  XOR2X1  g08086(.A(n11334), .B(n11327), .Y(n11335));
  NOR4X1  g08087(.A(n11264), .B(n11188), .C(n10929), .D(n11142), .Y(n11336));
  XOR2X1  g08088(.A(n11336), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .Y(n11337));
  AOI22X1 g08089(.A0(n11335), .A1(n11096), .B0(n10988), .B1(n11337), .Y(n11338));
  NAND2X1 g08090(.A(n11234), .B(n11188), .Y(n11339));
  INVX1   g08091(.A(n11283), .Y(n11340));
  OAI21X1 g08092(.A0(n11308), .A1(n11007), .B0(n11340), .Y(n11341));
  OAI21X1 g08093(.A0(n11341), .A1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B0(n11339), .Y(n11342));
  NOR2X1  g08094(.A(n11342), .B(n11213), .Y(n11343));
  OAI21X1 g08095(.A0(n11341), .A1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B0(n11273), .Y(n11344));
  OAI21X1 g08096(.A0(n11301), .A1(n11264), .B0(n11344), .Y(n11345));
  NOR2X1  g08097(.A(n11345), .B(n11343), .Y(n11346));
  INVX1   g08098(.A(n11346), .Y(n11347));
  NAND2X1 g08099(.A(n11280), .B(n11277), .Y(n11348));
  INVX1   g08100(.A(P2_EBX_REG_6__SCAN_IN), .Y(n11349));
  NAND2X1 g08101(.A(n9138), .B(n8825), .Y(n11350));
  OAI21X1 g08102(.A0(n8825), .A1(n11349), .B0(n11350), .Y(n11351));
  XOR2X1  g08103(.A(n11351), .B(n11348), .Y(n11352));
  NAND2X1 g08104(.A(n11352), .B(n11007), .Y(n11353));
  NAND3X1 g08105(.A(n11298), .B(n11232), .C(n11220), .Y(n11354));
  AOI22X1 g08106(.A0(n9754), .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B0(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(n9993), .Y(n11355));
  AOI22X1 g08107(.A0(n10053), .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B0(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(n10110), .Y(n11356));
  AOI22X1 g08108(.A0(n10168), .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B0(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(n10226), .Y(n11357));
  AOI22X1 g08109(.A0(n10286), .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B0(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(n10344), .Y(n11358));
  NAND4X1 g08110(.A(n11357), .B(n11356), .C(n11355), .D(n11358), .Y(n11359));
  AOI22X1 g08111(.A0(n10629), .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B0(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(n10685), .Y(n11360));
  AOI22X1 g08112(.A0(n10743), .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B0(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(n10799), .Y(n11361));
  AOI22X1 g08113(.A0(n10403), .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B0(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(n10459), .Y(n11362));
  AOI22X1 g08114(.A0(n10517), .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B0(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(n10573), .Y(n11363));
  NAND4X1 g08115(.A(n11362), .B(n11361), .C(n11360), .D(n11363), .Y(n11364));
  OAI21X1 g08116(.A0(n11364), .A1(n11359), .B0(n8975), .Y(n11365));
  OAI21X1 g08117(.A0(n11328), .A1(n8975), .B0(n11365), .Y(n11366));
  XOR2X1  g08118(.A(n11366), .B(n11354), .Y(n11367));
  OAI21X1 g08119(.A0(n11367), .A1(n11007), .B0(n11353), .Y(n11368));
  XOR2X1  g08120(.A(n11368), .B(n11331), .Y(n11369));
  XOR2X1  g08121(.A(n11369), .B(n11347), .Y(n11370));
  INVX1   g08122(.A(n11370), .Y(n11371));
  NAND2X1 g08123(.A(n11371), .B(n11035), .Y(n11372));
  AOI21X1 g08124(.A0(n11308), .A1(n11264), .B0(n11307), .Y(n11373));
  AOI21X1 g08125(.A0(n11300), .A1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B0(n11373), .Y(n11374));
  XOR2X1  g08126(.A(n11367), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .Y(n11375));
  XOR2X1  g08127(.A(n11375), .B(n11374), .Y(n11376));
  NOR3X1  g08128(.A(n11314), .B(n11249), .C(n11246), .Y(n11377));
  AOI22X1 g08129(.A0(P2_REIP_REG_6__SCAN_IN), .A1(n9488), .B0(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(P2_STATE2_REG_1__SCAN_IN), .Y(n11378));
  OAI21X1 g08130(.A0(n9485), .A1(n11349), .B0(n11378), .Y(n11379));
  AOI21X1 g08131(.A0(n9483), .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B0(n11379), .Y(n11380));
  XOR2X1  g08132(.A(n11380), .B(n11377), .Y(n11381));
  AOI22X1 g08133(.A0(n10979), .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B0(P2_REIP_REG_6__SCAN_IN), .B1(n10965), .Y(n11382));
  OAI21X1 g08134(.A0(n11381), .A1(n11042), .B0(n11382), .Y(n11383));
  AOI21X1 g08135(.A0(n11376), .A1(n12547), .B0(n11383), .Y(n11384));
  NAND4X1 g08136(.A(n11372), .B(n11338), .C(n11322), .D(n11384), .Y(P2_U3040));
  INVX1   g08137(.A(n11035), .Y(n11386));
  NAND2X1 g08138(.A(n11368), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .Y(n11387));
  NOR2X1  g08139(.A(n11368), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .Y(n11388));
  OAI21X1 g08140(.A0(n11388), .A1(n11346), .B0(n11387), .Y(n11389));
  INVX1   g08141(.A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .Y(n11390));
  NOR2X1  g08142(.A(n11351), .B(n11348), .Y(n11391));
  NOR3X1  g08143(.A(n11001), .B(n10996), .C(n8979), .Y(n11392));
  XOR2X1  g08144(.A(n9134), .B(n11392), .Y(n11395));
  NOR2X1  g08145(.A(n11395), .B(n9468), .Y(n11396));
  AOI21X1 g08146(.A0(n9468), .A1(P2_EBX_REG_7__SCAN_IN), .B0(n11396), .Y(n11397));
  XOR2X1  g08147(.A(n11397), .B(n11391), .Y(n11398));
  NAND2X1 g08148(.A(n11398), .B(n11007), .Y(n11399));
  INVX1   g08149(.A(n11366), .Y(n11400));
  NOR2X1  g08150(.A(n11400), .B(n11354), .Y(n11401));
  AOI22X1 g08151(.A0(n9754), .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B0(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(n9993), .Y(n11402));
  AOI22X1 g08152(.A0(n10053), .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B0(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(n10110), .Y(n11403));
  AOI22X1 g08153(.A0(n10168), .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B0(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(n10226), .Y(n11404));
  AOI22X1 g08154(.A0(n10286), .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B0(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(n10344), .Y(n11405));
  NAND4X1 g08155(.A(n11404), .B(n11403), .C(n11402), .D(n11405), .Y(n11406));
  AOI22X1 g08156(.A0(n10629), .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B0(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(n10685), .Y(n11407));
  AOI22X1 g08157(.A0(n10743), .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B0(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(n10799), .Y(n11408));
  AOI22X1 g08158(.A0(n10403), .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B0(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(n10459), .Y(n11409));
  AOI22X1 g08159(.A0(n10517), .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B0(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(n10573), .Y(n11410));
  NAND4X1 g08160(.A(n11409), .B(n11408), .C(n11407), .D(n11410), .Y(n11411));
  OAI21X1 g08161(.A0(n11411), .A1(n11406), .B0(n8975), .Y(n11412));
  OAI21X1 g08162(.A0(n11002), .A1(n8975), .B0(n11412), .Y(n11413));
  INVX1   g08163(.A(n11413), .Y(n11414));
  XOR2X1  g08164(.A(n11414), .B(n11401), .Y(n11415));
  OAI21X1 g08165(.A0(n11415), .A1(n11007), .B0(n11399), .Y(n11416));
  XOR2X1  g08166(.A(n11416), .B(n11390), .Y(n11417));
  XOR2X1  g08167(.A(n11417), .B(n11389), .Y(n11418));
  NOR2X1  g08168(.A(n11367), .B(n11331), .Y(n11419));
  AOI21X1 g08169(.A0(n11367), .A1(n11331), .B0(n11374), .Y(n11420));
  NOR2X1  g08170(.A(n11420), .B(n11419), .Y(n11421));
  XOR2X1  g08171(.A(n11413), .B(n11401), .Y(n11422));
  XOR2X1  g08172(.A(n11422), .B(n11390), .Y(n11423));
  XOR2X1  g08173(.A(n11423), .B(n11421), .Y(n11424));
  NOR4X1  g08174(.A(n11314), .B(n11249), .C(n11246), .D(n11380), .Y(n11425));
  NAND2X1 g08175(.A(n9483), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .Y(n11426));
  NAND2X1 g08176(.A(n9573), .B(P2_EBX_REG_7__SCAN_IN), .Y(n11427));
  AOI22X1 g08177(.A0(P2_REIP_REG_7__SCAN_IN), .A1(n9488), .B0(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(P2_STATE2_REG_1__SCAN_IN), .Y(n11428));
  NAND3X1 g08178(.A(n11428), .B(n11427), .C(n11426), .Y(n11429));
  XOR2X1  g08179(.A(n11429), .B(n11425), .Y(n11430));
  OAI22X1 g08180(.A0(n10978), .A1(n11390), .B0(n8593), .B1(n10966), .Y(n11432));
  AOI21X1 g08181(.A0(n11430), .A1(n11041), .B0(n11432), .Y(n11433));
  NOR4X1  g08182(.A(n11331), .B(n11264), .C(n11188), .D(n11189), .Y(n11434));
  XOR2X1  g08183(.A(n11434), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .Y(n11435));
  NAND2X1 g08184(.A(n11435), .B(n10983), .Y(n11436));
  INVX1   g08185(.A(n10892), .Y(n11437));
  NAND2X1 g08186(.A(n11437), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .Y(n11438));
  AOI21X1 g08187(.A0(n11332), .A1(n11438), .B0(n11330), .Y(n11439));
  INVX1   g08188(.A(n11439), .Y(n11440));
  NOR2X1  g08189(.A(n11333), .B(n11329), .Y(n11441));
  OAI21X1 g08190(.A0(n11441), .A1(n11327), .B0(n11440), .Y(n11442));
  NOR4X1  g08191(.A(n8975), .B(n9468), .C(P2_STATE2_REG_3__SCAN_IN), .D(n11002), .Y(n11443));
  INVX1   g08192(.A(n11443), .Y(n11444));
  AOI22X1 g08193(.A0(n10895), .A1(P2_REIP_REG_7__SCAN_IN), .B0(P2_EAX_REG_7__SCAN_IN), .B1(n10896), .Y(n11445));
  OAI21X1 g08194(.A0(n10892), .A1(n11390), .B0(n11445), .Y(n11446));
  XOR2X1  g08195(.A(n11446), .B(n11444), .Y(n11447));
  INVX1   g08196(.A(n11447), .Y(n11448));
  XOR2X1  g08197(.A(n11448), .B(n11442), .Y(n11449));
  NAND2X1 g08198(.A(n11336), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .Y(n11450));
  XOR2X1  g08199(.A(n11450), .B(n11390), .Y(n11451));
  AOI22X1 g08200(.A0(n11449), .A1(n11096), .B0(n10988), .B1(n11451), .Y(n11452));
  NAND3X1 g08201(.A(n11452), .B(n11436), .C(n11433), .Y(n11453));
  AOI21X1 g08202(.A0(n11424), .A1(n12547), .B0(n11453), .Y(n11454));
  OAI21X1 g08203(.A0(n11418), .A1(n11386), .B0(n11454), .Y(P2_U3039));
  NAND2X1 g08204(.A(n11422), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .Y(n11456));
  NOR2X1  g08205(.A(n11422), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .Y(n11457));
  OAI21X1 g08206(.A0(n11457), .A1(n11421), .B0(n11456), .Y(n11458));
  NOR3X1  g08207(.A(n11414), .B(n11400), .C(n11354), .Y(n11459));
  XOR2X1  g08208(.A(n11459), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .Y(n11460));
  XOR2X1  g08209(.A(n11460), .B(n11458), .Y(n11461));
  NAND2X1 g08210(.A(n11461), .B(n12547), .Y(n11462));
  INVX1   g08211(.A(n11399), .Y(n11463));
  AOI21X1 g08212(.A0(n11422), .A1(n11002), .B0(n11463), .Y(n11464));
  AOI21X1 g08213(.A0(n11464), .A1(n11390), .B0(n11388), .Y(n11465));
  OAI21X1 g08214(.A0(n11345), .A1(n11343), .B0(n11465), .Y(n11466));
  INVX1   g08215(.A(n11466), .Y(n11467));
  AOI21X1 g08216(.A0(n11464), .A1(n11390), .B0(n11387), .Y(n11468));
  AOI21X1 g08217(.A0(n11416), .A1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B0(n11468), .Y(n11469));
  INVX1   g08218(.A(n11469), .Y(n11470));
  NOR2X1  g08219(.A(n11470), .B(n11467), .Y(n11471));
  INVX1   g08220(.A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .Y(n11472));
  INVX1   g08221(.A(n11459), .Y(n11473));
  NAND2X1 g08222(.A(n11397), .B(n11391), .Y(n11474));
  NOR3X1  g08223(.A(n9134), .B(n11392), .C(n9468), .Y(n11477));
  AOI21X1 g08224(.A0(n9468), .A1(P2_EBX_REG_8__SCAN_IN), .B0(n11477), .Y(n11478));
  INVX1   g08225(.A(n11478), .Y(n11479));
  XOR2X1  g08226(.A(n11479), .B(n11474), .Y(n11480));
  NAND2X1 g08227(.A(n11480), .B(n11007), .Y(n11481));
  OAI21X1 g08228(.A0(n11473), .A1(n11007), .B0(n11481), .Y(n11482));
  XOR2X1  g08229(.A(n11482), .B(n11472), .Y(n11483));
  XOR2X1  g08230(.A(n11483), .B(n11471), .Y(n11484));
  NAND2X1 g08231(.A(n11484), .B(n11035), .Y(n11485));
  NAND2X1 g08232(.A(n11429), .B(n11425), .Y(n11486));
  NAND2X1 g08233(.A(n9483), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .Y(n11487));
  NAND2X1 g08234(.A(n9573), .B(P2_EBX_REG_8__SCAN_IN), .Y(n11488));
  AOI22X1 g08235(.A0(P2_REIP_REG_8__SCAN_IN), .A1(n9488), .B0(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(P2_STATE2_REG_1__SCAN_IN), .Y(n11489));
  NAND3X1 g08236(.A(n11489), .B(n11488), .C(n11487), .Y(n11490));
  XOR2X1  g08237(.A(n11490), .B(n11486), .Y(n11491));
  AOI22X1 g08238(.A0(n10979), .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B0(P2_REIP_REG_8__SCAN_IN), .B1(n10965), .Y(n11492));
  OAI21X1 g08239(.A0(n11491), .A1(n11042), .B0(n11492), .Y(n11493));
  INVX1   g08240(.A(n10983), .Y(n11494));
  NAND2X1 g08241(.A(n11434), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .Y(n11495));
  XOR2X1  g08242(.A(n11495), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .Y(n11496));
  NOR2X1  g08243(.A(n11496), .B(n11494), .Y(n11497));
  INVX1   g08244(.A(n11446), .Y(n11498));
  NOR2X1  g08245(.A(n11498), .B(n11444), .Y(n11499));
  NAND2X1 g08246(.A(n11498), .B(n11444), .Y(n11500));
  AOI21X1 g08247(.A0(n11500), .A1(n11442), .B0(n11499), .Y(n11501));
  AOI22X1 g08248(.A0(n8999), .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B0(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(n8980), .Y(n11504));
  AOI22X1 g08249(.A0(n8984), .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B0(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(n8981), .Y(n11507));
  AOI22X1 g08250(.A0(n8983), .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B0(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(n8986), .Y(n11510));
  AOI22X1 g08251(.A0(n8990), .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B0(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(n8987), .Y(n11513));
  NAND4X1 g08252(.A(n11510), .B(n11507), .C(n11504), .D(n11513), .Y(n11514));
  AOI22X1 g08253(.A0(n8993), .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B0(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(n9002), .Y(n11517));
  AOI22X1 g08254(.A0(n9000), .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B0(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(n9003), .Y(n11520));
  AOI22X1 g08255(.A0(n8989), .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B0(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(n8996), .Y(n11523));
  AOI22X1 g08256(.A0(n8994), .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B0(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(n8997), .Y(n11526));
  NAND4X1 g08257(.A(n11523), .B(n11520), .C(n11517), .D(n11526), .Y(n11527));
  NOR2X1  g08258(.A(n11527), .B(n11514), .Y(n11528));
  AOI22X1 g08259(.A0(n10895), .A1(P2_REIP_REG_8__SCAN_IN), .B0(P2_EAX_REG_8__SCAN_IN), .B1(n10896), .Y(n11529));
  OAI21X1 g08260(.A0(n11528), .A1(n10915), .B0(n11529), .Y(n11530));
  AOI21X1 g08261(.A0(n11437), .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B0(n11530), .Y(n11531));
  XOR2X1  g08262(.A(n11531), .B(n11501), .Y(n11532));
  INVX1   g08263(.A(n11532), .Y(n11533));
  NAND3X1 g08264(.A(n11336), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .Y(n11534));
  XOR2X1  g08265(.A(n11534), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .Y(n11535));
  OAI22X1 g08266(.A0(n11533), .A1(n10986), .B0(n10989), .B1(n11535), .Y(n11536));
  NOR3X1  g08267(.A(n11536), .B(n11497), .C(n11493), .Y(n11537));
  NAND3X1 g08268(.A(n11537), .B(n11485), .C(n11462), .Y(P2_U3038));
  NOR2X1  g08269(.A(n11482), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .Y(n11539));
  AOI21X1 g08270(.A0(n11469), .A1(n11466), .B0(n11539), .Y(n11540));
  AOI21X1 g08271(.A0(n11482), .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B0(n11540), .Y(n11541));
  NOR2X1  g08272(.A(n11479), .B(n11474), .Y(n11542));
  AOI21X1 g08273(.A0(n9468), .A1(P2_EBX_REG_9__SCAN_IN), .B0(n11477), .Y(n11543));
  INVX1   g08274(.A(n11543), .Y(n11544));
  NOR3X1  g08275(.A(n11544), .B(n11479), .C(n11474), .Y(n11545));
  INVX1   g08276(.A(n11545), .Y(n11546));
  OAI21X1 g08277(.A0(n11543), .A1(n11542), .B0(n11546), .Y(n11547));
  NOR2X1  g08278(.A(n11547), .B(n11002), .Y(n11548));
  XOR2X1  g08279(.A(n11548), .B(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .Y(n11549));
  XOR2X1  g08280(.A(n11549), .B(n11541), .Y(n11550));
  INVX1   g08281(.A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .Y(n11551));
  NOR2X1  g08282(.A(n11459), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .Y(n11552));
  NOR3X1  g08283(.A(n11552), .B(n11457), .C(n11421), .Y(n11553));
  NOR3X1  g08284(.A(n11552), .B(n11415), .C(n11390), .Y(n11554));
  AOI21X1 g08285(.A0(n11459), .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B0(n11554), .Y(n11555));
  INVX1   g08286(.A(n11555), .Y(n11556));
  NOR2X1  g08287(.A(n11556), .B(n11553), .Y(n11557));
  XOR2X1  g08288(.A(n11557), .B(n11551), .Y(n11558));
  NAND3X1 g08289(.A(n11490), .B(n11429), .C(n11425), .Y(n11559));
  AOI22X1 g08290(.A0(P2_REIP_REG_9__SCAN_IN), .A1(n9488), .B0(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .B1(P2_STATE2_REG_1__SCAN_IN), .Y(n11560));
  INVX1   g08291(.A(n11560), .Y(n11561));
  AOI21X1 g08292(.A0(n9573), .A1(P2_EBX_REG_9__SCAN_IN), .B0(n11561), .Y(n11562));
  OAI21X1 g08293(.A0(n9542), .A1(n11551), .B0(n11562), .Y(n11563));
  INVX1   g08294(.A(n11563), .Y(n11564));
  XOR2X1  g08295(.A(n11564), .B(n11559), .Y(n11565));
  OAI22X1 g08296(.A0(n10978), .A1(n11551), .B0(n8587), .B1(n10966), .Y(n11566));
  AOI21X1 g08297(.A0(n11565), .A1(n11041), .B0(n11566), .Y(n11567));
  NAND3X1 g08298(.A(n11434), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .C(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .Y(n11568));
  XOR2X1  g08299(.A(n11568), .B(n11551), .Y(n11569));
  NAND2X1 g08300(.A(n11569), .B(n10983), .Y(n11570));
  NOR2X1  g08301(.A(n11531), .B(n11501), .Y(n11571));
  AOI22X1 g08302(.A0(n8999), .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B0(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(n8980), .Y(n11572));
  AOI22X1 g08303(.A0(n8984), .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B0(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(n8981), .Y(n11573));
  AOI22X1 g08304(.A0(n8983), .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B0(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(n8986), .Y(n11574));
  AOI22X1 g08305(.A0(n8990), .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B0(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(n8987), .Y(n11575));
  NAND4X1 g08306(.A(n11574), .B(n11573), .C(n11572), .D(n11575), .Y(n11576));
  AOI22X1 g08307(.A0(n8993), .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B0(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(n9002), .Y(n11577));
  AOI22X1 g08308(.A0(n9000), .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B0(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(n9003), .Y(n11578));
  AOI22X1 g08309(.A0(n8989), .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B0(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(n8996), .Y(n11579));
  AOI22X1 g08310(.A0(n8994), .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B0(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(n8997), .Y(n11580));
  NAND4X1 g08311(.A(n11579), .B(n11578), .C(n11577), .D(n11580), .Y(n11581));
  NOR2X1  g08312(.A(n11581), .B(n11576), .Y(n11582));
  AOI22X1 g08313(.A0(n10895), .A1(P2_REIP_REG_9__SCAN_IN), .B0(P2_EAX_REG_9__SCAN_IN), .B1(n10896), .Y(n11583));
  OAI21X1 g08314(.A0(n11582), .A1(n10915), .B0(n11583), .Y(n11584));
  AOI21X1 g08315(.A0(n11437), .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B0(n11584), .Y(n11585));
  XOR2X1  g08316(.A(n11585), .B(n11571), .Y(n11586));
  INVX1   g08317(.A(n11586), .Y(n11587));
  NAND4X1 g08318(.A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .D(n11336), .Y(n11588));
  XOR2X1  g08319(.A(n11588), .B(n11551), .Y(n11589));
  AOI22X1 g08320(.A0(n11587), .A1(n11096), .B0(n10988), .B1(n11589), .Y(n11590));
  NAND3X1 g08321(.A(n11590), .B(n11570), .C(n11567), .Y(n11591));
  AOI21X1 g08322(.A0(n11558), .A1(n12547), .B0(n11591), .Y(n11592));
  OAI21X1 g08323(.A0(n11550), .A1(n11386), .B0(n11592), .Y(P2_U3037));
  INVX1   g08324(.A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .Y(n11594));
  OAI21X1 g08325(.A0(n11556), .A1(n11553), .B0(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .Y(n11595));
  NOR3X1  g08326(.A(n11557), .B(n11594), .C(n11551), .Y(n11596));
  AOI21X1 g08327(.A0(n11595), .A1(n11594), .B0(n11596), .Y(n11597));
  NAND2X1 g08328(.A(n11597), .B(n12547), .Y(n11598));
  OAI22X1 g08329(.A0(n11482), .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B0(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B1(n11548), .Y(n11599));
  AOI21X1 g08330(.A0(n11469), .A1(n11466), .B0(n11599), .Y(n11600));
  NAND2X1 g08331(.A(n11482), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .Y(n11601));
  NOR2X1  g08332(.A(n11548), .B(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .Y(n11602));
  NOR3X1  g08333(.A(n11547), .B(n11002), .C(n11551), .Y(n11603));
  INVX1   g08334(.A(n11603), .Y(n11604));
  OAI21X1 g08335(.A0(n11602), .A1(n11601), .B0(n11604), .Y(n11605));
  NOR2X1  g08336(.A(n11605), .B(n11600), .Y(n11606));
  AOI21X1 g08337(.A0(n9468), .A1(P2_EBX_REG_10__SCAN_IN), .B0(n11477), .Y(n11607));
  XOR2X1  g08338(.A(n11607), .B(n11545), .Y(n11608));
  NAND2X1 g08339(.A(n11608), .B(n11007), .Y(n11609));
  XOR2X1  g08340(.A(n11609), .B(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .Y(n11610));
  XOR2X1  g08341(.A(n11610), .B(n11606), .Y(n11611));
  NAND2X1 g08342(.A(n11611), .B(n11035), .Y(n11612));
  NAND4X1 g08343(.A(n11490), .B(n11429), .C(n11425), .D(n11563), .Y(n11613));
  AOI22X1 g08344(.A0(P2_REIP_REG_10__SCAN_IN), .A1(n9488), .B0(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(P2_STATE2_REG_1__SCAN_IN), .Y(n11614));
  INVX1   g08345(.A(n11614), .Y(n11615));
  AOI21X1 g08346(.A0(n9573), .A1(P2_EBX_REG_10__SCAN_IN), .B0(n11615), .Y(n11616));
  OAI21X1 g08347(.A0(n9542), .A1(n11594), .B0(n11616), .Y(n11617));
  XOR2X1  g08348(.A(n11617), .B(n11613), .Y(n11618));
  AOI22X1 g08349(.A0(n10979), .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B0(P2_REIP_REG_10__SCAN_IN), .B1(n10965), .Y(n11619));
  OAI21X1 g08350(.A0(n11618), .A1(n11042), .B0(n11619), .Y(n11620));
  NAND4X1 g08351(.A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .C(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .D(n11434), .Y(n11621));
  XOR2X1  g08352(.A(n11621), .B(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .Y(n11622));
  NOR2X1  g08353(.A(n11622), .B(n11494), .Y(n11623));
  NOR3X1  g08354(.A(n11585), .B(n11531), .C(n11501), .Y(n11624));
  AOI22X1 g08355(.A0(n8999), .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B0(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(n8980), .Y(n11625));
  AOI22X1 g08356(.A0(n8984), .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B0(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(n8981), .Y(n11626));
  AOI22X1 g08357(.A0(n8983), .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B0(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(n8986), .Y(n11627));
  AOI22X1 g08358(.A0(n8990), .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B0(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(n8987), .Y(n11628));
  NAND4X1 g08359(.A(n11627), .B(n11626), .C(n11625), .D(n11628), .Y(n11629));
  AOI22X1 g08360(.A0(n8993), .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B0(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(n9002), .Y(n11630));
  AOI22X1 g08361(.A0(n9000), .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B0(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(n9003), .Y(n11631));
  AOI22X1 g08362(.A0(n8989), .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B0(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(n8996), .Y(n11632));
  AOI22X1 g08363(.A0(n8994), .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B0(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(n8997), .Y(n11633));
  NAND4X1 g08364(.A(n11632), .B(n11631), .C(n11630), .D(n11633), .Y(n11634));
  NOR2X1  g08365(.A(n11634), .B(n11629), .Y(n11635));
  AOI22X1 g08366(.A0(n10895), .A1(P2_REIP_REG_10__SCAN_IN), .B0(P2_EAX_REG_10__SCAN_IN), .B1(n10896), .Y(n11636));
  OAI21X1 g08367(.A0(n11635), .A1(n10915), .B0(n11636), .Y(n11637));
  AOI21X1 g08368(.A0(n11437), .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B0(n11637), .Y(n11638));
  XOR2X1  g08369(.A(n11638), .B(n11624), .Y(n11639));
  NOR2X1  g08370(.A(n11588), .B(n11551), .Y(n11640));
  XOR2X1  g08371(.A(n11640), .B(n11594), .Y(n11641));
  OAI22X1 g08372(.A0(n11639), .A1(n10986), .B0(n10989), .B1(n11641), .Y(n11642));
  NOR3X1  g08373(.A(n11642), .B(n11623), .C(n11620), .Y(n11643));
  NAND3X1 g08374(.A(n11643), .B(n11612), .C(n11598), .Y(P2_U3036));
  NOR2X1  g08375(.A(n11609), .B(n11594), .Y(n11645));
  AOI21X1 g08376(.A0(n11609), .A1(n11594), .B0(n11606), .Y(n11646));
  NOR2X1  g08377(.A(n11646), .B(n11645), .Y(n11647));
  INVX1   g08378(.A(n11607), .Y(n11648));
  NOR4X1  g08379(.A(n11544), .B(n11479), .C(n11474), .D(n11648), .Y(n11649));
  AOI21X1 g08380(.A0(n9468), .A1(P2_EBX_REG_11__SCAN_IN), .B0(n11477), .Y(n11650));
  NAND3X1 g08381(.A(n11650), .B(n11607), .C(n11545), .Y(n11651));
  OAI21X1 g08382(.A0(n11650), .A1(n11649), .B0(n11651), .Y(n11652));
  NOR2X1  g08383(.A(n11652), .B(n11002), .Y(n11653));
  XOR2X1  g08384(.A(n11653), .B(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .Y(n11654));
  XOR2X1  g08385(.A(n11654), .B(n11647), .Y(n11655));
  NOR2X1  g08386(.A(n11596), .B(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .Y(n11656));
  INVX1   g08387(.A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .Y(n11657));
  NOR4X1  g08388(.A(n11657), .B(n11594), .C(n11551), .D(n11557), .Y(n11658));
  NOR2X1  g08389(.A(n11658), .B(n11656), .Y(n11659));
  INVX1   g08390(.A(n11617), .Y(n11660));
  NOR2X1  g08391(.A(n11660), .B(n11613), .Y(n11661));
  NAND2X1 g08392(.A(n9483), .B(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .Y(n11662));
  NAND2X1 g08393(.A(n9573), .B(P2_EBX_REG_11__SCAN_IN), .Y(n11663));
  AOI22X1 g08394(.A0(P2_REIP_REG_11__SCAN_IN), .A1(n9488), .B0(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(P2_STATE2_REG_1__SCAN_IN), .Y(n11664));
  NAND3X1 g08395(.A(n11664), .B(n11663), .C(n11662), .Y(n11665));
  XOR2X1  g08396(.A(n11665), .B(n11661), .Y(n11666));
  OAI22X1 g08397(.A0(n10978), .A1(n11657), .B0(n8581), .B1(n10966), .Y(n11667));
  AOI21X1 g08398(.A0(n11666), .A1(n11041), .B0(n11667), .Y(n11668));
  NOR2X1  g08399(.A(n11621), .B(n11594), .Y(n11669));
  XOR2X1  g08400(.A(n11669), .B(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .Y(n11670));
  NAND2X1 g08401(.A(n11670), .B(n10983), .Y(n11671));
  NOR4X1  g08402(.A(n11585), .B(n11531), .C(n11501), .D(n11638), .Y(n11672));
  AOI22X1 g08403(.A0(n8999), .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B0(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(n8980), .Y(n11673));
  AOI22X1 g08404(.A0(n8984), .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B0(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(n8981), .Y(n11674));
  AOI22X1 g08405(.A0(n8983), .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B0(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(n8986), .Y(n11675));
  AOI22X1 g08406(.A0(n8990), .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B0(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(n8987), .Y(n11676));
  NAND4X1 g08407(.A(n11675), .B(n11674), .C(n11673), .D(n11676), .Y(n11677));
  AOI22X1 g08408(.A0(n8993), .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B0(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(n9002), .Y(n11678));
  AOI22X1 g08409(.A0(n9000), .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B0(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(n9003), .Y(n11679));
  AOI22X1 g08410(.A0(n8989), .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B0(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(n8996), .Y(n11680));
  AOI22X1 g08411(.A0(n8994), .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B0(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(n8997), .Y(n11681));
  NAND4X1 g08412(.A(n11680), .B(n11679), .C(n11678), .D(n11681), .Y(n11682));
  NOR2X1  g08413(.A(n11682), .B(n11677), .Y(n11683));
  AOI22X1 g08414(.A0(n10895), .A1(P2_REIP_REG_11__SCAN_IN), .B0(P2_EAX_REG_11__SCAN_IN), .B1(n10896), .Y(n11684));
  OAI21X1 g08415(.A0(n11683), .A1(n10915), .B0(n11684), .Y(n11685));
  AOI21X1 g08416(.A0(n11437), .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B0(n11685), .Y(n11686));
  XOR2X1  g08417(.A(n11686), .B(n11672), .Y(n11687));
  INVX1   g08418(.A(n11687), .Y(n11688));
  NOR3X1  g08419(.A(n11588), .B(n11594), .C(n11551), .Y(n11689));
  XOR2X1  g08420(.A(n11689), .B(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .Y(n11690));
  AOI22X1 g08421(.A0(n11688), .A1(n11096), .B0(n10988), .B1(n11690), .Y(n11691));
  NAND3X1 g08422(.A(n11691), .B(n11671), .C(n11668), .Y(n11692));
  AOI21X1 g08423(.A0(n11659), .A1(n12547), .B0(n11692), .Y(n11693));
  OAI21X1 g08424(.A0(n11655), .A1(n11386), .B0(n11693), .Y(P2_U3035));
  NOR2X1  g08425(.A(n11653), .B(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .Y(n11695));
  AOI21X1 g08426(.A0(n11609), .A1(n11594), .B0(n11695), .Y(n11696));
  OAI21X1 g08427(.A0(n11605), .A1(n11600), .B0(n11696), .Y(n11697));
  INVX1   g08428(.A(n11697), .Y(n11698));
  INVX1   g08429(.A(n11695), .Y(n11699));
  NOR3X1  g08430(.A(n11652), .B(n11002), .C(n11657), .Y(n11700));
  AOI21X1 g08431(.A0(n11699), .A1(n11645), .B0(n11700), .Y(n11701));
  INVX1   g08432(.A(n11701), .Y(n11702));
  NOR2X1  g08433(.A(n11702), .B(n11698), .Y(n11703));
  INVX1   g08434(.A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .Y(n11704));
  AOI21X1 g08435(.A0(n9468), .A1(P2_EBX_REG_12__SCAN_IN), .B0(n11477), .Y(n11705));
  INVX1   g08436(.A(n11705), .Y(n11706));
  XOR2X1  g08437(.A(n11706), .B(n11651), .Y(n11707));
  NAND2X1 g08438(.A(n11707), .B(n11007), .Y(n11708));
  XOR2X1  g08439(.A(n11708), .B(n11704), .Y(n11709));
  XOR2X1  g08440(.A(n11709), .B(n11703), .Y(n11710));
  XOR2X1  g08441(.A(n11658), .B(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .Y(n11711));
  NAND2X1 g08442(.A(n11665), .B(n11661), .Y(n11712));
  AOI22X1 g08443(.A0(P2_REIP_REG_12__SCAN_IN), .A1(n9488), .B0(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(P2_STATE2_REG_1__SCAN_IN), .Y(n11713));
  INVX1   g08444(.A(n11713), .Y(n11714));
  AOI21X1 g08445(.A0(n9573), .A1(P2_EBX_REG_12__SCAN_IN), .B0(n11714), .Y(n11715));
  OAI21X1 g08446(.A0(n9542), .A1(n11704), .B0(n11715), .Y(n11716));
  INVX1   g08447(.A(n11716), .Y(n11717));
  XOR2X1  g08448(.A(n11717), .B(n11712), .Y(n11718));
  OAI22X1 g08449(.A0(n10978), .A1(n11704), .B0(n8578), .B1(n10966), .Y(n11719));
  AOI21X1 g08450(.A0(n11718), .A1(n11041), .B0(n11719), .Y(n11720));
  NOR3X1  g08451(.A(n11621), .B(n11657), .C(n11594), .Y(n11721));
  XOR2X1  g08452(.A(n11721), .B(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .Y(n11722));
  NAND2X1 g08453(.A(n11722), .B(n10983), .Y(n11723));
  INVX1   g08454(.A(n11686), .Y(n11724));
  NAND2X1 g08455(.A(n11724), .B(n11672), .Y(n11725));
  AOI22X1 g08456(.A0(n8999), .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B0(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(n8980), .Y(n11726));
  AOI22X1 g08457(.A0(n8984), .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B0(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(n8981), .Y(n11727));
  AOI22X1 g08458(.A0(n8983), .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B0(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(n8986), .Y(n11728));
  AOI22X1 g08459(.A0(n8990), .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B0(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(n8987), .Y(n11729));
  NAND4X1 g08460(.A(n11728), .B(n11727), .C(n11726), .D(n11729), .Y(n11730));
  AOI22X1 g08461(.A0(n8993), .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B0(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(n9002), .Y(n11731));
  AOI22X1 g08462(.A0(n9000), .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B0(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(n9003), .Y(n11732));
  AOI22X1 g08463(.A0(n8989), .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B0(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(n8996), .Y(n11733));
  AOI22X1 g08464(.A0(n8994), .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B0(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(n8997), .Y(n11734));
  NAND4X1 g08465(.A(n11733), .B(n11732), .C(n11731), .D(n11734), .Y(n11735));
  NOR2X1  g08466(.A(n11735), .B(n11730), .Y(n11736));
  AOI22X1 g08467(.A0(n10895), .A1(P2_REIP_REG_12__SCAN_IN), .B0(P2_EAX_REG_12__SCAN_IN), .B1(n10896), .Y(n11737));
  OAI21X1 g08468(.A0(n11736), .A1(n10915), .B0(n11737), .Y(n11738));
  AOI21X1 g08469(.A0(n11437), .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B0(n11738), .Y(n11739));
  INVX1   g08470(.A(n11739), .Y(n11740));
  XOR2X1  g08471(.A(n11740), .B(n11725), .Y(n11741));
  INVX1   g08472(.A(n11741), .Y(n11742));
  NOR4X1  g08473(.A(n11657), .B(n11594), .C(n11551), .D(n11588), .Y(n11743));
  XOR2X1  g08474(.A(n11743), .B(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .Y(n11744));
  AOI22X1 g08475(.A0(n11742), .A1(n11096), .B0(n10988), .B1(n11744), .Y(n11745));
  NAND3X1 g08476(.A(n11745), .B(n11723), .C(n11720), .Y(n11746));
  AOI21X1 g08477(.A0(n11711), .A1(n12547), .B0(n11746), .Y(n11747));
  OAI21X1 g08478(.A0(n11710), .A1(n11386), .B0(n11747), .Y(P2_U3034));
  NOR2X1  g08479(.A(n11708), .B(n11704), .Y(n11749));
  AOI22X1 g08480(.A0(n11701), .A1(n11697), .B0(n11704), .B1(n11708), .Y(n11750));
  NOR2X1  g08481(.A(n11750), .B(n11749), .Y(n11751));
  NOR2X1  g08482(.A(n11706), .B(n11651), .Y(n11752));
  AOI21X1 g08483(.A0(n9468), .A1(P2_EBX_REG_13__SCAN_IN), .B0(n11477), .Y(n11753));
  INVX1   g08484(.A(n11753), .Y(n11754));
  NOR3X1  g08485(.A(n11754), .B(n11706), .C(n11651), .Y(n11755));
  INVX1   g08486(.A(n11755), .Y(n11756));
  OAI21X1 g08487(.A0(n11753), .A1(n11752), .B0(n11756), .Y(n11757));
  NOR2X1  g08488(.A(n11757), .B(n11002), .Y(n11758));
  XOR2X1  g08489(.A(n11758), .B(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .Y(n11759));
  XOR2X1  g08490(.A(n11759), .B(n11751), .Y(n11760));
  INVX1   g08491(.A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .Y(n11761));
  INVX1   g08492(.A(n11557), .Y(n11762));
  NOR4X1  g08493(.A(n11657), .B(n11594), .C(n11551), .D(n11704), .Y(n11763));
  OAI21X1 g08494(.A0(n11556), .A1(n11553), .B0(n11763), .Y(n11764));
  INVX1   g08495(.A(n11763), .Y(n11765));
  NOR2X1  g08496(.A(n11765), .B(n11761), .Y(n11766));
  AOI22X1 g08497(.A0(n11764), .A1(n11761), .B0(n11762), .B1(n11766), .Y(n11767));
  NOR2X1  g08498(.A(n11717), .B(n11712), .Y(n11768));
  NAND2X1 g08499(.A(n9483), .B(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .Y(n11769));
  NAND2X1 g08500(.A(n9573), .B(P2_EBX_REG_13__SCAN_IN), .Y(n11770));
  AOI22X1 g08501(.A0(P2_REIP_REG_13__SCAN_IN), .A1(n9488), .B0(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .B1(P2_STATE2_REG_1__SCAN_IN), .Y(n11771));
  NAND3X1 g08502(.A(n11771), .B(n11770), .C(n11769), .Y(n11772));
  XOR2X1  g08503(.A(n11772), .B(n11768), .Y(n11773));
  OAI22X1 g08504(.A0(n10978), .A1(n11761), .B0(n8575), .B1(n10966), .Y(n11774));
  AOI21X1 g08505(.A0(n11773), .A1(n11041), .B0(n11774), .Y(n11775));
  NOR4X1  g08506(.A(n11704), .B(n11657), .C(n11594), .D(n11621), .Y(n11776));
  XOR2X1  g08507(.A(n11776), .B(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .Y(n11777));
  NAND2X1 g08508(.A(n11777), .B(n10983), .Y(n11778));
  NAND3X1 g08509(.A(n11740), .B(n11724), .C(n11672), .Y(n11779));
  AOI22X1 g08510(.A0(n8999), .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B0(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(n8980), .Y(n11780));
  AOI22X1 g08511(.A0(n8984), .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B0(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(n8981), .Y(n11781));
  AOI22X1 g08512(.A0(n8983), .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B0(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(n8986), .Y(n11782));
  AOI22X1 g08513(.A0(n8990), .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B0(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(n8987), .Y(n11783));
  NAND4X1 g08514(.A(n11782), .B(n11781), .C(n11780), .D(n11783), .Y(n11784));
  AOI22X1 g08515(.A0(n8993), .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B0(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(n9002), .Y(n11785));
  AOI22X1 g08516(.A0(n9000), .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B0(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(n9003), .Y(n11786));
  AOI22X1 g08517(.A0(n8989), .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B0(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(n8996), .Y(n11787));
  AOI22X1 g08518(.A0(n8994), .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B0(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(n8997), .Y(n11788));
  NAND4X1 g08519(.A(n11787), .B(n11786), .C(n11785), .D(n11788), .Y(n11789));
  NOR2X1  g08520(.A(n11789), .B(n11784), .Y(n11790));
  AOI22X1 g08521(.A0(n10895), .A1(P2_REIP_REG_13__SCAN_IN), .B0(P2_EAX_REG_13__SCAN_IN), .B1(n10896), .Y(n11791));
  OAI21X1 g08522(.A0(n11790), .A1(n10915), .B0(n11791), .Y(n11792));
  AOI21X1 g08523(.A0(n11437), .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .B0(n11792), .Y(n11793));
  INVX1   g08524(.A(n11793), .Y(n11794));
  XOR2X1  g08525(.A(n11794), .B(n11779), .Y(n11795));
  INVX1   g08526(.A(n11795), .Y(n11796));
  NAND2X1 g08527(.A(n11743), .B(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .Y(n11797));
  XOR2X1  g08528(.A(n11797), .B(n11761), .Y(n11798));
  AOI22X1 g08529(.A0(n11796), .A1(n11096), .B0(n10988), .B1(n11798), .Y(n11799));
  NAND3X1 g08530(.A(n11799), .B(n11778), .C(n11775), .Y(n11800));
  AOI21X1 g08531(.A0(n11767), .A1(n12547), .B0(n11800), .Y(n11801));
  OAI21X1 g08532(.A0(n11760), .A1(n11386), .B0(n11801), .Y(P2_U3033));
  NAND2X1 g08533(.A(n11708), .B(n11704), .Y(n11803));
  OAI21X1 g08534(.A0(n11758), .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .B0(n11803), .Y(n11804));
  AOI21X1 g08535(.A0(n11701), .A1(n11697), .B0(n11804), .Y(n11805));
  OAI21X1 g08536(.A0(n11758), .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .B0(n11749), .Y(n11806));
  NAND2X1 g08537(.A(n11758), .B(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .Y(n11807));
  NAND2X1 g08538(.A(n11807), .B(n11806), .Y(n11808));
  NOR2X1  g08539(.A(n11808), .B(n11805), .Y(n11809));
  INVX1   g08540(.A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .Y(n11810));
  AOI21X1 g08541(.A0(n9468), .A1(P2_EBX_REG_14__SCAN_IN), .B0(n11477), .Y(n11811));
  XOR2X1  g08542(.A(n11811), .B(n11755), .Y(n11812));
  NAND2X1 g08543(.A(n11812), .B(n11007), .Y(n11813));
  XOR2X1  g08544(.A(n11813), .B(n11810), .Y(n11814));
  XOR2X1  g08545(.A(n11814), .B(n11809), .Y(n11815));
  OAI21X1 g08546(.A0(n11556), .A1(n11553), .B0(n11766), .Y(n11816));
  NOR4X1  g08547(.A(n11557), .B(n11810), .C(n11761), .D(n11765), .Y(n11817));
  AOI21X1 g08548(.A0(n11816), .A1(n11810), .B0(n11817), .Y(n11818));
  NAND4X1 g08549(.A(n11716), .B(n11665), .C(n11661), .D(n11772), .Y(n11819));
  NAND2X1 g08550(.A(n9483), .B(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .Y(n11820));
  NAND2X1 g08551(.A(n9573), .B(P2_EBX_REG_14__SCAN_IN), .Y(n11821));
  AOI22X1 g08552(.A0(P2_REIP_REG_14__SCAN_IN), .A1(n9488), .B0(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(P2_STATE2_REG_1__SCAN_IN), .Y(n11822));
  NAND3X1 g08553(.A(n11822), .B(n11821), .C(n11820), .Y(n11823));
  INVX1   g08554(.A(n11823), .Y(n11824));
  XOR2X1  g08555(.A(n11824), .B(n11819), .Y(n11825));
  OAI22X1 g08556(.A0(n10978), .A1(n11810), .B0(n8572), .B1(n10966), .Y(n11826));
  AOI21X1 g08557(.A0(n11825), .A1(n11041), .B0(n11826), .Y(n11827));
  NAND2X1 g08558(.A(n11776), .B(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .Y(n11828));
  XOR2X1  g08559(.A(n11828), .B(n11810), .Y(n11829));
  NAND2X1 g08560(.A(n11829), .B(n10983), .Y(n11830));
  NAND4X1 g08561(.A(n11740), .B(n11724), .C(n11672), .D(n11794), .Y(n11831));
  AOI22X1 g08562(.A0(n8999), .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B0(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(n8980), .Y(n11832));
  AOI22X1 g08563(.A0(n8984), .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B0(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(n8981), .Y(n11833));
  AOI22X1 g08564(.A0(n8983), .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B0(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(n8986), .Y(n11834));
  AOI22X1 g08565(.A0(n8990), .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B0(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(n8987), .Y(n11835));
  NAND4X1 g08566(.A(n11834), .B(n11833), .C(n11832), .D(n11835), .Y(n11836));
  AOI22X1 g08567(.A0(n8993), .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B0(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(n9002), .Y(n11837));
  AOI22X1 g08568(.A0(n9000), .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B0(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(n9003), .Y(n11838));
  AOI22X1 g08569(.A0(n8989), .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B0(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(n8996), .Y(n11839));
  AOI22X1 g08570(.A0(n8994), .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B0(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(n8997), .Y(n11840));
  NAND4X1 g08571(.A(n11839), .B(n11838), .C(n11837), .D(n11840), .Y(n11841));
  NOR2X1  g08572(.A(n11841), .B(n11836), .Y(n11842));
  AOI22X1 g08573(.A0(n10895), .A1(P2_REIP_REG_14__SCAN_IN), .B0(P2_EAX_REG_14__SCAN_IN), .B1(n10896), .Y(n11843));
  OAI21X1 g08574(.A0(n11842), .A1(n10915), .B0(n11843), .Y(n11844));
  AOI21X1 g08575(.A0(n11437), .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B0(n11844), .Y(n11845));
  INVX1   g08576(.A(n11845), .Y(n11846));
  XOR2X1  g08577(.A(n11846), .B(n11831), .Y(n11847));
  INVX1   g08578(.A(n11847), .Y(n11848));
  NAND3X1 g08579(.A(n11743), .B(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .C(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .Y(n11849));
  XOR2X1  g08580(.A(n11849), .B(n11810), .Y(n11850));
  AOI22X1 g08581(.A0(n11848), .A1(n11096), .B0(n10988), .B1(n11850), .Y(n11851));
  NAND3X1 g08582(.A(n11851), .B(n11830), .C(n11827), .Y(n11852));
  AOI21X1 g08583(.A0(n11818), .A1(n12547), .B0(n11852), .Y(n11853));
  OAI21X1 g08584(.A0(n11815), .A1(n11386), .B0(n11853), .Y(P2_U3032));
  NOR2X1  g08585(.A(n11813), .B(n11810), .Y(n11855));
  INVX1   g08586(.A(n11855), .Y(n11856));
  AOI21X1 g08587(.A0(n11812), .A1(n11007), .B0(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .Y(n11857));
  OAI21X1 g08588(.A0(n11857), .A1(n11809), .B0(n11856), .Y(n11858));
  INVX1   g08589(.A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .Y(n11859));
  INVX1   g08590(.A(n11811), .Y(n11860));
  NOR4X1  g08591(.A(n11754), .B(n11706), .C(n11651), .D(n11860), .Y(n11861));
  AOI21X1 g08592(.A0(n9468), .A1(P2_EBX_REG_15__SCAN_IN), .B0(n11477), .Y(n11862));
  NAND3X1 g08593(.A(n11862), .B(n11811), .C(n11755), .Y(n11863));
  OAI21X1 g08594(.A0(n11862), .A1(n11861), .B0(n11863), .Y(n11864));
  NOR2X1  g08595(.A(n11864), .B(n11002), .Y(n11865));
  XOR2X1  g08596(.A(n11865), .B(n11859), .Y(n11866));
  XOR2X1  g08597(.A(n11866), .B(n11858), .Y(n11867));
  XOR2X1  g08598(.A(n11817), .B(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .Y(n11868));
  NOR2X1  g08599(.A(n11824), .B(n11819), .Y(n11869));
  NAND2X1 g08600(.A(n9483), .B(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .Y(n11870));
  NAND2X1 g08601(.A(n9573), .B(P2_EBX_REG_15__SCAN_IN), .Y(n11871));
  AOI22X1 g08602(.A0(P2_REIP_REG_15__SCAN_IN), .A1(n9488), .B0(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(P2_STATE2_REG_1__SCAN_IN), .Y(n11872));
  NAND3X1 g08603(.A(n11872), .B(n11871), .C(n11870), .Y(n11873));
  XOR2X1  g08604(.A(n11873), .B(n11869), .Y(n11874));
  OAI22X1 g08605(.A0(n10978), .A1(n11859), .B0(n8569), .B1(n10966), .Y(n11875));
  AOI21X1 g08606(.A0(n11874), .A1(n11041), .B0(n11875), .Y(n11876));
  NAND3X1 g08607(.A(n11776), .B(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .C(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .Y(n11877));
  XOR2X1  g08608(.A(n11877), .B(n11859), .Y(n11878));
  NAND2X1 g08609(.A(n11878), .B(n10983), .Y(n11879));
  NOR2X1  g08610(.A(n11845), .B(n11831), .Y(n11880));
  AOI22X1 g08611(.A0(n8999), .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B0(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(n8980), .Y(n11881));
  AOI22X1 g08612(.A0(n8984), .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B0(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(n8981), .Y(n11882));
  AOI22X1 g08613(.A0(n8983), .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B0(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(n8986), .Y(n11883));
  AOI22X1 g08614(.A0(n8990), .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B0(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(n8987), .Y(n11884));
  NAND4X1 g08615(.A(n11883), .B(n11882), .C(n11881), .D(n11884), .Y(n11885));
  AOI22X1 g08616(.A0(n8993), .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B0(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(n9002), .Y(n11886));
  AOI22X1 g08617(.A0(n9000), .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B0(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(n9003), .Y(n11887));
  AOI22X1 g08618(.A0(n8989), .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B0(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(n8996), .Y(n11888));
  AOI22X1 g08619(.A0(n8994), .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B0(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(n8997), .Y(n11889));
  NAND4X1 g08620(.A(n11888), .B(n11887), .C(n11886), .D(n11889), .Y(n11890));
  NOR2X1  g08621(.A(n11890), .B(n11885), .Y(n11891));
  AOI22X1 g08622(.A0(n10895), .A1(P2_REIP_REG_15__SCAN_IN), .B0(P2_EAX_REG_15__SCAN_IN), .B1(n10896), .Y(n11892));
  OAI21X1 g08623(.A0(n11891), .A1(n10915), .B0(n11892), .Y(n11893));
  AOI21X1 g08624(.A0(n11437), .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B0(n11893), .Y(n11894));
  XOR2X1  g08625(.A(n11894), .B(n11880), .Y(n11895));
  INVX1   g08626(.A(n11895), .Y(n11896));
  NAND4X1 g08627(.A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .C(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .D(n11743), .Y(n11897));
  XOR2X1  g08628(.A(n11897), .B(n11859), .Y(n11898));
  AOI22X1 g08629(.A0(n11896), .A1(n11096), .B0(n10988), .B1(n11898), .Y(n11899));
  NAND3X1 g08630(.A(n11899), .B(n11879), .C(n11876), .Y(n11900));
  AOI21X1 g08631(.A0(n11868), .A1(n12547), .B0(n11900), .Y(n11901));
  OAI21X1 g08632(.A0(n11867), .A1(n11386), .B0(n11901), .Y(P2_U3031));
  NOR2X1  g08633(.A(n11865), .B(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .Y(n11903));
  NOR2X1  g08634(.A(n11903), .B(n11857), .Y(n11904));
  OAI21X1 g08635(.A0(n11808), .A1(n11805), .B0(n11904), .Y(n11905));
  INVX1   g08636(.A(n11905), .Y(n11906));
  NOR2X1  g08637(.A(n11903), .B(n11856), .Y(n11907));
  NOR3X1  g08638(.A(n11864), .B(n11002), .C(n11859), .Y(n11908));
  NOR2X1  g08639(.A(n11908), .B(n11907), .Y(n11909));
  INVX1   g08640(.A(n11909), .Y(n11910));
  NOR2X1  g08641(.A(n11910), .B(n11906), .Y(n11911));
  AOI21X1 g08642(.A0(n9468), .A1(P2_EBX_REG_16__SCAN_IN), .B0(n11477), .Y(n11912));
  INVX1   g08643(.A(n11912), .Y(n11913));
  XOR2X1  g08644(.A(n11913), .B(n11863), .Y(n11914));
  INVX1   g08645(.A(n11914), .Y(n11915));
  NOR2X1  g08646(.A(n11915), .B(n11002), .Y(n11916));
  XOR2X1  g08647(.A(n11916), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .Y(n11917));
  XOR2X1  g08648(.A(n11917), .B(n11911), .Y(n11918));
  INVX1   g08649(.A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .Y(n11919));
  NOR4X1  g08650(.A(n11859), .B(n11810), .C(n11761), .D(n11765), .Y(n11920));
  OAI21X1 g08651(.A0(n11556), .A1(n11553), .B0(n11920), .Y(n11921));
  INVX1   g08652(.A(n11920), .Y(n11922));
  NOR3X1  g08653(.A(n11922), .B(n11557), .C(n11919), .Y(n11923));
  AOI21X1 g08654(.A0(n11921), .A1(n11919), .B0(n11923), .Y(n11924));
  NAND2X1 g08655(.A(n11873), .B(n11869), .Y(n11925));
  NAND2X1 g08656(.A(n9483), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .Y(n11926));
  NAND2X1 g08657(.A(n9573), .B(P2_EBX_REG_16__SCAN_IN), .Y(n11927));
  AOI22X1 g08658(.A0(P2_REIP_REG_16__SCAN_IN), .A1(n9488), .B0(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(P2_STATE2_REG_1__SCAN_IN), .Y(n11928));
  NAND3X1 g08659(.A(n11928), .B(n11927), .C(n11926), .Y(n11929));
  INVX1   g08660(.A(n11929), .Y(n11930));
  XOR2X1  g08661(.A(n11930), .B(n11925), .Y(n11931));
  OAI22X1 g08662(.A0(n10978), .A1(n11919), .B0(n8566), .B1(n10966), .Y(n11932));
  AOI21X1 g08663(.A0(n11931), .A1(n11041), .B0(n11932), .Y(n11933));
  NAND4X1 g08664(.A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .C(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .D(n11776), .Y(n11934));
  XOR2X1  g08665(.A(n11934), .B(n11919), .Y(n11935));
  NAND2X1 g08666(.A(n11935), .B(n10983), .Y(n11936));
  NOR3X1  g08667(.A(n11894), .B(n11845), .C(n11831), .Y(n11937));
  AOI22X1 g08668(.A0(n10895), .A1(P2_REIP_REG_16__SCAN_IN), .B0(P2_EAX_REG_16__SCAN_IN), .B1(n10896), .Y(n11938));
  OAI21X1 g08669(.A0(n10892), .A1(n11919), .B0(n11938), .Y(n11939));
  INVX1   g08670(.A(n11939), .Y(n11940));
  XOR2X1  g08671(.A(n11940), .B(n11937), .Y(n11941));
  INVX1   g08672(.A(n11941), .Y(n11942));
  NOR2X1  g08673(.A(n11897), .B(n11859), .Y(n11943));
  XOR2X1  g08674(.A(n11943), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .Y(n11944));
  AOI22X1 g08675(.A0(n11942), .A1(n11096), .B0(n10988), .B1(n11944), .Y(n11945));
  NAND3X1 g08676(.A(n11945), .B(n11936), .C(n11933), .Y(n11946));
  AOI21X1 g08677(.A0(n11924), .A1(n12547), .B0(n11946), .Y(n11947));
  OAI21X1 g08678(.A0(n11918), .A1(n11386), .B0(n11947), .Y(P2_U3030));
  NOR3X1  g08679(.A(n11915), .B(n11002), .C(n11919), .Y(n11949));
  INVX1   g08680(.A(n11949), .Y(n11950));
  OAI22X1 g08681(.A0(n11910), .A1(n11906), .B0(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B1(n11916), .Y(n11951));
  NAND2X1 g08682(.A(n11951), .B(n11950), .Y(n11952));
  INVX1   g08683(.A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .Y(n11953));
  AOI21X1 g08684(.A0(n9468), .A1(P2_EBX_REG_17__SCAN_IN), .B0(n11477), .Y(n11954));
  INVX1   g08685(.A(n11954), .Y(n11955));
  OAI21X1 g08686(.A0(n11913), .A1(n11863), .B0(n11955), .Y(n11956));
  NAND2X1 g08687(.A(n11954), .B(n11912), .Y(n11957));
  OAI21X1 g08688(.A0(n11957), .A1(n11863), .B0(n11956), .Y(n11958));
  NOR2X1  g08689(.A(n11958), .B(n11002), .Y(n11959));
  XOR2X1  g08690(.A(n11959), .B(n11953), .Y(n11960));
  XOR2X1  g08691(.A(n11960), .B(n11952), .Y(n11961));
  XOR2X1  g08692(.A(n11923), .B(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .Y(n11962));
  NOR2X1  g08693(.A(n11930), .B(n11925), .Y(n11963));
  INVX1   g08694(.A(P2_EBX_REG_17__SCAN_IN), .Y(n11964));
  AOI22X1 g08695(.A0(P2_REIP_REG_17__SCAN_IN), .A1(n9488), .B0(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(P2_STATE2_REG_1__SCAN_IN), .Y(n11965));
  OAI21X1 g08696(.A0(n9485), .A1(n11964), .B0(n11965), .Y(n11966));
  AOI21X1 g08697(.A0(n9483), .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .B0(n11966), .Y(n11967));
  XOR2X1  g08698(.A(n11967), .B(n11963), .Y(n11968));
  INVX1   g08699(.A(n11968), .Y(n11969));
  OAI22X1 g08700(.A0(n10978), .A1(n11953), .B0(n8563), .B1(n10966), .Y(n11970));
  AOI21X1 g08701(.A0(n11969), .A1(n11041), .B0(n11970), .Y(n11971));
  NOR2X1  g08702(.A(n11934), .B(n11919), .Y(n11972));
  XOR2X1  g08703(.A(n11972), .B(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .Y(n11973));
  NAND2X1 g08704(.A(n11973), .B(n10983), .Y(n11974));
  NOR4X1  g08705(.A(n11894), .B(n11845), .C(n11831), .D(n11940), .Y(n11975));
  AOI22X1 g08706(.A0(n10895), .A1(P2_REIP_REG_17__SCAN_IN), .B0(P2_EAX_REG_17__SCAN_IN), .B1(n10896), .Y(n11976));
  OAI21X1 g08707(.A0(n10892), .A1(n11953), .B0(n11976), .Y(n11977));
  INVX1   g08708(.A(n11977), .Y(n11978));
  XOR2X1  g08709(.A(n11978), .B(n11975), .Y(n11979));
  INVX1   g08710(.A(n11979), .Y(n11980));
  NOR3X1  g08711(.A(n11897), .B(n11919), .C(n11859), .Y(n11981));
  XOR2X1  g08712(.A(n11981), .B(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .Y(n11982));
  AOI22X1 g08713(.A0(n11980), .A1(n11096), .B0(n10988), .B1(n11982), .Y(n11983));
  NAND3X1 g08714(.A(n11983), .B(n11974), .C(n11971), .Y(n11984));
  AOI21X1 g08715(.A0(n11962), .A1(n12547), .B0(n11984), .Y(n11985));
  OAI21X1 g08716(.A0(n11961), .A1(n11386), .B0(n11985), .Y(P2_U3029));
  OAI22X1 g08717(.A0(n11916), .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B0(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .B1(n11959), .Y(n11987));
  AOI21X1 g08718(.A0(n11909), .A1(n11905), .B0(n11987), .Y(n11988));
  INVX1   g08719(.A(n11959), .Y(n11989));
  OAI21X1 g08720(.A0(n11959), .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .B0(n11949), .Y(n11990));
  OAI21X1 g08721(.A0(n11989), .A1(n11953), .B0(n11990), .Y(n11991));
  NOR2X1  g08722(.A(n11991), .B(n11988), .Y(n11992));
  NOR3X1  g08723(.A(n11955), .B(n11913), .C(n11863), .Y(n11993));
  AOI21X1 g08724(.A0(n9468), .A1(P2_EBX_REG_18__SCAN_IN), .B0(n11477), .Y(n11994));
  XOR2X1  g08725(.A(n11994), .B(n11993), .Y(n11995));
  INVX1   g08726(.A(n11995), .Y(n11996));
  NOR2X1  g08727(.A(n11996), .B(n11002), .Y(n11997));
  XOR2X1  g08728(.A(n11997), .B(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .Y(n11998));
  XOR2X1  g08729(.A(n11998), .B(n11992), .Y(n11999));
  NOR4X1  g08730(.A(n11557), .B(n11953), .C(n11919), .D(n11922), .Y(n12000));
  XOR2X1  g08731(.A(n12000), .B(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .Y(n12001));
  NOR3X1  g08732(.A(n11967), .B(n11930), .C(n11925), .Y(n12002));
  NAND2X1 g08733(.A(n9483), .B(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .Y(n12003));
  NAND2X1 g08734(.A(n9573), .B(P2_EBX_REG_18__SCAN_IN), .Y(n12004));
  AOI22X1 g08735(.A0(P2_REIP_REG_18__SCAN_IN), .A1(n9488), .B0(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(P2_STATE2_REG_1__SCAN_IN), .Y(n12005));
  NAND3X1 g08736(.A(n12005), .B(n12004), .C(n12003), .Y(n12006));
  XOR2X1  g08737(.A(n12006), .B(n12002), .Y(n12007));
  INVX1   g08738(.A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .Y(n12008));
  OAI22X1 g08739(.A0(n10978), .A1(n12008), .B0(n8560), .B1(n10966), .Y(n12009));
  AOI21X1 g08740(.A0(n12007), .A1(n11041), .B0(n12009), .Y(n12010));
  NOR3X1  g08741(.A(n11934), .B(n11953), .C(n11919), .Y(n12011));
  XOR2X1  g08742(.A(n12011), .B(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .Y(n12012));
  NAND2X1 g08743(.A(n12012), .B(n10983), .Y(n12013));
  NAND2X1 g08744(.A(n11977), .B(n11975), .Y(n12014));
  AOI22X1 g08745(.A0(n10895), .A1(P2_REIP_REG_18__SCAN_IN), .B0(P2_EAX_REG_18__SCAN_IN), .B1(n10896), .Y(n12015));
  OAI21X1 g08746(.A0(n10892), .A1(n12008), .B0(n12015), .Y(n12016));
  XOR2X1  g08747(.A(n12016), .B(n12014), .Y(n12017));
  INVX1   g08748(.A(n12017), .Y(n12018));
  NOR4X1  g08749(.A(n11953), .B(n11919), .C(n11859), .D(n11897), .Y(n12019));
  XOR2X1  g08750(.A(n12019), .B(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .Y(n12020));
  AOI22X1 g08751(.A0(n12018), .A1(n11096), .B0(n10988), .B1(n12020), .Y(n12021));
  NAND3X1 g08752(.A(n12021), .B(n12013), .C(n12010), .Y(n12022));
  AOI21X1 g08753(.A0(n12001), .A1(n12547), .B0(n12022), .Y(n12023));
  OAI21X1 g08754(.A0(n11999), .A1(n11386), .B0(n12023), .Y(P2_U3028));
  NAND3X1 g08755(.A(n11995), .B(n11007), .C(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .Y(n12025));
  OAI22X1 g08756(.A0(n11991), .A1(n11988), .B0(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .B1(n11997), .Y(n12026));
  NAND2X1 g08757(.A(n12026), .B(n12025), .Y(n12027));
  INVX1   g08758(.A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .Y(n12028));
  INVX1   g08759(.A(n11994), .Y(n12029));
  NOR3X1  g08760(.A(n12029), .B(n11957), .C(n11863), .Y(n12030));
  AOI21X1 g08761(.A0(n9468), .A1(P2_EBX_REG_19__SCAN_IN), .B0(n11477), .Y(n12031));
  NAND3X1 g08762(.A(n12031), .B(n11994), .C(n11993), .Y(n12032));
  OAI21X1 g08763(.A0(n12031), .A1(n12030), .B0(n12032), .Y(n12033));
  NOR2X1  g08764(.A(n12033), .B(n11002), .Y(n12034));
  XOR2X1  g08765(.A(n12034), .B(n12028), .Y(n12035));
  XOR2X1  g08766(.A(n12035), .B(n12027), .Y(n12036));
  NOR4X1  g08767(.A(n12008), .B(n11953), .C(n11919), .D(n11922), .Y(n12037));
  OAI21X1 g08768(.A0(n11556), .A1(n11553), .B0(n12037), .Y(n12038));
  INVX1   g08769(.A(n12037), .Y(n12039));
  NOR3X1  g08770(.A(n12039), .B(n11557), .C(n12028), .Y(n12040));
  AOI21X1 g08771(.A0(n12038), .A1(n12028), .B0(n12040), .Y(n12041));
  NAND2X1 g08772(.A(n12006), .B(n12002), .Y(n12042));
  NAND2X1 g08773(.A(n9483), .B(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .Y(n12043));
  NAND2X1 g08774(.A(n9573), .B(P2_EBX_REG_19__SCAN_IN), .Y(n12044));
  AOI22X1 g08775(.A0(P2_REIP_REG_19__SCAN_IN), .A1(n9488), .B0(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(P2_STATE2_REG_1__SCAN_IN), .Y(n12045));
  NAND3X1 g08776(.A(n12045), .B(n12044), .C(n12043), .Y(n12046));
  INVX1   g08777(.A(n12046), .Y(n12047));
  XOR2X1  g08778(.A(n12047), .B(n12042), .Y(n12048));
  OAI22X1 g08779(.A0(n10978), .A1(n12028), .B0(n8557), .B1(n10966), .Y(n12049));
  AOI21X1 g08780(.A0(n12048), .A1(n11041), .B0(n12049), .Y(n12050));
  NOR4X1  g08781(.A(n12008), .B(n11953), .C(n11919), .D(n11934), .Y(n12051));
  XOR2X1  g08782(.A(n12051), .B(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .Y(n12052));
  NAND2X1 g08783(.A(n12052), .B(n10983), .Y(n12053));
  NAND3X1 g08784(.A(n12016), .B(n11977), .C(n11975), .Y(n12054));
  AOI22X1 g08785(.A0(n10895), .A1(P2_REIP_REG_19__SCAN_IN), .B0(P2_EAX_REG_19__SCAN_IN), .B1(n10896), .Y(n12055));
  OAI21X1 g08786(.A0(n10892), .A1(n12028), .B0(n12055), .Y(n12056));
  XOR2X1  g08787(.A(n12056), .B(n12054), .Y(n12057));
  INVX1   g08788(.A(n12057), .Y(n12058));
  NAND2X1 g08789(.A(n12019), .B(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .Y(n12059));
  XOR2X1  g08790(.A(n12059), .B(n12028), .Y(n12060));
  AOI22X1 g08791(.A0(n12058), .A1(n11096), .B0(n10988), .B1(n12060), .Y(n12061));
  NAND3X1 g08792(.A(n12061), .B(n12053), .C(n12050), .Y(n12062));
  AOI21X1 g08793(.A0(n12041), .A1(n12547), .B0(n12062), .Y(n12063));
  OAI21X1 g08794(.A0(n12036), .A1(n11386), .B0(n12063), .Y(P2_U3027));
  NOR2X1  g08795(.A(n12034), .B(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .Y(n12065));
  AOI22X1 g08796(.A0(n11997), .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .B0(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .B1(n12034), .Y(n12066));
  OAI22X1 g08797(.A0(n11997), .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .B0(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .B1(n12034), .Y(n12067));
  OAI22X1 g08798(.A0(n12066), .A1(n12065), .B0(n11992), .B1(n12067), .Y(n12068));
  INVX1   g08799(.A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .Y(n12069));
  AOI21X1 g08800(.A0(n9468), .A1(P2_EBX_REG_20__SCAN_IN), .B0(n11477), .Y(n12070));
  INVX1   g08801(.A(n12070), .Y(n12071));
  XOR2X1  g08802(.A(n12071), .B(n12032), .Y(n12072));
  INVX1   g08803(.A(n12072), .Y(n12073));
  NOR2X1  g08804(.A(n12073), .B(n11002), .Y(n12074));
  XOR2X1  g08805(.A(n12074), .B(n12069), .Y(n12075));
  XOR2X1  g08806(.A(n12075), .B(n12068), .Y(n12076));
  NOR2X1  g08807(.A(n12040), .B(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .Y(n12077));
  NOR3X1  g08808(.A(n12039), .B(n12069), .C(n12028), .Y(n12078));
  INVX1   g08809(.A(n12078), .Y(n12079));
  NOR2X1  g08810(.A(n12079), .B(n11557), .Y(n12080));
  NOR2X1  g08811(.A(n12080), .B(n12077), .Y(n12081));
  NOR2X1  g08812(.A(n12047), .B(n12042), .Y(n12082));
  INVX1   g08813(.A(P2_EBX_REG_20__SCAN_IN), .Y(n12083));
  AOI22X1 g08814(.A0(P2_REIP_REG_20__SCAN_IN), .A1(n9488), .B0(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B1(P2_STATE2_REG_1__SCAN_IN), .Y(n12084));
  OAI21X1 g08815(.A0(n9485), .A1(n12083), .B0(n12084), .Y(n12085));
  AOI21X1 g08816(.A0(n9483), .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B0(n12085), .Y(n12086));
  INVX1   g08817(.A(n12086), .Y(n12087));
  XOR2X1  g08818(.A(n12087), .B(n12082), .Y(n12088));
  OAI22X1 g08819(.A0(n10978), .A1(n12069), .B0(n8554), .B1(n10966), .Y(n12089));
  AOI21X1 g08820(.A0(n12088), .A1(n11041), .B0(n12089), .Y(n12090));
  NAND2X1 g08821(.A(n12051), .B(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .Y(n12091));
  XOR2X1  g08822(.A(n12091), .B(n12069), .Y(n12092));
  NAND2X1 g08823(.A(n12092), .B(n10983), .Y(n12093));
  NAND4X1 g08824(.A(n12016), .B(n11977), .C(n11975), .D(n12056), .Y(n12094));
  AOI22X1 g08825(.A0(n10895), .A1(P2_REIP_REG_20__SCAN_IN), .B0(P2_EAX_REG_20__SCAN_IN), .B1(n10896), .Y(n12095));
  OAI21X1 g08826(.A0(n10892), .A1(n12069), .B0(n12095), .Y(n12096));
  XOR2X1  g08827(.A(n12096), .B(n12094), .Y(n12097));
  INVX1   g08828(.A(n12097), .Y(n12098));
  NAND3X1 g08829(.A(n12019), .B(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .C(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .Y(n12099));
  XOR2X1  g08830(.A(n12099), .B(n12069), .Y(n12100));
  AOI22X1 g08831(.A0(n12098), .A1(n11096), .B0(n10988), .B1(n12100), .Y(n12101));
  NAND3X1 g08832(.A(n12101), .B(n12093), .C(n12090), .Y(n12102));
  AOI21X1 g08833(.A0(n12081), .A1(n12547), .B0(n12102), .Y(n12103));
  OAI21X1 g08834(.A0(n12076), .A1(n11386), .B0(n12103), .Y(P2_U3026));
  OAI22X1 g08835(.A0(n12034), .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .B0(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(n12074), .Y(n12105));
  NAND3X1 g08836(.A(n12072), .B(n11007), .C(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .Y(n12106));
  OAI21X1 g08837(.A0(n12105), .A1(n12066), .B0(n12106), .Y(n12107));
  INVX1   g08838(.A(n12107), .Y(n12108));
  OAI21X1 g08839(.A0(n12105), .A1(n12026), .B0(n12108), .Y(n12109));
  INVX1   g08840(.A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .Y(n12110));
  AOI21X1 g08841(.A0(n9468), .A1(P2_EBX_REG_21__SCAN_IN), .B0(n11477), .Y(n12111));
  INVX1   g08842(.A(n12111), .Y(n12112));
  OAI21X1 g08843(.A0(n12071), .A1(n12032), .B0(n12112), .Y(n12113));
  NAND2X1 g08844(.A(n12111), .B(n12070), .Y(n12114));
  OAI21X1 g08845(.A0(n12114), .A1(n12032), .B0(n12113), .Y(n12115));
  NOR2X1  g08846(.A(n12115), .B(n11002), .Y(n12116));
  XOR2X1  g08847(.A(n12116), .B(n12110), .Y(n12117));
  XOR2X1  g08848(.A(n12117), .B(n12109), .Y(n12118));
  XOR2X1  g08849(.A(n12080), .B(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .Y(n12119));
  NOR3X1  g08850(.A(n12086), .B(n12047), .C(n12042), .Y(n12120));
  INVX1   g08851(.A(P2_EBX_REG_21__SCAN_IN), .Y(n12121));
  AOI22X1 g08852(.A0(P2_REIP_REG_21__SCAN_IN), .A1(n9488), .B0(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .B1(P2_STATE2_REG_1__SCAN_IN), .Y(n12122));
  OAI21X1 g08853(.A0(n9485), .A1(n12121), .B0(n12122), .Y(n12123));
  AOI21X1 g08854(.A0(n9483), .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .B0(n12123), .Y(n12124));
  INVX1   g08855(.A(n12124), .Y(n12125));
  XOR2X1  g08856(.A(n12125), .B(n12120), .Y(n12126));
  OAI22X1 g08857(.A0(n10978), .A1(n12110), .B0(n8551), .B1(n10966), .Y(n12127));
  AOI21X1 g08858(.A0(n12126), .A1(n11041), .B0(n12127), .Y(n12128));
  NAND3X1 g08859(.A(n12051), .B(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .C(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .Y(n12129));
  XOR2X1  g08860(.A(n12129), .B(n12110), .Y(n12130));
  NAND2X1 g08861(.A(n12130), .B(n10983), .Y(n12131));
  INVX1   g08862(.A(n12096), .Y(n12132));
  NOR2X1  g08863(.A(n12132), .B(n12094), .Y(n12133));
  AOI22X1 g08864(.A0(n10895), .A1(P2_REIP_REG_21__SCAN_IN), .B0(P2_EAX_REG_21__SCAN_IN), .B1(n10896), .Y(n12134));
  OAI21X1 g08865(.A0(n10892), .A1(n12110), .B0(n12134), .Y(n12135));
  INVX1   g08866(.A(n12135), .Y(n12136));
  XOR2X1  g08867(.A(n12136), .B(n12133), .Y(n12137));
  INVX1   g08868(.A(n12137), .Y(n12138));
  NAND4X1 g08869(.A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .C(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .D(n12019), .Y(n12139));
  XOR2X1  g08870(.A(n12139), .B(n12110), .Y(n12140));
  AOI22X1 g08871(.A0(n12138), .A1(n11096), .B0(n10988), .B1(n12140), .Y(n12141));
  NAND3X1 g08872(.A(n12141), .B(n12131), .C(n12128), .Y(n12142));
  AOI21X1 g08873(.A0(n12119), .A1(n12547), .B0(n12142), .Y(n12143));
  OAI21X1 g08874(.A0(n12118), .A1(n11386), .B0(n12143), .Y(P2_U3025));
  NOR3X1  g08875(.A(n12115), .B(n11002), .C(n12110), .Y(n12145));
  OAI21X1 g08876(.A0(n12115), .A1(n11002), .B0(n12110), .Y(n12146));
  AOI21X1 g08877(.A0(n12146), .A1(n12109), .B0(n12145), .Y(n12147));
  NOR3X1  g08878(.A(n12112), .B(n12071), .C(n12032), .Y(n12148));
  AOI21X1 g08879(.A0(n9468), .A1(P2_EBX_REG_22__SCAN_IN), .B0(n11477), .Y(n12149));
  XOR2X1  g08880(.A(n12149), .B(n12148), .Y(n12150));
  INVX1   g08881(.A(n12150), .Y(n12151));
  NOR2X1  g08882(.A(n12151), .B(n11002), .Y(n12152));
  XOR2X1  g08883(.A(n12152), .B(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .Y(n12153));
  XOR2X1  g08884(.A(n12153), .B(n12147), .Y(n12154));
  INVX1   g08885(.A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .Y(n12155));
  NAND3X1 g08886(.A(n12078), .B(n11762), .C(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .Y(n12156));
  NOR4X1  g08887(.A(n11557), .B(n12155), .C(n12110), .D(n12079), .Y(n12157));
  AOI21X1 g08888(.A0(n12156), .A1(n12155), .B0(n12157), .Y(n12158));
  NOR4X1  g08889(.A(n12086), .B(n12047), .C(n12042), .D(n12124), .Y(n12159));
  INVX1   g08890(.A(P2_EBX_REG_22__SCAN_IN), .Y(n12160));
  AOI22X1 g08891(.A0(P2_REIP_REG_22__SCAN_IN), .A1(n9488), .B0(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(P2_STATE2_REG_1__SCAN_IN), .Y(n12161));
  OAI21X1 g08892(.A0(n9485), .A1(n12160), .B0(n12161), .Y(n12162));
  AOI21X1 g08893(.A0(n9483), .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B0(n12162), .Y(n12163));
  INVX1   g08894(.A(n12163), .Y(n12164));
  XOR2X1  g08895(.A(n12164), .B(n12159), .Y(n12165));
  OAI22X1 g08896(.A0(n10978), .A1(n12155), .B0(n8548), .B1(n10966), .Y(n12166));
  AOI21X1 g08897(.A0(n12165), .A1(n11041), .B0(n12166), .Y(n12167));
  NAND4X1 g08898(.A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .B(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .C(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .D(n12051), .Y(n12168));
  XOR2X1  g08899(.A(n12168), .B(n12155), .Y(n12169));
  NAND2X1 g08900(.A(n12169), .B(n10983), .Y(n12170));
  NOR3X1  g08901(.A(n12136), .B(n12132), .C(n12094), .Y(n12171));
  AOI22X1 g08902(.A0(n10895), .A1(P2_REIP_REG_22__SCAN_IN), .B0(P2_EAX_REG_22__SCAN_IN), .B1(n10896), .Y(n12172));
  OAI21X1 g08903(.A0(n10892), .A1(n12155), .B0(n12172), .Y(n12173));
  INVX1   g08904(.A(n12173), .Y(n12174));
  XOR2X1  g08905(.A(n12174), .B(n12171), .Y(n12175));
  INVX1   g08906(.A(n12175), .Y(n12176));
  NOR2X1  g08907(.A(n12139), .B(n12110), .Y(n12177));
  XOR2X1  g08908(.A(n12177), .B(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .Y(n12178));
  AOI22X1 g08909(.A0(n12176), .A1(n11096), .B0(n10988), .B1(n12178), .Y(n12179));
  NAND3X1 g08910(.A(n12179), .B(n12170), .C(n12167), .Y(n12180));
  AOI21X1 g08911(.A0(n12158), .A1(n12547), .B0(n12180), .Y(n12181));
  OAI21X1 g08912(.A0(n12154), .A1(n11386), .B0(n12181), .Y(P2_U3024));
  AOI21X1 g08913(.A0(n12150), .A1(n11007), .B0(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .Y(n12183));
  INVX1   g08914(.A(n12183), .Y(n12184));
  NAND2X1 g08915(.A(n12184), .B(n12146), .Y(n12185));
  INVX1   g08916(.A(n12185), .Y(n12186));
  NOR3X1  g08917(.A(n12151), .B(n11002), .C(n12155), .Y(n12187));
  AOI21X1 g08918(.A0(n12184), .A1(n12145), .B0(n12187), .Y(n12188));
  INVX1   g08919(.A(n12188), .Y(n12189));
  AOI21X1 g08920(.A0(n12186), .A1(n12109), .B0(n12189), .Y(n12190));
  INVX1   g08921(.A(n12149), .Y(n12191));
  NOR3X1  g08922(.A(n12191), .B(n12114), .C(n12032), .Y(n12192));
  AOI21X1 g08923(.A0(n9468), .A1(P2_EBX_REG_23__SCAN_IN), .B0(n11477), .Y(n12193));
  NAND3X1 g08924(.A(n12193), .B(n12149), .C(n12148), .Y(n12194));
  OAI21X1 g08925(.A0(n12193), .A1(n12192), .B0(n12194), .Y(n12195));
  NOR2X1  g08926(.A(n12195), .B(n11002), .Y(n12196));
  XOR2X1  g08927(.A(n12196), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .Y(n12197));
  XOR2X1  g08928(.A(n12197), .B(n12190), .Y(n12198));
  NOR2X1  g08929(.A(n12157), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .Y(n12199));
  INVX1   g08930(.A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .Y(n12200));
  NOR4X1  g08931(.A(n12200), .B(n12155), .C(n12110), .D(n12079), .Y(n12201));
  INVX1   g08932(.A(n12201), .Y(n12202));
  NOR2X1  g08933(.A(n12202), .B(n11557), .Y(n12203));
  NOR2X1  g08934(.A(n12203), .B(n12199), .Y(n12204));
  NAND2X1 g08935(.A(n12164), .B(n12159), .Y(n12205));
  NAND2X1 g08936(.A(n9483), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .Y(n12206));
  NAND2X1 g08937(.A(n9573), .B(P2_EBX_REG_23__SCAN_IN), .Y(n12207));
  AOI22X1 g08938(.A0(P2_REIP_REG_23__SCAN_IN), .A1(n9488), .B0(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .B1(P2_STATE2_REG_1__SCAN_IN), .Y(n12208));
  NAND3X1 g08939(.A(n12208), .B(n12207), .C(n12206), .Y(n12209));
  INVX1   g08940(.A(n12209), .Y(n12210));
  XOR2X1  g08941(.A(n12210), .B(n12205), .Y(n12211));
  OAI22X1 g08942(.A0(n10978), .A1(n12200), .B0(n8545), .B1(n10966), .Y(n12212));
  AOI21X1 g08943(.A0(n12211), .A1(n11041), .B0(n12212), .Y(n12213));
  NOR2X1  g08944(.A(n12168), .B(n12155), .Y(n12214));
  XOR2X1  g08945(.A(n12214), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .Y(n12215));
  NAND2X1 g08946(.A(n12215), .B(n10983), .Y(n12216));
  NOR4X1  g08947(.A(n12136), .B(n12132), .C(n12094), .D(n12174), .Y(n12217));
  AOI22X1 g08948(.A0(n10895), .A1(P2_REIP_REG_23__SCAN_IN), .B0(P2_EAX_REG_23__SCAN_IN), .B1(n10896), .Y(n12218));
  OAI21X1 g08949(.A0(n10892), .A1(n12200), .B0(n12218), .Y(n12219));
  INVX1   g08950(.A(n12219), .Y(n12220));
  XOR2X1  g08951(.A(n12220), .B(n12217), .Y(n12221));
  INVX1   g08952(.A(n12221), .Y(n12222));
  NOR3X1  g08953(.A(n12139), .B(n12155), .C(n12110), .Y(n12223));
  XOR2X1  g08954(.A(n12223), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .Y(n12224));
  AOI22X1 g08955(.A0(n12222), .A1(n11096), .B0(n10988), .B1(n12224), .Y(n12225));
  NAND3X1 g08956(.A(n12225), .B(n12216), .C(n12213), .Y(n12226));
  AOI21X1 g08957(.A0(n12204), .A1(n12547), .B0(n12226), .Y(n12227));
  OAI21X1 g08958(.A0(n12198), .A1(n11386), .B0(n12227), .Y(P2_U3023));
  NOR3X1  g08959(.A(n12195), .B(n11002), .C(n12200), .Y(n12229));
  INVX1   g08960(.A(n12229), .Y(n12230));
  NOR2X1  g08961(.A(n12196), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .Y(n12231));
  OAI21X1 g08962(.A0(n12231), .A1(n12190), .B0(n12230), .Y(n12232));
  INVX1   g08963(.A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .Y(n12233));
  AOI21X1 g08964(.A0(n9468), .A1(P2_EBX_REG_24__SCAN_IN), .B0(n11477), .Y(n12234));
  INVX1   g08965(.A(n12234), .Y(n12235));
  XOR2X1  g08966(.A(n12235), .B(n12194), .Y(n12236));
  INVX1   g08967(.A(n12236), .Y(n12237));
  NOR2X1  g08968(.A(n12237), .B(n11002), .Y(n12238));
  XOR2X1  g08969(.A(n12238), .B(n12233), .Y(n12239));
  XOR2X1  g08970(.A(n12239), .B(n12232), .Y(n12240));
  XOR2X1  g08971(.A(n12203), .B(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .Y(n12241));
  NOR2X1  g08972(.A(n12210), .B(n12205), .Y(n12242));
  INVX1   g08973(.A(P2_EBX_REG_24__SCAN_IN), .Y(n12243));
  AOI22X1 g08974(.A0(P2_REIP_REG_24__SCAN_IN), .A1(n9488), .B0(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B1(P2_STATE2_REG_1__SCAN_IN), .Y(n12244));
  OAI21X1 g08975(.A0(n9485), .A1(n12243), .B0(n12244), .Y(n12245));
  AOI21X1 g08976(.A0(n9483), .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B0(n12245), .Y(n12246));
  INVX1   g08977(.A(n12246), .Y(n12247));
  XOR2X1  g08978(.A(n12247), .B(n12242), .Y(n12248));
  OAI22X1 g08979(.A0(n10978), .A1(n12233), .B0(n8542), .B1(n10966), .Y(n12249));
  AOI21X1 g08980(.A0(n12248), .A1(n11041), .B0(n12249), .Y(n12250));
  NOR3X1  g08981(.A(n12168), .B(n12200), .C(n12155), .Y(n12251));
  XOR2X1  g08982(.A(n12251), .B(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .Y(n12252));
  NAND2X1 g08983(.A(n12252), .B(n10983), .Y(n12253));
  NAND2X1 g08984(.A(n12219), .B(n12217), .Y(n12254));
  AOI22X1 g08985(.A0(n10895), .A1(P2_REIP_REG_24__SCAN_IN), .B0(P2_EAX_REG_24__SCAN_IN), .B1(n10896), .Y(n12255));
  OAI21X1 g08986(.A0(n10892), .A1(n12233), .B0(n12255), .Y(n12256));
  XOR2X1  g08987(.A(n12256), .B(n12254), .Y(n12257));
  INVX1   g08988(.A(n12257), .Y(n12258));
  NOR4X1  g08989(.A(n12200), .B(n12155), .C(n12110), .D(n12139), .Y(n12259));
  XOR2X1  g08990(.A(n12259), .B(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .Y(n12260));
  AOI22X1 g08991(.A0(n12258), .A1(n11096), .B0(n10988), .B1(n12260), .Y(n12261));
  NAND3X1 g08992(.A(n12261), .B(n12253), .C(n12250), .Y(n12262));
  AOI21X1 g08993(.A0(n12241), .A1(n12547), .B0(n12262), .Y(n12263));
  OAI21X1 g08994(.A0(n12240), .A1(n11386), .B0(n12263), .Y(P2_U3022));
  INVX1   g08995(.A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .Y(n12265));
  AOI21X1 g08996(.A0(n12236), .A1(n11007), .B0(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .Y(n12266));
  NOR2X1  g08997(.A(n12266), .B(n12231), .Y(n12267));
  INVX1   g08998(.A(n12267), .Y(n12268));
  NOR4X1  g08999(.A(n12195), .B(n11002), .C(n12200), .D(n12266), .Y(n12269));
  AOI21X1 g09000(.A0(n12238), .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B0(n12269), .Y(n12270));
  OAI21X1 g09001(.A0(n12268), .A1(n12190), .B0(n12270), .Y(n12271));
  XOR2X1  g09002(.A(n12271), .B(n12265), .Y(n12272));
  AOI21X1 g09003(.A0(n9468), .A1(P2_EBX_REG_25__SCAN_IN), .B0(n11477), .Y(n12273));
  INVX1   g09004(.A(n12273), .Y(n12274));
  OAI21X1 g09005(.A0(n12235), .A1(n12194), .B0(n12274), .Y(n12275));
  NAND2X1 g09006(.A(n12273), .B(n12234), .Y(n12276));
  OAI21X1 g09007(.A0(n12276), .A1(n12194), .B0(n12275), .Y(n12277));
  NOR2X1  g09008(.A(n12277), .B(n11002), .Y(n12278));
  XOR2X1  g09009(.A(n12278), .B(n12272), .Y(n12279));
  NOR3X1  g09010(.A(n12202), .B(n11557), .C(n12233), .Y(n12280));
  XOR2X1  g09011(.A(n12280), .B(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .Y(n12281));
  NOR3X1  g09012(.A(n12246), .B(n12210), .C(n12205), .Y(n12282));
  NAND2X1 g09013(.A(n9483), .B(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .Y(n12283));
  NAND2X1 g09014(.A(n9573), .B(P2_EBX_REG_25__SCAN_IN), .Y(n12284));
  AOI22X1 g09015(.A0(P2_REIP_REG_25__SCAN_IN), .A1(n9488), .B0(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .B1(P2_STATE2_REG_1__SCAN_IN), .Y(n12285));
  NAND3X1 g09016(.A(n12285), .B(n12284), .C(n12283), .Y(n12286));
  XOR2X1  g09017(.A(n12286), .B(n12282), .Y(n12287));
  OAI22X1 g09018(.A0(n10978), .A1(n12265), .B0(n8539), .B1(n10966), .Y(n12288));
  AOI21X1 g09019(.A0(n12287), .A1(n11041), .B0(n12288), .Y(n12289));
  NOR4X1  g09020(.A(n12233), .B(n12200), .C(n12155), .D(n12168), .Y(n12290));
  XOR2X1  g09021(.A(n12290), .B(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .Y(n12291));
  NAND2X1 g09022(.A(n12291), .B(n10983), .Y(n12292));
  NAND3X1 g09023(.A(n12256), .B(n12219), .C(n12217), .Y(n12293));
  AOI22X1 g09024(.A0(n10895), .A1(P2_REIP_REG_25__SCAN_IN), .B0(P2_EAX_REG_25__SCAN_IN), .B1(n10896), .Y(n12294));
  OAI21X1 g09025(.A0(n10892), .A1(n12265), .B0(n12294), .Y(n12295));
  XOR2X1  g09026(.A(n12295), .B(n12293), .Y(n12296));
  INVX1   g09027(.A(n12296), .Y(n12297));
  NAND2X1 g09028(.A(n12259), .B(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .Y(n12298));
  XOR2X1  g09029(.A(n12298), .B(n12265), .Y(n12299));
  AOI22X1 g09030(.A0(n12297), .A1(n11096), .B0(n10988), .B1(n12299), .Y(n12300));
  NAND3X1 g09031(.A(n12300), .B(n12292), .C(n12289), .Y(n12301));
  AOI21X1 g09032(.A0(n12281), .A1(n12547), .B0(n12301), .Y(n12302));
  OAI21X1 g09033(.A0(n12279), .A1(n11386), .B0(n12302), .Y(P2_U3021));
  NAND2X1 g09034(.A(n12271), .B(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .Y(n12304));
  OAI21X1 g09035(.A0(n12271), .A1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B0(n12278), .Y(n12305));
  NAND2X1 g09036(.A(n12305), .B(n12304), .Y(n12306));
  NOR3X1  g09037(.A(n12274), .B(n12235), .C(n12194), .Y(n12307));
  AOI21X1 g09038(.A0(n9468), .A1(P2_EBX_REG_26__SCAN_IN), .B0(n11477), .Y(n12308));
  XOR2X1  g09039(.A(n12308), .B(n12307), .Y(n12309));
  INVX1   g09040(.A(n12309), .Y(n12310));
  NOR2X1  g09041(.A(n12310), .B(n11002), .Y(n12311));
  XOR2X1  g09042(.A(n12311), .B(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .Y(n12312));
  XOR2X1  g09043(.A(n12312), .B(n12306), .Y(n12313));
  NAND2X1 g09044(.A(n12313), .B(n11035), .Y(n12314));
  INVX1   g09045(.A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .Y(n12315));
  NAND4X1 g09046(.A(n11762), .B(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .C(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .D(n12201), .Y(n12316));
  NOR4X1  g09047(.A(n12315), .B(n12265), .C(n12233), .D(n12202), .Y(n12317));
  INVX1   g09048(.A(n12317), .Y(n12318));
  NOR2X1  g09049(.A(n12318), .B(n11557), .Y(n12319));
  AOI21X1 g09050(.A0(n12316), .A1(n12315), .B0(n12319), .Y(n12320));
  NAND2X1 g09051(.A(n12320), .B(n12547), .Y(n12321));
  NAND2X1 g09052(.A(n12286), .B(n12282), .Y(n12322));
  INVX1   g09053(.A(P2_EBX_REG_26__SCAN_IN), .Y(n12323));
  AOI22X1 g09054(.A0(P2_REIP_REG_26__SCAN_IN), .A1(n9488), .B0(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .B1(P2_STATE2_REG_1__SCAN_IN), .Y(n12324));
  OAI21X1 g09055(.A0(n9485), .A1(n12323), .B0(n12324), .Y(n12325));
  AOI21X1 g09056(.A0(n9483), .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B0(n12325), .Y(n12326));
  XOR2X1  g09057(.A(n12326), .B(n12322), .Y(n12327));
  OAI22X1 g09058(.A0(n10978), .A1(n12315), .B0(n8536), .B1(n10966), .Y(n12328));
  AOI21X1 g09059(.A0(n12327), .A1(n11041), .B0(n12328), .Y(n12329));
  NAND2X1 g09060(.A(n12290), .B(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .Y(n12330));
  XOR2X1  g09061(.A(n12330), .B(n12315), .Y(n12331));
  NAND4X1 g09062(.A(n12256), .B(n12219), .C(n12217), .D(n12295), .Y(n12332));
  AOI22X1 g09063(.A0(n10895), .A1(P2_REIP_REG_26__SCAN_IN), .B0(P2_EAX_REG_26__SCAN_IN), .B1(n10896), .Y(n12333));
  OAI21X1 g09064(.A0(n10892), .A1(n12315), .B0(n12333), .Y(n12334));
  XOR2X1  g09065(.A(n12334), .B(n12332), .Y(n12335));
  NAND3X1 g09066(.A(n12259), .B(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .C(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .Y(n12336));
  XOR2X1  g09067(.A(n12336), .B(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .Y(n12337));
  OAI22X1 g09068(.A0(n12335), .A1(n10986), .B0(n10989), .B1(n12337), .Y(n12338));
  AOI21X1 g09069(.A0(n12331), .A1(n10983), .B0(n12338), .Y(n12339));
  NAND4X1 g09070(.A(n12329), .B(n12321), .C(n12314), .D(n12339), .Y(P2_U3020));
  NOR3X1  g09071(.A(n12310), .B(n11002), .C(n12315), .Y(n12341));
  OAI21X1 g09072(.A0(n12310), .A1(n11002), .B0(n12315), .Y(n12342));
  AOI21X1 g09073(.A0(n12342), .A1(n12306), .B0(n12341), .Y(n12343));
  INVX1   g09074(.A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .Y(n12344));
  INVX1   g09075(.A(n12308), .Y(n12345));
  NOR3X1  g09076(.A(n12345), .B(n12276), .C(n12194), .Y(n12346));
  AOI21X1 g09077(.A0(n9468), .A1(P2_EBX_REG_27__SCAN_IN), .B0(n11477), .Y(n12347));
  NAND3X1 g09078(.A(n12347), .B(n12308), .C(n12307), .Y(n12348));
  OAI21X1 g09079(.A0(n12347), .A1(n12346), .B0(n12348), .Y(n12349));
  NOR2X1  g09080(.A(n12349), .B(n11002), .Y(n12350));
  XOR2X1  g09081(.A(n12350), .B(n12344), .Y(n12351));
  XOR2X1  g09082(.A(n12351), .B(n12343), .Y(n12352));
  NAND2X1 g09083(.A(n12352), .B(n11035), .Y(n12353));
  XOR2X1  g09084(.A(n12319), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .Y(n12354));
  NAND2X1 g09085(.A(n12354), .B(n12547), .Y(n12355));
  NOR2X1  g09086(.A(n12326), .B(n12322), .Y(n12356));
  NAND2X1 g09087(.A(n9483), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .Y(n12357));
  NAND2X1 g09088(.A(n9573), .B(P2_EBX_REG_27__SCAN_IN), .Y(n12358));
  AOI22X1 g09089(.A0(P2_REIP_REG_27__SCAN_IN), .A1(n9488), .B0(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .B1(P2_STATE2_REG_1__SCAN_IN), .Y(n12359));
  NAND3X1 g09090(.A(n12359), .B(n12358), .C(n12357), .Y(n12360));
  XOR2X1  g09091(.A(n12360), .B(n12356), .Y(n12361));
  OAI22X1 g09092(.A0(n10978), .A1(n12344), .B0(n8533), .B1(n10966), .Y(n12362));
  AOI21X1 g09093(.A0(n12361), .A1(n11041), .B0(n12362), .Y(n12363));
  NAND3X1 g09094(.A(n12290), .B(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .C(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .Y(n12364));
  XOR2X1  g09095(.A(n12364), .B(n12344), .Y(n12365));
  INVX1   g09096(.A(n12334), .Y(n12366));
  NOR2X1  g09097(.A(n12366), .B(n12332), .Y(n12367));
  AOI22X1 g09098(.A0(n10895), .A1(P2_REIP_REG_27__SCAN_IN), .B0(P2_EAX_REG_27__SCAN_IN), .B1(n10896), .Y(n12368));
  OAI21X1 g09099(.A0(n10892), .A1(n12344), .B0(n12368), .Y(n12369));
  INVX1   g09100(.A(n12369), .Y(n12370));
  XOR2X1  g09101(.A(n12370), .B(n12367), .Y(n12371));
  NAND4X1 g09102(.A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .C(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .D(n12259), .Y(n12372));
  XOR2X1  g09103(.A(n12372), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .Y(n12373));
  OAI22X1 g09104(.A0(n12371), .A1(n10986), .B0(n10989), .B1(n12373), .Y(n12374));
  AOI21X1 g09105(.A0(n12365), .A1(n10983), .B0(n12374), .Y(n12375));
  NAND4X1 g09106(.A(n12363), .B(n12355), .C(n12353), .D(n12375), .Y(P2_U3019));
  INVX1   g09107(.A(n12350), .Y(n12377));
  OAI21X1 g09108(.A0(n12350), .A1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B0(n12341), .Y(n12378));
  OAI21X1 g09109(.A0(n12377), .A1(n12344), .B0(n12378), .Y(n12379));
  OAI21X1 g09110(.A0(n12350), .A1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B0(n12342), .Y(n12380));
  AOI21X1 g09111(.A0(n12305), .A1(n12304), .B0(n12380), .Y(n12381));
  NOR2X1  g09112(.A(n12381), .B(n12379), .Y(n12382));
  INVX1   g09113(.A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .Y(n12383));
  AOI21X1 g09114(.A0(n9468), .A1(P2_EBX_REG_28__SCAN_IN), .B0(n11477), .Y(n12384));
  INVX1   g09115(.A(n12384), .Y(n12385));
  XOR2X1  g09116(.A(n12385), .B(n12348), .Y(n12386));
  NAND2X1 g09117(.A(n12386), .B(n11007), .Y(n12387));
  XOR2X1  g09118(.A(n12387), .B(n12383), .Y(n12388));
  XOR2X1  g09119(.A(n12388), .B(n12382), .Y(n12389));
  NAND3X1 g09120(.A(n12317), .B(n11762), .C(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .Y(n12390));
  NAND2X1 g09121(.A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .Y(n12391));
  NOR3X1  g09122(.A(n12391), .B(n12318), .C(n11557), .Y(n12392));
  AOI21X1 g09123(.A0(n12390), .A1(n12383), .B0(n12392), .Y(n12393));
  NOR3X1  g09124(.A(n12370), .B(n12366), .C(n12332), .Y(n12394));
  AOI22X1 g09125(.A0(n10895), .A1(P2_REIP_REG_28__SCAN_IN), .B0(P2_EAX_REG_28__SCAN_IN), .B1(n10896), .Y(n12395));
  OAI21X1 g09126(.A0(n10892), .A1(n12383), .B0(n12395), .Y(n12396));
  INVX1   g09127(.A(n12396), .Y(n12397));
  XOR2X1  g09128(.A(n12397), .B(n12394), .Y(n12398));
  INVX1   g09129(.A(n12398), .Y(n12399));
  NAND2X1 g09130(.A(n12399), .B(n11096), .Y(n12400));
  NAND2X1 g09131(.A(n12360), .B(n12356), .Y(n12401));
  NAND2X1 g09132(.A(n9483), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .Y(n12402));
  NAND2X1 g09133(.A(n9573), .B(P2_EBX_REG_28__SCAN_IN), .Y(n12403));
  AOI22X1 g09134(.A0(P2_REIP_REG_28__SCAN_IN), .A1(n9488), .B0(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .B1(P2_STATE2_REG_1__SCAN_IN), .Y(n12404));
  NAND3X1 g09135(.A(n12404), .B(n12403), .C(n12402), .Y(n12405));
  XOR2X1  g09136(.A(n12405), .B(n12401), .Y(n12406));
  INVX1   g09137(.A(n12406), .Y(n12407));
  OAI22X1 g09138(.A0(n10978), .A1(n12383), .B0(n8530), .B1(n10966), .Y(n12408));
  AOI21X1 g09139(.A0(n12407), .A1(n11041), .B0(n12408), .Y(n12409));
  NOR2X1  g09140(.A(n12372), .B(n12344), .Y(n12410));
  XOR2X1  g09141(.A(n12410), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .Y(n12411));
  NAND4X1 g09142(.A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .C(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .D(n12290), .Y(n12412));
  XOR2X1  g09143(.A(n12412), .B(n12383), .Y(n12413));
  AOI22X1 g09144(.A0(n12411), .A1(n10988), .B0(n10983), .B1(n12413), .Y(n12414));
  NAND3X1 g09145(.A(n12414), .B(n12409), .C(n12400), .Y(n12415));
  AOI21X1 g09146(.A0(n12393), .A1(n12547), .B0(n12415), .Y(n12416));
  OAI21X1 g09147(.A0(n12389), .A1(n11386), .B0(n12416), .Y(P2_U3018));
  AOI21X1 g09148(.A0(n12387), .A1(n12383), .B0(n12380), .Y(n12418));
  INVX1   g09149(.A(n12418), .Y(n12419));
  AOI21X1 g09150(.A0(n12305), .A1(n12304), .B0(n12419), .Y(n12420));
  NAND2X1 g09151(.A(n12387), .B(n12383), .Y(n12421));
  NAND2X1 g09152(.A(n12421), .B(n12379), .Y(n12422));
  NAND3X1 g09153(.A(n12386), .B(n11007), .C(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .Y(n12423));
  NAND2X1 g09154(.A(n12423), .B(n12422), .Y(n12424));
  NOR2X1  g09155(.A(n12424), .B(n12420), .Y(n12425));
  AOI21X1 g09156(.A0(n9468), .A1(P2_EBX_REG_29__SCAN_IN), .B0(n11477), .Y(n12426));
  INVX1   g09157(.A(n12426), .Y(n12427));
  OAI21X1 g09158(.A0(n12385), .A1(n12348), .B0(n12427), .Y(n12428));
  NAND2X1 g09159(.A(n12426), .B(n12384), .Y(n12429));
  OAI21X1 g09160(.A0(n12429), .A1(n12348), .B0(n12428), .Y(n12430));
  NOR2X1  g09161(.A(n12430), .B(n11002), .Y(n12431));
  XOR2X1  g09162(.A(n12431), .B(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .Y(n12432));
  XOR2X1  g09163(.A(n12432), .B(n12425), .Y(n12433));
  NOR2X1  g09164(.A(n12392), .B(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .Y(n12434));
  INVX1   g09165(.A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .Y(n12435));
  NOR4X1  g09166(.A(n12318), .B(n11557), .C(n12435), .D(n12391), .Y(n12436));
  NOR2X1  g09167(.A(n12436), .B(n12434), .Y(n12437));
  NOR4X1  g09168(.A(n12370), .B(n12366), .C(n12332), .D(n12397), .Y(n12438));
  AOI22X1 g09169(.A0(n10895), .A1(P2_REIP_REG_29__SCAN_IN), .B0(P2_EAX_REG_29__SCAN_IN), .B1(n10896), .Y(n12439));
  OAI21X1 g09170(.A0(n10892), .A1(n12435), .B0(n12439), .Y(n12440));
  INVX1   g09171(.A(n12440), .Y(n12441));
  XOR2X1  g09172(.A(n12441), .B(n12438), .Y(n12442));
  NAND3X1 g09173(.A(n12405), .B(n12360), .C(n12356), .Y(n12443));
  NAND2X1 g09174(.A(n9483), .B(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .Y(n12444));
  NAND2X1 g09175(.A(n9573), .B(P2_EBX_REG_29__SCAN_IN), .Y(n12445));
  AOI22X1 g09176(.A0(P2_REIP_REG_29__SCAN_IN), .A1(n9488), .B0(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B1(P2_STATE2_REG_1__SCAN_IN), .Y(n12446));
  NAND3X1 g09177(.A(n12446), .B(n12445), .C(n12444), .Y(n12447));
  XOR2X1  g09178(.A(n12447), .B(n12443), .Y(n12448));
  NOR2X1  g09179(.A(n12448), .B(n11042), .Y(n12449));
  NOR2X1  g09180(.A(n12412), .B(n12383), .Y(n12450));
  XOR2X1  g09181(.A(n12450), .B(n12435), .Y(n12451));
  NOR2X1  g09182(.A(n12451), .B(n11494), .Y(n12452));
  NOR3X1  g09183(.A(n12372), .B(n12383), .C(n12344), .Y(n12453));
  XOR2X1  g09184(.A(n12453), .B(n12435), .Y(n12454));
  AOI22X1 g09185(.A0(n10979), .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .B0(P2_REIP_REG_29__SCAN_IN), .B1(n10965), .Y(n12455));
  OAI21X1 g09186(.A0(n12454), .A1(n10989), .B0(n12455), .Y(n12456));
  NOR3X1  g09187(.A(n12456), .B(n12452), .C(n12449), .Y(n12457));
  OAI21X1 g09188(.A0(n12442), .A1(n10986), .B0(n12457), .Y(n12458));
  AOI21X1 g09189(.A0(n12437), .A1(n12547), .B0(n12458), .Y(n12459));
  OAI21X1 g09190(.A0(n12433), .A1(n11386), .B0(n12459), .Y(P2_U3017));
  NOR3X1  g09191(.A(n12430), .B(n11002), .C(n12435), .Y(n12461));
  INVX1   g09192(.A(n12461), .Y(n12462));
  OAI22X1 g09193(.A0(n12424), .A1(n12420), .B0(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .B1(n12431), .Y(n12463));
  NAND2X1 g09194(.A(n12463), .B(n12462), .Y(n12464));
  NOR3X1  g09195(.A(n12427), .B(n12385), .C(n12348), .Y(n12465));
  AOI21X1 g09196(.A0(n9468), .A1(P2_EBX_REG_30__SCAN_IN), .B0(n11477), .Y(n12466));
  XOR2X1  g09197(.A(n12466), .B(n12465), .Y(n12467));
  NAND2X1 g09198(.A(n12467), .B(n11007), .Y(n12468));
  XOR2X1  g09199(.A(n12468), .B(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .Y(n12469));
  XOR2X1  g09200(.A(n12469), .B(n12464), .Y(n12470));
  XOR2X1  g09201(.A(n12436), .B(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .Y(n12471));
  INVX1   g09202(.A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .Y(n12472));
  AOI22X1 g09203(.A0(n10895), .A1(P2_REIP_REG_30__SCAN_IN), .B0(P2_EAX_REG_30__SCAN_IN), .B1(n10896), .Y(n12473));
  OAI21X1 g09204(.A0(n10892), .A1(n12472), .B0(n12473), .Y(n12474));
  NAND2X1 g09205(.A(n12440), .B(n12438), .Y(n12475));
  XOR2X1  g09206(.A(n12475), .B(n12474), .Y(n12476));
  NAND4X1 g09207(.A(n12405), .B(n12360), .C(n12356), .D(n12447), .Y(n12477));
  AOI22X1 g09208(.A0(P2_REIP_REG_30__SCAN_IN), .A1(n9488), .B0(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .B1(P2_STATE2_REG_1__SCAN_IN), .Y(n12478));
  INVX1   g09209(.A(n12478), .Y(n12479));
  AOI21X1 g09210(.A0(n9573), .A1(P2_EBX_REG_30__SCAN_IN), .B0(n12479), .Y(n12480));
  OAI21X1 g09211(.A0(n9542), .A1(n12472), .B0(n12480), .Y(n12481));
  XOR2X1  g09212(.A(n12481), .B(n12477), .Y(n12482));
  NOR2X1  g09213(.A(n12482), .B(n11042), .Y(n12483));
  NOR3X1  g09214(.A(n12412), .B(n12435), .C(n12383), .Y(n12484));
  XOR2X1  g09215(.A(n12484), .B(n12472), .Y(n12485));
  NOR2X1  g09216(.A(n12485), .B(n11494), .Y(n12486));
  NOR4X1  g09217(.A(n12435), .B(n12383), .C(n12344), .D(n12372), .Y(n12487));
  XOR2X1  g09218(.A(n12487), .B(n12472), .Y(n12488));
  AOI22X1 g09219(.A0(n10979), .A1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B0(P2_REIP_REG_30__SCAN_IN), .B1(n10965), .Y(n12489));
  OAI21X1 g09220(.A0(n12488), .A1(n10989), .B0(n12489), .Y(n12490));
  NOR3X1  g09221(.A(n12490), .B(n12486), .C(n12483), .Y(n12491));
  OAI21X1 g09222(.A0(n12476), .A1(n10986), .B0(n12491), .Y(n12492));
  AOI21X1 g09223(.A0(n12471), .A1(n12547), .B0(n12492), .Y(n12493));
  OAI21X1 g09224(.A0(n12470), .A1(n11386), .B0(n12493), .Y(P2_U3016));
  NAND2X1 g09225(.A(n12466), .B(n12465), .Y(n12495));
  AOI21X1 g09226(.A0(n9468), .A1(P2_EBX_REG_31__SCAN_IN), .B0(n11477), .Y(n12496));
  XOR2X1  g09227(.A(n12496), .B(n12495), .Y(n12497));
  NOR2X1  g09228(.A(n12497), .B(n11002), .Y(n12498));
  XOR2X1  g09229(.A(n12498), .B(n9163), .Y(n12499));
  NOR2X1  g09230(.A(n12468), .B(n12472), .Y(n12500));
  INVX1   g09231(.A(n12500), .Y(n12501));
  NAND4X1 g09232(.A(n12499), .B(n12463), .C(n12462), .D(n12501), .Y(n12502));
  NAND3X1 g09233(.A(n12462), .B(n12423), .C(n12422), .Y(n12503));
  NOR2X1  g09234(.A(n12431), .B(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .Y(n12504));
  AOI21X1 g09235(.A0(n12467), .A1(n11007), .B0(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .Y(n12505));
  NOR3X1  g09236(.A(n12505), .B(n12499), .C(n12504), .Y(n12506));
  OAI21X1 g09237(.A0(n12503), .A1(n12420), .B0(n12506), .Y(n12507));
  NOR2X1  g09238(.A(n12501), .B(n12499), .Y(n12508));
  AOI21X1 g09239(.A0(n12505), .A1(n12499), .B0(n12508), .Y(n12509));
  NAND3X1 g09240(.A(n12509), .B(n12507), .C(n12502), .Y(n12510));
  NOR4X1  g09241(.A(n12318), .B(n12472), .C(n12435), .D(n12391), .Y(n12511));
  OAI21X1 g09242(.A0(n11556), .A1(n11553), .B0(n12511), .Y(n12512));
  XOR2X1  g09243(.A(n12512), .B(n9163), .Y(n12513));
  AOI22X1 g09244(.A0(n10895), .A1(P2_REIP_REG_31__SCAN_IN), .B0(P2_EAX_REG_31__SCAN_IN), .B1(n10896), .Y(n12514));
  OAI21X1 g09245(.A0(n10892), .A1(n9163), .B0(n12514), .Y(n12515));
  NAND4X1 g09246(.A(n12474), .B(n12440), .C(n12438), .D(n12515), .Y(n12516));
  INVX1   g09247(.A(n12474), .Y(n12517));
  NOR2X1  g09248(.A(n12475), .B(n12517), .Y(n12518));
  OAI21X1 g09249(.A0(n12518), .A1(n12515), .B0(n12516), .Y(n12519));
  INVX1   g09250(.A(n12481), .Y(n12520));
  NOR2X1  g09251(.A(n12520), .B(n12477), .Y(n12521));
  INVX1   g09252(.A(P2_EBX_REG_31__SCAN_IN), .Y(n12522));
  AOI22X1 g09253(.A0(P2_REIP_REG_31__SCAN_IN), .A1(n9488), .B0(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B1(P2_STATE2_REG_1__SCAN_IN), .Y(n12523));
  OAI21X1 g09254(.A0(n9485), .A1(n12522), .B0(n12523), .Y(n12524));
  AOI21X1 g09255(.A0(n9483), .A1(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B0(n12524), .Y(n12525));
  XOR2X1  g09256(.A(n12525), .B(n12521), .Y(n12526));
  NOR2X1  g09257(.A(n12526), .B(n11042), .Y(n12527));
  NOR4X1  g09258(.A(n12472), .B(n12435), .C(n12383), .D(n12412), .Y(n12528));
  XOR2X1  g09259(.A(n12528), .B(n9163), .Y(n12529));
  NOR2X1  g09260(.A(n12529), .B(n11494), .Y(n12530));
  NAND2X1 g09261(.A(n12487), .B(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .Y(n12531));
  XOR2X1  g09262(.A(n12531), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .Y(n12532));
  AOI22X1 g09263(.A0(n10979), .A1(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B0(P2_REIP_REG_31__SCAN_IN), .B1(n10965), .Y(n12533));
  OAI21X1 g09264(.A0(n12532), .A1(n10989), .B0(n12533), .Y(n12534));
  NOR3X1  g09265(.A(n12534), .B(n12530), .C(n12527), .Y(n12535));
  OAI21X1 g09266(.A0(n12519), .A1(n10986), .B0(n12535), .Y(n12536));
  AOI21X1 g09267(.A0(n12513), .A1(n12547), .B0(n12536), .Y(n12537));
  OAI21X1 g09268(.A0(n12510), .A1(n11386), .B0(n12537), .Y(P2_U3015));
  NAND2X1 g09269(.A(n9724), .B(n8915), .Y(n12539));
  OAI22X1 g09270(.A0(n10958), .A1(P2_STATE2_REG_0__SCAN_IN), .B0(n9406), .B1(n12539), .Y(n12540));
  INVX1   g09271(.A(n12540), .Y(n12541));
  NOR2X1  g09272(.A(P2_STATEBS16_REG_SCAN_IN), .B(n9205), .Y(n12542));
  OAI21X1 g09273(.A0(n9765), .A1(n12542), .B0(n12540), .Y(n12543));
  INVX1   g09274(.A(n12543), .Y(n12544));
  OAI21X1 g09275(.A0(n12544), .A1(n12541), .B0(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .Y(n12545));
  NOR3X1  g09276(.A(n12541), .B(n9710), .C(n9205), .Y(n12546));
  NOR2X1  g09277(.A(n12541), .B(n9278), .Y(n12547));
  AOI22X1 g09278(.A0(n12546), .A1(n9752), .B0(n11037), .B1(n12547), .Y(n12548));
  NOR3X1  g09279(.A(n12541), .B(n9022), .C(n8720), .Y(n12549));
  AOI22X1 g09280(.A0(n12549), .A1(n11034), .B0(P2_REIP_REG_0__SCAN_IN), .B1(n10965), .Y(n12551));
  NAND3X1 g09281(.A(n12551), .B(n12548), .C(n12545), .Y(P2_U3014));
  NOR2X1  g09282(.A(n12540), .B(n9574), .Y(n12553));
  AOI21X1 g09283(.A0(n12544), .A1(n9574), .B0(n12553), .Y(n12554));
  AOI22X1 g09284(.A0(n12546), .A1(n9751), .B0(n11088), .B1(n12547), .Y(n12555));
  OAI21X1 g09285(.A0(n11079), .A1(n11075), .B0(n12549), .Y(n12556));
  NAND3X1 g09286(.A(n12540), .B(n9729), .C(P2_REIP_REG_1__SCAN_IN), .Y(n12557));
  NAND4X1 g09287(.A(n12556), .B(n12555), .C(n12554), .D(n12557), .Y(P2_U3013));
  XOR2X1  g09288(.A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .Y(n12559));
  AOI22X1 g09289(.A0(n12544), .A1(n12559), .B0(n12541), .B1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .Y(n12560));
  AOI22X1 g09290(.A0(n12546), .A1(n9794), .B0(n11133), .B1(n12547), .Y(n12561));
  AOI22X1 g09291(.A0(n12549), .A1(n11128), .B0(P2_REIP_REG_2__SCAN_IN), .B1(n10965), .Y(n12562));
  NAND3X1 g09292(.A(n12562), .B(n12561), .C(n12560), .Y(P2_U3012));
  NAND2X1 g09293(.A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .Y(n12564));
  XOR2X1  g09294(.A(n12564), .B(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .Y(n12565));
  INVX1   g09295(.A(n12565), .Y(n12566));
  AOI22X1 g09296(.A0(n12544), .A1(n12566), .B0(n12541), .B1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .Y(n12567));
  AOI22X1 g09297(.A0(n12546), .A1(n9815), .B0(n11183), .B1(n12547), .Y(n12568));
  AOI22X1 g09298(.A0(n12549), .A1(n11177), .B0(P2_REIP_REG_3__SCAN_IN), .B1(n10965), .Y(n12569));
  NAND3X1 g09299(.A(n12569), .B(n12568), .C(n12567), .Y(P2_U3011));
  NAND2X1 g09300(.A(n12549), .B(n11236), .Y(n12571));
  INVX1   g09301(.A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .Y(n12572));
  NAND3X1 g09302(.A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .C(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .Y(n12573));
  XOR2X1  g09303(.A(n12573), .B(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .Y(n12574));
  OAI22X1 g09304(.A0(n12543), .A1(n12574), .B0(n12540), .B1(n12572), .Y(n12575));
  NOR4X1  g09305(.A(n8602), .B(P2_STATE2_REG_1__SCAN_IN), .C(P2_STATE2_REG_2__SCAN_IN), .D(n12541), .Y(n12576));
  INVX1   g09306(.A(n12546), .Y(n12577));
  INVX1   g09307(.A(n12547), .Y(n12578));
  OAI22X1 g09308(.A0(n12577), .A1(n11251), .B0(n11242), .B1(n12578), .Y(n12579));
  NOR3X1  g09309(.A(n12579), .B(n12576), .C(n12575), .Y(n12580));
  NAND2X1 g09310(.A(n12580), .B(n12571), .Y(P2_U3010));
  NAND2X1 g09311(.A(n12549), .B(n11303), .Y(n12582));
  NAND2X1 g09312(.A(n12547), .B(n11310), .Y(n12583));
  XOR2X1  g09313(.A(n9180), .B(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .Y(n12584));
  INVX1   g09314(.A(n12584), .Y(n12585));
  AOI22X1 g09315(.A0(n12544), .A1(n12585), .B0(n12541), .B1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .Y(n12586));
  NOR4X1  g09316(.A(n11315), .B(n9710), .C(n9205), .D(n12541), .Y(n12587));
  AOI21X1 g09317(.A0(n10965), .A1(P2_REIP_REG_5__SCAN_IN), .B0(n12587), .Y(n12588));
  NAND4X1 g09318(.A(n12586), .B(n12583), .C(n12582), .D(n12588), .Y(P2_U3009));
  INVX1   g09319(.A(n12549), .Y(n12590));
  NOR2X1  g09320(.A(n9180), .B(n9177), .Y(n12591));
  XOR2X1  g09321(.A(n12591), .B(n9178), .Y(n12592));
  INVX1   g09322(.A(n12592), .Y(n12593));
  AOI22X1 g09323(.A0(n12544), .A1(n12593), .B0(n12541), .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .Y(n12594));
  INVX1   g09324(.A(n11381), .Y(n12595));
  AOI22X1 g09325(.A0(n12546), .A1(n12595), .B0(P2_REIP_REG_6__SCAN_IN), .B1(n10965), .Y(n12596));
  NAND2X1 g09326(.A(n12596), .B(n12594), .Y(n12597));
  AOI21X1 g09327(.A0(n12547), .A1(n11376), .B0(n12597), .Y(n12598));
  OAI21X1 g09328(.A0(n12590), .A1(n11370), .B0(n12598), .Y(P2_U3008));
  NOR3X1  g09329(.A(n9180), .B(n9178), .C(n9177), .Y(n12600));
  XOR2X1  g09330(.A(n12600), .B(n9179), .Y(n12601));
  INVX1   g09331(.A(n12601), .Y(n12602));
  AOI22X1 g09332(.A0(n12544), .A1(n12602), .B0(n12541), .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .Y(n12603));
  AOI22X1 g09333(.A0(n12546), .A1(n11430), .B0(P2_REIP_REG_7__SCAN_IN), .B1(n10965), .Y(n12604));
  NAND2X1 g09334(.A(n12604), .B(n12603), .Y(n12605));
  AOI21X1 g09335(.A0(n12547), .A1(n11424), .B0(n12605), .Y(n12606));
  OAI21X1 g09336(.A0(n12590), .A1(n11418), .B0(n12606), .Y(P2_U3007));
  NAND2X1 g09337(.A(n12549), .B(n11484), .Y(n12609));
  XOR2X1  g09338(.A(n9181), .B(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .Y(n12610));
  AOI22X1 g09339(.A0(n12544), .A1(n12610), .B0(n12541), .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .Y(n12611));
  INVX1   g09340(.A(n11491), .Y(n12612));
  AOI22X1 g09341(.A0(n12546), .A1(n12612), .B0(P2_REIP_REG_8__SCAN_IN), .B1(n10965), .Y(n12613));
  NAND4X1 g09342(.A(n12611), .B(n12609), .C(n11462), .D(n12613), .Y(P2_U3006));
  NAND2X1 g09343(.A(n9181), .B(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .Y(n12615));
  XOR2X1  g09344(.A(n12615), .B(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .Y(n12616));
  INVX1   g09345(.A(n12616), .Y(n12617));
  AOI22X1 g09346(.A0(n12544), .A1(n12617), .B0(n12541), .B1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .Y(n12618));
  AOI22X1 g09347(.A0(n12546), .A1(n11565), .B0(P2_REIP_REG_9__SCAN_IN), .B1(n10965), .Y(n12619));
  NAND2X1 g09348(.A(n12619), .B(n12618), .Y(n12620));
  AOI21X1 g09349(.A0(n12547), .A1(n11558), .B0(n12620), .Y(n12621));
  OAI21X1 g09350(.A0(n12590), .A1(n11550), .B0(n12621), .Y(P2_U3005));
  NAND2X1 g09351(.A(n12549), .B(n11611), .Y(n12624));
  NAND3X1 g09352(.A(n9181), .B(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .C(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .Y(n12625));
  XOR2X1  g09353(.A(n12625), .B(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .Y(n12626));
  INVX1   g09354(.A(n12626), .Y(n12627));
  AOI22X1 g09355(.A0(n12544), .A1(n12627), .B0(n12541), .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .Y(n12628));
  INVX1   g09356(.A(n11618), .Y(n12629));
  AOI22X1 g09357(.A0(n12546), .A1(n12629), .B0(P2_REIP_REG_10__SCAN_IN), .B1(n10965), .Y(n12630));
  NAND4X1 g09358(.A(n12628), .B(n12624), .C(n11598), .D(n12630), .Y(P2_U3004));
  XOR2X1  g09359(.A(n9182), .B(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .Y(n12632));
  INVX1   g09360(.A(n12632), .Y(n12633));
  AOI22X1 g09361(.A0(n12544), .A1(n12633), .B0(n12541), .B1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .Y(n12634));
  AOI22X1 g09362(.A0(n12546), .A1(n11666), .B0(P2_REIP_REG_11__SCAN_IN), .B1(n10965), .Y(n12635));
  NAND2X1 g09363(.A(n12635), .B(n12634), .Y(n12636));
  AOI21X1 g09364(.A0(n12547), .A1(n11659), .B0(n12636), .Y(n12637));
  OAI21X1 g09365(.A0(n12590), .A1(n11655), .B0(n12637), .Y(P2_U3003));
  NOR2X1  g09366(.A(n9182), .B(n9174), .Y(n12639));
  XOR2X1  g09367(.A(n12639), .B(n9175), .Y(n12640));
  INVX1   g09368(.A(n12640), .Y(n12641));
  AOI22X1 g09369(.A0(n12544), .A1(n12641), .B0(n12541), .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .Y(n12642));
  AOI22X1 g09370(.A0(n12546), .A1(n11718), .B0(P2_REIP_REG_12__SCAN_IN), .B1(n10965), .Y(n12643));
  NAND2X1 g09371(.A(n12643), .B(n12642), .Y(n12644));
  AOI21X1 g09372(.A0(n12547), .A1(n11711), .B0(n12644), .Y(n12645));
  OAI21X1 g09373(.A0(n12590), .A1(n11710), .B0(n12645), .Y(P2_U3002));
  NOR3X1  g09374(.A(n9182), .B(n9175), .C(n9174), .Y(n12647));
  XOR2X1  g09375(.A(n12647), .B(n9176), .Y(n12648));
  INVX1   g09376(.A(n12648), .Y(n12649));
  AOI22X1 g09377(.A0(n12544), .A1(n12649), .B0(n12541), .B1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .Y(n12650));
  AOI22X1 g09378(.A0(n12546), .A1(n11773), .B0(P2_REIP_REG_13__SCAN_IN), .B1(n10965), .Y(n12651));
  NAND2X1 g09379(.A(n12651), .B(n12650), .Y(n12652));
  AOI21X1 g09380(.A0(n12547), .A1(n11767), .B0(n12652), .Y(n12653));
  OAI21X1 g09381(.A0(n12590), .A1(n11760), .B0(n12653), .Y(P2_U3001));
  XOR2X1  g09382(.A(n9183), .B(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .Y(n12655));
  AOI22X1 g09383(.A0(n12544), .A1(n12655), .B0(n12541), .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .Y(n12656));
  AOI22X1 g09384(.A0(n12546), .A1(n11825), .B0(P2_REIP_REG_14__SCAN_IN), .B1(n10965), .Y(n12657));
  NAND2X1 g09385(.A(n12657), .B(n12656), .Y(n12658));
  AOI21X1 g09386(.A0(n12547), .A1(n11818), .B0(n12658), .Y(n12659));
  OAI21X1 g09387(.A0(n12590), .A1(n11815), .B0(n12659), .Y(P2_U3000));
  NAND2X1 g09388(.A(n9183), .B(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .Y(n12661));
  XOR2X1  g09389(.A(n12661), .B(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .Y(n12662));
  INVX1   g09390(.A(n12662), .Y(n12663));
  AOI22X1 g09391(.A0(n12544), .A1(n12663), .B0(n12541), .B1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .Y(n12664));
  AOI22X1 g09392(.A0(n12546), .A1(n11874), .B0(P2_REIP_REG_15__SCAN_IN), .B1(n10965), .Y(n12665));
  NAND2X1 g09393(.A(n12665), .B(n12664), .Y(n12666));
  AOI21X1 g09394(.A0(n12547), .A1(n11868), .B0(n12666), .Y(n12667));
  OAI21X1 g09395(.A0(n12590), .A1(n11867), .B0(n12667), .Y(P2_U2999));
  NAND3X1 g09396(.A(n9183), .B(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .C(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .Y(n12669));
  XOR2X1  g09397(.A(n12669), .B(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .Y(n12670));
  INVX1   g09398(.A(n12670), .Y(n12671));
  AOI22X1 g09399(.A0(n12544), .A1(n12671), .B0(n12541), .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .Y(n12672));
  AOI22X1 g09400(.A0(n12546), .A1(n11931), .B0(P2_REIP_REG_16__SCAN_IN), .B1(n10965), .Y(n12673));
  NAND2X1 g09401(.A(n12673), .B(n12672), .Y(n12674));
  AOI21X1 g09402(.A0(n12547), .A1(n11924), .B0(n12674), .Y(n12675));
  OAI21X1 g09403(.A0(n12590), .A1(n11918), .B0(n12675), .Y(P2_U2998));
  XOR2X1  g09404(.A(n9184), .B(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .Y(n12677));
  INVX1   g09405(.A(n12677), .Y(n12678));
  AOI22X1 g09406(.A0(n12544), .A1(n12678), .B0(n12541), .B1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .Y(n12679));
  AOI22X1 g09407(.A0(n12546), .A1(n11969), .B0(P2_REIP_REG_17__SCAN_IN), .B1(n10965), .Y(n12680));
  NAND2X1 g09408(.A(n12680), .B(n12679), .Y(n12681));
  AOI21X1 g09409(.A0(n12547), .A1(n11962), .B0(n12681), .Y(n12682));
  OAI21X1 g09410(.A0(n12590), .A1(n11961), .B0(n12682), .Y(P2_U2997));
  NOR2X1  g09411(.A(n9184), .B(n9171), .Y(n12684));
  XOR2X1  g09412(.A(n12684), .B(n9172), .Y(n12685));
  INVX1   g09413(.A(n12685), .Y(n12686));
  AOI22X1 g09414(.A0(n12544), .A1(n12686), .B0(n12541), .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .Y(n12687));
  AOI22X1 g09415(.A0(n12546), .A1(n12007), .B0(P2_REIP_REG_18__SCAN_IN), .B1(n10965), .Y(n12688));
  NAND2X1 g09416(.A(n12688), .B(n12687), .Y(n12689));
  AOI21X1 g09417(.A0(n12547), .A1(n12001), .B0(n12689), .Y(n12690));
  OAI21X1 g09418(.A0(n12590), .A1(n11999), .B0(n12690), .Y(P2_U2996));
  NOR3X1  g09419(.A(n9184), .B(n9172), .C(n9171), .Y(n12692));
  XOR2X1  g09420(.A(n12692), .B(n9173), .Y(n12693));
  INVX1   g09421(.A(n12693), .Y(n12694));
  AOI22X1 g09422(.A0(n12544), .A1(n12694), .B0(n12541), .B1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .Y(n12695));
  AOI22X1 g09423(.A0(n12546), .A1(n12048), .B0(P2_REIP_REG_19__SCAN_IN), .B1(n10965), .Y(n12696));
  NAND2X1 g09424(.A(n12696), .B(n12695), .Y(n12697));
  AOI21X1 g09425(.A0(n12547), .A1(n12041), .B0(n12697), .Y(n12698));
  OAI21X1 g09426(.A0(n12590), .A1(n12036), .B0(n12698), .Y(P2_U2995));
  XOR2X1  g09427(.A(n9185), .B(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .Y(n12700));
  AOI22X1 g09428(.A0(n12544), .A1(n12700), .B0(n12541), .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .Y(n12701));
  AOI22X1 g09429(.A0(n12546), .A1(n12088), .B0(P2_REIP_REG_20__SCAN_IN), .B1(n10965), .Y(n12702));
  NAND2X1 g09430(.A(n12702), .B(n12701), .Y(n12703));
  AOI21X1 g09431(.A0(n12547), .A1(n12081), .B0(n12703), .Y(n12704));
  OAI21X1 g09432(.A0(n12590), .A1(n12076), .B0(n12704), .Y(P2_U2994));
  NAND2X1 g09433(.A(n9185), .B(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .Y(n12706));
  XOR2X1  g09434(.A(n12706), .B(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .Y(n12707));
  INVX1   g09435(.A(n12707), .Y(n12708));
  AOI22X1 g09436(.A0(n12544), .A1(n12708), .B0(n12541), .B1(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .Y(n12709));
  AOI22X1 g09437(.A0(n12546), .A1(n12126), .B0(P2_REIP_REG_21__SCAN_IN), .B1(n10965), .Y(n12710));
  NAND2X1 g09438(.A(n12710), .B(n12709), .Y(n12711));
  AOI21X1 g09439(.A0(n12547), .A1(n12119), .B0(n12711), .Y(n12712));
  OAI21X1 g09440(.A0(n12590), .A1(n12118), .B0(n12712), .Y(P2_U2993));
  NAND3X1 g09441(.A(n9185), .B(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .C(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .Y(n12714));
  XOR2X1  g09442(.A(n12714), .B(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .Y(n12715));
  INVX1   g09443(.A(n12715), .Y(n12716));
  AOI22X1 g09444(.A0(n12544), .A1(n12716), .B0(n12541), .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .Y(n12717));
  AOI22X1 g09445(.A0(n12546), .A1(n12165), .B0(P2_REIP_REG_22__SCAN_IN), .B1(n10965), .Y(n12718));
  NAND2X1 g09446(.A(n12718), .B(n12717), .Y(n12719));
  AOI21X1 g09447(.A0(n12547), .A1(n12158), .B0(n12719), .Y(n12720));
  OAI21X1 g09448(.A0(n12590), .A1(n12154), .B0(n12720), .Y(P2_U2992));
  XOR2X1  g09449(.A(n9186), .B(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .Y(n12722));
  INVX1   g09450(.A(n12722), .Y(n12723));
  AOI22X1 g09451(.A0(n12544), .A1(n12723), .B0(n12541), .B1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .Y(n12724));
  AOI22X1 g09452(.A0(n12546), .A1(n12211), .B0(P2_REIP_REG_23__SCAN_IN), .B1(n10965), .Y(n12725));
  NAND2X1 g09453(.A(n12725), .B(n12724), .Y(n12726));
  AOI21X1 g09454(.A0(n12547), .A1(n12204), .B0(n12726), .Y(n12727));
  OAI21X1 g09455(.A0(n12590), .A1(n12198), .B0(n12727), .Y(P2_U2991));
  NOR2X1  g09456(.A(n9186), .B(n9168), .Y(n12729));
  XOR2X1  g09457(.A(n12729), .B(n9169), .Y(n12730));
  INVX1   g09458(.A(n12730), .Y(n12731));
  AOI22X1 g09459(.A0(n12544), .A1(n12731), .B0(n12541), .B1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .Y(n12732));
  AOI22X1 g09460(.A0(n12546), .A1(n12248), .B0(P2_REIP_REG_24__SCAN_IN), .B1(n10965), .Y(n12733));
  NAND2X1 g09461(.A(n12733), .B(n12732), .Y(n12734));
  AOI21X1 g09462(.A0(n12547), .A1(n12241), .B0(n12734), .Y(n12735));
  OAI21X1 g09463(.A0(n12590), .A1(n12240), .B0(n12735), .Y(P2_U2990));
  NOR3X1  g09464(.A(n9186), .B(n9169), .C(n9168), .Y(n12737));
  XOR2X1  g09465(.A(n12737), .B(n9170), .Y(n12738));
  INVX1   g09466(.A(n12738), .Y(n12739));
  AOI22X1 g09467(.A0(n12544), .A1(n12739), .B0(n12541), .B1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .Y(n12740));
  AOI22X1 g09468(.A0(n12546), .A1(n12287), .B0(P2_REIP_REG_25__SCAN_IN), .B1(n10965), .Y(n12741));
  NAND2X1 g09469(.A(n12741), .B(n12740), .Y(n12742));
  AOI21X1 g09470(.A0(n12547), .A1(n12281), .B0(n12742), .Y(n12743));
  OAI21X1 g09471(.A0(n12590), .A1(n12279), .B0(n12743), .Y(P2_U2989));
  NAND2X1 g09472(.A(n12549), .B(n12313), .Y(n12745));
  NAND2X1 g09473(.A(n12546), .B(n12327), .Y(n12746));
  NAND3X1 g09474(.A(n12540), .B(n9729), .C(P2_REIP_REG_26__SCAN_IN), .Y(n12747));
  XOR2X1  g09475(.A(n9187), .B(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .Y(n12748));
  AOI22X1 g09476(.A0(n12544), .A1(n12748), .B0(n12541), .B1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .Y(n12749));
  NAND3X1 g09477(.A(n12749), .B(n12747), .C(n12746), .Y(n12750));
  AOI21X1 g09478(.A0(n12547), .A1(n12320), .B0(n12750), .Y(n12751));
  NAND2X1 g09479(.A(n12751), .B(n12745), .Y(P2_U2988));
  NAND2X1 g09480(.A(n12549), .B(n12352), .Y(n12753));
  NAND2X1 g09481(.A(n12546), .B(n12361), .Y(n12755));
  INVX1   g09482(.A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .Y(n12756));
  NAND2X1 g09483(.A(n9187), .B(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .Y(n12757));
  XOR2X1  g09484(.A(n12757), .B(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .Y(n12758));
  OAI22X1 g09485(.A0(n12543), .A1(n12758), .B0(n12540), .B1(n12756), .Y(n12759));
  AOI21X1 g09486(.A0(n10965), .A1(P2_REIP_REG_27__SCAN_IN), .B0(n12759), .Y(n12760));
  NAND4X1 g09487(.A(n12755), .B(n12355), .C(n12753), .D(n12760), .Y(P2_U2987));
  INVX1   g09488(.A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .Y(n12762));
  NAND3X1 g09489(.A(n9187), .B(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .C(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .Y(n12763));
  XOR2X1  g09490(.A(n12763), .B(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .Y(n12764));
  OAI22X1 g09491(.A0(n12543), .A1(n12764), .B0(n12540), .B1(n12762), .Y(n12765));
  AOI21X1 g09492(.A0(n10965), .A1(P2_REIP_REG_28__SCAN_IN), .B0(n12765), .Y(n12766));
  OAI21X1 g09493(.A0(n12577), .A1(n12406), .B0(n12766), .Y(n12767));
  AOI21X1 g09494(.A0(n12547), .A1(n12393), .B0(n12767), .Y(n12768));
  OAI21X1 g09495(.A0(n12590), .A1(n12389), .B0(n12768), .Y(P2_U2986));
  XOR2X1  g09496(.A(n9188), .B(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .Y(n12770));
  OAI22X1 g09497(.A0(n12543), .A1(n12770), .B0(n12540), .B1(n9166), .Y(n12771));
  AOI21X1 g09498(.A0(n10965), .A1(P2_REIP_REG_29__SCAN_IN), .B0(n12771), .Y(n12772));
  OAI21X1 g09499(.A0(n12577), .A1(n12448), .B0(n12772), .Y(n12773));
  AOI21X1 g09500(.A0(n12547), .A1(n12437), .B0(n12773), .Y(n12774));
  OAI21X1 g09501(.A0(n12590), .A1(n12433), .B0(n12774), .Y(P2_U2985));
  NOR2X1  g09502(.A(n9188), .B(n9166), .Y(n12776));
  XOR2X1  g09503(.A(n12776), .B(n9167), .Y(n12777));
  OAI22X1 g09504(.A0(n12543), .A1(n12777), .B0(n12540), .B1(n9167), .Y(n12778));
  AOI21X1 g09505(.A0(n10965), .A1(P2_REIP_REG_30__SCAN_IN), .B0(n12778), .Y(n12779));
  OAI21X1 g09506(.A0(n12577), .A1(n12482), .B0(n12779), .Y(n12780));
  AOI21X1 g09507(.A0(n12547), .A1(n12471), .B0(n12780), .Y(n12781));
  OAI21X1 g09508(.A0(n12590), .A1(n12470), .B0(n12781), .Y(P2_U2984));
  OAI22X1 g09509(.A0(n12540), .A1(n9165), .B0(n9190), .B1(n12543), .Y(n12783));
  AOI21X1 g09510(.A0(n10965), .A1(P2_REIP_REG_31__SCAN_IN), .B0(n12783), .Y(n12784));
  OAI21X1 g09511(.A0(n12577), .A1(n12526), .B0(n12784), .Y(n12785));
  AOI21X1 g09512(.A0(n12547), .A1(n12513), .B0(n12785), .Y(n12786));
  OAI21X1 g09513(.A0(n12590), .A1(n12510), .B0(n12786), .Y(P2_U2983));
  INVX1   g09514(.A(BUF1_REG_15__SCAN_IN), .Y(n12788));
  NOR2X1  g09515(.A(n3086), .B(n12788), .Y(n12789));
  AOI21X1 g09516(.A0(n3086), .A1(BUF2_REG_15__SCAN_IN), .B0(n12789), .Y(n12790));
  NOR2X1  g09517(.A(n9487), .B(n9357), .Y(n12791));
  INVX1   g09518(.A(n12791), .Y(n12792));
  INVX1   g09519(.A(n9714), .Y(n12793));
  NOR2X1  g09520(.A(n9022), .B(n8620), .Y(n12794));
  NOR4X1  g09521(.A(n12793), .B(n12792), .C(n9262), .D(n12794), .Y(n12795));
  INVX1   g09522(.A(n12795), .Y(n12796));
  NOR2X1  g09523(.A(n12796), .B(n9022), .Y(n12797));
  INVX1   g09524(.A(n12797), .Y(n12798));
  NOR2X1  g09525(.A(n12796), .B(n8975), .Y(n12799));
  AOI22X1 g09526(.A0(n12796), .A1(P2_LWORD_REG_15__SCAN_IN), .B0(P2_EAX_REG_15__SCAN_IN), .B1(n12799), .Y(n12800));
  OAI21X1 g09527(.A0(n12798), .A1(n12790), .B0(n12800), .Y(P2_U2982));
  INVX1   g09528(.A(BUF1_REG_14__SCAN_IN), .Y(n12802));
  NOR2X1  g09529(.A(n3086), .B(n12802), .Y(n12803));
  AOI21X1 g09530(.A0(n3086), .A1(BUF2_REG_14__SCAN_IN), .B0(n12803), .Y(n12804));
  INVX1   g09531(.A(n12804), .Y(n12805));
  NAND3X1 g09532(.A(n12805), .B(n12795), .C(n8975), .Y(n12806));
  AOI22X1 g09533(.A0(n12796), .A1(P2_LWORD_REG_14__SCAN_IN), .B0(P2_EAX_REG_14__SCAN_IN), .B1(n12799), .Y(n12807));
  NAND2X1 g09534(.A(n12807), .B(n12806), .Y(P2_U2981));
  INVX1   g09535(.A(BUF1_REG_13__SCAN_IN), .Y(n12809));
  NOR2X1  g09536(.A(n3086), .B(n12809), .Y(n12810));
  AOI21X1 g09537(.A0(n3086), .A1(BUF2_REG_13__SCAN_IN), .B0(n12810), .Y(n12811));
  INVX1   g09538(.A(n12811), .Y(n12812));
  NAND3X1 g09539(.A(n12812), .B(n12795), .C(n8975), .Y(n12813));
  AOI22X1 g09540(.A0(n12796), .A1(P2_LWORD_REG_13__SCAN_IN), .B0(P2_EAX_REG_13__SCAN_IN), .B1(n12799), .Y(n12814));
  NAND2X1 g09541(.A(n12814), .B(n12813), .Y(P2_U2980));
  INVX1   g09542(.A(BUF1_REG_12__SCAN_IN), .Y(n12816));
  NAND2X1 g09543(.A(n3086), .B(BUF2_REG_12__SCAN_IN), .Y(n12817));
  OAI21X1 g09544(.A0(n3086), .A1(n12816), .B0(n12817), .Y(n12818));
  NAND3X1 g09545(.A(n12818), .B(n12795), .C(n8975), .Y(n12819));
  AOI22X1 g09546(.A0(n12796), .A1(P2_LWORD_REG_12__SCAN_IN), .B0(P2_EAX_REG_12__SCAN_IN), .B1(n12799), .Y(n12820));
  NAND2X1 g09547(.A(n12820), .B(n12819), .Y(P2_U2979));
  INVX1   g09548(.A(BUF1_REG_11__SCAN_IN), .Y(n12822));
  NAND2X1 g09549(.A(n3086), .B(BUF2_REG_11__SCAN_IN), .Y(n12823));
  OAI21X1 g09550(.A0(n3086), .A1(n12822), .B0(n12823), .Y(n12824));
  NAND3X1 g09551(.A(n12824), .B(n12795), .C(n8975), .Y(n12825));
  AOI22X1 g09552(.A0(n12796), .A1(P2_LWORD_REG_11__SCAN_IN), .B0(P2_EAX_REG_11__SCAN_IN), .B1(n12799), .Y(n12826));
  NAND2X1 g09553(.A(n12826), .B(n12825), .Y(P2_U2978));
  INVX1   g09554(.A(BUF1_REG_10__SCAN_IN), .Y(n12828));
  NAND2X1 g09555(.A(n3086), .B(BUF2_REG_10__SCAN_IN), .Y(n12829));
  OAI21X1 g09556(.A0(n3086), .A1(n12828), .B0(n12829), .Y(n12830));
  NAND3X1 g09557(.A(n12830), .B(n12795), .C(n8975), .Y(n12831));
  AOI22X1 g09558(.A0(n12796), .A1(P2_LWORD_REG_10__SCAN_IN), .B0(P2_EAX_REG_10__SCAN_IN), .B1(n12799), .Y(n12832));
  NAND2X1 g09559(.A(n12832), .B(n12831), .Y(P2_U2977));
  INVX1   g09560(.A(BUF1_REG_9__SCAN_IN), .Y(n12834));
  NAND2X1 g09561(.A(n3086), .B(BUF2_REG_9__SCAN_IN), .Y(n12835));
  OAI21X1 g09562(.A0(n3086), .A1(n12834), .B0(n12835), .Y(n12836));
  NAND3X1 g09563(.A(n12836), .B(n12795), .C(n8975), .Y(n12837));
  AOI22X1 g09564(.A0(n12796), .A1(P2_LWORD_REG_9__SCAN_IN), .B0(P2_EAX_REG_9__SCAN_IN), .B1(n12799), .Y(n12838));
  NAND2X1 g09565(.A(n12838), .B(n12837), .Y(P2_U2976));
  INVX1   g09566(.A(BUF1_REG_8__SCAN_IN), .Y(n12840));
  NAND2X1 g09567(.A(n3086), .B(BUF2_REG_8__SCAN_IN), .Y(n12841));
  OAI21X1 g09568(.A0(n3086), .A1(n12840), .B0(n12841), .Y(n12842));
  NAND3X1 g09569(.A(n12842), .B(n12795), .C(n8975), .Y(n12843));
  AOI22X1 g09570(.A0(n12796), .A1(P2_LWORD_REG_8__SCAN_IN), .B0(P2_EAX_REG_8__SCAN_IN), .B1(n12799), .Y(n12844));
  NAND2X1 g09571(.A(n12844), .B(n12843), .Y(P2_U2975));
  AOI22X1 g09572(.A0(n12796), .A1(P2_LWORD_REG_7__SCAN_IN), .B0(P2_EAX_REG_7__SCAN_IN), .B1(n12799), .Y(n12846));
  OAI21X1 g09573(.A0(n12798), .A1(n9743), .B0(n12846), .Y(P2_U2974));
  AOI22X1 g09574(.A0(n12796), .A1(P2_LWORD_REG_6__SCAN_IN), .B0(P2_EAX_REG_6__SCAN_IN), .B1(n12799), .Y(n12848));
  OAI21X1 g09575(.A0(n12798), .A1(n9860), .B0(n12848), .Y(P2_U2973));
  AOI22X1 g09576(.A0(n12796), .A1(P2_LWORD_REG_5__SCAN_IN), .B0(P2_EAX_REG_5__SCAN_IN), .B1(n12799), .Y(n12850));
  OAI21X1 g09577(.A0(n12798), .A1(n9879), .B0(n12850), .Y(P2_U2972));
  AOI22X1 g09578(.A0(n12796), .A1(P2_LWORD_REG_4__SCAN_IN), .B0(P2_EAX_REG_4__SCAN_IN), .B1(n12799), .Y(n12852));
  OAI21X1 g09579(.A0(n12798), .A1(n9898), .B0(n12852), .Y(P2_U2971));
  AOI22X1 g09580(.A0(n12796), .A1(P2_LWORD_REG_3__SCAN_IN), .B0(P2_EAX_REG_3__SCAN_IN), .B1(n12799), .Y(n12854));
  OAI21X1 g09581(.A0(n12798), .A1(n9917), .B0(n12854), .Y(P2_U2970));
  AOI22X1 g09582(.A0(n12796), .A1(P2_LWORD_REG_2__SCAN_IN), .B0(P2_EAX_REG_2__SCAN_IN), .B1(n12799), .Y(n12856));
  OAI21X1 g09583(.A0(n12798), .A1(n9936), .B0(n12856), .Y(P2_U2969));
  AOI22X1 g09584(.A0(n12796), .A1(P2_LWORD_REG_1__SCAN_IN), .B0(P2_EAX_REG_1__SCAN_IN), .B1(n12799), .Y(n12858));
  OAI21X1 g09585(.A0(n12798), .A1(n9955), .B0(n12858), .Y(P2_U2968));
  AOI22X1 g09586(.A0(n12796), .A1(P2_LWORD_REG_0__SCAN_IN), .B0(P2_EAX_REG_0__SCAN_IN), .B1(n12799), .Y(n12860));
  OAI21X1 g09587(.A0(n12798), .A1(n9974), .B0(n12860), .Y(P2_U2967));
  AOI22X1 g09588(.A0(n12796), .A1(P2_UWORD_REG_14__SCAN_IN), .B0(P2_EAX_REG_30__SCAN_IN), .B1(n12799), .Y(n12862));
  NAND2X1 g09589(.A(n12862), .B(n12806), .Y(P2_U2966));
  AOI22X1 g09590(.A0(n12796), .A1(P2_UWORD_REG_13__SCAN_IN), .B0(P2_EAX_REG_29__SCAN_IN), .B1(n12799), .Y(n12864));
  NAND2X1 g09591(.A(n12864), .B(n12813), .Y(P2_U2965));
  AOI22X1 g09592(.A0(n12796), .A1(P2_UWORD_REG_12__SCAN_IN), .B0(P2_EAX_REG_28__SCAN_IN), .B1(n12799), .Y(n12866));
  NAND2X1 g09593(.A(n12866), .B(n12819), .Y(P2_U2964));
  AOI22X1 g09594(.A0(n12796), .A1(P2_UWORD_REG_11__SCAN_IN), .B0(P2_EAX_REG_27__SCAN_IN), .B1(n12799), .Y(n12868));
  NAND2X1 g09595(.A(n12868), .B(n12825), .Y(P2_U2963));
  AOI22X1 g09596(.A0(n12796), .A1(P2_UWORD_REG_10__SCAN_IN), .B0(P2_EAX_REG_26__SCAN_IN), .B1(n12799), .Y(n12870));
  NAND2X1 g09597(.A(n12870), .B(n12831), .Y(P2_U2962));
  AOI22X1 g09598(.A0(n12796), .A1(P2_UWORD_REG_9__SCAN_IN), .B0(P2_EAX_REG_25__SCAN_IN), .B1(n12799), .Y(n12872));
  NAND2X1 g09599(.A(n12872), .B(n12837), .Y(P2_U2961));
  AOI22X1 g09600(.A0(n12796), .A1(P2_UWORD_REG_8__SCAN_IN), .B0(P2_EAX_REG_24__SCAN_IN), .B1(n12799), .Y(n12874));
  NAND2X1 g09601(.A(n12874), .B(n12843), .Y(P2_U2960));
  AOI22X1 g09602(.A0(n12796), .A1(P2_UWORD_REG_7__SCAN_IN), .B0(P2_EAX_REG_23__SCAN_IN), .B1(n12799), .Y(n12876));
  OAI21X1 g09603(.A0(n12798), .A1(n9743), .B0(n12876), .Y(P2_U2959));
  AOI22X1 g09604(.A0(n12796), .A1(P2_UWORD_REG_6__SCAN_IN), .B0(P2_EAX_REG_22__SCAN_IN), .B1(n12799), .Y(n12878));
  OAI21X1 g09605(.A0(n12798), .A1(n9860), .B0(n12878), .Y(P2_U2958));
  AOI22X1 g09606(.A0(n12796), .A1(P2_UWORD_REG_5__SCAN_IN), .B0(P2_EAX_REG_21__SCAN_IN), .B1(n12799), .Y(n12880));
  OAI21X1 g09607(.A0(n12798), .A1(n9879), .B0(n12880), .Y(P2_U2957));
  AOI22X1 g09608(.A0(n12796), .A1(P2_UWORD_REG_4__SCAN_IN), .B0(P2_EAX_REG_20__SCAN_IN), .B1(n12799), .Y(n12882));
  OAI21X1 g09609(.A0(n12798), .A1(n9898), .B0(n12882), .Y(P2_U2956));
  AOI22X1 g09610(.A0(n12796), .A1(P2_UWORD_REG_3__SCAN_IN), .B0(P2_EAX_REG_19__SCAN_IN), .B1(n12799), .Y(n12884));
  OAI21X1 g09611(.A0(n12798), .A1(n9917), .B0(n12884), .Y(P2_U2955));
  AOI22X1 g09612(.A0(n12796), .A1(P2_UWORD_REG_2__SCAN_IN), .B0(P2_EAX_REG_18__SCAN_IN), .B1(n12799), .Y(n12886));
  OAI21X1 g09613(.A0(n12798), .A1(n9936), .B0(n12886), .Y(P2_U2954));
  AOI22X1 g09614(.A0(n12796), .A1(P2_UWORD_REG_1__SCAN_IN), .B0(P2_EAX_REG_17__SCAN_IN), .B1(n12799), .Y(n12888));
  OAI21X1 g09615(.A0(n12798), .A1(n9955), .B0(n12888), .Y(P2_U2953));
  AOI22X1 g09616(.A0(n12796), .A1(P2_UWORD_REG_0__SCAN_IN), .B0(P2_EAX_REG_16__SCAN_IN), .B1(n12799), .Y(n12890));
  OAI21X1 g09617(.A0(n12798), .A1(n9974), .B0(n12890), .Y(P2_U2952));
  NOR2X1  g09618(.A(n9417), .B(P2_STATE_REG_0__SCAN_IN), .Y(n12892));
  NAND3X1 g09619(.A(n9724), .B(n12791), .C(n8976), .Y(n12893));
  NAND4X1 g09620(.A(n9518), .B(n9308), .C(n8975), .D(n9714), .Y(n12894));
  NAND2X1 g09621(.A(n12894), .B(n12893), .Y(n12895));
  AOI22X1 g09622(.A0(n9765), .A1(P2_STATE2_REG_1__SCAN_IN), .B0(n12892), .B1(n12895), .Y(n12896));
  INVX1   g09623(.A(n12896), .Y(n12897));
  NAND3X1 g09624(.A(n12897), .B(P2_LWORD_REG_0__SCAN_IN), .C(n8720), .Y(n12898));
  NOR2X1  g09625(.A(n12896), .B(n8720), .Y(n12899));
  AOI22X1 g09626(.A0(n12896), .A1(P2_DATAO_REG_0__SCAN_IN), .B0(P2_EAX_REG_0__SCAN_IN), .B1(n12899), .Y(n12900));
  NAND2X1 g09627(.A(n12900), .B(n12898), .Y(P2_U2951));
  NAND3X1 g09628(.A(n12897), .B(P2_LWORD_REG_1__SCAN_IN), .C(n8720), .Y(n12902));
  AOI22X1 g09629(.A0(n12896), .A1(P2_DATAO_REG_1__SCAN_IN), .B0(P2_EAX_REG_1__SCAN_IN), .B1(n12899), .Y(n12903));
  NAND2X1 g09630(.A(n12903), .B(n12902), .Y(P2_U2950));
  NAND3X1 g09631(.A(n12897), .B(P2_LWORD_REG_2__SCAN_IN), .C(n8720), .Y(n12905));
  AOI22X1 g09632(.A0(n12896), .A1(P2_DATAO_REG_2__SCAN_IN), .B0(P2_EAX_REG_2__SCAN_IN), .B1(n12899), .Y(n12906));
  NAND2X1 g09633(.A(n12906), .B(n12905), .Y(P2_U2949));
  NAND3X1 g09634(.A(n12897), .B(P2_LWORD_REG_3__SCAN_IN), .C(n8720), .Y(n12908));
  AOI22X1 g09635(.A0(n12896), .A1(P2_DATAO_REG_3__SCAN_IN), .B0(P2_EAX_REG_3__SCAN_IN), .B1(n12899), .Y(n12909));
  NAND2X1 g09636(.A(n12909), .B(n12908), .Y(P2_U2948));
  NAND3X1 g09637(.A(n12897), .B(P2_LWORD_REG_4__SCAN_IN), .C(n8720), .Y(n12911));
  AOI22X1 g09638(.A0(n12896), .A1(P2_DATAO_REG_4__SCAN_IN), .B0(P2_EAX_REG_4__SCAN_IN), .B1(n12899), .Y(n12912));
  NAND2X1 g09639(.A(n12912), .B(n12911), .Y(P2_U2947));
  NAND3X1 g09640(.A(n12897), .B(P2_LWORD_REG_5__SCAN_IN), .C(n8720), .Y(n12914));
  AOI22X1 g09641(.A0(n12896), .A1(P2_DATAO_REG_5__SCAN_IN), .B0(P2_EAX_REG_5__SCAN_IN), .B1(n12899), .Y(n12915));
  NAND2X1 g09642(.A(n12915), .B(n12914), .Y(P2_U2946));
  NAND3X1 g09643(.A(n12897), .B(P2_LWORD_REG_6__SCAN_IN), .C(n8720), .Y(n12917));
  AOI22X1 g09644(.A0(n12896), .A1(P2_DATAO_REG_6__SCAN_IN), .B0(P2_EAX_REG_6__SCAN_IN), .B1(n12899), .Y(n12918));
  NAND2X1 g09645(.A(n12918), .B(n12917), .Y(P2_U2945));
  NAND3X1 g09646(.A(n12897), .B(P2_LWORD_REG_7__SCAN_IN), .C(n8720), .Y(n12920));
  AOI22X1 g09647(.A0(n12896), .A1(P2_DATAO_REG_7__SCAN_IN), .B0(P2_EAX_REG_7__SCAN_IN), .B1(n12899), .Y(n12921));
  NAND2X1 g09648(.A(n12921), .B(n12920), .Y(P2_U2944));
  NAND3X1 g09649(.A(n12897), .B(P2_LWORD_REG_8__SCAN_IN), .C(n8720), .Y(n12923));
  AOI22X1 g09650(.A0(n12896), .A1(P2_DATAO_REG_8__SCAN_IN), .B0(P2_EAX_REG_8__SCAN_IN), .B1(n12899), .Y(n12924));
  NAND2X1 g09651(.A(n12924), .B(n12923), .Y(P2_U2943));
  NAND3X1 g09652(.A(n12897), .B(P2_LWORD_REG_9__SCAN_IN), .C(n8720), .Y(n12926));
  AOI22X1 g09653(.A0(n12896), .A1(P2_DATAO_REG_9__SCAN_IN), .B0(P2_EAX_REG_9__SCAN_IN), .B1(n12899), .Y(n12927));
  NAND2X1 g09654(.A(n12927), .B(n12926), .Y(P2_U2942));
  NAND3X1 g09655(.A(n12897), .B(P2_LWORD_REG_10__SCAN_IN), .C(n8720), .Y(n12929));
  AOI22X1 g09656(.A0(n12896), .A1(P2_DATAO_REG_10__SCAN_IN), .B0(P2_EAX_REG_10__SCAN_IN), .B1(n12899), .Y(n12930));
  NAND2X1 g09657(.A(n12930), .B(n12929), .Y(P2_U2941));
  NAND3X1 g09658(.A(n12897), .B(P2_LWORD_REG_11__SCAN_IN), .C(n8720), .Y(n12932));
  AOI22X1 g09659(.A0(n12896), .A1(P2_DATAO_REG_11__SCAN_IN), .B0(P2_EAX_REG_11__SCAN_IN), .B1(n12899), .Y(n12933));
  NAND2X1 g09660(.A(n12933), .B(n12932), .Y(P2_U2940));
  NAND3X1 g09661(.A(n12897), .B(P2_LWORD_REG_12__SCAN_IN), .C(n8720), .Y(n12935));
  AOI22X1 g09662(.A0(n12896), .A1(P2_DATAO_REG_12__SCAN_IN), .B0(P2_EAX_REG_12__SCAN_IN), .B1(n12899), .Y(n12936));
  NAND2X1 g09663(.A(n12936), .B(n12935), .Y(P2_U2939));
  NAND3X1 g09664(.A(n12897), .B(P2_LWORD_REG_13__SCAN_IN), .C(n8720), .Y(n12938));
  AOI22X1 g09665(.A0(n12896), .A1(P2_DATAO_REG_13__SCAN_IN), .B0(P2_EAX_REG_13__SCAN_IN), .B1(n12899), .Y(n12939));
  NAND2X1 g09666(.A(n12939), .B(n12938), .Y(P2_U2938));
  NAND3X1 g09667(.A(n12897), .B(P2_LWORD_REG_14__SCAN_IN), .C(n8720), .Y(n12941));
  AOI22X1 g09668(.A0(n12896), .A1(P2_DATAO_REG_14__SCAN_IN), .B0(P2_EAX_REG_14__SCAN_IN), .B1(n12899), .Y(n12942));
  NAND2X1 g09669(.A(n12942), .B(n12941), .Y(P2_U2937));
  NAND3X1 g09670(.A(n12897), .B(P2_LWORD_REG_15__SCAN_IN), .C(n8720), .Y(n12944));
  AOI22X1 g09671(.A0(n12896), .A1(P2_DATAO_REG_15__SCAN_IN), .B0(P2_EAX_REG_15__SCAN_IN), .B1(n12899), .Y(n12945));
  NAND2X1 g09672(.A(n12945), .B(n12944), .Y(P2_U2936));
  NAND3X1 g09673(.A(n12897), .B(P2_UWORD_REG_0__SCAN_IN), .C(n8720), .Y(n12947));
  NOR2X1  g09674(.A(n12896), .B(n9262), .Y(n12948));
  AOI22X1 g09675(.A0(n12896), .A1(P2_DATAO_REG_16__SCAN_IN), .B0(P2_EAX_REG_16__SCAN_IN), .B1(n12948), .Y(n12949));
  NAND2X1 g09676(.A(n12949), .B(n12947), .Y(P2_U2935));
  NAND3X1 g09677(.A(n12897), .B(P2_UWORD_REG_1__SCAN_IN), .C(n8720), .Y(n12951));
  AOI22X1 g09678(.A0(n12896), .A1(P2_DATAO_REG_17__SCAN_IN), .B0(P2_EAX_REG_17__SCAN_IN), .B1(n12948), .Y(n12952));
  NAND2X1 g09679(.A(n12952), .B(n12951), .Y(P2_U2934));
  NAND3X1 g09680(.A(n12897), .B(P2_UWORD_REG_2__SCAN_IN), .C(n8720), .Y(n12954));
  AOI22X1 g09681(.A0(n12896), .A1(P2_DATAO_REG_18__SCAN_IN), .B0(P2_EAX_REG_18__SCAN_IN), .B1(n12948), .Y(n12955));
  NAND2X1 g09682(.A(n12955), .B(n12954), .Y(P2_U2933));
  NAND3X1 g09683(.A(n12897), .B(P2_UWORD_REG_3__SCAN_IN), .C(n8720), .Y(n12957));
  AOI22X1 g09684(.A0(n12896), .A1(P2_DATAO_REG_19__SCAN_IN), .B0(P2_EAX_REG_19__SCAN_IN), .B1(n12948), .Y(n12958));
  NAND2X1 g09685(.A(n12958), .B(n12957), .Y(P2_U2932));
  NAND3X1 g09686(.A(n12897), .B(P2_UWORD_REG_4__SCAN_IN), .C(n8720), .Y(n12960));
  AOI22X1 g09687(.A0(n12896), .A1(P2_DATAO_REG_20__SCAN_IN), .B0(P2_EAX_REG_20__SCAN_IN), .B1(n12948), .Y(n12961));
  NAND2X1 g09688(.A(n12961), .B(n12960), .Y(P2_U2931));
  NAND3X1 g09689(.A(n12897), .B(P2_UWORD_REG_5__SCAN_IN), .C(n8720), .Y(n12963));
  AOI22X1 g09690(.A0(n12896), .A1(P2_DATAO_REG_21__SCAN_IN), .B0(P2_EAX_REG_21__SCAN_IN), .B1(n12948), .Y(n12964));
  NAND2X1 g09691(.A(n12964), .B(n12963), .Y(P2_U2930));
  NAND3X1 g09692(.A(n12897), .B(P2_UWORD_REG_6__SCAN_IN), .C(n8720), .Y(n12966));
  AOI22X1 g09693(.A0(n12896), .A1(P2_DATAO_REG_22__SCAN_IN), .B0(P2_EAX_REG_22__SCAN_IN), .B1(n12948), .Y(n12967));
  NAND2X1 g09694(.A(n12967), .B(n12966), .Y(P2_U2929));
  NAND3X1 g09695(.A(n12897), .B(P2_UWORD_REG_7__SCAN_IN), .C(n8720), .Y(n12969));
  AOI22X1 g09696(.A0(n12896), .A1(P2_DATAO_REG_23__SCAN_IN), .B0(P2_EAX_REG_23__SCAN_IN), .B1(n12948), .Y(n12970));
  NAND2X1 g09697(.A(n12970), .B(n12969), .Y(P2_U2928));
  NAND3X1 g09698(.A(n12897), .B(P2_UWORD_REG_8__SCAN_IN), .C(n8720), .Y(n12972));
  AOI22X1 g09699(.A0(n12896), .A1(P2_DATAO_REG_24__SCAN_IN), .B0(P2_EAX_REG_24__SCAN_IN), .B1(n12948), .Y(n12973));
  NAND2X1 g09700(.A(n12973), .B(n12972), .Y(P2_U2927));
  NAND3X1 g09701(.A(n12897), .B(P2_UWORD_REG_9__SCAN_IN), .C(n8720), .Y(n12975));
  AOI22X1 g09702(.A0(n12896), .A1(P2_DATAO_REG_25__SCAN_IN), .B0(P2_EAX_REG_25__SCAN_IN), .B1(n12948), .Y(n12976));
  NAND2X1 g09703(.A(n12976), .B(n12975), .Y(P2_U2926));
  NAND3X1 g09704(.A(n12897), .B(P2_UWORD_REG_10__SCAN_IN), .C(n8720), .Y(n12978));
  AOI22X1 g09705(.A0(n12896), .A1(P2_DATAO_REG_26__SCAN_IN), .B0(P2_EAX_REG_26__SCAN_IN), .B1(n12948), .Y(n12979));
  NAND2X1 g09706(.A(n12979), .B(n12978), .Y(P2_U2925));
  NAND3X1 g09707(.A(n12897), .B(P2_UWORD_REG_11__SCAN_IN), .C(n8720), .Y(n12981));
  AOI22X1 g09708(.A0(n12896), .A1(P2_DATAO_REG_27__SCAN_IN), .B0(P2_EAX_REG_27__SCAN_IN), .B1(n12948), .Y(n12982));
  NAND2X1 g09709(.A(n12982), .B(n12981), .Y(P2_U2924));
  NAND3X1 g09710(.A(n12897), .B(P2_UWORD_REG_12__SCAN_IN), .C(n8720), .Y(n12984));
  AOI22X1 g09711(.A0(n12896), .A1(P2_DATAO_REG_28__SCAN_IN), .B0(P2_EAX_REG_28__SCAN_IN), .B1(n12948), .Y(n12985));
  NAND2X1 g09712(.A(n12985), .B(n12984), .Y(P2_U2923));
  NAND3X1 g09713(.A(n12897), .B(P2_UWORD_REG_13__SCAN_IN), .C(n8720), .Y(n12987));
  AOI22X1 g09714(.A0(n12896), .A1(P2_DATAO_REG_29__SCAN_IN), .B0(P2_EAX_REG_29__SCAN_IN), .B1(n12948), .Y(n12988));
  NAND2X1 g09715(.A(n12988), .B(n12987), .Y(P2_U2922));
  NAND3X1 g09716(.A(n12897), .B(P2_UWORD_REG_14__SCAN_IN), .C(n8720), .Y(n12990));
  AOI22X1 g09717(.A0(n12896), .A1(P2_DATAO_REG_30__SCAN_IN), .B0(P2_EAX_REG_30__SCAN_IN), .B1(n12948), .Y(n12991));
  NAND2X1 g09718(.A(n12991), .B(n12990), .Y(P2_U2921));
  NOR2X1  g09719(.A(n12897), .B(n2967), .Y(P2_U2920));
  AOI21X1 g09720(.A0(n9464), .A1(n9411), .B0(n9732), .Y(n12994));
  NAND4X1 g09721(.A(n9975), .B(n9332), .C(n8884), .D(n12994), .Y(n12995));
  XOR2X1  g09722(.A(n10960), .B(n9771), .Y(n12996));
  NAND3X1 g09723(.A(n12996), .B(n12994), .C(n9434), .Y(n12997));
  INVX1   g09724(.A(n12994), .Y(n12998));
  NOR2X1  g09725(.A(n12998), .B(n8884), .Y(n12999));
  AOI22X1 g09726(.A0(n12998), .A1(P2_EAX_REG_0__SCAN_IN), .B0(n10959), .B1(n12999), .Y(n13000));
  NAND3X1 g09727(.A(n13000), .B(n12997), .C(n12995), .Y(P2_U2919));
  NAND4X1 g09728(.A(n9956), .B(n9332), .C(n8884), .D(n12994), .Y(n13002));
  NOR2X1  g09729(.A(n10960), .B(n9771), .Y(n13003));
  XOR2X1  g09730(.A(n13003), .B(n9784), .Y(n13004));
  NOR3X1  g09731(.A(n10960), .B(n10954), .C(n9771), .Y(n13005));
  NOR3X1  g09732(.A(n13003), .B(n10954), .C(n9996), .Y(n13006));
  AOI21X1 g09733(.A0(n13005), .A1(n9996), .B0(n13006), .Y(n13007));
  OAI21X1 g09734(.A0(n13004), .A1(n10953), .B0(n13007), .Y(n13008));
  NAND3X1 g09735(.A(n13008), .B(n12994), .C(n9434), .Y(n13009));
  AOI22X1 g09736(.A0(n12998), .A1(P2_EAX_REG_1__SCAN_IN), .B0(n10953), .B1(n12999), .Y(n13010));
  NAND3X1 g09737(.A(n13010), .B(n13009), .C(n13002), .Y(P2_U2918));
  NAND4X1 g09738(.A(n9937), .B(n9332), .C(n8884), .D(n12994), .Y(n13012));
  NAND2X1 g09739(.A(n13003), .B(n10953), .Y(n13013));
  NOR2X1  g09740(.A(n13003), .B(n10953), .Y(n13014));
  OAI21X1 g09741(.A0(n13014), .A1(n9784), .B0(n13013), .Y(n13015));
  XOR2X1  g09742(.A(n10940), .B(n9810), .Y(n13016));
  XOR2X1  g09743(.A(n13016), .B(n13015), .Y(n13017));
  NAND3X1 g09744(.A(n13017), .B(n12994), .C(n9434), .Y(n13018));
  AOI22X1 g09745(.A0(n12998), .A1(P2_EAX_REG_2__SCAN_IN), .B0(n10940), .B1(n12999), .Y(n13019));
  NAND3X1 g09746(.A(n13019), .B(n13018), .C(n13012), .Y(P2_U2917));
  NAND4X1 g09747(.A(n9918), .B(n9332), .C(n8884), .D(n12994), .Y(n13021));
  NOR3X1  g09748(.A(n10941), .B(n9809), .C(n9801), .Y(n13022));
  OAI21X1 g09749(.A0(n9809), .A1(n9801), .B0(n10941), .Y(n13023));
  AOI21X1 g09750(.A0(n13023), .A1(n13015), .B0(n13022), .Y(n13024));
  XOR2X1  g09751(.A(n11141), .B(n9827), .Y(n13025));
  XOR2X1  g09752(.A(n13025), .B(n13024), .Y(n13026));
  NAND3X1 g09753(.A(n13026), .B(n12994), .C(n9434), .Y(n13027));
  AOI22X1 g09754(.A0(n12998), .A1(P2_EAX_REG_3__SCAN_IN), .B0(n11141), .B1(n12999), .Y(n13028));
  NAND3X1 g09755(.A(n13028), .B(n13027), .C(n13021), .Y(P2_U2916));
  OAI21X1 g09756(.A0(n10960), .A1(n9771), .B0(n10954), .Y(n13030));
  AOI21X1 g09757(.A0(n13030), .A1(n9996), .B0(n13005), .Y(n13031));
  NAND3X1 g09758(.A(n9808), .B(n9812), .C(n10347), .Y(n13032));
  OAI21X1 g09759(.A0(n9760), .A1(n9791), .B0(n9789), .Y(n13033));
  NAND3X1 g09760(.A(n9796), .B(n9785), .C(P2_INSTQUEUE_REG_0__2__SCAN_IN), .Y(n13034));
  NAND3X1 g09761(.A(n9800), .B(n13034), .C(n13033), .Y(n13036));
  NAND3X1 g09762(.A(n10940), .B(n13036), .C(n13032), .Y(n13037));
  AOI21X1 g09763(.A0(n13036), .A1(n13032), .B0(n10940), .Y(n13038));
  OAI21X1 g09764(.A0(n13038), .A1(n13031), .B0(n13037), .Y(n13039));
  NOR2X1  g09765(.A(n10933), .B(n9827), .Y(n13040));
  NAND2X1 g09766(.A(n10933), .B(n9827), .Y(n13041));
  AOI21X1 g09767(.A0(n13041), .A1(n13039), .B0(n13040), .Y(n13042));
  INVX1   g09768(.A(n11201), .Y(n13043));
  NOR3X1  g09769(.A(n9823), .B(n9760), .C(n9824), .Y(n13044));
  OAI21X1 g09770(.A0(n9760), .A1(n9824), .B0(n9823), .Y(n13045));
  AOI21X1 g09771(.A0(n13045), .A1(n9813), .B0(n13044), .Y(n13046));
  NOR3X1  g09772(.A(n9470), .B(n9019), .C(n8720), .Y(n13047));
  INVX1   g09773(.A(n13047), .Y(n13048));
  INVX1   g09774(.A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .Y(n13049));
  NOR2X1  g09775(.A(n9760), .B(n13049), .Y(n13050));
  XOR2X1  g09776(.A(n13067), .B(n13046), .Y(n13052));
  XOR2X1  g09777(.A(n13052), .B(n13043), .Y(n13053));
  XOR2X1  g09778(.A(n13053), .B(n13042), .Y(n13054));
  NAND3X1 g09779(.A(n13054), .B(n12994), .C(n9434), .Y(n13055));
  NAND4X1 g09780(.A(n9899), .B(n9332), .C(n8884), .D(n12994), .Y(n13056));
  AOI22X1 g09781(.A0(n12998), .A1(P2_EAX_REG_4__SCAN_IN), .B0(n11201), .B1(n12999), .Y(n13057));
  NAND3X1 g09782(.A(n13057), .B(n13056), .C(n13055), .Y(P2_U2915));
  NAND2X1 g09783(.A(n13052), .B(n11201), .Y(n13059));
  NOR2X1  g09784(.A(n13052), .B(n11201), .Y(n13060));
  OAI21X1 g09785(.A0(n13060), .A1(n13042), .B0(n13059), .Y(n13061));
  OAI21X1 g09786(.A0(n9774), .A1(n9663), .B0(n9821), .Y(n13062));
  NAND2X1 g09787(.A(n9825), .B(n13062), .Y(n13063));
  NOR2X1  g09788(.A(n9825), .B(n13062), .Y(n13064));
  OAI21X1 g09789(.A0(n13064), .A1(n10349), .B0(n13063), .Y(n13065));
  NOR3X1  g09790(.A(n13048), .B(n9760), .C(n13049), .Y(n13066));
  NOR2X1  g09791(.A(n13050), .B(n13047), .Y(n13067));
  INVX1   g09792(.A(n13067), .Y(n13068));
  AOI21X1 g09793(.A0(n13068), .A1(n13065), .B0(n13066), .Y(n13069));
  INVX1   g09794(.A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .Y(n13070));
  NOR2X1  g09795(.A(n9760), .B(n13070), .Y(n13071));
  XOR2X1  g09796(.A(n13071), .B(n13069), .Y(n13072));
  NAND2X1 g09797(.A(n13072), .B(n11268), .Y(n13073));
  INVX1   g09798(.A(n13066), .Y(n13074));
  OAI21X1 g09799(.A0(n13067), .A1(n13046), .B0(n13074), .Y(n13075));
  XOR2X1  g09800(.A(n13071), .B(n13075), .Y(n13076));
  NAND2X1 g09801(.A(n13076), .B(n11269), .Y(n13077));
  NAND3X1 g09802(.A(n13077), .B(n13073), .C(n13061), .Y(n13078));
  NAND2X1 g09803(.A(n11141), .B(n10350), .Y(n13079));
  NOR2X1  g09804(.A(n11141), .B(n10350), .Y(n13080));
  OAI21X1 g09805(.A0(n13080), .A1(n13024), .B0(n13079), .Y(n13081));
  XOR2X1  g09806(.A(n13067), .B(n13065), .Y(n13082));
  NOR2X1  g09807(.A(n13082), .B(n13043), .Y(n13083));
  NAND2X1 g09808(.A(n13082), .B(n13043), .Y(n13084));
  AOI21X1 g09809(.A0(n13084), .A1(n13081), .B0(n13083), .Y(n13085));
  XOR2X1  g09810(.A(n13076), .B(n11268), .Y(n13086));
  NAND2X1 g09811(.A(n13086), .B(n13085), .Y(n13087));
  NAND4X1 g09812(.A(n13078), .B(n12994), .C(n9434), .D(n13087), .Y(n13088));
  NAND4X1 g09813(.A(n9880), .B(n9332), .C(n8884), .D(n12994), .Y(n13089));
  AOI22X1 g09814(.A0(n12998), .A1(P2_EAX_REG_5__SCAN_IN), .B0(n11269), .B1(n12999), .Y(n13090));
  NAND3X1 g09815(.A(n13090), .B(n13089), .C(n13088), .Y(P2_U2914));
  NAND2X1 g09816(.A(n13071), .B(n13075), .Y(n13092));
  INVX1   g09817(.A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .Y(n13093));
  NOR2X1  g09818(.A(n9760), .B(n13093), .Y(n13094));
  XOR2X1  g09819(.A(n13094), .B(n13092), .Y(n13095));
  XOR2X1  g09820(.A(n13095), .B(n11335), .Y(n13096));
  NOR2X1  g09821(.A(n13076), .B(n11269), .Y(n13097));
  OAI21X1 g09822(.A0(n13097), .A1(n13085), .B0(n13077), .Y(n13098));
  NAND2X1 g09823(.A(n13096), .B(n13098), .Y(n13100));
  OAI21X1 g09824(.A0(n13098), .A1(n13096), .B0(n13100), .Y(n13101));
  NAND3X1 g09825(.A(n13101), .B(n12994), .C(n9434), .Y(n13102));
  NAND4X1 g09826(.A(n9861), .B(n9332), .C(n8884), .D(n12994), .Y(n13103));
  AOI22X1 g09827(.A0(n12998), .A1(P2_EAX_REG_6__SCAN_IN), .B0(n11335), .B1(n12999), .Y(n13104));
  NAND3X1 g09828(.A(n13104), .B(n13103), .C(n13102), .Y(P2_U2913));
  INVX1   g09829(.A(n11335), .Y(n13106));
  NOR2X1  g09830(.A(n13095), .B(n13106), .Y(n13107));
  XOR2X1  g09831(.A(n11447), .B(n11442), .Y(n13108));
  NAND3X1 g09832(.A(n13094), .B(n13071), .C(n13075), .Y(n13109));
  INVX1   g09833(.A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .Y(n13110));
  NOR2X1  g09834(.A(n9760), .B(n13110), .Y(n13111));
  XOR2X1  g09835(.A(n13111), .B(n13109), .Y(n13112));
  AOI22X1 g09836(.A0(n13095), .A1(n13106), .B0(n13108), .B1(n13112), .Y(n13113));
  OAI21X1 g09837(.A0(n13107), .A1(n13098), .B0(n13113), .Y(n13114));
  NOR2X1  g09838(.A(n13112), .B(n13108), .Y(n13115));
  NOR2X1  g09839(.A(n12998), .B(n9332), .Y(n13116));
  INVX1   g09840(.A(n13116), .Y(n13117));
  NOR3X1  g09841(.A(n13069), .B(n9760), .C(n13070), .Y(n13118));
  XOR2X1  g09842(.A(n13094), .B(n13118), .Y(n13119));
  OAI21X1 g09843(.A0(n13119), .A1(n11335), .B0(n13098), .Y(n13120));
  OAI22X1 g09844(.A0(n13095), .A1(n13106), .B0(n11449), .B1(n13112), .Y(n13121));
  AOI21X1 g09845(.A0(n13112), .A1(n11449), .B0(n13121), .Y(n13122));
  AOI21X1 g09846(.A0(n13122), .A1(n13120), .B0(n13117), .Y(n13123));
  OAI21X1 g09847(.A0(n13115), .A1(n13114), .B0(n13123), .Y(n13124));
  NAND4X1 g09848(.A(n9744), .B(n9332), .C(n8884), .D(n12994), .Y(n13125));
  AOI22X1 g09849(.A0(n12998), .A1(P2_EAX_REG_7__SCAN_IN), .B0(n11449), .B1(n12999), .Y(n13126));
  NAND3X1 g09850(.A(n13126), .B(n13125), .C(n13124), .Y(P2_U2912));
  NOR2X1  g09851(.A(n13072), .B(n11268), .Y(n13128));
  AOI21X1 g09852(.A0(n13073), .A1(n13061), .B0(n13128), .Y(n13129));
  NAND2X1 g09853(.A(n13119), .B(n11335), .Y(n13130));
  INVX1   g09854(.A(n13111), .Y(n13131));
  XOR2X1  g09855(.A(n13131), .B(n13109), .Y(n13132));
  OAI22X1 g09856(.A0(n13119), .A1(n11335), .B0(n11449), .B1(n13132), .Y(n13133));
  AOI21X1 g09857(.A0(n13130), .A1(n13129), .B0(n13133), .Y(n13134));
  NOR2X1  g09858(.A(n13115), .B(n13134), .Y(n13135));
  NAND4X1 g09859(.A(n13094), .B(n13071), .C(n13075), .D(n13111), .Y(n13136));
  NOR2X1  g09860(.A(n11528), .B(n9760), .Y(n13137));
  INVX1   g09861(.A(n13137), .Y(n13138));
  XOR2X1  g09862(.A(n13138), .B(n13136), .Y(n13139));
  XOR2X1  g09863(.A(n13139), .B(n11533), .Y(n13140));
  XOR2X1  g09864(.A(n13140), .B(n13135), .Y(n13141));
  NAND3X1 g09865(.A(n13141), .B(n12994), .C(n9434), .Y(n13142));
  NAND4X1 g09866(.A(n12842), .B(n9332), .C(n8884), .D(n12994), .Y(n13143));
  AOI22X1 g09867(.A0(n12998), .A1(P2_EAX_REG_8__SCAN_IN), .B0(n11532), .B1(n12999), .Y(n13144));
  NAND3X1 g09868(.A(n13144), .B(n13143), .C(n13142), .Y(P2_U2911));
  NAND2X1 g09869(.A(n13139), .B(n11532), .Y(n13146));
  OAI22X1 g09870(.A0(n13115), .A1(n13134), .B0(n11532), .B1(n13139), .Y(n13147));
  NOR2X1  g09871(.A(n13138), .B(n13136), .Y(n13148));
  NOR2X1  g09872(.A(n11582), .B(n9760), .Y(n13149));
  XOR2X1  g09873(.A(n13149), .B(n13148), .Y(n13150));
  INVX1   g09874(.A(n13150), .Y(n13151));
  AOI22X1 g09875(.A0(n13147), .A1(n13146), .B0(n11586), .B1(n13151), .Y(n13152));
  NAND2X1 g09876(.A(n13150), .B(n11587), .Y(n13153));
  NAND2X1 g09877(.A(n13153), .B(n13152), .Y(n13154));
  XOR2X1  g09878(.A(n13150), .B(n11586), .Y(n13155));
  NAND3X1 g09879(.A(n13155), .B(n13147), .C(n13146), .Y(n13156));
  NAND3X1 g09880(.A(n13156), .B(n13154), .C(n13116), .Y(n13157));
  NAND4X1 g09881(.A(n12836), .B(n9332), .C(n8884), .D(n12994), .Y(n13158));
  AOI22X1 g09882(.A0(n12998), .A1(P2_EAX_REG_9__SCAN_IN), .B0(n11587), .B1(n12999), .Y(n13159));
  NAND3X1 g09883(.A(n13159), .B(n13158), .C(n13157), .Y(P2_U2910));
  NOR2X1  g09884(.A(n13151), .B(n11586), .Y(n13161));
  NOR4X1  g09885(.A(n11582), .B(n11528), .C(n9760), .D(n13136), .Y(n13162));
  NOR2X1  g09886(.A(n11635), .B(n9760), .Y(n13163));
  XOR2X1  g09887(.A(n13163), .B(n13162), .Y(n13164));
  XOR2X1  g09888(.A(n13164), .B(n11639), .Y(n13165));
  NOR3X1  g09889(.A(n13165), .B(n13161), .C(n13152), .Y(n13166));
  INVX1   g09890(.A(n13146), .Y(n13167));
  NAND2X1 g09891(.A(n13132), .B(n11449), .Y(n13168));
  INVX1   g09892(.A(n13139), .Y(n13169));
  AOI22X1 g09893(.A0(n13168), .A1(n13114), .B0(n11533), .B1(n13169), .Y(n13170));
  OAI22X1 g09894(.A0(n13170), .A1(n13167), .B0(n11587), .B1(n13150), .Y(n13171));
  INVX1   g09895(.A(n13164), .Y(n13172));
  NAND2X1 g09896(.A(n13172), .B(n11639), .Y(n13173));
  INVX1   g09897(.A(n11639), .Y(n13174));
  NAND2X1 g09898(.A(n13164), .B(n13174), .Y(n13175));
  AOI22X1 g09899(.A0(n13173), .A1(n13175), .B0(n13153), .B1(n13171), .Y(n13176));
  OAI21X1 g09900(.A0(n13176), .A1(n13166), .B0(n13116), .Y(n13177));
  NAND4X1 g09901(.A(n12830), .B(n9332), .C(n8884), .D(n12994), .Y(n13178));
  AOI22X1 g09902(.A0(n12998), .A1(P2_EAX_REG_10__SCAN_IN), .B0(n13174), .B1(n12999), .Y(n13179));
  NAND3X1 g09903(.A(n13179), .B(n13178), .C(n13177), .Y(P2_U2909));
  NOR2X1  g09904(.A(n13172), .B(n11639), .Y(n13181));
  NOR3X1  g09905(.A(n13181), .B(n13161), .C(n13152), .Y(n13182));
  NAND2X1 g09906(.A(n13163), .B(n13162), .Y(n13183));
  NOR2X1  g09907(.A(n11683), .B(n9760), .Y(n13184));
  XOR2X1  g09908(.A(n13184), .B(n13183), .Y(n13185));
  AOI22X1 g09909(.A0(n13172), .A1(n11639), .B0(n11687), .B1(n13185), .Y(n13186));
  INVX1   g09910(.A(n13186), .Y(n13187));
  NOR2X1  g09911(.A(n13185), .B(n11687), .Y(n13188));
  NOR3X1  g09912(.A(n13188), .B(n13187), .C(n13182), .Y(n13189));
  AOI22X1 g09913(.A0(n13153), .A1(n13171), .B0(n11639), .B1(n13172), .Y(n13190));
  INVX1   g09914(.A(n13185), .Y(n13191));
  AOI21X1 g09915(.A0(n13191), .A1(n11687), .B0(n13181), .Y(n13192));
  OAI21X1 g09916(.A0(n13191), .A1(n11687), .B0(n13192), .Y(n13193));
  OAI21X1 g09917(.A0(n13193), .A1(n13190), .B0(n13116), .Y(n13194));
  NAND2X1 g09918(.A(n12994), .B(n8884), .Y(n13195));
  NOR2X1  g09919(.A(n13195), .B(n9434), .Y(n13196));
  INVX1   g09920(.A(n12999), .Y(n13197));
  NAND2X1 g09921(.A(n12998), .B(P2_EAX_REG_11__SCAN_IN), .Y(n13198));
  OAI21X1 g09922(.A0(n13197), .A1(n11687), .B0(n13198), .Y(n13199));
  AOI21X1 g09923(.A0(n13196), .A1(n12824), .B0(n13199), .Y(n13200));
  OAI21X1 g09924(.A0(n13194), .A1(n13189), .B0(n13200), .Y(P2_U2908));
  NAND3X1 g09925(.A(n13175), .B(n13153), .C(n13171), .Y(n13202));
  AOI21X1 g09926(.A0(n13186), .A1(n13202), .B0(n13188), .Y(n13203));
  NAND3X1 g09927(.A(n13184), .B(n13163), .C(n13162), .Y(n13204));
  NOR2X1  g09928(.A(n11736), .B(n9760), .Y(n13205));
  XOR2X1  g09929(.A(n13205), .B(n13204), .Y(n13206));
  XOR2X1  g09930(.A(n13206), .B(n11741), .Y(n13207));
  XOR2X1  g09931(.A(n13207), .B(n13203), .Y(n13208));
  NAND2X1 g09932(.A(n12998), .B(P2_EAX_REG_12__SCAN_IN), .Y(n13209));
  OAI21X1 g09933(.A0(n13197), .A1(n11741), .B0(n13209), .Y(n13210));
  AOI21X1 g09934(.A0(n13196), .A1(n12818), .B0(n13210), .Y(n13211));
  OAI21X1 g09935(.A0(n13208), .A1(n13117), .B0(n13211), .Y(P2_U2907));
  OAI22X1 g09936(.A0(n13185), .A1(n11687), .B0(n13182), .B1(n13187), .Y(n13213));
  NOR2X1  g09937(.A(n13206), .B(n11741), .Y(n13214));
  NAND2X1 g09938(.A(n13206), .B(n11741), .Y(n13215));
  AOI21X1 g09939(.A0(n13215), .A1(n13213), .B0(n13214), .Y(n13216));
  NAND4X1 g09940(.A(n13184), .B(n13163), .C(n13162), .D(n13205), .Y(n13217));
  NOR2X1  g09941(.A(n11790), .B(n9760), .Y(n13218));
  XOR2X1  g09942(.A(n13218), .B(n13217), .Y(n13219));
  INVX1   g09943(.A(n13219), .Y(n13220));
  NOR2X1  g09944(.A(n13220), .B(n11796), .Y(n13221));
  NOR2X1  g09945(.A(n13219), .B(n11795), .Y(n13222));
  NOR3X1  g09946(.A(n13222), .B(n13221), .C(n13216), .Y(n13223));
  INVX1   g09947(.A(n13214), .Y(n13224));
  INVX1   g09948(.A(n13215), .Y(n13225));
  OAI21X1 g09949(.A0(n13225), .A1(n13203), .B0(n13224), .Y(n13226));
  XOR2X1  g09950(.A(n13219), .B(n11795), .Y(n13227));
  OAI21X1 g09951(.A0(n13227), .A1(n13226), .B0(n13116), .Y(n13228));
  INVX1   g09952(.A(n13196), .Y(n13229));
  NAND2X1 g09953(.A(n12998), .B(P2_EAX_REG_13__SCAN_IN), .Y(n13230));
  OAI21X1 g09954(.A0(n13229), .A1(n12811), .B0(n13230), .Y(n13231));
  AOI21X1 g09955(.A0(n12999), .A1(n11796), .B0(n13231), .Y(n13232));
  OAI21X1 g09956(.A0(n13228), .A1(n13223), .B0(n13232), .Y(P2_U2906));
  NOR3X1  g09957(.A(n13217), .B(n11790), .C(n9760), .Y(n13234));
  NOR2X1  g09958(.A(n11842), .B(n9760), .Y(n13235));
  INVX1   g09959(.A(n13235), .Y(n13236));
  XOR2X1  g09960(.A(n13236), .B(n13234), .Y(n13237));
  XOR2X1  g09961(.A(n13237), .B(n11847), .Y(n13238));
  INVX1   g09962(.A(n13221), .Y(n13239));
  AOI21X1 g09963(.A0(n13239), .A1(n13226), .B0(n13222), .Y(n13240));
  NOR2X1  g09964(.A(n13238), .B(n13240), .Y(n13242));
  AOI21X1 g09965(.A0(n13240), .A1(n13238), .B0(n13242), .Y(n13243));
  NAND2X1 g09966(.A(n12998), .B(P2_EAX_REG_14__SCAN_IN), .Y(n13244));
  OAI21X1 g09967(.A0(n13229), .A1(n12804), .B0(n13244), .Y(n13245));
  AOI21X1 g09968(.A0(n12999), .A1(n11848), .B0(n13245), .Y(n13246));
  OAI21X1 g09969(.A0(n13243), .A1(n13117), .B0(n13246), .Y(P2_U2905));
  INVX1   g09970(.A(n13222), .Y(n13248));
  OAI21X1 g09971(.A0(n13221), .A1(n13216), .B0(n13248), .Y(n13249));
  NOR2X1  g09972(.A(n13237), .B(n11847), .Y(n13250));
  NOR4X1  g09973(.A(n11842), .B(n11790), .C(n9760), .D(n13217), .Y(n13251));
  NOR2X1  g09974(.A(n11891), .B(n9760), .Y(n13252));
  INVX1   g09975(.A(n13252), .Y(n13253));
  XOR2X1  g09976(.A(n13253), .B(n13251), .Y(n13254));
  AOI22X1 g09977(.A0(n13237), .A1(n11847), .B0(n11895), .B1(n13254), .Y(n13255));
  OAI21X1 g09978(.A0(n13250), .A1(n13249), .B0(n13255), .Y(n13256));
  NOR2X1  g09979(.A(n13254), .B(n11895), .Y(n13257));
  NOR2X1  g09980(.A(n13257), .B(n13256), .Y(n13258));
  INVX1   g09981(.A(n13237), .Y(n13259));
  NOR2X1  g09982(.A(n13259), .B(n11848), .Y(n13260));
  OAI22X1 g09983(.A0(n13237), .A1(n11847), .B0(n11896), .B1(n13254), .Y(n13261));
  AOI21X1 g09984(.A0(n13254), .A1(n11896), .B0(n13261), .Y(n13262));
  OAI21X1 g09985(.A0(n13260), .A1(n13240), .B0(n13262), .Y(n13263));
  NAND2X1 g09986(.A(n13263), .B(n13116), .Y(n13264));
  NAND2X1 g09987(.A(n12998), .B(P2_EAX_REG_15__SCAN_IN), .Y(n13265));
  OAI21X1 g09988(.A0(n13229), .A1(n12790), .B0(n13265), .Y(n13266));
  AOI21X1 g09989(.A0(n12999), .A1(n11896), .B0(n13266), .Y(n13267));
  OAI21X1 g09990(.A0(n13264), .A1(n13258), .B0(n13267), .Y(P2_U2904));
  OAI21X1 g09991(.A0(n13254), .A1(n11895), .B0(n13256), .Y(n13269));
  INVX1   g09992(.A(n13234), .Y(n13270));
  NOR3X1  g09993(.A(n13253), .B(n13236), .C(n13270), .Y(n13271));
  AOI22X1 g09994(.A0(n9003), .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B0(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(n9002), .Y(n13274));
  AOI22X1 g09995(.A0(n8994), .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B0(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(n8993), .Y(n13277));
  AOI22X1 g09996(.A0(n8997), .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B0(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(n8996), .Y(n13280));
  AOI22X1 g09997(.A0(n8990), .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B0(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(n8989), .Y(n13283));
  NAND4X1 g09998(.A(n13280), .B(n13277), .C(n13274), .D(n13283), .Y(n13284));
  AOI22X1 g09999(.A0(n8981), .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B0(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(n8980), .Y(n13287));
  AOI22X1 g10000(.A0(n9000), .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B0(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(n8999), .Y(n13290));
  AOI22X1 g10001(.A0(n8987), .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B0(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(n8986), .Y(n13293));
  AOI22X1 g10002(.A0(n8984), .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B0(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(n8983), .Y(n13296));
  NAND4X1 g10003(.A(n13293), .B(n13290), .C(n13287), .D(n13296), .Y(n13297));
  OAI22X1 g10004(.A0(n13284), .A1(n13297), .B0(n9785), .B1(n9479), .Y(n13298));
  XOR2X1  g10005(.A(n13298), .B(n13271), .Y(n13299));
  XOR2X1  g10006(.A(n13299), .B(n11942), .Y(n13300));
  XOR2X1  g10007(.A(n13300), .B(n13269), .Y(n13301));
  NOR2X1  g10008(.A(n13195), .B(n9470), .Y(n13302));
  INVX1   g10009(.A(n13302), .Y(n13303));
  NOR2X1  g10010(.A(n13195), .B(n8825), .Y(n13304));
  AOI22X1 g10011(.A0(n12998), .A1(P2_EAX_REG_16__SCAN_IN), .B0(n9975), .B1(n13304), .Y(n13305));
  OAI21X1 g10012(.A0(n13303), .A1(n9984), .B0(n13305), .Y(n13306));
  AOI21X1 g10013(.A0(n12999), .A1(n11942), .B0(n13306), .Y(n13307));
  OAI21X1 g10014(.A0(n13301), .A1(n13117), .B0(n13307), .Y(P2_U2903));
  NOR2X1  g10015(.A(n13299), .B(n11941), .Y(n13309));
  NAND2X1 g10016(.A(n13299), .B(n11941), .Y(n13310));
  AOI21X1 g10017(.A0(n13310), .A1(n13269), .B0(n13309), .Y(n13311));
  NOR4X1  g10018(.A(n13253), .B(n13236), .C(n13270), .D(n13298), .Y(n13312));
  AOI22X1 g10019(.A0(n9003), .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B0(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(n9002), .Y(n13313));
  AOI22X1 g10020(.A0(n8994), .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B0(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(n8993), .Y(n13314));
  AOI22X1 g10021(.A0(n8997), .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B0(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(n8996), .Y(n13315));
  AOI22X1 g10022(.A0(n8990), .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B0(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(n8989), .Y(n13316));
  NAND4X1 g10023(.A(n13315), .B(n13314), .C(n13313), .D(n13316), .Y(n13317));
  AOI22X1 g10024(.A0(n8981), .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B0(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(n8980), .Y(n13318));
  AOI22X1 g10025(.A0(n9000), .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B0(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(n8999), .Y(n13319));
  AOI22X1 g10026(.A0(n8987), .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B0(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(n8986), .Y(n13320));
  AOI22X1 g10027(.A0(n8984), .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B0(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(n8983), .Y(n13321));
  NAND4X1 g10028(.A(n13320), .B(n13319), .C(n13318), .D(n13321), .Y(n13322));
  OAI22X1 g10029(.A0(n13317), .A1(n13322), .B0(n9785), .B1(n9479), .Y(n13323));
  XOR2X1  g10030(.A(n13323), .B(n13312), .Y(n13324));
  XOR2X1  g10031(.A(n13324), .B(n11979), .Y(n13325));
  XOR2X1  g10032(.A(n13325), .B(n13311), .Y(n13326));
  AOI22X1 g10033(.A0(n12998), .A1(P2_EAX_REG_17__SCAN_IN), .B0(n9956), .B1(n13304), .Y(n13327));
  OAI21X1 g10034(.A0(n13303), .A1(n9965), .B0(n13327), .Y(n13328));
  AOI21X1 g10035(.A0(n12999), .A1(n11980), .B0(n13328), .Y(n13329));
  OAI21X1 g10036(.A0(n13326), .A1(n13117), .B0(n13329), .Y(P2_U2902));
  NOR2X1  g10037(.A(n13324), .B(n11979), .Y(n13331));
  INVX1   g10038(.A(n13331), .Y(n13332));
  NAND2X1 g10039(.A(n13324), .B(n11979), .Y(n13333));
  INVX1   g10040(.A(n13333), .Y(n13334));
  OAI21X1 g10041(.A0(n13334), .A1(n13311), .B0(n13332), .Y(n13335));
  INVX1   g10042(.A(n13312), .Y(n13336));
  NOR2X1  g10043(.A(n13323), .B(n13336), .Y(n13337));
  AOI22X1 g10044(.A0(n9003), .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B0(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(n9002), .Y(n13338));
  AOI22X1 g10045(.A0(n8994), .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B0(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(n8993), .Y(n13339));
  AOI22X1 g10046(.A0(n8997), .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B0(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(n8996), .Y(n13340));
  AOI22X1 g10047(.A0(n8990), .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B0(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(n8989), .Y(n13341));
  NAND4X1 g10048(.A(n13340), .B(n13339), .C(n13338), .D(n13341), .Y(n13342));
  AOI22X1 g10049(.A0(n8981), .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B0(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(n8980), .Y(n13343));
  AOI22X1 g10050(.A0(n9000), .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B0(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(n8999), .Y(n13344));
  AOI22X1 g10051(.A0(n8987), .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B0(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(n8986), .Y(n13345));
  AOI22X1 g10052(.A0(n8984), .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B0(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(n8983), .Y(n13346));
  NAND4X1 g10053(.A(n13345), .B(n13344), .C(n13343), .D(n13346), .Y(n13347));
  OAI22X1 g10054(.A0(n13342), .A1(n13347), .B0(n9785), .B1(n9479), .Y(n13348));
  XOR2X1  g10055(.A(n13348), .B(n13337), .Y(n13349));
  XOR2X1  g10056(.A(n13349), .B(n12018), .Y(n13350));
  XOR2X1  g10057(.A(n13350), .B(n13335), .Y(n13351));
  AOI22X1 g10058(.A0(n12998), .A1(P2_EAX_REG_18__SCAN_IN), .B0(n9937), .B1(n13304), .Y(n13352));
  OAI21X1 g10059(.A0(n13303), .A1(n9946), .B0(n13352), .Y(n13353));
  AOI21X1 g10060(.A0(n12999), .A1(n12018), .B0(n13353), .Y(n13354));
  OAI21X1 g10061(.A0(n13351), .A1(n13117), .B0(n13354), .Y(P2_U2901));
  NOR2X1  g10062(.A(n13349), .B(n12017), .Y(n13356));
  INVX1   g10063(.A(n13349), .Y(n13357));
  NOR2X1  g10064(.A(n13357), .B(n12018), .Y(n13358));
  INVX1   g10065(.A(n13358), .Y(n13359));
  AOI21X1 g10066(.A0(n13359), .A1(n13335), .B0(n13356), .Y(n13360));
  NOR3X1  g10067(.A(n13348), .B(n13323), .C(n13336), .Y(n13361));
  AOI22X1 g10068(.A0(n9003), .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B0(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(n9002), .Y(n13362));
  AOI22X1 g10069(.A0(n8994), .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B0(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(n8993), .Y(n13363));
  AOI22X1 g10070(.A0(n8997), .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B0(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(n8996), .Y(n13364));
  AOI22X1 g10071(.A0(n8990), .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B0(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(n8989), .Y(n13365));
  NAND4X1 g10072(.A(n13364), .B(n13363), .C(n13362), .D(n13365), .Y(n13366));
  AOI22X1 g10073(.A0(n8981), .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B0(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(n8980), .Y(n13367));
  AOI22X1 g10074(.A0(n9000), .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B0(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(n8999), .Y(n13368));
  AOI22X1 g10075(.A0(n8987), .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B0(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(n8986), .Y(n13369));
  AOI22X1 g10076(.A0(n8984), .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B0(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(n8983), .Y(n13370));
  NAND4X1 g10077(.A(n13369), .B(n13368), .C(n13367), .D(n13370), .Y(n13371));
  OAI22X1 g10078(.A0(n13366), .A1(n13371), .B0(n9785), .B1(n9479), .Y(n13372));
  XOR2X1  g10079(.A(n13372), .B(n13361), .Y(n13373));
  XOR2X1  g10080(.A(n13373), .B(n12057), .Y(n13374));
  XOR2X1  g10081(.A(n13374), .B(n13360), .Y(n13375));
  AOI22X1 g10082(.A0(n12998), .A1(P2_EAX_REG_19__SCAN_IN), .B0(n9918), .B1(n13304), .Y(n13376));
  OAI21X1 g10083(.A0(n13303), .A1(n9927), .B0(n13376), .Y(n13377));
  AOI21X1 g10084(.A0(n12999), .A1(n12058), .B0(n13377), .Y(n13378));
  OAI21X1 g10085(.A0(n13375), .A1(n13117), .B0(n13378), .Y(P2_U2900));
  NOR2X1  g10086(.A(n13373), .B(n12057), .Y(n13380));
  INVX1   g10087(.A(n13380), .Y(n13381));
  NAND2X1 g10088(.A(n13373), .B(n12057), .Y(n13382));
  INVX1   g10089(.A(n13382), .Y(n13383));
  OAI21X1 g10090(.A0(n13383), .A1(n13360), .B0(n13381), .Y(n13384));
  NOR4X1  g10091(.A(n13348), .B(n13323), .C(n13336), .D(n13372), .Y(n13385));
  AOI22X1 g10092(.A0(n9003), .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B0(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(n9002), .Y(n13386));
  AOI22X1 g10093(.A0(n8994), .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B0(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(n8993), .Y(n13387));
  AOI22X1 g10094(.A0(n8997), .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B0(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(n8996), .Y(n13388));
  AOI22X1 g10095(.A0(n8990), .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B0(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(n8989), .Y(n13389));
  NAND4X1 g10096(.A(n13388), .B(n13387), .C(n13386), .D(n13389), .Y(n13390));
  AOI22X1 g10097(.A0(n8981), .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B0(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(n8980), .Y(n13391));
  AOI22X1 g10098(.A0(n9000), .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B0(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(n8999), .Y(n13392));
  AOI22X1 g10099(.A0(n8987), .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B0(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(n8986), .Y(n13393));
  AOI22X1 g10100(.A0(n8984), .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B0(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(n8983), .Y(n13394));
  NAND4X1 g10101(.A(n13393), .B(n13392), .C(n13391), .D(n13394), .Y(n13395));
  OAI22X1 g10102(.A0(n13390), .A1(n13395), .B0(n9785), .B1(n9479), .Y(n13396));
  XOR2X1  g10103(.A(n13396), .B(n13385), .Y(n13397));
  XOR2X1  g10104(.A(n13397), .B(n12098), .Y(n13398));
  XOR2X1  g10105(.A(n13398), .B(n13384), .Y(n13399));
  AOI22X1 g10106(.A0(n12998), .A1(P2_EAX_REG_20__SCAN_IN), .B0(n9899), .B1(n13304), .Y(n13400));
  OAI21X1 g10107(.A0(n13303), .A1(n9908), .B0(n13400), .Y(n13401));
  AOI21X1 g10108(.A0(n12999), .A1(n12098), .B0(n13401), .Y(n13402));
  OAI21X1 g10109(.A0(n13399), .A1(n13117), .B0(n13402), .Y(P2_U2899));
  NOR2X1  g10110(.A(n13397), .B(n12097), .Y(n13404));
  INVX1   g10111(.A(n13397), .Y(n13405));
  NOR2X1  g10112(.A(n13405), .B(n12098), .Y(n13406));
  INVX1   g10113(.A(n13406), .Y(n13407));
  AOI21X1 g10114(.A0(n13407), .A1(n13384), .B0(n13404), .Y(n13408));
  INVX1   g10115(.A(n13385), .Y(n13409));
  NOR2X1  g10116(.A(n13396), .B(n13409), .Y(n13410));
  AOI22X1 g10117(.A0(n9003), .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B0(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(n9002), .Y(n13411));
  AOI22X1 g10118(.A0(n8994), .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B0(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(n8993), .Y(n13412));
  AOI22X1 g10119(.A0(n8997), .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B0(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(n8996), .Y(n13413));
  AOI22X1 g10120(.A0(n8990), .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B0(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(n8989), .Y(n13414));
  NAND4X1 g10121(.A(n13413), .B(n13412), .C(n13411), .D(n13414), .Y(n13415));
  AOI22X1 g10122(.A0(n8981), .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B0(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(n8980), .Y(n13416));
  AOI22X1 g10123(.A0(n9000), .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B0(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(n8999), .Y(n13417));
  AOI22X1 g10124(.A0(n8987), .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B0(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(n8986), .Y(n13418));
  AOI22X1 g10125(.A0(n8984), .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B0(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(n8983), .Y(n13419));
  NAND4X1 g10126(.A(n13418), .B(n13417), .C(n13416), .D(n13419), .Y(n13420));
  OAI22X1 g10127(.A0(n13415), .A1(n13420), .B0(n9785), .B1(n9479), .Y(n13421));
  XOR2X1  g10128(.A(n13421), .B(n13410), .Y(n13422));
  XOR2X1  g10129(.A(n13422), .B(n12137), .Y(n13423));
  XOR2X1  g10130(.A(n13423), .B(n13408), .Y(n13424));
  AOI22X1 g10131(.A0(n12998), .A1(P2_EAX_REG_21__SCAN_IN), .B0(n9880), .B1(n13304), .Y(n13425));
  OAI21X1 g10132(.A0(n13303), .A1(n9889), .B0(n13425), .Y(n13426));
  AOI21X1 g10133(.A0(n12999), .A1(n12138), .B0(n13426), .Y(n13427));
  OAI21X1 g10134(.A0(n13424), .A1(n13117), .B0(n13427), .Y(P2_U2898));
  NOR2X1  g10135(.A(n13422), .B(n12137), .Y(n13429));
  INVX1   g10136(.A(n13429), .Y(n13430));
  NAND2X1 g10137(.A(n13422), .B(n12137), .Y(n13431));
  INVX1   g10138(.A(n13431), .Y(n13432));
  OAI21X1 g10139(.A0(n13432), .A1(n13408), .B0(n13430), .Y(n13433));
  NOR3X1  g10140(.A(n13421), .B(n13396), .C(n13409), .Y(n13434));
  AOI22X1 g10141(.A0(n9003), .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B0(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(n9002), .Y(n13435));
  AOI22X1 g10142(.A0(n8994), .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B0(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(n8993), .Y(n13436));
  AOI22X1 g10143(.A0(n8997), .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B0(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(n8996), .Y(n13437));
  AOI22X1 g10144(.A0(n8990), .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B0(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(n8989), .Y(n13438));
  NAND4X1 g10145(.A(n13437), .B(n13436), .C(n13435), .D(n13438), .Y(n13439));
  AOI22X1 g10146(.A0(n8981), .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B0(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(n8980), .Y(n13440));
  AOI22X1 g10147(.A0(n9000), .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B0(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(n8999), .Y(n13441));
  AOI22X1 g10148(.A0(n8987), .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B0(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(n8986), .Y(n13442));
  AOI22X1 g10149(.A0(n8984), .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B0(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(n8983), .Y(n13443));
  NAND4X1 g10150(.A(n13442), .B(n13441), .C(n13440), .D(n13443), .Y(n13444));
  OAI22X1 g10151(.A0(n13439), .A1(n13444), .B0(n9785), .B1(n9479), .Y(n13445));
  XOR2X1  g10152(.A(n13445), .B(n13434), .Y(n13446));
  XOR2X1  g10153(.A(n13446), .B(n12176), .Y(n13447));
  XOR2X1  g10154(.A(n13447), .B(n13433), .Y(n13448));
  AOI22X1 g10155(.A0(n12998), .A1(P2_EAX_REG_22__SCAN_IN), .B0(n9861), .B1(n13304), .Y(n13449));
  OAI21X1 g10156(.A0(n13303), .A1(n9870), .B0(n13449), .Y(n13450));
  AOI21X1 g10157(.A0(n12999), .A1(n12176), .B0(n13450), .Y(n13451));
  OAI21X1 g10158(.A0(n13448), .A1(n13117), .B0(n13451), .Y(P2_U2897));
  NOR2X1  g10159(.A(n13446), .B(n12175), .Y(n13453));
  INVX1   g10160(.A(n13446), .Y(n13454));
  NOR2X1  g10161(.A(n13454), .B(n12176), .Y(n13455));
  INVX1   g10162(.A(n13455), .Y(n13456));
  AOI21X1 g10163(.A0(n13456), .A1(n13433), .B0(n13453), .Y(n13457));
  NOR4X1  g10164(.A(n13421), .B(n13396), .C(n13409), .D(n13445), .Y(n13458));
  INVX1   g10165(.A(n9479), .Y(n13459));
  AOI22X1 g10166(.A0(n9003), .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B0(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(n9002), .Y(n13460));
  AOI22X1 g10167(.A0(n8994), .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B0(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(n8993), .Y(n13461));
  AOI22X1 g10168(.A0(n8997), .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B0(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(n8996), .Y(n13462));
  AOI22X1 g10169(.A0(n8990), .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B0(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(n8989), .Y(n13463));
  NAND4X1 g10170(.A(n13462), .B(n13461), .C(n13460), .D(n13463), .Y(n13464));
  AOI22X1 g10171(.A0(n8981), .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B0(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(n8980), .Y(n13465));
  AOI22X1 g10172(.A0(n9000), .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B0(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(n8999), .Y(n13466));
  AOI22X1 g10173(.A0(n8987), .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B0(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(n8986), .Y(n13467));
  AOI22X1 g10174(.A0(n8984), .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B0(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(n8983), .Y(n13468));
  NAND4X1 g10175(.A(n13467), .B(n13466), .C(n13465), .D(n13468), .Y(n13469));
  NOR2X1  g10176(.A(n13469), .B(n13464), .Y(n13470));
  INVX1   g10177(.A(n13470), .Y(n13471));
  XOR2X1  g10178(.A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n8724), .Y(n13472));
  INVX1   g10179(.A(n13472), .Y(n13473));
  AOI21X1 g10180(.A0(n13473), .A1(n8926), .B0(n8722), .Y(n13474));
  OAI21X1 g10181(.A0(n13473), .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B0(n13474), .Y(n13475));
  AOI21X1 g10182(.A0(n13473), .A1(n8931), .B0(n8728), .Y(n13476));
  OAI21X1 g10183(.A0(n13473), .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B0(n13476), .Y(n13477));
  AOI21X1 g10184(.A0(n13473), .A1(n8934), .B0(n8733), .Y(n13478));
  OAI21X1 g10185(.A0(n13473), .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B0(n13478), .Y(n13479));
  AOI21X1 g10186(.A0(n13473), .A1(n8916), .B0(n8737), .Y(n13480));
  OAI21X1 g10187(.A0(n13473), .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B0(n13480), .Y(n13481));
  NAND4X1 g10188(.A(n13479), .B(n13477), .C(n13475), .D(n13481), .Y(n13482));
  NAND2X1 g10189(.A(n13472), .B(n9102), .Y(n13483));
  AOI21X1 g10190(.A0(n13473), .A1(n8919), .B0(n8742), .Y(n13484));
  NAND2X1 g10191(.A(n13484), .B(n13483), .Y(n13485));
  AOI21X1 g10192(.A0(n13473), .A1(n8923), .B0(n8746), .Y(n13486));
  OAI21X1 g10193(.A0(n13473), .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B0(n13486), .Y(n13487));
  AOI21X1 g10194(.A0(n13473), .A1(n8941), .B0(n8750), .Y(n13488));
  OAI21X1 g10195(.A0(n13473), .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B0(n13488), .Y(n13489));
  AOI21X1 g10196(.A0(n13473), .A1(n8938), .B0(n8754), .Y(n13490));
  OAI21X1 g10197(.A0(n13473), .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B0(n13490), .Y(n13491));
  NAND4X1 g10198(.A(n13489), .B(n13487), .C(n13485), .D(n13491), .Y(n13492));
  NOR2X1  g10199(.A(n13492), .B(n13482), .Y(n13493));
  XOR2X1  g10200(.A(n13493), .B(n13471), .Y(n13494));
  OAI22X1 g10201(.A0(n13470), .A1(n13459), .B0(n9760), .B1(n13494), .Y(n13495));
  NOR2X1  g10202(.A(n13493), .B(n13459), .Y(n13496));
  INVX1   g10203(.A(n13496), .Y(n13497));
  XOR2X1  g10204(.A(n13497), .B(n13495), .Y(n13498));
  XOR2X1  g10205(.A(n13498), .B(n13458), .Y(n13499));
  XOR2X1  g10206(.A(n13499), .B(n12221), .Y(n13500));
  XOR2X1  g10207(.A(n13500), .B(n13457), .Y(n13501));
  AOI22X1 g10208(.A0(n12998), .A1(P2_EAX_REG_23__SCAN_IN), .B0(n9744), .B1(n13304), .Y(n13502));
  OAI21X1 g10209(.A0(n13303), .A1(n9851), .B0(n13502), .Y(n13503));
  AOI21X1 g10210(.A0(n12999), .A1(n12222), .B0(n13503), .Y(n13504));
  OAI21X1 g10211(.A0(n13501), .A1(n13117), .B0(n13504), .Y(P2_U2896));
  NOR2X1  g10212(.A(n13499), .B(n12221), .Y(n13506));
  INVX1   g10213(.A(n13506), .Y(n13507));
  NAND2X1 g10214(.A(n13499), .B(n12221), .Y(n13508));
  INVX1   g10215(.A(n13508), .Y(n13509));
  OAI21X1 g10216(.A0(n13509), .A1(n13457), .B0(n13507), .Y(n13510));
  INVX1   g10217(.A(n13495), .Y(n13511));
  NOR2X1  g10218(.A(n13497), .B(n13511), .Y(n13512));
  NOR2X1  g10219(.A(n13496), .B(n13495), .Y(n13513));
  INVX1   g10220(.A(n13513), .Y(n13514));
  AOI21X1 g10221(.A0(n13514), .A1(n13458), .B0(n13512), .Y(n13515));
  INVX1   g10222(.A(n13515), .Y(n13516));
  NOR2X1  g10223(.A(n13493), .B(n13470), .Y(n13517));
  AOI21X1 g10224(.A0(n13473), .A1(n8957), .B0(n8722), .Y(n13518));
  OAI21X1 g10225(.A0(n13473), .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B0(n13518), .Y(n13519));
  AOI21X1 g10226(.A0(n13473), .A1(n8961), .B0(n8728), .Y(n13520));
  OAI21X1 g10227(.A0(n13473), .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B0(n13520), .Y(n13521));
  AOI21X1 g10228(.A0(n13473), .A1(n8964), .B0(n8733), .Y(n13522));
  OAI21X1 g10229(.A0(n13473), .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B0(n13522), .Y(n13523));
  AOI21X1 g10230(.A0(n13473), .A1(n8947), .B0(n8737), .Y(n13524));
  OAI21X1 g10231(.A0(n13473), .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B0(n13524), .Y(n13525));
  NAND4X1 g10232(.A(n13523), .B(n13521), .C(n13519), .D(n13525), .Y(n13526));
  NAND2X1 g10233(.A(n13472), .B(n9074), .Y(n13527));
  AOI21X1 g10234(.A0(n13473), .A1(n8950), .B0(n8742), .Y(n13528));
  NAND2X1 g10235(.A(n13528), .B(n13527), .Y(n13529));
  AOI21X1 g10236(.A0(n13473), .A1(n8954), .B0(n8746), .Y(n13530));
  OAI21X1 g10237(.A0(n13473), .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B0(n13530), .Y(n13531));
  AOI21X1 g10238(.A0(n13473), .A1(n8971), .B0(n8750), .Y(n13532));
  OAI21X1 g10239(.A0(n13473), .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B0(n13532), .Y(n13533));
  AOI21X1 g10240(.A0(n13473), .A1(n8968), .B0(n8754), .Y(n13534));
  OAI21X1 g10241(.A0(n13473), .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B0(n13534), .Y(n13535));
  NAND4X1 g10242(.A(n13533), .B(n13531), .C(n13529), .D(n13535), .Y(n13536));
  NOR2X1  g10243(.A(n13536), .B(n13526), .Y(n13537));
  XOR2X1  g10244(.A(n13537), .B(n13517), .Y(n13538));
  NOR2X1  g10245(.A(n13538), .B(n9760), .Y(n13539));
  NOR2X1  g10246(.A(n13537), .B(n13459), .Y(n13540));
  INVX1   g10247(.A(n13540), .Y(n13541));
  XOR2X1  g10248(.A(n13541), .B(n13539), .Y(n13542));
  XOR2X1  g10249(.A(n13542), .B(n13516), .Y(n13543));
  XOR2X1  g10250(.A(n13543), .B(n12258), .Y(n13544));
  XOR2X1  g10251(.A(n13544), .B(n13510), .Y(n13545));
  AOI22X1 g10252(.A0(n12998), .A1(P2_EAX_REG_24__SCAN_IN), .B0(n12842), .B1(n13304), .Y(n13546));
  OAI21X1 g10253(.A0(n13303), .A1(n9980), .B0(n13546), .Y(n13547));
  AOI21X1 g10254(.A0(n12999), .A1(n12258), .B0(n13547), .Y(n13548));
  OAI21X1 g10255(.A0(n13545), .A1(n13117), .B0(n13548), .Y(P2_U2895));
  NOR2X1  g10256(.A(n13543), .B(n12257), .Y(n13550));
  INVX1   g10257(.A(n13543), .Y(n13551));
  NOR2X1  g10258(.A(n13551), .B(n12258), .Y(n13552));
  INVX1   g10259(.A(n13552), .Y(n13553));
  AOI21X1 g10260(.A0(n13553), .A1(n13510), .B0(n13550), .Y(n13554));
  NOR4X1  g10261(.A(n13517), .B(n9760), .C(n13459), .D(n13537), .Y(n13555));
  NOR2X1  g10262(.A(n13542), .B(n13515), .Y(n13557));
  NOR2X1  g10263(.A(n13557), .B(n13555), .Y(n13558));
  NOR3X1  g10264(.A(n13537), .B(n13493), .C(n13470), .Y(n13559));
  AOI21X1 g10265(.A0(n13473), .A1(n8837), .B0(n8722), .Y(n13560));
  OAI21X1 g10266(.A0(n13473), .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B0(n13560), .Y(n13561));
  AOI21X1 g10267(.A0(n13473), .A1(n8841), .B0(n8728), .Y(n13562));
  OAI21X1 g10268(.A0(n13473), .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B0(n13562), .Y(n13563));
  AOI21X1 g10269(.A0(n13473), .A1(n8844), .B0(n8733), .Y(n13564));
  OAI21X1 g10270(.A0(n13473), .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B0(n13564), .Y(n13565));
  AOI21X1 g10271(.A0(n13473), .A1(n8827), .B0(n8737), .Y(n13566));
  OAI21X1 g10272(.A0(n13473), .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B0(n13566), .Y(n13567));
  NAND4X1 g10273(.A(n13565), .B(n13563), .C(n13561), .D(n13567), .Y(n13568));
  INVX1   g10274(.A(P2_INSTQUEUE_REG_3__2__SCAN_IN), .Y(n13569));
  NAND2X1 g10275(.A(n13472), .B(n13569), .Y(n13570));
  AOI21X1 g10276(.A0(n13473), .A1(n8830), .B0(n8742), .Y(n13571));
  NAND2X1 g10277(.A(n13571), .B(n13570), .Y(n13572));
  AOI21X1 g10278(.A0(n13473), .A1(n8834), .B0(n8746), .Y(n13573));
  OAI21X1 g10279(.A0(n13473), .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B0(n13573), .Y(n13574));
  AOI21X1 g10280(.A0(n13473), .A1(n8851), .B0(n8750), .Y(n13575));
  OAI21X1 g10281(.A0(n13473), .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B0(n13575), .Y(n13576));
  AOI21X1 g10282(.A0(n13473), .A1(n8848), .B0(n8754), .Y(n13577));
  OAI21X1 g10283(.A0(n13473), .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B0(n13577), .Y(n13578));
  NAND4X1 g10284(.A(n13576), .B(n13574), .C(n13572), .D(n13578), .Y(n13579));
  NOR2X1  g10285(.A(n13579), .B(n13568), .Y(n13580));
  XOR2X1  g10286(.A(n13580), .B(n13559), .Y(n13581));
  NOR2X1  g10287(.A(n13581), .B(n9760), .Y(n13582));
  NOR2X1  g10288(.A(n13580), .B(n13459), .Y(n13583));
  INVX1   g10289(.A(n13583), .Y(n13584));
  XOR2X1  g10290(.A(n13584), .B(n13582), .Y(n13585));
  INVX1   g10291(.A(n13585), .Y(n13586));
  XOR2X1  g10292(.A(n13586), .B(n13558), .Y(n13587));
  XOR2X1  g10293(.A(n13587), .B(n12296), .Y(n13588));
  XOR2X1  g10294(.A(n13588), .B(n13554), .Y(n13589));
  AOI22X1 g10295(.A0(n12998), .A1(P2_EAX_REG_25__SCAN_IN), .B0(n12836), .B1(n13304), .Y(n13590));
  OAI21X1 g10296(.A0(n13303), .A1(n9961), .B0(n13590), .Y(n13591));
  AOI21X1 g10297(.A0(n12999), .A1(n12297), .B0(n13591), .Y(n13592));
  OAI21X1 g10298(.A0(n13589), .A1(n13117), .B0(n13592), .Y(P2_U2894));
  NOR2X1  g10299(.A(n13587), .B(n12296), .Y(n13594));
  INVX1   g10300(.A(n13594), .Y(n13595));
  NAND2X1 g10301(.A(n13587), .B(n12296), .Y(n13596));
  INVX1   g10302(.A(n13596), .Y(n13597));
  OAI21X1 g10303(.A0(n13597), .A1(n13554), .B0(n13595), .Y(n13598));
  INVX1   g10304(.A(n12335), .Y(n13599));
  NOR4X1  g10305(.A(n13559), .B(n9760), .C(n13459), .D(n13580), .Y(n13600));
  NOR2X1  g10306(.A(n13585), .B(n13558), .Y(n13602));
  NOR2X1  g10307(.A(n13602), .B(n13600), .Y(n13603));
  NOR4X1  g10308(.A(n13537), .B(n13493), .C(n13470), .D(n13580), .Y(n13604));
  AOI21X1 g10309(.A0(n13473), .A1(n8895), .B0(n8722), .Y(n13605));
  OAI21X1 g10310(.A0(n13473), .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B0(n13605), .Y(n13606));
  AOI21X1 g10311(.A0(n13473), .A1(n8899), .B0(n8728), .Y(n13607));
  OAI21X1 g10312(.A0(n13473), .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B0(n13607), .Y(n13608));
  AOI21X1 g10313(.A0(n13473), .A1(n8902), .B0(n8733), .Y(n13609));
  OAI21X1 g10314(.A0(n13473), .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B0(n13609), .Y(n13610));
  AOI21X1 g10315(.A0(n13473), .A1(n8885), .B0(n8737), .Y(n13611));
  OAI21X1 g10316(.A0(n13473), .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B0(n13611), .Y(n13612));
  NAND4X1 g10317(.A(n13610), .B(n13608), .C(n13606), .D(n13612), .Y(n13613));
  NAND2X1 g10318(.A(n13472), .B(n11162), .Y(n13614));
  AOI21X1 g10319(.A0(n13473), .A1(n8888), .B0(n8742), .Y(n13615));
  NAND2X1 g10320(.A(n13615), .B(n13614), .Y(n13616));
  AOI21X1 g10321(.A0(n13473), .A1(n8892), .B0(n8746), .Y(n13617));
  OAI21X1 g10322(.A0(n13473), .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B0(n13617), .Y(n13618));
  AOI21X1 g10323(.A0(n13473), .A1(n8909), .B0(n8750), .Y(n13619));
  OAI21X1 g10324(.A0(n13473), .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B0(n13619), .Y(n13620));
  AOI21X1 g10325(.A0(n13473), .A1(n8906), .B0(n8754), .Y(n13621));
  OAI21X1 g10326(.A0(n13473), .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B0(n13621), .Y(n13622));
  NAND4X1 g10327(.A(n13620), .B(n13618), .C(n13616), .D(n13622), .Y(n13623));
  NOR2X1  g10328(.A(n13623), .B(n13613), .Y(n13624));
  XOR2X1  g10329(.A(n13624), .B(n13604), .Y(n13625));
  NOR2X1  g10330(.A(n13625), .B(n9760), .Y(n13626));
  NOR2X1  g10331(.A(n13624), .B(n13459), .Y(n13627));
  INVX1   g10332(.A(n13627), .Y(n13628));
  XOR2X1  g10333(.A(n13628), .B(n13626), .Y(n13629));
  INVX1   g10334(.A(n13629), .Y(n13630));
  XOR2X1  g10335(.A(n13630), .B(n13603), .Y(n13631));
  XOR2X1  g10336(.A(n13631), .B(n13599), .Y(n13632));
  XOR2X1  g10337(.A(n13632), .B(n13598), .Y(n13633));
  AOI22X1 g10338(.A0(n12998), .A1(P2_EAX_REG_26__SCAN_IN), .B0(n12830), .B1(n13304), .Y(n13634));
  OAI21X1 g10339(.A0(n13303), .A1(n9942), .B0(n13634), .Y(n13635));
  AOI21X1 g10340(.A0(n12999), .A1(n13599), .B0(n13635), .Y(n13636));
  OAI21X1 g10341(.A0(n13633), .A1(n13117), .B0(n13636), .Y(P2_U2893));
  NOR2X1  g10342(.A(n13631), .B(n12335), .Y(n13638));
  NAND2X1 g10343(.A(n13631), .B(n12335), .Y(n13639));
  AOI21X1 g10344(.A0(n13639), .A1(n13598), .B0(n13638), .Y(n13640));
  INVX1   g10345(.A(n13626), .Y(n13641));
  OAI22X1 g10346(.A0(n13626), .A1(n13627), .B0(n13602), .B1(n13600), .Y(n13642));
  OAI21X1 g10347(.A0(n13628), .A1(n13641), .B0(n13642), .Y(n13643));
  INVX1   g10348(.A(n13604), .Y(n13644));
  NOR2X1  g10349(.A(n13624), .B(n13644), .Y(n13645));
  AOI21X1 g10350(.A0(n13473), .A1(n9365), .B0(n8722), .Y(n13646));
  OAI21X1 g10351(.A0(n13473), .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B0(n13646), .Y(n13647));
  AOI21X1 g10352(.A0(n13473), .A1(n9368), .B0(n8728), .Y(n13648));
  OAI21X1 g10353(.A0(n13473), .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B0(n13648), .Y(n13649));
  AOI21X1 g10354(.A0(n13473), .A1(n9370), .B0(n8733), .Y(n13650));
  OAI21X1 g10355(.A0(n13473), .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B0(n13650), .Y(n13651));
  AOI21X1 g10356(.A0(n13473), .A1(n9358), .B0(n8737), .Y(n13652));
  OAI21X1 g10357(.A0(n13473), .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B0(n13652), .Y(n13653));
  NAND4X1 g10358(.A(n13651), .B(n13649), .C(n13647), .D(n13653), .Y(n13654));
  INVX1   g10359(.A(P2_INSTQUEUE_REG_3__4__SCAN_IN), .Y(n13655));
  NAND2X1 g10360(.A(n13472), .B(n13655), .Y(n13656));
  AOI21X1 g10361(.A0(n13473), .A1(n9360), .B0(n8742), .Y(n13657));
  NAND2X1 g10362(.A(n13657), .B(n13656), .Y(n13658));
  AOI21X1 g10363(.A0(n13473), .A1(n9363), .B0(n8746), .Y(n13659));
  OAI21X1 g10364(.A0(n13473), .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B0(n13659), .Y(n13660));
  AOI21X1 g10365(.A0(n13473), .A1(n9375), .B0(n8750), .Y(n13661));
  OAI21X1 g10366(.A0(n13473), .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B0(n13661), .Y(n13662));
  AOI21X1 g10367(.A0(n13473), .A1(n9373), .B0(n8754), .Y(n13663));
  OAI21X1 g10368(.A0(n13473), .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B0(n13663), .Y(n13664));
  NAND4X1 g10369(.A(n13662), .B(n13660), .C(n13658), .D(n13664), .Y(n13665));
  NOR2X1  g10370(.A(n13665), .B(n13654), .Y(n13666));
  XOR2X1  g10371(.A(n13666), .B(n13645), .Y(n13667));
  NOR2X1  g10372(.A(n13667), .B(n9760), .Y(n13668));
  NOR2X1  g10373(.A(n13666), .B(n13459), .Y(n13669));
  INVX1   g10374(.A(n13669), .Y(n13670));
  XOR2X1  g10375(.A(n13670), .B(n13668), .Y(n13671));
  XOR2X1  g10376(.A(n13671), .B(n13643), .Y(n13672));
  XOR2X1  g10377(.A(n13672), .B(n12371), .Y(n13673));
  XOR2X1  g10378(.A(n13673), .B(n13640), .Y(n13674));
  NOR2X1  g10379(.A(n13197), .B(n12371), .Y(n13675));
  AOI22X1 g10380(.A0(n12998), .A1(P2_EAX_REG_27__SCAN_IN), .B0(n12824), .B1(n13304), .Y(n13676));
  OAI21X1 g10381(.A0(n13303), .A1(n9923), .B0(n13676), .Y(n13677));
  NOR2X1  g10382(.A(n13677), .B(n13675), .Y(n13678));
  OAI21X1 g10383(.A0(n13674), .A1(n13117), .B0(n13678), .Y(P2_U2892));
  NOR2X1  g10384(.A(n13672), .B(n12371), .Y(n13680));
  INVX1   g10385(.A(n13680), .Y(n13681));
  NAND2X1 g10386(.A(n13672), .B(n12371), .Y(n13682));
  INVX1   g10387(.A(n13682), .Y(n13683));
  OAI21X1 g10388(.A0(n13683), .A1(n13640), .B0(n13681), .Y(n13684));
  NOR4X1  g10389(.A(n13645), .B(n9760), .C(n13459), .D(n13666), .Y(n13685));
  INVX1   g10390(.A(n13671), .Y(n13687));
  AOI21X1 g10391(.A0(n13687), .A1(n13643), .B0(n13685), .Y(n13688));
  NOR3X1  g10392(.A(n13666), .B(n13624), .C(n13644), .Y(n13689));
  AOI21X1 g10393(.A0(n13473), .A1(n8807), .B0(n8722), .Y(n13690));
  OAI21X1 g10394(.A0(n13473), .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B0(n13690), .Y(n13691));
  AOI21X1 g10395(.A0(n13473), .A1(n8811), .B0(n8728), .Y(n13692));
  OAI21X1 g10396(.A0(n13473), .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B0(n13692), .Y(n13693));
  AOI21X1 g10397(.A0(n13473), .A1(n8814), .B0(n8733), .Y(n13694));
  OAI21X1 g10398(.A0(n13473), .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B0(n13694), .Y(n13695));
  AOI21X1 g10399(.A0(n13473), .A1(n8797), .B0(n8737), .Y(n13696));
  OAI21X1 g10400(.A0(n13473), .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B0(n13696), .Y(n13697));
  NAND4X1 g10401(.A(n13695), .B(n13693), .C(n13691), .D(n13697), .Y(n13698));
  INVX1   g10402(.A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .Y(n13699));
  NAND2X1 g10403(.A(n13472), .B(n13699), .Y(n13700));
  AOI21X1 g10404(.A0(n13473), .A1(n8800), .B0(n8742), .Y(n13701));
  NAND2X1 g10405(.A(n13701), .B(n13700), .Y(n13702));
  AOI21X1 g10406(.A0(n13473), .A1(n8804), .B0(n8746), .Y(n13703));
  OAI21X1 g10407(.A0(n13473), .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B0(n13703), .Y(n13704));
  AOI21X1 g10408(.A0(n13473), .A1(n8821), .B0(n8750), .Y(n13705));
  OAI21X1 g10409(.A0(n13473), .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B0(n13705), .Y(n13706));
  AOI21X1 g10410(.A0(n13473), .A1(n8818), .B0(n8754), .Y(n13707));
  OAI21X1 g10411(.A0(n13473), .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B0(n13707), .Y(n13708));
  NAND4X1 g10412(.A(n13706), .B(n13704), .C(n13702), .D(n13708), .Y(n13709));
  NOR2X1  g10413(.A(n13709), .B(n13698), .Y(n13710));
  XOR2X1  g10414(.A(n13710), .B(n13689), .Y(n13711));
  NOR2X1  g10415(.A(n13711), .B(n9760), .Y(n13712));
  NOR2X1  g10416(.A(n13710), .B(n13459), .Y(n13713));
  XOR2X1  g10417(.A(n13713), .B(n13712), .Y(n13714));
  XOR2X1  g10418(.A(n13714), .B(n13688), .Y(n13715));
  XOR2X1  g10419(.A(n13715), .B(n12399), .Y(n13716));
  XOR2X1  g10420(.A(n13716), .B(n13684), .Y(n13717));
  AOI22X1 g10421(.A0(n12998), .A1(P2_EAX_REG_28__SCAN_IN), .B0(n12818), .B1(n13304), .Y(n13718));
  OAI21X1 g10422(.A0(n13303), .A1(n9904), .B0(n13718), .Y(n13719));
  AOI21X1 g10423(.A0(n12999), .A1(n12399), .B0(n13719), .Y(n13720));
  OAI21X1 g10424(.A0(n13717), .A1(n13117), .B0(n13720), .Y(P2_U2891));
  NOR4X1  g10425(.A(n13666), .B(n13624), .C(n13644), .D(n13710), .Y(n13722));
  AOI21X1 g10426(.A0(n13473), .A1(n8773), .B0(n8722), .Y(n13723));
  OAI21X1 g10427(.A0(n13473), .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B0(n13723), .Y(n13724));
  AOI21X1 g10428(.A0(n13473), .A1(n8780), .B0(n8728), .Y(n13725));
  OAI21X1 g10429(.A0(n13473), .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B0(n13725), .Y(n13726));
  AOI21X1 g10430(.A0(n13473), .A1(n8783), .B0(n8733), .Y(n13727));
  OAI21X1 g10431(.A0(n13473), .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B0(n13727), .Y(n13728));
  AOI21X1 g10432(.A0(n13473), .A1(n8761), .B0(n8737), .Y(n13729));
  OAI21X1 g10433(.A0(n13473), .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B0(n13729), .Y(n13730));
  NAND4X1 g10434(.A(n13728), .B(n13726), .C(n13724), .D(n13730), .Y(n13731));
  INVX1   g10435(.A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .Y(n13732));
  NAND2X1 g10436(.A(n13472), .B(n13732), .Y(n13733));
  AOI21X1 g10437(.A0(n13473), .A1(n8764), .B0(n8742), .Y(n13734));
  NAND2X1 g10438(.A(n13734), .B(n13733), .Y(n13735));
  AOI21X1 g10439(.A0(n13473), .A1(n8770), .B0(n8746), .Y(n13736));
  OAI21X1 g10440(.A0(n13473), .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B0(n13736), .Y(n13737));
  AOI21X1 g10441(.A0(n13473), .A1(n8792), .B0(n8750), .Y(n13738));
  OAI21X1 g10442(.A0(n13473), .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B0(n13738), .Y(n13739));
  AOI21X1 g10443(.A0(n13473), .A1(n8789), .B0(n8754), .Y(n13740));
  OAI21X1 g10444(.A0(n13473), .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B0(n13740), .Y(n13741));
  NAND4X1 g10445(.A(n13739), .B(n13737), .C(n13735), .D(n13741), .Y(n13742));
  NOR2X1  g10446(.A(n13742), .B(n13731), .Y(n13743));
  XOR2X1  g10447(.A(n13743), .B(n13722), .Y(n13744));
  NOR2X1  g10448(.A(n13744), .B(n9760), .Y(n13745));
  NOR2X1  g10449(.A(n13743), .B(n13459), .Y(n13746));
  INVX1   g10450(.A(n13746), .Y(n13747));
  XOR2X1  g10451(.A(n13747), .B(n13745), .Y(n13748));
  NOR4X1  g10452(.A(n13689), .B(n9760), .C(n13459), .D(n13710), .Y(n13749));
  INVX1   g10453(.A(n13749), .Y(n13750));
  NOR2X1  g10454(.A(n13713), .B(n13712), .Y(n13751));
  OAI21X1 g10455(.A0(n13751), .A1(n13688), .B0(n13750), .Y(n13752));
  XOR2X1  g10456(.A(n13752), .B(n13748), .Y(n13753));
  XOR2X1  g10457(.A(n13753), .B(n12442), .Y(n13754));
  NOR2X1  g10458(.A(n13715), .B(n12398), .Y(n13755));
  INVX1   g10459(.A(n13715), .Y(n13756));
  NOR2X1  g10460(.A(n13756), .B(n12399), .Y(n13757));
  INVX1   g10461(.A(n13757), .Y(n13758));
  AOI21X1 g10462(.A0(n13758), .A1(n13684), .B0(n13755), .Y(n13759));
  XOR2X1  g10463(.A(n13759), .B(n13754), .Y(n13760));
  INVX1   g10464(.A(n12442), .Y(n13761));
  AOI22X1 g10465(.A0(n12998), .A1(P2_EAX_REG_29__SCAN_IN), .B0(n12812), .B1(n13304), .Y(n13762));
  OAI21X1 g10466(.A0(n13303), .A1(n9885), .B0(n13762), .Y(n13763));
  AOI21X1 g10467(.A0(n12999), .A1(n13761), .B0(n13763), .Y(n13764));
  OAI21X1 g10468(.A0(n13760), .A1(n13117), .B0(n13764), .Y(P2_U2890));
  INVX1   g10469(.A(n13753), .Y(n13766));
  NAND2X1 g10470(.A(n13766), .B(n13761), .Y(n13767));
  INVX1   g10471(.A(n12476), .Y(n13768));
  NOR4X1  g10472(.A(n13722), .B(n9760), .C(n13459), .D(n13743), .Y(n13769));
  INVX1   g10473(.A(n13722), .Y(n13771));
  NOR2X1  g10474(.A(n13743), .B(n13771), .Y(n13772));
  NOR2X1  g10475(.A(n13473), .B(P2_INSTQUEUE_REG_2__7__SCAN_IN), .Y(n13773));
  OAI21X1 g10476(.A0(n13472), .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B0(n8759), .Y(n13774));
  NOR2X1  g10477(.A(n13473), .B(P2_INSTQUEUE_REG_7__7__SCAN_IN), .Y(n13775));
  OAI21X1 g10478(.A0(n13472), .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B0(n8760), .Y(n13776));
  OAI22X1 g10479(.A0(n13775), .A1(n13776), .B0(n13774), .B1(n13773), .Y(n13777));
  NOR2X1  g10480(.A(n13473), .B(P2_INSTQUEUE_REG_1__7__SCAN_IN), .Y(n13778));
  OAI21X1 g10481(.A0(n13472), .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B0(n8768), .Y(n13779));
  NOR2X1  g10482(.A(n13473), .B(P2_INSTQUEUE_REG_6__7__SCAN_IN), .Y(n13780));
  OAI21X1 g10483(.A0(n13472), .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B0(n8769), .Y(n13781));
  OAI22X1 g10484(.A0(n13780), .A1(n13781), .B0(n13779), .B1(n13778), .Y(n13782));
  NOR2X1  g10485(.A(n13782), .B(n13777), .Y(n13783));
  AOI21X1 g10486(.A0(n13473), .A1(n8859), .B0(n8742), .Y(n13784));
  OAI21X1 g10487(.A0(n13473), .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B0(n13784), .Y(n13785));
  AOI21X1 g10488(.A0(n13473), .A1(n8863), .B0(n8746), .Y(n13786));
  OAI21X1 g10489(.A0(n13473), .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B0(n13786), .Y(n13787));
  INVX1   g10490(.A(P2_INSTQUEUE_REG_4__7__SCAN_IN), .Y(n13788));
  OAI21X1 g10491(.A0(n13472), .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B0(n8787), .Y(n13789));
  AOI21X1 g10492(.A0(n13472), .A1(n13788), .B0(n13789), .Y(n13790));
  OAI21X1 g10493(.A0(n13472), .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B0(n8788), .Y(n13791));
  AOI21X1 g10494(.A0(n13472), .A1(n13110), .B0(n13791), .Y(n13792));
  NOR2X1  g10495(.A(n13792), .B(n13790), .Y(n13793));
  NAND4X1 g10496(.A(n13787), .B(n13785), .C(n13783), .D(n13793), .Y(n13794));
  XOR2X1  g10497(.A(n13794), .B(n13772), .Y(n13795));
  NAND2X1 g10498(.A(n13795), .B(n9785), .Y(n13796));
  NAND2X1 g10499(.A(n13794), .B(n9479), .Y(n13797));
  XOR2X1  g10500(.A(n13797), .B(n13796), .Y(n13798));
  INVX1   g10501(.A(n13798), .Y(n13799));
  NOR2X1  g10502(.A(n13799), .B(n13748), .Y(n13800));
  OAI21X1 g10503(.A0(n13769), .A1(n13752), .B0(n13800), .Y(n13801));
  INVX1   g10504(.A(n13801), .Y(n13802));
  INVX1   g10505(.A(n13748), .Y(n13803));
  AOI21X1 g10506(.A0(n13803), .A1(n13752), .B0(n13798), .Y(n13806));
  OAI21X1 g10507(.A0(n13806), .A1(n13802), .B0(n13768), .Y(n13807));
  INVX1   g10508(.A(n13806), .Y(n13808));
  NAND3X1 g10509(.A(n13808), .B(n13801), .C(n12476), .Y(n13809));
  NAND2X1 g10510(.A(n13809), .B(n13807), .Y(n13810));
  OAI21X1 g10511(.A0(n13766), .A1(n13761), .B0(n13810), .Y(n13811));
  AOI21X1 g10512(.A0(n13767), .A1(n13759), .B0(n13811), .Y(n13812));
  INVX1   g10513(.A(n13755), .Y(n13813));
  INVX1   g10514(.A(n13638), .Y(n13814));
  INVX1   g10515(.A(n13550), .Y(n13815));
  INVX1   g10516(.A(n13453), .Y(n13816));
  INVX1   g10517(.A(n13404), .Y(n13817));
  INVX1   g10518(.A(n13356), .Y(n13818));
  INVX1   g10519(.A(n13309), .Y(n13819));
  INVX1   g10520(.A(n13250), .Y(n13820));
  INVX1   g10521(.A(n13255), .Y(n13821));
  AOI21X1 g10522(.A0(n13820), .A1(n13240), .B0(n13821), .Y(n13822));
  OAI21X1 g10523(.A0(n13257), .A1(n13822), .B0(n13310), .Y(n13823));
  AOI21X1 g10524(.A0(n13823), .A1(n13819), .B0(n13334), .Y(n13824));
  OAI21X1 g10525(.A0(n13824), .A1(n13331), .B0(n13359), .Y(n13825));
  AOI21X1 g10526(.A0(n13825), .A1(n13818), .B0(n13383), .Y(n13826));
  OAI21X1 g10527(.A0(n13826), .A1(n13380), .B0(n13407), .Y(n13827));
  AOI21X1 g10528(.A0(n13827), .A1(n13817), .B0(n13432), .Y(n13828));
  OAI21X1 g10529(.A0(n13828), .A1(n13429), .B0(n13456), .Y(n13829));
  AOI21X1 g10530(.A0(n13829), .A1(n13816), .B0(n13509), .Y(n13830));
  OAI21X1 g10531(.A0(n13830), .A1(n13506), .B0(n13553), .Y(n13831));
  AOI21X1 g10532(.A0(n13831), .A1(n13815), .B0(n13597), .Y(n13832));
  OAI21X1 g10533(.A0(n13832), .A1(n13594), .B0(n13639), .Y(n13833));
  AOI21X1 g10534(.A0(n13833), .A1(n13814), .B0(n13683), .Y(n13834));
  OAI21X1 g10535(.A0(n13834), .A1(n13680), .B0(n13758), .Y(n13835));
  AOI22X1 g10536(.A0(n13813), .A1(n13835), .B0(n13753), .B1(n12442), .Y(n13836));
  NAND3X1 g10537(.A(n13809), .B(n13807), .C(n13767), .Y(n13837));
  OAI21X1 g10538(.A0(n13837), .A1(n13836), .B0(n13116), .Y(n13838));
  AOI22X1 g10539(.A0(n12998), .A1(P2_EAX_REG_30__SCAN_IN), .B0(n12805), .B1(n13304), .Y(n13839));
  OAI21X1 g10540(.A0(n13303), .A1(n9866), .B0(n13839), .Y(n13840));
  AOI21X1 g10541(.A0(n12999), .A1(n13768), .B0(n13840), .Y(n13841));
  OAI21X1 g10542(.A0(n13838), .A1(n13812), .B0(n13841), .Y(P2_U2889));
  NOR3X1  g10543(.A(n13195), .B(n9846), .C(n9470), .Y(n13843));
  AOI21X1 g10544(.A0(n12998), .A1(P2_EAX_REG_31__SCAN_IN), .B0(n13843), .Y(n13844));
  OAI21X1 g10545(.A0(n13197), .A1(n12519), .B0(n13844), .Y(P2_U2888));
  OAI21X1 g10546(.A0(n9639), .A1(n9413), .B0(n9724), .Y(n13846));
  NOR2X1  g10547(.A(n13846), .B(n8884), .Y(n13847));
  INVX1   g10548(.A(n13847), .Y(n13848));
  NOR2X1  g10549(.A(n13846), .B(n9339), .Y(n13849));
  AOI22X1 g10550(.A0(n13846), .A1(P2_EBX_REG_0__SCAN_IN), .B0(n9772), .B1(n13849), .Y(n13850));
  OAI21X1 g10551(.A0(n13848), .A1(n9614), .B0(n13850), .Y(P2_U2887));
  AOI22X1 g10552(.A0(n13846), .A1(P2_EBX_REG_1__SCAN_IN), .B0(n9996), .B1(n13849), .Y(n13852));
  OAI21X1 g10553(.A0(n13848), .A1(n9595), .B0(n13852), .Y(P2_U2886));
  AOI22X1 g10554(.A0(n13846), .A1(P2_EBX_REG_2__SCAN_IN), .B0(n9810), .B1(n13849), .Y(n13854));
  OAI21X1 g10555(.A0(n13848), .A1(n9633), .B0(n13854), .Y(P2_U2885));
  AOI22X1 g10556(.A0(n13846), .A1(P2_EBX_REG_3__SCAN_IN), .B0(n10350), .B1(n13849), .Y(n13856));
  OAI21X1 g10557(.A0(n13848), .A1(n9663), .B0(n13856), .Y(P2_U2884));
  AOI22X1 g10558(.A0(n13846), .A1(P2_EBX_REG_4__SCAN_IN), .B0(n13052), .B1(n13849), .Y(n13858));
  OAI21X1 g10559(.A0(n13848), .A1(n11251), .B0(n13858), .Y(P2_U2883));
  AOI22X1 g10560(.A0(n13846), .A1(P2_EBX_REG_5__SCAN_IN), .B0(n13076), .B1(n13849), .Y(n13860));
  OAI21X1 g10561(.A0(n13848), .A1(n11315), .B0(n13860), .Y(P2_U2882));
  INVX1   g10562(.A(n13849), .Y(n13862));
  AOI22X1 g10563(.A0(n13846), .A1(P2_EBX_REG_6__SCAN_IN), .B0(n12595), .B1(n13847), .Y(n13863));
  OAI21X1 g10564(.A0(n13862), .A1(n13095), .B0(n13863), .Y(P2_U2881));
  AOI22X1 g10565(.A0(n13846), .A1(P2_EBX_REG_7__SCAN_IN), .B0(n11430), .B1(n13847), .Y(n13865));
  OAI21X1 g10566(.A0(n13862), .A1(n13112), .B0(n13865), .Y(P2_U2880));
  AOI22X1 g10567(.A0(n13846), .A1(P2_EBX_REG_8__SCAN_IN), .B0(n12612), .B1(n13847), .Y(n13867));
  OAI21X1 g10568(.A0(n13862), .A1(n13169), .B0(n13867), .Y(P2_U2879));
  AOI22X1 g10569(.A0(n13846), .A1(P2_EBX_REG_9__SCAN_IN), .B0(n11565), .B1(n13847), .Y(n13869));
  OAI21X1 g10570(.A0(n13862), .A1(n13151), .B0(n13869), .Y(P2_U2878));
  AOI22X1 g10571(.A0(n13846), .A1(P2_EBX_REG_10__SCAN_IN), .B0(n12629), .B1(n13847), .Y(n13871));
  OAI21X1 g10572(.A0(n13862), .A1(n13172), .B0(n13871), .Y(P2_U2877));
  AOI22X1 g10573(.A0(n13846), .A1(P2_EBX_REG_11__SCAN_IN), .B0(n11666), .B1(n13847), .Y(n13873));
  OAI21X1 g10574(.A0(n13862), .A1(n13185), .B0(n13873), .Y(P2_U2876));
  AOI22X1 g10575(.A0(n13846), .A1(P2_EBX_REG_12__SCAN_IN), .B0(n11718), .B1(n13847), .Y(n13875));
  OAI21X1 g10576(.A0(n13862), .A1(n13206), .B0(n13875), .Y(P2_U2875));
  AOI22X1 g10577(.A0(n13846), .A1(P2_EBX_REG_13__SCAN_IN), .B0(n11773), .B1(n13847), .Y(n13877));
  OAI21X1 g10578(.A0(n13862), .A1(n13219), .B0(n13877), .Y(P2_U2874));
  AOI22X1 g10579(.A0(n13846), .A1(P2_EBX_REG_14__SCAN_IN), .B0(n11825), .B1(n13847), .Y(n13879));
  OAI21X1 g10580(.A0(n13862), .A1(n13237), .B0(n13879), .Y(P2_U2873));
  AOI22X1 g10581(.A0(n13846), .A1(P2_EBX_REG_15__SCAN_IN), .B0(n11874), .B1(n13847), .Y(n13881));
  OAI21X1 g10582(.A0(n13862), .A1(n13254), .B0(n13881), .Y(P2_U2872));
  AOI22X1 g10583(.A0(n13846), .A1(P2_EBX_REG_16__SCAN_IN), .B0(n11931), .B1(n13847), .Y(n13883));
  OAI21X1 g10584(.A0(n13862), .A1(n13299), .B0(n13883), .Y(P2_U2871));
  AOI22X1 g10585(.A0(n13846), .A1(P2_EBX_REG_17__SCAN_IN), .B0(n11969), .B1(n13847), .Y(n13885));
  OAI21X1 g10586(.A0(n13862), .A1(n13324), .B0(n13885), .Y(P2_U2870));
  AOI22X1 g10587(.A0(n13846), .A1(P2_EBX_REG_18__SCAN_IN), .B0(n12007), .B1(n13847), .Y(n13887));
  OAI21X1 g10588(.A0(n13862), .A1(n13349), .B0(n13887), .Y(P2_U2869));
  AOI22X1 g10589(.A0(n13846), .A1(P2_EBX_REG_19__SCAN_IN), .B0(n12048), .B1(n13847), .Y(n13889));
  OAI21X1 g10590(.A0(n13862), .A1(n13373), .B0(n13889), .Y(P2_U2868));
  AOI22X1 g10591(.A0(n13846), .A1(P2_EBX_REG_20__SCAN_IN), .B0(n12088), .B1(n13847), .Y(n13891));
  OAI21X1 g10592(.A0(n13862), .A1(n13397), .B0(n13891), .Y(P2_U2867));
  AOI22X1 g10593(.A0(n13846), .A1(P2_EBX_REG_21__SCAN_IN), .B0(n12126), .B1(n13847), .Y(n13893));
  OAI21X1 g10594(.A0(n13862), .A1(n13422), .B0(n13893), .Y(P2_U2866));
  AOI22X1 g10595(.A0(n13846), .A1(P2_EBX_REG_22__SCAN_IN), .B0(n12165), .B1(n13847), .Y(n13895));
  OAI21X1 g10596(.A0(n13862), .A1(n13446), .B0(n13895), .Y(P2_U2865));
  AOI22X1 g10597(.A0(n13846), .A1(P2_EBX_REG_23__SCAN_IN), .B0(n12211), .B1(n13847), .Y(n13897));
  OAI21X1 g10598(.A0(n13862), .A1(n13499), .B0(n13897), .Y(P2_U2864));
  AOI22X1 g10599(.A0(n13846), .A1(P2_EBX_REG_24__SCAN_IN), .B0(n12248), .B1(n13847), .Y(n13899));
  OAI21X1 g10600(.A0(n13862), .A1(n13543), .B0(n13899), .Y(P2_U2863));
  AOI22X1 g10601(.A0(n13846), .A1(P2_EBX_REG_25__SCAN_IN), .B0(n12287), .B1(n13847), .Y(n13901));
  OAI21X1 g10602(.A0(n13862), .A1(n13587), .B0(n13901), .Y(P2_U2862));
  AOI22X1 g10603(.A0(n13846), .A1(P2_EBX_REG_26__SCAN_IN), .B0(n12327), .B1(n13847), .Y(n13903));
  OAI21X1 g10604(.A0(n13862), .A1(n13631), .B0(n13903), .Y(P2_U2861));
  AOI22X1 g10605(.A0(n13846), .A1(P2_EBX_REG_27__SCAN_IN), .B0(n12361), .B1(n13847), .Y(n13905));
  OAI21X1 g10606(.A0(n13862), .A1(n13672), .B0(n13905), .Y(P2_U2860));
  AOI22X1 g10607(.A0(n13846), .A1(P2_EBX_REG_28__SCAN_IN), .B0(n12407), .B1(n13847), .Y(n13907));
  OAI21X1 g10608(.A0(n13862), .A1(n13715), .B0(n13907), .Y(P2_U2859));
  INVX1   g10609(.A(n12448), .Y(n13909));
  AOI22X1 g10610(.A0(n13846), .A1(P2_EBX_REG_29__SCAN_IN), .B0(n13909), .B1(n13847), .Y(n13910));
  OAI21X1 g10611(.A0(n13862), .A1(n13753), .B0(n13910), .Y(P2_U2858));
  NAND3X1 g10612(.A(n13849), .B(n13808), .C(n13801), .Y(n13912));
  INVX1   g10613(.A(n12482), .Y(n13913));
  AOI22X1 g10614(.A0(n13846), .A1(P2_EBX_REG_30__SCAN_IN), .B0(n13913), .B1(n13847), .Y(n13914));
  NAND2X1 g10615(.A(n13914), .B(n13912), .Y(P2_U2857));
  NAND2X1 g10616(.A(n13846), .B(P2_EBX_REG_31__SCAN_IN), .Y(n13916));
  OAI21X1 g10617(.A0(n13848), .A1(n12526), .B0(n13916), .Y(P2_U2856));
  AOI22X1 g10618(.A0(n9687), .A1(n9400), .B0(n10984), .B1(n9308), .Y(n13918));
  NOR2X1  g10619(.A(n13918), .B(n9732), .Y(n13919));
  NOR4X1  g10620(.A(n10965), .B(n9733), .C(n9723), .D(n13919), .Y(n13920));
  NOR4X1  g10621(.A(n9701), .B(n8979), .C(n9700), .D(n13920), .Y(n13921));
  INVX1   g10622(.A(n12892), .Y(n13922));
  OAI21X1 g10623(.A0(n9702), .A1(n13922), .B0(n12799), .Y(n13924));
  INVX1   g10624(.A(n13924), .Y(n13925));
  AOI21X1 g10625(.A0(n13921), .A1(n12522), .B0(n13925), .Y(n13926));
  NOR4X1  g10626(.A(n9702), .B(n8979), .C(n9700), .D(n13920), .Y(n13927));
  NAND2X1 g10627(.A(n13927), .B(n9752), .Y(n13928));
  INVX1   g10628(.A(n9195), .Y(n13929));
  NOR3X1  g10629(.A(n13920), .B(n9192), .C(n9205), .Y(n13930));
  NAND2X1 g10630(.A(n13930), .B(n13929), .Y(n13931));
  NOR2X1  g10631(.A(n13920), .B(n8719), .Y(n13932));
  AOI22X1 g10632(.A0(n13920), .A1(P2_REIP_REG_0__SCAN_IN), .B0(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B1(n13932), .Y(n13933));
  INVX1   g10633(.A(n9192), .Y(n13934));
  NOR3X1  g10634(.A(n13920), .B(n13934), .C(n9205), .Y(n13935));
  NOR3X1  g10635(.A(n13920), .B(n8978), .C(n9700), .Y(n13936));
  AOI22X1 g10636(.A0(n13935), .A1(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B0(n9772), .B1(n13936), .Y(n13937));
  NAND4X1 g10637(.A(n13933), .B(n13931), .C(n13928), .D(n13937), .Y(n13938));
  INVX1   g10638(.A(n13919), .Y(n13940));
  NOR4X1  g10639(.A(n9702), .B(n13922), .C(n8977), .D(n13940), .Y(n13941));
  INVX1   g10640(.A(n13941), .Y(n13942));
  NOR4X1  g10641(.A(n9701), .B(n8979), .C(n12522), .D(n13940), .Y(n13943));
  INVX1   g10642(.A(n13943), .Y(n13944));
  OAI22X1 g10643(.A0(n13942), .A1(n10960), .B0(n11005), .B1(n13944), .Y(n13945));
  NOR2X1  g10644(.A(n13945), .B(n13938), .Y(n13946));
  OAI21X1 g10645(.A0(n13926), .A1(n9532), .B0(n13946), .Y(P2_U2855));
  INVX1   g10646(.A(n13927), .Y(n13948));
  NOR2X1  g10647(.A(n13948), .B(n9595), .Y(n13949));
  INVX1   g10648(.A(n13930), .Y(n13950));
  AOI22X1 g10649(.A0(n13920), .A1(P2_REIP_REG_1__SCAN_IN), .B0(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(n13932), .Y(n13951));
  OAI21X1 g10650(.A0(n13950), .A1(n9201), .B0(n13951), .Y(n13952));
  INVX1   g10651(.A(n13935), .Y(n13953));
  INVX1   g10652(.A(n13936), .Y(n13954));
  OAI22X1 g10653(.A0(n13953), .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B0(n9784), .B1(n13954), .Y(n13955));
  OAI22X1 g10654(.A0(n13942), .A1(n10954), .B0(n11056), .B1(n13944), .Y(n13956));
  NOR4X1  g10655(.A(n13955), .B(n13952), .C(n13949), .D(n13956), .Y(n13957));
  OAI21X1 g10656(.A0(n13926), .A1(n9484), .B0(n13957), .Y(P2_U2854));
  INVX1   g10657(.A(n13926), .Y(n13959));
  NAND2X1 g10658(.A(n13959), .B(P2_EBX_REG_2__SCAN_IN), .Y(n13960));
  NOR2X1  g10659(.A(n10888), .B(n8720), .Y(n13961));
  AOI21X1 g10660(.A0(n12559), .A1(n8720), .B0(n13961), .Y(n13962));
  NOR2X1  g10661(.A(n9200), .B(n13929), .Y(n13963));
  XOR2X1  g10662(.A(n13963), .B(n13962), .Y(n13964));
  NAND2X1 g10663(.A(n13964), .B(n13930), .Y(n13965));
  AOI22X1 g10664(.A0(n13920), .A1(P2_REIP_REG_2__SCAN_IN), .B0(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(n13932), .Y(n13966));
  AOI22X1 g10665(.A0(n13935), .A1(n12559), .B0(n9810), .B1(n13936), .Y(n13967));
  NAND3X1 g10666(.A(n13967), .B(n13966), .C(n13965), .Y(n13968));
  AOI21X1 g10667(.A0(n13927), .A1(n9794), .B0(n13968), .Y(n13969));
  AOI22X1 g10668(.A0(n13941), .A1(n10940), .B0(n11106), .B1(n13943), .Y(n13970));
  NAND3X1 g10669(.A(n13970), .B(n13969), .C(n13960), .Y(P2_U2853));
  NAND2X1 g10670(.A(n13927), .B(n9815), .Y(n13972));
  NAND3X1 g10671(.A(n13962), .B(n9199), .C(n9195), .Y(n13973));
  NOR2X1  g10672(.A(n10929), .B(n8720), .Y(n13974));
  AOI21X1 g10673(.A0(n12566), .A1(n8720), .B0(n13974), .Y(n13975));
  INVX1   g10674(.A(n13975), .Y(n13976));
  XOR2X1  g10675(.A(n13976), .B(n13973), .Y(n13977));
  NAND2X1 g10676(.A(n13977), .B(n13930), .Y(n13978));
  AOI22X1 g10677(.A0(n13920), .A1(P2_REIP_REG_3__SCAN_IN), .B0(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(n13932), .Y(n13979));
  AOI22X1 g10678(.A0(n13935), .A1(n12566), .B0(n10350), .B1(n13936), .Y(n13980));
  NAND4X1 g10679(.A(n13979), .B(n13978), .C(n13972), .D(n13980), .Y(n13981));
  OAI22X1 g10680(.A0(n13942), .A1(n10933), .B0(n11151), .B1(n13944), .Y(n13982));
  NOR2X1  g10681(.A(n13982), .B(n13981), .Y(n13983));
  OAI21X1 g10682(.A0(n13926), .A1(n9658), .B0(n13983), .Y(P2_U2852));
  INVX1   g10683(.A(n13973), .Y(n13985));
  NOR2X1  g10684(.A(n11188), .B(n8720), .Y(n13986));
  NOR2X1  g10685(.A(n12574), .B(P2_STATE2_REG_0__SCAN_IN), .Y(n13987));
  NOR2X1  g10686(.A(n13987), .B(n13986), .Y(n13988));
  AOI21X1 g10687(.A0(n13975), .A1(n13985), .B0(n13988), .Y(n13989));
  NOR4X1  g10688(.A(n13986), .B(n13976), .C(n13973), .D(n13987), .Y(n13990));
  NOR3X1  g10689(.A(n13990), .B(n13989), .C(n13950), .Y(n13991));
  INVX1   g10690(.A(n13932), .Y(n13992));
  NOR3X1  g10691(.A(P2_STATE2_REG_1__SCAN_IN), .B(P2_STATE2_REG_2__SCAN_IN), .C(P2_STATE2_REG_3__SCAN_IN), .Y(n13993));
  INVX1   g10692(.A(n13993), .Y(n13994));
  AOI21X1 g10693(.A0(n13920), .A1(P2_REIP_REG_4__SCAN_IN), .B0(n10965), .Y(n13996));
  OAI21X1 g10694(.A0(n13992), .A1(n12572), .B0(n13996), .Y(n13997));
  OAI22X1 g10695(.A0(n13953), .A1(n12574), .B0(n13082), .B1(n13954), .Y(n13998));
  NOR3X1  g10696(.A(n13998), .B(n13997), .C(n13991), .Y(n13999));
  OAI21X1 g10697(.A0(n13948), .A1(n11251), .B0(n13999), .Y(n14000));
  OAI22X1 g10698(.A0(n13942), .A1(n13043), .B0(n11218), .B1(n13944), .Y(n14001));
  NOR2X1  g10699(.A(n14001), .B(n14000), .Y(n14002));
  OAI21X1 g10700(.A0(n13926), .A1(n11215), .B0(n14002), .Y(P2_U2851));
  NOR2X1  g10701(.A(n13948), .B(n11315), .Y(n14004));
  NOR2X1  g10702(.A(n11264), .B(n8720), .Y(n14005));
  AOI21X1 g10703(.A0(n12585), .A1(n8720), .B0(n14005), .Y(n14006));
  XOR2X1  g10704(.A(n14006), .B(n13990), .Y(n14007));
  NAND2X1 g10705(.A(n14007), .B(n13930), .Y(n14008));
  NAND2X1 g10706(.A(n13932), .B(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .Y(n14009));
  AOI21X1 g10707(.A0(n13920), .A1(P2_REIP_REG_5__SCAN_IN), .B0(n10965), .Y(n14010));
  AOI22X1 g10708(.A0(n13935), .A1(n12585), .B0(n13076), .B1(n13936), .Y(n14011));
  NAND4X1 g10709(.A(n14010), .B(n14009), .C(n14008), .D(n14011), .Y(n14012));
  OAI22X1 g10710(.A0(n13942), .A1(n11268), .B0(n11282), .B1(n13944), .Y(n14013));
  NOR3X1  g10711(.A(n14013), .B(n14012), .C(n14004), .Y(n14014));
  OAI21X1 g10712(.A0(n13926), .A1(n11278), .B0(n14014), .Y(P2_U2850));
  NAND2X1 g10713(.A(n13959), .B(P2_EBX_REG_6__SCAN_IN), .Y(n14016));
  NAND2X1 g10714(.A(n13935), .B(n12593), .Y(n14017));
  NOR2X1  g10715(.A(n11331), .B(n8720), .Y(n14018));
  AOI21X1 g10716(.A0(n12593), .A1(n8720), .B0(n14018), .Y(n14019));
  AOI21X1 g10717(.A0(n14006), .A1(n13990), .B0(n14019), .Y(n14020));
  NAND3X1 g10718(.A(n14019), .B(n14006), .C(n13990), .Y(n14021));
  INVX1   g10719(.A(n14021), .Y(n14022));
  NOR2X1  g10720(.A(n14022), .B(n14020), .Y(n14023));
  NAND2X1 g10721(.A(n14023), .B(n13930), .Y(n14024));
  NAND2X1 g10722(.A(n13932), .B(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .Y(n14025));
  AOI21X1 g10723(.A0(n13920), .A1(P2_REIP_REG_6__SCAN_IN), .B0(n10965), .Y(n14026));
  NAND4X1 g10724(.A(n14025), .B(n14024), .C(n14017), .D(n14026), .Y(n14027));
  AOI21X1 g10725(.A0(n13927), .A1(n12595), .B0(n14027), .Y(n14028));
  AOI22X1 g10726(.A0(n13941), .A1(n11335), .B0(n11352), .B1(n13943), .Y(n14029));
  NAND3X1 g10727(.A(n14029), .B(n14028), .C(n14016), .Y(P2_U2849));
  NAND2X1 g10728(.A(n13959), .B(P2_EBX_REG_7__SCAN_IN), .Y(n14031));
  NAND2X1 g10729(.A(n13935), .B(n12602), .Y(n14032));
  NOR2X1  g10730(.A(n11390), .B(n8720), .Y(n14033));
  AOI21X1 g10731(.A0(n12602), .A1(n8720), .B0(n14033), .Y(n14034));
  XOR2X1  g10732(.A(n14034), .B(n14022), .Y(n14035));
  NAND2X1 g10733(.A(n14035), .B(n13930), .Y(n14036));
  NAND2X1 g10734(.A(n13932), .B(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .Y(n14037));
  AOI21X1 g10735(.A0(n13920), .A1(P2_REIP_REG_7__SCAN_IN), .B0(n10965), .Y(n14038));
  NAND4X1 g10736(.A(n14037), .B(n14036), .C(n14032), .D(n14038), .Y(n14039));
  AOI21X1 g10737(.A0(n13927), .A1(n11430), .B0(n14039), .Y(n14040));
  AOI22X1 g10738(.A0(n13941), .A1(n11449), .B0(n11398), .B1(n13943), .Y(n14041));
  NAND3X1 g10739(.A(n14041), .B(n14040), .C(n14031), .Y(P2_U2848));
  NAND2X1 g10740(.A(n13959), .B(P2_EBX_REG_8__SCAN_IN), .Y(n14043));
  NAND2X1 g10741(.A(n13935), .B(n12610), .Y(n14044));
  NAND4X1 g10742(.A(n14019), .B(n14006), .C(n13990), .D(n14034), .Y(n14045));
  INVX1   g10743(.A(n14045), .Y(n14046));
  NOR2X1  g10744(.A(n11472), .B(n8720), .Y(n14047));
  AOI21X1 g10745(.A0(n12610), .A1(n8720), .B0(n14047), .Y(n14048));
  XOR2X1  g10746(.A(n14048), .B(n14046), .Y(n14049));
  NAND2X1 g10747(.A(n14049), .B(n13930), .Y(n14050));
  NAND2X1 g10748(.A(n13932), .B(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .Y(n14051));
  AOI21X1 g10749(.A0(n13920), .A1(P2_REIP_REG_8__SCAN_IN), .B0(n10965), .Y(n14052));
  NAND4X1 g10750(.A(n14051), .B(n14050), .C(n14044), .D(n14052), .Y(n14053));
  AOI21X1 g10751(.A0(n13927), .A1(n12612), .B0(n14053), .Y(n14054));
  AOI22X1 g10752(.A0(n13941), .A1(n11532), .B0(n11480), .B1(n13943), .Y(n14055));
  NAND3X1 g10753(.A(n14055), .B(n14054), .C(n14043), .Y(P2_U2847));
  NAND2X1 g10754(.A(n13959), .B(P2_EBX_REG_9__SCAN_IN), .Y(n14057));
  NAND2X1 g10755(.A(n13935), .B(n12617), .Y(n14058));
  NAND2X1 g10756(.A(n14048), .B(n14046), .Y(n14059));
  NOR2X1  g10757(.A(n11551), .B(n8720), .Y(n14060));
  AOI21X1 g10758(.A0(n12617), .A1(n8720), .B0(n14060), .Y(n14061));
  INVX1   g10759(.A(n14061), .Y(n14062));
  XOR2X1  g10760(.A(n14062), .B(n14059), .Y(n14063));
  NAND2X1 g10761(.A(n14063), .B(n13930), .Y(n14064));
  NAND2X1 g10762(.A(n13932), .B(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .Y(n14065));
  AOI21X1 g10763(.A0(n13920), .A1(P2_REIP_REG_9__SCAN_IN), .B0(n10965), .Y(n14066));
  NAND4X1 g10764(.A(n14065), .B(n14064), .C(n14058), .D(n14066), .Y(n14067));
  AOI21X1 g10765(.A0(n13927), .A1(n11565), .B0(n14067), .Y(n14068));
  INVX1   g10766(.A(n11547), .Y(n14069));
  AOI22X1 g10767(.A0(n13941), .A1(n11587), .B0(n14069), .B1(n13943), .Y(n14070));
  NAND3X1 g10768(.A(n14070), .B(n14068), .C(n14057), .Y(P2_U2846));
  NAND2X1 g10769(.A(n13959), .B(P2_EBX_REG_10__SCAN_IN), .Y(n14072));
  NAND2X1 g10770(.A(n13935), .B(n12627), .Y(n14073));
  NOR2X1  g10771(.A(n11594), .B(n8720), .Y(n14074));
  AOI21X1 g10772(.A0(n12627), .A1(n8720), .B0(n14074), .Y(n14075));
  INVX1   g10773(.A(n14075), .Y(n14076));
  OAI21X1 g10774(.A0(n14062), .A1(n14059), .B0(n14076), .Y(n14077));
  NOR3X1  g10775(.A(n14076), .B(n14062), .C(n14059), .Y(n14078));
  INVX1   g10776(.A(n14078), .Y(n14079));
  NAND3X1 g10777(.A(n14079), .B(n14077), .C(n13930), .Y(n14080));
  NAND2X1 g10778(.A(n13932), .B(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .Y(n14081));
  AOI21X1 g10779(.A0(n13920), .A1(P2_REIP_REG_10__SCAN_IN), .B0(n10965), .Y(n14082));
  NAND4X1 g10780(.A(n14081), .B(n14080), .C(n14073), .D(n14082), .Y(n14083));
  AOI21X1 g10781(.A0(n13927), .A1(n12629), .B0(n14083), .Y(n14084));
  AOI22X1 g10782(.A0(n13941), .A1(n13174), .B0(n11608), .B1(n13943), .Y(n14085));
  NAND3X1 g10783(.A(n14085), .B(n14084), .C(n14072), .Y(P2_U2845));
  NAND2X1 g10784(.A(n13959), .B(P2_EBX_REG_11__SCAN_IN), .Y(n14087));
  NOR2X1  g10785(.A(n11657), .B(n8720), .Y(n14088));
  AOI21X1 g10786(.A0(n12633), .A1(n8720), .B0(n14088), .Y(n14089));
  XOR2X1  g10787(.A(n14089), .B(n14079), .Y(n14090));
  NOR4X1  g10788(.A(n13920), .B(n9192), .C(n9205), .D(n14090), .Y(n14091));
  AOI21X1 g10789(.A0(n13920), .A1(P2_REIP_REG_11__SCAN_IN), .B0(n10965), .Y(n14092));
  OAI21X1 g10790(.A0(n13992), .A1(n9174), .B0(n14092), .Y(n14093));
  NOR2X1  g10791(.A(n14093), .B(n14091), .Y(n14094));
  OAI21X1 g10792(.A0(n13953), .A1(n12632), .B0(n14094), .Y(n14095));
  AOI21X1 g10793(.A0(n13927), .A1(n11666), .B0(n14095), .Y(n14096));
  INVX1   g10794(.A(n11652), .Y(n14097));
  AOI22X1 g10795(.A0(n13941), .A1(n11688), .B0(n14097), .B1(n13943), .Y(n14098));
  NAND3X1 g10796(.A(n14098), .B(n14096), .C(n14087), .Y(P2_U2844));
  NAND2X1 g10797(.A(n13959), .B(P2_EBX_REG_12__SCAN_IN), .Y(n14100));
  NAND2X1 g10798(.A(n13927), .B(n11718), .Y(n14101));
  NOR4X1  g10799(.A(n12640), .B(n13934), .C(n9205), .D(n13920), .Y(n14102));
  NAND2X1 g10800(.A(n14089), .B(n14078), .Y(n14103));
  NOR2X1  g10801(.A(n11704), .B(n8720), .Y(n14104));
  AOI21X1 g10802(.A0(n12641), .A1(n8720), .B0(n14104), .Y(n14105));
  XOR2X1  g10803(.A(n14105), .B(n14103), .Y(n14106));
  NOR4X1  g10804(.A(n13920), .B(n9192), .C(n9205), .D(n14106), .Y(n14107));
  AOI21X1 g10805(.A0(n13920), .A1(P2_REIP_REG_12__SCAN_IN), .B0(n10965), .Y(n14108));
  OAI21X1 g10806(.A0(n13992), .A1(n9175), .B0(n14108), .Y(n14109));
  NOR3X1  g10807(.A(n14109), .B(n14107), .C(n14102), .Y(n14110));
  AOI22X1 g10808(.A0(n13941), .A1(n11742), .B0(n11707), .B1(n13943), .Y(n14111));
  NAND4X1 g10809(.A(n14110), .B(n14101), .C(n14100), .D(n14111), .Y(P2_U2843));
  NAND2X1 g10810(.A(n13959), .B(P2_EBX_REG_13__SCAN_IN), .Y(n14113));
  INVX1   g10811(.A(n14105), .Y(n14114));
  NOR2X1  g10812(.A(n14114), .B(n14103), .Y(n14115));
  NOR2X1  g10813(.A(n11761), .B(n8720), .Y(n14116));
  AOI21X1 g10814(.A0(n12649), .A1(n8720), .B0(n14116), .Y(n14117));
  INVX1   g10815(.A(n14117), .Y(n14118));
  XOR2X1  g10816(.A(n14118), .B(n14115), .Y(n14119));
  NOR4X1  g10817(.A(n13920), .B(n9192), .C(n9205), .D(n14119), .Y(n14120));
  AOI21X1 g10818(.A0(n13920), .A1(P2_REIP_REG_13__SCAN_IN), .B0(n10965), .Y(n14121));
  OAI21X1 g10819(.A0(n13992), .A1(n9176), .B0(n14121), .Y(n14122));
  NOR2X1  g10820(.A(n14122), .B(n14120), .Y(n14123));
  OAI21X1 g10821(.A0(n13953), .A1(n12648), .B0(n14123), .Y(n14124));
  AOI21X1 g10822(.A0(n13927), .A1(n11773), .B0(n14124), .Y(n14125));
  INVX1   g10823(.A(n11757), .Y(n14126));
  AOI22X1 g10824(.A0(n13941), .A1(n11796), .B0(n14126), .B1(n13943), .Y(n14127));
  NAND3X1 g10825(.A(n14127), .B(n14125), .C(n14113), .Y(P2_U2842));
  NAND2X1 g10826(.A(n13959), .B(P2_EBX_REG_14__SCAN_IN), .Y(n14129));
  NAND2X1 g10827(.A(n13935), .B(n12655), .Y(n14130));
  NOR3X1  g10828(.A(n14118), .B(n14114), .C(n14103), .Y(n14131));
  NOR2X1  g10829(.A(n11810), .B(n8720), .Y(n14132));
  AOI21X1 g10830(.A0(n12655), .A1(n8720), .B0(n14132), .Y(n14133));
  XOR2X1  g10831(.A(n14133), .B(n14131), .Y(n14134));
  NAND2X1 g10832(.A(n14134), .B(n13930), .Y(n14135));
  NAND2X1 g10833(.A(n13932), .B(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .Y(n14136));
  AOI21X1 g10834(.A0(n13920), .A1(P2_REIP_REG_14__SCAN_IN), .B0(n10965), .Y(n14137));
  NAND4X1 g10835(.A(n14136), .B(n14135), .C(n14130), .D(n14137), .Y(n14138));
  AOI21X1 g10836(.A0(n13927), .A1(n11825), .B0(n14138), .Y(n14139));
  AOI22X1 g10837(.A0(n13941), .A1(n11848), .B0(n11812), .B1(n13943), .Y(n14140));
  NAND3X1 g10838(.A(n14140), .B(n14139), .C(n14129), .Y(P2_U2841));
  NAND2X1 g10839(.A(n13959), .B(P2_EBX_REG_15__SCAN_IN), .Y(n14142));
  NAND4X1 g10840(.A(n11896), .B(n9701), .C(n12892), .D(n12799), .Y(n14143));
  NOR2X1  g10841(.A(n11859), .B(n8720), .Y(n14144));
  AOI21X1 g10842(.A0(n12663), .A1(n8720), .B0(n14144), .Y(n14145));
  NAND3X1 g10843(.A(n14145), .B(n14133), .C(n14131), .Y(n14146));
  INVX1   g10844(.A(n14146), .Y(n14147));
  AOI21X1 g10845(.A0(n14133), .A1(n14131), .B0(n14145), .Y(n14148));
  NOR3X1  g10846(.A(n14148), .B(n14147), .C(n13950), .Y(n14149));
  NAND2X1 g10847(.A(n13935), .B(n12663), .Y(n14150));
  NAND2X1 g10848(.A(n13932), .B(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .Y(n14151));
  AOI21X1 g10849(.A0(n13920), .A1(P2_REIP_REG_15__SCAN_IN), .B0(n10965), .Y(n14152));
  NAND3X1 g10850(.A(n14152), .B(n14151), .C(n14150), .Y(n14153));
  NOR2X1  g10851(.A(n14153), .B(n14149), .Y(n14154));
  OAI21X1 g10852(.A0(n13944), .A1(n11864), .B0(n14154), .Y(n14155));
  AOI21X1 g10853(.A0(n13927), .A1(n11874), .B0(n14155), .Y(n14156));
  NAND3X1 g10854(.A(n14156), .B(n14143), .C(n14142), .Y(P2_U2840));
  NAND4X1 g10855(.A(n11942), .B(n9701), .C(n12892), .D(n12799), .Y(n14158));
  NAND2X1 g10856(.A(n13959), .B(P2_EBX_REG_16__SCAN_IN), .Y(n14159));
  NOR2X1  g10857(.A(n11919), .B(n8720), .Y(n14160));
  AOI21X1 g10858(.A0(n12671), .A1(n8720), .B0(n14160), .Y(n14161));
  XOR2X1  g10859(.A(n14161), .B(n14147), .Y(n14162));
  NAND2X1 g10860(.A(n13935), .B(n12671), .Y(n14163));
  NAND2X1 g10861(.A(n13932), .B(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .Y(n14164));
  AOI21X1 g10862(.A0(n13920), .A1(P2_REIP_REG_16__SCAN_IN), .B0(n10965), .Y(n14165));
  NAND3X1 g10863(.A(n14165), .B(n14164), .C(n14163), .Y(n14166));
  AOI21X1 g10864(.A0(n14162), .A1(n13930), .B0(n14166), .Y(n14167));
  OAI21X1 g10865(.A0(n13944), .A1(n11915), .B0(n14167), .Y(n14168));
  AOI21X1 g10866(.A0(n13927), .A1(n11931), .B0(n14168), .Y(n14169));
  NAND3X1 g10867(.A(n14169), .B(n14159), .C(n14158), .Y(P2_U2839));
  NOR2X1  g10868(.A(n13944), .B(n11958), .Y(n14171));
  NAND4X1 g10869(.A(n14145), .B(n14133), .C(n14131), .D(n14161), .Y(n14172));
  NOR2X1  g10870(.A(n11953), .B(n8720), .Y(n14173));
  AOI21X1 g10871(.A0(n12678), .A1(n8720), .B0(n14173), .Y(n14174));
  XOR2X1  g10872(.A(n14174), .B(n14172), .Y(n14175));
  NOR4X1  g10873(.A(n13920), .B(n9192), .C(n9205), .D(n14175), .Y(n14176));
  NOR4X1  g10874(.A(n12677), .B(n13934), .C(n9205), .D(n13920), .Y(n14177));
  AOI21X1 g10875(.A0(n13920), .A1(P2_REIP_REG_17__SCAN_IN), .B0(n10965), .Y(n14178));
  OAI21X1 g10876(.A0(n13992), .A1(n9171), .B0(n14178), .Y(n14179));
  NOR4X1  g10877(.A(n14177), .B(n14176), .C(n14171), .D(n14179), .Y(n14180));
  OAI21X1 g10878(.A0(n13926), .A1(n11964), .B0(n14180), .Y(n14181));
  AOI21X1 g10879(.A0(n13927), .A1(n11969), .B0(n14181), .Y(n14182));
  OAI21X1 g10880(.A0(n13942), .A1(n11979), .B0(n14182), .Y(P2_U2838));
  NAND4X1 g10881(.A(n12018), .B(n9701), .C(n12892), .D(n12799), .Y(n14184));
  NAND2X1 g10882(.A(n13927), .B(n12007), .Y(n14185));
  NAND3X1 g10883(.A(n14174), .B(n14161), .C(n14147), .Y(n14186));
  NOR2X1  g10884(.A(n12008), .B(n8720), .Y(n14187));
  AOI21X1 g10885(.A0(n12686), .A1(n8720), .B0(n14187), .Y(n14188));
  XOR2X1  g10886(.A(n14188), .B(n14186), .Y(n14189));
  NOR4X1  g10887(.A(n13920), .B(n9192), .C(n9205), .D(n14189), .Y(n14190));
  NOR4X1  g10888(.A(n12685), .B(n13934), .C(n9205), .D(n13920), .Y(n14191));
  AOI21X1 g10889(.A0(n13920), .A1(P2_REIP_REG_18__SCAN_IN), .B0(n10965), .Y(n14192));
  OAI21X1 g10890(.A0(n13992), .A1(n9172), .B0(n14192), .Y(n14193));
  NOR3X1  g10891(.A(n14193), .B(n14191), .C(n14190), .Y(n14194));
  OAI21X1 g10892(.A0(n13944), .A1(n11996), .B0(n14194), .Y(n14195));
  AOI21X1 g10893(.A0(n13959), .A1(P2_EBX_REG_18__SCAN_IN), .B0(n14195), .Y(n14196));
  NAND3X1 g10894(.A(n14196), .B(n14185), .C(n14184), .Y(P2_U2837));
  NAND4X1 g10895(.A(n12058), .B(n9701), .C(n12892), .D(n12799), .Y(n14198));
  NAND2X1 g10896(.A(n13927), .B(n12048), .Y(n14199));
  INVX1   g10897(.A(n14188), .Y(n14200));
  NOR2X1  g10898(.A(n14200), .B(n14186), .Y(n14201));
  NOR2X1  g10899(.A(n12028), .B(n8720), .Y(n14202));
  AOI21X1 g10900(.A0(n12694), .A1(n8720), .B0(n14202), .Y(n14203));
  INVX1   g10901(.A(n14203), .Y(n14204));
  XOR2X1  g10902(.A(n14204), .B(n14201), .Y(n14205));
  NOR4X1  g10903(.A(n13920), .B(n9192), .C(n9205), .D(n14205), .Y(n14206));
  NOR4X1  g10904(.A(n12693), .B(n13934), .C(n9205), .D(n13920), .Y(n14207));
  AOI21X1 g10905(.A0(n13920), .A1(P2_REIP_REG_19__SCAN_IN), .B0(n10965), .Y(n14208));
  OAI21X1 g10906(.A0(n13992), .A1(n9173), .B0(n14208), .Y(n14209));
  NOR3X1  g10907(.A(n14209), .B(n14207), .C(n14206), .Y(n14210));
  OAI21X1 g10908(.A0(n13944), .A1(n12033), .B0(n14210), .Y(n14211));
  AOI21X1 g10909(.A0(n13959), .A1(P2_EBX_REG_19__SCAN_IN), .B0(n14211), .Y(n14212));
  NAND3X1 g10910(.A(n14212), .B(n14199), .C(n14198), .Y(P2_U2836));
  NAND2X1 g10911(.A(n13935), .B(n12700), .Y(n14214));
  NOR3X1  g10912(.A(n14204), .B(n14200), .C(n14186), .Y(n14215));
  NOR2X1  g10913(.A(n12069), .B(n8720), .Y(n14216));
  AOI21X1 g10914(.A0(n12700), .A1(n8720), .B0(n14216), .Y(n14217));
  XOR2X1  g10915(.A(n14217), .B(n14215), .Y(n14218));
  NAND2X1 g10916(.A(n14218), .B(n13930), .Y(n14219));
  AOI22X1 g10917(.A0(n13920), .A1(P2_REIP_REG_20__SCAN_IN), .B0(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B1(n13932), .Y(n14220));
  NAND3X1 g10918(.A(n14220), .B(n14219), .C(n14214), .Y(n14221));
  AOI21X1 g10919(.A0(n13943), .A1(n12072), .B0(n14221), .Y(n14222));
  OAI21X1 g10920(.A0(n13926), .A1(n12083), .B0(n14222), .Y(n14223));
  AOI21X1 g10921(.A0(n13927), .A1(n12088), .B0(n14223), .Y(n14224));
  OAI21X1 g10922(.A0(n13942), .A1(n12097), .B0(n14224), .Y(P2_U2835));
  NOR2X1  g10923(.A(n13944), .B(n12115), .Y(n14226));
  NAND2X1 g10924(.A(n13935), .B(n12708), .Y(n14227));
  INVX1   g10925(.A(n14217), .Y(n14228));
  NOR4X1  g10926(.A(n14204), .B(n14200), .C(n14186), .D(n14228), .Y(n14229));
  NOR2X1  g10927(.A(n12110), .B(n8720), .Y(n14230));
  AOI21X1 g10928(.A0(n12708), .A1(n8720), .B0(n14230), .Y(n14231));
  XOR2X1  g10929(.A(n14231), .B(n14229), .Y(n14232));
  NAND2X1 g10930(.A(n14232), .B(n13930), .Y(n14233));
  AOI22X1 g10931(.A0(n13920), .A1(P2_REIP_REG_21__SCAN_IN), .B0(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .B1(n13932), .Y(n14234));
  NAND3X1 g10932(.A(n14234), .B(n14233), .C(n14227), .Y(n14235));
  NOR2X1  g10933(.A(n14235), .B(n14226), .Y(n14236));
  OAI21X1 g10934(.A0(n13926), .A1(n12121), .B0(n14236), .Y(n14237));
  AOI21X1 g10935(.A0(n13927), .A1(n12126), .B0(n14237), .Y(n14238));
  OAI21X1 g10936(.A0(n13942), .A1(n12137), .B0(n14238), .Y(P2_U2834));
  NOR2X1  g10937(.A(n13944), .B(n12151), .Y(n14240));
  NOR4X1  g10938(.A(n12715), .B(n13934), .C(n9205), .D(n13920), .Y(n14241));
  NAND2X1 g10939(.A(n14231), .B(n14229), .Y(n14242));
  NOR2X1  g10940(.A(n12155), .B(n8720), .Y(n14243));
  AOI21X1 g10941(.A0(n12716), .A1(n8720), .B0(n14243), .Y(n14244));
  XOR2X1  g10942(.A(n14244), .B(n14242), .Y(n14245));
  AOI22X1 g10943(.A0(n13920), .A1(P2_REIP_REG_22__SCAN_IN), .B0(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(n13932), .Y(n14246));
  OAI21X1 g10944(.A0(n14245), .A1(n13950), .B0(n14246), .Y(n14247));
  NOR3X1  g10945(.A(n14247), .B(n14241), .C(n14240), .Y(n14248));
  OAI21X1 g10946(.A0(n13926), .A1(n12160), .B0(n14248), .Y(n14249));
  AOI21X1 g10947(.A0(n13927), .A1(n12165), .B0(n14249), .Y(n14250));
  OAI21X1 g10948(.A0(n13942), .A1(n12175), .B0(n14250), .Y(P2_U2833));
  NAND4X1 g10949(.A(n12222), .B(n9701), .C(n12892), .D(n12799), .Y(n14252));
  NAND2X1 g10950(.A(n13927), .B(n12211), .Y(n14253));
  NAND3X1 g10951(.A(n14244), .B(n14231), .C(n14229), .Y(n14254));
  NOR2X1  g10952(.A(n12200), .B(n8720), .Y(n14255));
  AOI21X1 g10953(.A0(n12723), .A1(n8720), .B0(n14255), .Y(n14256));
  XOR2X1  g10954(.A(n14256), .B(n14254), .Y(n14257));
  NOR4X1  g10955(.A(n13920), .B(n9192), .C(n9205), .D(n14257), .Y(n14258));
  AOI22X1 g10956(.A0(n13920), .A1(P2_REIP_REG_23__SCAN_IN), .B0(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .B1(n13932), .Y(n14259));
  OAI21X1 g10957(.A0(n13953), .A1(n12722), .B0(n14259), .Y(n14260));
  NOR2X1  g10958(.A(n14260), .B(n14258), .Y(n14261));
  OAI21X1 g10959(.A0(n13944), .A1(n12195), .B0(n14261), .Y(n14262));
  AOI21X1 g10960(.A0(n13959), .A1(P2_EBX_REG_23__SCAN_IN), .B0(n14262), .Y(n14263));
  NAND3X1 g10961(.A(n14263), .B(n14253), .C(n14252), .Y(P2_U2832));
  NAND4X1 g10962(.A(n14244), .B(n14231), .C(n14229), .D(n14256), .Y(n14265));
  NOR2X1  g10963(.A(n12233), .B(n8720), .Y(n14266));
  AOI21X1 g10964(.A0(n12731), .A1(n8720), .B0(n14266), .Y(n14267));
  XOR2X1  g10965(.A(n14267), .B(n14265), .Y(n14268));
  INVX1   g10966(.A(n13920), .Y(n14269));
  OAI22X1 g10967(.A0(n14269), .A1(n8542), .B0(n9169), .B1(n13992), .Y(n14270));
  AOI21X1 g10968(.A0(n13935), .A1(n12731), .B0(n14270), .Y(n14271));
  OAI21X1 g10969(.A0(n14268), .A1(n13950), .B0(n14271), .Y(n14272));
  AOI21X1 g10970(.A0(n13943), .A1(n12236), .B0(n14272), .Y(n14273));
  OAI21X1 g10971(.A0(n13926), .A1(n12243), .B0(n14273), .Y(n14274));
  AOI21X1 g10972(.A0(n13927), .A1(n12248), .B0(n14274), .Y(n14275));
  OAI21X1 g10973(.A0(n13942), .A1(n12257), .B0(n14275), .Y(P2_U2831));
  INVX1   g10974(.A(n14267), .Y(n14277));
  NOR2X1  g10975(.A(n14277), .B(n14265), .Y(n14278));
  NOR2X1  g10976(.A(n12265), .B(n8720), .Y(n14279));
  AOI21X1 g10977(.A0(n12739), .A1(n8720), .B0(n14279), .Y(n14280));
  XOR2X1  g10978(.A(n14280), .B(n14278), .Y(n14281));
  OAI22X1 g10979(.A0(n14269), .A1(n8539), .B0(n9170), .B1(n13992), .Y(n14282));
  AOI21X1 g10980(.A0(n14281), .A1(n13930), .B0(n14282), .Y(n14283));
  OAI21X1 g10981(.A0(n13953), .A1(n12738), .B0(n14283), .Y(n14284));
  AOI21X1 g10982(.A0(n13959), .A1(P2_EBX_REG_25__SCAN_IN), .B0(n14284), .Y(n14285));
  OAI21X1 g10983(.A0(n13944), .A1(n12277), .B0(n14285), .Y(n14286));
  AOI21X1 g10984(.A0(n13927), .A1(n12287), .B0(n14286), .Y(n14287));
  OAI21X1 g10985(.A0(n13942), .A1(n12296), .B0(n14287), .Y(P2_U2830));
  NAND2X1 g10986(.A(n13935), .B(n12748), .Y(n14289));
  NAND2X1 g10987(.A(n14280), .B(n14278), .Y(n14290));
  NOR2X1  g10988(.A(n12315), .B(n8720), .Y(n14291));
  AOI21X1 g10989(.A0(n12748), .A1(n8720), .B0(n14291), .Y(n14292));
  INVX1   g10990(.A(n14292), .Y(n14293));
  XOR2X1  g10991(.A(n14293), .B(n14290), .Y(n14294));
  NAND2X1 g10992(.A(n14294), .B(n13930), .Y(n14295));
  AOI22X1 g10993(.A0(n13920), .A1(P2_REIP_REG_26__SCAN_IN), .B0(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .B1(n13932), .Y(n14296));
  NAND3X1 g10994(.A(n14296), .B(n14295), .C(n14289), .Y(n14297));
  AOI21X1 g10995(.A0(n13943), .A1(n12309), .B0(n14297), .Y(n14298));
  OAI21X1 g10996(.A0(n13926), .A1(n12323), .B0(n14298), .Y(n14299));
  AOI21X1 g10997(.A0(n13927), .A1(n12327), .B0(n14299), .Y(n14300));
  OAI21X1 g10998(.A0(n13942), .A1(n12335), .B0(n14300), .Y(P2_U2829));
  NAND3X1 g10999(.A(n14292), .B(n14280), .C(n14278), .Y(n14302));
  INVX1   g11000(.A(n12758), .Y(n14303));
  NOR2X1  g11001(.A(n12344), .B(n8720), .Y(n14304));
  AOI21X1 g11002(.A0(n14303), .A1(n8720), .B0(n14304), .Y(n14305));
  XOR2X1  g11003(.A(n14305), .B(n14302), .Y(n14306));
  NOR4X1  g11004(.A(n13920), .B(n9192), .C(n9205), .D(n14306), .Y(n14307));
  OAI22X1 g11005(.A0(n14269), .A1(n8533), .B0(n12756), .B1(n13992), .Y(n14308));
  NOR2X1  g11006(.A(n14308), .B(n14307), .Y(n14309));
  OAI21X1 g11007(.A0(n13953), .A1(n12758), .B0(n14309), .Y(n14310));
  AOI21X1 g11008(.A0(n13959), .A1(P2_EBX_REG_27__SCAN_IN), .B0(n14310), .Y(n14311));
  OAI21X1 g11009(.A0(n13944), .A1(n12349), .B0(n14311), .Y(n14312));
  AOI21X1 g11010(.A0(n13927), .A1(n12361), .B0(n14312), .Y(n14313));
  OAI21X1 g11011(.A0(n13942), .A1(n12371), .B0(n14313), .Y(P2_U2828));
  NAND2X1 g11012(.A(n13943), .B(n12386), .Y(n14315));
  NAND2X1 g11013(.A(n13959), .B(P2_EBX_REG_28__SCAN_IN), .Y(n14316));
  INVX1   g11014(.A(n12764), .Y(n14317));
  NAND2X1 g11015(.A(n13935), .B(n14317), .Y(n14318));
  NAND4X1 g11016(.A(n14292), .B(n14280), .C(n14278), .D(n14305), .Y(n14319));
  INVX1   g11017(.A(n14319), .Y(n14320));
  NOR2X1  g11018(.A(n12383), .B(n8720), .Y(n14321));
  AOI21X1 g11019(.A0(n14317), .A1(n8720), .B0(n14321), .Y(n14322));
  XOR2X1  g11020(.A(n14322), .B(n14320), .Y(n14323));
  OAI22X1 g11021(.A0(n14269), .A1(n8530), .B0(n12762), .B1(n13992), .Y(n14324));
  AOI21X1 g11022(.A0(n14323), .A1(n13930), .B0(n14324), .Y(n14325));
  NAND4X1 g11023(.A(n14318), .B(n14316), .C(n14315), .D(n14325), .Y(n14326));
  AOI21X1 g11024(.A0(n13927), .A1(n12407), .B0(n14326), .Y(n14327));
  OAI21X1 g11025(.A0(n13942), .A1(n12398), .B0(n14327), .Y(P2_U2827));
  NAND2X1 g11026(.A(n14322), .B(n14320), .Y(n14329));
  INVX1   g11027(.A(n12770), .Y(n14330));
  NOR2X1  g11028(.A(n12435), .B(n8720), .Y(n14331));
  AOI21X1 g11029(.A0(n14330), .A1(n8720), .B0(n14331), .Y(n14332));
  INVX1   g11030(.A(n14332), .Y(n14333));
  XOR2X1  g11031(.A(n14333), .B(n14329), .Y(n14334));
  OAI22X1 g11032(.A0(n14269), .A1(n8527), .B0(n9166), .B1(n13992), .Y(n14335));
  AOI21X1 g11033(.A0(n14334), .A1(n13930), .B0(n14335), .Y(n14336));
  OAI21X1 g11034(.A0(n13953), .A1(n12770), .B0(n14336), .Y(n14337));
  AOI21X1 g11035(.A0(n13959), .A1(P2_EBX_REG_29__SCAN_IN), .B0(n14337), .Y(n14338));
  OAI21X1 g11036(.A0(n13944), .A1(n12430), .B0(n14338), .Y(n14339));
  AOI21X1 g11037(.A0(n13927), .A1(n13909), .B0(n14339), .Y(n14340));
  OAI21X1 g11038(.A0(n13942), .A1(n12442), .B0(n14340), .Y(P2_U2826));
  NAND2X1 g11039(.A(n13943), .B(n12467), .Y(n14342));
  NAND2X1 g11040(.A(n13959), .B(P2_EBX_REG_30__SCAN_IN), .Y(n14343));
  INVX1   g11041(.A(n12777), .Y(n14344));
  NAND2X1 g11042(.A(n13935), .B(n14344), .Y(n14345));
  NOR2X1  g11043(.A(n14333), .B(n14329), .Y(n14346));
  NOR2X1  g11044(.A(n12472), .B(n8720), .Y(n14347));
  AOI21X1 g11045(.A0(n14344), .A1(n8720), .B0(n14347), .Y(n14348));
  XOR2X1  g11046(.A(n14348), .B(n14346), .Y(n14349));
  OAI22X1 g11047(.A0(n14269), .A1(n8522), .B0(n9167), .B1(n13992), .Y(n14350));
  AOI21X1 g11048(.A0(n14349), .A1(n13930), .B0(n14350), .Y(n14351));
  NAND4X1 g11049(.A(n14345), .B(n14343), .C(n14342), .D(n14351), .Y(n14352));
  AOI21X1 g11050(.A0(n13927), .A1(n13913), .B0(n14352), .Y(n14353));
  OAI21X1 g11051(.A0(n13942), .A1(n12476), .B0(n14353), .Y(P2_U2825));
  NOR2X1  g11052(.A(n13948), .B(n12526), .Y(n14355));
  NAND2X1 g11053(.A(n13935), .B(n9191), .Y(n14356));
  NAND4X1 g11054(.A(n14346), .B(n9723), .C(n13934), .D(n14348), .Y(n14358));
  AOI22X1 g11055(.A0(n13920), .A1(P2_REIP_REG_31__SCAN_IN), .B0(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B1(n13932), .Y(n14359));
  NAND3X1 g11056(.A(n14359), .B(n14358), .C(n14356), .Y(n14360));
  AOI21X1 g11057(.A0(n13959), .A1(P2_EBX_REG_31__SCAN_IN), .B0(n14360), .Y(n14361));
  OAI21X1 g11058(.A0(n13944), .A1(n12497), .B0(n14361), .Y(n14362));
  NOR2X1  g11059(.A(n14362), .B(n14355), .Y(n14363));
  OAI21X1 g11060(.A0(n13942), .A1(n12519), .B0(n14363), .Y(P2_U2824));
  NOR4X1  g11061(.A(P2_DATAWIDTH_REG_15__SCAN_IN), .B(P2_DATAWIDTH_REG_14__SCAN_IN), .C(P2_DATAWIDTH_REG_13__SCAN_IN), .D(P2_DATAWIDTH_REG_16__SCAN_IN), .Y(n14365));
  NOR4X1  g11062(.A(P2_DATAWIDTH_REG_12__SCAN_IN), .B(P2_DATAWIDTH_REG_11__SCAN_IN), .C(P2_DATAWIDTH_REG_10__SCAN_IN), .D(P2_DATAWIDTH_REG_26__SCAN_IN), .Y(n14366));
  NOR4X1  g11063(.A(P2_DATAWIDTH_REG_7__SCAN_IN), .B(P2_DATAWIDTH_REG_6__SCAN_IN), .C(P2_DATAWIDTH_REG_5__SCAN_IN), .D(P2_DATAWIDTH_REG_8__SCAN_IN), .Y(n14367));
  NOR4X1  g11064(.A(P2_DATAWIDTH_REG_4__SCAN_IN), .B(P2_DATAWIDTH_REG_3__SCAN_IN), .C(P2_DATAWIDTH_REG_2__SCAN_IN), .D(P2_DATAWIDTH_REG_17__SCAN_IN), .Y(n14368));
  NAND4X1 g11065(.A(n14367), .B(n14366), .C(n14365), .D(n14368), .Y(n14369));
  NOR4X1  g11066(.A(P2_DATAWIDTH_REG_22__SCAN_IN), .B(P2_DATAWIDTH_REG_21__SCAN_IN), .C(P2_DATAWIDTH_REG_20__SCAN_IN), .D(P2_DATAWIDTH_REG_23__SCAN_IN), .Y(n14370));
  INVX1   g11067(.A(P2_DATAWIDTH_REG_0__SCAN_IN), .Y(n14371));
  NOR2X1  g11068(.A(n8655), .B(n14371), .Y(n14372));
  NOR3X1  g11069(.A(n14372), .B(P2_DATAWIDTH_REG_19__SCAN_IN), .C(P2_DATAWIDTH_REG_18__SCAN_IN), .Y(n14373));
  NOR4X1  g11070(.A(P2_DATAWIDTH_REG_29__SCAN_IN), .B(P2_DATAWIDTH_REG_28__SCAN_IN), .C(P2_DATAWIDTH_REG_27__SCAN_IN), .D(P2_DATAWIDTH_REG_30__SCAN_IN), .Y(n14374));
  NOR4X1  g11071(.A(P2_DATAWIDTH_REG_25__SCAN_IN), .B(P2_DATAWIDTH_REG_24__SCAN_IN), .C(P2_DATAWIDTH_REG_9__SCAN_IN), .D(P2_DATAWIDTH_REG_31__SCAN_IN), .Y(n14375));
  NAND4X1 g11072(.A(n14374), .B(n14373), .C(n14370), .D(n14375), .Y(n14376));
  NOR2X1  g11073(.A(n14376), .B(n14369), .Y(n14377));
  NAND3X1 g11074(.A(n14377), .B(n8611), .C(n8655), .Y(n14378));
  NAND4X1 g11075(.A(n9582), .B(n8655), .C(n14371), .D(n14377), .Y(n14379));
  OAI21X1 g11076(.A0(n14376), .A1(n14369), .B0(P2_BYTEENABLE_REG_3__SCAN_IN), .Y(n14380));
  NAND3X1 g11077(.A(n14380), .B(n14379), .C(n14378), .Y(P2_U2823));
  NAND2X1 g11078(.A(n14377), .B(P2_REIP_REG_1__SCAN_IN), .Y(n14382));
  NAND2X1 g11079(.A(n8611), .B(n8655), .Y(n14383));
  AOI21X1 g11080(.A0(P2_REIP_REG_0__SCAN_IN), .A1(P2_DATAWIDTH_REG_0__SCAN_IN), .B0(n14383), .Y(n14384));
  NOR2X1  g11081(.A(n14377), .B(n8511), .Y(n14385));
  AOI21X1 g11082(.A0(n14384), .A1(n14377), .B0(n14385), .Y(n14386));
  OAI21X1 g11083(.A0(n14382), .A1(n9582), .B0(n14386), .Y(P2_U2822));
  OAI21X1 g11084(.A0(n14376), .A1(n14369), .B0(P2_BYTEENABLE_REG_1__SCAN_IN), .Y(n14388));
  NAND3X1 g11085(.A(n14388), .B(n14382), .C(n14379), .Y(P2_U2821));
  NAND2X1 g11086(.A(n14377), .B(P2_REIP_REG_0__SCAN_IN), .Y(n14390));
  OAI21X1 g11087(.A0(n14376), .A1(n14369), .B0(P2_BYTEENABLE_REG_0__SCAN_IN), .Y(n14391));
  NAND3X1 g11088(.A(n14391), .B(n14390), .C(n14382), .Y(P2_U2820));
  INVX1   g11089(.A(P2_READREQUEST_REG_SCAN_IN), .Y(n14393));
  NAND3X1 g11090(.A(n14393), .B(n8506), .C(P2_STATE_REG_1__SCAN_IN), .Y(n14394));
  OAI21X1 g11091(.A0(n8512), .A1(n3087), .B0(n14394), .Y(P2_U3608));
  NOR2X1  g11092(.A(n9732), .B(n9694), .Y(n14396));
  NOR2X1  g11093(.A(n9259), .B(n9022), .Y(n14397));
  NOR3X1  g11094(.A(n12793), .B(n9262), .C(n9404), .Y(n14398));
  OAI21X1 g11095(.A0(n9161), .A1(n8975), .B0(n14398), .Y(n14399));
  OAI22X1 g11096(.A0(n14397), .A1(n14399), .B0(n14396), .B1(n9162), .Y(P2_U2819));
  OAI21X1 g11097(.A0(n9732), .A1(n9694), .B0(P2_MORE_REG_SCAN_IN), .Y(n14401));
  NAND2X1 g11098(.A(n14396), .B(n9403), .Y(n14402));
  NAND2X1 g11099(.A(n14402), .B(n14401), .Y(P2_U3609));
  AOI22X1 g11100(.A0(n8628), .A1(n8506), .B0(P2_STATEBS16_REG_SCAN_IN), .B1(n8652), .Y(n14404));
  OAI21X1 g11101(.A0(n8652), .A1(n3439), .B0(n14404), .Y(P2_U2818));
  AOI21X1 g11102(.A0(n9486), .A1(n9278), .B0(n8620), .Y(n14406));
  NOR4X1  g11103(.A(n9022), .B(n8978), .C(n8720), .D(n9418), .Y(n14407));
  NOR3X1  g11104(.A(n9417), .B(n9710), .C(P2_STATE_REG_0__SCAN_IN), .Y(n14408));
  NOR3X1  g11105(.A(n14408), .B(n9262), .C(n8975), .Y(n14409));
  AOI21X1 g11106(.A0(n8720), .A1(P2_STATE2_REG_1__SCAN_IN), .B0(P2_STATE2_REG_2__SCAN_IN), .Y(n14410));
  NOR4X1  g11107(.A(n14409), .B(n14407), .C(n14406), .D(n14410), .Y(n14411));
  NOR4X1  g11108(.A(P2_STATE2_REG_0__SCAN_IN), .B(n9205), .C(n9700), .D(n8619), .Y(n14412));
  OAI21X1 g11109(.A0(n10857), .A1(P2_STATE2_REG_0__SCAN_IN), .B0(n9767), .Y(n14413));
  NOR3X1  g11110(.A(n14413), .B(n14412), .C(n13919), .Y(n14414));
  NAND2X1 g11111(.A(n14414), .B(P2_REQUESTPENDING_REG_SCAN_IN), .Y(n14415));
  OAI21X1 g11112(.A0(n14414), .A1(n14411), .B0(n14415), .Y(P2_U3610));
  OAI21X1 g11113(.A0(P2_STATE_REG_0__SCAN_IN), .A1(n8508), .B0(P2_D_C_N_REG_SCAN_IN), .Y(n14417));
  NOR3X1  g11114(.A(P2_CODEFETCH_REG_SCAN_IN), .B(P2_STATE_REG_0__SCAN_IN), .C(n8508), .Y(n14418));
  AOI21X1 g11115(.A0(n8628), .A1(n8506), .B0(n14418), .Y(n14419));
  NAND2X1 g11116(.A(n14419), .B(n14417), .Y(P2_U2817));
  NAND3X1 g11117(.A(P2_MEMORYFETCH_REG_SCAN_IN), .B(n8506), .C(P2_STATE_REG_1__SCAN_IN), .Y(n14421));
  OAI21X1 g11118(.A0(n8512), .A1(n3089), .B0(n14421), .Y(P2_U3611));
  OAI21X1 g11119(.A0(n9732), .A1(n13918), .B0(P2_CODEFETCH_REG_SCAN_IN), .Y(n14423));
  OAI21X1 g11120(.A0(n13994), .A1(n8720), .B0(n14423), .Y(P2_U2816));
  NAND2X1 g11121(.A(P2_ADS_N_REG_SCAN_IN), .B(P2_STATE_REG_0__SCAN_IN), .Y(n14425));
  NAND2X1 g11122(.A(n14425), .B(n8652), .Y(P2_U2815));
  OAI21X1 g11123(.A0(n13918), .A1(n9732), .B0(n13994), .Y(n14427));
  OAI21X1 g11124(.A0(n9458), .A1(n9700), .B0(n14427), .Y(n14428));
  OAI21X1 g11125(.A0(n14427), .A1(n14393), .B0(n14428), .Y(P2_U3612));
  AOI21X1 g11126(.A0(n9356), .A1(n9230), .B0(n8975), .Y(n14430));
  NOR3X1  g11127(.A(n14430), .B(n12793), .C(n9478), .Y(n14431));
  OAI21X1 g11128(.A0(n9308), .A1(n9022), .B0(n14431), .Y(n14432));
  NAND2X1 g11129(.A(n14432), .B(P2_MEMORYFETCH_REG_SCAN_IN), .Y(n14433));
  NAND3X1 g11130(.A(n9724), .B(n12791), .C(n8978), .Y(n14434));
  NAND3X1 g11131(.A(n14434), .B(n14433), .C(n13994), .Y(P2_U2814));
  INVX1   g11132(.A(P1_STATE_REG_0__SCAN_IN), .Y(n14436));
  NAND3X1 g11133(.A(n14436), .B(P1_STATE_REG_1__SCAN_IN), .C(P1_BYTEENABLE_REG_3__SCAN_IN), .Y(n14437));
  INVX1   g11134(.A(P1_STATE_REG_1__SCAN_IN), .Y(n14438));
  OAI21X1 g11135(.A0(P1_STATE_REG_0__SCAN_IN), .A1(n14438), .B0(P1_BE_N_REG_3__SCAN_IN), .Y(n14439));
  NAND2X1 g11136(.A(n14439), .B(n14437), .Y(P1_U3458));
  INVX1   g11137(.A(P1_BYTEENABLE_REG_2__SCAN_IN), .Y(n14441));
  NOR2X1  g11138(.A(P1_STATE_REG_0__SCAN_IN), .B(n14438), .Y(n14442));
  INVX1   g11139(.A(n14442), .Y(n14443));
  OAI21X1 g11140(.A0(P1_STATE_REG_0__SCAN_IN), .A1(n14438), .B0(P1_BE_N_REG_2__SCAN_IN), .Y(n14444));
  OAI21X1 g11141(.A0(n14443), .A1(n14441), .B0(n14444), .Y(P1_U3459));
  NAND3X1 g11142(.A(n14436), .B(P1_STATE_REG_1__SCAN_IN), .C(P1_BYTEENABLE_REG_1__SCAN_IN), .Y(n14446));
  OAI21X1 g11143(.A0(P1_STATE_REG_0__SCAN_IN), .A1(n14438), .B0(P1_BE_N_REG_1__SCAN_IN), .Y(n14447));
  NAND2X1 g11144(.A(n14447), .B(n14446), .Y(P1_U3460));
  INVX1   g11145(.A(P1_BYTEENABLE_REG_0__SCAN_IN), .Y(n14449));
  OAI21X1 g11146(.A0(P1_STATE_REG_0__SCAN_IN), .A1(n14438), .B0(P1_BE_N_REG_0__SCAN_IN), .Y(n14450));
  OAI21X1 g11147(.A0(n14443), .A1(n14449), .B0(n14450), .Y(P1_U3461));
  INVX1   g11148(.A(P1_REIP_REG_30__SCAN_IN), .Y(n14452));
  NAND3X1 g11149(.A(n14436), .B(P1_STATE_REG_1__SCAN_IN), .C(P1_STATE_REG_2__SCAN_IN), .Y(n14453));
  NOR3X1  g11150(.A(P1_STATE_REG_0__SCAN_IN), .B(n14438), .C(P1_STATE_REG_2__SCAN_IN), .Y(n14454));
  AOI22X1 g11151(.A0(n14443), .A1(P1_ADDRESS_REG_29__SCAN_IN), .B0(P1_REIP_REG_31__SCAN_IN), .B1(n14454), .Y(n14455));
  OAI21X1 g11152(.A0(n14453), .A1(n14452), .B0(n14455), .Y(P1_U3226));
  INVX1   g11153(.A(P1_REIP_REG_29__SCAN_IN), .Y(n14457));
  AOI22X1 g11154(.A0(n14443), .A1(P1_ADDRESS_REG_28__SCAN_IN), .B0(P1_REIP_REG_30__SCAN_IN), .B1(n14454), .Y(n14458));
  OAI21X1 g11155(.A0(n14453), .A1(n14457), .B0(n14458), .Y(P1_U3225));
  INVX1   g11156(.A(P1_REIP_REG_28__SCAN_IN), .Y(n14460));
  AOI22X1 g11157(.A0(n14443), .A1(P1_ADDRESS_REG_27__SCAN_IN), .B0(P1_REIP_REG_29__SCAN_IN), .B1(n14454), .Y(n14461));
  OAI21X1 g11158(.A0(n14453), .A1(n14460), .B0(n14461), .Y(P1_U3224));
  INVX1   g11159(.A(P1_REIP_REG_27__SCAN_IN), .Y(n14463));
  AOI22X1 g11160(.A0(n14443), .A1(P1_ADDRESS_REG_26__SCAN_IN), .B0(P1_REIP_REG_28__SCAN_IN), .B1(n14454), .Y(n14464));
  OAI21X1 g11161(.A0(n14453), .A1(n14463), .B0(n14464), .Y(P1_U3223));
  NAND4X1 g11162(.A(P1_STATE_REG_1__SCAN_IN), .B(P1_STATE_REG_2__SCAN_IN), .C(P1_REIP_REG_26__SCAN_IN), .D(n14436), .Y(n14466));
  AOI22X1 g11163(.A0(n14443), .A1(P1_ADDRESS_REG_25__SCAN_IN), .B0(P1_REIP_REG_27__SCAN_IN), .B1(n14454), .Y(n14467));
  NAND2X1 g11164(.A(n14467), .B(n14466), .Y(P1_U3222));
  INVX1   g11165(.A(P1_REIP_REG_25__SCAN_IN), .Y(n14469));
  AOI22X1 g11166(.A0(n14443), .A1(P1_ADDRESS_REG_24__SCAN_IN), .B0(P1_REIP_REG_26__SCAN_IN), .B1(n14454), .Y(n14470));
  OAI21X1 g11167(.A0(n14453), .A1(n14469), .B0(n14470), .Y(P1_U3221));
  INVX1   g11168(.A(P1_REIP_REG_24__SCAN_IN), .Y(n14472));
  AOI22X1 g11169(.A0(n14443), .A1(P1_ADDRESS_REG_23__SCAN_IN), .B0(P1_REIP_REG_25__SCAN_IN), .B1(n14454), .Y(n14473));
  OAI21X1 g11170(.A0(n14453), .A1(n14472), .B0(n14473), .Y(P1_U3220));
  INVX1   g11171(.A(P1_REIP_REG_23__SCAN_IN), .Y(n14475));
  AOI22X1 g11172(.A0(n14443), .A1(P1_ADDRESS_REG_22__SCAN_IN), .B0(P1_REIP_REG_24__SCAN_IN), .B1(n14454), .Y(n14476));
  OAI21X1 g11173(.A0(n14453), .A1(n14475), .B0(n14476), .Y(P1_U3219));
  INVX1   g11174(.A(P1_REIP_REG_22__SCAN_IN), .Y(n14478));
  AOI22X1 g11175(.A0(n14443), .A1(P1_ADDRESS_REG_21__SCAN_IN), .B0(P1_REIP_REG_23__SCAN_IN), .B1(n14454), .Y(n14479));
  OAI21X1 g11176(.A0(n14453), .A1(n14478), .B0(n14479), .Y(P1_U3218));
  INVX1   g11177(.A(P1_REIP_REG_21__SCAN_IN), .Y(n14481));
  AOI22X1 g11178(.A0(n14443), .A1(P1_ADDRESS_REG_20__SCAN_IN), .B0(P1_REIP_REG_22__SCAN_IN), .B1(n14454), .Y(n14482));
  OAI21X1 g11179(.A0(n14453), .A1(n14481), .B0(n14482), .Y(P1_U3217));
  INVX1   g11180(.A(P1_REIP_REG_20__SCAN_IN), .Y(n14484));
  AOI22X1 g11181(.A0(n14443), .A1(P1_ADDRESS_REG_19__SCAN_IN), .B0(P1_REIP_REG_21__SCAN_IN), .B1(n14454), .Y(n14485));
  OAI21X1 g11182(.A0(n14453), .A1(n14484), .B0(n14485), .Y(P1_U3216));
  INVX1   g11183(.A(P1_REIP_REG_19__SCAN_IN), .Y(n14487));
  AOI22X1 g11184(.A0(n14443), .A1(P1_ADDRESS_REG_18__SCAN_IN), .B0(P1_REIP_REG_20__SCAN_IN), .B1(n14454), .Y(n14488));
  OAI21X1 g11185(.A0(n14453), .A1(n14487), .B0(n14488), .Y(P1_U3215));
  INVX1   g11186(.A(P1_REIP_REG_18__SCAN_IN), .Y(n14490));
  AOI22X1 g11187(.A0(n14443), .A1(P1_ADDRESS_REG_17__SCAN_IN), .B0(P1_REIP_REG_19__SCAN_IN), .B1(n14454), .Y(n14491));
  OAI21X1 g11188(.A0(n14453), .A1(n14490), .B0(n14491), .Y(P1_U3214));
  INVX1   g11189(.A(P1_REIP_REG_17__SCAN_IN), .Y(n14493));
  AOI22X1 g11190(.A0(n14443), .A1(P1_ADDRESS_REG_16__SCAN_IN), .B0(P1_REIP_REG_18__SCAN_IN), .B1(n14454), .Y(n14494));
  OAI21X1 g11191(.A0(n14453), .A1(n14493), .B0(n14494), .Y(P1_U3213));
  INVX1   g11192(.A(P1_REIP_REG_16__SCAN_IN), .Y(n14496));
  AOI22X1 g11193(.A0(n14443), .A1(P1_ADDRESS_REG_15__SCAN_IN), .B0(P1_REIP_REG_17__SCAN_IN), .B1(n14454), .Y(n14497));
  OAI21X1 g11194(.A0(n14453), .A1(n14496), .B0(n14497), .Y(P1_U3212));
  INVX1   g11195(.A(P1_REIP_REG_15__SCAN_IN), .Y(n14499));
  AOI22X1 g11196(.A0(n14443), .A1(P1_ADDRESS_REG_14__SCAN_IN), .B0(P1_REIP_REG_16__SCAN_IN), .B1(n14454), .Y(n14500));
  OAI21X1 g11197(.A0(n14453), .A1(n14499), .B0(n14500), .Y(P1_U3211));
  INVX1   g11198(.A(P1_REIP_REG_14__SCAN_IN), .Y(n14502));
  AOI22X1 g11199(.A0(n14443), .A1(P1_ADDRESS_REG_13__SCAN_IN), .B0(P1_REIP_REG_15__SCAN_IN), .B1(n14454), .Y(n14503));
  OAI21X1 g11200(.A0(n14453), .A1(n14502), .B0(n14503), .Y(P1_U3210));
  INVX1   g11201(.A(P1_REIP_REG_13__SCAN_IN), .Y(n14505));
  AOI22X1 g11202(.A0(n14443), .A1(P1_ADDRESS_REG_12__SCAN_IN), .B0(P1_REIP_REG_14__SCAN_IN), .B1(n14454), .Y(n14506));
  OAI21X1 g11203(.A0(n14453), .A1(n14505), .B0(n14506), .Y(P1_U3209));
  INVX1   g11204(.A(P1_REIP_REG_12__SCAN_IN), .Y(n14508));
  AOI22X1 g11205(.A0(n14443), .A1(P1_ADDRESS_REG_11__SCAN_IN), .B0(P1_REIP_REG_13__SCAN_IN), .B1(n14454), .Y(n14509));
  OAI21X1 g11206(.A0(n14453), .A1(n14508), .B0(n14509), .Y(P1_U3208));
  INVX1   g11207(.A(P1_REIP_REG_11__SCAN_IN), .Y(n14511));
  AOI22X1 g11208(.A0(n14443), .A1(P1_ADDRESS_REG_10__SCAN_IN), .B0(P1_REIP_REG_12__SCAN_IN), .B1(n14454), .Y(n14512));
  OAI21X1 g11209(.A0(n14453), .A1(n14511), .B0(n14512), .Y(P1_U3207));
  INVX1   g11210(.A(P1_REIP_REG_10__SCAN_IN), .Y(n14514));
  AOI22X1 g11211(.A0(n14443), .A1(P1_ADDRESS_REG_9__SCAN_IN), .B0(P1_REIP_REG_11__SCAN_IN), .B1(n14454), .Y(n14515));
  OAI21X1 g11212(.A0(n14453), .A1(n14514), .B0(n14515), .Y(P1_U3206));
  INVX1   g11213(.A(P1_REIP_REG_9__SCAN_IN), .Y(n14517));
  AOI22X1 g11214(.A0(n14443), .A1(P1_ADDRESS_REG_8__SCAN_IN), .B0(P1_REIP_REG_10__SCAN_IN), .B1(n14454), .Y(n14518));
  OAI21X1 g11215(.A0(n14453), .A1(n14517), .B0(n14518), .Y(P1_U3205));
  INVX1   g11216(.A(P1_REIP_REG_8__SCAN_IN), .Y(n14520));
  AOI22X1 g11217(.A0(n14443), .A1(P1_ADDRESS_REG_7__SCAN_IN), .B0(P1_REIP_REG_9__SCAN_IN), .B1(n14454), .Y(n14521));
  OAI21X1 g11218(.A0(n14453), .A1(n14520), .B0(n14521), .Y(P1_U3204));
  INVX1   g11219(.A(P1_REIP_REG_7__SCAN_IN), .Y(n14523));
  AOI22X1 g11220(.A0(n14443), .A1(P1_ADDRESS_REG_6__SCAN_IN), .B0(P1_REIP_REG_8__SCAN_IN), .B1(n14454), .Y(n14524));
  OAI21X1 g11221(.A0(n14453), .A1(n14523), .B0(n14524), .Y(P1_U3203));
  INVX1   g11222(.A(P1_REIP_REG_6__SCAN_IN), .Y(n14526));
  AOI22X1 g11223(.A0(n14443), .A1(P1_ADDRESS_REG_5__SCAN_IN), .B0(P1_REIP_REG_7__SCAN_IN), .B1(n14454), .Y(n14527));
  OAI21X1 g11224(.A0(n14453), .A1(n14526), .B0(n14527), .Y(P1_U3202));
  INVX1   g11225(.A(P1_REIP_REG_5__SCAN_IN), .Y(n14529));
  AOI22X1 g11226(.A0(n14443), .A1(P1_ADDRESS_REG_4__SCAN_IN), .B0(P1_REIP_REG_6__SCAN_IN), .B1(n14454), .Y(n14530));
  OAI21X1 g11227(.A0(n14453), .A1(n14529), .B0(n14530), .Y(P1_U3201));
  INVX1   g11228(.A(P1_REIP_REG_4__SCAN_IN), .Y(n14532));
  AOI22X1 g11229(.A0(n14443), .A1(P1_ADDRESS_REG_3__SCAN_IN), .B0(P1_REIP_REG_5__SCAN_IN), .B1(n14454), .Y(n14533));
  OAI21X1 g11230(.A0(n14453), .A1(n14532), .B0(n14533), .Y(P1_U3200));
  NAND4X1 g11231(.A(P1_STATE_REG_1__SCAN_IN), .B(P1_STATE_REG_2__SCAN_IN), .C(P1_REIP_REG_3__SCAN_IN), .D(n14436), .Y(n14535));
  AOI22X1 g11232(.A0(n14443), .A1(P1_ADDRESS_REG_2__SCAN_IN), .B0(P1_REIP_REG_4__SCAN_IN), .B1(n14454), .Y(n14536));
  NAND2X1 g11233(.A(n14536), .B(n14535), .Y(P1_U3199));
  INVX1   g11234(.A(P1_REIP_REG_2__SCAN_IN), .Y(n14538));
  AOI22X1 g11235(.A0(n14443), .A1(P1_ADDRESS_REG_1__SCAN_IN), .B0(P1_REIP_REG_3__SCAN_IN), .B1(n14454), .Y(n14539));
  OAI21X1 g11236(.A0(n14453), .A1(n14538), .B0(n14539), .Y(P1_U3198));
  INVX1   g11237(.A(P1_REIP_REG_1__SCAN_IN), .Y(n14541));
  AOI22X1 g11238(.A0(n14443), .A1(P1_ADDRESS_REG_0__SCAN_IN), .B0(P1_REIP_REG_2__SCAN_IN), .B1(n14454), .Y(n14542));
  OAI21X1 g11239(.A0(n14453), .A1(n14541), .B0(n14542), .Y(P1_U3197));
  INVX1   g11240(.A(P1_STATE_REG_2__SCAN_IN), .Y(n14544));
  INVX1   g11241(.A(READY1), .Y(n14545));
  INVX1   g11242(.A(READY11_REG_SCAN_IN), .Y(n14546));
  NOR2X1  g11243(.A(P1_REQUESTPENDING_REG_SCAN_IN), .B(HOLD), .Y(n14547));
  OAI21X1 g11244(.A0(n14546), .A1(n14545), .B0(n14547), .Y(n14548));
  NOR2X1  g11245(.A(n14546), .B(n14545), .Y(n14549));
  INVX1   g11246(.A(n14549), .Y(n14550));
  INVX1   g11247(.A(P1_REQUESTPENDING_REG_SCAN_IN), .Y(n14551));
  NOR2X1  g11248(.A(n14551), .B(HOLD), .Y(n14552));
  AOI21X1 g11249(.A0(n14552), .A1(n14550), .B0(n14438), .Y(n14553));
  AOI21X1 g11250(.A0(P1_REQUESTPENDING_REG_SCAN_IN), .A1(n3428), .B0(n14436), .Y(n14554));
  OAI21X1 g11251(.A0(P1_REQUESTPENDING_REG_SCAN_IN), .A1(HOLD), .B0(n14554), .Y(n14555));
  OAI21X1 g11252(.A0(P1_STATE_REG_0__SCAN_IN), .A1(NA), .B0(n14555), .Y(n14556));
  AOI21X1 g11253(.A0(n14553), .A1(n14548), .B0(n14556), .Y(n14557));
  NAND3X1 g11254(.A(P1_STATE_REG_1__SCAN_IN), .B(READY11_REG_SCAN_IN), .C(READY1), .Y(n14558));
  NOR2X1  g11255(.A(P1_STATE_REG_1__SCAN_IN), .B(P1_STATE_REG_2__SCAN_IN), .Y(n14559));
  NAND3X1 g11256(.A(n14559), .B(n14551), .C(HOLD), .Y(n14560));
  OAI21X1 g11257(.A0(n14558), .A1(n14547), .B0(n14560), .Y(n14561));
  NOR3X1  g11258(.A(n14438), .B(P1_STATE_REG_2__SCAN_IN), .C(n3419), .Y(n14562));
  NOR2X1  g11259(.A(n14562), .B(n14436), .Y(n14563));
  AOI22X1 g11260(.A0(n14561), .A1(n14563), .B0(n14442), .B1(P1_STATE_REG_2__SCAN_IN), .Y(n14564));
  OAI21X1 g11261(.A0(n14557), .A1(n14544), .B0(n14564), .Y(P1_U3196));
  NAND3X1 g11262(.A(P1_STATE_REG_0__SCAN_IN), .B(n14544), .C(P1_REQUESTPENDING_REG_SCAN_IN), .Y(n14566));
  OAI21X1 g11263(.A0(n14554), .A1(n14544), .B0(n14566), .Y(n14567));
  NAND2X1 g11264(.A(n14567), .B(n14438), .Y(n14568));
  AOI21X1 g11265(.A0(READY11_REG_SCAN_IN), .A1(READY1), .B0(n3428), .Y(n14569));
  OAI21X1 g11266(.A0(n14569), .A1(n14436), .B0(P1_STATE_REG_2__SCAN_IN), .Y(n14570));
  NAND3X1 g11267(.A(n14570), .B(n14548), .C(P1_STATE_REG_1__SCAN_IN), .Y(n14571));
  OAI21X1 g11268(.A0(n14549), .A1(n14544), .B0(n14442), .Y(n14572));
  NAND3X1 g11269(.A(n14572), .B(n14571), .C(n14568), .Y(P1_U3195));
  NAND2X1 g11270(.A(P1_STATE_REG_0__SCAN_IN), .B(P1_REQUESTPENDING_REG_SCAN_IN), .Y(n14574));
  OAI21X1 g11271(.A0(n14574), .A1(n14553), .B0(n14544), .Y(n14575));
  OAI22X1 g11272(.A0(P1_STATE_REG_0__SCAN_IN), .A1(n3419), .B0(n14544), .B1(n14552), .Y(n14576));
  NOR3X1  g11273(.A(n14552), .B(n14436), .C(n14544), .Y(n14577));
  AOI21X1 g11274(.A0(n14576), .A1(n14438), .B0(n14577), .Y(n14578));
  NAND2X1 g11275(.A(n14578), .B(n14575), .Y(P1_U3194));
  OAI21X1 g11276(.A0(P1_STATE_REG_1__SCAN_IN), .A1(P1_STATE_REG_2__SCAN_IN), .B0(n3439), .Y(n14580));
  NOR3X1  g11277(.A(n14436), .B(n14438), .C(P1_STATE_REG_2__SCAN_IN), .Y(n14581));
  AOI21X1 g11278(.A0(n14436), .A1(n14438), .B0(n14581), .Y(n14582));
  NAND2X1 g11279(.A(n14582), .B(P1_DATAWIDTH_REG_0__SCAN_IN), .Y(n14583));
  OAI21X1 g11280(.A0(n14582), .A1(n14580), .B0(n14583), .Y(P1_U3464));
  INVX1   g11281(.A(P1_DATAWIDTH_REG_1__SCAN_IN), .Y(n14585));
  INVX1   g11282(.A(n14582), .Y(n14586));
  NAND2X1 g11283(.A(n14586), .B(n14580), .Y(n14587));
  OAI21X1 g11284(.A0(n14586), .A1(n14585), .B0(n14587), .Y(P1_U3465));
  INVX1   g11285(.A(P1_DATAWIDTH_REG_2__SCAN_IN), .Y(n14589));
  NOR2X1  g11286(.A(n14586), .B(n14589), .Y(P1_U3193));
  INVX1   g11287(.A(P1_DATAWIDTH_REG_3__SCAN_IN), .Y(n14591));
  NOR2X1  g11288(.A(n14586), .B(n14591), .Y(P1_U3192));
  INVX1   g11289(.A(P1_DATAWIDTH_REG_4__SCAN_IN), .Y(n14593));
  NOR2X1  g11290(.A(n14586), .B(n14593), .Y(P1_U3191));
  INVX1   g11291(.A(P1_DATAWIDTH_REG_5__SCAN_IN), .Y(n14595));
  NOR2X1  g11292(.A(n14586), .B(n14595), .Y(P1_U3190));
  INVX1   g11293(.A(P1_DATAWIDTH_REG_6__SCAN_IN), .Y(n14597));
  NOR2X1  g11294(.A(n14586), .B(n14597), .Y(P1_U3189));
  INVX1   g11295(.A(P1_DATAWIDTH_REG_7__SCAN_IN), .Y(n14599));
  NOR2X1  g11296(.A(n14586), .B(n14599), .Y(P1_U3188));
  INVX1   g11297(.A(P1_DATAWIDTH_REG_8__SCAN_IN), .Y(n14601));
  NOR2X1  g11298(.A(n14586), .B(n14601), .Y(P1_U3187));
  INVX1   g11299(.A(P1_DATAWIDTH_REG_9__SCAN_IN), .Y(n14603));
  NOR2X1  g11300(.A(n14586), .B(n14603), .Y(P1_U3186));
  INVX1   g11301(.A(P1_DATAWIDTH_REG_10__SCAN_IN), .Y(n14605));
  NOR2X1  g11302(.A(n14586), .B(n14605), .Y(P1_U3185));
  INVX1   g11303(.A(P1_DATAWIDTH_REG_11__SCAN_IN), .Y(n14607));
  NOR2X1  g11304(.A(n14586), .B(n14607), .Y(P1_U3184));
  INVX1   g11305(.A(P1_DATAWIDTH_REG_12__SCAN_IN), .Y(n14609));
  NOR2X1  g11306(.A(n14586), .B(n14609), .Y(P1_U3183));
  INVX1   g11307(.A(P1_DATAWIDTH_REG_13__SCAN_IN), .Y(n14611));
  NOR2X1  g11308(.A(n14586), .B(n14611), .Y(P1_U3182));
  INVX1   g11309(.A(P1_DATAWIDTH_REG_14__SCAN_IN), .Y(n14613));
  NOR2X1  g11310(.A(n14586), .B(n14613), .Y(P1_U3181));
  INVX1   g11311(.A(P1_DATAWIDTH_REG_15__SCAN_IN), .Y(n14615));
  NOR2X1  g11312(.A(n14586), .B(n14615), .Y(P1_U3180));
  INVX1   g11313(.A(P1_DATAWIDTH_REG_16__SCAN_IN), .Y(n14617));
  NOR2X1  g11314(.A(n14586), .B(n14617), .Y(P1_U3179));
  INVX1   g11315(.A(P1_DATAWIDTH_REG_17__SCAN_IN), .Y(n14619));
  NOR2X1  g11316(.A(n14586), .B(n14619), .Y(P1_U3178));
  INVX1   g11317(.A(P1_DATAWIDTH_REG_18__SCAN_IN), .Y(n14621));
  NOR2X1  g11318(.A(n14586), .B(n14621), .Y(P1_U3177));
  INVX1   g11319(.A(P1_DATAWIDTH_REG_19__SCAN_IN), .Y(n14623));
  NOR2X1  g11320(.A(n14586), .B(n14623), .Y(P1_U3176));
  INVX1   g11321(.A(P1_DATAWIDTH_REG_20__SCAN_IN), .Y(n14625));
  NOR2X1  g11322(.A(n14586), .B(n14625), .Y(P1_U3175));
  INVX1   g11323(.A(P1_DATAWIDTH_REG_21__SCAN_IN), .Y(n14627));
  NOR2X1  g11324(.A(n14586), .B(n14627), .Y(P1_U3174));
  INVX1   g11325(.A(P1_DATAWIDTH_REG_22__SCAN_IN), .Y(n14629));
  NOR2X1  g11326(.A(n14586), .B(n14629), .Y(P1_U3173));
  INVX1   g11327(.A(P1_DATAWIDTH_REG_23__SCAN_IN), .Y(n14631));
  NOR2X1  g11328(.A(n14586), .B(n14631), .Y(P1_U3172));
  INVX1   g11329(.A(P1_DATAWIDTH_REG_24__SCAN_IN), .Y(n14633));
  NOR2X1  g11330(.A(n14586), .B(n14633), .Y(P1_U3171));
  INVX1   g11331(.A(P1_DATAWIDTH_REG_25__SCAN_IN), .Y(n14635));
  NOR2X1  g11332(.A(n14586), .B(n14635), .Y(P1_U3170));
  INVX1   g11333(.A(P1_DATAWIDTH_REG_26__SCAN_IN), .Y(n14637));
  NOR2X1  g11334(.A(n14586), .B(n14637), .Y(P1_U3169));
  INVX1   g11335(.A(P1_DATAWIDTH_REG_27__SCAN_IN), .Y(n14639));
  NOR2X1  g11336(.A(n14586), .B(n14639), .Y(P1_U3168));
  INVX1   g11337(.A(P1_DATAWIDTH_REG_28__SCAN_IN), .Y(n14641));
  NOR2X1  g11338(.A(n14586), .B(n14641), .Y(P1_U3167));
  INVX1   g11339(.A(P1_DATAWIDTH_REG_29__SCAN_IN), .Y(n14643));
  NOR2X1  g11340(.A(n14586), .B(n14643), .Y(P1_U3166));
  INVX1   g11341(.A(P1_DATAWIDTH_REG_30__SCAN_IN), .Y(n14645));
  NOR2X1  g11342(.A(n14586), .B(n14645), .Y(P1_U3165));
  INVX1   g11343(.A(P1_DATAWIDTH_REG_31__SCAN_IN), .Y(n14647));
  NOR2X1  g11344(.A(n14586), .B(n14647), .Y(P1_U3164));
  INVX1   g11345(.A(P1_STATE2_REG_3__SCAN_IN), .Y(n14649));
  INVX1   g11346(.A(P1_STATE2_REG_0__SCAN_IN), .Y(n14650));
  INVX1   g11347(.A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .Y(n14651));
  NOR2X1  g11348(.A(n14651), .B(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .Y(n14652));
  INVX1   g11349(.A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .Y(n14653));
  NOR2X1  g11350(.A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n14653), .Y(n14654));
  INVX1   g11351(.A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Y(n14655));
  INVX1   g11352(.A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .Y(n14656));
  INVX1   g11353(.A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Y(n14657));
  INVX1   g11354(.A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Y(n14658));
  INVX1   g11355(.A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Y(n14659));
  AOI21X1 g11356(.A0(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A1(n14658), .B0(n14659), .Y(n14660));
  NAND3X1 g11357(.A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(n14659), .C(n14658), .Y(n14661));
  AOI21X1 g11358(.A0(n14661), .A1(n14657), .B0(n14660), .Y(n14662));
  AOI21X1 g11359(.A0(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A1(n14656), .B0(n14662), .Y(n14663));
  AOI21X1 g11360(.A0(n14655), .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B0(n14663), .Y(n14664));
  AOI21X1 g11361(.A0(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A1(n14653), .B0(n14664), .Y(n14665));
  INVX1   g11362(.A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .Y(n14666));
  NOR2X1  g11363(.A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n14666), .Y(n14667));
  NOR3X1  g11364(.A(n14667), .B(n14665), .C(n14654), .Y(n14668));
  NOR2X1  g11365(.A(n14668), .B(n14652), .Y(n14669));
  INVX1   g11366(.A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n14670));
  NOR4X1  g11367(.A(n14655), .B(n14657), .C(n14670), .D(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n14671));
  NAND2X1 g11368(.A(n14671), .B(P1_INSTQUEUE_REG_7__0__SCAN_IN), .Y(n14672));
  NOR4X1  g11369(.A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .D(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n14673));
  NOR4X1  g11370(.A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n14657), .C(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .D(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n14674));
  AOI22X1 g11371(.A0(n14673), .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B0(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(n14674), .Y(n14675));
  NAND2X1 g11372(.A(n14675), .B(n14672), .Y(n14676));
  INVX1   g11373(.A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n14677));
  NOR2X1  g11374(.A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n14678));
  NAND4X1 g11375(.A(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B(n14677), .C(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .D(n14678), .Y(n14679));
  NOR4X1  g11376(.A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n14657), .C(n14670), .D(n14677), .Y(n14680));
  NAND2X1 g11377(.A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Y(n14681));
  NOR3X1  g11378(.A(n14681), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n14682));
  AOI22X1 g11379(.A0(n14680), .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B0(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(n14682), .Y(n14683));
  NAND2X1 g11380(.A(n14683), .B(n14679), .Y(n14684));
  NOR2X1  g11381(.A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Y(n14685));
  NAND4X1 g11382(.A(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B(n14657), .C(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .D(n14685), .Y(n14686));
  NOR3X1  g11383(.A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n14687));
  NAND3X1 g11384(.A(n14687), .B(P1_INSTQUEUE_REG_8__0__SCAN_IN), .C(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n14688));
  NAND2X1 g11385(.A(n14688), .B(n14686), .Y(n14689));
  INVX1   g11386(.A(P1_INSTQUEUE_REG_15__0__SCAN_IN), .Y(n14690));
  INVX1   g11387(.A(P1_INSTQUEUE_REG_13__0__SCAN_IN), .Y(n14691));
  NAND4X1 g11388(.A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n14657), .C(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .D(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n14692));
  NAND4X1 g11389(.A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .D(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n14693));
  OAI22X1 g11390(.A0(n14692), .A1(n14691), .B0(n14690), .B1(n14693), .Y(n14694));
  INVX1   g11391(.A(P1_INSTQUEUE_REG_5__0__SCAN_IN), .Y(n14695));
  NAND4X1 g11392(.A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n14657), .C(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .D(n14677), .Y(n14696));
  NAND4X1 g11393(.A(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .D(n14678), .Y(n14697));
  OAI21X1 g11394(.A0(n14696), .A1(n14695), .B0(n14697), .Y(n14698));
  NOR2X1  g11395(.A(n14698), .B(n14694), .Y(n14699));
  NAND4X1 g11396(.A(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .D(n14685), .Y(n14700));
  NOR2X1  g11397(.A(n14677), .B(n14670), .Y(n14701));
  NAND4X1 g11398(.A(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B(n14655), .C(n14657), .D(n14701), .Y(n14702));
  NOR4X1  g11399(.A(n14655), .B(n14657), .C(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .D(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n14703));
  NOR4X1  g11400(.A(n14655), .B(n14657), .C(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .D(n14677), .Y(n14704));
  AOI22X1 g11401(.A0(n14703), .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B0(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(n14704), .Y(n14705));
  NAND4X1 g11402(.A(n14702), .B(n14700), .C(n14699), .D(n14705), .Y(n14706));
  NOR4X1  g11403(.A(n14689), .B(n14684), .C(n14676), .D(n14706), .Y(n14707));
  INVX1   g11404(.A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .Y(n14708));
  INVX1   g11405(.A(n14673), .Y(n14709));
  NOR2X1  g11406(.A(n14709), .B(n14708), .Y(n14710));
  NAND4X1 g11407(.A(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B(n14657), .C(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .D(n14685), .Y(n14711));
  NAND3X1 g11408(.A(n14687), .B(P1_INSTQUEUE_REG_8__4__SCAN_IN), .C(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n14712));
  NOR2X1  g11409(.A(n14655), .B(n14657), .Y(n14713));
  NAND4X1 g11410(.A(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C(n14670), .D(n14713), .Y(n14714));
  NAND4X1 g11411(.A(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .D(n14701), .Y(n14715));
  NAND4X1 g11412(.A(n14714), .B(n14712), .C(n14711), .D(n14715), .Y(n14716));
  INVX1   g11413(.A(P1_INSTQUEUE_REG_7__4__SCAN_IN), .Y(n14717));
  NAND2X1 g11414(.A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n14718));
  NOR4X1  g11415(.A(n14717), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C(n14657), .D(n14718), .Y(n14719));
  NAND2X1 g11416(.A(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Y(n14720));
  NOR4X1  g11417(.A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .D(n14720), .Y(n14721));
  NAND3X1 g11418(.A(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n14722));
  NOR3X1  g11419(.A(n14722), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Y(n14723));
  NOR3X1  g11420(.A(n14723), .B(n14721), .C(n14719), .Y(n14724));
  NAND2X1 g11421(.A(n14677), .B(n14670), .Y(n14725));
  NAND3X1 g11422(.A(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Y(n14726));
  NAND3X1 g11423(.A(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C(n14657), .Y(n14727));
  OAI22X1 g11424(.A0(n14726), .A1(n14725), .B0(n14718), .B1(n14727), .Y(n14728));
  INVX1   g11425(.A(n14678), .Y(n14729));
  NAND3X1 g11426(.A(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B(n14677), .C(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Y(n14730));
  NAND3X1 g11427(.A(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Y(n14731));
  AOI21X1 g11428(.A0(n14731), .A1(n14730), .B0(n14729), .Y(n14732));
  NOR2X1  g11429(.A(n14732), .B(n14728), .Y(n14733));
  INVX1   g11430(.A(n14685), .Y(n14734));
  INVX1   g11431(.A(n14701), .Y(n14735));
  NAND3X1 g11432(.A(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B(n14655), .C(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Y(n14736));
  NAND3X1 g11433(.A(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n14737));
  OAI22X1 g11434(.A0(n14736), .A1(n14735), .B0(n14734), .B1(n14737), .Y(n14738));
  NAND2X1 g11435(.A(n14655), .B(n14657), .Y(n14739));
  NOR2X1  g11436(.A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n14740));
  NAND4X1 g11437(.A(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .D(n14740), .Y(n14741));
  NAND3X1 g11438(.A(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n14742));
  OAI21X1 g11439(.A0(n14742), .A1(n14739), .B0(n14741), .Y(n14743));
  NOR2X1  g11440(.A(n14743), .B(n14738), .Y(n14744));
  NAND3X1 g11441(.A(n14744), .B(n14733), .C(n14724), .Y(n14745));
  NOR3X1  g11442(.A(n14745), .B(n14716), .C(n14710), .Y(n14746));
  NOR4X1  g11443(.A(n14707), .B(n14669), .C(n14650), .D(n14746), .Y(n14747));
  INVX1   g11444(.A(n14669), .Y(n14748));
  NAND2X1 g11445(.A(n14671), .B(P1_INSTQUEUE_REG_7__1__SCAN_IN), .Y(n14749));
  AOI22X1 g11446(.A0(n14673), .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B0(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(n14674), .Y(n14750));
  NAND2X1 g11447(.A(n14750), .B(n14749), .Y(n14751));
  NAND4X1 g11448(.A(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B(n14677), .C(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .D(n14678), .Y(n14752));
  AOI22X1 g11449(.A0(n14680), .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B0(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(n14682), .Y(n14753));
  NAND2X1 g11450(.A(n14753), .B(n14752), .Y(n14754));
  NAND4X1 g11451(.A(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B(n14657), .C(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .D(n14685), .Y(n14755));
  NAND3X1 g11452(.A(n14687), .B(P1_INSTQUEUE_REG_8__1__SCAN_IN), .C(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n14756));
  NAND2X1 g11453(.A(n14756), .B(n14755), .Y(n14757));
  INVX1   g11454(.A(P1_INSTQUEUE_REG_15__1__SCAN_IN), .Y(n14758));
  INVX1   g11455(.A(P1_INSTQUEUE_REG_13__1__SCAN_IN), .Y(n14759));
  OAI22X1 g11456(.A0(n14692), .A1(n14759), .B0(n14758), .B1(n14693), .Y(n14760));
  INVX1   g11457(.A(P1_INSTQUEUE_REG_5__1__SCAN_IN), .Y(n14761));
  NAND4X1 g11458(.A(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .D(n14678), .Y(n14762));
  OAI21X1 g11459(.A0(n14696), .A1(n14761), .B0(n14762), .Y(n14763));
  NOR2X1  g11460(.A(n14763), .B(n14760), .Y(n14764));
  NAND4X1 g11461(.A(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .D(n14685), .Y(n14765));
  NAND4X1 g11462(.A(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B(n14655), .C(n14657), .D(n14701), .Y(n14766));
  AOI22X1 g11463(.A0(n14703), .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B0(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(n14704), .Y(n14767));
  NAND4X1 g11464(.A(n14766), .B(n14765), .C(n14764), .D(n14767), .Y(n14768));
  NOR4X1  g11465(.A(n14757), .B(n14754), .C(n14751), .D(n14768), .Y(n14769));
  INVX1   g11466(.A(n14769), .Y(n14770));
  NAND4X1 g11467(.A(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .D(n14678), .Y(n14771));
  NAND4X1 g11468(.A(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .D(n14701), .Y(n14772));
  NAND2X1 g11469(.A(n14772), .B(n14771), .Y(n14773));
  NAND4X1 g11470(.A(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B(n14655), .C(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .D(n14701), .Y(n14774));
  NAND4X1 g11471(.A(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(n14657), .D(n14701), .Y(n14775));
  NAND2X1 g11472(.A(n14775), .B(n14774), .Y(n14776));
  NAND4X1 g11473(.A(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .D(n14740), .Y(n14777));
  NAND4X1 g11474(.A(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .D(n14685), .Y(n14778));
  NAND2X1 g11475(.A(n14778), .B(n14777), .Y(n14779));
  NAND3X1 g11476(.A(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(n14670), .Y(n14780));
  NAND3X1 g11477(.A(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n14781));
  OAI22X1 g11478(.A0(n14780), .A1(n14681), .B0(n14739), .B1(n14781), .Y(n14782));
  NOR4X1  g11479(.A(n14779), .B(n14776), .C(n14773), .D(n14782), .Y(n14783));
  INVX1   g11480(.A(P1_INSTQUEUE_REG_2__5__SCAN_IN), .Y(n14784));
  NOR4X1  g11481(.A(n14784), .B(n14657), .C(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .D(n14734), .Y(n14785));
  INVX1   g11482(.A(P1_INSTQUEUE_REG_1__5__SCAN_IN), .Y(n14786));
  NOR4X1  g11483(.A(n14786), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C(n14670), .D(n14734), .Y(n14787));
  INVX1   g11484(.A(P1_INSTQUEUE_REG_4__5__SCAN_IN), .Y(n14788));
  NOR4X1  g11485(.A(n14788), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C(n14655), .D(n14729), .Y(n14789));
  NOR3X1  g11486(.A(n14789), .B(n14787), .C(n14785), .Y(n14790));
  NAND2X1 g11487(.A(n14673), .B(P1_INSTQUEUE_REG_0__5__SCAN_IN), .Y(n14791));
  INVX1   g11488(.A(P1_INSTQUEUE_REG_7__5__SCAN_IN), .Y(n14792));
  NOR4X1  g11489(.A(n14792), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C(n14657), .D(n14718), .Y(n14793));
  INVX1   g11490(.A(P1_INSTQUEUE_REG_6__5__SCAN_IN), .Y(n14794));
  NOR4X1  g11491(.A(n14794), .B(n14655), .C(n14657), .D(n14725), .Y(n14795));
  INVX1   g11492(.A(P1_INSTQUEUE_REG_5__5__SCAN_IN), .Y(n14796));
  NOR4X1  g11493(.A(n14796), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .D(n14718), .Y(n14797));
  NAND2X1 g11494(.A(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n14798));
  NOR4X1  g11495(.A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .D(n14798), .Y(n14799));
  NOR4X1  g11496(.A(n14797), .B(n14795), .C(n14793), .D(n14799), .Y(n14800));
  NAND4X1 g11497(.A(n14791), .B(n14790), .C(n14783), .D(n14800), .Y(n14801));
  NOR3X1  g11498(.A(n14801), .B(n14770), .C(n14650), .Y(n14802));
  NAND2X1 g11499(.A(n14801), .B(n14746), .Y(n14803));
  NOR2X1  g11500(.A(n14803), .B(n14650), .Y(n14804));
  INVX1   g11501(.A(n14804), .Y(n14805));
  INVX1   g11502(.A(n14707), .Y(n14806));
  NAND2X1 g11503(.A(n14770), .B(n14806), .Y(n14807));
  INVX1   g11504(.A(n14801), .Y(n14808));
  NOR4X1  g11505(.A(n14770), .B(n14707), .C(n14650), .D(n14808), .Y(n14809));
  NOR3X1  g11506(.A(n14769), .B(n14806), .C(n14650), .Y(n14810));
  NOR3X1  g11507(.A(n14801), .B(n14769), .C(n14650), .Y(n14811));
  NOR3X1  g11508(.A(n14770), .B(n14806), .C(n14650), .Y(n14812));
  NOR4X1  g11509(.A(n14811), .B(n14810), .C(n14809), .D(n14812), .Y(n14813));
  OAI21X1 g11510(.A0(n14807), .A1(n14805), .B0(n14813), .Y(n14814));
  OAI21X1 g11511(.A0(n14814), .A1(n14802), .B0(n14748), .Y(n14815));
  INVX1   g11512(.A(n14747), .Y(n14816));
  INVX1   g11513(.A(n14815), .Y(n14817));
  NOR3X1  g11514(.A(n14746), .B(n14707), .C(n14650), .Y(n14818));
  INVX1   g11515(.A(n14818), .Y(n14819));
  NOR2X1  g11516(.A(n14808), .B(n14769), .Y(n14820));
  INVX1   g11517(.A(n14820), .Y(n14821));
  NOR2X1  g11518(.A(n14821), .B(n14819), .Y(n14822));
  NOR2X1  g11519(.A(n14808), .B(n14650), .Y(n14823));
  NOR2X1  g11520(.A(n14806), .B(n14650), .Y(n14824));
  OAI21X1 g11521(.A0(n14824), .A1(n14823), .B0(n14769), .Y(n14825));
  INVX1   g11522(.A(n14825), .Y(n14826));
  XOR2X1  g11523(.A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B(n14658), .Y(n14827));
  AOI22X1 g11524(.A0(n14806), .A1(n14804), .B0(n14650), .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n14828));
  OAI21X1 g11525(.A0(n14827), .A1(n14819), .B0(n14828), .Y(n14829));
  NOR2X1  g11526(.A(n14829), .B(n14826), .Y(n14830));
  INVX1   g11527(.A(n14830), .Y(n14831));
  INVX1   g11528(.A(n14814), .Y(n14832));
  NOR2X1  g11529(.A(n14746), .B(n14707), .Y(n14833));
  NOR4X1  g11530(.A(n14801), .B(n14770), .C(n14650), .D(n14827), .Y(n14834));
  NOR3X1  g11531(.A(n14834), .B(n14833), .C(n14650), .Y(n14835));
  OAI21X1 g11532(.A0(n14827), .A1(n14832), .B0(n14835), .Y(n14836));
  INVX1   g11533(.A(n14836), .Y(n14837));
  OAI21X1 g11534(.A0(n14837), .A1(n14831), .B0(n14822), .Y(n14838));
  NOR2X1  g11535(.A(n14670), .B(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Y(n14839));
  XOR2X1  g11536(.A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n14659), .Y(n14840));
  XOR2X1  g11537(.A(n14840), .B(n14839), .Y(n14841));
  INVX1   g11538(.A(n14841), .Y(n14842));
  AOI21X1 g11539(.A0(n14842), .A1(n14802), .B0(n14650), .Y(n14843));
  OAI21X1 g11540(.A0(n14841), .A1(n14832), .B0(n14843), .Y(n14844));
  NOR4X1  g11541(.A(n14746), .B(n14707), .C(n14650), .D(n14841), .Y(n14845));
  INVX1   g11542(.A(n14746), .Y(n14846));
  NOR3X1  g11543(.A(n14769), .B(n14846), .C(n14650), .Y(n14847));
  NOR2X1  g11544(.A(n14801), .B(n14650), .Y(n14848));
  AOI21X1 g11545(.A0(n14650), .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B0(n14848), .Y(n14849));
  INVX1   g11546(.A(n14849), .Y(n14850));
  NOR4X1  g11547(.A(n14847), .B(n14845), .C(n14810), .D(n14850), .Y(n14851));
  NOR2X1  g11548(.A(n14851), .B(n14844), .Y(n14852));
  AOI21X1 g11549(.A0(n14837), .A1(n14831), .B0(n14852), .Y(n14853));
  XOR2X1  g11550(.A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n14656), .Y(n14854));
  XOR2X1  g11551(.A(n14854), .B(n14662), .Y(n14855));
  INVX1   g11552(.A(n14855), .Y(n14856));
  AOI22X1 g11553(.A0(n14818), .A1(n14856), .B0(n14650), .B1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Y(n14857));
  NAND2X1 g11554(.A(n14857), .B(n14825), .Y(n14858));
  INVX1   g11555(.A(n14858), .Y(n14859));
  NOR4X1  g11556(.A(n14801), .B(n14770), .C(n14650), .D(n14855), .Y(n14860));
  NOR3X1  g11557(.A(n14860), .B(n14833), .C(n14650), .Y(n14861));
  OAI21X1 g11558(.A0(n14855), .A1(n14832), .B0(n14861), .Y(n14862));
  AOI22X1 g11559(.A0(n14859), .A1(n14862), .B0(n14851), .B1(n14844), .Y(n14863));
  INVX1   g11560(.A(n14863), .Y(n14864));
  AOI21X1 g11561(.A0(n14853), .A1(n14838), .B0(n14864), .Y(n14865));
  XOR2X1  g11562(.A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n14653), .Y(n14866));
  XOR2X1  g11563(.A(n14866), .B(n14664), .Y(n14867));
  INVX1   g11564(.A(n14867), .Y(n14868));
  AOI21X1 g11565(.A0(n14868), .A1(n14802), .B0(n14650), .Y(n14869));
  OAI21X1 g11566(.A0(n14867), .A1(n14832), .B0(n14869), .Y(n14870));
  AOI22X1 g11567(.A0(n14818), .A1(n14868), .B0(n14650), .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n14871));
  OAI22X1 g11568(.A0(n14870), .A1(n14871), .B0(n14862), .B1(n14859), .Y(n14872));
  NOR2X1  g11569(.A(n14665), .B(n14654), .Y(n14873));
  XOR2X1  g11570(.A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n14666), .Y(n14874));
  XOR2X1  g11571(.A(n14874), .B(n14873), .Y(n14875));
  INVX1   g11572(.A(n14875), .Y(n14876));
  AOI22X1 g11573(.A0(n14818), .A1(n14876), .B0(n14650), .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .Y(n14877));
  OAI21X1 g11574(.A0(n14814), .A1(n14802), .B0(n14876), .Y(n14878));
  INVX1   g11575(.A(n14878), .Y(n14879));
  AOI22X1 g11576(.A0(n14877), .A1(n14879), .B0(n14871), .B1(n14870), .Y(n14880));
  OAI21X1 g11577(.A0(n14872), .A1(n14865), .B0(n14880), .Y(n14881));
  OAI22X1 g11578(.A0(n14877), .A1(n14879), .B0(n14817), .B1(n14816), .Y(n14882));
  INVX1   g11579(.A(n14882), .Y(n14883));
  AOI22X1 g11580(.A0(n14881), .A1(n14883), .B0(n14817), .B1(n14816), .Y(n14884));
  NAND2X1 g11581(.A(n14815), .B(P1_STATE2_REG_0__SCAN_IN), .Y(n14885));
  OAI21X1 g11582(.A0(n14884), .A1(n14815), .B0(n14885), .Y(n14886));
  NAND2X1 g11583(.A(n14886), .B(n14747), .Y(n14887));
  NOR2X1  g11584(.A(n14884), .B(n14817), .Y(n14888));
  NOR2X1  g11585(.A(n14815), .B(P1_STATE2_REG_0__SCAN_IN), .Y(n14889));
  OAI21X1 g11586(.A0(n14889), .A1(n14888), .B0(n14816), .Y(n14890));
  INVX1   g11587(.A(P1_INSTQUEUE_REG_0__6__SCAN_IN), .Y(n14891));
  NOR2X1  g11588(.A(n14709), .B(n14891), .Y(n14892));
  NAND4X1 g11589(.A(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .D(n14685), .Y(n14893));
  NAND4X1 g11590(.A(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B(n14655), .C(n14657), .D(n14701), .Y(n14894));
  NOR2X1  g11591(.A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n14655), .Y(n14895));
  NOR2X1  g11592(.A(n14657), .B(n14670), .Y(n14896));
  NAND3X1 g11593(.A(n14896), .B(n14895), .C(P1_INSTQUEUE_REG_7__6__SCAN_IN), .Y(n14897));
  NAND3X1 g11594(.A(n14687), .B(P1_INSTQUEUE_REG_8__6__SCAN_IN), .C(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n14898));
  NAND4X1 g11595(.A(n14897), .B(n14894), .C(n14893), .D(n14898), .Y(n14899));
  NAND4X1 g11596(.A(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B(n14657), .C(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .D(n14685), .Y(n14900));
  NAND4X1 g11597(.A(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B(n14677), .C(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .D(n14678), .Y(n14901));
  NAND4X1 g11598(.A(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C(n14670), .D(n14685), .Y(n14902));
  NAND3X1 g11599(.A(n14902), .B(n14901), .C(n14900), .Y(n14903));
  NAND4X1 g11600(.A(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B(n14657), .C(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .D(n14895), .Y(n14904));
  NAND4X1 g11601(.A(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .D(n14896), .Y(n14905));
  NAND2X1 g11602(.A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Y(n14906));
  NOR3X1  g11603(.A(n14906), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n14907));
  INVX1   g11604(.A(P1_INSTQUEUE_REG_6__6__SCAN_IN), .Y(n14908));
  NOR3X1  g11605(.A(n14908), .B(n14657), .C(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n14909));
  AOI22X1 g11606(.A0(n14907), .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B0(n14895), .B1(n14909), .Y(n14910));
  NAND4X1 g11607(.A(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .D(n14740), .Y(n14911));
  NAND3X1 g11608(.A(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B(n14655), .C(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Y(n14912));
  OAI21X1 g11609(.A0(n14912), .A1(n14735), .B0(n14911), .Y(n14913));
  NAND3X1 g11610(.A(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C(n14670), .Y(n14914));
  NAND3X1 g11611(.A(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B(n14657), .C(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n14915));
  AOI21X1 g11612(.A0(n14915), .A1(n14914), .B0(n14906), .Y(n14916));
  NOR2X1  g11613(.A(n14916), .B(n14913), .Y(n14917));
  NAND4X1 g11614(.A(n14910), .B(n14905), .C(n14904), .D(n14917), .Y(n14918));
  NOR4X1  g11615(.A(n14903), .B(n14899), .C(n14892), .D(n14918), .Y(n14919));
  NAND2X1 g11616(.A(n14671), .B(P1_INSTQUEUE_REG_7__3__SCAN_IN), .Y(n14920));
  AOI22X1 g11617(.A0(n14673), .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B0(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(n14674), .Y(n14921));
  NAND2X1 g11618(.A(n14921), .B(n14920), .Y(n14922));
  NAND4X1 g11619(.A(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B(n14677), .C(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .D(n14678), .Y(n14923));
  AOI22X1 g11620(.A0(n14680), .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B0(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(n14682), .Y(n14924));
  NAND2X1 g11621(.A(n14924), .B(n14923), .Y(n14925));
  NAND4X1 g11622(.A(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B(n14657), .C(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .D(n14685), .Y(n14926));
  NAND3X1 g11623(.A(n14687), .B(P1_INSTQUEUE_REG_8__3__SCAN_IN), .C(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n14927));
  NAND2X1 g11624(.A(n14927), .B(n14926), .Y(n14928));
  INVX1   g11625(.A(P1_INSTQUEUE_REG_15__3__SCAN_IN), .Y(n14929));
  INVX1   g11626(.A(P1_INSTQUEUE_REG_13__3__SCAN_IN), .Y(n14930));
  OAI22X1 g11627(.A0(n14692), .A1(n14930), .B0(n14929), .B1(n14693), .Y(n14931));
  INVX1   g11628(.A(P1_INSTQUEUE_REG_5__3__SCAN_IN), .Y(n14932));
  NAND4X1 g11629(.A(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .D(n14678), .Y(n14933));
  OAI21X1 g11630(.A0(n14696), .A1(n14932), .B0(n14933), .Y(n14934));
  NOR2X1  g11631(.A(n14934), .B(n14931), .Y(n14935));
  NAND4X1 g11632(.A(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .D(n14685), .Y(n14936));
  NAND4X1 g11633(.A(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B(n14655), .C(n14657), .D(n14701), .Y(n14937));
  AOI22X1 g11634(.A0(n14703), .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B0(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(n14704), .Y(n14938));
  NAND4X1 g11635(.A(n14937), .B(n14936), .C(n14935), .D(n14938), .Y(n14939));
  NOR4X1  g11636(.A(n14928), .B(n14925), .C(n14922), .D(n14939), .Y(n14940));
  NAND2X1 g11637(.A(n14671), .B(P1_INSTQUEUE_REG_7__7__SCAN_IN), .Y(n14941));
  AOI22X1 g11638(.A0(n14673), .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B0(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(n14674), .Y(n14942));
  NAND2X1 g11639(.A(n14942), .B(n14941), .Y(n14943));
  NAND4X1 g11640(.A(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B(n14677), .C(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .D(n14678), .Y(n14944));
  AOI22X1 g11641(.A0(n14680), .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B0(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(n14682), .Y(n14945));
  NAND2X1 g11642(.A(n14945), .B(n14944), .Y(n14946));
  INVX1   g11643(.A(P1_INSTQUEUE_REG_1__7__SCAN_IN), .Y(n14947));
  NAND3X1 g11644(.A(n14685), .B(n14657), .C(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n14948));
  NAND3X1 g11645(.A(n14687), .B(P1_INSTQUEUE_REG_8__7__SCAN_IN), .C(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n14949));
  OAI21X1 g11646(.A0(n14948), .A1(n14947), .B0(n14949), .Y(n14950));
  INVX1   g11647(.A(P1_INSTQUEUE_REG_15__7__SCAN_IN), .Y(n14951));
  INVX1   g11648(.A(P1_INSTQUEUE_REG_13__7__SCAN_IN), .Y(n14952));
  OAI22X1 g11649(.A0(n14692), .A1(n14952), .B0(n14951), .B1(n14693), .Y(n14953));
  INVX1   g11650(.A(P1_INSTQUEUE_REG_5__7__SCAN_IN), .Y(n14954));
  NAND4X1 g11651(.A(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .D(n14678), .Y(n14955));
  OAI21X1 g11652(.A0(n14696), .A1(n14954), .B0(n14955), .Y(n14956));
  NOR2X1  g11653(.A(n14956), .B(n14953), .Y(n14957));
  NAND4X1 g11654(.A(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .D(n14685), .Y(n14958));
  NAND4X1 g11655(.A(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B(n14655), .C(n14657), .D(n14701), .Y(n14959));
  AOI22X1 g11656(.A0(n14703), .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B0(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(n14704), .Y(n14960));
  NAND4X1 g11657(.A(n14959), .B(n14958), .C(n14957), .D(n14960), .Y(n14961));
  NOR4X1  g11658(.A(n14950), .B(n14946), .C(n14943), .D(n14961), .Y(n14962));
  NOR2X1  g11659(.A(n14962), .B(n14940), .Y(n14963));
  NAND2X1 g11660(.A(n14671), .B(P1_INSTQUEUE_REG_7__2__SCAN_IN), .Y(n14964));
  AOI22X1 g11661(.A0(n14673), .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B0(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(n14674), .Y(n14965));
  NAND2X1 g11662(.A(n14965), .B(n14964), .Y(n14966));
  NAND4X1 g11663(.A(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B(n14677), .C(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .D(n14678), .Y(n14967));
  AOI22X1 g11664(.A0(n14680), .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B0(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(n14682), .Y(n14968));
  NAND2X1 g11665(.A(n14968), .B(n14967), .Y(n14969));
  NAND4X1 g11666(.A(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B(n14657), .C(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .D(n14685), .Y(n14970));
  NAND3X1 g11667(.A(n14687), .B(P1_INSTQUEUE_REG_8__2__SCAN_IN), .C(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n14971));
  NAND2X1 g11668(.A(n14971), .B(n14970), .Y(n14972));
  INVX1   g11669(.A(P1_INSTQUEUE_REG_15__2__SCAN_IN), .Y(n14973));
  INVX1   g11670(.A(P1_INSTQUEUE_REG_13__2__SCAN_IN), .Y(n14974));
  OAI22X1 g11671(.A0(n14692), .A1(n14974), .B0(n14973), .B1(n14693), .Y(n14975));
  INVX1   g11672(.A(P1_INSTQUEUE_REG_5__2__SCAN_IN), .Y(n14976));
  NAND4X1 g11673(.A(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .D(n14678), .Y(n14977));
  OAI21X1 g11674(.A0(n14696), .A1(n14976), .B0(n14977), .Y(n14978));
  NOR2X1  g11675(.A(n14978), .B(n14975), .Y(n14979));
  NAND4X1 g11676(.A(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .D(n14685), .Y(n14980));
  NAND4X1 g11677(.A(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B(n14655), .C(n14657), .D(n14701), .Y(n14981));
  AOI22X1 g11678(.A0(n14703), .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B0(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(n14704), .Y(n14982));
  NAND4X1 g11679(.A(n14981), .B(n14980), .C(n14979), .D(n14982), .Y(n14983));
  NOR4X1  g11680(.A(n14972), .B(n14969), .C(n14966), .D(n14983), .Y(n14984));
  INVX1   g11681(.A(n14984), .Y(n14985));
  NOR4X1  g11682(.A(n14745), .B(n14716), .C(n14710), .D(n14985), .Y(n14986));
  NAND4X1 g11683(.A(n14963), .B(n14919), .C(n14808), .D(n14986), .Y(n14987));
  INVX1   g11684(.A(n14987), .Y(n14988));
  NOR2X1  g11685(.A(n14769), .B(n14806), .Y(n14989));
  INVX1   g11686(.A(n14989), .Y(n14990));
  NAND2X1 g11687(.A(n14985), .B(n14940), .Y(n14991));
  NOR2X1  g11688(.A(n14962), .B(n14919), .Y(n14992));
  INVX1   g11689(.A(n14992), .Y(n14993));
  NOR4X1  g11690(.A(n14991), .B(n14990), .C(n14803), .D(n14993), .Y(n14994));
  XOR2X1  g11691(.A(P1_STATE_REG_1__SCAN_IN), .B(n14544), .Y(n14995));
  NOR3X1  g11692(.A(n14995), .B(n14549), .C(P1_STATE_REG_0__SCAN_IN), .Y(n14996));
  OAI21X1 g11693(.A0(n14994), .A1(n14988), .B0(n14996), .Y(n14997));
  INVX1   g11694(.A(n14919), .Y(n14998));
  NOR4X1  g11695(.A(n14998), .B(n14808), .C(n14746), .D(n14962), .Y(n14999));
  INVX1   g11696(.A(n14999), .Y(n15000));
  NOR2X1  g11697(.A(n14770), .B(n14806), .Y(n15001));
  INVX1   g11698(.A(n15001), .Y(n15002));
  NOR4X1  g11699(.A(n15000), .B(n14985), .C(n14940), .D(n15002), .Y(n15003));
  NOR3X1  g11700(.A(n14987), .B(n14807), .C(n14549), .Y(n15004));
  NOR2X1  g11701(.A(n15004), .B(n15003), .Y(n15005));
  AOI22X1 g11702(.A0(n14997), .A1(n15005), .B0(n14890), .B1(n14887), .Y(n15006));
  NAND2X1 g11703(.A(n14890), .B(n14887), .Y(n15007));
  NOR3X1  g11704(.A(n14940), .B(n14769), .C(n14707), .Y(n15008));
  INVX1   g11705(.A(n15008), .Y(n15009));
  NOR3X1  g11706(.A(n15009), .B(n15000), .C(n14985), .Y(n15010));
  INVX1   g11707(.A(n15010), .Y(n15011));
  NOR2X1  g11708(.A(n15011), .B(n15007), .Y(n15012));
  NOR2X1  g11709(.A(n14999), .B(n14806), .Y(n15013));
  NOR2X1  g11710(.A(n14919), .B(n14801), .Y(n15014));
  NOR2X1  g11711(.A(n15014), .B(n14962), .Y(n15015));
  NAND3X1 g11712(.A(n14919), .B(n14801), .C(n14746), .Y(n15016));
  NAND2X1 g11713(.A(n15016), .B(n15015), .Y(n15017));
  NOR3X1  g11714(.A(n15017), .B(n15013), .C(n14940), .Y(n15018));
  NOR2X1  g11715(.A(n15018), .B(n14985), .Y(n15019));
  NOR2X1  g11716(.A(n14770), .B(n14707), .Y(n15020));
  INVX1   g11717(.A(n15020), .Y(n15021));
  NOR2X1  g11718(.A(n14998), .B(n14808), .Y(n15022));
  NOR3X1  g11719(.A(n15022), .B(n15014), .C(n14962), .Y(n15023));
  INVX1   g11720(.A(n14940), .Y(n15024));
  NOR4X1  g11721(.A(n15024), .B(n14803), .C(n14806), .D(n14993), .Y(n15025));
  OAI22X1 g11722(.A0(n15023), .A1(n15021), .B0(n14984), .B1(n15025), .Y(n15026));
  NOR4X1  g11723(.A(n14993), .B(n14991), .C(n14803), .D(n15002), .Y(n15027));
  INVX1   g11724(.A(n15027), .Y(n15028));
  NOR3X1  g11725(.A(n14868), .B(n14856), .C(n14842), .Y(n15029));
  AOI21X1 g11726(.A0(n15029), .A1(n14875), .B0(n14748), .Y(n15030));
  NAND2X1 g11727(.A(n15030), .B(n14550), .Y(n15031));
  INVX1   g11728(.A(n15022), .Y(n15032));
  AOI22X1 g11729(.A0(n14989), .A1(n14984), .B0(n14833), .B1(n15032), .Y(n15033));
  OAI21X1 g11730(.A0(n15031), .A1(n15028), .B0(n15033), .Y(n15034));
  NOR3X1  g11731(.A(n15034), .B(n15026), .C(n15019), .Y(n15035));
  INVX1   g11732(.A(n15035), .Y(n15036));
  NOR3X1  g11733(.A(n15036), .B(n15012), .C(n15006), .Y(n15037));
  INVX1   g11734(.A(n15037), .Y(n15038));
  NOR4X1  g11735(.A(n14745), .B(n14716), .C(n14710), .D(n14808), .Y(n15039));
  OAI21X1 g11736(.A0(n14998), .A1(n14746), .B0(n14984), .Y(n15040));
  NOR2X1  g11737(.A(n14999), .B(n14940), .Y(n15041));
  INVX1   g11738(.A(n14962), .Y(n15042));
  AOI21X1 g11739(.A0(n14808), .A1(n14746), .B0(n15042), .Y(n15043));
  NOR2X1  g11740(.A(n15043), .B(n15041), .Y(n15044));
  OAI21X1 g11741(.A0(n15040), .A1(n15014), .B0(n15044), .Y(n15045));
  INVX1   g11742(.A(n15014), .Y(n15046));
  AOI21X1 g11743(.A0(n15042), .A1(n14919), .B0(n14846), .Y(n15047));
  AOI21X1 g11744(.A0(n15047), .A1(n15046), .B0(n14984), .Y(n15048));
  OAI21X1 g11745(.A0(n15048), .A1(n15045), .B0(n14769), .Y(n15049));
  OAI21X1 g11746(.A0(n15039), .A1(n14769), .B0(n15049), .Y(n15050));
  NOR3X1  g11747(.A(n14985), .B(n15024), .C(n14806), .Y(n15051));
  NOR2X1  g11748(.A(n14984), .B(n14998), .Y(n15052));
  OAI21X1 g11749(.A0(n15052), .A1(n15051), .B0(n14770), .Y(n15053));
  NOR2X1  g11750(.A(n14940), .B(n14769), .Y(n15054));
  OAI21X1 g11751(.A0(n15054), .A1(n14806), .B0(n14985), .Y(n15055));
  NOR2X1  g11752(.A(n15024), .B(n14707), .Y(n15056));
  AOI21X1 g11753(.A0(n15032), .A1(n14833), .B0(n15056), .Y(n15057));
  OAI21X1 g11754(.A0(n14998), .A1(n14808), .B0(n15015), .Y(n15058));
  AOI22X1 g11755(.A0(n15017), .A1(n15054), .B0(n15020), .B1(n15058), .Y(n15059));
  NAND4X1 g11756(.A(n15057), .B(n15055), .C(n15053), .D(n15059), .Y(n15060));
  AOI21X1 g11757(.A0(n15050), .A1(n14707), .B0(n15060), .Y(n15061));
  NAND3X1 g11758(.A(n15054), .B(n14992), .C(n15039), .Y(n15062));
  INVX1   g11759(.A(n15062), .Y(n15063));
  NOR2X1  g11760(.A(n14985), .B(n15024), .Y(n15064));
  INVX1   g11761(.A(n15064), .Y(n15065));
  NOR3X1  g11762(.A(n15065), .B(n15002), .C(n14801), .Y(n15066));
  NOR3X1  g11763(.A(n15066), .B(n15063), .C(n14988), .Y(n15067));
  NOR2X1  g11764(.A(n14998), .B(n14801), .Y(n15068));
  INVX1   g11765(.A(n15068), .Y(n15069));
  NAND2X1 g11766(.A(n14962), .B(n14746), .Y(n15070));
  NOR4X1  g11767(.A(n14984), .B(n15024), .C(n15069), .D(n15070), .Y(n15071));
  NOR3X1  g11768(.A(n15070), .B(n14919), .C(n14801), .Y(n15072));
  AOI22X1 g11769(.A0(n15051), .A1(n15072), .B0(n14962), .B1(n14770), .Y(n15073));
  INVX1   g11770(.A(n15073), .Y(n15074));
  NOR3X1  g11771(.A(n15074), .B(n15071), .C(n15027), .Y(n15075));
  NAND3X1 g11772(.A(n15075), .B(n15067), .C(n15061), .Y(n15076));
  INVX1   g11773(.A(n15076), .Y(n15077));
  NAND2X1 g11774(.A(n15050), .B(n14707), .Y(n15078));
  OAI21X1 g11775(.A0(n14998), .A1(n14808), .B0(n14846), .Y(n15079));
  NAND3X1 g11776(.A(n15079), .B(n15016), .C(n15015), .Y(n15080));
  OAI21X1 g11777(.A0(n14985), .A1(n15024), .B0(n14806), .Y(n15081));
  OAI21X1 g11778(.A0(n15081), .A1(n15080), .B0(n14770), .Y(n15082));
  NOR3X1  g11779(.A(n14650), .B(P1_STATE2_REG_1__SCAN_IN), .C(P1_STATE2_REG_3__SCAN_IN), .Y(n15083));
  OAI21X1 g11780(.A0(n14984), .A1(n14707), .B0(n15083), .Y(n15084));
  INVX1   g11781(.A(n15051), .Y(n15085));
  NOR3X1  g11782(.A(n14962), .B(n14998), .C(n14746), .Y(n15086));
  NOR2X1  g11783(.A(n15086), .B(n15072), .Y(n15087));
  NAND4X1 g11784(.A(n15046), .B(n14963), .C(n14746), .D(n15032), .Y(n15088));
  NAND2X1 g11785(.A(n15088), .B(n15020), .Y(n15089));
  OAI21X1 g11786(.A0(n15087), .A1(n15085), .B0(n15089), .Y(n15090));
  NOR4X1  g11787(.A(n15084), .B(n15071), .C(n15063), .D(n15090), .Y(n15091));
  NAND3X1 g11788(.A(n15091), .B(n15082), .C(n15078), .Y(n15092));
  INVX1   g11789(.A(P1_STATE2_REG_1__SCAN_IN), .Y(n15093));
  AOI21X1 g11790(.A0(n15093), .A1(P1_STATE2_REG_2__SCAN_IN), .B0(n14658), .Y(n15094));
  NOR3X1  g11791(.A(P1_STATE2_REG_0__SCAN_IN), .B(P1_STATE2_REG_1__SCAN_IN), .C(P1_STATE2_REG_3__SCAN_IN), .Y(n15095));
  AOI21X1 g11792(.A0(n15095), .A1(n14658), .B0(n15094), .Y(n15096));
  INVX1   g11793(.A(n15048), .Y(n15097));
  NOR4X1  g11794(.A(n14962), .B(n14998), .C(n14746), .D(n15065), .Y(n15098));
  INVX1   g11795(.A(n15098), .Y(n15099));
  NAND2X1 g11796(.A(n15099), .B(n15097), .Y(n15100));
  OAI21X1 g11797(.A0(n15100), .A1(n15045), .B0(n14812), .Y(n15101));
  NAND3X1 g11798(.A(n15080), .B(n15008), .C(P1_STATE2_REG_0__SCAN_IN), .Y(n15102));
  NAND3X1 g11799(.A(n15066), .B(n14992), .C(n14746), .Y(n15103));
  NOR2X1  g11800(.A(n15103), .B(n14650), .Y(n15104));
  NOR4X1  g11801(.A(n15085), .B(n15046), .C(n14650), .D(n15070), .Y(n15105));
  INVX1   g11802(.A(n14810), .Y(n15106));
  NAND3X1 g11803(.A(n14940), .B(n14806), .C(P1_STATE2_REG_0__SCAN_IN), .Y(n15107));
  NAND2X1 g11804(.A(n15107), .B(n15106), .Y(n15108));
  NOR3X1  g11805(.A(n15108), .B(n15105), .C(n15104), .Y(n15109));
  NAND3X1 g11806(.A(n15109), .B(n15102), .C(n15101), .Y(n15110));
  NAND3X1 g11807(.A(n14800), .B(n14790), .C(n14783), .Y(n15111));
  NAND2X1 g11808(.A(n15111), .B(n14919), .Y(n15112));
  NAND3X1 g11809(.A(n15112), .B(n15042), .C(n14746), .Y(n15113));
  OAI21X1 g11810(.A0(n15113), .A1(n15014), .B0(n15020), .Y(n15114));
  AOI21X1 g11811(.A0(n15114), .A1(n15055), .B0(n14650), .Y(n15115));
  NAND2X1 g11812(.A(n14992), .B(n14846), .Y(n15116));
  NOR4X1  g11813(.A(n15065), .B(n15002), .C(n14801), .D(n15116), .Y(n15117));
  NAND2X1 g11814(.A(n15117), .B(P1_STATE2_REG_0__SCAN_IN), .Y(n15118));
  NOR4X1  g11815(.A(n14984), .B(n14998), .C(n14801), .D(n15070), .Y(n15119));
  OAI21X1 g11816(.A0(n15119), .A1(n15063), .B0(P1_STATE2_REG_0__SCAN_IN), .Y(n15120));
  NOR3X1  g11817(.A(n14962), .B(n14919), .C(n14803), .Y(n15121));
  INVX1   g11818(.A(n15121), .Y(n15122));
  NOR4X1  g11819(.A(n15122), .B(n14991), .C(n14650), .D(n15002), .Y(n15123));
  INVX1   g11820(.A(n14995), .Y(n15124));
  NAND4X1 g11821(.A(n14769), .B(n14806), .C(P1_STATE2_REG_0__SCAN_IN), .D(n15124), .Y(n15125));
  OAI21X1 g11822(.A0(n14807), .A1(n14650), .B0(n15125), .Y(n15126));
  AOI21X1 g11823(.A0(n15126), .A1(n14988), .B0(n15123), .Y(n15127));
  NAND4X1 g11824(.A(n15127), .B(n15120), .C(n15118), .D(n15096), .Y(n15128));
  NOR3X1  g11825(.A(n15128), .B(n15115), .C(n15110), .Y(n15129));
  AOI21X1 g11826(.A0(n15096), .A1(n14670), .B0(n15129), .Y(n15130));
  XOR2X1  g11827(.A(n15130), .B(n15092), .Y(n15131));
  INVX1   g11828(.A(n15131), .Y(n15132));
  NOR2X1  g11829(.A(n15000), .B(n14985), .Y(n15133));
  AOI21X1 g11830(.A0(n15001), .A1(n15133), .B0(n15010), .Y(n15134));
  INVX1   g11831(.A(n15134), .Y(n15135));
  NOR4X1  g11832(.A(n14962), .B(n14919), .C(n14803), .D(n14991), .Y(n15136));
  INVX1   g11833(.A(n15136), .Y(n15137));
  NOR3X1  g11834(.A(n15137), .B(n14990), .C(n14670), .Y(n15138));
  AOI21X1 g11835(.A0(n15135), .A1(n14670), .B0(n15138), .Y(n15139));
  OAI21X1 g11836(.A0(n15132), .A1(n15077), .B0(n15139), .Y(n15140));
  NOR4X1  g11837(.A(n15012), .B(n15006), .C(n14670), .D(n15036), .Y(n15141));
  AOI21X1 g11838(.A0(n15140), .A1(n15038), .B0(n15141), .Y(n15142));
  NAND2X1 g11839(.A(n15130), .B(n15092), .Y(n15143));
  NAND3X1 g11840(.A(n15051), .B(n14992), .C(n14802), .Y(n15144));
  NAND2X1 g11841(.A(n15144), .B(n15127), .Y(n15145));
  INVX1   g11842(.A(n15095), .Y(n15146));
  XOR2X1  g11843(.A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n14658), .Y(n15147));
  NOR2X1  g11844(.A(n15147), .B(n15146), .Y(n15148));
  OAI21X1 g11845(.A0(n15103), .A1(n14650), .B0(n15102), .Y(n15149));
  INVX1   g11846(.A(n14812), .Y(n15150));
  OAI21X1 g11847(.A0(n15097), .A1(n15150), .B0(n15118), .Y(n15151));
  NOR2X1  g11848(.A(n15151), .B(n15149), .Y(n15152));
  NOR4X1  g11849(.A(n14984), .B(n15069), .C(n14650), .D(n15070), .Y(n15153));
  NOR2X1  g11850(.A(n15062), .B(n14650), .Y(n15154));
  INVX1   g11851(.A(P1_STATE2_REG_2__SCAN_IN), .Y(n15155));
  NOR2X1  g11852(.A(P1_STATE2_REG_1__SCAN_IN), .B(n15155), .Y(n15156));
  INVX1   g11853(.A(n15156), .Y(n15157));
  AOI21X1 g11854(.A0(n15157), .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B0(n15148), .Y(n15158));
  NAND3X1 g11855(.A(n15158), .B(n15107), .C(n15106), .Y(n15159));
  AOI21X1 g11856(.A0(n15098), .A1(n14812), .B0(n15159), .Y(n15160));
  NAND2X1 g11857(.A(n15160), .B(n15127), .Y(n15161));
  NOR4X1  g11858(.A(n15154), .B(n15153), .C(n15105), .D(n15161), .Y(n15162));
  AOI21X1 g11859(.A0(n15045), .A1(n14812), .B0(n15115), .Y(n15163));
  NAND3X1 g11860(.A(n15163), .B(n15162), .C(n15152), .Y(n15164));
  OAI21X1 g11861(.A0(n15156), .A1(n14659), .B0(n14657), .Y(n15165));
  OAI21X1 g11862(.A0(n15165), .A1(n15148), .B0(n15164), .Y(n15166));
  XOR2X1  g11863(.A(n15166), .B(n15145), .Y(n15167));
  XOR2X1  g11864(.A(n15167), .B(n15143), .Y(n15168));
  INVX1   g11865(.A(n15168), .Y(n15169));
  XOR2X1  g11866(.A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Y(n15170));
  AOI22X1 g11867(.A0(n15135), .A1(n15170), .B0(n14994), .B1(n14657), .Y(n15171));
  OAI21X1 g11868(.A0(n15169), .A1(n15077), .B0(n15171), .Y(n15172));
  NOR4X1  g11869(.A(n15012), .B(n15006), .C(n14657), .D(n15036), .Y(n15173));
  AOI21X1 g11870(.A0(n15172), .A1(n15038), .B0(n15173), .Y(n15174));
  NAND3X1 g11871(.A(n15174), .B(n15142), .C(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Y(n15175));
  NOR2X1  g11872(.A(n14659), .B(n14658), .Y(n15176));
  NAND2X1 g11873(.A(n15174), .B(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Y(n15177));
  INVX1   g11874(.A(n15166), .Y(n15178));
  NAND2X1 g11875(.A(n15178), .B(n15145), .Y(n15179));
  NOR2X1  g11876(.A(n15178), .B(n15145), .Y(n15180));
  OAI21X1 g11877(.A0(n15180), .A1(n15143), .B0(n15179), .Y(n15181));
  NAND2X1 g11878(.A(n15120), .B(n15118), .Y(n15182));
  INVX1   g11879(.A(n15127), .Y(n15183));
  NOR4X1  g11880(.A(n15182), .B(n15115), .C(n15110), .D(n15183), .Y(n15184));
  XOR2X1  g11881(.A(n15176), .B(n14656), .Y(n15185));
  NOR2X1  g11882(.A(n15185), .B(n15146), .Y(n15186));
  INVX1   g11883(.A(n15186), .Y(n15187));
  AOI21X1 g11884(.A0(n15157), .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B0(n15186), .Y(n15188));
  AOI21X1 g11885(.A0(n15157), .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B0(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Y(n15189));
  AOI22X1 g11886(.A0(n15188), .A1(n15184), .B0(n15187), .B1(n15189), .Y(n15190));
  INVX1   g11887(.A(n15190), .Y(n15191));
  XOR2X1  g11888(.A(n15191), .B(n15181), .Y(n15192));
  NOR2X1  g11889(.A(n15010), .B(n15003), .Y(n15193));
  INVX1   g11890(.A(n15193), .Y(n15194));
  INVX1   g11891(.A(n14896), .Y(n15195));
  NOR3X1  g11892(.A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n14657), .C(n14670), .Y(n15196));
  AOI21X1 g11893(.A0(n15195), .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B0(n15196), .Y(n15197));
  INVX1   g11894(.A(n14994), .Y(n15198));
  XOR2X1  g11895(.A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n14657), .Y(n15199));
  NOR3X1  g11896(.A(n15085), .B(n15000), .C(n14770), .Y(n15200));
  INVX1   g11897(.A(n15200), .Y(n15201));
  OAI22X1 g11898(.A0(n15199), .A1(n15198), .B0(n15197), .B1(n15201), .Y(n15202));
  AOI21X1 g11899(.A0(n15197), .A1(n15194), .B0(n15202), .Y(n15203));
  OAI21X1 g11900(.A0(n15192), .A1(n15077), .B0(n15203), .Y(n15204));
  NOR4X1  g11901(.A(n15012), .B(n15006), .C(n14655), .D(n15036), .Y(n15205));
  AOI21X1 g11902(.A0(n15204), .A1(n15038), .B0(n15205), .Y(n15206));
  NAND2X1 g11903(.A(n15206), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .Y(n15207));
  NAND2X1 g11904(.A(n15207), .B(n15177), .Y(n15208));
  AOI21X1 g11905(.A0(n15176), .A1(n15142), .B0(n15208), .Y(n15209));
  NAND2X1 g11906(.A(n15190), .B(n15181), .Y(n15210));
  NOR2X1  g11907(.A(n15184), .B(n14677), .Y(n15211));
  AOI21X1 g11908(.A0(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B0(n14653), .Y(n15212));
  NOR4X1  g11909(.A(n14656), .B(n14659), .C(n14658), .D(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .Y(n15213));
  NOR2X1  g11910(.A(n14653), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .Y(n15214));
  NOR3X1  g11911(.A(n15214), .B(n15213), .C(n15212), .Y(n15215));
  OAI22X1 g11912(.A0(n15146), .A1(n15215), .B0(n15156), .B1(n14653), .Y(n15216));
  NOR2X1  g11913(.A(n15216), .B(n15211), .Y(n15217));
  XOR2X1  g11914(.A(n15217), .B(n15210), .Y(n15218));
  INVX1   g11915(.A(n15218), .Y(n15219));
  OAI21X1 g11916(.A0(n14657), .A1(n14670), .B0(n14655), .Y(n15220));
  AOI22X1 g11917(.A0(n15195), .A1(n14685), .B0(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(n15220), .Y(n15221));
  AOI21X1 g11918(.A0(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B0(n14677), .Y(n15222));
  AOI21X1 g11919(.A0(n14895), .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B0(n15222), .Y(n15223));
  NOR3X1  g11920(.A(n15223), .B(n15137), .C(n14990), .Y(n15224));
  NAND3X1 g11921(.A(n14677), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Y(n15225));
  NOR3X1  g11922(.A(n14655), .B(n14657), .C(n14670), .Y(n15226));
  OAI22X1 g11923(.A0(n15225), .A1(n14670), .B0(n14677), .B1(n15226), .Y(n15227));
  AOI21X1 g11924(.A0(n15227), .A1(n15200), .B0(n15224), .Y(n15228));
  INVX1   g11925(.A(n15228), .Y(n15229));
  AOI21X1 g11926(.A0(n15221), .A1(n15194), .B0(n15229), .Y(n15230));
  OAI21X1 g11927(.A0(n15219), .A1(n15077), .B0(n15230), .Y(n15231));
  NOR4X1  g11928(.A(n15012), .B(n15006), .C(n14677), .D(n15036), .Y(n15232));
  AOI21X1 g11929(.A0(n15231), .A1(n15038), .B0(n15232), .Y(n15233));
  OAI22X1 g11930(.A0(n15206), .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B0(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B1(n15233), .Y(n15234));
  AOI21X1 g11931(.A0(n15209), .A1(n15175), .B0(n15234), .Y(n15235));
  INVX1   g11932(.A(n15233), .Y(n15236));
  NOR3X1  g11933(.A(n15137), .B(n14990), .C(n14650), .Y(n15237));
  NOR2X1  g11934(.A(n15237), .B(n15123), .Y(n15238));
  NOR2X1  g11935(.A(n15238), .B(n14651), .Y(n15239));
  INVX1   g11936(.A(n15239), .Y(n15240));
  INVX1   g11937(.A(n15181), .Y(n15241));
  NOR3X1  g11938(.A(n15217), .B(n15191), .C(n15241), .Y(n15242));
  XOR2X1  g11939(.A(n15242), .B(n15240), .Y(n15243));
  NOR3X1  g11940(.A(n15243), .B(n15037), .C(n15028), .Y(n15244));
  AOI21X1 g11941(.A0(n15037), .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B0(n15244), .Y(n15245));
  INVX1   g11942(.A(n15245), .Y(n15246));
  OAI22X1 g11943(.A0(n15236), .A1(n14653), .B0(n14666), .B1(n15246), .Y(n15247));
  NOR2X1  g11944(.A(n15247), .B(n15235), .Y(n15248));
  NOR2X1  g11945(.A(n15093), .B(P1_FLUSH_REG_SCAN_IN), .Y(n15249));
  INVX1   g11946(.A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .Y(n15250));
  INVX1   g11947(.A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .Y(n15251));
  NOR2X1  g11948(.A(n15251), .B(n15250), .Y(n15252));
  NOR2X1  g11949(.A(n15251), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .Y(n15253));
  INVX1   g11950(.A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .Y(n15255));
  XOR2X1  g11951(.A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n15255), .Y(n15256));
  INVX1   g11952(.A(n15256), .Y(n15257));
  NOR2X1  g11953(.A(n15255), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .Y(n15258));
  AOI21X1 g11954(.A0(n15257), .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B0(n15258), .Y(n15259));
  NOR3X1  g11955(.A(n15259), .B(n15251), .C(n15093), .Y(n15260));
  AOI22X1 g11956(.A0(n15249), .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B0(P1_FLUSH_REG_SCAN_IN), .B1(n15260), .Y(n15261));
  OAI21X1 g11957(.A0(n15206), .A1(P1_STATE2_REG_1__SCAN_IN), .B0(n15261), .Y(n15262));
  INVX1   g11958(.A(n15262), .Y(n15263));
  AOI22X1 g11959(.A0(n15246), .A1(n15093), .B0(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B1(n15249), .Y(n15264));
  AOI22X1 g11960(.A0(n15236), .A1(n15093), .B0(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(n15249), .Y(n15265));
  OAI21X1 g11961(.A0(n15265), .A1(n15263), .B0(n15264), .Y(n15266));
  NAND2X1 g11962(.A(n15246), .B(n14666), .Y(n15267));
  INVX1   g11963(.A(n15007), .Y(n15268));
  OAI21X1 g11964(.A0(n14987), .A1(n15268), .B0(n14806), .Y(n15269));
  NOR2X1  g11965(.A(n15007), .B(n14769), .Y(n15270));
  INVX1   g11966(.A(n15270), .Y(n15271));
  NOR2X1  g11967(.A(n15030), .B(n14770), .Y(n15272));
  OAI21X1 g11968(.A0(n15272), .A1(n15137), .B0(n14707), .Y(n15273));
  NAND3X1 g11969(.A(n15273), .B(n15271), .C(n15269), .Y(n15274));
  NOR2X1  g11970(.A(n14995), .B(P1_STATE_REG_0__SCAN_IN), .Y(n15275));
  INVX1   g11971(.A(n15275), .Y(n15276));
  NAND3X1 g11972(.A(n15002), .B(n15276), .C(n14807), .Y(n15277));
  AOI21X1 g11973(.A0(n15277), .A1(n14550), .B0(n15274), .Y(n15278));
  OAI21X1 g11974(.A0(P1_FLUSH_REG_SCAN_IN), .A1(P1_MORE_REG_SCAN_IN), .B0(n15278), .Y(n15279));
  NOR4X1  g11975(.A(n14985), .B(n14940), .C(n14803), .D(n14993), .Y(n15280));
  NOR4X1  g11976(.A(n14940), .B(n14846), .C(n14707), .D(n14985), .Y(n15281));
  OAI21X1 g11977(.A0(n15280), .A1(n15068), .B0(n15281), .Y(n15282));
  NOR2X1  g11978(.A(n15003), .B(n14994), .Y(n15283));
  NAND2X1 g11979(.A(n15283), .B(n15282), .Y(n15284));
  NAND3X1 g11980(.A(n15284), .B(n14890), .C(n14887), .Y(n15285));
  INVX1   g11981(.A(n15030), .Y(n15286));
  AOI22X1 g11982(.A0(n15027), .A1(n15286), .B0(n15010), .B1(n15007), .Y(n15287));
  AOI21X1 g11983(.A0(n15287), .A1(n15285), .B0(n14962), .Y(n15288));
  AOI21X1 g11984(.A0(n14890), .A1(n14887), .B0(n14707), .Y(n15289));
  AOI21X1 g11985(.A0(n15289), .A1(n15280), .B0(n15288), .Y(n15290));
  NAND3X1 g11986(.A(n15290), .B(n15279), .C(n15267), .Y(n15291));
  NOR4X1  g11987(.A(n15266), .B(n15248), .C(P1_STATE2_REG_1__SCAN_IN), .D(n15291), .Y(n15292));
  AOI21X1 g11988(.A0(n14890), .A1(n14887), .B0(n15276), .Y(n15293));
  AOI21X1 g11989(.A0(READY11_REG_SCAN_IN), .A1(READY1), .B0(P1_STATEBS16_REG_SCAN_IN), .Y(n15294));
  INVX1   g11990(.A(n15294), .Y(n15295));
  NOR3X1  g11991(.A(n15295), .B(n14987), .C(n15021), .Y(n15296));
  NOR3X1  g11992(.A(n15093), .B(n14546), .C(n14545), .Y(n15297));
  OAI21X1 g11993(.A0(n15297), .A1(P1_STATE2_REG_0__SCAN_IN), .B0(P1_STATE2_REG_2__SCAN_IN), .Y(n15298));
  AOI21X1 g11994(.A0(n15296), .A1(n15293), .B0(n15298), .Y(n15299));
  AOI21X1 g11995(.A0(n15299), .A1(n15292), .B0(n14650), .Y(n15300));
  NOR3X1  g11996(.A(n15291), .B(n15266), .C(n15248), .Y(n15301));
  NAND3X1 g11997(.A(P1_STATE2_REG_0__SCAN_IN), .B(P1_STATE2_REG_1__SCAN_IN), .C(P1_STATE2_REG_2__SCAN_IN), .Y(n15302));
  OAI21X1 g11998(.A0(n15300), .A1(n14649), .B0(n15302), .Y(P1_U3466));
  OAI21X1 g11999(.A0(n14549), .A1(P1_STATE2_REG_2__SCAN_IN), .B0(P1_STATE2_REG_0__SCAN_IN), .Y(n15304));
  INVX1   g12000(.A(P1_STATEBS16_REG_SCAN_IN), .Y(n15305));
  AOI21X1 g12001(.A0(n14650), .A1(n15305), .B0(n15093), .Y(n15306));
  AOI21X1 g12002(.A0(n15306), .A1(n15304), .B0(n15156), .Y(n15307));
  OAI21X1 g12003(.A0(n15300), .A1(n15155), .B0(n15307), .Y(P1_U3163));
  NOR2X1  g12004(.A(P1_STATE2_REG_1__SCAN_IN), .B(P1_STATE2_REG_3__SCAN_IN), .Y(n15309));
  NAND3X1 g12005(.A(n15300), .B(n15309), .C(n14550), .Y(n15310));
  OAI21X1 g12006(.A0(n15292), .A1(n14650), .B0(n15299), .Y(n15311));
  INVX1   g12007(.A(n15311), .Y(n15312));
  NOR4X1  g12008(.A(P1_STATE2_REG_2__SCAN_IN), .B(n14546), .C(n14545), .D(n14650), .Y(n15313));
  OAI21X1 g12009(.A0(n15313), .A1(n15312), .B0(P1_STATE2_REG_1__SCAN_IN), .Y(n15314));
  NOR4X1  g12010(.A(n15093), .B(P1_STATE2_REG_2__SCAN_IN), .C(P1_STATEBS16_REG_SCAN_IN), .D(P1_STATE2_REG_0__SCAN_IN), .Y(n15315));
  NOR3X1  g12011(.A(n14650), .B(P1_STATE2_REG_1__SCAN_IN), .C(n15155), .Y(n15316));
  AOI21X1 g12012(.A0(n15316), .A1(n15311), .B0(n15315), .Y(n15317));
  NAND3X1 g12013(.A(n15317), .B(n15314), .C(n15310), .Y(P1_U3162));
  INVX1   g12014(.A(n15264), .Y(n15319));
  NOR2X1  g12015(.A(n15142), .B(P1_STATE2_REG_1__SCAN_IN), .Y(n15320));
  NOR2X1  g12016(.A(n15174), .B(P1_STATE2_REG_1__SCAN_IN), .Y(n15321));
  INVX1   g12017(.A(P1_FLUSH_REG_SCAN_IN), .Y(n15322));
  INVX1   g12018(.A(n15252), .Y(n15323));
  INVX1   g12019(.A(n15253), .Y(n15324));
  AOI21X1 g12020(.A0(n15324), .A1(n15323), .B0(n15093), .Y(n15325));
  NAND2X1 g12021(.A(n15259), .B(n15325), .Y(n15326));
  NOR2X1  g12022(.A(n15326), .B(n15322), .Y(n15327));
  NOR3X1  g12023(.A(n15253), .B(n15252), .C(n15093), .Y(n15328));
  NAND2X1 g12024(.A(n15328), .B(P1_FLUSH_REG_SCAN_IN), .Y(n15329));
  OAI21X1 g12025(.A0(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B0(n15249), .Y(n15330));
  NAND2X1 g12026(.A(n15330), .B(n15329), .Y(n15331));
  NOR4X1  g12027(.A(n15327), .B(n15321), .C(n15320), .D(n15331), .Y(n15332));
  NOR3X1  g12028(.A(n15332), .B(n15265), .C(n15263), .Y(n15333));
  NOR4X1  g12029(.A(n15319), .B(n15093), .C(n15155), .D(n15333), .Y(n15334));
  OAI21X1 g12030(.A0(n15334), .A1(n15312), .B0(P1_STATE2_REG_0__SCAN_IN), .Y(n15335));
  AOI21X1 g12031(.A0(n14890), .A1(n14887), .B0(n14649), .Y(n15336));
  NAND3X1 g12032(.A(n15336), .B(n15093), .C(n15155), .Y(n15337));
  NAND3X1 g12033(.A(n15337), .B(n15311), .C(n14650), .Y(n15338));
  INVX1   g12034(.A(n15316), .Y(n15339));
  NOR2X1  g12035(.A(n15339), .B(n15301), .Y(n15340));
  NOR4X1  g12036(.A(P1_STATE2_REG_1__SCAN_IN), .B(P1_STATE2_REG_2__SCAN_IN), .C(n14649), .D(n14650), .Y(n15341));
  NOR3X1  g12037(.A(n15341), .B(n15340), .C(n15313), .Y(n15342));
  NAND3X1 g12038(.A(n15342), .B(n15338), .C(n15335), .Y(P1_U3161));
  INVX1   g12039(.A(n15336), .Y(n15344));
  XOR2X1  g12040(.A(P1_STATE2_REG_1__SCAN_IN), .B(n15155), .Y(n15345));
  AOI21X1 g12041(.A0(n15345), .A1(n15344), .B0(P1_STATE2_REG_0__SCAN_IN), .Y(n15346));
  NOR4X1  g12042(.A(n14656), .B(n14659), .C(n14658), .D(n14653), .Y(n15347));
  NOR2X1  g12043(.A(n15219), .B(n15192), .Y(n15348));
  NOR2X1  g12044(.A(n15169), .B(n15132), .Y(n15349));
  AOI21X1 g12045(.A0(n15349), .A1(n15348), .B0(n15347), .Y(n15350));
  NOR3X1  g12046(.A(P1_STATE2_REG_2__SCAN_IN), .B(P1_STATE2_REG_3__SCAN_IN), .C(P1_STATEBS16_REG_SCAN_IN), .Y(n15351));
  NOR3X1  g12047(.A(P1_STATE2_REG_2__SCAN_IN), .B(P1_STATE2_REG_3__SCAN_IN), .C(n15305), .Y(n15352));
  INVX1   g12048(.A(n15352), .Y(n15353));
  INVX1   g12049(.A(n15346), .Y(n15354));
  NOR4X1  g12050(.A(n14655), .B(n14657), .C(n14670), .D(n14677), .Y(n15355));
  AOI22X1 g12051(.A0(n15355), .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B0(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(n14673), .Y(n15357));
  NOR4X1  g12052(.A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C(n14670), .D(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n15359));
  AOI22X1 g12053(.A0(n14674), .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B0(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(n15359), .Y(n15360));
  NOR4X1  g12054(.A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n14657), .C(n14670), .D(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n15361));
  NOR4X1  g12055(.A(n14655), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .D(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n15362));
  AOI22X1 g12056(.A0(n15361), .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B0(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(n15362), .Y(n15363));
  NOR4X1  g12057(.A(n14655), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C(n14670), .D(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n15365));
  AOI22X1 g12058(.A0(n14703), .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B0(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(n15365), .Y(n15366));
  NAND4X1 g12059(.A(n15363), .B(n15360), .C(n15357), .D(n15366), .Y(n15367));
  AOI22X1 g12060(.A0(n14680), .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B0(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(n14907), .Y(n15370));
  NOR4X1  g12061(.A(n14655), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C(n14670), .D(n14677), .Y(n15372));
  AOI22X1 g12062(.A0(n14704), .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B0(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(n15372), .Y(n15373));
  NOR4X1  g12063(.A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .D(n14677), .Y(n15375));
  AOI22X1 g12064(.A0(n14671), .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B0(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(n15375), .Y(n15376));
  NOR4X1  g12065(.A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C(n14670), .D(n14677), .Y(n15378));
  AOI22X1 g12066(.A0(n14682), .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B0(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(n15378), .Y(n15379));
  NAND4X1 g12067(.A(n15376), .B(n15373), .C(n15370), .D(n15379), .Y(n15380));
  NOR2X1  g12068(.A(n15380), .B(n15367), .Y(n15381));
  NOR3X1  g12069(.A(n15381), .B(n14846), .C(n14650), .Y(n15382));
  AOI22X1 g12070(.A0(n15355), .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B0(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(n14673), .Y(n15384));
  AOI22X1 g12071(.A0(n14674), .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B0(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(n15359), .Y(n15385));
  AOI22X1 g12072(.A0(n15361), .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B0(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(n15362), .Y(n15386));
  AOI22X1 g12073(.A0(n14703), .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B0(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(n15365), .Y(n15387));
  NAND4X1 g12074(.A(n15386), .B(n15385), .C(n15384), .D(n15387), .Y(n15388));
  AOI22X1 g12075(.A0(n14680), .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B0(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(n14907), .Y(n15389));
  AOI22X1 g12076(.A0(n14704), .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B0(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(n15372), .Y(n15390));
  AOI22X1 g12077(.A0(n14671), .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B0(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(n15375), .Y(n15391));
  AOI22X1 g12078(.A0(n14682), .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B0(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(n15378), .Y(n15392));
  NAND4X1 g12079(.A(n15391), .B(n15390), .C(n15389), .D(n15392), .Y(n15393));
  NOR2X1  g12080(.A(n15393), .B(n15388), .Y(n15394));
  NOR3X1  g12081(.A(n15394), .B(n14806), .C(n14650), .Y(n15395));
  NOR4X1  g12082(.A(n14745), .B(n14716), .C(n14710), .D(n15381), .Y(n15396));
  INVX1   g12083(.A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .Y(n15397));
  NOR4X1  g12084(.A(n14707), .B(n14650), .C(n15397), .D(n14746), .Y(n15398));
  NOR4X1  g12085(.A(n15396), .B(n15395), .C(n14650), .D(n15398), .Y(n15399));
  INVX1   g12086(.A(n15394), .Y(n15400));
  NOR4X1  g12087(.A(n14716), .B(n14710), .C(n14650), .D(n14745), .Y(n15401));
  NAND3X1 g12088(.A(n15400), .B(n15381), .C(n15401), .Y(n15402));
  OAI21X1 g12089(.A0(n15400), .A1(n16815), .B0(n15402), .Y(n15403));
  AOI21X1 g12090(.A0(n15131), .A1(n14650), .B0(n15403), .Y(n15404));
  XOR2X1  g12091(.A(n15404), .B(n15382), .Y(n15405));
  XOR2X1  g12092(.A(n15405), .B(n15399), .Y(n15406));
  XOR2X1  g12093(.A(n15406), .B(n16815), .Y(n15407));
  INVX1   g12094(.A(n15407), .Y(n15408));
  OAI21X1 g12095(.A0(n15405), .A1(n15399), .B0(n16815), .Y(n15411));
  INVX1   g12096(.A(n15381), .Y(n15412));
  NOR3X1  g12097(.A(n15412), .B(n14846), .C(n14650), .Y(n15413));
  INVX1   g12098(.A(n15413), .Y(n15414));
  AOI22X1 g12099(.A0(n15355), .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B0(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(n14673), .Y(n15415));
  AOI22X1 g12100(.A0(n14674), .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B0(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(n15359), .Y(n15416));
  AOI22X1 g12101(.A0(n15361), .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B0(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(n15362), .Y(n15417));
  AOI22X1 g12102(.A0(n14703), .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B0(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(n15365), .Y(n15418));
  NAND4X1 g12103(.A(n15417), .B(n15416), .C(n15415), .D(n15418), .Y(n15419));
  AOI22X1 g12104(.A0(n14680), .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B0(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(n14907), .Y(n15420));
  AOI22X1 g12105(.A0(n14704), .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B0(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(n15372), .Y(n15421));
  AOI22X1 g12106(.A0(n14671), .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B0(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(n15375), .Y(n15422));
  AOI22X1 g12107(.A0(n14682), .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B0(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(n15378), .Y(n15423));
  NAND4X1 g12108(.A(n15422), .B(n15421), .C(n15420), .D(n15423), .Y(n15424));
  NOR2X1  g12109(.A(n15424), .B(n15419), .Y(n15425));
  NAND3X1 g12110(.A(n15425), .B(n15412), .C(n15401), .Y(n15426));
  OAI21X1 g12111(.A0(n15425), .A1(n15414), .B0(n15426), .Y(n15427));
  AOI21X1 g12112(.A0(n15168), .A1(n14650), .B0(n15427), .Y(n15428));
  XOR2X1  g12113(.A(n15428), .B(n15382), .Y(n15429));
  INVX1   g12114(.A(n14824), .Y(n15430));
  AOI22X1 g12115(.A0(n15401), .A1(n15381), .B0(n14818), .B1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .Y(n15431));
  OAI21X1 g12116(.A0(n15425), .A1(n15430), .B0(n15431), .Y(n15432));
  XOR2X1  g12117(.A(n15432), .B(n15429), .Y(n15433));
  XOR2X1  g12118(.A(n15433), .B(n15411), .Y(n15434));
  AOI22X1 g12119(.A0(n15355), .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B0(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(n14673), .Y(n15435));
  AOI22X1 g12120(.A0(n14674), .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B0(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(n15359), .Y(n15436));
  AOI22X1 g12121(.A0(n15361), .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B0(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(n15362), .Y(n15437));
  AOI22X1 g12122(.A0(n14703), .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B0(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(n15365), .Y(n15438));
  NAND4X1 g12123(.A(n15437), .B(n15436), .C(n15435), .D(n15438), .Y(n15439));
  AOI22X1 g12124(.A0(n14680), .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B0(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(n14907), .Y(n15440));
  AOI22X1 g12125(.A0(n14704), .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B0(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(n15372), .Y(n15441));
  AOI22X1 g12126(.A0(n14671), .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B0(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(n15375), .Y(n15442));
  AOI22X1 g12127(.A0(n14682), .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B0(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(n15378), .Y(n15443));
  NAND4X1 g12128(.A(n15442), .B(n15441), .C(n15440), .D(n15443), .Y(n15444));
  NOR2X1  g12129(.A(n15444), .B(n15439), .Y(n15445));
  INVX1   g12130(.A(n15445), .Y(n15446));
  AOI22X1 g12131(.A0(n14824), .A1(n15446), .B0(n14818), .B1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .Y(n15447));
  NOR4X1  g12132(.A(n15412), .B(n14846), .C(n14650), .D(n15445), .Y(n15448));
  AOI21X1 g12133(.A0(n15445), .A1(n15382), .B0(n15448), .Y(n15449));
  OAI21X1 g12134(.A0(n15192), .A1(P1_STATE2_REG_0__SCAN_IN), .B0(n15449), .Y(n15450));
  XOR2X1  g12135(.A(n15450), .B(n16815), .Y(n15451));
  XOR2X1  g12136(.A(n15451), .B(n15447), .Y(n15452));
  INVX1   g12137(.A(n15432), .Y(n15453));
  NOR2X1  g12138(.A(n15453), .B(n15429), .Y(n15454));
  INVX1   g12139(.A(n15429), .Y(n15455));
  NOR2X1  g12140(.A(n15432), .B(n15455), .Y(n15456));
  INVX1   g12141(.A(n15456), .Y(n15457));
  AOI21X1 g12142(.A0(n15457), .A1(n15411), .B0(n15454), .Y(n15458));
  XOR2X1  g12143(.A(n15458), .B(n15452), .Y(n15459));
  AOI22X1 g12144(.A0(n15355), .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B0(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(n14673), .Y(n15460));
  AOI22X1 g12145(.A0(n14674), .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B0(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(n15359), .Y(n15461));
  AOI22X1 g12146(.A0(n15361), .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B0(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(n15362), .Y(n15462));
  AOI22X1 g12147(.A0(n14703), .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B0(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(n15365), .Y(n15463));
  NAND4X1 g12148(.A(n15462), .B(n15461), .C(n15460), .D(n15463), .Y(n15464));
  AOI22X1 g12149(.A0(n14680), .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B0(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(n14907), .Y(n15465));
  AOI22X1 g12150(.A0(n14704), .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B0(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(n15372), .Y(n15466));
  AOI22X1 g12151(.A0(n14671), .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B0(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(n15375), .Y(n15467));
  AOI22X1 g12152(.A0(n14682), .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B0(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(n15378), .Y(n15468));
  NAND4X1 g12153(.A(n15467), .B(n15466), .C(n15465), .D(n15468), .Y(n15469));
  NOR2X1  g12154(.A(n15469), .B(n15464), .Y(n15470));
  INVX1   g12155(.A(n15470), .Y(n15471));
  AOI22X1 g12156(.A0(n14824), .A1(n15471), .B0(n14818), .B1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .Y(n15472));
  NAND3X1 g12157(.A(n15471), .B(n15381), .C(n15401), .Y(n15473));
  OAI21X1 g12158(.A0(n15471), .A1(n16815), .B0(n15473), .Y(n15474));
  AOI21X1 g12159(.A0(n15218), .A1(n14650), .B0(n15474), .Y(n15475));
  XOR2X1  g12160(.A(n15475), .B(n15382), .Y(n15476));
  XOR2X1  g12161(.A(n15476), .B(n15472), .Y(n15477));
  INVX1   g12162(.A(n15447), .Y(n15478));
  INVX1   g12163(.A(n15451), .Y(n15479));
  NAND2X1 g12164(.A(n15479), .B(n15478), .Y(n15480));
  NOR2X1  g12165(.A(n15479), .B(n15478), .Y(n15481));
  OAI21X1 g12166(.A0(n15458), .A1(n15481), .B0(n15480), .Y(n15482));
  XOR2X1  g12167(.A(n15482), .B(n15477), .Y(n15483));
  INVX1   g12168(.A(n15483), .Y(n15484));
  NOR4X1  g12169(.A(n15459), .B(n15434), .C(n15408), .D(n15484), .Y(n15485));
  NOR2X1  g12170(.A(n15434), .B(n15407), .Y(n15486));
  INVX1   g12171(.A(n15486), .Y(n15487));
  NOR3X1  g12172(.A(n15484), .B(n15459), .C(n15487), .Y(n15488));
  NOR4X1  g12173(.A(n15485), .B(n15354), .C(n15353), .D(n15488), .Y(n15489));
  OAI21X1 g12174(.A0(n15489), .A1(n15351), .B0(n15350), .Y(n15490));
  INVX1   g12175(.A(n15347), .Y(n15491));
  NOR2X1  g12176(.A(n15215), .B(n15185), .Y(n15492));
  NOR2X1  g12177(.A(n14659), .B(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Y(n15493));
  AOI21X1 g12178(.A0(n15493), .A1(n15492), .B0(n15347), .Y(n15494));
  AOI22X1 g12179(.A0(n15491), .A1(P1_STATE2_REG_3__SCAN_IN), .B0(P1_STATE2_REG_2__SCAN_IN), .B1(n15494), .Y(n15495));
  NAND3X1 g12180(.A(n15495), .B(n15490), .C(n15346), .Y(n15496));
  NAND2X1 g12181(.A(n15496), .B(P1_INSTQUEUE_REG_15__7__SCAN_IN), .Y(n15497));
  NOR2X1  g12182(.A(n3070), .B(n9741), .Y(n15498));
  AOI21X1 g12183(.A0(n3070), .A1(DATAI_7_), .B0(n15498), .Y(n15499));
  NOR2X1  g12184(.A(n15499), .B(n15354), .Y(n15500));
  NOR3X1  g12185(.A(n15488), .B(n15485), .C(n15353), .Y(n15501));
  NOR2X1  g12186(.A(n15501), .B(n15351), .Y(n15502));
  OAI22X1 g12187(.A0(n15494), .A1(n15155), .B0(n15350), .B1(n15502), .Y(n15503));
  NAND2X1 g12188(.A(n15503), .B(n15500), .Y(n15504));
  NOR2X1  g12189(.A(n3070), .B(n9844), .Y(n15505));
  AOI21X1 g12190(.A0(n3070), .A1(DATAI_31_), .B0(n15505), .Y(n15506));
  NOR3X1  g12191(.A(n15506), .B(n15354), .C(n15353), .Y(n15507));
  INVX1   g12192(.A(n15488), .Y(n15508));
  NOR2X1  g12193(.A(n3070), .B(n9849), .Y(n15509));
  AOI21X1 g12194(.A0(n3070), .A1(DATAI_23_), .B0(n15509), .Y(n15510));
  INVX1   g12195(.A(n15510), .Y(n15511));
  NAND3X1 g12196(.A(n15511), .B(n15346), .C(n15352), .Y(n15512));
  NAND3X1 g12197(.A(n15346), .B(n15042), .C(P1_STATE2_REG_3__SCAN_IN), .Y(n15513));
  OAI22X1 g12198(.A0(n15512), .A1(n15508), .B0(n15491), .B1(n15513), .Y(n15514));
  AOI21X1 g12199(.A0(n15507), .A1(n15485), .B0(n15514), .Y(n15515));
  NAND3X1 g12200(.A(n15515), .B(n15504), .C(n15497), .Y(P1_U3160));
  NAND2X1 g12201(.A(n15496), .B(P1_INSTQUEUE_REG_15__6__SCAN_IN), .Y(n15517));
  NOR2X1  g12202(.A(n3070), .B(n9858), .Y(n15518));
  AOI21X1 g12203(.A0(n3070), .A1(DATAI_6_), .B0(n15518), .Y(n15519));
  NOR2X1  g12204(.A(n15519), .B(n15354), .Y(n15520));
  NAND2X1 g12205(.A(n15520), .B(n15503), .Y(n15521));
  NOR2X1  g12206(.A(n3070), .B(n9864), .Y(n15522));
  AOI21X1 g12207(.A0(n3070), .A1(DATAI_30_), .B0(n15522), .Y(n15523));
  NOR3X1  g12208(.A(n15523), .B(n15354), .C(n15353), .Y(n15524));
  NAND2X1 g12209(.A(n15524), .B(n15485), .Y(n15525));
  NOR2X1  g12210(.A(n3070), .B(n9868), .Y(n15526));
  AOI21X1 g12211(.A0(n3070), .A1(DATAI_22_), .B0(n15526), .Y(n15527));
  NOR3X1  g12212(.A(n15527), .B(n15354), .C(n15353), .Y(n15528));
  NOR3X1  g12213(.A(n15354), .B(n14919), .C(n14649), .Y(n15529));
  AOI22X1 g12214(.A0(n15528), .A1(n15488), .B0(n15347), .B1(n15529), .Y(n15530));
  NAND4X1 g12215(.A(n15525), .B(n15521), .C(n15517), .D(n15530), .Y(P1_U3159));
  NAND2X1 g12216(.A(n15496), .B(P1_INSTQUEUE_REG_15__5__SCAN_IN), .Y(n15532));
  NOR2X1  g12217(.A(n3070), .B(n9877), .Y(n15533));
  AOI21X1 g12218(.A0(n3070), .A1(DATAI_5_), .B0(n15533), .Y(n15534));
  NOR2X1  g12219(.A(n15534), .B(n15354), .Y(n15535));
  NAND2X1 g12220(.A(n15535), .B(n15503), .Y(n15536));
  NOR2X1  g12221(.A(n3070), .B(n9883), .Y(n15537));
  AOI21X1 g12222(.A0(n3070), .A1(DATAI_29_), .B0(n15537), .Y(n15538));
  NOR3X1  g12223(.A(n15538), .B(n15354), .C(n15353), .Y(n15539));
  NAND2X1 g12224(.A(n15539), .B(n15485), .Y(n15540));
  NOR2X1  g12225(.A(n3070), .B(n9887), .Y(n15541));
  AOI21X1 g12226(.A0(n3070), .A1(DATAI_21_), .B0(n15541), .Y(n15542));
  NOR3X1  g12227(.A(n15542), .B(n15354), .C(n15353), .Y(n15543));
  NOR3X1  g12228(.A(n15354), .B(n14808), .C(n14649), .Y(n15544));
  AOI22X1 g12229(.A0(n15543), .A1(n15488), .B0(n15347), .B1(n15544), .Y(n15545));
  NAND4X1 g12230(.A(n15540), .B(n15536), .C(n15532), .D(n15545), .Y(P1_U3158));
  NAND2X1 g12231(.A(n15496), .B(P1_INSTQUEUE_REG_15__4__SCAN_IN), .Y(n15547));
  NOR2X1  g12232(.A(n3070), .B(n9896), .Y(n15548));
  AOI21X1 g12233(.A0(n3070), .A1(DATAI_4_), .B0(n15548), .Y(n15549));
  NOR2X1  g12234(.A(n15549), .B(n15354), .Y(n15550));
  NAND2X1 g12235(.A(n15550), .B(n15503), .Y(n15551));
  NOR2X1  g12236(.A(n3070), .B(n9902), .Y(n15552));
  AOI21X1 g12237(.A0(n3070), .A1(DATAI_28_), .B0(n15552), .Y(n15553));
  NOR3X1  g12238(.A(n15553), .B(n15354), .C(n15353), .Y(n15554));
  NAND2X1 g12239(.A(n15554), .B(n15485), .Y(n15555));
  NOR2X1  g12240(.A(n3070), .B(n9906), .Y(n15556));
  AOI21X1 g12241(.A0(n3070), .A1(DATAI_20_), .B0(n15556), .Y(n15557));
  NOR3X1  g12242(.A(n15557), .B(n15354), .C(n15353), .Y(n15558));
  NOR3X1  g12243(.A(n15354), .B(n14746), .C(n14649), .Y(n15559));
  AOI22X1 g12244(.A0(n15558), .A1(n15488), .B0(n15347), .B1(n15559), .Y(n15560));
  NAND4X1 g12245(.A(n15555), .B(n15551), .C(n15547), .D(n15560), .Y(P1_U3157));
  NAND2X1 g12246(.A(n15496), .B(P1_INSTQUEUE_REG_15__3__SCAN_IN), .Y(n15562));
  NOR2X1  g12247(.A(n3070), .B(n9915), .Y(n15563));
  AOI21X1 g12248(.A0(n3070), .A1(DATAI_3_), .B0(n15563), .Y(n15564));
  NOR2X1  g12249(.A(n15564), .B(n15354), .Y(n15565));
  NAND2X1 g12250(.A(n15565), .B(n15503), .Y(n15566));
  NOR2X1  g12251(.A(n3070), .B(n9921), .Y(n15567));
  AOI21X1 g12252(.A0(n3070), .A1(DATAI_27_), .B0(n15567), .Y(n15568));
  NOR3X1  g12253(.A(n15568), .B(n15354), .C(n15353), .Y(n15569));
  NOR2X1  g12254(.A(n3070), .B(n9925), .Y(n15570));
  AOI21X1 g12255(.A0(n3070), .A1(DATAI_19_), .B0(n15570), .Y(n15571));
  INVX1   g12256(.A(n15571), .Y(n15572));
  NAND3X1 g12257(.A(n15572), .B(n15346), .C(n15352), .Y(n15573));
  NAND3X1 g12258(.A(n15346), .B(n15024), .C(P1_STATE2_REG_3__SCAN_IN), .Y(n15574));
  OAI22X1 g12259(.A0(n15573), .A1(n15508), .B0(n15491), .B1(n15574), .Y(n15575));
  AOI21X1 g12260(.A0(n15569), .A1(n15485), .B0(n15575), .Y(n15576));
  NAND3X1 g12261(.A(n15576), .B(n15566), .C(n15562), .Y(P1_U3156));
  NAND2X1 g12262(.A(n15496), .B(P1_INSTQUEUE_REG_15__2__SCAN_IN), .Y(n15578));
  NOR2X1  g12263(.A(n3070), .B(n9934), .Y(n15579));
  AOI21X1 g12264(.A0(n3070), .A1(DATAI_2_), .B0(n15579), .Y(n15580));
  NOR2X1  g12265(.A(n15580), .B(n15354), .Y(n15581));
  NAND2X1 g12266(.A(n15581), .B(n15503), .Y(n15582));
  NOR2X1  g12267(.A(n3070), .B(n9940), .Y(n15583));
  AOI21X1 g12268(.A0(n3070), .A1(DATAI_26_), .B0(n15583), .Y(n15584));
  NOR3X1  g12269(.A(n15584), .B(n15354), .C(n15353), .Y(n15585));
  NOR2X1  g12270(.A(n3070), .B(n9944), .Y(n15586));
  AOI21X1 g12271(.A0(n3070), .A1(DATAI_18_), .B0(n15586), .Y(n15587));
  INVX1   g12272(.A(n15587), .Y(n15588));
  NAND3X1 g12273(.A(n15588), .B(n15346), .C(n15352), .Y(n15589));
  NAND3X1 g12274(.A(n15346), .B(n14985), .C(P1_STATE2_REG_3__SCAN_IN), .Y(n15590));
  OAI22X1 g12275(.A0(n15589), .A1(n15508), .B0(n15491), .B1(n15590), .Y(n15591));
  AOI21X1 g12276(.A0(n15585), .A1(n15485), .B0(n15591), .Y(n15592));
  NAND3X1 g12277(.A(n15592), .B(n15582), .C(n15578), .Y(P1_U3155));
  NAND2X1 g12278(.A(n15496), .B(P1_INSTQUEUE_REG_15__1__SCAN_IN), .Y(n15594));
  NOR2X1  g12279(.A(n3070), .B(n9953), .Y(n15595));
  AOI21X1 g12280(.A0(n3070), .A1(DATAI_1_), .B0(n15595), .Y(n15596));
  NOR2X1  g12281(.A(n15596), .B(n15354), .Y(n15597));
  NAND2X1 g12282(.A(n15597), .B(n15503), .Y(n15598));
  NOR2X1  g12283(.A(n3070), .B(n9959), .Y(n15599));
  AOI21X1 g12284(.A0(n3070), .A1(DATAI_25_), .B0(n15599), .Y(n15600));
  NOR3X1  g12285(.A(n15600), .B(n15354), .C(n15353), .Y(n15601));
  NOR2X1  g12286(.A(n3070), .B(n9963), .Y(n15602));
  AOI21X1 g12287(.A0(n3070), .A1(DATAI_17_), .B0(n15602), .Y(n15603));
  INVX1   g12288(.A(n15603), .Y(n15604));
  NAND3X1 g12289(.A(n15604), .B(n15346), .C(n15352), .Y(n15605));
  NAND3X1 g12290(.A(n15346), .B(n14770), .C(P1_STATE2_REG_3__SCAN_IN), .Y(n15606));
  OAI22X1 g12291(.A0(n15605), .A1(n15508), .B0(n15491), .B1(n15606), .Y(n15607));
  AOI21X1 g12292(.A0(n15601), .A1(n15485), .B0(n15607), .Y(n15608));
  NAND3X1 g12293(.A(n15608), .B(n15598), .C(n15594), .Y(P1_U3154));
  NAND2X1 g12294(.A(n15496), .B(P1_INSTQUEUE_REG_15__0__SCAN_IN), .Y(n15610));
  NOR2X1  g12295(.A(n3070), .B(n9972), .Y(n15611));
  AOI21X1 g12296(.A0(n3070), .A1(DATAI_0_), .B0(n15611), .Y(n15612));
  NOR2X1  g12297(.A(n15612), .B(n15354), .Y(n15613));
  NAND2X1 g12298(.A(n15613), .B(n15503), .Y(n15614));
  NOR2X1  g12299(.A(n3070), .B(n9978), .Y(n15615));
  AOI21X1 g12300(.A0(n3070), .A1(DATAI_24_), .B0(n15615), .Y(n15616));
  NOR3X1  g12301(.A(n15616), .B(n15354), .C(n15353), .Y(n15617));
  NOR2X1  g12302(.A(n3070), .B(n9982), .Y(n15618));
  AOI21X1 g12303(.A0(n3070), .A1(DATAI_16_), .B0(n15618), .Y(n15619));
  INVX1   g12304(.A(n15619), .Y(n15620));
  NAND3X1 g12305(.A(n15620), .B(n15346), .C(n15352), .Y(n15621));
  NAND3X1 g12306(.A(n15346), .B(n14806), .C(P1_STATE2_REG_3__SCAN_IN), .Y(n15622));
  OAI22X1 g12307(.A0(n15621), .A1(n15508), .B0(n15491), .B1(n15622), .Y(n15623));
  AOI21X1 g12308(.A0(n15617), .A1(n15485), .B0(n15623), .Y(n15624));
  NAND3X1 g12309(.A(n15624), .B(n15614), .C(n15610), .Y(P1_U3153));
  NOR4X1  g12310(.A(n14656), .B(n14659), .C(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .D(n14653), .Y(n15626));
  NOR2X1  g12311(.A(n15169), .B(n15131), .Y(n15627));
  AOI21X1 g12312(.A0(n15627), .A1(n15348), .B0(n15626), .Y(n15628));
  INVX1   g12313(.A(n15434), .Y(n15629));
  NOR4X1  g12314(.A(n15459), .B(n15629), .C(n15407), .D(n15484), .Y(n15630));
  NOR2X1  g12315(.A(n15434), .B(n15408), .Y(n15631));
  NOR4X1  g12316(.A(n15630), .B(n15354), .C(n15353), .D(n15485), .Y(n15634));
  OAI21X1 g12317(.A0(n15634), .A1(n15351), .B0(n15628), .Y(n15635));
  INVX1   g12318(.A(n15626), .Y(n15636));
  INVX1   g12319(.A(n15147), .Y(n15637));
  NAND2X1 g12320(.A(n15492), .B(n15637), .Y(n15638));
  AOI22X1 g12321(.A0(n15636), .A1(P1_STATE2_REG_3__SCAN_IN), .B0(P1_STATE2_REG_2__SCAN_IN), .B1(n15638), .Y(n15639));
  NAND3X1 g12322(.A(n15639), .B(n15635), .C(n15346), .Y(n15640));
  NAND2X1 g12323(.A(n15640), .B(P1_INSTQUEUE_REG_14__7__SCAN_IN), .Y(n15641));
  NOR3X1  g12324(.A(n15485), .B(n15630), .C(n15353), .Y(n15642));
  NOR2X1  g12325(.A(n15642), .B(n15351), .Y(n15643));
  OAI22X1 g12326(.A0(n15638), .A1(n15155), .B0(n15628), .B1(n15643), .Y(n15644));
  NAND2X1 g12327(.A(n15644), .B(n15500), .Y(n15645));
  INVX1   g12328(.A(n15485), .Y(n15646));
  OAI22X1 g12329(.A0(n15636), .A1(n15513), .B0(n15512), .B1(n15646), .Y(n15647));
  AOI21X1 g12330(.A0(n15630), .A1(n15507), .B0(n15647), .Y(n15648));
  NAND3X1 g12331(.A(n15648), .B(n15645), .C(n15641), .Y(P1_U3152));
  NAND2X1 g12332(.A(n15640), .B(P1_INSTQUEUE_REG_14__6__SCAN_IN), .Y(n15650));
  NAND2X1 g12333(.A(n15644), .B(n15520), .Y(n15651));
  NAND2X1 g12334(.A(n15630), .B(n15524), .Y(n15652));
  AOI22X1 g12335(.A0(n15626), .A1(n15529), .B0(n15528), .B1(n15485), .Y(n15653));
  NAND4X1 g12336(.A(n15652), .B(n15651), .C(n15650), .D(n15653), .Y(P1_U3151));
  NAND2X1 g12337(.A(n15640), .B(P1_INSTQUEUE_REG_14__5__SCAN_IN), .Y(n15655));
  NAND2X1 g12338(.A(n15644), .B(n15535), .Y(n15656));
  NAND2X1 g12339(.A(n15630), .B(n15539), .Y(n15657));
  AOI22X1 g12340(.A0(n15626), .A1(n15544), .B0(n15543), .B1(n15485), .Y(n15658));
  NAND4X1 g12341(.A(n15657), .B(n15656), .C(n15655), .D(n15658), .Y(P1_U3150));
  NAND2X1 g12342(.A(n15640), .B(P1_INSTQUEUE_REG_14__4__SCAN_IN), .Y(n15660));
  NAND2X1 g12343(.A(n15644), .B(n15550), .Y(n15661));
  NAND2X1 g12344(.A(n15630), .B(n15554), .Y(n15662));
  AOI22X1 g12345(.A0(n15626), .A1(n15559), .B0(n15558), .B1(n15485), .Y(n15663));
  NAND4X1 g12346(.A(n15662), .B(n15661), .C(n15660), .D(n15663), .Y(P1_U3149));
  NAND2X1 g12347(.A(n15640), .B(P1_INSTQUEUE_REG_14__3__SCAN_IN), .Y(n15665));
  NAND2X1 g12348(.A(n15644), .B(n15565), .Y(n15666));
  OAI22X1 g12349(.A0(n15636), .A1(n15574), .B0(n15573), .B1(n15646), .Y(n15667));
  AOI21X1 g12350(.A0(n15630), .A1(n15569), .B0(n15667), .Y(n15668));
  NAND3X1 g12351(.A(n15668), .B(n15666), .C(n15665), .Y(P1_U3148));
  NAND2X1 g12352(.A(n15640), .B(P1_INSTQUEUE_REG_14__2__SCAN_IN), .Y(n15670));
  NAND2X1 g12353(.A(n15644), .B(n15581), .Y(n15671));
  OAI22X1 g12354(.A0(n15636), .A1(n15590), .B0(n15589), .B1(n15646), .Y(n15672));
  AOI21X1 g12355(.A0(n15630), .A1(n15585), .B0(n15672), .Y(n15673));
  NAND3X1 g12356(.A(n15673), .B(n15671), .C(n15670), .Y(P1_U3147));
  NAND2X1 g12357(.A(n15640), .B(P1_INSTQUEUE_REG_14__1__SCAN_IN), .Y(n15675));
  NAND2X1 g12358(.A(n15644), .B(n15597), .Y(n15676));
  OAI22X1 g12359(.A0(n15636), .A1(n15606), .B0(n15605), .B1(n15646), .Y(n15677));
  AOI21X1 g12360(.A0(n15630), .A1(n15601), .B0(n15677), .Y(n15678));
  NAND3X1 g12361(.A(n15678), .B(n15676), .C(n15675), .Y(P1_U3146));
  NAND2X1 g12362(.A(n15640), .B(P1_INSTQUEUE_REG_14__0__SCAN_IN), .Y(n15680));
  NAND2X1 g12363(.A(n15644), .B(n15613), .Y(n15681));
  OAI22X1 g12364(.A0(n15636), .A1(n15622), .B0(n15621), .B1(n15646), .Y(n15682));
  AOI21X1 g12365(.A0(n15630), .A1(n15617), .B0(n15682), .Y(n15683));
  NAND3X1 g12366(.A(n15683), .B(n15681), .C(n15680), .Y(P1_U3145));
  NOR4X1  g12367(.A(n14656), .B(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C(n14658), .D(n14653), .Y(n15685));
  NOR2X1  g12368(.A(n15168), .B(n15132), .Y(n15686));
  AOI21X1 g12369(.A0(n15686), .A1(n15348), .B0(n15685), .Y(n15687));
  NOR4X1  g12370(.A(n15459), .B(n15629), .C(n15408), .D(n15484), .Y(n15688));
  NOR4X1  g12371(.A(n15688), .B(n15354), .C(n15353), .D(n15630), .Y(n15692));
  OAI21X1 g12372(.A0(n15692), .A1(n15351), .B0(n15687), .Y(n15693));
  INVX1   g12373(.A(n15685), .Y(n15694));
  NOR2X1  g12374(.A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Y(n15695));
  AOI21X1 g12375(.A0(n15695), .A1(n15492), .B0(n15685), .Y(n15696));
  AOI22X1 g12376(.A0(n15694), .A1(P1_STATE2_REG_3__SCAN_IN), .B0(P1_STATE2_REG_2__SCAN_IN), .B1(n15696), .Y(n15697));
  NAND3X1 g12377(.A(n15697), .B(n15693), .C(n15346), .Y(n15698));
  NAND2X1 g12378(.A(n15698), .B(P1_INSTQUEUE_REG_13__7__SCAN_IN), .Y(n15699));
  NOR3X1  g12379(.A(n15630), .B(n15688), .C(n15353), .Y(n15700));
  NOR2X1  g12380(.A(n15700), .B(n15351), .Y(n15701));
  OAI22X1 g12381(.A0(n15696), .A1(n15155), .B0(n15687), .B1(n15701), .Y(n15702));
  NAND2X1 g12382(.A(n15702), .B(n15500), .Y(n15703));
  INVX1   g12383(.A(n15630), .Y(n15704));
  OAI22X1 g12384(.A0(n15694), .A1(n15513), .B0(n15512), .B1(n15704), .Y(n15705));
  AOI21X1 g12385(.A0(n15688), .A1(n15507), .B0(n15705), .Y(n15706));
  NAND3X1 g12386(.A(n15706), .B(n15703), .C(n15699), .Y(P1_U3144));
  NAND2X1 g12387(.A(n15698), .B(P1_INSTQUEUE_REG_13__6__SCAN_IN), .Y(n15708));
  NAND2X1 g12388(.A(n15702), .B(n15520), .Y(n15709));
  NAND2X1 g12389(.A(n15688), .B(n15524), .Y(n15710));
  AOI22X1 g12390(.A0(n15685), .A1(n15529), .B0(n15528), .B1(n15630), .Y(n15711));
  NAND4X1 g12391(.A(n15710), .B(n15709), .C(n15708), .D(n15711), .Y(P1_U3143));
  NAND2X1 g12392(.A(n15698), .B(P1_INSTQUEUE_REG_13__5__SCAN_IN), .Y(n15713));
  NAND2X1 g12393(.A(n15702), .B(n15535), .Y(n15714));
  NAND2X1 g12394(.A(n15688), .B(n15539), .Y(n15715));
  AOI22X1 g12395(.A0(n15685), .A1(n15544), .B0(n15543), .B1(n15630), .Y(n15716));
  NAND4X1 g12396(.A(n15715), .B(n15714), .C(n15713), .D(n15716), .Y(P1_U3142));
  NAND2X1 g12397(.A(n15698), .B(P1_INSTQUEUE_REG_13__4__SCAN_IN), .Y(n15718));
  NAND2X1 g12398(.A(n15702), .B(n15550), .Y(n15719));
  NAND2X1 g12399(.A(n15688), .B(n15554), .Y(n15720));
  AOI22X1 g12400(.A0(n15685), .A1(n15559), .B0(n15558), .B1(n15630), .Y(n15721));
  NAND4X1 g12401(.A(n15720), .B(n15719), .C(n15718), .D(n15721), .Y(P1_U3141));
  NAND2X1 g12402(.A(n15698), .B(P1_INSTQUEUE_REG_13__3__SCAN_IN), .Y(n15723));
  NAND2X1 g12403(.A(n15702), .B(n15565), .Y(n15724));
  OAI22X1 g12404(.A0(n15694), .A1(n15574), .B0(n15573), .B1(n15704), .Y(n15725));
  AOI21X1 g12405(.A0(n15688), .A1(n15569), .B0(n15725), .Y(n15726));
  NAND3X1 g12406(.A(n15726), .B(n15724), .C(n15723), .Y(P1_U3140));
  NAND2X1 g12407(.A(n15698), .B(P1_INSTQUEUE_REG_13__2__SCAN_IN), .Y(n15728));
  NAND2X1 g12408(.A(n15702), .B(n15581), .Y(n15729));
  OAI22X1 g12409(.A0(n15694), .A1(n15590), .B0(n15589), .B1(n15704), .Y(n15730));
  AOI21X1 g12410(.A0(n15688), .A1(n15585), .B0(n15730), .Y(n15731));
  NAND3X1 g12411(.A(n15731), .B(n15729), .C(n15728), .Y(P1_U3139));
  NAND2X1 g12412(.A(n15698), .B(P1_INSTQUEUE_REG_13__1__SCAN_IN), .Y(n15733));
  NAND2X1 g12413(.A(n15702), .B(n15597), .Y(n15734));
  OAI22X1 g12414(.A0(n15694), .A1(n15606), .B0(n15605), .B1(n15704), .Y(n15735));
  AOI21X1 g12415(.A0(n15688), .A1(n15601), .B0(n15735), .Y(n15736));
  NAND3X1 g12416(.A(n15736), .B(n15734), .C(n15733), .Y(P1_U3138));
  NAND2X1 g12417(.A(n15698), .B(P1_INSTQUEUE_REG_13__0__SCAN_IN), .Y(n15738));
  NAND2X1 g12418(.A(n15702), .B(n15613), .Y(n15739));
  OAI22X1 g12419(.A0(n15694), .A1(n15622), .B0(n15621), .B1(n15704), .Y(n15740));
  AOI21X1 g12420(.A0(n15688), .A1(n15617), .B0(n15740), .Y(n15741));
  NAND3X1 g12421(.A(n15741), .B(n15739), .C(n15738), .Y(P1_U3137));
  NOR4X1  g12422(.A(n14656), .B(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .D(n14653), .Y(n15743));
  NOR2X1  g12423(.A(n15168), .B(n15131), .Y(n15744));
  AOI21X1 g12424(.A0(n15744), .A1(n15348), .B0(n15743), .Y(n15745));
  INVX1   g12425(.A(n15459), .Y(n15746));
  NOR4X1  g12426(.A(n15746), .B(n15434), .C(n15407), .D(n15484), .Y(n15747));
  NOR4X1  g12427(.A(n15747), .B(n15354), .C(n15353), .D(n15688), .Y(n15751));
  OAI21X1 g12428(.A0(n15751), .A1(n15351), .B0(n15745), .Y(n15752));
  INVX1   g12429(.A(n15743), .Y(n15753));
  NAND2X1 g12430(.A(n15492), .B(n15147), .Y(n15754));
  AOI22X1 g12431(.A0(n15753), .A1(P1_STATE2_REG_3__SCAN_IN), .B0(P1_STATE2_REG_2__SCAN_IN), .B1(n15754), .Y(n15755));
  NAND3X1 g12432(.A(n15755), .B(n15752), .C(n15346), .Y(n15756));
  NAND2X1 g12433(.A(n15756), .B(P1_INSTQUEUE_REG_12__7__SCAN_IN), .Y(n15757));
  NOR3X1  g12434(.A(n15688), .B(n15747), .C(n15353), .Y(n15758));
  NOR2X1  g12435(.A(n15758), .B(n15351), .Y(n15759));
  OAI22X1 g12436(.A0(n15754), .A1(n15155), .B0(n15745), .B1(n15759), .Y(n15760));
  NAND2X1 g12437(.A(n15760), .B(n15500), .Y(n15761));
  INVX1   g12438(.A(n15688), .Y(n15762));
  OAI22X1 g12439(.A0(n15753), .A1(n15513), .B0(n15512), .B1(n15762), .Y(n15763));
  AOI21X1 g12440(.A0(n15747), .A1(n15507), .B0(n15763), .Y(n15764));
  NAND3X1 g12441(.A(n15764), .B(n15761), .C(n15757), .Y(P1_U3136));
  NAND2X1 g12442(.A(n15756), .B(P1_INSTQUEUE_REG_12__6__SCAN_IN), .Y(n15766));
  NAND2X1 g12443(.A(n15760), .B(n15520), .Y(n15767));
  NAND2X1 g12444(.A(n15747), .B(n15524), .Y(n15768));
  AOI22X1 g12445(.A0(n15743), .A1(n15529), .B0(n15528), .B1(n15688), .Y(n15769));
  NAND4X1 g12446(.A(n15768), .B(n15767), .C(n15766), .D(n15769), .Y(P1_U3135));
  NAND2X1 g12447(.A(n15756), .B(P1_INSTQUEUE_REG_12__5__SCAN_IN), .Y(n15771));
  NAND2X1 g12448(.A(n15760), .B(n15535), .Y(n15772));
  NAND2X1 g12449(.A(n15747), .B(n15539), .Y(n15773));
  AOI22X1 g12450(.A0(n15743), .A1(n15544), .B0(n15543), .B1(n15688), .Y(n15774));
  NAND4X1 g12451(.A(n15773), .B(n15772), .C(n15771), .D(n15774), .Y(P1_U3134));
  NAND2X1 g12452(.A(n15756), .B(P1_INSTQUEUE_REG_12__4__SCAN_IN), .Y(n15776));
  NAND2X1 g12453(.A(n15760), .B(n15550), .Y(n15777));
  NAND2X1 g12454(.A(n15747), .B(n15554), .Y(n15778));
  AOI22X1 g12455(.A0(n15743), .A1(n15559), .B0(n15558), .B1(n15688), .Y(n15779));
  NAND4X1 g12456(.A(n15778), .B(n15777), .C(n15776), .D(n15779), .Y(P1_U3133));
  NAND2X1 g12457(.A(n15756), .B(P1_INSTQUEUE_REG_12__3__SCAN_IN), .Y(n15781));
  NAND2X1 g12458(.A(n15760), .B(n15565), .Y(n15782));
  OAI22X1 g12459(.A0(n15753), .A1(n15574), .B0(n15573), .B1(n15762), .Y(n15783));
  AOI21X1 g12460(.A0(n15747), .A1(n15569), .B0(n15783), .Y(n15784));
  NAND3X1 g12461(.A(n15784), .B(n15782), .C(n15781), .Y(P1_U3132));
  NAND2X1 g12462(.A(n15756), .B(P1_INSTQUEUE_REG_12__2__SCAN_IN), .Y(n15786));
  NAND2X1 g12463(.A(n15760), .B(n15581), .Y(n15787));
  OAI22X1 g12464(.A0(n15753), .A1(n15590), .B0(n15589), .B1(n15762), .Y(n15788));
  AOI21X1 g12465(.A0(n15747), .A1(n15585), .B0(n15788), .Y(n15789));
  NAND3X1 g12466(.A(n15789), .B(n15787), .C(n15786), .Y(P1_U3131));
  NAND2X1 g12467(.A(n15756), .B(P1_INSTQUEUE_REG_12__1__SCAN_IN), .Y(n15791));
  NAND2X1 g12468(.A(n15760), .B(n15597), .Y(n15792));
  OAI22X1 g12469(.A0(n15753), .A1(n15606), .B0(n15605), .B1(n15762), .Y(n15793));
  AOI21X1 g12470(.A0(n15747), .A1(n15601), .B0(n15793), .Y(n15794));
  NAND3X1 g12471(.A(n15794), .B(n15792), .C(n15791), .Y(P1_U3130));
  NAND2X1 g12472(.A(n15756), .B(P1_INSTQUEUE_REG_12__0__SCAN_IN), .Y(n15796));
  NAND2X1 g12473(.A(n15760), .B(n15613), .Y(n15797));
  OAI22X1 g12474(.A0(n15753), .A1(n15622), .B0(n15621), .B1(n15762), .Y(n15798));
  AOI21X1 g12475(.A0(n15747), .A1(n15617), .B0(n15798), .Y(n15799));
  NAND3X1 g12476(.A(n15799), .B(n15797), .C(n15796), .Y(P1_U3129));
  NOR4X1  g12477(.A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n14659), .C(n14658), .D(n14653), .Y(n15801));
  INVX1   g12478(.A(n15192), .Y(n15802));
  NOR2X1  g12479(.A(n15219), .B(n15802), .Y(n15803));
  AOI21X1 g12480(.A0(n15803), .A1(n15349), .B0(n15801), .Y(n15804));
  NOR4X1  g12481(.A(n15746), .B(n15434), .C(n15408), .D(n15484), .Y(n15805));
  NOR4X1  g12482(.A(n15805), .B(n15354), .C(n15353), .D(n15747), .Y(n15807));
  OAI21X1 g12483(.A0(n15807), .A1(n15351), .B0(n15804), .Y(n15808));
  INVX1   g12484(.A(n15801), .Y(n15809));
  INVX1   g12485(.A(n15185), .Y(n15810));
  NOR2X1  g12486(.A(n15215), .B(n15810), .Y(n15811));
  AOI21X1 g12487(.A0(n15811), .A1(n15493), .B0(n15801), .Y(n15812));
  AOI22X1 g12488(.A0(n15809), .A1(P1_STATE2_REG_3__SCAN_IN), .B0(P1_STATE2_REG_2__SCAN_IN), .B1(n15812), .Y(n15813));
  NAND3X1 g12489(.A(n15813), .B(n15808), .C(n15346), .Y(n15814));
  NAND2X1 g12490(.A(n15814), .B(P1_INSTQUEUE_REG_11__7__SCAN_IN), .Y(n15815));
  NOR3X1  g12491(.A(n15747), .B(n15805), .C(n15353), .Y(n15816));
  NOR2X1  g12492(.A(n15816), .B(n15351), .Y(n15817));
  OAI22X1 g12493(.A0(n15812), .A1(n15155), .B0(n15804), .B1(n15817), .Y(n15818));
  NAND2X1 g12494(.A(n15818), .B(n15500), .Y(n15819));
  INVX1   g12495(.A(n15747), .Y(n15820));
  OAI22X1 g12496(.A0(n15809), .A1(n15513), .B0(n15512), .B1(n15820), .Y(n15821));
  AOI21X1 g12497(.A0(n15805), .A1(n15507), .B0(n15821), .Y(n15822));
  NAND3X1 g12498(.A(n15822), .B(n15819), .C(n15815), .Y(P1_U3128));
  NAND2X1 g12499(.A(n15814), .B(P1_INSTQUEUE_REG_11__6__SCAN_IN), .Y(n15824));
  NAND2X1 g12500(.A(n15818), .B(n15520), .Y(n15825));
  NAND2X1 g12501(.A(n15805), .B(n15524), .Y(n15826));
  AOI22X1 g12502(.A0(n15801), .A1(n15529), .B0(n15528), .B1(n15747), .Y(n15827));
  NAND4X1 g12503(.A(n15826), .B(n15825), .C(n15824), .D(n15827), .Y(P1_U3127));
  NAND2X1 g12504(.A(n15814), .B(P1_INSTQUEUE_REG_11__5__SCAN_IN), .Y(n15829));
  NAND2X1 g12505(.A(n15818), .B(n15535), .Y(n15830));
  NAND2X1 g12506(.A(n15805), .B(n15539), .Y(n15831));
  AOI22X1 g12507(.A0(n15801), .A1(n15544), .B0(n15543), .B1(n15747), .Y(n15832));
  NAND4X1 g12508(.A(n15831), .B(n15830), .C(n15829), .D(n15832), .Y(P1_U3126));
  NAND2X1 g12509(.A(n15814), .B(P1_INSTQUEUE_REG_11__4__SCAN_IN), .Y(n15834));
  NAND2X1 g12510(.A(n15818), .B(n15550), .Y(n15835));
  NAND2X1 g12511(.A(n15805), .B(n15554), .Y(n15836));
  AOI22X1 g12512(.A0(n15801), .A1(n15559), .B0(n15558), .B1(n15747), .Y(n15837));
  NAND4X1 g12513(.A(n15836), .B(n15835), .C(n15834), .D(n15837), .Y(P1_U3125));
  NAND2X1 g12514(.A(n15814), .B(P1_INSTQUEUE_REG_11__3__SCAN_IN), .Y(n15839));
  NAND2X1 g12515(.A(n15818), .B(n15565), .Y(n15840));
  OAI22X1 g12516(.A0(n15809), .A1(n15574), .B0(n15573), .B1(n15820), .Y(n15841));
  AOI21X1 g12517(.A0(n15805), .A1(n15569), .B0(n15841), .Y(n15842));
  NAND3X1 g12518(.A(n15842), .B(n15840), .C(n15839), .Y(P1_U3124));
  NAND2X1 g12519(.A(n15814), .B(P1_INSTQUEUE_REG_11__2__SCAN_IN), .Y(n15844));
  NAND2X1 g12520(.A(n15818), .B(n15581), .Y(n15845));
  OAI22X1 g12521(.A0(n15809), .A1(n15590), .B0(n15589), .B1(n15820), .Y(n15846));
  AOI21X1 g12522(.A0(n15805), .A1(n15585), .B0(n15846), .Y(n15847));
  NAND3X1 g12523(.A(n15847), .B(n15845), .C(n15844), .Y(P1_U3123));
  NAND2X1 g12524(.A(n15814), .B(P1_INSTQUEUE_REG_11__1__SCAN_IN), .Y(n15849));
  NAND2X1 g12525(.A(n15818), .B(n15597), .Y(n15850));
  OAI22X1 g12526(.A0(n15809), .A1(n15606), .B0(n15605), .B1(n15820), .Y(n15851));
  AOI21X1 g12527(.A0(n15805), .A1(n15601), .B0(n15851), .Y(n15852));
  NAND3X1 g12528(.A(n15852), .B(n15850), .C(n15849), .Y(P1_U3122));
  NAND2X1 g12529(.A(n15814), .B(P1_INSTQUEUE_REG_11__0__SCAN_IN), .Y(n15854));
  NAND2X1 g12530(.A(n15818), .B(n15613), .Y(n15855));
  OAI22X1 g12531(.A0(n15809), .A1(n15622), .B0(n15621), .B1(n15820), .Y(n15856));
  AOI21X1 g12532(.A0(n15805), .A1(n15617), .B0(n15856), .Y(n15857));
  NAND3X1 g12533(.A(n15857), .B(n15855), .C(n15854), .Y(P1_U3121));
  NOR4X1  g12534(.A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n14659), .C(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .D(n14653), .Y(n15859));
  AOI21X1 g12535(.A0(n15803), .A1(n15627), .B0(n15859), .Y(n15860));
  NOR4X1  g12536(.A(n15746), .B(n15629), .C(n15407), .D(n15484), .Y(n15861));
  NOR4X1  g12537(.A(n15861), .B(n15354), .C(n15353), .D(n15805), .Y(n15863));
  OAI21X1 g12538(.A0(n15863), .A1(n15351), .B0(n15860), .Y(n15864));
  INVX1   g12539(.A(n15859), .Y(n15865));
  INVX1   g12540(.A(n15215), .Y(n15866));
  NAND3X1 g12541(.A(n15866), .B(n15185), .C(n15637), .Y(n15867));
  AOI22X1 g12542(.A0(n15865), .A1(P1_STATE2_REG_3__SCAN_IN), .B0(P1_STATE2_REG_2__SCAN_IN), .B1(n15867), .Y(n15868));
  NAND3X1 g12543(.A(n15868), .B(n15864), .C(n15346), .Y(n15869));
  NAND2X1 g12544(.A(n15869), .B(P1_INSTQUEUE_REG_10__7__SCAN_IN), .Y(n15870));
  NOR3X1  g12545(.A(n15805), .B(n15861), .C(n15353), .Y(n15871));
  NOR2X1  g12546(.A(n15871), .B(n15351), .Y(n15872));
  OAI22X1 g12547(.A0(n15867), .A1(n15155), .B0(n15860), .B1(n15872), .Y(n15873));
  NAND2X1 g12548(.A(n15873), .B(n15500), .Y(n15874));
  INVX1   g12549(.A(n15805), .Y(n15875));
  OAI22X1 g12550(.A0(n15865), .A1(n15513), .B0(n15512), .B1(n15875), .Y(n15876));
  AOI21X1 g12551(.A0(n15861), .A1(n15507), .B0(n15876), .Y(n15877));
  NAND3X1 g12552(.A(n15877), .B(n15874), .C(n15870), .Y(P1_U3120));
  NAND2X1 g12553(.A(n15869), .B(P1_INSTQUEUE_REG_10__6__SCAN_IN), .Y(n15879));
  NAND2X1 g12554(.A(n15873), .B(n15520), .Y(n15880));
  NAND2X1 g12555(.A(n15861), .B(n15524), .Y(n15881));
  AOI22X1 g12556(.A0(n15859), .A1(n15529), .B0(n15528), .B1(n15805), .Y(n15882));
  NAND4X1 g12557(.A(n15881), .B(n15880), .C(n15879), .D(n15882), .Y(P1_U3119));
  NAND2X1 g12558(.A(n15869), .B(P1_INSTQUEUE_REG_10__5__SCAN_IN), .Y(n15884));
  NAND2X1 g12559(.A(n15873), .B(n15535), .Y(n15885));
  NAND2X1 g12560(.A(n15861), .B(n15539), .Y(n15886));
  AOI22X1 g12561(.A0(n15859), .A1(n15544), .B0(n15543), .B1(n15805), .Y(n15887));
  NAND4X1 g12562(.A(n15886), .B(n15885), .C(n15884), .D(n15887), .Y(P1_U3118));
  NAND2X1 g12563(.A(n15869), .B(P1_INSTQUEUE_REG_10__4__SCAN_IN), .Y(n15889));
  NAND2X1 g12564(.A(n15873), .B(n15550), .Y(n15890));
  NAND2X1 g12565(.A(n15861), .B(n15554), .Y(n15891));
  AOI22X1 g12566(.A0(n15859), .A1(n15559), .B0(n15558), .B1(n15805), .Y(n15892));
  NAND4X1 g12567(.A(n15891), .B(n15890), .C(n15889), .D(n15892), .Y(P1_U3117));
  NAND2X1 g12568(.A(n15869), .B(P1_INSTQUEUE_REG_10__3__SCAN_IN), .Y(n15894));
  NAND2X1 g12569(.A(n15873), .B(n15565), .Y(n15895));
  OAI22X1 g12570(.A0(n15865), .A1(n15574), .B0(n15573), .B1(n15875), .Y(n15896));
  AOI21X1 g12571(.A0(n15861), .A1(n15569), .B0(n15896), .Y(n15897));
  NAND3X1 g12572(.A(n15897), .B(n15895), .C(n15894), .Y(P1_U3116));
  NAND2X1 g12573(.A(n15869), .B(P1_INSTQUEUE_REG_10__2__SCAN_IN), .Y(n15899));
  NAND2X1 g12574(.A(n15873), .B(n15581), .Y(n15900));
  OAI22X1 g12575(.A0(n15865), .A1(n15590), .B0(n15589), .B1(n15875), .Y(n15901));
  AOI21X1 g12576(.A0(n15861), .A1(n15585), .B0(n15901), .Y(n15902));
  NAND3X1 g12577(.A(n15902), .B(n15900), .C(n15899), .Y(P1_U3115));
  NAND2X1 g12578(.A(n15869), .B(P1_INSTQUEUE_REG_10__1__SCAN_IN), .Y(n15904));
  NAND2X1 g12579(.A(n15873), .B(n15597), .Y(n15905));
  OAI22X1 g12580(.A0(n15865), .A1(n15606), .B0(n15605), .B1(n15875), .Y(n15906));
  AOI21X1 g12581(.A0(n15861), .A1(n15601), .B0(n15906), .Y(n15907));
  NAND3X1 g12582(.A(n15907), .B(n15905), .C(n15904), .Y(P1_U3114));
  NAND2X1 g12583(.A(n15869), .B(P1_INSTQUEUE_REG_10__0__SCAN_IN), .Y(n15909));
  NAND2X1 g12584(.A(n15873), .B(n15613), .Y(n15910));
  OAI22X1 g12585(.A0(n15865), .A1(n15622), .B0(n15621), .B1(n15875), .Y(n15911));
  AOI21X1 g12586(.A0(n15861), .A1(n15617), .B0(n15911), .Y(n15912));
  NAND3X1 g12587(.A(n15912), .B(n15910), .C(n15909), .Y(P1_U3113));
  NOR4X1  g12588(.A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C(n14658), .D(n14653), .Y(n15914));
  AOI21X1 g12589(.A0(n15803), .A1(n15686), .B0(n15914), .Y(n15915));
  NOR4X1  g12590(.A(n15746), .B(n15629), .C(n15408), .D(n15484), .Y(n15916));
  NOR4X1  g12591(.A(n15916), .B(n15354), .C(n15353), .D(n15861), .Y(n15918));
  OAI21X1 g12592(.A0(n15918), .A1(n15351), .B0(n15915), .Y(n15919));
  INVX1   g12593(.A(n15914), .Y(n15920));
  AOI21X1 g12594(.A0(n15811), .A1(n15695), .B0(n15914), .Y(n15921));
  AOI22X1 g12595(.A0(n15920), .A1(P1_STATE2_REG_3__SCAN_IN), .B0(P1_STATE2_REG_2__SCAN_IN), .B1(n15921), .Y(n15922));
  NAND3X1 g12596(.A(n15922), .B(n15919), .C(n15346), .Y(n15923));
  NAND2X1 g12597(.A(n15923), .B(P1_INSTQUEUE_REG_9__7__SCAN_IN), .Y(n15924));
  NOR3X1  g12598(.A(n15861), .B(n15916), .C(n15353), .Y(n15925));
  NOR2X1  g12599(.A(n15925), .B(n15351), .Y(n15926));
  OAI22X1 g12600(.A0(n15921), .A1(n15155), .B0(n15915), .B1(n15926), .Y(n15927));
  NAND2X1 g12601(.A(n15927), .B(n15500), .Y(n15928));
  INVX1   g12602(.A(n15861), .Y(n15929));
  OAI22X1 g12603(.A0(n15920), .A1(n15513), .B0(n15512), .B1(n15929), .Y(n15930));
  AOI21X1 g12604(.A0(n15916), .A1(n15507), .B0(n15930), .Y(n15931));
  NAND3X1 g12605(.A(n15931), .B(n15928), .C(n15924), .Y(P1_U3112));
  NAND2X1 g12606(.A(n15923), .B(P1_INSTQUEUE_REG_9__6__SCAN_IN), .Y(n15933));
  NAND2X1 g12607(.A(n15927), .B(n15520), .Y(n15934));
  NAND2X1 g12608(.A(n15916), .B(n15524), .Y(n15935));
  AOI22X1 g12609(.A0(n15914), .A1(n15529), .B0(n15528), .B1(n15861), .Y(n15936));
  NAND4X1 g12610(.A(n15935), .B(n15934), .C(n15933), .D(n15936), .Y(P1_U3111));
  NAND2X1 g12611(.A(n15923), .B(P1_INSTQUEUE_REG_9__5__SCAN_IN), .Y(n15938));
  NAND2X1 g12612(.A(n15927), .B(n15535), .Y(n15939));
  NAND2X1 g12613(.A(n15916), .B(n15539), .Y(n15940));
  AOI22X1 g12614(.A0(n15914), .A1(n15544), .B0(n15543), .B1(n15861), .Y(n15941));
  NAND4X1 g12615(.A(n15940), .B(n15939), .C(n15938), .D(n15941), .Y(P1_U3110));
  NAND2X1 g12616(.A(n15923), .B(P1_INSTQUEUE_REG_9__4__SCAN_IN), .Y(n15943));
  NAND2X1 g12617(.A(n15927), .B(n15550), .Y(n15944));
  NAND2X1 g12618(.A(n15916), .B(n15554), .Y(n15945));
  AOI22X1 g12619(.A0(n15914), .A1(n15559), .B0(n15558), .B1(n15861), .Y(n15946));
  NAND4X1 g12620(.A(n15945), .B(n15944), .C(n15943), .D(n15946), .Y(P1_U3109));
  NAND2X1 g12621(.A(n15923), .B(P1_INSTQUEUE_REG_9__3__SCAN_IN), .Y(n15948));
  NAND2X1 g12622(.A(n15927), .B(n15565), .Y(n15949));
  OAI22X1 g12623(.A0(n15920), .A1(n15574), .B0(n15573), .B1(n15929), .Y(n15950));
  AOI21X1 g12624(.A0(n15916), .A1(n15569), .B0(n15950), .Y(n15951));
  NAND3X1 g12625(.A(n15951), .B(n15949), .C(n15948), .Y(P1_U3108));
  NAND2X1 g12626(.A(n15923), .B(P1_INSTQUEUE_REG_9__2__SCAN_IN), .Y(n15953));
  NAND2X1 g12627(.A(n15927), .B(n15581), .Y(n15954));
  OAI22X1 g12628(.A0(n15920), .A1(n15590), .B0(n15589), .B1(n15929), .Y(n15955));
  AOI21X1 g12629(.A0(n15916), .A1(n15585), .B0(n15955), .Y(n15956));
  NAND3X1 g12630(.A(n15956), .B(n15954), .C(n15953), .Y(P1_U3107));
  NAND2X1 g12631(.A(n15923), .B(P1_INSTQUEUE_REG_9__1__SCAN_IN), .Y(n15958));
  NAND2X1 g12632(.A(n15927), .B(n15597), .Y(n15959));
  OAI22X1 g12633(.A0(n15920), .A1(n15606), .B0(n15605), .B1(n15929), .Y(n15960));
  AOI21X1 g12634(.A0(n15916), .A1(n15601), .B0(n15960), .Y(n15961));
  NAND3X1 g12635(.A(n15961), .B(n15959), .C(n15958), .Y(P1_U3106));
  NAND2X1 g12636(.A(n15923), .B(P1_INSTQUEUE_REG_9__0__SCAN_IN), .Y(n15963));
  NAND2X1 g12637(.A(n15927), .B(n15613), .Y(n15964));
  OAI22X1 g12638(.A0(n15920), .A1(n15622), .B0(n15621), .B1(n15929), .Y(n15965));
  AOI21X1 g12639(.A0(n15916), .A1(n15617), .B0(n15965), .Y(n15966));
  NAND3X1 g12640(.A(n15966), .B(n15964), .C(n15963), .Y(P1_U3105));
  NOR4X1  g12641(.A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .D(n14653), .Y(n15968));
  AOI21X1 g12642(.A0(n15803), .A1(n15744), .B0(n15968), .Y(n15969));
  NOR4X1  g12643(.A(n15459), .B(n15434), .C(n15407), .D(n15483), .Y(n15970));
  NOR4X1  g12644(.A(n15970), .B(n15354), .C(n15353), .D(n15916), .Y(n15972));
  OAI21X1 g12645(.A0(n15972), .A1(n15351), .B0(n15969), .Y(n15973));
  INVX1   g12646(.A(n15968), .Y(n15974));
  NAND3X1 g12647(.A(n15866), .B(n15185), .C(n15147), .Y(n15975));
  AOI22X1 g12648(.A0(n15974), .A1(P1_STATE2_REG_3__SCAN_IN), .B0(P1_STATE2_REG_2__SCAN_IN), .B1(n15975), .Y(n15976));
  NAND3X1 g12649(.A(n15976), .B(n15973), .C(n15346), .Y(n15977));
  NAND2X1 g12650(.A(n15977), .B(P1_INSTQUEUE_REG_8__7__SCAN_IN), .Y(n15978));
  NOR3X1  g12651(.A(n15916), .B(n15970), .C(n15353), .Y(n15979));
  NOR2X1  g12652(.A(n15979), .B(n15351), .Y(n15980));
  OAI22X1 g12653(.A0(n15975), .A1(n15155), .B0(n15969), .B1(n15980), .Y(n15981));
  NAND2X1 g12654(.A(n15981), .B(n15500), .Y(n15982));
  INVX1   g12655(.A(n15916), .Y(n15983));
  OAI22X1 g12656(.A0(n15974), .A1(n15513), .B0(n15512), .B1(n15983), .Y(n15984));
  AOI21X1 g12657(.A0(n15970), .A1(n15507), .B0(n15984), .Y(n15985));
  NAND3X1 g12658(.A(n15985), .B(n15982), .C(n15978), .Y(P1_U3104));
  NAND2X1 g12659(.A(n15977), .B(P1_INSTQUEUE_REG_8__6__SCAN_IN), .Y(n15987));
  NAND2X1 g12660(.A(n15981), .B(n15520), .Y(n15988));
  NAND2X1 g12661(.A(n15970), .B(n15524), .Y(n15989));
  AOI22X1 g12662(.A0(n15968), .A1(n15529), .B0(n15528), .B1(n15916), .Y(n15990));
  NAND4X1 g12663(.A(n15989), .B(n15988), .C(n15987), .D(n15990), .Y(P1_U3103));
  NAND2X1 g12664(.A(n15977), .B(P1_INSTQUEUE_REG_8__5__SCAN_IN), .Y(n15992));
  NAND2X1 g12665(.A(n15981), .B(n15535), .Y(n15993));
  NAND2X1 g12666(.A(n15970), .B(n15539), .Y(n15994));
  AOI22X1 g12667(.A0(n15968), .A1(n15544), .B0(n15543), .B1(n15916), .Y(n15995));
  NAND4X1 g12668(.A(n15994), .B(n15993), .C(n15992), .D(n15995), .Y(P1_U3102));
  NAND2X1 g12669(.A(n15977), .B(P1_INSTQUEUE_REG_8__4__SCAN_IN), .Y(n15997));
  NAND2X1 g12670(.A(n15981), .B(n15550), .Y(n15998));
  NAND2X1 g12671(.A(n15970), .B(n15554), .Y(n15999));
  AOI22X1 g12672(.A0(n15968), .A1(n15559), .B0(n15558), .B1(n15916), .Y(n16000));
  NAND4X1 g12673(.A(n15999), .B(n15998), .C(n15997), .D(n16000), .Y(P1_U3101));
  NAND2X1 g12674(.A(n15977), .B(P1_INSTQUEUE_REG_8__3__SCAN_IN), .Y(n16002));
  NAND2X1 g12675(.A(n15981), .B(n15565), .Y(n16003));
  OAI22X1 g12676(.A0(n15974), .A1(n15574), .B0(n15573), .B1(n15983), .Y(n16004));
  AOI21X1 g12677(.A0(n15970), .A1(n15569), .B0(n16004), .Y(n16005));
  NAND3X1 g12678(.A(n16005), .B(n16003), .C(n16002), .Y(P1_U3100));
  NAND2X1 g12679(.A(n15977), .B(P1_INSTQUEUE_REG_8__2__SCAN_IN), .Y(n16007));
  NAND2X1 g12680(.A(n15981), .B(n15581), .Y(n16008));
  OAI22X1 g12681(.A0(n15974), .A1(n15590), .B0(n15589), .B1(n15983), .Y(n16009));
  AOI21X1 g12682(.A0(n15970), .A1(n15585), .B0(n16009), .Y(n16010));
  NAND3X1 g12683(.A(n16010), .B(n16008), .C(n16007), .Y(P1_U3099));
  NAND2X1 g12684(.A(n15977), .B(P1_INSTQUEUE_REG_8__1__SCAN_IN), .Y(n16012));
  NAND2X1 g12685(.A(n15981), .B(n15597), .Y(n16013));
  OAI22X1 g12686(.A0(n15974), .A1(n15606), .B0(n15605), .B1(n15983), .Y(n16014));
  AOI21X1 g12687(.A0(n15970), .A1(n15601), .B0(n16014), .Y(n16015));
  NAND3X1 g12688(.A(n16015), .B(n16013), .C(n16012), .Y(P1_U3098));
  NAND2X1 g12689(.A(n15977), .B(P1_INSTQUEUE_REG_8__0__SCAN_IN), .Y(n16017));
  NAND2X1 g12690(.A(n15981), .B(n15613), .Y(n16018));
  OAI22X1 g12691(.A0(n15974), .A1(n15622), .B0(n15621), .B1(n15983), .Y(n16019));
  AOI21X1 g12692(.A0(n15970), .A1(n15617), .B0(n16019), .Y(n16020));
  NAND3X1 g12693(.A(n16020), .B(n16018), .C(n16017), .Y(P1_U3097));
  NOR2X1  g12694(.A(n15218), .B(n15192), .Y(n16022));
  AOI21X1 g12695(.A0(n16022), .A1(n15349), .B0(n15213), .Y(n16023));
  NOR4X1  g12696(.A(n15459), .B(n15434), .C(n15408), .D(n15483), .Y(n16025));
  NOR4X1  g12697(.A(n15970), .B(n15354), .C(n15353), .D(n16025), .Y(n16026));
  OAI21X1 g12698(.A0(n16026), .A1(n15351), .B0(n16023), .Y(n16027));
  INVX1   g12699(.A(n15213), .Y(n16028));
  NOR4X1  g12700(.A(n15213), .B(n15212), .C(n15185), .D(n15214), .Y(n16029));
  AOI21X1 g12701(.A0(n16029), .A1(n15493), .B0(n15213), .Y(n16030));
  AOI22X1 g12702(.A0(n16028), .A1(P1_STATE2_REG_3__SCAN_IN), .B0(P1_STATE2_REG_2__SCAN_IN), .B1(n16030), .Y(n16031));
  NAND3X1 g12703(.A(n16031), .B(n16027), .C(n15346), .Y(n16032));
  NAND2X1 g12704(.A(n16032), .B(P1_INSTQUEUE_REG_7__7__SCAN_IN), .Y(n16033));
  NOR3X1  g12705(.A(n16025), .B(n15970), .C(n15353), .Y(n16034));
  NOR2X1  g12706(.A(n16034), .B(n15351), .Y(n16035));
  OAI22X1 g12707(.A0(n16030), .A1(n15155), .B0(n16023), .B1(n16035), .Y(n16036));
  NAND2X1 g12708(.A(n16036), .B(n15500), .Y(n16037));
  INVX1   g12709(.A(n15970), .Y(n16038));
  OAI22X1 g12710(.A0(n15512), .A1(n16038), .B0(n16028), .B1(n15513), .Y(n16039));
  AOI21X1 g12711(.A0(n16025), .A1(n15507), .B0(n16039), .Y(n16040));
  NAND3X1 g12712(.A(n16040), .B(n16037), .C(n16033), .Y(P1_U3096));
  NAND2X1 g12713(.A(n16032), .B(P1_INSTQUEUE_REG_7__6__SCAN_IN), .Y(n16042));
  NAND2X1 g12714(.A(n16036), .B(n15520), .Y(n16043));
  NAND2X1 g12715(.A(n16025), .B(n15524), .Y(n16044));
  AOI22X1 g12716(.A0(n15528), .A1(n15970), .B0(n15213), .B1(n15529), .Y(n16045));
  NAND4X1 g12717(.A(n16044), .B(n16043), .C(n16042), .D(n16045), .Y(P1_U3095));
  NAND2X1 g12718(.A(n16032), .B(P1_INSTQUEUE_REG_7__5__SCAN_IN), .Y(n16047));
  NAND2X1 g12719(.A(n16036), .B(n15535), .Y(n16048));
  NAND2X1 g12720(.A(n16025), .B(n15539), .Y(n16049));
  AOI22X1 g12721(.A0(n15543), .A1(n15970), .B0(n15213), .B1(n15544), .Y(n16050));
  NAND4X1 g12722(.A(n16049), .B(n16048), .C(n16047), .D(n16050), .Y(P1_U3094));
  NAND2X1 g12723(.A(n16032), .B(P1_INSTQUEUE_REG_7__4__SCAN_IN), .Y(n16052));
  NAND2X1 g12724(.A(n16036), .B(n15550), .Y(n16053));
  NAND2X1 g12725(.A(n16025), .B(n15554), .Y(n16054));
  AOI22X1 g12726(.A0(n15558), .A1(n15970), .B0(n15213), .B1(n15559), .Y(n16055));
  NAND4X1 g12727(.A(n16054), .B(n16053), .C(n16052), .D(n16055), .Y(P1_U3093));
  NAND2X1 g12728(.A(n16032), .B(P1_INSTQUEUE_REG_7__3__SCAN_IN), .Y(n16057));
  NAND2X1 g12729(.A(n16036), .B(n15565), .Y(n16058));
  OAI22X1 g12730(.A0(n15573), .A1(n16038), .B0(n16028), .B1(n15574), .Y(n16059));
  AOI21X1 g12731(.A0(n16025), .A1(n15569), .B0(n16059), .Y(n16060));
  NAND3X1 g12732(.A(n16060), .B(n16058), .C(n16057), .Y(P1_U3092));
  NAND2X1 g12733(.A(n16032), .B(P1_INSTQUEUE_REG_7__2__SCAN_IN), .Y(n16062));
  NAND2X1 g12734(.A(n16036), .B(n15581), .Y(n16063));
  OAI22X1 g12735(.A0(n15589), .A1(n16038), .B0(n16028), .B1(n15590), .Y(n16064));
  AOI21X1 g12736(.A0(n16025), .A1(n15585), .B0(n16064), .Y(n16065));
  NAND3X1 g12737(.A(n16065), .B(n16063), .C(n16062), .Y(P1_U3091));
  NAND2X1 g12738(.A(n16032), .B(P1_INSTQUEUE_REG_7__1__SCAN_IN), .Y(n16067));
  NAND2X1 g12739(.A(n16036), .B(n15597), .Y(n16068));
  OAI22X1 g12740(.A0(n15605), .A1(n16038), .B0(n16028), .B1(n15606), .Y(n16069));
  AOI21X1 g12741(.A0(n16025), .A1(n15601), .B0(n16069), .Y(n16070));
  NAND3X1 g12742(.A(n16070), .B(n16068), .C(n16067), .Y(P1_U3090));
  NAND2X1 g12743(.A(n16032), .B(P1_INSTQUEUE_REG_7__0__SCAN_IN), .Y(n16072));
  NAND2X1 g12744(.A(n16036), .B(n15613), .Y(n16073));
  OAI22X1 g12745(.A0(n15621), .A1(n16038), .B0(n16028), .B1(n15622), .Y(n16074));
  AOI21X1 g12746(.A0(n16025), .A1(n15617), .B0(n16074), .Y(n16075));
  NAND3X1 g12747(.A(n16075), .B(n16073), .C(n16072), .Y(P1_U3089));
  NOR4X1  g12748(.A(n14656), .B(n14659), .C(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .D(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .Y(n16077));
  AOI21X1 g12749(.A0(n16022), .A1(n15627), .B0(n16077), .Y(n16078));
  NOR4X1  g12750(.A(n15459), .B(n15629), .C(n15407), .D(n15483), .Y(n16079));
  NOR4X1  g12751(.A(n16079), .B(n15354), .C(n15353), .D(n16025), .Y(n16081));
  OAI21X1 g12752(.A0(n16081), .A1(n15351), .B0(n16078), .Y(n16082));
  INVX1   g12753(.A(n16077), .Y(n16083));
  NAND2X1 g12754(.A(n16029), .B(n15637), .Y(n16084));
  AOI22X1 g12755(.A0(n16083), .A1(P1_STATE2_REG_3__SCAN_IN), .B0(P1_STATE2_REG_2__SCAN_IN), .B1(n16084), .Y(n16085));
  NAND3X1 g12756(.A(n16085), .B(n16082), .C(n15346), .Y(n16086));
  NAND2X1 g12757(.A(n16086), .B(P1_INSTQUEUE_REG_6__7__SCAN_IN), .Y(n16087));
  NOR3X1  g12758(.A(n16025), .B(n16079), .C(n15353), .Y(n16088));
  NOR2X1  g12759(.A(n16088), .B(n15351), .Y(n16089));
  OAI22X1 g12760(.A0(n16084), .A1(n15155), .B0(n16078), .B1(n16089), .Y(n16090));
  NAND2X1 g12761(.A(n16090), .B(n15500), .Y(n16091));
  INVX1   g12762(.A(n16025), .Y(n16092));
  OAI22X1 g12763(.A0(n16083), .A1(n15513), .B0(n15512), .B1(n16092), .Y(n16093));
  AOI21X1 g12764(.A0(n16079), .A1(n15507), .B0(n16093), .Y(n16094));
  NAND3X1 g12765(.A(n16094), .B(n16091), .C(n16087), .Y(P1_U3088));
  NAND2X1 g12766(.A(n16086), .B(P1_INSTQUEUE_REG_6__6__SCAN_IN), .Y(n16096));
  NAND2X1 g12767(.A(n16090), .B(n15520), .Y(n16097));
  NAND2X1 g12768(.A(n16079), .B(n15524), .Y(n16098));
  AOI22X1 g12769(.A0(n16077), .A1(n15529), .B0(n15528), .B1(n16025), .Y(n16099));
  NAND4X1 g12770(.A(n16098), .B(n16097), .C(n16096), .D(n16099), .Y(P1_U3087));
  NAND2X1 g12771(.A(n16086), .B(P1_INSTQUEUE_REG_6__5__SCAN_IN), .Y(n16101));
  NAND2X1 g12772(.A(n16090), .B(n15535), .Y(n16102));
  NAND2X1 g12773(.A(n16079), .B(n15539), .Y(n16103));
  AOI22X1 g12774(.A0(n16077), .A1(n15544), .B0(n15543), .B1(n16025), .Y(n16104));
  NAND4X1 g12775(.A(n16103), .B(n16102), .C(n16101), .D(n16104), .Y(P1_U3086));
  NAND2X1 g12776(.A(n16086), .B(P1_INSTQUEUE_REG_6__4__SCAN_IN), .Y(n16106));
  NAND2X1 g12777(.A(n16090), .B(n15550), .Y(n16107));
  NAND2X1 g12778(.A(n16079), .B(n15554), .Y(n16108));
  AOI22X1 g12779(.A0(n16077), .A1(n15559), .B0(n15558), .B1(n16025), .Y(n16109));
  NAND4X1 g12780(.A(n16108), .B(n16107), .C(n16106), .D(n16109), .Y(P1_U3085));
  NAND2X1 g12781(.A(n16086), .B(P1_INSTQUEUE_REG_6__3__SCAN_IN), .Y(n16111));
  NAND2X1 g12782(.A(n16090), .B(n15565), .Y(n16112));
  OAI22X1 g12783(.A0(n16083), .A1(n15574), .B0(n15573), .B1(n16092), .Y(n16113));
  AOI21X1 g12784(.A0(n16079), .A1(n15569), .B0(n16113), .Y(n16114));
  NAND3X1 g12785(.A(n16114), .B(n16112), .C(n16111), .Y(P1_U3084));
  NAND2X1 g12786(.A(n16086), .B(P1_INSTQUEUE_REG_6__2__SCAN_IN), .Y(n16116));
  NAND2X1 g12787(.A(n16090), .B(n15581), .Y(n16117));
  OAI22X1 g12788(.A0(n16083), .A1(n15590), .B0(n15589), .B1(n16092), .Y(n16118));
  AOI21X1 g12789(.A0(n16079), .A1(n15585), .B0(n16118), .Y(n16119));
  NAND3X1 g12790(.A(n16119), .B(n16117), .C(n16116), .Y(P1_U3083));
  NAND2X1 g12791(.A(n16086), .B(P1_INSTQUEUE_REG_6__1__SCAN_IN), .Y(n16121));
  NAND2X1 g12792(.A(n16090), .B(n15597), .Y(n16122));
  OAI22X1 g12793(.A0(n16083), .A1(n15606), .B0(n15605), .B1(n16092), .Y(n16123));
  AOI21X1 g12794(.A0(n16079), .A1(n15601), .B0(n16123), .Y(n16124));
  NAND3X1 g12795(.A(n16124), .B(n16122), .C(n16121), .Y(P1_U3082));
  NAND2X1 g12796(.A(n16086), .B(P1_INSTQUEUE_REG_6__0__SCAN_IN), .Y(n16126));
  NAND2X1 g12797(.A(n16090), .B(n15613), .Y(n16127));
  OAI22X1 g12798(.A0(n16083), .A1(n15622), .B0(n15621), .B1(n16092), .Y(n16128));
  AOI21X1 g12799(.A0(n16079), .A1(n15617), .B0(n16128), .Y(n16129));
  NAND3X1 g12800(.A(n16129), .B(n16127), .C(n16126), .Y(P1_U3081));
  NOR4X1  g12801(.A(n14656), .B(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C(n14658), .D(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .Y(n16131));
  AOI21X1 g12802(.A0(n16022), .A1(n15686), .B0(n16131), .Y(n16132));
  NOR4X1  g12803(.A(n15459), .B(n15629), .C(n15408), .D(n15483), .Y(n16133));
  NOR4X1  g12804(.A(n16133), .B(n15354), .C(n15353), .D(n16079), .Y(n16135));
  OAI21X1 g12805(.A0(n16135), .A1(n15351), .B0(n16132), .Y(n16136));
  INVX1   g12806(.A(n16131), .Y(n16137));
  AOI21X1 g12807(.A0(n16029), .A1(n15695), .B0(n16131), .Y(n16138));
  AOI22X1 g12808(.A0(n16137), .A1(P1_STATE2_REG_3__SCAN_IN), .B0(P1_STATE2_REG_2__SCAN_IN), .B1(n16138), .Y(n16139));
  NAND3X1 g12809(.A(n16139), .B(n16136), .C(n15346), .Y(n16140));
  NAND2X1 g12810(.A(n16140), .B(P1_INSTQUEUE_REG_5__7__SCAN_IN), .Y(n16141));
  NOR3X1  g12811(.A(n16079), .B(n16133), .C(n15353), .Y(n16142));
  NOR2X1  g12812(.A(n16142), .B(n15351), .Y(n16143));
  OAI22X1 g12813(.A0(n16138), .A1(n15155), .B0(n16132), .B1(n16143), .Y(n16144));
  NAND2X1 g12814(.A(n16144), .B(n15500), .Y(n16145));
  INVX1   g12815(.A(n16079), .Y(n16146));
  OAI22X1 g12816(.A0(n16137), .A1(n15513), .B0(n15512), .B1(n16146), .Y(n16147));
  AOI21X1 g12817(.A0(n16133), .A1(n15507), .B0(n16147), .Y(n16148));
  NAND3X1 g12818(.A(n16148), .B(n16145), .C(n16141), .Y(P1_U3080));
  NAND2X1 g12819(.A(n16140), .B(P1_INSTQUEUE_REG_5__6__SCAN_IN), .Y(n16150));
  NAND2X1 g12820(.A(n16144), .B(n15520), .Y(n16151));
  NAND2X1 g12821(.A(n16133), .B(n15524), .Y(n16152));
  AOI22X1 g12822(.A0(n16131), .A1(n15529), .B0(n15528), .B1(n16079), .Y(n16153));
  NAND4X1 g12823(.A(n16152), .B(n16151), .C(n16150), .D(n16153), .Y(P1_U3079));
  NAND2X1 g12824(.A(n16140), .B(P1_INSTQUEUE_REG_5__5__SCAN_IN), .Y(n16155));
  NAND2X1 g12825(.A(n16144), .B(n15535), .Y(n16156));
  NAND2X1 g12826(.A(n16133), .B(n15539), .Y(n16157));
  AOI22X1 g12827(.A0(n16131), .A1(n15544), .B0(n15543), .B1(n16079), .Y(n16158));
  NAND4X1 g12828(.A(n16157), .B(n16156), .C(n16155), .D(n16158), .Y(P1_U3078));
  NAND2X1 g12829(.A(n16140), .B(P1_INSTQUEUE_REG_5__4__SCAN_IN), .Y(n16160));
  NAND2X1 g12830(.A(n16144), .B(n15550), .Y(n16161));
  NAND2X1 g12831(.A(n16133), .B(n15554), .Y(n16162));
  AOI22X1 g12832(.A0(n16131), .A1(n15559), .B0(n15558), .B1(n16079), .Y(n16163));
  NAND4X1 g12833(.A(n16162), .B(n16161), .C(n16160), .D(n16163), .Y(P1_U3077));
  NAND2X1 g12834(.A(n16140), .B(P1_INSTQUEUE_REG_5__3__SCAN_IN), .Y(n16165));
  NAND2X1 g12835(.A(n16144), .B(n15565), .Y(n16166));
  OAI22X1 g12836(.A0(n16137), .A1(n15574), .B0(n15573), .B1(n16146), .Y(n16167));
  AOI21X1 g12837(.A0(n16133), .A1(n15569), .B0(n16167), .Y(n16168));
  NAND3X1 g12838(.A(n16168), .B(n16166), .C(n16165), .Y(P1_U3076));
  NAND2X1 g12839(.A(n16140), .B(P1_INSTQUEUE_REG_5__2__SCAN_IN), .Y(n16170));
  NAND2X1 g12840(.A(n16144), .B(n15581), .Y(n16171));
  OAI22X1 g12841(.A0(n16137), .A1(n15590), .B0(n15589), .B1(n16146), .Y(n16172));
  AOI21X1 g12842(.A0(n16133), .A1(n15585), .B0(n16172), .Y(n16173));
  NAND3X1 g12843(.A(n16173), .B(n16171), .C(n16170), .Y(P1_U3075));
  NAND2X1 g12844(.A(n16140), .B(P1_INSTQUEUE_REG_5__1__SCAN_IN), .Y(n16175));
  NAND2X1 g12845(.A(n16144), .B(n15597), .Y(n16176));
  OAI22X1 g12846(.A0(n16137), .A1(n15606), .B0(n15605), .B1(n16146), .Y(n16177));
  AOI21X1 g12847(.A0(n16133), .A1(n15601), .B0(n16177), .Y(n16178));
  NAND3X1 g12848(.A(n16178), .B(n16176), .C(n16175), .Y(P1_U3074));
  NAND2X1 g12849(.A(n16140), .B(P1_INSTQUEUE_REG_5__0__SCAN_IN), .Y(n16180));
  NAND2X1 g12850(.A(n16144), .B(n15613), .Y(n16181));
  OAI22X1 g12851(.A0(n16137), .A1(n15622), .B0(n15621), .B1(n16146), .Y(n16182));
  AOI21X1 g12852(.A0(n16133), .A1(n15617), .B0(n16182), .Y(n16183));
  NAND3X1 g12853(.A(n16183), .B(n16181), .C(n16180), .Y(P1_U3073));
  NOR4X1  g12854(.A(n14656), .B(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .D(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .Y(n16185));
  AOI21X1 g12855(.A0(n16022), .A1(n15744), .B0(n16185), .Y(n16186));
  NOR4X1  g12856(.A(n15746), .B(n15434), .C(n15407), .D(n15483), .Y(n16187));
  NOR4X1  g12857(.A(n16187), .B(n15354), .C(n15353), .D(n16133), .Y(n16189));
  OAI21X1 g12858(.A0(n16189), .A1(n15351), .B0(n16186), .Y(n16190));
  INVX1   g12859(.A(n16185), .Y(n16191));
  NAND2X1 g12860(.A(n16029), .B(n15147), .Y(n16192));
  AOI22X1 g12861(.A0(n16191), .A1(P1_STATE2_REG_3__SCAN_IN), .B0(P1_STATE2_REG_2__SCAN_IN), .B1(n16192), .Y(n16193));
  NAND3X1 g12862(.A(n16193), .B(n16190), .C(n15346), .Y(n16194));
  NAND2X1 g12863(.A(n16194), .B(P1_INSTQUEUE_REG_4__7__SCAN_IN), .Y(n16195));
  NOR3X1  g12864(.A(n16133), .B(n16187), .C(n15353), .Y(n16196));
  NOR2X1  g12865(.A(n16196), .B(n15351), .Y(n16197));
  OAI22X1 g12866(.A0(n16192), .A1(n15155), .B0(n16186), .B1(n16197), .Y(n16198));
  NAND2X1 g12867(.A(n16198), .B(n15500), .Y(n16199));
  INVX1   g12868(.A(n16133), .Y(n16200));
  OAI22X1 g12869(.A0(n16191), .A1(n15513), .B0(n15512), .B1(n16200), .Y(n16201));
  AOI21X1 g12870(.A0(n16187), .A1(n15507), .B0(n16201), .Y(n16202));
  NAND3X1 g12871(.A(n16202), .B(n16199), .C(n16195), .Y(P1_U3072));
  NAND2X1 g12872(.A(n16194), .B(P1_INSTQUEUE_REG_4__6__SCAN_IN), .Y(n16204));
  NAND2X1 g12873(.A(n16198), .B(n15520), .Y(n16205));
  NAND2X1 g12874(.A(n16187), .B(n15524), .Y(n16206));
  AOI22X1 g12875(.A0(n16185), .A1(n15529), .B0(n15528), .B1(n16133), .Y(n16207));
  NAND4X1 g12876(.A(n16206), .B(n16205), .C(n16204), .D(n16207), .Y(P1_U3071));
  NAND2X1 g12877(.A(n16194), .B(P1_INSTQUEUE_REG_4__5__SCAN_IN), .Y(n16209));
  NAND2X1 g12878(.A(n16198), .B(n15535), .Y(n16210));
  NAND2X1 g12879(.A(n16187), .B(n15539), .Y(n16211));
  AOI22X1 g12880(.A0(n16185), .A1(n15544), .B0(n15543), .B1(n16133), .Y(n16212));
  NAND4X1 g12881(.A(n16211), .B(n16210), .C(n16209), .D(n16212), .Y(P1_U3070));
  NAND2X1 g12882(.A(n16194), .B(P1_INSTQUEUE_REG_4__4__SCAN_IN), .Y(n16214));
  NAND2X1 g12883(.A(n16198), .B(n15550), .Y(n16215));
  NAND2X1 g12884(.A(n16187), .B(n15554), .Y(n16216));
  AOI22X1 g12885(.A0(n16185), .A1(n15559), .B0(n15558), .B1(n16133), .Y(n16217));
  NAND4X1 g12886(.A(n16216), .B(n16215), .C(n16214), .D(n16217), .Y(P1_U3069));
  NAND2X1 g12887(.A(n16194), .B(P1_INSTQUEUE_REG_4__3__SCAN_IN), .Y(n16219));
  NAND2X1 g12888(.A(n16198), .B(n15565), .Y(n16220));
  OAI22X1 g12889(.A0(n16191), .A1(n15574), .B0(n15573), .B1(n16200), .Y(n16221));
  AOI21X1 g12890(.A0(n16187), .A1(n15569), .B0(n16221), .Y(n16222));
  NAND3X1 g12891(.A(n16222), .B(n16220), .C(n16219), .Y(P1_U3068));
  NAND2X1 g12892(.A(n16194), .B(P1_INSTQUEUE_REG_4__2__SCAN_IN), .Y(n16224));
  NAND2X1 g12893(.A(n16198), .B(n15581), .Y(n16225));
  OAI22X1 g12894(.A0(n16191), .A1(n15590), .B0(n15589), .B1(n16200), .Y(n16226));
  AOI21X1 g12895(.A0(n16187), .A1(n15585), .B0(n16226), .Y(n16227));
  NAND3X1 g12896(.A(n16227), .B(n16225), .C(n16224), .Y(P1_U3067));
  NAND2X1 g12897(.A(n16194), .B(P1_INSTQUEUE_REG_4__1__SCAN_IN), .Y(n16229));
  NAND2X1 g12898(.A(n16198), .B(n15597), .Y(n16230));
  OAI22X1 g12899(.A0(n16191), .A1(n15606), .B0(n15605), .B1(n16200), .Y(n16231));
  AOI21X1 g12900(.A0(n16187), .A1(n15601), .B0(n16231), .Y(n16232));
  NAND3X1 g12901(.A(n16232), .B(n16230), .C(n16229), .Y(P1_U3066));
  NAND2X1 g12902(.A(n16194), .B(P1_INSTQUEUE_REG_4__0__SCAN_IN), .Y(n16234));
  NAND2X1 g12903(.A(n16198), .B(n15613), .Y(n16235));
  OAI22X1 g12904(.A0(n16191), .A1(n15622), .B0(n15621), .B1(n16200), .Y(n16236));
  AOI21X1 g12905(.A0(n16187), .A1(n15617), .B0(n16236), .Y(n16237));
  NAND3X1 g12906(.A(n16237), .B(n16235), .C(n16234), .Y(P1_U3065));
  NOR4X1  g12907(.A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n14659), .C(n14658), .D(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .Y(n16239));
  NOR2X1  g12908(.A(n15218), .B(n15802), .Y(n16240));
  AOI21X1 g12909(.A0(n16240), .A1(n15349), .B0(n16239), .Y(n16241));
  NOR4X1  g12910(.A(n15746), .B(n15434), .C(n15408), .D(n15483), .Y(n16242));
  NOR4X1  g12911(.A(n16242), .B(n15354), .C(n15353), .D(n16187), .Y(n16244));
  OAI21X1 g12912(.A0(n16244), .A1(n15351), .B0(n16241), .Y(n16245));
  INVX1   g12913(.A(n16239), .Y(n16246));
  NOR2X1  g12914(.A(n15866), .B(n15810), .Y(n16247));
  AOI21X1 g12915(.A0(n16247), .A1(n15493), .B0(n16239), .Y(n16248));
  AOI22X1 g12916(.A0(n16246), .A1(P1_STATE2_REG_3__SCAN_IN), .B0(P1_STATE2_REG_2__SCAN_IN), .B1(n16248), .Y(n16249));
  NAND3X1 g12917(.A(n16249), .B(n16245), .C(n15346), .Y(n16250));
  NAND2X1 g12918(.A(n16250), .B(P1_INSTQUEUE_REG_3__7__SCAN_IN), .Y(n16251));
  NOR3X1  g12919(.A(n16187), .B(n16242), .C(n15353), .Y(n16252));
  NOR2X1  g12920(.A(n16252), .B(n15351), .Y(n16253));
  OAI22X1 g12921(.A0(n16248), .A1(n15155), .B0(n16241), .B1(n16253), .Y(n16254));
  NAND2X1 g12922(.A(n16254), .B(n15500), .Y(n16255));
  INVX1   g12923(.A(n16187), .Y(n16256));
  OAI22X1 g12924(.A0(n16246), .A1(n15513), .B0(n15512), .B1(n16256), .Y(n16257));
  AOI21X1 g12925(.A0(n16242), .A1(n15507), .B0(n16257), .Y(n16258));
  NAND3X1 g12926(.A(n16258), .B(n16255), .C(n16251), .Y(P1_U3064));
  NAND2X1 g12927(.A(n16250), .B(P1_INSTQUEUE_REG_3__6__SCAN_IN), .Y(n16260));
  NAND2X1 g12928(.A(n16254), .B(n15520), .Y(n16261));
  NAND2X1 g12929(.A(n16242), .B(n15524), .Y(n16262));
  AOI22X1 g12930(.A0(n16239), .A1(n15529), .B0(n15528), .B1(n16187), .Y(n16263));
  NAND4X1 g12931(.A(n16262), .B(n16261), .C(n16260), .D(n16263), .Y(P1_U3063));
  NAND2X1 g12932(.A(n16250), .B(P1_INSTQUEUE_REG_3__5__SCAN_IN), .Y(n16265));
  NAND2X1 g12933(.A(n16254), .B(n15535), .Y(n16266));
  NAND2X1 g12934(.A(n16242), .B(n15539), .Y(n16267));
  AOI22X1 g12935(.A0(n16239), .A1(n15544), .B0(n15543), .B1(n16187), .Y(n16268));
  NAND4X1 g12936(.A(n16267), .B(n16266), .C(n16265), .D(n16268), .Y(P1_U3062));
  NAND2X1 g12937(.A(n16250), .B(P1_INSTQUEUE_REG_3__4__SCAN_IN), .Y(n16270));
  NAND2X1 g12938(.A(n16254), .B(n15550), .Y(n16271));
  NAND2X1 g12939(.A(n16242), .B(n15554), .Y(n16272));
  AOI22X1 g12940(.A0(n16239), .A1(n15559), .B0(n15558), .B1(n16187), .Y(n16273));
  NAND4X1 g12941(.A(n16272), .B(n16271), .C(n16270), .D(n16273), .Y(P1_U3061));
  NAND2X1 g12942(.A(n16250), .B(P1_INSTQUEUE_REG_3__3__SCAN_IN), .Y(n16275));
  NAND2X1 g12943(.A(n16254), .B(n15565), .Y(n16276));
  OAI22X1 g12944(.A0(n16246), .A1(n15574), .B0(n15573), .B1(n16256), .Y(n16277));
  AOI21X1 g12945(.A0(n16242), .A1(n15569), .B0(n16277), .Y(n16278));
  NAND3X1 g12946(.A(n16278), .B(n16276), .C(n16275), .Y(P1_U3060));
  NAND2X1 g12947(.A(n16250), .B(P1_INSTQUEUE_REG_3__2__SCAN_IN), .Y(n16280));
  NAND2X1 g12948(.A(n16254), .B(n15581), .Y(n16281));
  OAI22X1 g12949(.A0(n16246), .A1(n15590), .B0(n15589), .B1(n16256), .Y(n16282));
  AOI21X1 g12950(.A0(n16242), .A1(n15585), .B0(n16282), .Y(n16283));
  NAND3X1 g12951(.A(n16283), .B(n16281), .C(n16280), .Y(P1_U3059));
  NAND2X1 g12952(.A(n16250), .B(P1_INSTQUEUE_REG_3__1__SCAN_IN), .Y(n16285));
  NAND2X1 g12953(.A(n16254), .B(n15597), .Y(n16286));
  OAI22X1 g12954(.A0(n16246), .A1(n15606), .B0(n15605), .B1(n16256), .Y(n16287));
  AOI21X1 g12955(.A0(n16242), .A1(n15601), .B0(n16287), .Y(n16288));
  NAND3X1 g12956(.A(n16288), .B(n16286), .C(n16285), .Y(P1_U3058));
  NAND2X1 g12957(.A(n16250), .B(P1_INSTQUEUE_REG_3__0__SCAN_IN), .Y(n16290));
  NAND2X1 g12958(.A(n16254), .B(n15613), .Y(n16291));
  OAI22X1 g12959(.A0(n16246), .A1(n15622), .B0(n15621), .B1(n16256), .Y(n16292));
  AOI21X1 g12960(.A0(n16242), .A1(n15617), .B0(n16292), .Y(n16293));
  NAND3X1 g12961(.A(n16293), .B(n16291), .C(n16290), .Y(P1_U3057));
  NOR4X1  g12962(.A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n14659), .C(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .D(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .Y(n16295));
  AOI21X1 g12963(.A0(n16240), .A1(n15627), .B0(n16295), .Y(n16296));
  NOR4X1  g12964(.A(n15746), .B(n15629), .C(n15407), .D(n15483), .Y(n16297));
  NOR4X1  g12965(.A(n16297), .B(n15354), .C(n15353), .D(n16242), .Y(n16299));
  OAI21X1 g12966(.A0(n16299), .A1(n15351), .B0(n16296), .Y(n16300));
  INVX1   g12967(.A(n16295), .Y(n16301));
  NAND3X1 g12968(.A(n15215), .B(n15185), .C(n15637), .Y(n16302));
  AOI22X1 g12969(.A0(n16301), .A1(P1_STATE2_REG_3__SCAN_IN), .B0(P1_STATE2_REG_2__SCAN_IN), .B1(n16302), .Y(n16303));
  NAND3X1 g12970(.A(n16303), .B(n16300), .C(n15346), .Y(n16304));
  NAND2X1 g12971(.A(n16304), .B(P1_INSTQUEUE_REG_2__7__SCAN_IN), .Y(n16305));
  NOR3X1  g12972(.A(n16242), .B(n16297), .C(n15353), .Y(n16306));
  NOR2X1  g12973(.A(n16306), .B(n15351), .Y(n16307));
  OAI22X1 g12974(.A0(n16302), .A1(n15155), .B0(n16296), .B1(n16307), .Y(n16308));
  NAND2X1 g12975(.A(n16308), .B(n15500), .Y(n16309));
  INVX1   g12976(.A(n16242), .Y(n16310));
  OAI22X1 g12977(.A0(n16301), .A1(n15513), .B0(n15512), .B1(n16310), .Y(n16311));
  AOI21X1 g12978(.A0(n16297), .A1(n15507), .B0(n16311), .Y(n16312));
  NAND3X1 g12979(.A(n16312), .B(n16309), .C(n16305), .Y(P1_U3056));
  NAND2X1 g12980(.A(n16304), .B(P1_INSTQUEUE_REG_2__6__SCAN_IN), .Y(n16314));
  NAND2X1 g12981(.A(n16308), .B(n15520), .Y(n16315));
  NAND2X1 g12982(.A(n16297), .B(n15524), .Y(n16316));
  AOI22X1 g12983(.A0(n16295), .A1(n15529), .B0(n15528), .B1(n16242), .Y(n16317));
  NAND4X1 g12984(.A(n16316), .B(n16315), .C(n16314), .D(n16317), .Y(P1_U3055));
  NAND2X1 g12985(.A(n16304), .B(P1_INSTQUEUE_REG_2__5__SCAN_IN), .Y(n16319));
  NAND2X1 g12986(.A(n16308), .B(n15535), .Y(n16320));
  NAND2X1 g12987(.A(n16297), .B(n15539), .Y(n16321));
  AOI22X1 g12988(.A0(n16295), .A1(n15544), .B0(n15543), .B1(n16242), .Y(n16322));
  NAND4X1 g12989(.A(n16321), .B(n16320), .C(n16319), .D(n16322), .Y(P1_U3054));
  NAND2X1 g12990(.A(n16304), .B(P1_INSTQUEUE_REG_2__4__SCAN_IN), .Y(n16324));
  NAND2X1 g12991(.A(n16308), .B(n15550), .Y(n16325));
  NAND2X1 g12992(.A(n16297), .B(n15554), .Y(n16326));
  AOI22X1 g12993(.A0(n16295), .A1(n15559), .B0(n15558), .B1(n16242), .Y(n16327));
  NAND4X1 g12994(.A(n16326), .B(n16325), .C(n16324), .D(n16327), .Y(P1_U3053));
  NAND2X1 g12995(.A(n16304), .B(P1_INSTQUEUE_REG_2__3__SCAN_IN), .Y(n16329));
  NAND2X1 g12996(.A(n16308), .B(n15565), .Y(n16330));
  OAI22X1 g12997(.A0(n16301), .A1(n15574), .B0(n15573), .B1(n16310), .Y(n16331));
  AOI21X1 g12998(.A0(n16297), .A1(n15569), .B0(n16331), .Y(n16332));
  NAND3X1 g12999(.A(n16332), .B(n16330), .C(n16329), .Y(P1_U3052));
  NAND2X1 g13000(.A(n16304), .B(P1_INSTQUEUE_REG_2__2__SCAN_IN), .Y(n16334));
  NAND2X1 g13001(.A(n16308), .B(n15581), .Y(n16335));
  OAI22X1 g13002(.A0(n16301), .A1(n15590), .B0(n15589), .B1(n16310), .Y(n16336));
  AOI21X1 g13003(.A0(n16297), .A1(n15585), .B0(n16336), .Y(n16337));
  NAND3X1 g13004(.A(n16337), .B(n16335), .C(n16334), .Y(P1_U3051));
  NAND2X1 g13005(.A(n16304), .B(P1_INSTQUEUE_REG_2__1__SCAN_IN), .Y(n16339));
  NAND2X1 g13006(.A(n16308), .B(n15597), .Y(n16340));
  OAI22X1 g13007(.A0(n16301), .A1(n15606), .B0(n15605), .B1(n16310), .Y(n16341));
  AOI21X1 g13008(.A0(n16297), .A1(n15601), .B0(n16341), .Y(n16342));
  NAND3X1 g13009(.A(n16342), .B(n16340), .C(n16339), .Y(P1_U3050));
  NAND2X1 g13010(.A(n16304), .B(P1_INSTQUEUE_REG_2__0__SCAN_IN), .Y(n16344));
  NAND2X1 g13011(.A(n16308), .B(n15613), .Y(n16345));
  OAI22X1 g13012(.A0(n16301), .A1(n15622), .B0(n15621), .B1(n16310), .Y(n16346));
  AOI21X1 g13013(.A0(n16297), .A1(n15617), .B0(n16346), .Y(n16347));
  NAND3X1 g13014(.A(n16347), .B(n16345), .C(n16344), .Y(P1_U3049));
  NOR4X1  g13015(.A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C(n14658), .D(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .Y(n16349));
  AOI21X1 g13016(.A0(n16240), .A1(n15686), .B0(n16349), .Y(n16350));
  NOR4X1  g13017(.A(n15746), .B(n15629), .C(n15408), .D(n15483), .Y(n16351));
  NOR4X1  g13018(.A(n16351), .B(n15354), .C(n15353), .D(n16297), .Y(n16353));
  OAI21X1 g13019(.A0(n16353), .A1(n15351), .B0(n16350), .Y(n16354));
  INVX1   g13020(.A(n16349), .Y(n16355));
  AOI21X1 g13021(.A0(n16247), .A1(n15695), .B0(n16349), .Y(n16356));
  AOI22X1 g13022(.A0(n16355), .A1(P1_STATE2_REG_3__SCAN_IN), .B0(P1_STATE2_REG_2__SCAN_IN), .B1(n16356), .Y(n16357));
  NAND3X1 g13023(.A(n16357), .B(n16354), .C(n15346), .Y(n16358));
  NAND2X1 g13024(.A(n16358), .B(P1_INSTQUEUE_REG_1__7__SCAN_IN), .Y(n16359));
  NOR3X1  g13025(.A(n16297), .B(n16351), .C(n15353), .Y(n16360));
  NOR2X1  g13026(.A(n16360), .B(n15351), .Y(n16361));
  OAI22X1 g13027(.A0(n16356), .A1(n15155), .B0(n16350), .B1(n16361), .Y(n16362));
  NAND2X1 g13028(.A(n16362), .B(n15500), .Y(n16363));
  INVX1   g13029(.A(n16297), .Y(n16364));
  OAI22X1 g13030(.A0(n16355), .A1(n15513), .B0(n15512), .B1(n16364), .Y(n16365));
  AOI21X1 g13031(.A0(n16351), .A1(n15507), .B0(n16365), .Y(n16366));
  NAND3X1 g13032(.A(n16366), .B(n16363), .C(n16359), .Y(P1_U3048));
  NAND2X1 g13033(.A(n16358), .B(P1_INSTQUEUE_REG_1__6__SCAN_IN), .Y(n16368));
  NAND2X1 g13034(.A(n16362), .B(n15520), .Y(n16369));
  NAND2X1 g13035(.A(n16351), .B(n15524), .Y(n16370));
  AOI22X1 g13036(.A0(n16349), .A1(n15529), .B0(n15528), .B1(n16297), .Y(n16371));
  NAND4X1 g13037(.A(n16370), .B(n16369), .C(n16368), .D(n16371), .Y(P1_U3047));
  NAND2X1 g13038(.A(n16358), .B(P1_INSTQUEUE_REG_1__5__SCAN_IN), .Y(n16373));
  NAND2X1 g13039(.A(n16362), .B(n15535), .Y(n16374));
  NAND2X1 g13040(.A(n16351), .B(n15539), .Y(n16375));
  AOI22X1 g13041(.A0(n16349), .A1(n15544), .B0(n15543), .B1(n16297), .Y(n16376));
  NAND4X1 g13042(.A(n16375), .B(n16374), .C(n16373), .D(n16376), .Y(P1_U3046));
  NAND2X1 g13043(.A(n16358), .B(P1_INSTQUEUE_REG_1__4__SCAN_IN), .Y(n16378));
  NAND2X1 g13044(.A(n16362), .B(n15550), .Y(n16379));
  NAND2X1 g13045(.A(n16351), .B(n15554), .Y(n16380));
  AOI22X1 g13046(.A0(n16349), .A1(n15559), .B0(n15558), .B1(n16297), .Y(n16381));
  NAND4X1 g13047(.A(n16380), .B(n16379), .C(n16378), .D(n16381), .Y(P1_U3045));
  NAND2X1 g13048(.A(n16358), .B(P1_INSTQUEUE_REG_1__3__SCAN_IN), .Y(n16383));
  NAND2X1 g13049(.A(n16362), .B(n15565), .Y(n16384));
  OAI22X1 g13050(.A0(n16355), .A1(n15574), .B0(n15573), .B1(n16364), .Y(n16385));
  AOI21X1 g13051(.A0(n16351), .A1(n15569), .B0(n16385), .Y(n16386));
  NAND3X1 g13052(.A(n16386), .B(n16384), .C(n16383), .Y(P1_U3044));
  NAND2X1 g13053(.A(n16358), .B(P1_INSTQUEUE_REG_1__2__SCAN_IN), .Y(n16388));
  NAND2X1 g13054(.A(n16362), .B(n15581), .Y(n16389));
  OAI22X1 g13055(.A0(n16355), .A1(n15590), .B0(n15589), .B1(n16364), .Y(n16390));
  AOI21X1 g13056(.A0(n16351), .A1(n15585), .B0(n16390), .Y(n16391));
  NAND3X1 g13057(.A(n16391), .B(n16389), .C(n16388), .Y(P1_U3043));
  NAND2X1 g13058(.A(n16358), .B(P1_INSTQUEUE_REG_1__1__SCAN_IN), .Y(n16393));
  NAND2X1 g13059(.A(n16362), .B(n15597), .Y(n16394));
  OAI22X1 g13060(.A0(n16355), .A1(n15606), .B0(n15605), .B1(n16364), .Y(n16395));
  AOI21X1 g13061(.A0(n16351), .A1(n15601), .B0(n16395), .Y(n16396));
  NAND3X1 g13062(.A(n16396), .B(n16394), .C(n16393), .Y(P1_U3042));
  NAND2X1 g13063(.A(n16358), .B(P1_INSTQUEUE_REG_1__0__SCAN_IN), .Y(n16398));
  NAND2X1 g13064(.A(n16362), .B(n15613), .Y(n16399));
  OAI22X1 g13065(.A0(n16355), .A1(n15622), .B0(n15621), .B1(n16364), .Y(n16400));
  AOI21X1 g13066(.A0(n16351), .A1(n15617), .B0(n16400), .Y(n16401));
  NAND3X1 g13067(.A(n16401), .B(n16399), .C(n16398), .Y(P1_U3041));
  NOR4X1  g13068(.A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .D(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .Y(n16403));
  AOI21X1 g13069(.A0(n16240), .A1(n15744), .B0(n16403), .Y(n16404));
  NOR4X1  g13070(.A(n15488), .B(n15354), .C(n15353), .D(n16351), .Y(n16407));
  OAI21X1 g13071(.A0(n16407), .A1(n15351), .B0(n16404), .Y(n16408));
  INVX1   g13072(.A(n16403), .Y(n16409));
  NAND3X1 g13073(.A(n15215), .B(n15185), .C(n15147), .Y(n16410));
  AOI22X1 g13074(.A0(n16409), .A1(P1_STATE2_REG_3__SCAN_IN), .B0(P1_STATE2_REG_2__SCAN_IN), .B1(n16410), .Y(n16411));
  NAND3X1 g13075(.A(n16411), .B(n16408), .C(n15346), .Y(n16412));
  NAND2X1 g13076(.A(n16412), .B(P1_INSTQUEUE_REG_0__7__SCAN_IN), .Y(n16413));
  NOR3X1  g13077(.A(n16351), .B(n15488), .C(n15353), .Y(n16414));
  NOR2X1  g13078(.A(n16414), .B(n15351), .Y(n16415));
  OAI22X1 g13079(.A0(n16410), .A1(n15155), .B0(n16404), .B1(n16415), .Y(n16416));
  NAND2X1 g13080(.A(n16416), .B(n15500), .Y(n16417));
  INVX1   g13081(.A(n16351), .Y(n16418));
  OAI22X1 g13082(.A0(n16409), .A1(n15513), .B0(n15512), .B1(n16418), .Y(n16419));
  AOI21X1 g13083(.A0(n15488), .A1(n15507), .B0(n16419), .Y(n16420));
  NAND3X1 g13084(.A(n16420), .B(n16417), .C(n16413), .Y(P1_U3040));
  NAND2X1 g13085(.A(n16412), .B(P1_INSTQUEUE_REG_0__6__SCAN_IN), .Y(n16422));
  NAND2X1 g13086(.A(n16416), .B(n15520), .Y(n16423));
  NAND2X1 g13087(.A(n15488), .B(n15524), .Y(n16424));
  AOI22X1 g13088(.A0(n16403), .A1(n15529), .B0(n15528), .B1(n16351), .Y(n16425));
  NAND4X1 g13089(.A(n16424), .B(n16423), .C(n16422), .D(n16425), .Y(P1_U3039));
  NAND2X1 g13090(.A(n16412), .B(P1_INSTQUEUE_REG_0__5__SCAN_IN), .Y(n16427));
  NAND2X1 g13091(.A(n16416), .B(n15535), .Y(n16428));
  NAND2X1 g13092(.A(n15488), .B(n15539), .Y(n16429));
  AOI22X1 g13093(.A0(n16403), .A1(n15544), .B0(n15543), .B1(n16351), .Y(n16430));
  NAND4X1 g13094(.A(n16429), .B(n16428), .C(n16427), .D(n16430), .Y(P1_U3038));
  NAND2X1 g13095(.A(n16412), .B(P1_INSTQUEUE_REG_0__4__SCAN_IN), .Y(n16432));
  NAND2X1 g13096(.A(n16416), .B(n15550), .Y(n16433));
  NAND2X1 g13097(.A(n15488), .B(n15554), .Y(n16434));
  AOI22X1 g13098(.A0(n16403), .A1(n15559), .B0(n15558), .B1(n16351), .Y(n16435));
  NAND4X1 g13099(.A(n16434), .B(n16433), .C(n16432), .D(n16435), .Y(P1_U3037));
  NAND2X1 g13100(.A(n16412), .B(P1_INSTQUEUE_REG_0__3__SCAN_IN), .Y(n16437));
  NAND2X1 g13101(.A(n16416), .B(n15565), .Y(n16438));
  OAI22X1 g13102(.A0(n16409), .A1(n15574), .B0(n15573), .B1(n16418), .Y(n16439));
  AOI21X1 g13103(.A0(n15488), .A1(n15569), .B0(n16439), .Y(n16440));
  NAND3X1 g13104(.A(n16440), .B(n16438), .C(n16437), .Y(P1_U3036));
  NAND2X1 g13105(.A(n16412), .B(P1_INSTQUEUE_REG_0__2__SCAN_IN), .Y(n16442));
  NAND2X1 g13106(.A(n16416), .B(n15581), .Y(n16443));
  OAI22X1 g13107(.A0(n16409), .A1(n15590), .B0(n15589), .B1(n16418), .Y(n16444));
  AOI21X1 g13108(.A0(n15488), .A1(n15585), .B0(n16444), .Y(n16445));
  NAND3X1 g13109(.A(n16445), .B(n16443), .C(n16442), .Y(P1_U3035));
  NAND2X1 g13110(.A(n16412), .B(P1_INSTQUEUE_REG_0__1__SCAN_IN), .Y(n16447));
  NAND2X1 g13111(.A(n16416), .B(n15597), .Y(n16448));
  OAI22X1 g13112(.A0(n16409), .A1(n15606), .B0(n15605), .B1(n16418), .Y(n16449));
  AOI21X1 g13113(.A0(n15488), .A1(n15601), .B0(n16449), .Y(n16450));
  NAND3X1 g13114(.A(n16450), .B(n16448), .C(n16447), .Y(P1_U3034));
  NAND2X1 g13115(.A(n16412), .B(P1_INSTQUEUE_REG_0__0__SCAN_IN), .Y(n16452));
  NAND2X1 g13116(.A(n16416), .B(n15613), .Y(n16453));
  OAI22X1 g13117(.A0(n16409), .A1(n15622), .B0(n15621), .B1(n16418), .Y(n16454));
  AOI21X1 g13118(.A0(n15488), .A1(n15617), .B0(n16454), .Y(n16455));
  NAND3X1 g13119(.A(n16455), .B(n16453), .C(n16452), .Y(P1_U3033));
  NOR4X1  g13120(.A(n15093), .B(n15155), .C(n15322), .D(n14650), .Y(n16457));
  AOI21X1 g13121(.A0(n14650), .A1(P1_STATE2_REG_3__SCAN_IN), .B0(n16457), .Y(n16458));
  OAI21X1 g13122(.A0(n15339), .A1(n15037), .B0(n16458), .Y(n16459));
  INVX1   g13123(.A(n15243), .Y(n16460));
  NAND4X1 g13124(.A(n16460), .B(n15309), .C(n15027), .D(n16459), .Y(n16461));
  OAI21X1 g13125(.A0(n16459), .A1(n14651), .B0(n16461), .Y(P1_U3468));
  INVX1   g13126(.A(n16459), .Y(n16463));
  AOI22X1 g13127(.A0(n15231), .A1(n15309), .B0(n15227), .B1(n15336), .Y(n16464));
  NAND2X1 g13128(.A(n16463), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n16465));
  OAI21X1 g13129(.A0(n16464), .A1(n16463), .B0(n16465), .Y(P1_U3469));
  AOI21X1 g13130(.A0(n15204), .A1(n15309), .B0(n15260), .Y(n16467));
  OAI21X1 g13131(.A0(n15344), .A1(n15197), .B0(n16467), .Y(n16468));
  NAND2X1 g13132(.A(n16468), .B(n16459), .Y(n16469));
  OAI21X1 g13133(.A0(n16459), .A1(n14655), .B0(n16469), .Y(P1_U3472));
  NAND2X1 g13134(.A(n15336), .B(n15170), .Y(n16471));
  AOI22X1 g13135(.A0(n15325), .A1(n15259), .B0(n15172), .B1(n15309), .Y(n16472));
  NAND2X1 g13136(.A(n16472), .B(n16471), .Y(n16473));
  NAND2X1 g13137(.A(n16473), .B(n16459), .Y(n16474));
  OAI21X1 g13138(.A0(n16459), .A1(n14657), .B0(n16474), .Y(P1_U3473));
  AOI21X1 g13139(.A0(n15140), .A1(n15309), .B0(n15328), .Y(n16476));
  OAI21X1 g13140(.A0(n15344), .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B0(n16476), .Y(n16477));
  NAND2X1 g13141(.A(n16477), .B(n16459), .Y(n16478));
  OAI21X1 g13142(.A0(n16459), .A1(n14670), .B0(n16478), .Y(P1_U3474));
  NOR2X1  g13143(.A(n15333), .B(n15319), .Y(n16480));
  NOR4X1  g13144(.A(n14650), .B(n15093), .C(n15155), .D(n16480), .Y(n16481));
  NOR4X1  g13145(.A(n16457), .B(n15346), .C(n14666), .D(n16481), .Y(P1_U3032));
  NOR3X1  g13146(.A(n16481), .B(n16457), .C(n15346), .Y(n16483));
  INVX1   g13147(.A(n16483), .Y(n16484));
  AOI21X1 g13148(.A0(n15746), .A1(n15486), .B0(n15484), .Y(n16486));
  NAND3X1 g13149(.A(n15746), .B(n15629), .C(n15407), .Y(n16487));
  OAI21X1 g13150(.A0(n16486), .A1(n15970), .B0(n16487), .Y(n16488));
  AOI21X1 g13151(.A0(n16488), .A1(n16092), .B0(n15353), .Y(n16489));
  INVX1   g13152(.A(n15351), .Y(n16490));
  NOR2X1  g13153(.A(n15093), .B(P1_STATE2_REG_3__SCAN_IN), .Y(n16491));
  OAI22X1 g13154(.A0(n15484), .A1(n16490), .B0(n15219), .B1(n16491), .Y(n16492));
  OAI21X1 g13155(.A0(n16492), .A1(n16489), .B0(n16484), .Y(n16493));
  OAI21X1 g13156(.A0(n16484), .A1(n14653), .B0(n16493), .Y(P1_U3475));
  XOR2X1  g13157(.A(n15459), .B(n15486), .Y(n16496));
  XOR2X1  g13158(.A(n16496), .B(n15631), .Y(n16497));
  NOR2X1  g13159(.A(n16497), .B(n15353), .Y(n16498));
  OAI22X1 g13160(.A0(n15459), .A1(n16490), .B0(n15192), .B1(n16491), .Y(n16499));
  OAI21X1 g13161(.A0(n16499), .A1(n16498), .B0(n16484), .Y(n16500));
  OAI21X1 g13162(.A0(n16484), .A1(n14656), .B0(n16500), .Y(P1_U3476));
  NAND2X1 g13163(.A(n15434), .B(n15408), .Y(n16502));
  NAND2X1 g13164(.A(n15434), .B(n15407), .Y(n16503));
  AOI21X1 g13165(.A0(n16503), .A1(n16502), .B0(n15353), .Y(n16504));
  OAI22X1 g13166(.A0(n15434), .A1(n16490), .B0(n15169), .B1(n16491), .Y(n16505));
  OAI21X1 g13167(.A0(n16505), .A1(n16504), .B0(n16484), .Y(n16506));
  OAI21X1 g13168(.A0(n16484), .A1(n14659), .B0(n16506), .Y(P1_U3477));
  NOR2X1  g13169(.A(P1_STATE2_REG_2__SCAN_IN), .B(P1_STATE2_REG_3__SCAN_IN), .Y(n16508));
  INVX1   g13170(.A(n16508), .Y(n16509));
  OAI22X1 g13171(.A0(n15407), .A1(n16509), .B0(n15132), .B1(n16491), .Y(n16510));
  OAI21X1 g13172(.A0(n16510), .A1(n15334), .B0(n16484), .Y(n16511));
  OAI21X1 g13173(.A0(n16484), .A1(n14658), .B0(n16511), .Y(P1_U3478));
  AOI22X1 g13174(.A0(n15024), .A1(n14707), .B0(n15020), .B1(n15394), .Y(n16513));
  OAI21X1 g13175(.A0(n15407), .A1(n14821), .B0(n16513), .Y(n16514));
  XOR2X1  g13176(.A(n16514), .B(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .Y(n16515));
  OAI21X1 g13177(.A0(n15276), .A1(n15268), .B0(n14770), .Y(n16516));
  NOR3X1  g13178(.A(n15272), .B(n14984), .C(n14549), .Y(n16517));
  NOR2X1  g13179(.A(n15026), .B(n15019), .Y(n16518));
  NAND4X1 g13180(.A(n14890), .B(n14887), .C(n14770), .D(n15133), .Y(n16519));
  AOI21X1 g13181(.A0(n15276), .A1(n14769), .B0(n14549), .Y(n16520));
  NAND4X1 g13182(.A(n14986), .B(n14963), .C(n15068), .D(n16520), .Y(n16521));
  NOR2X1  g13183(.A(n14992), .B(n14707), .Y(n16522));
  AOI21X1 g13184(.A0(n16522), .A1(n16521), .B0(n14985), .Y(n16523));
  NAND2X1 g13185(.A(n16523), .B(n15007), .Y(n16524));
  NAND3X1 g13186(.A(n16524), .B(n16519), .C(n16518), .Y(n16525));
  AOI21X1 g13187(.A0(n16517), .A1(n16516), .B0(n16525), .Y(n16526));
  NOR4X1  g13188(.A(P1_STATE2_REG_1__SCAN_IN), .B(P1_STATE2_REG_2__SCAN_IN), .C(P1_STATE2_REG_3__SCAN_IN), .D(P1_STATE2_REG_0__SCAN_IN), .Y(n16527));
  AOI21X1 g13189(.A0(n14919), .A1(n14801), .B0(n15157), .Y(n16528));
  AOI21X1 g13190(.A0(n16528), .A1(n14818), .B0(n16527), .Y(n16529));
  OAI21X1 g13191(.A0(n16526), .A1(n15339), .B0(n16529), .Y(n16530));
  NOR4X1  g13192(.A(n14993), .B(n14985), .C(n14803), .D(n15009), .Y(n16531));
  NOR4X1  g13193(.A(n14769), .B(n14707), .C(n15155), .D(n14987), .Y(n16532));
  NOR3X1  g13194(.A(n16532), .B(n16531), .C(n15027), .Y(n16533));
  NOR4X1  g13195(.A(n14985), .B(n14940), .C(n15021), .D(n15122), .Y(n16534));
  NOR3X1  g13196(.A(n16534), .B(n15117), .C(n15003), .Y(n16535));
  AOI21X1 g13197(.A0(n16535), .A1(n16533), .B0(n15155), .Y(n16536));
  NAND3X1 g13198(.A(n16536), .B(n16530), .C(n16515), .Y(n16537));
  INVX1   g13199(.A(n16530), .Y(n16538));
  AOI22X1 g13200(.A0(n16538), .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B0(P1_REIP_REG_0__SCAN_IN), .B1(n16527), .Y(n16540));
  NOR3X1  g13201(.A(n16538), .B(n15011), .C(n15155), .Y(n16541));
  AOI21X1 g13202(.A0(n15086), .A1(n15066), .B0(n15119), .Y(n16542));
  AOI21X1 g13203(.A0(n15063), .A1(n14707), .B0(n15074), .Y(n16543));
  NAND4X1 g13204(.A(n16542), .B(n15201), .C(n15061), .D(n16543), .Y(n16544));
  NAND3X1 g13205(.A(n16544), .B(n16530), .C(P1_STATE2_REG_2__SCAN_IN), .Y(n16545));
  INVX1   g13206(.A(n16545), .Y(n16546));
  OAI21X1 g13207(.A0(n16546), .A1(n16541), .B0(n15251), .Y(n16547));
  NOR3X1  g13208(.A(n16538), .B(n15198), .C(n15155), .Y(n16548));
  INVX1   g13209(.A(n15054), .Y(n16549));
  XOR2X1  g13210(.A(n15056), .B(n16549), .Y(n16550));
  OAI21X1 g13211(.A0(n15024), .A1(n14707), .B0(n16549), .Y(n16551));
  AOI21X1 g13212(.A0(n15124), .A1(n14769), .B0(n14707), .Y(n16552));
  INVX1   g13213(.A(n16552), .Y(n16553));
  AOI22X1 g13214(.A0(n16551), .A1(P1_EBX_REG_0__SCAN_IN), .B0(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(n16553), .Y(n16554));
  XOR2X1  g13215(.A(n16554), .B(n15054), .Y(n16555));
  XOR2X1  g13216(.A(n16555), .B(n16550), .Y(n16556));
  OAI21X1 g13217(.A0(n14987), .A1(n15021), .B0(n15103), .Y(n16557));
  NAND3X1 g13218(.A(n16557), .B(n16530), .C(P1_STATE2_REG_2__SCAN_IN), .Y(n16558));
  INVX1   g13219(.A(n16558), .Y(n16559));
  AOI22X1 g13220(.A0(n16556), .A1(n16559), .B0(n16548), .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .Y(n16560));
  NAND4X1 g13221(.A(n16547), .B(n16540), .C(n16537), .D(n16560), .Y(P1_U3031));
  NAND4X1 g13222(.A(n14994), .B(P1_STATE2_REG_2__SCAN_IN), .C(n15255), .D(n16530), .Y(n16562));
  INVX1   g13223(.A(n16555), .Y(n16563));
  NOR3X1  g13224(.A(n16549), .B(n15024), .C(n14707), .Y(n16564));
  AOI21X1 g13225(.A0(n16563), .A1(n16551), .B0(n16564), .Y(n16565));
  AOI22X1 g13226(.A0(n16551), .A1(P1_EBX_REG_1__SCAN_IN), .B0(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n16553), .Y(n16566));
  XOR2X1  g13227(.A(n16566), .B(n15054), .Y(n16567));
  XOR2X1  g13228(.A(n16567), .B(n16553), .Y(n16568));
  XOR2X1  g13229(.A(n16568), .B(n16565), .Y(n16569));
  AOI22X1 g13230(.A0(n16559), .A1(n16569), .B0(n16541), .B1(n15257), .Y(n16570));
  NAND2X1 g13231(.A(n16536), .B(n16530), .Y(n16571));
  INVX1   g13232(.A(n16571), .Y(n16572));
  XOR2X1  g13233(.A(n15425), .B(n15400), .Y(n16573));
  NOR2X1  g13234(.A(n14801), .B(n14707), .Y(n16574));
  NOR3X1  g13235(.A(n16574), .B(n14985), .C(n14940), .Y(n16575));
  OAI21X1 g13236(.A0(n16573), .A1(n15021), .B0(n16575), .Y(n16576));
  INVX1   g13237(.A(n16576), .Y(n16577));
  OAI21X1 g13238(.A0(n15434), .A1(n14821), .B0(n16577), .Y(n16578));
  NAND2X1 g13239(.A(n16514), .B(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .Y(n16579));
  XOR2X1  g13240(.A(n16579), .B(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .Y(n16580));
  NOR2X1  g13241(.A(n16580), .B(n16578), .Y(n16581));
  NAND3X1 g13242(.A(n16578), .B(n16514), .C(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .Y(n16582));
  NAND3X1 g13243(.A(n16579), .B(n16578), .C(n15255), .Y(n16583));
  OAI21X1 g13244(.A0(n16582), .A1(n15255), .B0(n16583), .Y(n16584));
  OAI21X1 g13245(.A0(n16584), .A1(n16581), .B0(n16572), .Y(n16585));
  INVX1   g13246(.A(n16527), .Y(n16586));
  OAI22X1 g13247(.A0(n16530), .A1(n15255), .B0(n14541), .B1(n16586), .Y(n16587));
  AOI21X1 g13248(.A0(n16546), .A1(n15257), .B0(n16587), .Y(n16588));
  NAND4X1 g13249(.A(n16585), .B(n16570), .C(n16562), .D(n16588), .Y(P1_U3030));
  AOI21X1 g13250(.A0(n16514), .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B0(n16578), .Y(n16590));
  OAI21X1 g13251(.A0(n16590), .A1(n15255), .B0(n16582), .Y(n16591));
  NOR2X1  g13252(.A(n15425), .B(n15394), .Y(n16592));
  XOR2X1  g13253(.A(n16592), .B(n15446), .Y(n16593));
  OAI22X1 g13254(.A0(n14940), .A1(n14806), .B0(n15021), .B1(n16593), .Y(n16594));
  INVX1   g13255(.A(n16594), .Y(n16595));
  OAI21X1 g13256(.A0(n15459), .A1(n14821), .B0(n16595), .Y(n16596));
  XOR2X1  g13257(.A(n16596), .B(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .Y(n16597));
  XOR2X1  g13258(.A(n16597), .B(n16591), .Y(n16598));
  NAND2X1 g13259(.A(n16598), .B(n16572), .Y(n16599));
  INVX1   g13260(.A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .Y(n16600));
  NAND2X1 g13261(.A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .Y(n16601));
  XOR2X1  g13262(.A(n16601), .B(n16600), .Y(n16602));
  OAI22X1 g13263(.A0(n16530), .A1(n16600), .B0(n14538), .B1(n16586), .Y(n16603));
  AOI21X1 g13264(.A0(n16602), .A1(n16546), .B0(n16603), .Y(n16604));
  XOR2X1  g13265(.A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .Y(n16605));
  NAND4X1 g13266(.A(n16530), .B(n14994), .C(P1_STATE2_REG_2__SCAN_IN), .D(n16605), .Y(n16606));
  XOR2X1  g13267(.A(n16601), .B(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .Y(n16607));
  AOI22X1 g13268(.A0(n16551), .A1(P1_EBX_REG_2__SCAN_IN), .B0(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B1(n16553), .Y(n16608));
  XOR2X1  g13269(.A(n16608), .B(n15054), .Y(n16609));
  NOR2X1  g13270(.A(n16567), .B(n16552), .Y(n16610));
  AOI21X1 g13271(.A0(n16567), .A1(n16552), .B0(n16565), .Y(n16611));
  NOR2X1  g13272(.A(n16611), .B(n16610), .Y(n16612));
  XOR2X1  g13273(.A(n16612), .B(n16609), .Y(n16613));
  AOI22X1 g13274(.A0(n16607), .A1(n16541), .B0(n16559), .B1(n16613), .Y(n16614));
  NAND4X1 g13275(.A(n16606), .B(n16604), .C(n16599), .D(n16614), .Y(P1_U3029));
  NAND2X1 g13276(.A(n16596), .B(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .Y(n16616));
  OAI21X1 g13277(.A0(n16596), .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B0(n16591), .Y(n16617));
  NAND2X1 g13278(.A(n16617), .B(n16616), .Y(n16618));
  NOR3X1  g13279(.A(n16592), .B(n15471), .C(n15446), .Y(n16619));
  OAI21X1 g13280(.A0(n16592), .A1(n15446), .B0(n15471), .Y(n16620));
  NAND3X1 g13281(.A(n16620), .B(n14769), .C(n14806), .Y(n16621));
  NOR2X1  g13282(.A(n16621), .B(n16619), .Y(n16622));
  AOI21X1 g13283(.A0(n15483), .A1(n14820), .B0(n16622), .Y(n16623));
  XOR2X1  g13284(.A(n16623), .B(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .Y(n16624));
  XOR2X1  g13285(.A(n16624), .B(n16618), .Y(n16625));
  AOI21X1 g13286(.A0(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B0(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .Y(n16627));
  XOR2X1  g13287(.A(n16627), .B(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .Y(n16628));
  AOI22X1 g13288(.A0(n16538), .A1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B0(P1_REIP_REG_3__SCAN_IN), .B1(n16527), .Y(n16629));
  OAI21X1 g13289(.A0(n16628), .A1(n18937), .B0(n16629), .Y(n16630));
  NOR2X1  g13290(.A(n16612), .B(n16609), .Y(n16631));
  AOI22X1 g13291(.A0(n16551), .A1(P1_EBX_REG_3__SCAN_IN), .B0(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(n16553), .Y(n16632));
  XOR2X1  g13292(.A(n16632), .B(n15054), .Y(n16633));
  XOR2X1  g13293(.A(n16633), .B(n16631), .Y(n16634));
  NOR2X1  g13294(.A(n16634), .B(n16558), .Y(n16635));
  INVX1   g13295(.A(n16548), .Y(n16636));
  INVX1   g13296(.A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .Y(n16637));
  NOR2X1  g13297(.A(n16601), .B(n16600), .Y(n16638));
  XOR2X1  g13298(.A(n16638), .B(n16637), .Y(n16639));
  NAND2X1 g13299(.A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .Y(n16640));
  XOR2X1  g13300(.A(n16640), .B(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .Y(n16641));
  OAI22X1 g13301(.A0(n16639), .A1(n16545), .B0(n16636), .B1(n16641), .Y(n16642));
  NOR3X1  g13302(.A(n16642), .B(n16635), .C(n16630), .Y(n16643));
  OAI21X1 g13303(.A0(n16625), .A1(n16571), .B0(n16643), .Y(P1_U3028));
  NAND2X1 g13304(.A(n16623), .B(n16637), .Y(n16645));
  NAND2X1 g13305(.A(n16645), .B(n16618), .Y(n16646));
  OAI21X1 g13306(.A0(n16623), .A1(n16637), .B0(n16646), .Y(n16647));
  AOI22X1 g13307(.A0(n15355), .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B0(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(n14673), .Y(n16648));
  AOI22X1 g13308(.A0(n14674), .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B0(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(n15359), .Y(n16649));
  AOI22X1 g13309(.A0(n15361), .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B0(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(n15362), .Y(n16650));
  AOI22X1 g13310(.A0(n14703), .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B0(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(n15365), .Y(n16651));
  NAND4X1 g13311(.A(n16650), .B(n16649), .C(n16648), .D(n16651), .Y(n16652));
  AOI22X1 g13312(.A0(n14680), .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B0(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(n14907), .Y(n16653));
  AOI22X1 g13313(.A0(n14704), .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B0(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(n15372), .Y(n16654));
  AOI22X1 g13314(.A0(n14671), .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B0(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(n15375), .Y(n16655));
  AOI22X1 g13315(.A0(n14682), .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B0(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(n15378), .Y(n16656));
  NAND4X1 g13316(.A(n16655), .B(n16654), .C(n16653), .D(n16656), .Y(n16657));
  NOR2X1  g13317(.A(n16657), .B(n16652), .Y(n16658));
  INVX1   g13318(.A(n16658), .Y(n16659));
  XOR2X1  g13319(.A(n16659), .B(n16620), .Y(n16660));
  NOR3X1  g13320(.A(n16660), .B(n14770), .C(n14707), .Y(n16661));
  AOI22X1 g13321(.A0(n14824), .A1(n16659), .B0(n14818), .B1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .Y(n16662));
  NOR4X1  g13322(.A(n15412), .B(n14846), .C(n14650), .D(n16658), .Y(n16663));
  NOR4X1  g13323(.A(n15381), .B(n14846), .C(n14650), .D(n16658), .Y(n16664));
  NOR2X1  g13324(.A(n16664), .B(n16663), .Y(n16665));
  XOR2X1  g13325(.A(n16665), .B(n16662), .Y(n16666));
  INVX1   g13326(.A(n15472), .Y(n16667));
  INVX1   g13327(.A(n15476), .Y(n16668));
  NOR2X1  g13328(.A(n15454), .B(n15411), .Y(n16669));
  OAI22X1 g13329(.A0(n15456), .A1(n16669), .B0(n15451), .B1(n15447), .Y(n16670));
  AOI22X1 g13330(.A0(n15472), .A1(n15476), .B0(n15451), .B1(n15447), .Y(n16671));
  AOI22X1 g13331(.A0(n16670), .A1(n16671), .B0(n16668), .B1(n16667), .Y(n16672));
  XOR2X1  g13332(.A(n16672), .B(n16666), .Y(n16673));
  INVX1   g13333(.A(n16673), .Y(n16674));
  AOI21X1 g13334(.A0(n16674), .A1(n14820), .B0(n16661), .Y(n16675));
  XOR2X1  g13335(.A(n16675), .B(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .Y(n16676));
  XOR2X1  g13336(.A(n16676), .B(n16647), .Y(n16677));
  INVX1   g13337(.A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .Y(n16678));
  NOR2X1  g13338(.A(n16627), .B(n16637), .Y(n16679));
  XOR2X1  g13339(.A(n16679), .B(n16678), .Y(n16680));
  AOI22X1 g13340(.A0(n16538), .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B0(P1_REIP_REG_4__SCAN_IN), .B1(n16527), .Y(n16681));
  OAI21X1 g13341(.A0(n16680), .A1(n18937), .B0(n16681), .Y(n16682));
  NAND4X1 g13342(.A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .C(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .D(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .Y(n16683));
  XOR2X1  g13343(.A(n16683), .B(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .Y(n16684));
  NOR2X1  g13344(.A(n16684), .B(n16545), .Y(n16685));
  AOI22X1 g13345(.A0(n16551), .A1(P1_EBX_REG_4__SCAN_IN), .B0(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .B1(n16553), .Y(n16686));
  XOR2X1  g13346(.A(n16686), .B(n15054), .Y(n16687));
  NOR3X1  g13347(.A(n16633), .B(n16612), .C(n16609), .Y(n16688));
  XOR2X1  g13348(.A(n16688), .B(n16687), .Y(n16689));
  NAND3X1 g13349(.A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .C(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .Y(n16690));
  XOR2X1  g13350(.A(n16690), .B(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .Y(n16691));
  OAI22X1 g13351(.A0(n16689), .A1(n16558), .B0(n16636), .B1(n16691), .Y(n16692));
  NOR3X1  g13352(.A(n16692), .B(n16685), .C(n16682), .Y(n16693));
  OAI21X1 g13353(.A0(n16677), .A1(n16571), .B0(n16693), .Y(P1_U3027));
  NAND2X1 g13354(.A(n16675), .B(n16678), .Y(n16695));
  NAND2X1 g13355(.A(n16695), .B(n16647), .Y(n16696));
  OAI21X1 g13356(.A0(n16675), .A1(n16678), .B0(n16696), .Y(n16697));
  INVX1   g13357(.A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .Y(n16698));
  NOR2X1  g13358(.A(n16658), .B(n16620), .Y(n16699));
  AOI22X1 g13359(.A0(n15355), .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B0(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(n14673), .Y(n16700));
  AOI22X1 g13360(.A0(n14674), .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B0(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(n15359), .Y(n16701));
  AOI22X1 g13361(.A0(n15361), .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B0(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(n15362), .Y(n16702));
  AOI22X1 g13362(.A0(n14703), .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B0(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(n15365), .Y(n16703));
  NAND4X1 g13363(.A(n16702), .B(n16701), .C(n16700), .D(n16703), .Y(n16704));
  AOI22X1 g13364(.A0(n14680), .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B0(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(n14907), .Y(n16705));
  AOI22X1 g13365(.A0(n14704), .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B0(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(n15372), .Y(n16706));
  AOI22X1 g13366(.A0(n14671), .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B0(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(n15375), .Y(n16707));
  AOI22X1 g13367(.A0(n14682), .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B0(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(n15378), .Y(n16708));
  NAND4X1 g13368(.A(n16707), .B(n16706), .C(n16705), .D(n16708), .Y(n16709));
  NOR2X1  g13369(.A(n16709), .B(n16704), .Y(n16710));
  XOR2X1  g13370(.A(n16710), .B(n16699), .Y(n16711));
  NOR3X1  g13371(.A(n16710), .B(n14806), .C(n14650), .Y(n16712));
  AOI21X1 g13372(.A0(n14818), .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B0(n16712), .Y(n16713));
  NOR4X1  g13373(.A(n15412), .B(n14846), .C(n14650), .D(n16710), .Y(n16714));
  NOR4X1  g13374(.A(n15381), .B(n14846), .C(n14650), .D(n16710), .Y(n16715));
  NOR2X1  g13375(.A(n16715), .B(n16714), .Y(n16716));
  XOR2X1  g13376(.A(n16716), .B(n16713), .Y(n16717));
  NOR2X1  g13377(.A(n16668), .B(n16667), .Y(n16718));
  NAND2X1 g13378(.A(n16665), .B(n16662), .Y(n16719));
  INVX1   g13379(.A(n16719), .Y(n16720));
  INVX1   g13380(.A(n16670), .Y(n16721));
  NOR4X1  g13381(.A(n16720), .B(n16718), .C(n15481), .D(n16721), .Y(n16722));
  NOR2X1  g13382(.A(n16665), .B(n16662), .Y(n16723));
  INVX1   g13383(.A(n16723), .Y(n16724));
  NOR3X1  g13384(.A(n16720), .B(n15476), .C(n15472), .Y(n16725));
  NOR2X1  g13385(.A(n16723), .B(n16722), .Y(n16728));
  XOR2X1  g13386(.A(n16728), .B(n16717), .Y(n16729));
  OAI22X1 g13387(.A0(n16711), .A1(n15021), .B0(n14821), .B1(n16729), .Y(n16730));
  INVX1   g13388(.A(n16730), .Y(n16731));
  NAND2X1 g13389(.A(n16731), .B(n16698), .Y(n16732));
  NAND2X1 g13390(.A(n16732), .B(n16697), .Y(n16733));
  NAND2X1 g13391(.A(n16730), .B(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .Y(n16734));
  INVX1   g13392(.A(n16734), .Y(n16735));
  XOR2X1  g13393(.A(n16730), .B(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .Y(n16736));
  OAI22X1 g13394(.A0(n16735), .A1(n16733), .B0(n16697), .B1(n16736), .Y(n16737));
  NOR3X1  g13395(.A(n16627), .B(n16637), .C(n16678), .Y(n16738));
  XOR2X1  g13396(.A(n16738), .B(n16698), .Y(n16739));
  AOI22X1 g13397(.A0(n16538), .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .B0(P1_REIP_REG_5__SCAN_IN), .B1(n16527), .Y(n16740));
  OAI21X1 g13398(.A0(n16739), .A1(n18937), .B0(n16740), .Y(n16741));
  NOR4X1  g13399(.A(n16600), .B(n16637), .C(n16678), .D(n16601), .Y(n16742));
  XOR2X1  g13400(.A(n16742), .B(n16698), .Y(n16743));
  NOR2X1  g13401(.A(n16743), .B(n16545), .Y(n16744));
  AOI22X1 g13402(.A0(n16551), .A1(P1_EBX_REG_5__SCAN_IN), .B0(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .B1(n16553), .Y(n16745));
  XOR2X1  g13403(.A(n16745), .B(n15054), .Y(n16746));
  NOR4X1  g13404(.A(n16633), .B(n16612), .C(n16609), .D(n16687), .Y(n16747));
  XOR2X1  g13405(.A(n16747), .B(n16746), .Y(n16748));
  NAND4X1 g13406(.A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .C(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .D(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .Y(n16749));
  XOR2X1  g13407(.A(n16749), .B(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .Y(n16750));
  OAI22X1 g13408(.A0(n16748), .A1(n16558), .B0(n16636), .B1(n16750), .Y(n16751));
  NOR3X1  g13409(.A(n16751), .B(n16744), .C(n16741), .Y(n16752));
  OAI21X1 g13410(.A0(n16737), .A1(n16571), .B0(n16752), .Y(P1_U3026));
  NOR3X1  g13411(.A(n16710), .B(n16658), .C(n16620), .Y(n16754));
  AOI22X1 g13412(.A0(n15355), .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B0(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(n14673), .Y(n16755));
  AOI22X1 g13413(.A0(n14674), .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B0(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(n15359), .Y(n16756));
  AOI22X1 g13414(.A0(n15361), .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B0(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(n15362), .Y(n16757));
  AOI22X1 g13415(.A0(n14703), .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B0(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(n15365), .Y(n16758));
  NAND4X1 g13416(.A(n16757), .B(n16756), .C(n16755), .D(n16758), .Y(n16759));
  AOI22X1 g13417(.A0(n14680), .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B0(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(n14907), .Y(n16760));
  AOI22X1 g13418(.A0(n14704), .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B0(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(n15372), .Y(n16761));
  AOI22X1 g13419(.A0(n14671), .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B0(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(n15375), .Y(n16762));
  AOI22X1 g13420(.A0(n14682), .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B0(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(n15378), .Y(n16763));
  NAND4X1 g13421(.A(n16762), .B(n16761), .C(n16760), .D(n16763), .Y(n16764));
  NOR2X1  g13422(.A(n16764), .B(n16759), .Y(n16765));
  XOR2X1  g13423(.A(n16765), .B(n16754), .Y(n16766));
  NOR2X1  g13424(.A(n16766), .B(n15021), .Y(n16767));
  NOR3X1  g13425(.A(n16765), .B(n14806), .C(n14650), .Y(n16768));
  AOI21X1 g13426(.A0(n14818), .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B0(n16768), .Y(n16769));
  NOR4X1  g13427(.A(n15412), .B(n14846), .C(n14650), .D(n16765), .Y(n16770));
  NOR4X1  g13428(.A(n15381), .B(n14846), .C(n14650), .D(n16765), .Y(n16771));
  NOR2X1  g13429(.A(n16771), .B(n16770), .Y(n16772));
  XOR2X1  g13430(.A(n16772), .B(n16769), .Y(n16773));
  NAND2X1 g13431(.A(n16716), .B(n16713), .Y(n16774));
  OAI21X1 g13432(.A0(n16723), .A1(n16722), .B0(n16774), .Y(n16775));
  NOR2X1  g13433(.A(n16716), .B(n16713), .Y(n16776));
  INVX1   g13434(.A(n16776), .Y(n16777));
  NAND2X1 g13435(.A(n16775), .B(n16777), .Y(n16778));
  NOR2X1  g13436(.A(n16773), .B(n16776), .Y(n16779));
  AOI22X1 g13437(.A0(n16778), .A1(n16773), .B0(n16775), .B1(n16779), .Y(n16780));
  AOI21X1 g13438(.A0(n16780), .A1(n14820), .B0(n16767), .Y(n16781));
  XOR2X1  g13439(.A(n16781), .B(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .Y(n16782));
  INVX1   g13440(.A(n16782), .Y(n16783));
  AOI21X1 g13441(.A0(n16732), .A1(n16697), .B0(n16735), .Y(n16784));
  INVX1   g13442(.A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .Y(n16785));
  NAND2X1 g13443(.A(n16781), .B(n16785), .Y(n16786));
  NOR2X1  g13444(.A(n16781), .B(n16785), .Y(n16787));
  INVX1   g13445(.A(n16787), .Y(n16788));
  AOI21X1 g13446(.A0(n16788), .A1(n16786), .B0(n16784), .Y(n16789));
  AOI21X1 g13447(.A0(n16784), .A1(n16783), .B0(n16789), .Y(n16790));
  NOR4X1  g13448(.A(n16637), .B(n16678), .C(n16698), .D(n16627), .Y(n16791));
  XOR2X1  g13449(.A(n16791), .B(n16785), .Y(n16792));
  AOI22X1 g13450(.A0(n16538), .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B0(P1_REIP_REG_6__SCAN_IN), .B1(n16527), .Y(n16793));
  OAI21X1 g13451(.A0(n16792), .A1(n18937), .B0(n16793), .Y(n16794));
  NAND2X1 g13452(.A(n16742), .B(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .Y(n16795));
  XOR2X1  g13453(.A(n16795), .B(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .Y(n16796));
  NOR2X1  g13454(.A(n16796), .B(n16545), .Y(n16797));
  AOI22X1 g13455(.A0(n16551), .A1(P1_EBX_REG_6__SCAN_IN), .B0(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B1(n16553), .Y(n16798));
  XOR2X1  g13456(.A(n16798), .B(n15054), .Y(n16799));
  INVX1   g13457(.A(n16688), .Y(n16800));
  NOR3X1  g13458(.A(n16746), .B(n16800), .C(n16687), .Y(n16801));
  XOR2X1  g13459(.A(n16801), .B(n16799), .Y(n16802));
  NOR2X1  g13460(.A(n16749), .B(n16698), .Y(n16803));
  XOR2X1  g13461(.A(n16803), .B(n16785), .Y(n16804));
  OAI22X1 g13462(.A0(n16802), .A1(n16558), .B0(n16636), .B1(n16804), .Y(n16805));
  NOR3X1  g13463(.A(n16805), .B(n16797), .C(n16794), .Y(n16806));
  OAI21X1 g13464(.A0(n16790), .A1(n16571), .B0(n16806), .Y(P1_U3025));
  INVX1   g13465(.A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .Y(n16808));
  NOR4X1  g13466(.A(n16710), .B(n16658), .C(n16620), .D(n16765), .Y(n16809));
  XOR2X1  g13467(.A(n16809), .B(n15381), .Y(n16810));
  NOR2X1  g13468(.A(n16810), .B(n15021), .Y(n16811));
  NOR2X1  g13469(.A(n16772), .B(n16769), .Y(n16812));
  INVX1   g13470(.A(n16812), .Y(n16813));
  AOI22X1 g13471(.A0(n14824), .A1(n15412), .B0(n14818), .B1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .Y(n16814));
  NAND2X1 g13472(.A(n15412), .B(n15401), .Y(n16815));
  XOR2X1  g13473(.A(n16815), .B(n16814), .Y(n16816));
  INVX1   g13474(.A(n16816), .Y(n16817));
  NAND4X1 g13475(.A(n16775), .B(n16813), .C(n16777), .D(n16817), .Y(n16818));
  INVX1   g13476(.A(n16818), .Y(n16819));
  NOR4X1  g13477(.A(n16722), .B(n16776), .C(n16723), .D(n16725), .Y(n16820));
  NAND2X1 g13478(.A(n16772), .B(n16769), .Y(n16821));
  NAND2X1 g13479(.A(n16821), .B(n16774), .Y(n16822));
  NOR3X1  g13480(.A(n16822), .B(n16820), .C(n16817), .Y(n16823));
  NOR2X1  g13481(.A(n16816), .B(n16821), .Y(n16824));
  NOR4X1  g13482(.A(n16823), .B(n16819), .C(n14821), .D(n16824), .Y(n16827));
  NOR2X1  g13483(.A(n16827), .B(n16811), .Y(n16828));
  AOI22X1 g13484(.A0(n16781), .A1(n16785), .B0(n16808), .B1(n16828), .Y(n16829));
  INVX1   g13485(.A(n16829), .Y(n16830));
  AOI21X1 g13486(.A0(n16788), .A1(n16784), .B0(n16830), .Y(n16831));
  OAI21X1 g13487(.A0(n16827), .A1(n16811), .B0(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .Y(n16832));
  AOI21X1 g13488(.A0(n16781), .A1(n16785), .B0(n16784), .Y(n16833));
  XOR2X1  g13489(.A(n16828), .B(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .Y(n16834));
  NAND2X1 g13490(.A(n16834), .B(n16788), .Y(n16835));
  NOR2X1  g13491(.A(n16835), .B(n16833), .Y(n16836));
  AOI21X1 g13492(.A0(n16832), .A1(n16831), .B0(n16836), .Y(n16837));
  NAND2X1 g13493(.A(n16837), .B(n16572), .Y(n16838));
  NAND2X1 g13494(.A(n16791), .B(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .Y(n16839));
  XOR2X1  g13495(.A(n16839), .B(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .Y(n16840));
  AOI22X1 g13496(.A0(n16538), .A1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B0(P1_REIP_REG_7__SCAN_IN), .B1(n16527), .Y(n16841));
  OAI21X1 g13497(.A0(n16840), .A1(n18937), .B0(n16841), .Y(n16842));
  INVX1   g13498(.A(n16742), .Y(n16843));
  NOR3X1  g13499(.A(n16843), .B(n16698), .C(n16785), .Y(n16844));
  XOR2X1  g13500(.A(n16844), .B(n16808), .Y(n16845));
  NOR2X1  g13501(.A(n16845), .B(n16545), .Y(n16846));
  AOI22X1 g13502(.A0(n16551), .A1(P1_EBX_REG_7__SCAN_IN), .B0(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B1(n16553), .Y(n16847));
  XOR2X1  g13503(.A(n16847), .B(n15054), .Y(n16848));
  NOR4X1  g13504(.A(n16746), .B(n16800), .C(n16687), .D(n16799), .Y(n16849));
  XOR2X1  g13505(.A(n16849), .B(n16848), .Y(n16850));
  NOR3X1  g13506(.A(n16749), .B(n16698), .C(n16785), .Y(n16851));
  XOR2X1  g13507(.A(n16851), .B(n16808), .Y(n16852));
  OAI22X1 g13508(.A0(n16850), .A1(n16558), .B0(n16636), .B1(n16852), .Y(n16853));
  NOR3X1  g13509(.A(n16853), .B(n16846), .C(n16842), .Y(n16854));
  NAND2X1 g13510(.A(n16854), .B(n16838), .Y(P1_U3024));
  INVX1   g13511(.A(n16832), .Y(n16856));
  NOR2X1  g13512(.A(n16856), .B(n16831), .Y(n16857));
  INVX1   g13513(.A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .Y(n16858));
  NOR4X1  g13514(.A(n15381), .B(n14770), .C(n14707), .D(n16765), .Y(n16859));
  AOI22X1 g13515(.A0(n14704), .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B0(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(n15355), .Y(n16862));
  AOI22X1 g13516(.A0(n15359), .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B0(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(n14673), .Y(n16865));
  AOI22X1 g13517(.A0(n14674), .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B0(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(n15361), .Y(n16868));
  AOI22X1 g13518(.A0(n15365), .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B0(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(n15362), .Y(n16871));
  NAND4X1 g13519(.A(n16868), .B(n16865), .C(n16862), .D(n16871), .Y(n16872));
  AOI22X1 g13520(.A0(n14682), .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B0(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(n14680), .Y(n16875));
  AOI22X1 g13521(.A0(n15372), .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B0(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(n14907), .Y(n16878));
  AOI22X1 g13522(.A0(n14703), .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B0(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(n14671), .Y(n16881));
  AOI22X1 g13523(.A0(n15378), .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B0(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(n15375), .Y(n16884));
  NAND4X1 g13524(.A(n16881), .B(n16878), .C(n16875), .D(n16884), .Y(n16885));
  AOI21X1 g13525(.A0(n14746), .A1(n14806), .B0(n14650), .Y(n16886));
  OAI21X1 g13526(.A0(n16885), .A1(n16872), .B0(n16886), .Y(n16887));
  XOR2X1  g13527(.A(n16887), .B(n15382), .Y(n16888));
  INVX1   g13528(.A(n16774), .Y(n16889));
  AOI22X1 g13529(.A0(n16814), .A1(n16815), .B0(n16772), .B1(n16769), .Y(n16890));
  INVX1   g13530(.A(n16890), .Y(n16891));
  NOR3X1  g13531(.A(n16891), .B(n16889), .C(n16720), .Y(n16892));
  INVX1   g13532(.A(n16892), .Y(n16893));
  NOR2X1  g13533(.A(n16815), .B(n16814), .Y(n16894));
  NOR2X1  g13534(.A(n16891), .B(n16777), .Y(n16895));
  NOR2X1  g13535(.A(n16891), .B(n16813), .Y(n16896));
  NOR3X1  g13536(.A(n16891), .B(n16889), .C(n16724), .Y(n16897));
  NOR4X1  g13537(.A(n16896), .B(n16895), .C(n16894), .D(n16897), .Y(n16898));
  OAI21X1 g13538(.A0(n16893), .A1(n16672), .B0(n16898), .Y(n16899));
  INVX1   g13539(.A(n16899), .Y(n16900));
  XOR2X1  g13540(.A(n16900), .B(n16888), .Y(n16901));
  AOI22X1 g13541(.A0(n16859), .A1(n16754), .B0(n14820), .B1(n16901), .Y(n16902));
  XOR2X1  g13542(.A(n16902), .B(n16858), .Y(n16903));
  XOR2X1  g13543(.A(n16903), .B(n16857), .Y(n16904));
  NAND3X1 g13544(.A(n16791), .B(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .C(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .Y(n16905));
  XOR2X1  g13545(.A(n16905), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .Y(n16906));
  AOI22X1 g13546(.A0(n16538), .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B0(P1_REIP_REG_8__SCAN_IN), .B1(n16527), .Y(n16907));
  OAI21X1 g13547(.A0(n16906), .A1(n18937), .B0(n16907), .Y(n16908));
  NAND4X1 g13548(.A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .B(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .C(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .D(n16742), .Y(n16909));
  XOR2X1  g13549(.A(n16909), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .Y(n16910));
  NOR2X1  g13550(.A(n16910), .B(n16545), .Y(n16911));
  AOI22X1 g13551(.A0(n16551), .A1(P1_EBX_REG_8__SCAN_IN), .B0(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(n16553), .Y(n16912));
  XOR2X1  g13552(.A(n16912), .B(n15054), .Y(n16913));
  INVX1   g13553(.A(n16913), .Y(n16914));
  NOR2X1  g13554(.A(n16848), .B(n16799), .Y(n16915));
  NAND2X1 g13555(.A(n16915), .B(n16801), .Y(n16916));
  XOR2X1  g13556(.A(n16916), .B(n16914), .Y(n16917));
  NOR4X1  g13557(.A(n16698), .B(n16785), .C(n16808), .D(n16749), .Y(n16918));
  XOR2X1  g13558(.A(n16918), .B(n16858), .Y(n16919));
  OAI22X1 g13559(.A0(n16917), .A1(n16558), .B0(n16636), .B1(n16919), .Y(n16920));
  NOR3X1  g13560(.A(n16920), .B(n16911), .C(n16908), .Y(n16921));
  OAI21X1 g13561(.A0(n16904), .A1(n16571), .B0(n16921), .Y(P1_U3023));
  NOR2X1  g13562(.A(n16900), .B(n16888), .Y(n16923));
  AOI22X1 g13563(.A0(n14704), .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B0(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(n15355), .Y(n16924));
  AOI22X1 g13564(.A0(n15359), .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B0(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(n14673), .Y(n16925));
  AOI22X1 g13565(.A0(n14674), .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B0(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(n15361), .Y(n16926));
  AOI22X1 g13566(.A0(n15365), .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B0(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(n15362), .Y(n16927));
  NAND4X1 g13567(.A(n16926), .B(n16925), .C(n16924), .D(n16927), .Y(n16928));
  AOI22X1 g13568(.A0(n14682), .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B0(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(n14680), .Y(n16929));
  AOI22X1 g13569(.A0(n15372), .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B0(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(n14907), .Y(n16930));
  AOI22X1 g13570(.A0(n14703), .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B0(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(n14671), .Y(n16931));
  AOI22X1 g13571(.A0(n15378), .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B0(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(n15375), .Y(n16932));
  NAND4X1 g13572(.A(n16931), .B(n16930), .C(n16929), .D(n16932), .Y(n16933));
  OAI21X1 g13573(.A0(n16933), .A1(n16928), .B0(n16886), .Y(n16934));
  XOR2X1  g13574(.A(n16934), .B(n15382), .Y(n16935));
  XOR2X1  g13575(.A(n16935), .B(n16923), .Y(n16936));
  NOR2X1  g13576(.A(n16936), .B(n14821), .Y(n16937));
  XOR2X1  g13577(.A(n16937), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .Y(n16938));
  INVX1   g13578(.A(n16902), .Y(n16939));
  OAI21X1 g13579(.A0(n16939), .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B0(n16829), .Y(n16940));
  AOI21X1 g13580(.A0(n16788), .A1(n16784), .B0(n16940), .Y(n16941));
  AOI21X1 g13581(.A0(n16902), .A1(n16858), .B0(n16832), .Y(n16942));
  NOR2X1  g13582(.A(n16902), .B(n16858), .Y(n16943));
  NOR3X1  g13583(.A(n16943), .B(n16942), .C(n16941), .Y(n16944));
  XOR2X1  g13584(.A(n16944), .B(n16938), .Y(n16945));
  NAND4X1 g13585(.A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .D(n16791), .Y(n16946));
  XOR2X1  g13586(.A(n16946), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .Y(n16947));
  AOI22X1 g13587(.A0(n16538), .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B0(P1_REIP_REG_9__SCAN_IN), .B1(n16527), .Y(n16948));
  OAI21X1 g13588(.A0(n16947), .A1(n18937), .B0(n16948), .Y(n16949));
  NAND3X1 g13589(.A(n16844), .B(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .Y(n16950));
  XOR2X1  g13590(.A(n16950), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .Y(n16951));
  NOR2X1  g13591(.A(n16951), .B(n16545), .Y(n16952));
  AOI22X1 g13592(.A0(n16551), .A1(P1_EBX_REG_9__SCAN_IN), .B0(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B1(n16553), .Y(n16953));
  XOR2X1  g13593(.A(n16953), .B(n15054), .Y(n16954));
  NOR2X1  g13594(.A(n16916), .B(n16913), .Y(n16955));
  XOR2X1  g13595(.A(n16955), .B(n16954), .Y(n16956));
  NAND2X1 g13596(.A(n16918), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .Y(n16957));
  XOR2X1  g13597(.A(n16957), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .Y(n16958));
  OAI22X1 g13598(.A0(n16956), .A1(n16558), .B0(n16636), .B1(n16958), .Y(n16959));
  NOR3X1  g13599(.A(n16959), .B(n16952), .C(n16949), .Y(n16960));
  OAI21X1 g13600(.A0(n16945), .A1(n16571), .B0(n16960), .Y(P1_U3022));
  INVX1   g13601(.A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .Y(n16962));
  NOR3X1  g13602(.A(n16936), .B(n14821), .C(n16962), .Y(n16963));
  INVX1   g13603(.A(n16963), .Y(n16964));
  NOR2X1  g13604(.A(n16937), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .Y(n16965));
  OAI21X1 g13605(.A0(n16944), .A1(n16965), .B0(n16964), .Y(n16966));
  INVX1   g13606(.A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .Y(n16967));
  AOI22X1 g13607(.A0(n14704), .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B0(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(n15355), .Y(n16968));
  AOI22X1 g13608(.A0(n15359), .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B0(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(n14673), .Y(n16969));
  AOI22X1 g13609(.A0(n14674), .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B0(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(n15361), .Y(n16970));
  AOI22X1 g13610(.A0(n15365), .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B0(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(n15362), .Y(n16971));
  NAND4X1 g13611(.A(n16970), .B(n16969), .C(n16968), .D(n16971), .Y(n16972));
  AOI22X1 g13612(.A0(n14682), .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B0(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(n14680), .Y(n16973));
  AOI22X1 g13613(.A0(n15372), .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B0(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(n14907), .Y(n16974));
  AOI22X1 g13614(.A0(n14703), .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B0(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(n14671), .Y(n16975));
  AOI22X1 g13615(.A0(n15378), .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B0(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(n15375), .Y(n16976));
  NAND4X1 g13616(.A(n16975), .B(n16974), .C(n16973), .D(n16976), .Y(n16977));
  OAI21X1 g13617(.A0(n16977), .A1(n16972), .B0(n16886), .Y(n16978));
  XOR2X1  g13618(.A(n16978), .B(n15382), .Y(n16979));
  INVX1   g13619(.A(n16979), .Y(n16980));
  NOR2X1  g13620(.A(n16935), .B(n16888), .Y(n16981));
  NAND2X1 g13621(.A(n16981), .B(n16899), .Y(n16982));
  XOR2X1  g13622(.A(n16982), .B(n16980), .Y(n16983));
  NOR2X1  g13623(.A(n16983), .B(n14821), .Y(n16984));
  XOR2X1  g13624(.A(n16984), .B(n16967), .Y(n16985));
  NOR2X1  g13625(.A(n16985), .B(n16966), .Y(n16986));
  AOI21X1 g13626(.A0(n16985), .A1(n16966), .B0(n16986), .Y(n16988));
  NOR2X1  g13627(.A(n16946), .B(n16962), .Y(n16989));
  XOR2X1  g13628(.A(n16989), .B(n16967), .Y(n16990));
  AOI22X1 g13629(.A0(n16538), .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B0(P1_REIP_REG_10__SCAN_IN), .B1(n16527), .Y(n16991));
  OAI21X1 g13630(.A0(n16990), .A1(n18937), .B0(n16991), .Y(n16992));
  NAND4X1 g13631(.A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .C(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .D(n16844), .Y(n16993));
  XOR2X1  g13632(.A(n16993), .B(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .Y(n16994));
  NOR2X1  g13633(.A(n16994), .B(n16545), .Y(n16995));
  AOI22X1 g13634(.A0(n16551), .A1(P1_EBX_REG_10__SCAN_IN), .B0(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B1(n16553), .Y(n16996));
  XOR2X1  g13635(.A(n16996), .B(n15054), .Y(n16997));
  NOR3X1  g13636(.A(n16954), .B(n16916), .C(n16913), .Y(n16998));
  XOR2X1  g13637(.A(n16998), .B(n16997), .Y(n16999));
  NAND3X1 g13638(.A(n16918), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .C(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .Y(n17000));
  XOR2X1  g13639(.A(n17000), .B(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .Y(n17001));
  OAI22X1 g13640(.A0(n16999), .A1(n16558), .B0(n16636), .B1(n17001), .Y(n17002));
  NOR3X1  g13641(.A(n17002), .B(n16995), .C(n16992), .Y(n17003));
  OAI21X1 g13642(.A0(n16988), .A1(n16571), .B0(n17003), .Y(P1_U3021));
  NOR3X1  g13643(.A(n16983), .B(n14821), .C(n16967), .Y(n17005));
  NOR4X1  g13644(.A(n16943), .B(n16942), .C(n16963), .D(n17005), .Y(n17006));
  INVX1   g13645(.A(n17006), .Y(n17007));
  NOR2X1  g13646(.A(n16984), .B(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .Y(n17008));
  NOR2X1  g13647(.A(n17008), .B(n16965), .Y(n17009));
  AOI22X1 g13648(.A0(n14704), .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B0(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(n15355), .Y(n17010));
  AOI22X1 g13649(.A0(n15359), .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B0(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(n14673), .Y(n17011));
  AOI22X1 g13650(.A0(n14674), .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B0(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(n15361), .Y(n17012));
  AOI22X1 g13651(.A0(n15365), .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B0(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(n15362), .Y(n17013));
  NAND4X1 g13652(.A(n17012), .B(n17011), .C(n17010), .D(n17013), .Y(n17014));
  AOI22X1 g13653(.A0(n14682), .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B0(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(n14680), .Y(n17015));
  AOI22X1 g13654(.A0(n15372), .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B0(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(n14907), .Y(n17016));
  AOI22X1 g13655(.A0(n14703), .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B0(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(n14671), .Y(n17017));
  AOI22X1 g13656(.A0(n15378), .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B0(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(n15375), .Y(n17018));
  NAND4X1 g13657(.A(n17017), .B(n17016), .C(n17015), .D(n17018), .Y(n17019));
  OAI21X1 g13658(.A0(n17019), .A1(n17014), .B0(n16886), .Y(n17020));
  XOR2X1  g13659(.A(n17020), .B(n15382), .Y(n17021));
  NOR4X1  g13660(.A(n16935), .B(n16900), .C(n16888), .D(n16979), .Y(n17022));
  XOR2X1  g13661(.A(n17022), .B(n17021), .Y(n17023));
  NOR2X1  g13662(.A(n17023), .B(n14821), .Y(n17024));
  OAI22X1 g13663(.A0(n17009), .A1(n17005), .B0(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B1(n17024), .Y(n17025));
  INVX1   g13664(.A(n17025), .Y(n17026));
  OAI21X1 g13665(.A0(n17007), .A1(n16941), .B0(n17026), .Y(n17027));
  INVX1   g13666(.A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .Y(n17028));
  NOR3X1  g13667(.A(n17023), .B(n14821), .C(n17028), .Y(n17029));
  INVX1   g13668(.A(n16966), .Y(n17030));
  NOR2X1  g13669(.A(n17008), .B(n17030), .Y(n17031));
  INVX1   g13670(.A(n17024), .Y(n17032));
  AOI21X1 g13671(.A0(n17032), .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B0(n17005), .Y(n17033));
  OAI21X1 g13672(.A0(n17032), .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B0(n17033), .Y(n17034));
  OAI22X1 g13673(.A0(n17031), .A1(n17034), .B0(n17029), .B1(n17027), .Y(n17035));
  NOR3X1  g13674(.A(n16946), .B(n16962), .C(n16967), .Y(n17036));
  XOR2X1  g13675(.A(n17036), .B(n17028), .Y(n17037));
  AOI22X1 g13676(.A0(n16538), .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B0(P1_REIP_REG_11__SCAN_IN), .B1(n16527), .Y(n17038));
  OAI21X1 g13677(.A0(n17037), .A1(n18937), .B0(n17038), .Y(n17039));
  NOR3X1  g13678(.A(n16950), .B(n16962), .C(n16967), .Y(n17040));
  XOR2X1  g13679(.A(n17040), .B(n17028), .Y(n17041));
  NOR2X1  g13680(.A(n17041), .B(n16545), .Y(n17042));
  AOI22X1 g13681(.A0(n16551), .A1(P1_EBX_REG_11__SCAN_IN), .B0(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B1(n16553), .Y(n17043));
  XOR2X1  g13682(.A(n17043), .B(n15054), .Y(n17044));
  NOR4X1  g13683(.A(n16954), .B(n16916), .C(n16913), .D(n16997), .Y(n17045));
  XOR2X1  g13684(.A(n17045), .B(n17044), .Y(n17046));
  NAND4X1 g13685(.A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .D(n16918), .Y(n17047));
  XOR2X1  g13686(.A(n17047), .B(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .Y(n17048));
  OAI22X1 g13687(.A0(n17046), .A1(n16558), .B0(n16636), .B1(n17048), .Y(n17049));
  NOR3X1  g13688(.A(n17049), .B(n17042), .C(n17039), .Y(n17050));
  OAI21X1 g13689(.A0(n17035), .A1(n16571), .B0(n17050), .Y(P1_U3020));
  INVX1   g13690(.A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .Y(n17052));
  AOI22X1 g13691(.A0(n14704), .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B0(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(n15355), .Y(n17053));
  AOI22X1 g13692(.A0(n15359), .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B0(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(n14673), .Y(n17054));
  AOI22X1 g13693(.A0(n14674), .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B0(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(n15361), .Y(n17055));
  AOI22X1 g13694(.A0(n15365), .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B0(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(n15362), .Y(n17056));
  NAND4X1 g13695(.A(n17055), .B(n17054), .C(n17053), .D(n17056), .Y(n17057));
  AOI22X1 g13696(.A0(n14682), .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B0(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(n14680), .Y(n17058));
  AOI22X1 g13697(.A0(n15372), .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B0(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(n14907), .Y(n17059));
  AOI22X1 g13698(.A0(n14703), .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B0(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(n14671), .Y(n17060));
  AOI22X1 g13699(.A0(n15378), .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B0(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(n15375), .Y(n17061));
  NAND4X1 g13700(.A(n17060), .B(n17059), .C(n17058), .D(n17061), .Y(n17062));
  OAI21X1 g13701(.A0(n17062), .A1(n17057), .B0(n16886), .Y(n17063));
  XOR2X1  g13702(.A(n17063), .B(n15382), .Y(n17064));
  NOR4X1  g13703(.A(n16979), .B(n16935), .C(n16888), .D(n17021), .Y(n17065));
  INVX1   g13704(.A(n17065), .Y(n17066));
  NOR2X1  g13705(.A(n17066), .B(n16900), .Y(n17067));
  XOR2X1  g13706(.A(n17067), .B(n17064), .Y(n17068));
  NOR3X1  g13707(.A(n17068), .B(n14821), .C(n17052), .Y(n17069));
  INVX1   g13708(.A(n17069), .Y(n17070));
  INVX1   g13709(.A(n17068), .Y(n17071));
  AOI21X1 g13710(.A0(n17071), .A1(n14820), .B0(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .Y(n17072));
  INVX1   g13711(.A(n17072), .Y(n17073));
  NAND2X1 g13712(.A(n17073), .B(n17070), .Y(n17074));
  INVX1   g13713(.A(n17029), .Y(n17075));
  NAND2X1 g13714(.A(n17075), .B(n17027), .Y(n17076));
  XOR2X1  g13715(.A(n17076), .B(n17074), .Y(n17077));
  NOR4X1  g13716(.A(n16962), .B(n16967), .C(n17028), .D(n16946), .Y(n17078));
  XOR2X1  g13717(.A(n17078), .B(n17052), .Y(n17079));
  AOI22X1 g13718(.A0(n16538), .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .B0(P1_REIP_REG_12__SCAN_IN), .B1(n16527), .Y(n17080));
  OAI21X1 g13719(.A0(n17079), .A1(n18937), .B0(n17080), .Y(n17081));
  NOR4X1  g13720(.A(n16962), .B(n16967), .C(n17028), .D(n16950), .Y(n17082));
  XOR2X1  g13721(.A(n17082), .B(n17052), .Y(n17083));
  NOR2X1  g13722(.A(n17083), .B(n16545), .Y(n17084));
  AOI22X1 g13723(.A0(n16551), .A1(P1_EBX_REG_12__SCAN_IN), .B0(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .B1(n16553), .Y(n17085));
  XOR2X1  g13724(.A(n17085), .B(n15054), .Y(n17086));
  INVX1   g13725(.A(n17086), .Y(n17087));
  NOR2X1  g13726(.A(n17044), .B(n16997), .Y(n17088));
  NAND2X1 g13727(.A(n17088), .B(n16998), .Y(n17089));
  XOR2X1  g13728(.A(n17089), .B(n17087), .Y(n17090));
  NOR2X1  g13729(.A(n17047), .B(n17028), .Y(n17091));
  XOR2X1  g13730(.A(n17091), .B(n17052), .Y(n17092));
  OAI22X1 g13731(.A0(n17090), .A1(n16558), .B0(n16636), .B1(n17092), .Y(n17093));
  NOR3X1  g13732(.A(n17093), .B(n17084), .C(n17081), .Y(n17094));
  OAI21X1 g13733(.A0(n17077), .A1(n16571), .B0(n17094), .Y(P1_U3019));
  AOI21X1 g13734(.A0(n17076), .A1(n17073), .B0(n17069), .Y(n17096));
  AOI22X1 g13735(.A0(n14704), .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B0(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(n15355), .Y(n17097));
  AOI22X1 g13736(.A0(n15359), .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B0(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(n14673), .Y(n17098));
  AOI22X1 g13737(.A0(n14674), .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B0(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(n15361), .Y(n17099));
  AOI22X1 g13738(.A0(n15365), .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B0(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(n15362), .Y(n17100));
  NAND4X1 g13739(.A(n17099), .B(n17098), .C(n17097), .D(n17100), .Y(n17101));
  AOI22X1 g13740(.A0(n14682), .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B0(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(n14680), .Y(n17102));
  AOI22X1 g13741(.A0(n15372), .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B0(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(n14907), .Y(n17103));
  AOI22X1 g13742(.A0(n14703), .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B0(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(n14671), .Y(n17104));
  AOI22X1 g13743(.A0(n15378), .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B0(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(n15375), .Y(n17105));
  NAND4X1 g13744(.A(n17104), .B(n17103), .C(n17102), .D(n17105), .Y(n17106));
  OAI21X1 g13745(.A0(n17106), .A1(n17101), .B0(n16886), .Y(n17107));
  XOR2X1  g13746(.A(n17107), .B(n15382), .Y(n17108));
  NOR3X1  g13747(.A(n17066), .B(n17064), .C(n16900), .Y(n17109));
  XOR2X1  g13748(.A(n17109), .B(n17108), .Y(n17110));
  NOR2X1  g13749(.A(n17110), .B(n14821), .Y(n17111));
  XOR2X1  g13750(.A(n17111), .B(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .Y(n17112));
  NOR2X1  g13751(.A(n17112), .B(n17096), .Y(n17114));
  AOI21X1 g13752(.A0(n17112), .A1(n17096), .B0(n17114), .Y(n17115));
  AOI22X1 g13753(.A0(n16551), .A1(P1_EBX_REG_13__SCAN_IN), .B0(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B1(n16553), .Y(n17116));
  XOR2X1  g13754(.A(n17116), .B(n15054), .Y(n17117));
  NOR2X1  g13755(.A(n17089), .B(n17086), .Y(n17118));
  XOR2X1  g13756(.A(n17118), .B(n17117), .Y(n17119));
  AOI22X1 g13757(.A0(n16538), .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B0(P1_REIP_REG_13__SCAN_IN), .B1(n16527), .Y(n17120));
  OAI21X1 g13758(.A0(n17119), .A1(n16558), .B0(n17120), .Y(n17121));
  NAND3X1 g13759(.A(n17040), .B(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .C(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .Y(n17122));
  XOR2X1  g13760(.A(n17122), .B(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .Y(n17123));
  NOR2X1  g13761(.A(n17123), .B(n16545), .Y(n17124));
  INVX1   g13762(.A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .Y(n17125));
  NOR3X1  g13763(.A(n17047), .B(n17028), .C(n17052), .Y(n17126));
  XOR2X1  g13764(.A(n17126), .B(n17125), .Y(n17127));
  NAND2X1 g13765(.A(n17078), .B(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .Y(n17128));
  XOR2X1  g13766(.A(n17128), .B(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .Y(n17129));
  OAI22X1 g13767(.A0(n17127), .A1(n16636), .B0(n18937), .B1(n17129), .Y(n17130));
  NOR3X1  g13768(.A(n17130), .B(n17124), .C(n17121), .Y(n17131));
  OAI21X1 g13769(.A0(n17115), .A1(n16571), .B0(n17131), .Y(P1_U3018));
  NOR2X1  g13770(.A(n17111), .B(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .Y(n17133));
  NOR3X1  g13771(.A(n17110), .B(n14821), .C(n17125), .Y(n17134));
  INVX1   g13772(.A(n17134), .Y(n17135));
  OAI21X1 g13773(.A0(n17133), .A1(n17096), .B0(n17135), .Y(n17136));
  INVX1   g13774(.A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .Y(n17137));
  AOI22X1 g13775(.A0(n14704), .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B0(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(n15355), .Y(n17138));
  AOI22X1 g13776(.A0(n15359), .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B0(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(n14673), .Y(n17139));
  AOI22X1 g13777(.A0(n14674), .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B0(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(n15361), .Y(n17140));
  AOI22X1 g13778(.A0(n15365), .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B0(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(n15362), .Y(n17141));
  NAND4X1 g13779(.A(n17140), .B(n17139), .C(n17138), .D(n17141), .Y(n17142));
  AOI22X1 g13780(.A0(n14682), .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B0(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(n14680), .Y(n17143));
  AOI22X1 g13781(.A0(n15372), .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B0(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(n14907), .Y(n17144));
  AOI22X1 g13782(.A0(n14703), .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B0(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(n14671), .Y(n17145));
  AOI22X1 g13783(.A0(n15378), .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B0(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(n15375), .Y(n17146));
  NAND4X1 g13784(.A(n17145), .B(n17144), .C(n17143), .D(n17146), .Y(n17147));
  OAI21X1 g13785(.A0(n17147), .A1(n17142), .B0(n16886), .Y(n17148));
  XOR2X1  g13786(.A(n17148), .B(n15382), .Y(n17149));
  INVX1   g13787(.A(n17149), .Y(n17150));
  NOR2X1  g13788(.A(n17108), .B(n17064), .Y(n17151));
  NAND3X1 g13789(.A(n17151), .B(n17065), .C(n16899), .Y(n17152));
  XOR2X1  g13790(.A(n17152), .B(n17150), .Y(n17153));
  NOR2X1  g13791(.A(n17153), .B(n14821), .Y(n17154));
  XOR2X1  g13792(.A(n17154), .B(n17137), .Y(n17155));
  NOR2X1  g13793(.A(n17136), .B(n17155), .Y(n17156));
  AOI21X1 g13794(.A0(n17155), .A1(n17136), .B0(n17156), .Y(n17158));
  AOI22X1 g13795(.A0(n16551), .A1(P1_EBX_REG_14__SCAN_IN), .B0(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B1(n16553), .Y(n17159));
  XOR2X1  g13796(.A(n17159), .B(n15054), .Y(n17160));
  NOR3X1  g13797(.A(n17117), .B(n17089), .C(n17086), .Y(n17161));
  XOR2X1  g13798(.A(n17161), .B(n17160), .Y(n17162));
  AOI22X1 g13799(.A0(n16538), .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B0(P1_REIP_REG_14__SCAN_IN), .B1(n16527), .Y(n17163));
  OAI21X1 g13800(.A0(n17162), .A1(n16558), .B0(n17163), .Y(n17164));
  NAND4X1 g13801(.A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .C(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .D(n17040), .Y(n17165));
  XOR2X1  g13802(.A(n17165), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .Y(n17166));
  NOR2X1  g13803(.A(n17166), .B(n16545), .Y(n17167));
  NOR4X1  g13804(.A(n17028), .B(n17052), .C(n17125), .D(n17047), .Y(n17168));
  XOR2X1  g13805(.A(n17168), .B(n17137), .Y(n17169));
  NAND3X1 g13806(.A(n17078), .B(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .C(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .Y(n17170));
  XOR2X1  g13807(.A(n17170), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .Y(n17171));
  OAI22X1 g13808(.A0(n17169), .A1(n16636), .B0(n18937), .B1(n17171), .Y(n17172));
  NOR3X1  g13809(.A(n17172), .B(n17167), .C(n17164), .Y(n17173));
  OAI21X1 g13810(.A0(n17158), .A1(n16571), .B0(n17173), .Y(P1_U3017));
  NOR3X1  g13811(.A(n17153), .B(n14821), .C(n17137), .Y(n17175));
  AOI22X1 g13812(.A0(n14704), .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B0(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(n15355), .Y(n17176));
  AOI22X1 g13813(.A0(n15359), .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B0(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(n14673), .Y(n17177));
  AOI22X1 g13814(.A0(n14674), .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B0(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(n15361), .Y(n17178));
  AOI22X1 g13815(.A0(n15365), .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B0(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(n15362), .Y(n17179));
  NAND4X1 g13816(.A(n17178), .B(n17177), .C(n17176), .D(n17179), .Y(n17180));
  AOI22X1 g13817(.A0(n14682), .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B0(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(n14680), .Y(n17181));
  AOI22X1 g13818(.A0(n15372), .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B0(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(n14907), .Y(n17182));
  AOI22X1 g13819(.A0(n14703), .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B0(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(n14671), .Y(n17183));
  AOI22X1 g13820(.A0(n15378), .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B0(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(n15375), .Y(n17184));
  NAND4X1 g13821(.A(n17183), .B(n17182), .C(n17181), .D(n17184), .Y(n17185));
  OAI21X1 g13822(.A0(n17185), .A1(n17180), .B0(n16886), .Y(n17186));
  XOR2X1  g13823(.A(n17186), .B(n15382), .Y(n17187));
  NOR2X1  g13824(.A(n17152), .B(n17149), .Y(n17188));
  XOR2X1  g13825(.A(n17188), .B(n17187), .Y(n17189));
  NOR2X1  g13826(.A(n17189), .B(n14821), .Y(n17190));
  OAI22X1 g13827(.A0(n17154), .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B0(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B1(n17190), .Y(n17191));
  AOI21X1 g13828(.A0(n17190), .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B0(n17191), .Y(n17192));
  OAI21X1 g13829(.A0(n17175), .A1(n17136), .B0(n17192), .Y(n17193));
  OAI21X1 g13830(.A0(n17154), .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B0(n17136), .Y(n17194));
  INVX1   g13831(.A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .Y(n17195));
  INVX1   g13832(.A(n17175), .Y(n17196));
  OAI21X1 g13833(.A0(n17190), .A1(n17195), .B0(n17196), .Y(n17197));
  AOI21X1 g13834(.A0(n17190), .A1(n17195), .B0(n17197), .Y(n17198));
  NAND2X1 g13835(.A(n17198), .B(n17194), .Y(n17199));
  NAND2X1 g13836(.A(n17199), .B(n17193), .Y(n17200));
  AOI22X1 g13837(.A0(n16551), .A1(P1_EBX_REG_15__SCAN_IN), .B0(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B1(n16553), .Y(n17201));
  XOR2X1  g13838(.A(n17201), .B(n15054), .Y(n17202));
  NOR4X1  g13839(.A(n17117), .B(n17089), .C(n17086), .D(n17160), .Y(n17203));
  XOR2X1  g13840(.A(n17203), .B(n17202), .Y(n17204));
  AOI22X1 g13841(.A0(n16538), .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B0(P1_REIP_REG_15__SCAN_IN), .B1(n16527), .Y(n17205));
  OAI21X1 g13842(.A0(n17204), .A1(n16558), .B0(n17205), .Y(n17206));
  NOR3X1  g13843(.A(n17122), .B(n17125), .C(n17137), .Y(n17207));
  XOR2X1  g13844(.A(n17207), .B(n17195), .Y(n17208));
  NOR2X1  g13845(.A(n17208), .B(n16545), .Y(n17209));
  NAND2X1 g13846(.A(n17168), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .Y(n17210));
  XOR2X1  g13847(.A(n17210), .B(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .Y(n17211));
  NAND4X1 g13848(.A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .B(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .C(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .D(n17078), .Y(n17212));
  XOR2X1  g13849(.A(n17212), .B(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .Y(n17213));
  OAI22X1 g13850(.A0(n17211), .A1(n16636), .B0(n18937), .B1(n17213), .Y(n17214));
  NOR3X1  g13851(.A(n17214), .B(n17209), .C(n17206), .Y(n17215));
  OAI21X1 g13852(.A0(n17200), .A1(n16571), .B0(n17215), .Y(P1_U3016));
  NOR2X1  g13853(.A(n17154), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .Y(n17217));
  OAI22X1 g13854(.A0(n17217), .A1(n17195), .B0(n14821), .B1(n17189), .Y(n17218));
  NOR3X1  g13855(.A(n17217), .B(n17133), .C(n17072), .Y(n17219));
  NAND2X1 g13856(.A(n17219), .B(n17218), .Y(n17220));
  AOI21X1 g13857(.A0(n17075), .A1(n17027), .B0(n17220), .Y(n17221));
  OAI21X1 g13858(.A0(n17111), .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B0(n17069), .Y(n17222));
  NOR2X1  g13859(.A(n17175), .B(n17134), .Y(n17223));
  AOI21X1 g13860(.A0(n17223), .A1(n17222), .B0(n17191), .Y(n17224));
  AOI21X1 g13861(.A0(n17190), .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B0(n17224), .Y(n17225));
  INVX1   g13862(.A(n17225), .Y(n17226));
  NOR2X1  g13863(.A(n17226), .B(n17221), .Y(n17227));
  NOR4X1  g13864(.A(n17149), .B(n17108), .C(n17064), .D(n17187), .Y(n17228));
  NAND3X1 g13865(.A(n17228), .B(n17065), .C(n16899), .Y(n17229));
  XOR2X1  g13866(.A(n17229), .B(n15382), .Y(n17230));
  NOR2X1  g13867(.A(n17230), .B(n14821), .Y(n17231));
  XOR2X1  g13868(.A(n17231), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .Y(n17232));
  XOR2X1  g13869(.A(n17232), .B(n17227), .Y(n17233));
  AOI22X1 g13870(.A0(n16551), .A1(P1_EBX_REG_16__SCAN_IN), .B0(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B1(n16553), .Y(n17234));
  XOR2X1  g13871(.A(n17234), .B(n15054), .Y(n17235));
  INVX1   g13872(.A(n17235), .Y(n17236));
  NOR2X1  g13873(.A(n17202), .B(n17160), .Y(n17237));
  NAND2X1 g13874(.A(n17237), .B(n17161), .Y(n17238));
  XOR2X1  g13875(.A(n17238), .B(n17236), .Y(n17239));
  AOI22X1 g13876(.A0(n16538), .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B0(P1_REIP_REG_16__SCAN_IN), .B1(n16527), .Y(n17240));
  OAI21X1 g13877(.A0(n17239), .A1(n16558), .B0(n17240), .Y(n17241));
  INVX1   g13878(.A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .Y(n17242));
  NOR4X1  g13879(.A(n17125), .B(n17137), .C(n17195), .D(n17122), .Y(n17243));
  XOR2X1  g13880(.A(n17243), .B(n17242), .Y(n17244));
  NOR2X1  g13881(.A(n17244), .B(n16545), .Y(n17245));
  NAND3X1 g13882(.A(n17168), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .C(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .Y(n17246));
  XOR2X1  g13883(.A(n17246), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .Y(n17247));
  NOR2X1  g13884(.A(n17212), .B(n17195), .Y(n17248));
  XOR2X1  g13885(.A(n17248), .B(n17242), .Y(n17249));
  OAI22X1 g13886(.A0(n17247), .A1(n16636), .B0(n18937), .B1(n17249), .Y(n17250));
  NOR3X1  g13887(.A(n17250), .B(n17245), .C(n17241), .Y(n17251));
  OAI21X1 g13888(.A0(n17233), .A1(n16571), .B0(n17251), .Y(P1_U3015));
  INVX1   g13889(.A(n17231), .Y(n17253));
  OAI22X1 g13890(.A0(n17226), .A1(n17221), .B0(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B1(n17231), .Y(n17254));
  OAI21X1 g13891(.A0(n17253), .A1(n17242), .B0(n17254), .Y(n17255));
  INVX1   g13892(.A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .Y(n17256));
  INVX1   g13893(.A(n17229), .Y(n17257));
  XOR2X1  g13894(.A(n17231), .B(n17256), .Y(n17259));
  XOR2X1  g13895(.A(n17259), .B(n17255), .Y(n17260));
  AOI22X1 g13896(.A0(n16551), .A1(P1_EBX_REG_17__SCAN_IN), .B0(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B1(n16553), .Y(n17261));
  XOR2X1  g13897(.A(n17261), .B(n15054), .Y(n17262));
  NOR2X1  g13898(.A(n17238), .B(n17235), .Y(n17263));
  XOR2X1  g13899(.A(n17263), .B(n17262), .Y(n17264));
  AOI22X1 g13900(.A0(n16538), .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B0(P1_REIP_REG_17__SCAN_IN), .B1(n16527), .Y(n17265));
  OAI21X1 g13901(.A0(n17264), .A1(n16558), .B0(n17265), .Y(n17266));
  NAND2X1 g13902(.A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .Y(n17267));
  NOR4X1  g13903(.A(n17122), .B(n17125), .C(n17137), .D(n17267), .Y(n17268));
  XOR2X1  g13904(.A(n17268), .B(n17256), .Y(n17269));
  NOR2X1  g13905(.A(n17269), .B(n16545), .Y(n17270));
  NAND4X1 g13906(.A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .C(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .D(n17168), .Y(n17271));
  XOR2X1  g13907(.A(n17271), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .Y(n17272));
  NOR3X1  g13908(.A(n17212), .B(n17195), .C(n17242), .Y(n17273));
  XOR2X1  g13909(.A(n17273), .B(n17256), .Y(n17274));
  OAI22X1 g13910(.A0(n17272), .A1(n16636), .B0(n18937), .B1(n17274), .Y(n17275));
  NOR3X1  g13911(.A(n17275), .B(n17270), .C(n17266), .Y(n17276));
  OAI21X1 g13912(.A0(n17260), .A1(n16571), .B0(n17276), .Y(P1_U3014));
  AOI22X1 g13913(.A0(n17231), .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B0(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B1(n17231), .Y(n17278));
  NOR2X1  g13914(.A(n17231), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .Y(n17279));
  AOI21X1 g13915(.A0(n17253), .A1(n17242), .B0(n17279), .Y(n17280));
  INVX1   g13916(.A(n17280), .Y(n17281));
  OAI22X1 g13917(.A0(n17279), .A1(n17278), .B0(n17227), .B1(n17281), .Y(n17282));
  INVX1   g13918(.A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .Y(n17283));
  XOR2X1  g13919(.A(n17231), .B(n17283), .Y(n17284));
  XOR2X1  g13920(.A(n17284), .B(n17282), .Y(n17285));
  AOI22X1 g13921(.A0(n16551), .A1(P1_EBX_REG_18__SCAN_IN), .B0(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .B1(n16553), .Y(n17286));
  XOR2X1  g13922(.A(n17286), .B(n15054), .Y(n17287));
  NOR3X1  g13923(.A(n17262), .B(n17238), .C(n17235), .Y(n17288));
  XOR2X1  g13924(.A(n17288), .B(n17287), .Y(n17289));
  AOI22X1 g13925(.A0(n16538), .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .B0(P1_REIP_REG_18__SCAN_IN), .B1(n16527), .Y(n17290));
  OAI21X1 g13926(.A0(n17289), .A1(n16558), .B0(n17290), .Y(n17291));
  NAND2X1 g13927(.A(n17268), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .Y(n17292));
  XOR2X1  g13928(.A(n17292), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .Y(n17293));
  NOR2X1  g13929(.A(n17293), .B(n16545), .Y(n17294));
  NOR2X1  g13930(.A(n17271), .B(n17256), .Y(n17295));
  XOR2X1  g13931(.A(n17295), .B(n17283), .Y(n17296));
  NOR4X1  g13932(.A(n17195), .B(n17242), .C(n17256), .D(n17212), .Y(n17297));
  XOR2X1  g13933(.A(n17297), .B(n17283), .Y(n17298));
  OAI22X1 g13934(.A0(n17296), .A1(n16636), .B0(n18937), .B1(n17298), .Y(n17299));
  NOR3X1  g13935(.A(n17299), .B(n17294), .C(n17291), .Y(n17300));
  OAI21X1 g13936(.A0(n17285), .A1(n16571), .B0(n17300), .Y(P1_U3013));
  AOI21X1 g13937(.A0(n17253), .A1(n17283), .B0(n17281), .Y(n17303));
  INVX1   g13938(.A(n17303), .Y(n17304));
  INVX1   g13939(.A(n17278), .Y(n17305));
  OAI21X1 g13940(.A0(n17256), .A1(n17283), .B0(n17253), .Y(n17306));
  AOI22X1 g13941(.A0(n17305), .A1(n17306), .B0(n17231), .B1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .Y(n17307));
  OAI21X1 g13942(.A0(n17304), .A1(n17227), .B0(n17307), .Y(n17308));
  INVX1   g13943(.A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .Y(n17309));
  XOR2X1  g13944(.A(n17231), .B(n17309), .Y(n17310));
  XOR2X1  g13945(.A(n17310), .B(n17308), .Y(n17311));
  AOI22X1 g13946(.A0(n16551), .A1(P1_EBX_REG_19__SCAN_IN), .B0(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B1(n16553), .Y(n17312));
  XOR2X1  g13947(.A(n17312), .B(n15054), .Y(n17313));
  NOR4X1  g13948(.A(n17262), .B(n17238), .C(n17235), .D(n17287), .Y(n17314));
  XOR2X1  g13949(.A(n17314), .B(n17313), .Y(n17315));
  AOI22X1 g13950(.A0(n16538), .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B0(P1_REIP_REG_19__SCAN_IN), .B1(n16527), .Y(n17316));
  OAI21X1 g13951(.A0(n17315), .A1(n16558), .B0(n17316), .Y(n17317));
  NAND3X1 g13952(.A(n17268), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .C(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .Y(n17318));
  XOR2X1  g13953(.A(n17318), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .Y(n17319));
  NOR2X1  g13954(.A(n17319), .B(n16545), .Y(n17320));
  NOR3X1  g13955(.A(n17271), .B(n17256), .C(n17283), .Y(n17321));
  XOR2X1  g13956(.A(n17321), .B(n17309), .Y(n17322));
  NAND2X1 g13957(.A(n17297), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .Y(n17323));
  XOR2X1  g13958(.A(n17323), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .Y(n17324));
  OAI22X1 g13959(.A0(n17322), .A1(n16636), .B0(n18937), .B1(n17324), .Y(n17325));
  NOR3X1  g13960(.A(n17325), .B(n17320), .C(n17317), .Y(n17326));
  OAI21X1 g13961(.A0(n17311), .A1(n16571), .B0(n17326), .Y(P1_U3012));
  OAI21X1 g13962(.A0(n17231), .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B0(n17308), .Y(n17328));
  OAI21X1 g13963(.A0(n17253), .A1(n17309), .B0(n17328), .Y(n17329));
  INVX1   g13964(.A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .Y(n17330));
  XOR2X1  g13965(.A(n17231), .B(n17330), .Y(n17331));
  XOR2X1  g13966(.A(n17331), .B(n17329), .Y(n17332));
  AOI22X1 g13967(.A0(n16551), .A1(P1_EBX_REG_20__SCAN_IN), .B0(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(n16553), .Y(n17333));
  XOR2X1  g13968(.A(n17333), .B(n15054), .Y(n17334));
  INVX1   g13969(.A(n17314), .Y(n17335));
  NOR2X1  g13970(.A(n17335), .B(n17313), .Y(n17336));
  XOR2X1  g13971(.A(n17336), .B(n17334), .Y(n17337));
  AOI22X1 g13972(.A0(n16538), .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B0(P1_REIP_REG_20__SCAN_IN), .B1(n16527), .Y(n17338));
  OAI21X1 g13973(.A0(n17337), .A1(n16558), .B0(n17338), .Y(n17339));
  NAND4X1 g13974(.A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .C(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .D(n17268), .Y(n17340));
  XOR2X1  g13975(.A(n17340), .B(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .Y(n17341));
  NOR2X1  g13976(.A(n17341), .B(n16545), .Y(n17342));
  NOR4X1  g13977(.A(n17256), .B(n17283), .C(n17309), .D(n17271), .Y(n17343));
  XOR2X1  g13978(.A(n17343), .B(n17330), .Y(n17344));
  NAND3X1 g13979(.A(n17297), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .C(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .Y(n17345));
  XOR2X1  g13980(.A(n17345), .B(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .Y(n17346));
  OAI22X1 g13981(.A0(n17344), .A1(n16636), .B0(n18937), .B1(n17346), .Y(n17347));
  NOR3X1  g13982(.A(n17347), .B(n17342), .C(n17339), .Y(n17348));
  OAI21X1 g13983(.A0(n17332), .A1(n16571), .B0(n17348), .Y(P1_U3011));
  OAI21X1 g13984(.A0(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B0(n17231), .Y(n17350));
  INVX1   g13985(.A(n17350), .Y(n17351));
  OAI21X1 g13986(.A0(n17309), .A1(n17330), .B0(n17253), .Y(n17352));
  AOI21X1 g13987(.A0(n17352), .A1(n17308), .B0(n17351), .Y(n17353));
  XOR2X1  g13988(.A(n17231), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .Y(n17354));
  XOR2X1  g13989(.A(n17354), .B(n17353), .Y(n17355));
  AOI22X1 g13990(.A0(n16551), .A1(P1_EBX_REG_21__SCAN_IN), .B0(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B1(n16553), .Y(n17356));
  XOR2X1  g13991(.A(n17356), .B(n15054), .Y(n17357));
  NOR3X1  g13992(.A(n17334), .B(n17335), .C(n17313), .Y(n17358));
  XOR2X1  g13993(.A(n17358), .B(n17357), .Y(n17359));
  AOI22X1 g13994(.A0(n16538), .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B0(P1_REIP_REG_21__SCAN_IN), .B1(n16527), .Y(n17360));
  OAI21X1 g13995(.A0(n17359), .A1(n16558), .B0(n17360), .Y(n17361));
  INVX1   g13996(.A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .Y(n17362));
  NOR3X1  g13997(.A(n17318), .B(n17309), .C(n17330), .Y(n17363));
  XOR2X1  g13998(.A(n17363), .B(n17362), .Y(n17364));
  NOR2X1  g13999(.A(n17364), .B(n16545), .Y(n17365));
  NAND2X1 g14000(.A(n17343), .B(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .Y(n17366));
  XOR2X1  g14001(.A(n17366), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .Y(n17367));
  NAND4X1 g14002(.A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .D(n17297), .Y(n17368));
  XOR2X1  g14003(.A(n17368), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .Y(n17369));
  OAI22X1 g14004(.A0(n17367), .A1(n16636), .B0(n18937), .B1(n17369), .Y(n17370));
  NOR3X1  g14005(.A(n17370), .B(n17365), .C(n17361), .Y(n17371));
  OAI21X1 g14006(.A0(n17355), .A1(n16571), .B0(n17371), .Y(P1_U3010));
  NOR4X1  g14007(.A(n16815), .B(n14821), .C(n17362), .D(n17257), .Y(n17374));
  NOR2X1  g14008(.A(n17374), .B(n17351), .Y(n17375));
  INVX1   g14009(.A(n17375), .Y(n17376));
  OAI21X1 g14010(.A0(n17231), .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B0(n17352), .Y(n17377));
  INVX1   g14011(.A(n17377), .Y(n17378));
  AOI21X1 g14012(.A0(n17378), .A1(n17308), .B0(n17376), .Y(n17379));
  XOR2X1  g14013(.A(n17231), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .Y(n17380));
  XOR2X1  g14014(.A(n17380), .B(n17379), .Y(n17381));
  AOI22X1 g14015(.A0(n16551), .A1(P1_EBX_REG_22__SCAN_IN), .B0(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B1(n16553), .Y(n17382));
  XOR2X1  g14016(.A(n17382), .B(n15054), .Y(n17383));
  NOR4X1  g14017(.A(n17334), .B(n17335), .C(n17313), .D(n17357), .Y(n17384));
  XOR2X1  g14018(.A(n17384), .B(n17383), .Y(n17385));
  AOI22X1 g14019(.A0(n16538), .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B0(P1_REIP_REG_22__SCAN_IN), .B1(n16527), .Y(n17386));
  OAI21X1 g14020(.A0(n17385), .A1(n16558), .B0(n17386), .Y(n17387));
  INVX1   g14021(.A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .Y(n17388));
  NOR4X1  g14022(.A(n17309), .B(n17330), .C(n17362), .D(n17318), .Y(n17389));
  XOR2X1  g14023(.A(n17389), .B(n17388), .Y(n17390));
  NOR2X1  g14024(.A(n17390), .B(n16545), .Y(n17391));
  NAND3X1 g14025(.A(n17343), .B(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .C(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .Y(n17392));
  XOR2X1  g14026(.A(n17392), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .Y(n17393));
  NOR2X1  g14027(.A(n17368), .B(n17362), .Y(n17394));
  XOR2X1  g14028(.A(n17394), .B(n17388), .Y(n17395));
  OAI22X1 g14029(.A0(n17393), .A1(n16636), .B0(n18937), .B1(n17395), .Y(n17396));
  NOR3X1  g14030(.A(n17396), .B(n17391), .C(n17387), .Y(n17397));
  OAI21X1 g14031(.A0(n17381), .A1(n16571), .B0(n17397), .Y(P1_U3009));
  NOR2X1  g14032(.A(n17231), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .Y(n17399));
  INVX1   g14033(.A(n17399), .Y(n17400));
  NAND3X1 g14034(.A(n17400), .B(n17378), .C(n17303), .Y(n17401));
  NOR4X1  g14035(.A(n16815), .B(n14821), .C(n17388), .D(n17257), .Y(n17405));
  NOR4X1  g14036(.A(n17377), .B(n17253), .C(n17283), .D(n17399), .Y(n17406));
  NOR4X1  g14037(.A(n17405), .B(n17305), .C(n17376), .D(n17406), .Y(n17407));
  OAI21X1 g14038(.A0(n17401), .A1(n17227), .B0(n17407), .Y(n17408));
  INVX1   g14039(.A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .Y(n17409));
  XOR2X1  g14040(.A(n17231), .B(n17409), .Y(n17410));
  XOR2X1  g14041(.A(n17410), .B(n17408), .Y(n17411));
  AOI22X1 g14042(.A0(n16551), .A1(P1_EBX_REG_23__SCAN_IN), .B0(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B1(n16553), .Y(n17412));
  XOR2X1  g14043(.A(n17412), .B(n15054), .Y(n17413));
  INVX1   g14044(.A(n17384), .Y(n17414));
  NOR2X1  g14045(.A(n17414), .B(n17383), .Y(n17415));
  XOR2X1  g14046(.A(n17415), .B(n17413), .Y(n17416));
  AOI22X1 g14047(.A0(n16538), .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B0(P1_REIP_REG_23__SCAN_IN), .B1(n16527), .Y(n17417));
  OAI21X1 g14048(.A0(n17416), .A1(n16558), .B0(n17417), .Y(n17418));
  NAND3X1 g14049(.A(n17363), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .Y(n17419));
  XOR2X1  g14050(.A(n17419), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .Y(n17420));
  NOR2X1  g14051(.A(n17420), .B(n16545), .Y(n17421));
  NAND4X1 g14052(.A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .D(n17343), .Y(n17422));
  XOR2X1  g14053(.A(n17422), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .Y(n17423));
  NOR3X1  g14054(.A(n17368), .B(n17362), .C(n17388), .Y(n17424));
  XOR2X1  g14055(.A(n17424), .B(n17409), .Y(n17425));
  OAI22X1 g14056(.A0(n17423), .A1(n16636), .B0(n18937), .B1(n17425), .Y(n17426));
  NOR3X1  g14057(.A(n17426), .B(n17421), .C(n17418), .Y(n17427));
  OAI21X1 g14058(.A0(n17411), .A1(n16571), .B0(n17427), .Y(P1_U3008));
  OAI21X1 g14059(.A0(n17231), .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B0(n17408), .Y(n17429));
  OAI21X1 g14060(.A0(n17253), .A1(n17409), .B0(n17429), .Y(n17430));
  INVX1   g14061(.A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .Y(n17431));
  XOR2X1  g14062(.A(n17231), .B(n17431), .Y(n17432));
  XOR2X1  g14063(.A(n17432), .B(n17430), .Y(n17433));
  AOI22X1 g14064(.A0(n16551), .A1(P1_EBX_REG_24__SCAN_IN), .B0(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B1(n16553), .Y(n17434));
  XOR2X1  g14065(.A(n17434), .B(n15054), .Y(n17435));
  NOR3X1  g14066(.A(n17413), .B(n17414), .C(n17383), .Y(n17436));
  XOR2X1  g14067(.A(n17436), .B(n17435), .Y(n17437));
  AOI22X1 g14068(.A0(n16538), .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B0(P1_REIP_REG_24__SCAN_IN), .B1(n16527), .Y(n17438));
  OAI21X1 g14069(.A0(n17437), .A1(n16558), .B0(n17438), .Y(n17439));
  NAND4X1 g14070(.A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .C(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .D(n17363), .Y(n17440));
  XOR2X1  g14071(.A(n17440), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .Y(n17441));
  NOR2X1  g14072(.A(n17441), .B(n16545), .Y(n17442));
  NOR2X1  g14073(.A(n17422), .B(n17409), .Y(n17443));
  XOR2X1  g14074(.A(n17443), .B(n17431), .Y(n17444));
  NOR4X1  g14075(.A(n17362), .B(n17388), .C(n17409), .D(n17368), .Y(n17445));
  XOR2X1  g14076(.A(n17445), .B(n17431), .Y(n17446));
  OAI22X1 g14077(.A0(n17444), .A1(n16636), .B0(n18937), .B1(n17446), .Y(n17447));
  NOR3X1  g14078(.A(n17447), .B(n17442), .C(n17439), .Y(n17448));
  OAI21X1 g14079(.A0(n17433), .A1(n16571), .B0(n17448), .Y(P1_U3007));
  OAI21X1 g14080(.A0(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B0(n17231), .Y(n17450));
  OAI21X1 g14081(.A0(n17409), .A1(n17431), .B0(n17253), .Y(n17451));
  NAND2X1 g14082(.A(n17451), .B(n17408), .Y(n17452));
  NAND2X1 g14083(.A(n17452), .B(n17450), .Y(n17453));
  INVX1   g14084(.A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .Y(n17454));
  XOR2X1  g14085(.A(n17231), .B(n17454), .Y(n17455));
  XOR2X1  g14086(.A(n17455), .B(n17453), .Y(n17456));
  AOI22X1 g14087(.A0(n16551), .A1(P1_EBX_REG_25__SCAN_IN), .B0(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B1(n16553), .Y(n17457));
  XOR2X1  g14088(.A(n17457), .B(n15054), .Y(n17458));
  NOR4X1  g14089(.A(n17413), .B(n17414), .C(n17383), .D(n17435), .Y(n17459));
  XOR2X1  g14090(.A(n17459), .B(n17458), .Y(n17460));
  AOI22X1 g14091(.A0(n16538), .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B0(P1_REIP_REG_25__SCAN_IN), .B1(n16527), .Y(n17461));
  OAI21X1 g14092(.A0(n17460), .A1(n16558), .B0(n17461), .Y(n17462));
  NOR3X1  g14093(.A(n17419), .B(n17409), .C(n17431), .Y(n17463));
  XOR2X1  g14094(.A(n17463), .B(n17454), .Y(n17464));
  NOR2X1  g14095(.A(n17464), .B(n16545), .Y(n17465));
  NOR3X1  g14096(.A(n17422), .B(n17409), .C(n17431), .Y(n17466));
  XOR2X1  g14097(.A(n17466), .B(n17454), .Y(n17467));
  NAND2X1 g14098(.A(n17445), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .Y(n17468));
  XOR2X1  g14099(.A(n17468), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .Y(n17469));
  OAI22X1 g14100(.A0(n17467), .A1(n16636), .B0(n18937), .B1(n17469), .Y(n17470));
  NOR3X1  g14101(.A(n17470), .B(n17465), .C(n17462), .Y(n17471));
  OAI21X1 g14102(.A0(n17456), .A1(n16571), .B0(n17471), .Y(P1_U3006));
  OAI21X1 g14103(.A0(n17231), .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B0(n17451), .Y(n17473));
  INVX1   g14104(.A(n17473), .Y(n17474));
  OAI21X1 g14105(.A0(n17253), .A1(n17454), .B0(n17450), .Y(n17477));
  AOI21X1 g14106(.A0(n17474), .A1(n17408), .B0(n17477), .Y(n17478));
  INVX1   g14107(.A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .Y(n17479));
  XOR2X1  g14108(.A(n17231), .B(n17479), .Y(n17480));
  XOR2X1  g14109(.A(n17480), .B(n17478), .Y(n17481));
  NAND2X1 g14110(.A(n17481), .B(n16572), .Y(n17482));
  AOI22X1 g14111(.A0(n16551), .A1(P1_EBX_REG_26__SCAN_IN), .B0(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B1(n16553), .Y(n17483));
  XOR2X1  g14112(.A(n17483), .B(n15054), .Y(n17484));
  INVX1   g14113(.A(n17459), .Y(n17485));
  NOR2X1  g14114(.A(n17485), .B(n17458), .Y(n17486));
  XOR2X1  g14115(.A(n17486), .B(n17484), .Y(n17487));
  NOR2X1  g14116(.A(n17487), .B(n16558), .Y(n17488));
  NOR4X1  g14117(.A(n17409), .B(n17431), .C(n17454), .D(n17419), .Y(n17489));
  XOR2X1  g14118(.A(n17489), .B(n17479), .Y(n17490));
  AOI22X1 g14119(.A0(n16538), .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B0(P1_REIP_REG_26__SCAN_IN), .B1(n16527), .Y(n17491));
  OAI21X1 g14120(.A0(n17490), .A1(n16545), .B0(n17491), .Y(n17492));
  NOR4X1  g14121(.A(n17409), .B(n17431), .C(n17454), .D(n17422), .Y(n17493));
  XOR2X1  g14122(.A(n17493), .B(n17479), .Y(n17494));
  NAND3X1 g14123(.A(n17445), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .C(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .Y(n17495));
  XOR2X1  g14124(.A(n17495), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .Y(n17496));
  OAI22X1 g14125(.A0(n17494), .A1(n16636), .B0(n18937), .B1(n17496), .Y(n17497));
  NOR3X1  g14126(.A(n17497), .B(n17492), .C(n17488), .Y(n17498));
  NAND2X1 g14127(.A(n17498), .B(n17482), .Y(P1_U3005));
  AOI21X1 g14128(.A0(n17253), .A1(n17479), .B0(n17473), .Y(n17500));
  OAI21X1 g14129(.A0(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B0(n17231), .Y(n17501));
  AOI22X1 g14130(.A0(n17450), .A1(n17501), .B0(n17253), .B1(n17479), .Y(n17502));
  AOI21X1 g14131(.A0(n17500), .A1(n17408), .B0(n17502), .Y(n17503));
  INVX1   g14132(.A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .Y(n17504));
  XOR2X1  g14133(.A(n17231), .B(n17504), .Y(n17505));
  XOR2X1  g14134(.A(n17505), .B(n17503), .Y(n17506));
  NAND2X1 g14135(.A(n17506), .B(n16572), .Y(n17507));
  AOI22X1 g14136(.A0(n16551), .A1(P1_EBX_REG_27__SCAN_IN), .B0(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B1(n16553), .Y(n17508));
  XOR2X1  g14137(.A(n17508), .B(n15054), .Y(n17509));
  NOR3X1  g14138(.A(n17484), .B(n17485), .C(n17458), .Y(n17510));
  XOR2X1  g14139(.A(n17510), .B(n17509), .Y(n17511));
  NOR2X1  g14140(.A(n17511), .B(n16558), .Y(n17512));
  NAND3X1 g14141(.A(n17463), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .C(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .Y(n17513));
  XOR2X1  g14142(.A(n17513), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .Y(n17514));
  AOI22X1 g14143(.A0(n16538), .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B0(P1_REIP_REG_27__SCAN_IN), .B1(n16527), .Y(n17515));
  OAI21X1 g14144(.A0(n17514), .A1(n16545), .B0(n17515), .Y(n17516));
  NAND2X1 g14145(.A(n17493), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .Y(n17517));
  XOR2X1  g14146(.A(n17517), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .Y(n17518));
  NAND4X1 g14147(.A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .C(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .D(n17445), .Y(n17519));
  XOR2X1  g14148(.A(n17519), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .Y(n17520));
  OAI22X1 g14149(.A0(n17518), .A1(n16636), .B0(n18937), .B1(n17520), .Y(n17521));
  NOR3X1  g14150(.A(n17521), .B(n17516), .C(n17512), .Y(n17522));
  NAND2X1 g14151(.A(n17522), .B(n17507), .Y(P1_U3004));
  NOR2X1  g14152(.A(n17231), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .Y(n17524));
  OAI21X1 g14153(.A0(n17479), .A1(n17504), .B0(n17253), .Y(n17525));
  INVX1   g14154(.A(n17525), .Y(n17526));
  NOR2X1  g14155(.A(n17526), .B(n17473), .Y(n17527));
  NAND2X1 g14156(.A(n17527), .B(n17408), .Y(n17528));
  AOI21X1 g14157(.A0(n17231), .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B0(n17502), .Y(n17529));
  OAI21X1 g14158(.A0(n17529), .A1(n17524), .B0(n17528), .Y(n17530));
  INVX1   g14159(.A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .Y(n17531));
  XOR2X1  g14160(.A(n17231), .B(n17531), .Y(n17532));
  XOR2X1  g14161(.A(n17532), .B(n17530), .Y(n17533));
  AOI22X1 g14162(.A0(n16551), .A1(P1_EBX_REG_28__SCAN_IN), .B0(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B1(n16553), .Y(n17534));
  XOR2X1  g14163(.A(n17534), .B(n15054), .Y(n17535));
  NOR4X1  g14164(.A(n17484), .B(n17485), .C(n17458), .D(n17509), .Y(n17536));
  XOR2X1  g14165(.A(n17536), .B(n17535), .Y(n17537));
  NOR2X1  g14166(.A(n17537), .B(n16558), .Y(n17538));
  NAND4X1 g14167(.A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .C(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .D(n17463), .Y(n17539));
  XOR2X1  g14168(.A(n17539), .B(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .Y(n17540));
  AOI22X1 g14169(.A0(n16538), .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B0(P1_REIP_REG_28__SCAN_IN), .B1(n16527), .Y(n17541));
  OAI21X1 g14170(.A0(n17540), .A1(n16545), .B0(n17541), .Y(n17542));
  NAND3X1 g14171(.A(n17493), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .C(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .Y(n17543));
  XOR2X1  g14172(.A(n17543), .B(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .Y(n17544));
  NOR2X1  g14173(.A(n17519), .B(n17504), .Y(n17545));
  XOR2X1  g14174(.A(n17545), .B(n17531), .Y(n17546));
  OAI22X1 g14175(.A0(n17544), .A1(n16636), .B0(n18937), .B1(n17546), .Y(n17547));
  NOR3X1  g14176(.A(n17547), .B(n17542), .C(n17538), .Y(n17548));
  OAI21X1 g14177(.A0(n17533), .A1(n16571), .B0(n17548), .Y(P1_U3003));
  INVX1   g14178(.A(n17527), .Y(n17550));
  NOR2X1  g14179(.A(n17231), .B(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .Y(n17551));
  NOR4X1  g14180(.A(n17399), .B(n17377), .C(n17304), .D(n17551), .Y(n17552));
  INVX1   g14181(.A(n17552), .Y(n17553));
  NOR3X1  g14182(.A(n17553), .B(n17550), .C(n17227), .Y(n17554));
  INVX1   g14183(.A(n17551), .Y(n17555));
  NAND3X1 g14184(.A(n17555), .B(n17527), .C(n17406), .Y(n17556));
  OAI21X1 g14185(.A0(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B0(n17231), .Y(n17558));
  INVX1   g14186(.A(n17558), .Y(n17559));
  NOR3X1  g14187(.A(n17405), .B(n17559), .C(n17406), .Y(n17561));
  INVX1   g14188(.A(n17502), .Y(n17563));
  NAND4X1 g14189(.A(n17278), .B(n17563), .C(n17561), .D(n17375), .Y(n17570));
  NOR2X1  g14190(.A(n17570), .B(n17554), .Y(n17571));
  INVX1   g14191(.A(n17571), .Y(n17572));
  INVX1   g14192(.A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .Y(n17573));
  XOR2X1  g14193(.A(n17231), .B(n17573), .Y(n17574));
  XOR2X1  g14194(.A(n17574), .B(n17572), .Y(n17575));
  AOI22X1 g14195(.A0(n16551), .A1(P1_EBX_REG_29__SCAN_IN), .B0(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .B1(n16553), .Y(n17576));
  XOR2X1  g14196(.A(n17576), .B(n15054), .Y(n17577));
  INVX1   g14197(.A(n17536), .Y(n17578));
  NOR2X1  g14198(.A(n17578), .B(n17535), .Y(n17579));
  XOR2X1  g14199(.A(n17579), .B(n17577), .Y(n17580));
  NOR2X1  g14200(.A(n17580), .B(n16558), .Y(n17581));
  NOR3X1  g14201(.A(n17513), .B(n17504), .C(n17531), .Y(n17582));
  XOR2X1  g14202(.A(n17582), .B(n17573), .Y(n17583));
  AOI22X1 g14203(.A0(n16538), .A1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .B0(P1_REIP_REG_29__SCAN_IN), .B1(n16527), .Y(n17584));
  OAI21X1 g14204(.A0(n17583), .A1(n16545), .B0(n17584), .Y(n17585));
  NAND4X1 g14205(.A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .C(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .D(n17493), .Y(n17586));
  XOR2X1  g14206(.A(n17586), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .Y(n17587));
  NOR3X1  g14207(.A(n17519), .B(n17504), .C(n17531), .Y(n17588));
  XOR2X1  g14208(.A(n17588), .B(n17573), .Y(n17589));
  OAI22X1 g14209(.A0(n17587), .A1(n16636), .B0(n18937), .B1(n17589), .Y(n17590));
  NOR3X1  g14210(.A(n17590), .B(n17585), .C(n17581), .Y(n17591));
  OAI21X1 g14211(.A0(n17575), .A1(n16571), .B0(n17591), .Y(P1_U3002));
  NOR2X1  g14212(.A(n17231), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .Y(n17593));
  NOR4X1  g14213(.A(n17553), .B(n17550), .C(n17227), .D(n17593), .Y(n17594));
  NOR2X1  g14214(.A(n17593), .B(n17561), .Y(n17595));
  NOR4X1  g14215(.A(n16815), .B(n14821), .C(n17573), .D(n17257), .Y(n17596));
  INVX1   g14216(.A(n17596), .Y(n17597));
  OAI21X1 g14217(.A0(n17593), .A1(n17375), .B0(n17597), .Y(n17598));
  AOI21X1 g14218(.A0(n17278), .A1(n17563), .B0(n17593), .Y(n17599));
  NOR4X1  g14219(.A(n17598), .B(n17595), .C(n17594), .D(n17599), .Y(n17600));
  INVX1   g14220(.A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .Y(n17601));
  XOR2X1  g14221(.A(n17231), .B(n17601), .Y(n17602));
  INVX1   g14222(.A(n17602), .Y(n17603));
  XOR2X1  g14223(.A(n17603), .B(n17600), .Y(n17604));
  AOI22X1 g14224(.A0(n16551), .A1(P1_EBX_REG_30__SCAN_IN), .B0(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B1(n16553), .Y(n17605));
  XOR2X1  g14225(.A(n17605), .B(n15054), .Y(n17606));
  NOR3X1  g14226(.A(n17577), .B(n17578), .C(n17535), .Y(n17607));
  XOR2X1  g14227(.A(n17607), .B(n17606), .Y(n17608));
  NOR2X1  g14228(.A(n17608), .B(n16558), .Y(n17609));
  NOR4X1  g14229(.A(n17504), .B(n17531), .C(n17573), .D(n17513), .Y(n17610));
  XOR2X1  g14230(.A(n17610), .B(n17601), .Y(n17611));
  AOI22X1 g14231(.A0(n16538), .A1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B0(P1_REIP_REG_30__SCAN_IN), .B1(n16527), .Y(n17612));
  OAI21X1 g14232(.A0(n17611), .A1(n16545), .B0(n17612), .Y(n17613));
  NOR2X1  g14233(.A(n17586), .B(n17573), .Y(n17614));
  XOR2X1  g14234(.A(n17614), .B(n17601), .Y(n17615));
  NOR4X1  g14235(.A(n17504), .B(n17531), .C(n17573), .D(n17519), .Y(n17616));
  XOR2X1  g14236(.A(n17616), .B(n17601), .Y(n17617));
  OAI22X1 g14237(.A0(n17615), .A1(n16636), .B0(n18937), .B1(n17617), .Y(n17618));
  NOR3X1  g14238(.A(n17618), .B(n17613), .C(n17609), .Y(n17619));
  OAI21X1 g14239(.A0(n17604), .A1(n16571), .B0(n17619), .Y(P1_U3001));
  XOR2X1  g14240(.A(n17231), .B(n15250), .Y(n17621));
  NOR2X1  g14241(.A(n17231), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .Y(n17622));
  NOR4X1  g14242(.A(n17621), .B(n17593), .C(n17571), .D(n17622), .Y(n17623));
  INVX1   g14243(.A(n17621), .Y(n17628));
  AOI21X1 g14244(.A0(n17573), .A1(n17601), .B0(n17253), .Y(n17633));
  NOR4X1  g14245(.A(n17559), .B(n17376), .C(n17628), .D(n17633), .Y(n17634));
  OAI21X1 g14246(.A0(n17593), .A1(n17556), .B0(n17634), .Y(n17635));
  NOR4X1  g14247(.A(n17405), .B(n17305), .C(n17502), .D(n17635), .Y(n17636));
  INVX1   g14248(.A(n17636), .Y(n17637));
  NOR2X1  g14249(.A(n17637), .B(n17594), .Y(n17638));
  NOR3X1  g14250(.A(n17622), .B(n17621), .C(n17597), .Y(n17639));
  NOR3X1  g14251(.A(n17253), .B(n17601), .C(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .Y(n17640));
  NOR3X1  g14252(.A(n17231), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .C(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .Y(n17641));
  NOR3X1  g14253(.A(n17641), .B(n17640), .C(n17639), .Y(n17642));
  INVX1   g14254(.A(n17642), .Y(n17643));
  NOR3X1  g14255(.A(n17643), .B(n17638), .C(n17623), .Y(n17644));
  NAND2X1 g14256(.A(n17644), .B(n16572), .Y(n17645));
  AOI22X1 g14257(.A0(n16551), .A1(P1_EBX_REG_31__SCAN_IN), .B0(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(n16553), .Y(n17646));
  XOR2X1  g14258(.A(n17646), .B(n15054), .Y(n17647));
  NOR4X1  g14259(.A(n17577), .B(n17578), .C(n17535), .D(n17606), .Y(n17648));
  XOR2X1  g14260(.A(n17648), .B(n17647), .Y(n17649));
  NOR2X1  g14261(.A(n17649), .B(n16558), .Y(n17650));
  NAND2X1 g14262(.A(n17610), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .Y(n17651));
  XOR2X1  g14263(.A(n17651), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .Y(n17652));
  AOI22X1 g14264(.A0(n16538), .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B0(P1_REIP_REG_31__SCAN_IN), .B1(n16527), .Y(n17653));
  OAI21X1 g14265(.A0(n17652), .A1(n16545), .B0(n17653), .Y(n17654));
  NOR3X1  g14266(.A(n17586), .B(n17573), .C(n17601), .Y(n17655));
  XOR2X1  g14267(.A(n17655), .B(n15250), .Y(n17656));
  NAND2X1 g14268(.A(n17616), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .Y(n17657));
  XOR2X1  g14269(.A(n17657), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .Y(n17658));
  OAI22X1 g14270(.A0(n17656), .A1(n16636), .B0(n18937), .B1(n17658), .Y(n17659));
  NOR3X1  g14271(.A(n17659), .B(n17654), .C(n17650), .Y(n17660));
  NAND2X1 g14272(.A(n17660), .B(n17645), .Y(P1_U3000));
  NOR2X1  g14273(.A(P1_STATE2_REG_2__SCAN_IN), .B(P1_STATEBS16_REG_SCAN_IN), .Y(n17662));
  INVX1   g14274(.A(n17662), .Y(n17663));
  NOR2X1  g14275(.A(n15042), .B(n15155), .Y(n17664));
  NOR2X1  g14276(.A(n17664), .B(n14998), .Y(n17665));
  AOI21X1 g14277(.A0(n17665), .A1(n15407), .B0(n15155), .Y(n17666));
  OAI21X1 g14278(.A0(n14919), .A1(n14770), .B0(P1_STATE2_REG_2__SCAN_IN), .Y(n17667));
  NOR3X1  g14279(.A(n14962), .B(n14919), .C(n15155), .Y(n17668));
  INVX1   g14280(.A(P1_EAX_REG_0__SCAN_IN), .Y(n17669));
  INVX1   g14281(.A(n17664), .Y(n17670));
  NOR2X1  g14282(.A(P1_STATE2_REG_2__SCAN_IN), .B(n15305), .Y(n17671));
  OAI21X1 g14283(.A0(n17671), .A1(n17662), .B0(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .Y(n17672));
  OAI21X1 g14284(.A0(n17670), .A1(n17669), .B0(n17672), .Y(n17673));
  AOI21X1 g14285(.A0(n17668), .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B0(n17673), .Y(n17674));
  OAI21X1 g14286(.A0(n17667), .A1(n15132), .B0(n17674), .Y(n17675));
  XOR2X1  g14287(.A(n17675), .B(n17663), .Y(n17676));
  INVX1   g14288(.A(n17676), .Y(n17677));
  XOR2X1  g14289(.A(n17677), .B(n17666), .Y(n17678));
  XOR2X1  g14290(.A(n17678), .B(n17663), .Y(n17679));
  INVX1   g14291(.A(n15289), .Y(n17680));
  NAND4X1 g14292(.A(n15024), .B(n14804), .C(n15093), .D(n14984), .Y(n17681));
  NOR4X1  g14293(.A(n17680), .B(n14993), .C(n15155), .D(n17681), .Y(n17682));
  INVX1   g14294(.A(n17682), .Y(n17683));
  OAI21X1 g14295(.A0(n16508), .A1(n15309), .B0(n14650), .Y(n17684));
  NAND2X1 g14296(.A(n17684), .B(n17683), .Y(n17685));
  INVX1   g14297(.A(n17685), .Y(n17686));
  NOR3X1  g14298(.A(n17686), .B(n15093), .C(n15305), .Y(n17687));
  INVX1   g14299(.A(n17687), .Y(n17688));
  INVX1   g14300(.A(P1_REIP_REG_0__SCAN_IN), .Y(n17690));
  AOI22X1 g14301(.A0(P1_STATE2_REG_1__SCAN_IN), .A1(n15305), .B0(P1_STATE2_REG_2__SCAN_IN), .B1(n14650), .Y(n17693));
  AOI21X1 g14302(.A0(n17684), .A1(n17683), .B0(n17693), .Y(n17694));
  OAI21X1 g14303(.A0(n17694), .A1(n17686), .B0(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .Y(n17695));
  OAI21X1 g14304(.A0(n16586), .A1(n17690), .B0(n17695), .Y(n17696));
  AOI21X1 g14305(.A0(n17682), .A1(n16515), .B0(n17696), .Y(n17697));
  OAI21X1 g14306(.A0(n17688), .A1(n17679), .B0(n17697), .Y(P1_U2999));
  OAI21X1 g14307(.A0(n16584), .A1(n16581), .B0(n17682), .Y(n17699));
  INVX1   g14308(.A(P1_EAX_REG_1__SCAN_IN), .Y(n17700));
  INVX1   g14309(.A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .Y(n17701));
  NOR3X1  g14310(.A(P1_STATE2_REG_2__SCAN_IN), .B(n17701), .C(n15305), .Y(n17702));
  AOI21X1 g14311(.A0(n17662), .A1(n17701), .B0(n17702), .Y(n17703));
  OAI21X1 g14312(.A0(n17670), .A1(n17700), .B0(n17703), .Y(n17704));
  AOI21X1 g14313(.A0(n17668), .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B0(n17704), .Y(n17705));
  OAI21X1 g14314(.A0(n17667), .A1(n15169), .B0(n17705), .Y(n17706));
  XOR2X1  g14315(.A(n17706), .B(n17663), .Y(n17707));
  NOR3X1  g14316(.A(n17707), .B(n17667), .C(n15434), .Y(n17708));
  OAI21X1 g14317(.A0(n17667), .A1(n15434), .B0(n17707), .Y(n17709));
  INVX1   g14318(.A(n17709), .Y(n17710));
  NOR2X1  g14319(.A(n17710), .B(n17708), .Y(n17711));
  NOR2X1  g14320(.A(n17677), .B(n17666), .Y(n17712));
  NOR2X1  g14321(.A(n17712), .B(n17663), .Y(n17713));
  AOI21X1 g14322(.A0(n17677), .A1(n17666), .B0(n17713), .Y(n17714));
  XOR2X1  g14323(.A(n17714), .B(n17711), .Y(n17715));
  INVX1   g14324(.A(n17715), .Y(n17716));
  NAND2X1 g14325(.A(n17716), .B(n17687), .Y(n17717));
  NAND4X1 g14326(.A(n15093), .B(n15155), .C(P1_REIP_REG_1__SCAN_IN), .D(n17685), .Y(n17718));
  NOR2X1  g14327(.A(n17685), .B(n17701), .Y(n17719));
  AOI21X1 g14328(.A0(n17694), .A1(n17701), .B0(n17719), .Y(n17720));
  NAND4X1 g14329(.A(n17718), .B(n17717), .C(n17699), .D(n17720), .Y(P1_U2998));
  INVX1   g14330(.A(n17708), .Y(n17722));
  OAI21X1 g14331(.A0(n17714), .A1(n17710), .B0(n17722), .Y(n17723));
  INVX1   g14332(.A(n17723), .Y(n17724));
  INVX1   g14333(.A(n17671), .Y(n17725));
  OAI21X1 g14334(.A0(n17667), .A1(n15459), .B0(n17725), .Y(n17726));
  INVX1   g14335(.A(P1_EAX_REG_2__SCAN_IN), .Y(n17727));
  XOR2X1  g14336(.A(n17701), .B(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .Y(n17728));
  INVX1   g14337(.A(n17728), .Y(n17729));
  AOI22X1 g14338(.A0(n17671), .A1(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B0(n17662), .B1(n17729), .Y(n17730));
  OAI21X1 g14339(.A0(n17670), .A1(n17727), .B0(n17730), .Y(n17731));
  AOI21X1 g14340(.A0(n17668), .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B0(n17731), .Y(n17732));
  OAI21X1 g14341(.A0(n17667), .A1(n15192), .B0(n17732), .Y(n17733));
  XOR2X1  g14342(.A(n17733), .B(n17663), .Y(n17734));
  INVX1   g14343(.A(n17734), .Y(n17735));
  NOR2X1  g14344(.A(n17735), .B(n17726), .Y(n17736));
  NOR2X1  g14345(.A(n17736), .B(n17724), .Y(n17737));
  NAND2X1 g14346(.A(n17735), .B(n17726), .Y(n17738));
  XOR2X1  g14347(.A(n17734), .B(n17726), .Y(n17739));
  AOI22X1 g14348(.A0(n17738), .A1(n17737), .B0(n17724), .B1(n17739), .Y(n17740));
  INVX1   g14349(.A(n17740), .Y(n17741));
  AOI22X1 g14350(.A0(n17694), .A1(n17729), .B0(n17686), .B1(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .Y(n17742));
  OAI21X1 g14351(.A0(n16586), .A1(n14538), .B0(n17742), .Y(n17743));
  AOI21X1 g14352(.A0(n17682), .A1(n16598), .B0(n17743), .Y(n17744));
  OAI21X1 g14353(.A0(n17741), .A1(n17688), .B0(n17744), .Y(P1_U2997));
  INVX1   g14354(.A(n17667), .Y(n17747));
  NAND2X1 g14355(.A(n17668), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Y(n17748));
  NAND3X1 g14356(.A(n14962), .B(P1_STATE2_REG_2__SCAN_IN), .C(P1_EAX_REG_3__SCAN_IN), .Y(n17749));
  NAND2X1 g14357(.A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .Y(n17750));
  XOR2X1  g14358(.A(n17750), .B(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .Y(n17751));
  INVX1   g14359(.A(n17751), .Y(n17752));
  AOI22X1 g14360(.A0(n17671), .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B0(n17662), .B1(n17752), .Y(n17753));
  NAND3X1 g14361(.A(n17753), .B(n17749), .C(n17748), .Y(n17754));
  AOI21X1 g14362(.A0(n17747), .A1(n15218), .B0(n17754), .Y(n17755));
  XOR2X1  g14363(.A(n17755), .B(n17662), .Y(n17756));
  INVX1   g14364(.A(n17756), .Y(n17757));
  AOI21X1 g14365(.A0(n17747), .A1(n15483), .B0(n17757), .Y(n17758));
  NOR3X1  g14366(.A(n17756), .B(n17667), .C(n15484), .Y(n17759));
  NOR2X1  g14367(.A(n17759), .B(n17758), .Y(n17760));
  OAI21X1 g14368(.A0(n17736), .A1(n17724), .B0(n17738), .Y(n17761));
  XOR2X1  g14369(.A(n17761), .B(n17760), .Y(n17762));
  NAND4X1 g14370(.A(n15093), .B(n15155), .C(P1_REIP_REG_3__SCAN_IN), .D(n17685), .Y(n17763));
  AOI22X1 g14371(.A0(n17694), .A1(n17752), .B0(n17686), .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .Y(n17764));
  NAND2X1 g14372(.A(n17764), .B(n17763), .Y(n17765));
  AOI21X1 g14373(.A0(n17762), .A1(n17687), .B0(n17765), .Y(n17766));
  OAI21X1 g14374(.A0(n17683), .A1(n16625), .B0(n17766), .Y(P1_U2996));
  NOR2X1  g14375(.A(n17667), .B(n16673), .Y(n17768));
  INVX1   g14376(.A(P1_EAX_REG_4__SCAN_IN), .Y(n17769));
  INVX1   g14377(.A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .Y(n17770));
  NAND3X1 g14378(.A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .C(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .Y(n17771));
  XOR2X1  g14379(.A(n17771), .B(n17770), .Y(n17772));
  AOI22X1 g14380(.A0(n17671), .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B0(n17662), .B1(n17772), .Y(n17773));
  OAI21X1 g14381(.A0(n17670), .A1(n17769), .B0(n17773), .Y(n17774));
  AOI21X1 g14382(.A0(n17668), .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B0(n17774), .Y(n17775));
  OAI21X1 g14383(.A0(n17667), .A1(n15243), .B0(n17775), .Y(n17776));
  XOR2X1  g14384(.A(n17776), .B(n17663), .Y(n17777));
  INVX1   g14385(.A(n17777), .Y(n17778));
  XOR2X1  g14386(.A(n17778), .B(n17768), .Y(n17779));
  AOI21X1 g14387(.A0(n17677), .A1(n17666), .B0(n17662), .Y(n17780));
  NOR3X1  g14388(.A(n17780), .B(n17710), .C(n17712), .Y(n17781));
  INVX1   g14389(.A(n17781), .Y(n17782));
  NAND3X1 g14390(.A(n17782), .B(n17738), .C(n17722), .Y(n17783));
  NOR2X1  g14391(.A(n17758), .B(n17736), .Y(n17784));
  AOI21X1 g14392(.A0(n17784), .A1(n17783), .B0(n17759), .Y(n17785));
  XOR2X1  g14393(.A(n17785), .B(n17779), .Y(n17786));
  NOR2X1  g14394(.A(n17786), .B(n17688), .Y(n17787));
  AOI22X1 g14395(.A0(n17694), .A1(n17772), .B0(n17686), .B1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .Y(n17788));
  OAI21X1 g14396(.A0(n16586), .A1(n14532), .B0(n17788), .Y(n17789));
  NOR2X1  g14397(.A(n17789), .B(n17787), .Y(n17790));
  OAI21X1 g14398(.A0(n17683), .A1(n16677), .B0(n17790), .Y(P1_U2995));
  NOR4X1  g14399(.A(n15217), .B(n15191), .C(n15241), .D(n15240), .Y(n17792));
  NAND2X1 g14400(.A(n17792), .B(n17747), .Y(n17793));
  INVX1   g14401(.A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .Y(n17794));
  NAND4X1 g14402(.A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .C(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .D(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .Y(n17795));
  XOR2X1  g14403(.A(n17795), .B(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .Y(n17796));
  OAI22X1 g14404(.A0(n17725), .A1(n17794), .B0(n17663), .B1(n17796), .Y(n17797));
  AOI21X1 g14405(.A0(n17664), .A1(P1_EAX_REG_5__SCAN_IN), .B0(n17797), .Y(n17798));
  NAND2X1 g14406(.A(n17798), .B(n17793), .Y(n17799));
  XOR2X1  g14407(.A(n17799), .B(n17663), .Y(n17800));
  NOR3X1  g14408(.A(n17800), .B(n17667), .C(n16729), .Y(n17801));
  OAI21X1 g14409(.A0(n17667), .A1(n16729), .B0(n17800), .Y(n17802));
  INVX1   g14410(.A(n17802), .Y(n17803));
  NOR2X1  g14411(.A(n17803), .B(n17801), .Y(n17804));
  NOR3X1  g14412(.A(n17777), .B(n17667), .C(n16673), .Y(n17805));
  NOR2X1  g14413(.A(n17778), .B(n17768), .Y(n17806));
  NOR2X1  g14414(.A(n17785), .B(n17806), .Y(n17807));
  NOR2X1  g14415(.A(n17807), .B(n17805), .Y(n17808));
  XOR2X1  g14416(.A(n17808), .B(n17804), .Y(n17809));
  NOR2X1  g14417(.A(n17809), .B(n17688), .Y(n17810));
  INVX1   g14418(.A(n17796), .Y(n17811));
  AOI22X1 g14419(.A0(n17694), .A1(n17811), .B0(n17686), .B1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .Y(n17812));
  OAI21X1 g14420(.A0(n16586), .A1(n14529), .B0(n17812), .Y(n17813));
  NOR2X1  g14421(.A(n17813), .B(n17810), .Y(n17814));
  OAI21X1 g14422(.A0(n17683), .A1(n16737), .B0(n17814), .Y(P1_U2994));
  INVX1   g14423(.A(n17801), .Y(n17816));
  OAI21X1 g14424(.A0(n17808), .A1(n17803), .B0(n17816), .Y(n17817));
  INVX1   g14425(.A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .Y(n17818));
  NOR2X1  g14426(.A(n17795), .B(n17794), .Y(n17819));
  XOR2X1  g14427(.A(n17819), .B(n17818), .Y(n17820));
  OAI22X1 g14428(.A0(n17725), .A1(n17818), .B0(n17663), .B1(n17820), .Y(n17821));
  AOI21X1 g14429(.A0(n17664), .A1(P1_EAX_REG_6__SCAN_IN), .B0(n17821), .Y(n17822));
  XOR2X1  g14430(.A(n17822), .B(n17662), .Y(n17823));
  INVX1   g14431(.A(n17823), .Y(n17824));
  AOI21X1 g14432(.A0(n17747), .A1(n16780), .B0(n17824), .Y(n17825));
  INVX1   g14433(.A(n17825), .Y(n17826));
  NAND3X1 g14434(.A(n17824), .B(n17747), .C(n16780), .Y(n17827));
  NAND3X1 g14435(.A(n17827), .B(n17826), .C(n17817), .Y(n17828));
  INVX1   g14436(.A(n17827), .Y(n17829));
  NOR2X1  g14437(.A(n17829), .B(n17825), .Y(n17830));
  OAI21X1 g14438(.A0(n17830), .A1(n17817), .B0(n17828), .Y(n17831));
  NOR2X1  g14439(.A(n17831), .B(n17688), .Y(n17832));
  INVX1   g14440(.A(n17820), .Y(n17833));
  AOI22X1 g14441(.A0(n17694), .A1(n17833), .B0(n17686), .B1(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .Y(n17834));
  OAI21X1 g14442(.A0(n16586), .A1(n14526), .B0(n17834), .Y(n17835));
  NOR2X1  g14443(.A(n17835), .B(n17832), .Y(n17836));
  OAI21X1 g14444(.A0(n17683), .A1(n16790), .B0(n17836), .Y(P1_U2993));
  NAND2X1 g14445(.A(n17682), .B(n16837), .Y(n17838));
  NOR2X1  g14446(.A(n16824), .B(n16823), .Y(n17839));
  NAND3X1 g14447(.A(n17747), .B(n17839), .C(n16818), .Y(n17840));
  INVX1   g14448(.A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .Y(n17841));
  NOR3X1  g14449(.A(n17795), .B(n17794), .C(n17818), .Y(n17842));
  XOR2X1  g14450(.A(n17842), .B(n17841), .Y(n17843));
  OAI22X1 g14451(.A0(n17725), .A1(n17841), .B0(n17663), .B1(n17843), .Y(n17844));
  AOI21X1 g14452(.A0(n17664), .A1(P1_EAX_REG_7__SCAN_IN), .B0(n17844), .Y(n17845));
  XOR2X1  g14453(.A(n17845), .B(n17662), .Y(n17846));
  XOR2X1  g14454(.A(n17846), .B(n17840), .Y(n17847));
  AOI21X1 g14455(.A0(n17826), .A1(n17817), .B0(n17829), .Y(n17848));
  XOR2X1  g14456(.A(n17848), .B(n17847), .Y(n17849));
  INVX1   g14457(.A(n17849), .Y(n17850));
  NAND2X1 g14458(.A(n17850), .B(n17687), .Y(n17851));
  NAND4X1 g14459(.A(n15093), .B(n15155), .C(P1_REIP_REG_7__SCAN_IN), .D(n17685), .Y(n17852));
  INVX1   g14460(.A(n17843), .Y(n17853));
  AOI22X1 g14461(.A0(n17694), .A1(n17853), .B0(n17686), .B1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .Y(n17854));
  NAND4X1 g14462(.A(n17852), .B(n17851), .C(n17838), .D(n17854), .Y(P1_U2992));
  INVX1   g14463(.A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .Y(n17856));
  NOR4X1  g14464(.A(n17794), .B(n17818), .C(n17841), .D(n17795), .Y(n17857));
  XOR2X1  g14465(.A(n17857), .B(n17856), .Y(n17858));
  OAI22X1 g14466(.A0(n17725), .A1(n17856), .B0(n17663), .B1(n17858), .Y(n17859));
  AOI21X1 g14467(.A0(n17664), .A1(P1_EAX_REG_8__SCAN_IN), .B0(n17859), .Y(n17860));
  XOR2X1  g14468(.A(n17860), .B(n17662), .Y(n17861));
  INVX1   g14469(.A(n17861), .Y(n17862));
  AOI21X1 g14470(.A0(n17747), .A1(n16901), .B0(n17862), .Y(n17863));
  NAND3X1 g14471(.A(n17862), .B(n17747), .C(n16901), .Y(n17864));
  INVX1   g14472(.A(n17864), .Y(n17865));
  NOR2X1  g14473(.A(n17865), .B(n17863), .Y(n17866));
  NAND2X1 g14474(.A(n17846), .B(n17840), .Y(n17867));
  NAND4X1 g14475(.A(n17826), .B(n17807), .C(n17802), .D(n17867), .Y(n17868));
  NOR2X1  g14476(.A(n17846), .B(n17840), .Y(n17869));
  AOI21X1 g14477(.A0(n17802), .A1(n17805), .B0(n17801), .Y(n17870));
  NAND2X1 g14478(.A(n17870), .B(n17827), .Y(n17871));
  AOI21X1 g14479(.A0(n17846), .A1(n17840), .B0(n17825), .Y(n17872));
  AOI21X1 g14480(.A0(n17872), .A1(n17871), .B0(n17869), .Y(n17873));
  NAND2X1 g14481(.A(n17873), .B(n17868), .Y(n17874));
  INVX1   g14482(.A(n17874), .Y(n17875));
  XOR2X1  g14483(.A(n17875), .B(n17866), .Y(n17876));
  NOR2X1  g14484(.A(n17876), .B(n17688), .Y(n17877));
  INVX1   g14485(.A(n17858), .Y(n17878));
  AOI22X1 g14486(.A0(n17694), .A1(n17878), .B0(n17686), .B1(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .Y(n17879));
  OAI21X1 g14487(.A0(n16586), .A1(n14520), .B0(n17879), .Y(n17880));
  NOR2X1  g14488(.A(n17880), .B(n17877), .Y(n17881));
  OAI21X1 g14489(.A0(n17683), .A1(n16904), .B0(n17881), .Y(P1_U2991));
  INVX1   g14490(.A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .Y(n17883));
  NAND2X1 g14491(.A(n17857), .B(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .Y(n17884));
  XOR2X1  g14492(.A(n17884), .B(n17883), .Y(n17885));
  INVX1   g14493(.A(P1_EAX_REG_9__SCAN_IN), .Y(n17886));
  OAI22X1 g14494(.A0(n17670), .A1(n17886), .B0(n17883), .B1(n17725), .Y(n17887));
  AOI21X1 g14495(.A0(n17885), .A1(n17662), .B0(n17887), .Y(n17888));
  XOR2X1  g14496(.A(n17888), .B(n17662), .Y(n17889));
  NOR3X1  g14497(.A(n17889), .B(n17667), .C(n16936), .Y(n17890));
  OAI21X1 g14498(.A0(n17667), .A1(n16936), .B0(n17889), .Y(n17891));
  INVX1   g14499(.A(n17891), .Y(n17892));
  NOR2X1  g14500(.A(n17892), .B(n17890), .Y(n17893));
  INVX1   g14501(.A(n17863), .Y(n17894));
  AOI21X1 g14502(.A0(n17874), .A1(n17894), .B0(n17865), .Y(n17895));
  XOR2X1  g14503(.A(n17895), .B(n17893), .Y(n17896));
  NOR2X1  g14504(.A(n17896), .B(n17688), .Y(n17897));
  AOI22X1 g14505(.A0(n17694), .A1(n17885), .B0(n17686), .B1(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .Y(n17898));
  OAI21X1 g14506(.A0(n16586), .A1(n14517), .B0(n17898), .Y(n17899));
  NOR2X1  g14507(.A(n17899), .B(n17897), .Y(n17900));
  OAI21X1 g14508(.A0(n17683), .A1(n16945), .B0(n17900), .Y(P1_U2990));
  INVX1   g14509(.A(n17890), .Y(n17902));
  OAI21X1 g14510(.A0(n17895), .A1(n17892), .B0(n17902), .Y(n17903));
  INVX1   g14511(.A(n17903), .Y(n17904));
  INVX1   g14512(.A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .Y(n17905));
  NAND3X1 g14513(.A(n17857), .B(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .C(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .Y(n17906));
  XOR2X1  g14514(.A(n17906), .B(n17905), .Y(n17907));
  INVX1   g14515(.A(P1_EAX_REG_10__SCAN_IN), .Y(n17908));
  OAI22X1 g14516(.A0(n17670), .A1(n17908), .B0(n17905), .B1(n17725), .Y(n17909));
  AOI21X1 g14517(.A0(n17907), .A1(n17662), .B0(n17909), .Y(n17910));
  XOR2X1  g14518(.A(n17910), .B(n17662), .Y(n17911));
  OAI21X1 g14519(.A0(n17667), .A1(n16983), .B0(n17911), .Y(n17912));
  INVX1   g14520(.A(n17912), .Y(n17913));
  NOR2X1  g14521(.A(n17913), .B(n17904), .Y(n17914));
  INVX1   g14522(.A(n17914), .Y(n17915));
  NOR3X1  g14523(.A(n17911), .B(n17667), .C(n16983), .Y(n17916));
  OAI21X1 g14524(.A0(n17916), .A1(n17913), .B0(n17904), .Y(n17917));
  OAI21X1 g14525(.A0(n17916), .A1(n17915), .B0(n17917), .Y(n17918));
  NOR2X1  g14526(.A(n17918), .B(n17688), .Y(n17919));
  AOI22X1 g14527(.A0(n17694), .A1(n17907), .B0(n17686), .B1(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .Y(n17920));
  OAI21X1 g14528(.A0(n16586), .A1(n14514), .B0(n17920), .Y(n17921));
  NOR2X1  g14529(.A(n17921), .B(n17919), .Y(n17922));
  OAI21X1 g14530(.A0(n17683), .A1(n16988), .B0(n17922), .Y(P1_U2989));
  INVX1   g14531(.A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .Y(n17924));
  NAND4X1 g14532(.A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .C(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .D(n17857), .Y(n17925));
  XOR2X1  g14533(.A(n17925), .B(n17924), .Y(n17926));
  INVX1   g14534(.A(P1_EAX_REG_11__SCAN_IN), .Y(n17927));
  OAI22X1 g14535(.A0(n17670), .A1(n17927), .B0(n17924), .B1(n17725), .Y(n17928));
  AOI21X1 g14536(.A0(n17926), .A1(n17662), .B0(n17928), .Y(n17929));
  XOR2X1  g14537(.A(n17929), .B(n17662), .Y(n17930));
  INVX1   g14538(.A(n17930), .Y(n17931));
  NOR2X1  g14539(.A(n17667), .B(n17023), .Y(n17932));
  XOR2X1  g14540(.A(n17932), .B(n17931), .Y(n17933));
  NOR2X1  g14541(.A(n17933), .B(n17916), .Y(n17934));
  INVX1   g14542(.A(n17916), .Y(n17935));
  OAI21X1 g14543(.A0(n17913), .A1(n17904), .B0(n17935), .Y(n17936));
  AOI22X1 g14544(.A0(n17934), .A1(n17915), .B0(n17933), .B1(n17936), .Y(n17937));
  AOI22X1 g14545(.A0(n17694), .A1(n17926), .B0(n17686), .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .Y(n17938));
  OAI21X1 g14546(.A0(n16586), .A1(n14511), .B0(n17938), .Y(n17939));
  AOI21X1 g14547(.A0(n17937), .A1(n17687), .B0(n17939), .Y(n17940));
  OAI21X1 g14548(.A0(n17683), .A1(n17035), .B0(n17940), .Y(P1_U2988));
  NOR2X1  g14549(.A(n17925), .B(n17924), .Y(n17942));
  XOR2X1  g14550(.A(n17942), .B(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .Y(n17943));
  INVX1   g14551(.A(P1_EAX_REG_12__SCAN_IN), .Y(n17944));
  INVX1   g14552(.A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .Y(n17945));
  OAI22X1 g14553(.A0(n17670), .A1(n17944), .B0(n17945), .B1(n17725), .Y(n17946));
  AOI21X1 g14554(.A0(n17943), .A1(n17662), .B0(n17946), .Y(n17947));
  XOR2X1  g14555(.A(n17947), .B(n17662), .Y(n17948));
  NOR3X1  g14556(.A(n17948), .B(n17667), .C(n17068), .Y(n17949));
  INVX1   g14557(.A(n17949), .Y(n17950));
  OAI21X1 g14558(.A0(n17667), .A1(n17068), .B0(n17948), .Y(n17951));
  NAND2X1 g14559(.A(n17951), .B(n17950), .Y(n17952));
  OAI21X1 g14560(.A0(n17667), .A1(n17023), .B0(n17930), .Y(n17953));
  NAND4X1 g14561(.A(n17912), .B(n17891), .C(n17894), .D(n17953), .Y(n17954));
  NOR3X1  g14562(.A(n17930), .B(n17667), .C(n17023), .Y(n17955));
  NOR3X1  g14563(.A(n17916), .B(n17890), .C(n17865), .Y(n17956));
  INVX1   g14564(.A(n17956), .Y(n17957));
  NAND2X1 g14565(.A(n17953), .B(n17912), .Y(n17958));
  AOI21X1 g14566(.A0(n17935), .A1(n17892), .B0(n17958), .Y(n17959));
  AOI21X1 g14567(.A0(n17959), .A1(n17957), .B0(n17955), .Y(n17960));
  OAI21X1 g14568(.A0(n17954), .A1(n17875), .B0(n17960), .Y(n17961));
  XOR2X1  g14569(.A(n17961), .B(n17952), .Y(n17962));
  NOR2X1  g14570(.A(n17962), .B(n17688), .Y(n17963));
  AOI22X1 g14571(.A0(n17694), .A1(n17943), .B0(n17686), .B1(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .Y(n17964));
  OAI21X1 g14572(.A0(n16586), .A1(n14508), .B0(n17964), .Y(n17965));
  NOR2X1  g14573(.A(n17965), .B(n17963), .Y(n17966));
  OAI21X1 g14574(.A0(n17683), .A1(n17077), .B0(n17966), .Y(P1_U2987));
  NOR3X1  g14575(.A(n17925), .B(n17924), .C(n17945), .Y(n17968));
  XOR2X1  g14576(.A(n17968), .B(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .Y(n17969));
  INVX1   g14577(.A(P1_EAX_REG_13__SCAN_IN), .Y(n17970));
  INVX1   g14578(.A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .Y(n17971));
  OAI22X1 g14579(.A0(n17670), .A1(n17970), .B0(n17971), .B1(n17725), .Y(n17972));
  AOI21X1 g14580(.A0(n17969), .A1(n17662), .B0(n17972), .Y(n17973));
  XOR2X1  g14581(.A(n17973), .B(n17662), .Y(n17974));
  NOR3X1  g14582(.A(n17974), .B(n17667), .C(n17110), .Y(n17975));
  OAI21X1 g14583(.A0(n17667), .A1(n17110), .B0(n17974), .Y(n17976));
  INVX1   g14584(.A(n17976), .Y(n17977));
  NOR2X1  g14585(.A(n17977), .B(n17975), .Y(n17978));
  AOI21X1 g14586(.A0(n17961), .A1(n17951), .B0(n17949), .Y(n17979));
  XOR2X1  g14587(.A(n17979), .B(n17978), .Y(n17980));
  NOR2X1  g14588(.A(n17980), .B(n17688), .Y(n17981));
  AOI22X1 g14589(.A0(n17694), .A1(n17969), .B0(n17686), .B1(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .Y(n17982));
  OAI21X1 g14590(.A0(n16586), .A1(n14505), .B0(n17982), .Y(n17983));
  NOR2X1  g14591(.A(n17983), .B(n17981), .Y(n17984));
  OAI21X1 g14592(.A0(n17683), .A1(n17115), .B0(n17984), .Y(P1_U2986));
  INVX1   g14593(.A(n17975), .Y(n17986));
  OAI21X1 g14594(.A0(n17979), .A1(n17977), .B0(n17986), .Y(n17987));
  INVX1   g14595(.A(n17987), .Y(n17988));
  INVX1   g14596(.A(n17153), .Y(n17989));
  NOR4X1  g14597(.A(n17924), .B(n17945), .C(n17971), .D(n17925), .Y(n17990));
  XOR2X1  g14598(.A(n17990), .B(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .Y(n17991));
  INVX1   g14599(.A(P1_EAX_REG_14__SCAN_IN), .Y(n17992));
  NAND3X1 g14600(.A(n15155), .B(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .C(P1_STATEBS16_REG_SCAN_IN), .Y(n17993));
  OAI21X1 g14601(.A0(n17670), .A1(n17992), .B0(n17993), .Y(n17994));
  AOI21X1 g14602(.A0(n17991), .A1(n17662), .B0(n17994), .Y(n17995));
  XOR2X1  g14603(.A(n17995), .B(n17662), .Y(n17996));
  INVX1   g14604(.A(n17996), .Y(n17997));
  AOI21X1 g14605(.A0(n17747), .A1(n17989), .B0(n17997), .Y(n17998));
  NOR2X1  g14606(.A(n17998), .B(n17988), .Y(n17999));
  INVX1   g14607(.A(n17999), .Y(n18000));
  NOR3X1  g14608(.A(n17996), .B(n17667), .C(n17153), .Y(n18001));
  OAI21X1 g14609(.A0(n18001), .A1(n17998), .B0(n17988), .Y(n18002));
  OAI21X1 g14610(.A0(n18001), .A1(n18000), .B0(n18002), .Y(n18003));
  NOR2X1  g14611(.A(n18003), .B(n17688), .Y(n18004));
  AOI22X1 g14612(.A0(n17694), .A1(n17991), .B0(n17686), .B1(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .Y(n18005));
  OAI21X1 g14613(.A0(n16586), .A1(n14502), .B0(n18005), .Y(n18006));
  NOR2X1  g14614(.A(n18006), .B(n18004), .Y(n18007));
  OAI21X1 g14615(.A0(n17683), .A1(n17158), .B0(n18007), .Y(P1_U2985));
  INVX1   g14616(.A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .Y(n18009));
  NAND2X1 g14617(.A(n17990), .B(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .Y(n18010));
  XOR2X1  g14618(.A(n18010), .B(n18009), .Y(n18011));
  INVX1   g14619(.A(P1_EAX_REG_15__SCAN_IN), .Y(n18012));
  OAI22X1 g14620(.A0(n17670), .A1(n18012), .B0(n18009), .B1(n17725), .Y(n18013));
  AOI21X1 g14621(.A0(n18011), .A1(n17662), .B0(n18013), .Y(n18014));
  XOR2X1  g14622(.A(n18014), .B(n17662), .Y(n18015));
  INVX1   g14623(.A(n18015), .Y(n18016));
  NOR2X1  g14624(.A(n17667), .B(n17189), .Y(n18017));
  XOR2X1  g14625(.A(n18017), .B(n18016), .Y(n18018));
  NOR2X1  g14626(.A(n18018), .B(n18001), .Y(n18019));
  NOR2X1  g14627(.A(n18017), .B(n18016), .Y(n18020));
  NOR3X1  g14628(.A(n18015), .B(n17667), .C(n17189), .Y(n18021));
  INVX1   g14629(.A(n17998), .Y(n18022));
  AOI21X1 g14630(.A0(n18022), .A1(n17987), .B0(n18001), .Y(n18023));
  NOR3X1  g14631(.A(n18023), .B(n18021), .C(n18020), .Y(n18024));
  AOI21X1 g14632(.A0(n18019), .A1(n18000), .B0(n18024), .Y(n18025));
  AOI22X1 g14633(.A0(n17694), .A1(n18011), .B0(n17686), .B1(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .Y(n18026));
  OAI21X1 g14634(.A0(n16586), .A1(n14499), .B0(n18026), .Y(n18027));
  AOI21X1 g14635(.A0(n18025), .A1(n17687), .B0(n18027), .Y(n18028));
  OAI21X1 g14636(.A0(n17683), .A1(n17200), .B0(n18028), .Y(P1_U2984));
  NAND3X1 g14637(.A(n17990), .B(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .C(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .Y(n18030));
  XOR2X1  g14638(.A(n18030), .B(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .Y(n18031));
  INVX1   g14639(.A(n18031), .Y(n18032));
  NOR3X1  g14640(.A(n15000), .B(n14985), .C(n15150), .Y(n18033));
  AOI21X1 g14641(.A0(n15010), .A1(P1_STATE2_REG_0__SCAN_IN), .B0(n18033), .Y(n18034));
  AOI22X1 g14642(.A0(n15362), .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B0(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(n15361), .Y(n18037));
  AOI22X1 g14643(.A0(n15359), .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B0(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(n14674), .Y(n18040));
  AOI22X1 g14644(.A0(n14673), .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B0(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(n15355), .Y(n18043));
  AOI22X1 g14645(.A0(n15372), .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B0(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(n14704), .Y(n18046));
  NAND4X1 g14646(.A(n18043), .B(n18040), .C(n18037), .D(n18046), .Y(n18047));
  AOI22X1 g14647(.A0(n15375), .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B0(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(n14671), .Y(n18050));
  AOI22X1 g14648(.A0(n15365), .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B0(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(n14703), .Y(n18053));
  AOI22X1 g14649(.A0(n14907), .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B0(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(n14680), .Y(n18056));
  AOI22X1 g14650(.A0(n15378), .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B0(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(n14682), .Y(n18059));
  NAND4X1 g14651(.A(n18056), .B(n18053), .C(n18050), .D(n18059), .Y(n18060));
  OAI21X1 g14652(.A0(n18060), .A1(n18047), .B0(n17747), .Y(n18061));
  AOI22X1 g14653(.A0(n17664), .A1(P1_EAX_REG_16__SCAN_IN), .B0(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(n17671), .Y(n18062));
  OAI21X1 g14654(.A0(n18061), .A1(n18034), .B0(n18062), .Y(n18063));
  AOI21X1 g14655(.A0(n18032), .A1(n17662), .B0(n18063), .Y(n18064));
  XOR2X1  g14656(.A(n18064), .B(n17662), .Y(n18065));
  NOR3X1  g14657(.A(n18065), .B(n17667), .C(n17230), .Y(n18066));
  OAI21X1 g14658(.A0(n17667), .A1(n17230), .B0(n18065), .Y(n18067));
  INVX1   g14659(.A(n18067), .Y(n18068));
  NOR2X1  g14660(.A(n18068), .B(n18066), .Y(n18069));
  INVX1   g14661(.A(n18020), .Y(n18070));
  NAND4X1 g14662(.A(n18022), .B(n17976), .C(n17951), .D(n18070), .Y(n18071));
  INVX1   g14663(.A(n18071), .Y(n18072));
  NAND2X1 g14664(.A(n18072), .B(n17961), .Y(n18073));
  NOR4X1  g14665(.A(n17998), .B(n17977), .C(n17950), .D(n18020), .Y(n18074));
  NOR4X1  g14666(.A(n17996), .B(n17667), .C(n17153), .D(n18020), .Y(n18075));
  NOR3X1  g14667(.A(n18020), .B(n17998), .C(n17986), .Y(n18076));
  NOR4X1  g14668(.A(n18075), .B(n18074), .C(n18021), .D(n18076), .Y(n18077));
  NAND2X1 g14669(.A(n18077), .B(n18073), .Y(n18078));
  INVX1   g14670(.A(n18078), .Y(n18079));
  XOR2X1  g14671(.A(n18079), .B(n18069), .Y(n18080));
  NOR2X1  g14672(.A(n18080), .B(n17688), .Y(n18081));
  AOI22X1 g14673(.A0(n17694), .A1(n18032), .B0(n17686), .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .Y(n18082));
  OAI21X1 g14674(.A0(n16586), .A1(n14496), .B0(n18082), .Y(n18083));
  NOR2X1  g14675(.A(n18083), .B(n18081), .Y(n18084));
  OAI21X1 g14676(.A0(n17683), .A1(n17233), .B0(n18084), .Y(P1_U2983));
  NOR3X1  g14677(.A(n17667), .B(n17257), .C(n16815), .Y(n18086));
  INVX1   g14678(.A(n18086), .Y(n18087));
  NAND4X1 g14679(.A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .C(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .D(n17990), .Y(n18088));
  XOR2X1  g14680(.A(n18088), .B(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .Y(n18089));
  INVX1   g14681(.A(n18089), .Y(n18090));
  AOI22X1 g14682(.A0(n15362), .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B0(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(n15361), .Y(n18091));
  AOI22X1 g14683(.A0(n15359), .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B0(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(n14674), .Y(n18092));
  AOI22X1 g14684(.A0(n14673), .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B0(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(n15355), .Y(n18093));
  AOI22X1 g14685(.A0(n15372), .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B0(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(n14704), .Y(n18094));
  NAND4X1 g14686(.A(n18093), .B(n18092), .C(n18091), .D(n18094), .Y(n18095));
  AOI22X1 g14687(.A0(n15375), .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B0(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(n14671), .Y(n18096));
  AOI22X1 g14688(.A0(n15365), .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B0(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(n14703), .Y(n18097));
  AOI22X1 g14689(.A0(n14907), .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B0(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(n14680), .Y(n18098));
  AOI22X1 g14690(.A0(n15378), .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B0(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(n14682), .Y(n18099));
  NAND4X1 g14691(.A(n18098), .B(n18097), .C(n18096), .D(n18099), .Y(n18100));
  OAI21X1 g14692(.A0(n18100), .A1(n18095), .B0(n17747), .Y(n18101));
  AOI22X1 g14693(.A0(n17664), .A1(P1_EAX_REG_17__SCAN_IN), .B0(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(n17671), .Y(n18102));
  OAI21X1 g14694(.A0(n18101), .A1(n18034), .B0(n18102), .Y(n18103));
  AOI21X1 g14695(.A0(n18090), .A1(n17662), .B0(n18103), .Y(n18104));
  XOR2X1  g14696(.A(n18104), .B(n17662), .Y(n18105));
  XOR2X1  g14697(.A(n18105), .B(n18087), .Y(n18106));
  AOI21X1 g14698(.A0(n18078), .A1(n18067), .B0(n18066), .Y(n18107));
  XOR2X1  g14699(.A(n18107), .B(n18106), .Y(n18108));
  NOR2X1  g14700(.A(n18108), .B(n17688), .Y(n18109));
  AOI22X1 g14701(.A0(n17694), .A1(n18090), .B0(n17686), .B1(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .Y(n18110));
  OAI21X1 g14702(.A0(n16586), .A1(n14493), .B0(n18110), .Y(n18111));
  NOR2X1  g14703(.A(n18111), .B(n18109), .Y(n18112));
  OAI21X1 g14704(.A0(n17683), .A1(n17260), .B0(n18112), .Y(P1_U2982));
  INVX1   g14705(.A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .Y(n18114));
  INVX1   g14706(.A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .Y(n18115));
  NOR2X1  g14707(.A(n18088), .B(n18115), .Y(n18116));
  XOR2X1  g14708(.A(n18116), .B(n18114), .Y(n18117));
  INVX1   g14709(.A(n18117), .Y(n18118));
  AOI22X1 g14710(.A0(n15362), .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B0(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(n15361), .Y(n18119));
  AOI22X1 g14711(.A0(n15359), .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B0(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(n14674), .Y(n18120));
  AOI22X1 g14712(.A0(n14673), .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B0(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(n15355), .Y(n18121));
  AOI22X1 g14713(.A0(n15372), .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B0(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(n14704), .Y(n18122));
  NAND4X1 g14714(.A(n18121), .B(n18120), .C(n18119), .D(n18122), .Y(n18123));
  AOI22X1 g14715(.A0(n15375), .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B0(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(n14671), .Y(n18124));
  AOI22X1 g14716(.A0(n15365), .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B0(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(n14703), .Y(n18125));
  AOI22X1 g14717(.A0(n14907), .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B0(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(n14680), .Y(n18126));
  AOI22X1 g14718(.A0(n15378), .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B0(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(n14682), .Y(n18127));
  NAND4X1 g14719(.A(n18126), .B(n18125), .C(n18124), .D(n18127), .Y(n18128));
  OAI21X1 g14720(.A0(n18128), .A1(n18123), .B0(n17747), .Y(n18129));
  AOI22X1 g14721(.A0(n17664), .A1(P1_EAX_REG_18__SCAN_IN), .B0(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(n17671), .Y(n18130));
  OAI21X1 g14722(.A0(n18129), .A1(n18034), .B0(n18130), .Y(n18131));
  AOI21X1 g14723(.A0(n18118), .A1(n17662), .B0(n18131), .Y(n18132));
  XOR2X1  g14724(.A(n18132), .B(n17662), .Y(n18133));
  XOR2X1  g14725(.A(n18133), .B(n18087), .Y(n18134));
  NOR4X1  g14726(.A(n17667), .B(n17257), .C(n16815), .D(n18105), .Y(n18135));
  NAND2X1 g14727(.A(n18105), .B(n18087), .Y(n18136));
  AOI21X1 g14728(.A0(n18136), .A1(n18066), .B0(n18135), .Y(n18137));
  AOI21X1 g14729(.A0(n18105), .A1(n18087), .B0(n18068), .Y(n18138));
  INVX1   g14730(.A(n18138), .Y(n18139));
  OAI21X1 g14731(.A0(n18139), .A1(n18079), .B0(n18137), .Y(n18140));
  XOR2X1  g14732(.A(n18140), .B(n18134), .Y(n18141));
  AOI22X1 g14733(.A0(n17694), .A1(n18118), .B0(n17686), .B1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .Y(n18142));
  OAI21X1 g14734(.A0(n16586), .A1(n14490), .B0(n18142), .Y(n18143));
  AOI21X1 g14735(.A0(n18141), .A1(n17687), .B0(n18143), .Y(n18144));
  OAI21X1 g14736(.A0(n17683), .A1(n17285), .B0(n18144), .Y(P1_U2981));
  INVX1   g14737(.A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .Y(n18146));
  NOR3X1  g14738(.A(n18088), .B(n18115), .C(n18114), .Y(n18147));
  XOR2X1  g14739(.A(n18147), .B(n18146), .Y(n18148));
  INVX1   g14740(.A(n18148), .Y(n18149));
  AOI22X1 g14741(.A0(n15362), .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B0(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(n15361), .Y(n18150));
  AOI22X1 g14742(.A0(n15359), .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B0(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(n14674), .Y(n18151));
  AOI22X1 g14743(.A0(n14673), .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B0(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(n15355), .Y(n18152));
  AOI22X1 g14744(.A0(n15372), .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B0(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(n14704), .Y(n18153));
  NAND4X1 g14745(.A(n18152), .B(n18151), .C(n18150), .D(n18153), .Y(n18154));
  AOI22X1 g14746(.A0(n15375), .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B0(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(n14671), .Y(n18155));
  AOI22X1 g14747(.A0(n15365), .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B0(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(n14703), .Y(n18156));
  AOI22X1 g14748(.A0(n14907), .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B0(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(n14680), .Y(n18157));
  AOI22X1 g14749(.A0(n15378), .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B0(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(n14682), .Y(n18158));
  NAND4X1 g14750(.A(n18157), .B(n18156), .C(n18155), .D(n18158), .Y(n18159));
  OAI21X1 g14751(.A0(n18159), .A1(n18154), .B0(n17747), .Y(n18160));
  AOI22X1 g14752(.A0(n17664), .A1(P1_EAX_REG_19__SCAN_IN), .B0(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(n17671), .Y(n18161));
  OAI21X1 g14753(.A0(n18160), .A1(n18034), .B0(n18161), .Y(n18162));
  AOI21X1 g14754(.A0(n18149), .A1(n17662), .B0(n18162), .Y(n18163));
  XOR2X1  g14755(.A(n18163), .B(n17662), .Y(n18164));
  XOR2X1  g14756(.A(n18164), .B(n18087), .Y(n18165));
  NAND2X1 g14757(.A(n18133), .B(n18087), .Y(n18166));
  INVX1   g14758(.A(n18166), .Y(n18167));
  NOR2X1  g14759(.A(n18139), .B(n18167), .Y(n18168));
  NOR4X1  g14760(.A(n17667), .B(n17257), .C(n16815), .D(n18133), .Y(n18169));
  INVX1   g14761(.A(n18169), .Y(n18170));
  OAI21X1 g14762(.A0(n18137), .A1(n18167), .B0(n18170), .Y(n18171));
  AOI21X1 g14763(.A0(n18168), .A1(n18078), .B0(n18171), .Y(n18172));
  XOR2X1  g14764(.A(n18172), .B(n18165), .Y(n18173));
  NOR2X1  g14765(.A(n18173), .B(n17688), .Y(n18174));
  AOI22X1 g14766(.A0(n17694), .A1(n18149), .B0(n17686), .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .Y(n18175));
  OAI21X1 g14767(.A0(n16586), .A1(n14487), .B0(n18175), .Y(n18176));
  NOR2X1  g14768(.A(n18176), .B(n18174), .Y(n18177));
  OAI21X1 g14769(.A0(n17683), .A1(n17311), .B0(n18177), .Y(P1_U2980));
  INVX1   g14770(.A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .Y(n18179));
  NOR4X1  g14771(.A(n18115), .B(n18114), .C(n18146), .D(n18088), .Y(n18180));
  XOR2X1  g14772(.A(n18180), .B(n18179), .Y(n18181));
  INVX1   g14773(.A(n18181), .Y(n18182));
  AOI22X1 g14774(.A0(n15362), .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B0(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(n15372), .Y(n18183));
  AOI22X1 g14775(.A0(n15361), .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B0(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(n14674), .Y(n18184));
  AOI22X1 g14776(.A0(n15359), .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B0(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(n14673), .Y(n18185));
  AOI22X1 g14777(.A0(n15355), .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B0(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(n14704), .Y(n18186));
  NAND4X1 g14778(.A(n18185), .B(n18184), .C(n18183), .D(n18186), .Y(n18187));
  AOI22X1 g14779(.A0(n15375), .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B0(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(n14671), .Y(n18188));
  AOI22X1 g14780(.A0(n15365), .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B0(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(n14703), .Y(n18189));
  AOI22X1 g14781(.A0(n14907), .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B0(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(n14680), .Y(n18190));
  AOI22X1 g14782(.A0(n15378), .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B0(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(n14682), .Y(n18191));
  NAND4X1 g14783(.A(n18190), .B(n18189), .C(n18188), .D(n18191), .Y(n18192));
  OAI21X1 g14784(.A0(n18192), .A1(n18187), .B0(n17747), .Y(n18193));
  AOI22X1 g14785(.A0(n17664), .A1(P1_EAX_REG_20__SCAN_IN), .B0(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B1(n17671), .Y(n18194));
  OAI21X1 g14786(.A0(n18193), .A1(n18034), .B0(n18194), .Y(n18195));
  AOI21X1 g14787(.A0(n18182), .A1(n17662), .B0(n18195), .Y(n18196));
  XOR2X1  g14788(.A(n18196), .B(n17662), .Y(n18197));
  XOR2X1  g14789(.A(n18197), .B(n18087), .Y(n18198));
  NOR4X1  g14790(.A(n17667), .B(n17257), .C(n16815), .D(n18164), .Y(n18199));
  AOI21X1 g14791(.A0(n18164), .A1(n18087), .B0(n18172), .Y(n18200));
  NOR2X1  g14792(.A(n18200), .B(n18199), .Y(n18201));
  XOR2X1  g14793(.A(n18201), .B(n18198), .Y(n18202));
  NOR2X1  g14794(.A(n18202), .B(n17688), .Y(n18203));
  AOI22X1 g14795(.A0(n17694), .A1(n18182), .B0(n17686), .B1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .Y(n18204));
  OAI21X1 g14796(.A0(n16586), .A1(n14484), .B0(n18204), .Y(n18205));
  NOR2X1  g14797(.A(n18205), .B(n18203), .Y(n18206));
  OAI21X1 g14798(.A0(n17683), .A1(n17332), .B0(n18206), .Y(P1_U2979));
  NAND2X1 g14799(.A(n18180), .B(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .Y(n18208));
  XOR2X1  g14800(.A(n18208), .B(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .Y(n18209));
  INVX1   g14801(.A(n18034), .Y(n18210));
  INVX1   g14802(.A(n15362), .Y(n18211));
  INVX1   g14803(.A(n15361), .Y(n18212));
  OAI22X1 g14804(.A0(n18211), .A1(n14792), .B0(n14794), .B1(n18212), .Y(n18213));
  INVX1   g14805(.A(n14674), .Y(n18215));
  OAI22X1 g14806(.A0(n14948), .A1(n14788), .B0(n14796), .B1(n18215), .Y(n18216));
  INVX1   g14807(.A(P1_INSTQUEUE_REG_3__5__SCAN_IN), .Y(n18217));
  OAI22X1 g14808(.A0(n14709), .A1(n18217), .B0(n14784), .B1(n14693), .Y(n18220));
  INVX1   g14809(.A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .Y(n18221));
  INVX1   g14810(.A(n14704), .Y(n18223));
  OAI22X1 g14811(.A0(n14692), .A1(n18221), .B0(n14786), .B1(n18223), .Y(n18224));
  NOR4X1  g14812(.A(n18220), .B(n18216), .C(n18213), .D(n18224), .Y(n18225));
  AOI22X1 g14813(.A0(n15375), .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B0(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(n14671), .Y(n18226));
  AOI22X1 g14814(.A0(n15365), .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B0(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(n14703), .Y(n18227));
  NAND2X1 g14815(.A(n18227), .B(n18226), .Y(n18228));
  AOI22X1 g14816(.A0(n14907), .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B0(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(n14680), .Y(n18229));
  AOI22X1 g14817(.A0(n15378), .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B0(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(n14682), .Y(n18230));
  NAND2X1 g14818(.A(n18230), .B(n18229), .Y(n18231));
  NOR2X1  g14819(.A(n18231), .B(n18228), .Y(n18232));
  AOI21X1 g14820(.A0(n18232), .A1(n18225), .B0(n17667), .Y(n18233));
  INVX1   g14821(.A(P1_EAX_REG_21__SCAN_IN), .Y(n18234));
  NAND3X1 g14822(.A(n15155), .B(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .C(P1_STATEBS16_REG_SCAN_IN), .Y(n18235));
  OAI21X1 g14823(.A0(n17670), .A1(n18234), .B0(n18235), .Y(n18236));
  AOI21X1 g14824(.A0(n18233), .A1(n18210), .B0(n18236), .Y(n18237));
  OAI21X1 g14825(.A0(n18209), .A1(n17663), .B0(n18237), .Y(n18238));
  XOR2X1  g14826(.A(n18238), .B(n17663), .Y(n18239));
  XOR2X1  g14827(.A(n18239), .B(n18087), .Y(n18240));
  INVX1   g14828(.A(n18172), .Y(n18241));
  AOI21X1 g14829(.A0(n18197), .A1(n18164), .B0(n18087), .Y(n18242));
  OAI21X1 g14830(.A0(n18197), .A1(n18164), .B0(n18087), .Y(n18243));
  AOI21X1 g14831(.A0(n18243), .A1(n18241), .B0(n18242), .Y(n18244));
  XOR2X1  g14832(.A(n18244), .B(n18240), .Y(n18245));
  NOR2X1  g14833(.A(n18245), .B(n17688), .Y(n18246));
  INVX1   g14834(.A(n18209), .Y(n18247));
  AOI22X1 g14835(.A0(n17694), .A1(n18247), .B0(n17686), .B1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .Y(n18248));
  OAI21X1 g14836(.A0(n16586), .A1(n14481), .B0(n18248), .Y(n18249));
  NOR2X1  g14837(.A(n18249), .B(n18246), .Y(n18250));
  OAI21X1 g14838(.A0(n17683), .A1(n17355), .B0(n18250), .Y(P1_U2978));
  NAND3X1 g14839(.A(n18180), .B(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .C(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .Y(n18252));
  XOR2X1  g14840(.A(n18252), .B(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .Y(n18253));
  NOR2X1  g14841(.A(n18253), .B(n17663), .Y(n18254));
  AOI22X1 g14842(.A0(n15362), .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B0(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(n15361), .Y(n18255));
  NAND2X1 g14843(.A(n15359), .B(P1_INSTQUEUE_REG_4__6__SCAN_IN), .Y(n18256));
  NAND2X1 g14844(.A(n14674), .B(P1_INSTQUEUE_REG_5__6__SCAN_IN), .Y(n18257));
  NAND3X1 g14845(.A(n18257), .B(n18256), .C(n18255), .Y(n18258));
  NAND2X1 g14846(.A(n14673), .B(P1_INSTQUEUE_REG_3__6__SCAN_IN), .Y(n18259));
  NAND2X1 g14847(.A(n15355), .B(P1_INSTQUEUE_REG_2__6__SCAN_IN), .Y(n18260));
  AOI22X1 g14848(.A0(n15372), .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B0(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(n14704), .Y(n18261));
  NAND3X1 g14849(.A(n18261), .B(n18260), .C(n18259), .Y(n18262));
  AOI22X1 g14850(.A0(n15375), .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B0(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(n14671), .Y(n18263));
  AOI22X1 g14851(.A0(n15365), .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B0(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(n14703), .Y(n18264));
  NAND2X1 g14852(.A(n18264), .B(n18263), .Y(n18265));
  AOI22X1 g14853(.A0(n14907), .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B0(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(n14680), .Y(n18266));
  AOI22X1 g14854(.A0(n15378), .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B0(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(n14682), .Y(n18267));
  NAND2X1 g14855(.A(n18267), .B(n18266), .Y(n18268));
  NOR4X1  g14856(.A(n18265), .B(n18262), .C(n18258), .D(n18268), .Y(n18269));
  NOR3X1  g14857(.A(n18269), .B(n18034), .C(n17667), .Y(n18270));
  INVX1   g14858(.A(P1_EAX_REG_22__SCAN_IN), .Y(n18271));
  NAND3X1 g14859(.A(n15155), .B(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .C(P1_STATEBS16_REG_SCAN_IN), .Y(n18272));
  OAI21X1 g14860(.A0(n17670), .A1(n18271), .B0(n18272), .Y(n18273));
  NOR3X1  g14861(.A(n18273), .B(n18270), .C(n18254), .Y(n18274));
  XOR2X1  g14862(.A(n18274), .B(n17662), .Y(n18275));
  XOR2X1  g14863(.A(n18275), .B(n18087), .Y(n18276));
  NAND2X1 g14864(.A(n18239), .B(n18087), .Y(n18277));
  NAND2X1 g14865(.A(n18242), .B(n18277), .Y(n18278));
  OAI21X1 g14866(.A0(n18239), .A1(n18087), .B0(n18278), .Y(n18279));
  NAND2X1 g14867(.A(n18243), .B(n18277), .Y(n18280));
  NOR2X1  g14868(.A(n18280), .B(n18172), .Y(n18281));
  NOR2X1  g14869(.A(n18281), .B(n18279), .Y(n18282));
  XOR2X1  g14870(.A(n18282), .B(n18276), .Y(n18283));
  NOR2X1  g14871(.A(n18283), .B(n17688), .Y(n18284));
  INVX1   g14872(.A(n18253), .Y(n18285));
  AOI22X1 g14873(.A0(n17694), .A1(n18285), .B0(n17686), .B1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .Y(n18286));
  OAI21X1 g14874(.A0(n16586), .A1(n14478), .B0(n18286), .Y(n18287));
  NOR2X1  g14875(.A(n18287), .B(n18284), .Y(n18288));
  OAI21X1 g14876(.A0(n17683), .A1(n17381), .B0(n18288), .Y(P1_U2977));
  INVX1   g14877(.A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .Y(n18290));
  NAND4X1 g14878(.A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .C(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .D(n18180), .Y(n18291));
  XOR2X1  g14879(.A(n18291), .B(n18290), .Y(n18292));
  NAND2X1 g14880(.A(n18292), .B(n17662), .Y(n18293));
  AOI22X1 g14881(.A0(n14671), .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B0(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(n14703), .Y(n18296));
  AOI22X1 g14882(.A0(n15362), .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B0(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(n15365), .Y(n18299));
  NAND2X1 g14883(.A(n18299), .B(n18296), .Y(n18300));
  AOI22X1 g14884(.A0(n14907), .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B0(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(n14704), .Y(n18303));
  AOI22X1 g14885(.A0(n15372), .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B0(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(n15355), .Y(n18306));
  NAND2X1 g14886(.A(n18306), .B(n18303), .Y(n18307));
  AOI22X1 g14887(.A0(n14680), .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B0(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(n14674), .Y(n18310));
  AOI22X1 g14888(.A0(n15359), .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B0(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(n15361), .Y(n18313));
  AOI22X1 g14889(.A0(n14682), .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B0(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(n14673), .Y(n18316));
  AOI22X1 g14890(.A0(n15375), .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B0(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(n15378), .Y(n18319));
  NAND4X1 g14891(.A(n18316), .B(n18313), .C(n18310), .D(n18319), .Y(n18320));
  NOR3X1  g14892(.A(n18320), .B(n18307), .C(n18300), .Y(n18321));
  AOI22X1 g14893(.A0(n15362), .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B0(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(n15361), .Y(n18322));
  AOI22X1 g14894(.A0(n15359), .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B0(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(n14674), .Y(n18323));
  AOI22X1 g14895(.A0(n14673), .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B0(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(n15355), .Y(n18324));
  AOI22X1 g14896(.A0(n15372), .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B0(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(n14704), .Y(n18325));
  NAND4X1 g14897(.A(n18324), .B(n18323), .C(n18322), .D(n18325), .Y(n18326));
  AOI22X1 g14898(.A0(n15375), .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B0(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(n14671), .Y(n18327));
  AOI22X1 g14899(.A0(n15365), .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B0(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(n14703), .Y(n18328));
  AOI22X1 g14900(.A0(n14907), .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B0(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(n14680), .Y(n18329));
  AOI22X1 g14901(.A0(n15378), .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B0(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(n14682), .Y(n18330));
  NAND4X1 g14902(.A(n18329), .B(n18328), .C(n18327), .D(n18330), .Y(n18331));
  OAI21X1 g14903(.A0(n18331), .A1(n18326), .B0(n18210), .Y(n18332));
  OAI21X1 g14904(.A0(n18321), .A1(n18034), .B0(n18332), .Y(n18333));
  NOR3X1  g14905(.A(n18332), .B(n18321), .C(n18034), .Y(n18334));
  NOR2X1  g14906(.A(n18334), .B(n17667), .Y(n18335));
  INVX1   g14907(.A(P1_EAX_REG_23__SCAN_IN), .Y(n18336));
  OAI22X1 g14908(.A0(n17670), .A1(n18336), .B0(n18290), .B1(n17725), .Y(n18337));
  AOI21X1 g14909(.A0(n18335), .A1(n18333), .B0(n18337), .Y(n18338));
  NAND2X1 g14910(.A(n18338), .B(n18293), .Y(n18339));
  XOR2X1  g14911(.A(n18339), .B(n17663), .Y(n18340));
  XOR2X1  g14912(.A(n18340), .B(n18087), .Y(n18341));
  NAND2X1 g14913(.A(n18275), .B(n18087), .Y(n18342));
  NAND3X1 g14914(.A(n18342), .B(n18243), .C(n18277), .Y(n18343));
  NOR4X1  g14915(.A(n17667), .B(n17257), .C(n16815), .D(n18275), .Y(n18344));
  AOI21X1 g14916(.A0(n18279), .A1(n18342), .B0(n18344), .Y(n18345));
  OAI21X1 g14917(.A0(n18343), .A1(n18172), .B0(n18345), .Y(n18346));
  INVX1   g14918(.A(n18346), .Y(n18347));
  XOR2X1  g14919(.A(n18347), .B(n18341), .Y(n18348));
  NOR2X1  g14920(.A(n18348), .B(n17688), .Y(n18349));
  AOI22X1 g14921(.A0(n17694), .A1(n18292), .B0(n17686), .B1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .Y(n18350));
  OAI21X1 g14922(.A0(n16586), .A1(n14475), .B0(n18350), .Y(n18351));
  NOR2X1  g14923(.A(n18351), .B(n18349), .Y(n18352));
  OAI21X1 g14924(.A0(n17683), .A1(n17411), .B0(n18352), .Y(P1_U2976));
  INVX1   g14925(.A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .Y(n18354));
  NOR2X1  g14926(.A(n18291), .B(n18290), .Y(n18355));
  XOR2X1  g14927(.A(n18355), .B(n18354), .Y(n18356));
  AOI22X1 g14928(.A0(n14671), .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B0(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(n14703), .Y(n18357));
  AOI22X1 g14929(.A0(n15362), .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B0(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(n15365), .Y(n18358));
  NAND2X1 g14930(.A(n18358), .B(n18357), .Y(n18359));
  AOI22X1 g14931(.A0(n14907), .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B0(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(n14704), .Y(n18360));
  AOI22X1 g14932(.A0(n15372), .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B0(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(n15355), .Y(n18361));
  NAND2X1 g14933(.A(n18361), .B(n18360), .Y(n18362));
  AOI22X1 g14934(.A0(n14680), .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B0(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(n14674), .Y(n18363));
  AOI22X1 g14935(.A0(n15359), .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B0(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(n15361), .Y(n18364));
  AOI22X1 g14936(.A0(n14682), .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B0(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(n14673), .Y(n18365));
  AOI22X1 g14937(.A0(n15375), .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B0(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(n15378), .Y(n18366));
  NAND4X1 g14938(.A(n18365), .B(n18364), .C(n18363), .D(n18366), .Y(n18367));
  NOR3X1  g14939(.A(n18367), .B(n18362), .C(n18359), .Y(n18368));
  NOR2X1  g14940(.A(n18368), .B(n18034), .Y(n18369));
  XOR2X1  g14941(.A(n18369), .B(n18334), .Y(n18370));
  INVX1   g14942(.A(P1_EAX_REG_24__SCAN_IN), .Y(n18371));
  OAI22X1 g14943(.A0(n17670), .A1(n18371), .B0(n18354), .B1(n17725), .Y(n18372));
  AOI21X1 g14944(.A0(n18370), .A1(n17747), .B0(n18372), .Y(n18373));
  OAI21X1 g14945(.A0(n18356), .A1(n17663), .B0(n18373), .Y(n18374));
  XOR2X1  g14946(.A(n18374), .B(n17663), .Y(n18375));
  XOR2X1  g14947(.A(n18375), .B(n18087), .Y(n18376));
  NOR4X1  g14948(.A(n17667), .B(n17257), .C(n16815), .D(n18340), .Y(n18377));
  NAND2X1 g14949(.A(n18340), .B(n18087), .Y(n18378));
  AOI21X1 g14950(.A0(n18346), .A1(n18378), .B0(n18377), .Y(n18379));
  XOR2X1  g14951(.A(n18379), .B(n18376), .Y(n18380));
  NOR2X1  g14952(.A(n18380), .B(n17688), .Y(n18381));
  INVX1   g14953(.A(n18356), .Y(n18382));
  AOI22X1 g14954(.A0(n17694), .A1(n18382), .B0(n17686), .B1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .Y(n18383));
  OAI21X1 g14955(.A0(n16586), .A1(n14472), .B0(n18383), .Y(n18384));
  NOR2X1  g14956(.A(n18384), .B(n18381), .Y(n18385));
  OAI21X1 g14957(.A0(n17683), .A1(n17433), .B0(n18385), .Y(P1_U2975));
  NOR3X1  g14958(.A(n18291), .B(n18290), .C(n18354), .Y(n18387));
  XOR2X1  g14959(.A(n18387), .B(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .Y(n18388));
  NAND2X1 g14960(.A(n18369), .B(n18334), .Y(n18389));
  AOI22X1 g14961(.A0(n14671), .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B0(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(n14703), .Y(n18390));
  AOI22X1 g14962(.A0(n15362), .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B0(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(n15365), .Y(n18391));
  NAND2X1 g14963(.A(n18391), .B(n18390), .Y(n18392));
  AOI22X1 g14964(.A0(n14907), .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B0(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(n14704), .Y(n18393));
  AOI22X1 g14965(.A0(n15372), .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B0(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(n15355), .Y(n18394));
  NAND2X1 g14966(.A(n18394), .B(n18393), .Y(n18395));
  AOI22X1 g14967(.A0(n14680), .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B0(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(n14674), .Y(n18396));
  AOI22X1 g14968(.A0(n15359), .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B0(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(n15361), .Y(n18397));
  AOI22X1 g14969(.A0(n14682), .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B0(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(n14673), .Y(n18398));
  AOI22X1 g14970(.A0(n15375), .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B0(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(n15378), .Y(n18399));
  NAND4X1 g14971(.A(n18398), .B(n18397), .C(n18396), .D(n18399), .Y(n18400));
  NOR3X1  g14972(.A(n18400), .B(n18395), .C(n18392), .Y(n18401));
  NOR2X1  g14973(.A(n18401), .B(n18034), .Y(n18402));
  XOR2X1  g14974(.A(n18402), .B(n18389), .Y(n18403));
  AOI22X1 g14975(.A0(n17664), .A1(P1_EAX_REG_25__SCAN_IN), .B0(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B1(n17671), .Y(n18404));
  OAI21X1 g14976(.A0(n18403), .A1(n17667), .B0(n18404), .Y(n18405));
  AOI21X1 g14977(.A0(n18388), .A1(n17662), .B0(n18405), .Y(n18406));
  XOR2X1  g14978(.A(n18406), .B(n17662), .Y(n18407));
  XOR2X1  g14979(.A(n18407), .B(n18087), .Y(n18408));
  AOI21X1 g14980(.A0(n18375), .A1(n18340), .B0(n18087), .Y(n18409));
  OAI21X1 g14981(.A0(n18375), .A1(n18340), .B0(n18087), .Y(n18410));
  AOI21X1 g14982(.A0(n18410), .A1(n18346), .B0(n18409), .Y(n18411));
  XOR2X1  g14983(.A(n18411), .B(n18408), .Y(n18412));
  NOR2X1  g14984(.A(n18412), .B(n17688), .Y(n18413));
  AOI22X1 g14985(.A0(n17694), .A1(n18388), .B0(n17686), .B1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .Y(n18414));
  OAI21X1 g14986(.A0(n16586), .A1(n14469), .B0(n18414), .Y(n18415));
  NOR2X1  g14987(.A(n18415), .B(n18413), .Y(n18416));
  OAI21X1 g14988(.A0(n17683), .A1(n17456), .B0(n18416), .Y(P1_U2974));
  NAND2X1 g14989(.A(n17682), .B(n17481), .Y(n18418));
  INVX1   g14990(.A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .Y(n18419));
  NOR4X1  g14991(.A(n18290), .B(n18354), .C(n18419), .D(n18291), .Y(n18420));
  XOR2X1  g14992(.A(n18420), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .Y(n18421));
  AOI22X1 g14993(.A0(n14671), .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B0(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(n14703), .Y(n18422));
  AOI22X1 g14994(.A0(n15362), .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B0(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(n15365), .Y(n18423));
  NAND2X1 g14995(.A(n18423), .B(n18422), .Y(n18424));
  AOI22X1 g14996(.A0(n14907), .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B0(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(n14704), .Y(n18425));
  AOI22X1 g14997(.A0(n15372), .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B0(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(n15355), .Y(n18426));
  NAND2X1 g14998(.A(n18426), .B(n18425), .Y(n18427));
  AOI22X1 g14999(.A0(n14680), .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B0(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(n14674), .Y(n18428));
  AOI22X1 g15000(.A0(n15359), .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B0(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(n15361), .Y(n18429));
  AOI22X1 g15001(.A0(n14682), .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B0(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(n14673), .Y(n18430));
  AOI22X1 g15002(.A0(n15375), .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B0(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(n15378), .Y(n18431));
  NAND4X1 g15003(.A(n18430), .B(n18429), .C(n18428), .D(n18431), .Y(n18432));
  NOR3X1  g15004(.A(n18432), .B(n18427), .C(n18424), .Y(n18433));
  NOR2X1  g15005(.A(n18433), .B(n18034), .Y(n18434));
  NAND3X1 g15006(.A(n18402), .B(n18369), .C(n18334), .Y(n18435));
  XOR2X1  g15007(.A(n18435), .B(n18434), .Y(n18436));
  AOI22X1 g15008(.A0(n17664), .A1(P1_EAX_REG_26__SCAN_IN), .B0(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B1(n17671), .Y(n18437));
  OAI21X1 g15009(.A0(n18436), .A1(n17667), .B0(n18437), .Y(n18438));
  AOI21X1 g15010(.A0(n18421), .A1(n17662), .B0(n18438), .Y(n18439));
  XOR2X1  g15011(.A(n18439), .B(n17662), .Y(n18440));
  XOR2X1  g15012(.A(n18440), .B(n18087), .Y(n18441));
  NOR4X1  g15013(.A(n17667), .B(n17257), .C(n16815), .D(n18407), .Y(n18442));
  NAND2X1 g15014(.A(n18407), .B(n18087), .Y(n18443));
  AOI21X1 g15015(.A0(n18409), .A1(n18443), .B0(n18442), .Y(n18444));
  INVX1   g15016(.A(n18444), .Y(n18445));
  NAND2X1 g15017(.A(n18410), .B(n18443), .Y(n18446));
  INVX1   g15018(.A(n18446), .Y(n18447));
  AOI21X1 g15019(.A0(n18447), .A1(n18346), .B0(n18445), .Y(n18448));
  XOR2X1  g15020(.A(n18448), .B(n18441), .Y(n18449));
  INVX1   g15021(.A(n18449), .Y(n18450));
  NAND2X1 g15022(.A(n18450), .B(n17687), .Y(n18451));
  NAND4X1 g15023(.A(n15093), .B(n15155), .C(P1_REIP_REG_26__SCAN_IN), .D(n17685), .Y(n18452));
  AOI22X1 g15024(.A0(n17694), .A1(n18421), .B0(n17686), .B1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .Y(n18453));
  NAND4X1 g15025(.A(n18452), .B(n18451), .C(n18418), .D(n18453), .Y(P1_U2973));
  NAND2X1 g15026(.A(n17682), .B(n17506), .Y(n18455));
  NAND2X1 g15027(.A(n18420), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .Y(n18456));
  XOR2X1  g15028(.A(n18456), .B(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .Y(n18457));
  INVX1   g15029(.A(n18457), .Y(n18458));
  NAND4X1 g15030(.A(n18402), .B(n18369), .C(n18334), .D(n18434), .Y(n18459));
  AOI22X1 g15031(.A0(n14671), .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B0(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(n14703), .Y(n18460));
  AOI22X1 g15032(.A0(n15362), .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B0(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(n15365), .Y(n18461));
  NAND2X1 g15033(.A(n18461), .B(n18460), .Y(n18462));
  AOI22X1 g15034(.A0(n14907), .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B0(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(n15355), .Y(n18463));
  AOI22X1 g15035(.A0(n14704), .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B0(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(n15372), .Y(n18464));
  NAND2X1 g15036(.A(n18464), .B(n18463), .Y(n18465));
  AOI22X1 g15037(.A0(n15361), .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B0(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(n15378), .Y(n18466));
  AOI22X1 g15038(.A0(n14680), .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B0(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(n15359), .Y(n18467));
  AOI22X1 g15039(.A0(n14674), .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B0(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(n14682), .Y(n18468));
  AOI22X1 g15040(.A0(n14673), .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B0(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(n15375), .Y(n18469));
  NAND4X1 g15041(.A(n18468), .B(n18467), .C(n18466), .D(n18469), .Y(n18470));
  NOR3X1  g15042(.A(n18470), .B(n18465), .C(n18462), .Y(n18471));
  NOR2X1  g15043(.A(n18471), .B(n18034), .Y(n18472));
  XOR2X1  g15044(.A(n18472), .B(n18459), .Y(n18473));
  AOI22X1 g15045(.A0(n17664), .A1(P1_EAX_REG_27__SCAN_IN), .B0(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B1(n17671), .Y(n18474));
  OAI21X1 g15046(.A0(n18473), .A1(n17667), .B0(n18474), .Y(n18475));
  AOI21X1 g15047(.A0(n18458), .A1(n17662), .B0(n18475), .Y(n18476));
  XOR2X1  g15048(.A(n18476), .B(n17662), .Y(n18477));
  XOR2X1  g15049(.A(n18477), .B(n18087), .Y(n18478));
  NOR4X1  g15050(.A(n17667), .B(n17257), .C(n16815), .D(n18440), .Y(n18479));
  NOR2X1  g15051(.A(n18445), .B(n18479), .Y(n18481));
  AOI21X1 g15052(.A0(n18440), .A1(n18087), .B0(n18446), .Y(n18482));
  INVX1   g15053(.A(n18482), .Y(n18483));
  OAI21X1 g15054(.A0(n18483), .A1(n18347), .B0(n18481), .Y(n18484));
  XOR2X1  g15055(.A(n18484), .B(n18478), .Y(n18485));
  NAND2X1 g15056(.A(n18485), .B(n17687), .Y(n18486));
  NAND4X1 g15057(.A(n15093), .B(n15155), .C(P1_REIP_REG_27__SCAN_IN), .D(n17685), .Y(n18487));
  AOI22X1 g15058(.A0(n17694), .A1(n18458), .B0(n17686), .B1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .Y(n18488));
  NAND4X1 g15059(.A(n18487), .B(n18486), .C(n18455), .D(n18488), .Y(P1_U2972));
  NAND3X1 g15060(.A(n18420), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .C(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .Y(n18490));
  XOR2X1  g15061(.A(n18490), .B(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .Y(n18491));
  INVX1   g15062(.A(n18491), .Y(n18492));
  NAND2X1 g15063(.A(n18492), .B(n17662), .Y(n18493));
  AOI22X1 g15064(.A0(n14671), .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B0(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(n14703), .Y(n18494));
  AOI22X1 g15065(.A0(n15362), .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B0(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(n15365), .Y(n18495));
  NAND2X1 g15066(.A(n18495), .B(n18494), .Y(n18496));
  NAND4X1 g15067(.A(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .D(n14678), .Y(n18497));
  NAND2X1 g15068(.A(n14704), .B(P1_INSTQUEUE_REG_2__5__SCAN_IN), .Y(n18498));
  AOI22X1 g15069(.A0(n15372), .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B0(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(n15355), .Y(n18499));
  NAND3X1 g15070(.A(n18499), .B(n18498), .C(n18497), .Y(n18500));
  AOI22X1 g15071(.A0(n14680), .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B0(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(n14674), .Y(n18501));
  AOI22X1 g15072(.A0(n15359), .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B0(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(n15361), .Y(n18502));
  AOI22X1 g15073(.A0(n14682), .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B0(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(n14673), .Y(n18503));
  AOI22X1 g15074(.A0(n15375), .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B0(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(n15378), .Y(n18504));
  NAND4X1 g15075(.A(n18503), .B(n18502), .C(n18501), .D(n18504), .Y(n18505));
  NOR3X1  g15076(.A(n18505), .B(n18500), .C(n18496), .Y(n18506));
  NOR2X1  g15077(.A(n18506), .B(n18034), .Y(n18507));
  NOR4X1  g15078(.A(n18435), .B(n18433), .C(n18034), .D(n18471), .Y(n18508));
  XOR2X1  g15079(.A(n18508), .B(n18507), .Y(n18509));
  NAND2X1 g15080(.A(n18509), .B(n17747), .Y(n18510));
  AOI22X1 g15081(.A0(n17664), .A1(P1_EAX_REG_28__SCAN_IN), .B0(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B1(n17671), .Y(n18511));
  NAND3X1 g15082(.A(n18511), .B(n18510), .C(n18493), .Y(n18512));
  XOR2X1  g15083(.A(n18512), .B(n17663), .Y(n18513));
  XOR2X1  g15084(.A(n18513), .B(n18087), .Y(n18514));
  NAND2X1 g15085(.A(n18477), .B(n18087), .Y(n18515));
  INVX1   g15086(.A(n18515), .Y(n18516));
  NOR2X1  g15087(.A(n18483), .B(n18516), .Y(n18517));
  NOR4X1  g15088(.A(n17667), .B(n17257), .C(n16815), .D(n18477), .Y(n18518));
  NOR2X1  g15089(.A(n18481), .B(n18516), .Y(n18519));
  NOR2X1  g15090(.A(n18519), .B(n18518), .Y(n18520));
  INVX1   g15091(.A(n18520), .Y(n18521));
  AOI21X1 g15092(.A0(n18517), .A1(n18346), .B0(n18521), .Y(n18522));
  XOR2X1  g15093(.A(n18522), .B(n18514), .Y(n18523));
  NOR2X1  g15094(.A(n18523), .B(n17688), .Y(n18524));
  AOI22X1 g15095(.A0(n17694), .A1(n18492), .B0(n17686), .B1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .Y(n18525));
  OAI21X1 g15096(.A0(n16586), .A1(n14460), .B0(n18525), .Y(n18526));
  NOR2X1  g15097(.A(n18526), .B(n18524), .Y(n18527));
  OAI21X1 g15098(.A0(n17683), .A1(n17533), .B0(n18527), .Y(P1_U2971));
  NAND4X1 g15099(.A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .C(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .D(n18420), .Y(n18529));
  XOR2X1  g15100(.A(n18529), .B(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .Y(n18530));
  INVX1   g15101(.A(n18530), .Y(n18531));
  NAND2X1 g15102(.A(n18508), .B(n18507), .Y(n18532));
  AOI22X1 g15103(.A0(n14671), .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B0(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(n14703), .Y(n18533));
  AOI22X1 g15104(.A0(n15362), .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B0(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(n15365), .Y(n18534));
  NAND2X1 g15105(.A(n18534), .B(n18533), .Y(n18535));
  AOI22X1 g15106(.A0(n14907), .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B0(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(n14704), .Y(n18536));
  AOI22X1 g15107(.A0(n15372), .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B0(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(n15355), .Y(n18537));
  NAND2X1 g15108(.A(n18537), .B(n18536), .Y(n18538));
  AOI22X1 g15109(.A0(n14680), .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B0(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(n14674), .Y(n18539));
  AOI22X1 g15110(.A0(n15359), .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B0(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(n15361), .Y(n18540));
  AOI22X1 g15111(.A0(n14682), .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B0(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(n14673), .Y(n18541));
  AOI22X1 g15112(.A0(n15375), .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B0(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(n15378), .Y(n18542));
  NAND4X1 g15113(.A(n18541), .B(n18540), .C(n18539), .D(n18542), .Y(n18543));
  NOR3X1  g15114(.A(n18543), .B(n18538), .C(n18535), .Y(n18544));
  NOR2X1  g15115(.A(n18544), .B(n18034), .Y(n18545));
  XOR2X1  g15116(.A(n18545), .B(n18532), .Y(n18546));
  AOI22X1 g15117(.A0(n17664), .A1(P1_EAX_REG_29__SCAN_IN), .B0(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B1(n17671), .Y(n18547));
  OAI21X1 g15118(.A0(n18546), .A1(n17667), .B0(n18547), .Y(n18548));
  AOI21X1 g15119(.A0(n18531), .A1(n17662), .B0(n18548), .Y(n18549));
  XOR2X1  g15120(.A(n18549), .B(n17662), .Y(n18550));
  XOR2X1  g15121(.A(n18550), .B(n18087), .Y(n18551));
  NOR4X1  g15122(.A(n17667), .B(n17257), .C(n16815), .D(n18513), .Y(n18552));
  AOI21X1 g15123(.A0(n18513), .A1(n18087), .B0(n18522), .Y(n18553));
  NOR2X1  g15124(.A(n18553), .B(n18552), .Y(n18554));
  XOR2X1  g15125(.A(n18554), .B(n18551), .Y(n18555));
  NOR2X1  g15126(.A(n17683), .B(n17575), .Y(n18556));
  AOI22X1 g15127(.A0(n17694), .A1(n18531), .B0(n17686), .B1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .Y(n18557));
  OAI21X1 g15128(.A0(n16586), .A1(n14457), .B0(n18557), .Y(n18558));
  NOR2X1  g15129(.A(n18558), .B(n18556), .Y(n18559));
  OAI21X1 g15130(.A0(n18555), .A1(n17688), .B0(n18559), .Y(P1_U2970));
  NAND2X1 g15131(.A(n18550), .B(n18087), .Y(n18561));
  OAI21X1 g15132(.A0(n18553), .A1(n18552), .B0(n18561), .Y(n18562));
  OAI21X1 g15133(.A0(n18550), .A1(n18087), .B0(n18562), .Y(n18563));
  INVX1   g15134(.A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .Y(n18564));
  INVX1   g15135(.A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .Y(n18565));
  NOR2X1  g15136(.A(n18529), .B(n18565), .Y(n18566));
  XOR2X1  g15137(.A(n18566), .B(n18564), .Y(n18567));
  NAND3X1 g15138(.A(n18545), .B(n18508), .C(n18507), .Y(n18568));
  AOI22X1 g15139(.A0(n14671), .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B0(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(n14703), .Y(n18569));
  AOI22X1 g15140(.A0(n15362), .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B0(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(n15365), .Y(n18570));
  NAND4X1 g15141(.A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .D(n14678), .Y(n18571));
  NAND2X1 g15142(.A(n14704), .B(P1_INSTQUEUE_REG_2__7__SCAN_IN), .Y(n18572));
  NAND2X1 g15143(.A(n15372), .B(P1_INSTQUEUE_REG_1__7__SCAN_IN), .Y(n18573));
  NAND2X1 g15144(.A(n15355), .B(P1_INSTQUEUE_REG_3__7__SCAN_IN), .Y(n18574));
  NAND4X1 g15145(.A(n18573), .B(n18572), .C(n18571), .D(n18574), .Y(n18575));
  AOI22X1 g15146(.A0(n14680), .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B0(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(n14674), .Y(n18576));
  AOI22X1 g15147(.A0(n15359), .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B0(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(n15361), .Y(n18577));
  AOI22X1 g15148(.A0(n14682), .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B0(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(n14673), .Y(n18578));
  AOI22X1 g15149(.A0(n15375), .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B0(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(n15378), .Y(n18579));
  NAND4X1 g15150(.A(n18578), .B(n18577), .C(n18576), .D(n18579), .Y(n18580));
  NOR2X1  g15151(.A(n18580), .B(n18575), .Y(n18581));
  NAND3X1 g15152(.A(n18581), .B(n18570), .C(n18569), .Y(n18582));
  NAND2X1 g15153(.A(n18582), .B(n18210), .Y(n18583));
  XOR2X1  g15154(.A(n18583), .B(n18568), .Y(n18584));
  INVX1   g15155(.A(P1_EAX_REG_30__SCAN_IN), .Y(n18585));
  OAI22X1 g15156(.A0(n17670), .A1(n18585), .B0(n18564), .B1(n17725), .Y(n18586));
  AOI21X1 g15157(.A0(n18584), .A1(n17747), .B0(n18586), .Y(n18587));
  OAI21X1 g15158(.A0(n18567), .A1(n17663), .B0(n18587), .Y(n18588));
  XOR2X1  g15159(.A(n18588), .B(n17663), .Y(n18589));
  XOR2X1  g15160(.A(n18589), .B(n18086), .Y(n18590));
  XOR2X1  g15161(.A(n18590), .B(n18563), .Y(n18591));
  NOR2X1  g15162(.A(n17683), .B(n17604), .Y(n18592));
  INVX1   g15163(.A(n18567), .Y(n18593));
  AOI22X1 g15164(.A0(n17694), .A1(n18593), .B0(n17686), .B1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .Y(n18594));
  OAI21X1 g15165(.A0(n16586), .A1(n14452), .B0(n18594), .Y(n18595));
  NOR2X1  g15166(.A(n18595), .B(n18592), .Y(n18596));
  OAI21X1 g15167(.A0(n18591), .A1(n17688), .B0(n18596), .Y(P1_U2969));
  INVX1   g15168(.A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .Y(n18598));
  NOR3X1  g15169(.A(n18529), .B(n18565), .C(n18564), .Y(n18599));
  XOR2X1  g15170(.A(n18599), .B(n18598), .Y(n18600));
  INVX1   g15171(.A(n18600), .Y(n18601));
  NAND3X1 g15172(.A(n14962), .B(P1_STATE2_REG_2__SCAN_IN), .C(P1_EAX_REG_31__SCAN_IN), .Y(n18602));
  OAI21X1 g15173(.A0(n17725), .A1(n18598), .B0(n18602), .Y(n18603));
  AOI21X1 g15174(.A0(n18601), .A1(n17662), .B0(n18603), .Y(n18604));
  XOR2X1  g15175(.A(n18604), .B(n17662), .Y(n18605));
  AOI21X1 g15176(.A0(n18589), .A1(n18087), .B0(n18605), .Y(n18606));
  INVX1   g15177(.A(n18606), .Y(n18607));
  NOR4X1  g15178(.A(n17667), .B(n17257), .C(n16815), .D(n18550), .Y(n18608));
  INVX1   g15179(.A(n18605), .Y(n18609));
  NOR4X1  g15180(.A(n17667), .B(n17257), .C(n16815), .D(n18589), .Y(n18610));
  NOR3X1  g15181(.A(n18610), .B(n18609), .C(n18608), .Y(n18611));
  NAND2X1 g15182(.A(n18606), .B(n18608), .Y(n18612));
  NOR2X1  g15183(.A(n18605), .B(n18589), .Y(n18613));
  NAND4X1 g15184(.A(n17747), .B(n17229), .C(n15382), .D(n18613), .Y(n18614));
  NAND3X1 g15185(.A(n18605), .B(n18589), .C(n18087), .Y(n18615));
  NAND3X1 g15186(.A(n18615), .B(n18614), .C(n18612), .Y(n18616));
  AOI21X1 g15187(.A0(n18611), .A1(n18562), .B0(n18616), .Y(n18617));
  OAI21X1 g15188(.A0(n18607), .A1(n18562), .B0(n18617), .Y(n18618));
  INVX1   g15189(.A(P1_REIP_REG_31__SCAN_IN), .Y(n18619));
  AOI22X1 g15190(.A0(n17694), .A1(n18601), .B0(n17686), .B1(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .Y(n18620));
  OAI21X1 g15191(.A0(n16586), .A1(n18619), .B0(n18620), .Y(n18621));
  AOI21X1 g15192(.A0(n17682), .A1(n17644), .B0(n18621), .Y(n18622));
  OAI21X1 g15193(.A0(n18618), .A1(n17688), .B0(n18622), .Y(P1_U2968));
  NAND2X1 g15194(.A(n3070), .B(DATAI_15_), .Y(n18624));
  OAI21X1 g15195(.A0(n3070), .A1(n12788), .B0(n18624), .Y(n18625));
  OAI21X1 g15196(.A0(n14770), .A1(n14707), .B0(n14549), .Y(n18626));
  NAND4X1 g15197(.A(n15316), .B(n15007), .C(n14806), .D(n18626), .Y(n18627));
  NOR2X1  g15198(.A(n18627), .B(n14769), .Y(n18628));
  NOR2X1  g15199(.A(n18627), .B(n14770), .Y(n18629));
  AOI22X1 g15200(.A0(n18628), .A1(n18625), .B0(P1_EAX_REG_15__SCAN_IN), .B1(n18629), .Y(n18630));
  OAI21X1 g15201(.A0(n18627), .A1(n14987), .B0(P1_LWORD_REG_15__SCAN_IN), .Y(n18631));
  OAI21X1 g15202(.A0(n18630), .A1(n14987), .B0(n18631), .Y(P1_U2967));
  NAND2X1 g15203(.A(n3070), .B(DATAI_14_), .Y(n18633));
  OAI21X1 g15204(.A0(n3070), .A1(n12802), .B0(n18633), .Y(n18634));
  AOI22X1 g15205(.A0(n18629), .A1(P1_EAX_REG_14__SCAN_IN), .B0(n18628), .B1(n18634), .Y(n18635));
  OAI21X1 g15206(.A0(n18627), .A1(n14987), .B0(P1_LWORD_REG_14__SCAN_IN), .Y(n18636));
  OAI21X1 g15207(.A0(n18635), .A1(n14987), .B0(n18636), .Y(P1_U2966));
  NAND2X1 g15208(.A(n3070), .B(DATAI_13_), .Y(n18638));
  OAI21X1 g15209(.A0(n3070), .A1(n12809), .B0(n18638), .Y(n18639));
  AOI22X1 g15210(.A0(n18629), .A1(P1_EAX_REG_13__SCAN_IN), .B0(n18628), .B1(n18639), .Y(n18640));
  OAI21X1 g15211(.A0(n18627), .A1(n14987), .B0(P1_LWORD_REG_13__SCAN_IN), .Y(n18641));
  OAI21X1 g15212(.A0(n18640), .A1(n14987), .B0(n18641), .Y(P1_U2965));
  NAND2X1 g15213(.A(n3070), .B(DATAI_12_), .Y(n18643));
  OAI21X1 g15214(.A0(n3070), .A1(n12816), .B0(n18643), .Y(n18644));
  AOI22X1 g15215(.A0(n18629), .A1(P1_EAX_REG_12__SCAN_IN), .B0(n18628), .B1(n18644), .Y(n18645));
  OAI21X1 g15216(.A0(n18627), .A1(n14987), .B0(P1_LWORD_REG_12__SCAN_IN), .Y(n18646));
  OAI21X1 g15217(.A0(n18645), .A1(n14987), .B0(n18646), .Y(P1_U2964));
  NAND2X1 g15218(.A(n3070), .B(DATAI_11_), .Y(n18648));
  OAI21X1 g15219(.A0(n3070), .A1(n12822), .B0(n18648), .Y(n18649));
  AOI22X1 g15220(.A0(n18629), .A1(P1_EAX_REG_11__SCAN_IN), .B0(n18628), .B1(n18649), .Y(n18650));
  OAI21X1 g15221(.A0(n18627), .A1(n14987), .B0(P1_LWORD_REG_11__SCAN_IN), .Y(n18651));
  OAI21X1 g15222(.A0(n18650), .A1(n14987), .B0(n18651), .Y(P1_U2963));
  NAND2X1 g15223(.A(n3070), .B(DATAI_10_), .Y(n18653));
  OAI21X1 g15224(.A0(n3070), .A1(n12828), .B0(n18653), .Y(n18654));
  AOI22X1 g15225(.A0(n18629), .A1(P1_EAX_REG_10__SCAN_IN), .B0(n18628), .B1(n18654), .Y(n18655));
  OAI21X1 g15226(.A0(n18627), .A1(n14987), .B0(P1_LWORD_REG_10__SCAN_IN), .Y(n18656));
  OAI21X1 g15227(.A0(n18655), .A1(n14987), .B0(n18656), .Y(P1_U2962));
  NAND2X1 g15228(.A(n3070), .B(DATAI_9_), .Y(n18658));
  OAI21X1 g15229(.A0(n3070), .A1(n12834), .B0(n18658), .Y(n18659));
  AOI22X1 g15230(.A0(n18629), .A1(P1_EAX_REG_9__SCAN_IN), .B0(n18628), .B1(n18659), .Y(n18660));
  OAI21X1 g15231(.A0(n18627), .A1(n14987), .B0(P1_LWORD_REG_9__SCAN_IN), .Y(n18661));
  OAI21X1 g15232(.A0(n18660), .A1(n14987), .B0(n18661), .Y(P1_U2961));
  NAND2X1 g15233(.A(n3070), .B(DATAI_8_), .Y(n18663));
  OAI21X1 g15234(.A0(n3070), .A1(n12840), .B0(n18663), .Y(n18664));
  AOI22X1 g15235(.A0(n18629), .A1(P1_EAX_REG_8__SCAN_IN), .B0(n18628), .B1(n18664), .Y(n18665));
  OAI21X1 g15236(.A0(n18627), .A1(n14987), .B0(P1_LWORD_REG_8__SCAN_IN), .Y(n18666));
  OAI21X1 g15237(.A0(n18665), .A1(n14987), .B0(n18666), .Y(P1_U2960));
  INVX1   g15238(.A(n15499), .Y(n18668));
  AOI22X1 g15239(.A0(n18628), .A1(n18668), .B0(P1_EAX_REG_7__SCAN_IN), .B1(n18629), .Y(n18669));
  OAI21X1 g15240(.A0(n18627), .A1(n14987), .B0(P1_LWORD_REG_7__SCAN_IN), .Y(n18670));
  OAI21X1 g15241(.A0(n18669), .A1(n14987), .B0(n18670), .Y(P1_U2959));
  INVX1   g15242(.A(n15519), .Y(n18672));
  AOI22X1 g15243(.A0(n18628), .A1(n18672), .B0(P1_EAX_REG_6__SCAN_IN), .B1(n18629), .Y(n18673));
  OAI21X1 g15244(.A0(n18627), .A1(n14987), .B0(P1_LWORD_REG_6__SCAN_IN), .Y(n18674));
  OAI21X1 g15245(.A0(n18673), .A1(n14987), .B0(n18674), .Y(P1_U2958));
  INVX1   g15246(.A(n15534), .Y(n18676));
  AOI22X1 g15247(.A0(n18628), .A1(n18676), .B0(P1_EAX_REG_5__SCAN_IN), .B1(n18629), .Y(n18677));
  OAI21X1 g15248(.A0(n18627), .A1(n14987), .B0(P1_LWORD_REG_5__SCAN_IN), .Y(n18678));
  OAI21X1 g15249(.A0(n18677), .A1(n14987), .B0(n18678), .Y(P1_U2957));
  INVX1   g15250(.A(n15549), .Y(n18680));
  AOI22X1 g15251(.A0(n18628), .A1(n18680), .B0(P1_EAX_REG_4__SCAN_IN), .B1(n18629), .Y(n18681));
  OAI21X1 g15252(.A0(n18627), .A1(n14987), .B0(P1_LWORD_REG_4__SCAN_IN), .Y(n18682));
  OAI21X1 g15253(.A0(n18681), .A1(n14987), .B0(n18682), .Y(P1_U2956));
  INVX1   g15254(.A(n15564), .Y(n18684));
  AOI22X1 g15255(.A0(n18628), .A1(n18684), .B0(P1_EAX_REG_3__SCAN_IN), .B1(n18629), .Y(n18685));
  OAI21X1 g15256(.A0(n18627), .A1(n14987), .B0(P1_LWORD_REG_3__SCAN_IN), .Y(n18686));
  OAI21X1 g15257(.A0(n18685), .A1(n14987), .B0(n18686), .Y(P1_U2955));
  INVX1   g15258(.A(n15580), .Y(n18688));
  AOI22X1 g15259(.A0(n18628), .A1(n18688), .B0(P1_EAX_REG_2__SCAN_IN), .B1(n18629), .Y(n18689));
  OAI21X1 g15260(.A0(n18627), .A1(n14987), .B0(P1_LWORD_REG_2__SCAN_IN), .Y(n18690));
  OAI21X1 g15261(.A0(n18689), .A1(n14987), .B0(n18690), .Y(P1_U2954));
  INVX1   g15262(.A(n15596), .Y(n18692));
  AOI22X1 g15263(.A0(n18628), .A1(n18692), .B0(P1_EAX_REG_1__SCAN_IN), .B1(n18629), .Y(n18693));
  OAI21X1 g15264(.A0(n18627), .A1(n14987), .B0(P1_LWORD_REG_1__SCAN_IN), .Y(n18694));
  OAI21X1 g15265(.A0(n18693), .A1(n14987), .B0(n18694), .Y(P1_U2953));
  INVX1   g15266(.A(n15612), .Y(n18696));
  AOI22X1 g15267(.A0(n18628), .A1(n18696), .B0(P1_EAX_REG_0__SCAN_IN), .B1(n18629), .Y(n18697));
  OAI21X1 g15268(.A0(n18627), .A1(n14987), .B0(P1_LWORD_REG_0__SCAN_IN), .Y(n18698));
  OAI21X1 g15269(.A0(n18697), .A1(n14987), .B0(n18698), .Y(P1_U2952));
  AOI22X1 g15270(.A0(n18629), .A1(P1_EAX_REG_30__SCAN_IN), .B0(n18628), .B1(n18634), .Y(n18700));
  OAI21X1 g15271(.A0(n18627), .A1(n14987), .B0(P1_UWORD_REG_14__SCAN_IN), .Y(n18701));
  OAI21X1 g15272(.A0(n18700), .A1(n14987), .B0(n18701), .Y(P1_U2951));
  AOI22X1 g15273(.A0(n18629), .A1(P1_EAX_REG_29__SCAN_IN), .B0(n18628), .B1(n18639), .Y(n18703));
  OAI21X1 g15274(.A0(n18627), .A1(n14987), .B0(P1_UWORD_REG_13__SCAN_IN), .Y(n18704));
  OAI21X1 g15275(.A0(n18703), .A1(n14987), .B0(n18704), .Y(P1_U2950));
  AOI22X1 g15276(.A0(n18629), .A1(P1_EAX_REG_28__SCAN_IN), .B0(n18628), .B1(n18644), .Y(n18706));
  OAI21X1 g15277(.A0(n18627), .A1(n14987), .B0(P1_UWORD_REG_12__SCAN_IN), .Y(n18707));
  OAI21X1 g15278(.A0(n18706), .A1(n14987), .B0(n18707), .Y(P1_U2949));
  AOI22X1 g15279(.A0(n18629), .A1(P1_EAX_REG_27__SCAN_IN), .B0(n18628), .B1(n18649), .Y(n18709));
  OAI21X1 g15280(.A0(n18627), .A1(n14987), .B0(P1_UWORD_REG_11__SCAN_IN), .Y(n18710));
  OAI21X1 g15281(.A0(n18709), .A1(n14987), .B0(n18710), .Y(P1_U2948));
  AOI22X1 g15282(.A0(n18629), .A1(P1_EAX_REG_26__SCAN_IN), .B0(n18628), .B1(n18654), .Y(n18712));
  OAI21X1 g15283(.A0(n18627), .A1(n14987), .B0(P1_UWORD_REG_10__SCAN_IN), .Y(n18713));
  OAI21X1 g15284(.A0(n18712), .A1(n14987), .B0(n18713), .Y(P1_U2947));
  AOI22X1 g15285(.A0(n18629), .A1(P1_EAX_REG_25__SCAN_IN), .B0(n18628), .B1(n18659), .Y(n18715));
  OAI21X1 g15286(.A0(n18627), .A1(n14987), .B0(P1_UWORD_REG_9__SCAN_IN), .Y(n18716));
  OAI21X1 g15287(.A0(n18715), .A1(n14987), .B0(n18716), .Y(P1_U2946));
  AOI22X1 g15288(.A0(n18629), .A1(P1_EAX_REG_24__SCAN_IN), .B0(n18628), .B1(n18664), .Y(n18718));
  OAI21X1 g15289(.A0(n18627), .A1(n14987), .B0(P1_UWORD_REG_8__SCAN_IN), .Y(n18719));
  OAI21X1 g15290(.A0(n18718), .A1(n14987), .B0(n18719), .Y(P1_U2945));
  AOI22X1 g15291(.A0(n18628), .A1(n18668), .B0(P1_EAX_REG_23__SCAN_IN), .B1(n18629), .Y(n18721));
  OAI21X1 g15292(.A0(n18627), .A1(n14987), .B0(P1_UWORD_REG_7__SCAN_IN), .Y(n18722));
  OAI21X1 g15293(.A0(n18721), .A1(n14987), .B0(n18722), .Y(P1_U2944));
  AOI22X1 g15294(.A0(n18628), .A1(n18672), .B0(P1_EAX_REG_22__SCAN_IN), .B1(n18629), .Y(n18724));
  OAI21X1 g15295(.A0(n18627), .A1(n14987), .B0(P1_UWORD_REG_6__SCAN_IN), .Y(n18725));
  OAI21X1 g15296(.A0(n18724), .A1(n14987), .B0(n18725), .Y(P1_U2943));
  AOI22X1 g15297(.A0(n18628), .A1(n18676), .B0(P1_EAX_REG_21__SCAN_IN), .B1(n18629), .Y(n18727));
  OAI21X1 g15298(.A0(n18627), .A1(n14987), .B0(P1_UWORD_REG_5__SCAN_IN), .Y(n18728));
  OAI21X1 g15299(.A0(n18727), .A1(n14987), .B0(n18728), .Y(P1_U2942));
  AOI22X1 g15300(.A0(n18628), .A1(n18680), .B0(P1_EAX_REG_20__SCAN_IN), .B1(n18629), .Y(n18730));
  OAI21X1 g15301(.A0(n18627), .A1(n14987), .B0(P1_UWORD_REG_4__SCAN_IN), .Y(n18731));
  OAI21X1 g15302(.A0(n18730), .A1(n14987), .B0(n18731), .Y(P1_U2941));
  AOI22X1 g15303(.A0(n18628), .A1(n18684), .B0(P1_EAX_REG_19__SCAN_IN), .B1(n18629), .Y(n18733));
  OAI21X1 g15304(.A0(n18627), .A1(n14987), .B0(P1_UWORD_REG_3__SCAN_IN), .Y(n18734));
  OAI21X1 g15305(.A0(n18733), .A1(n14987), .B0(n18734), .Y(P1_U2940));
  AOI22X1 g15306(.A0(n18628), .A1(n18688), .B0(P1_EAX_REG_18__SCAN_IN), .B1(n18629), .Y(n18736));
  OAI21X1 g15307(.A0(n18627), .A1(n14987), .B0(P1_UWORD_REG_2__SCAN_IN), .Y(n18737));
  OAI21X1 g15308(.A0(n18736), .A1(n14987), .B0(n18737), .Y(P1_U2939));
  AOI22X1 g15309(.A0(n18628), .A1(n18692), .B0(P1_EAX_REG_17__SCAN_IN), .B1(n18629), .Y(n18739));
  OAI21X1 g15310(.A0(n18627), .A1(n14987), .B0(P1_UWORD_REG_1__SCAN_IN), .Y(n18740));
  OAI21X1 g15311(.A0(n18739), .A1(n14987), .B0(n18740), .Y(P1_U2938));
  AOI22X1 g15312(.A0(n18628), .A1(n18696), .B0(P1_EAX_REG_16__SCAN_IN), .B1(n18629), .Y(n18742));
  OAI21X1 g15313(.A0(n18627), .A1(n14987), .B0(P1_UWORD_REG_0__SCAN_IN), .Y(n18743));
  OAI21X1 g15314(.A0(n18742), .A1(n14987), .B0(n18743), .Y(P1_U2937));
  NOR2X1  g15315(.A(n15093), .B(n15155), .Y(n18745));
  NOR3X1  g15316(.A(n15339), .B(n14987), .C(n15021), .Y(n18746));
  OAI21X1 g15317(.A0(n18746), .A1(n15237), .B0(n15156), .Y(n18747));
  INVX1   g15318(.A(n18747), .Y(n18748));
  AOI22X1 g15319(.A0(n15293), .A1(n18748), .B0(n18745), .B1(n14650), .Y(n18749));
  NOR2X1  g15320(.A(n18749), .B(n14650), .Y(n18750));
  INVX1   g15321(.A(n18750), .Y(n18751));
  NOR2X1  g15322(.A(n18749), .B(P1_STATE2_REG_0__SCAN_IN), .Y(n18752));
  AOI22X1 g15323(.A0(n18749), .A1(P1_DATAO_REG_0__SCAN_IN), .B0(P1_LWORD_REG_0__SCAN_IN), .B1(n18752), .Y(n18753));
  OAI21X1 g15324(.A0(n18751), .A1(n17669), .B0(n18753), .Y(P1_U2936));
  AOI22X1 g15325(.A0(n18749), .A1(P1_DATAO_REG_1__SCAN_IN), .B0(P1_LWORD_REG_1__SCAN_IN), .B1(n18752), .Y(n18755));
  OAI21X1 g15326(.A0(n18751), .A1(n17700), .B0(n18755), .Y(P1_U2935));
  AOI22X1 g15327(.A0(n18749), .A1(P1_DATAO_REG_2__SCAN_IN), .B0(P1_LWORD_REG_2__SCAN_IN), .B1(n18752), .Y(n18757));
  OAI21X1 g15328(.A0(n18751), .A1(n17727), .B0(n18757), .Y(P1_U2934));
  NAND2X1 g15329(.A(n18750), .B(P1_EAX_REG_3__SCAN_IN), .Y(n18759));
  AOI22X1 g15330(.A0(n18749), .A1(P1_DATAO_REG_3__SCAN_IN), .B0(P1_LWORD_REG_3__SCAN_IN), .B1(n18752), .Y(n18760));
  NAND2X1 g15331(.A(n18760), .B(n18759), .Y(P1_U2933));
  AOI22X1 g15332(.A0(n18749), .A1(P1_DATAO_REG_4__SCAN_IN), .B0(P1_LWORD_REG_4__SCAN_IN), .B1(n18752), .Y(n18762));
  OAI21X1 g15333(.A0(n18751), .A1(n17769), .B0(n18762), .Y(P1_U2932));
  NAND2X1 g15334(.A(n18750), .B(P1_EAX_REG_5__SCAN_IN), .Y(n18764));
  AOI22X1 g15335(.A0(n18749), .A1(P1_DATAO_REG_5__SCAN_IN), .B0(P1_LWORD_REG_5__SCAN_IN), .B1(n18752), .Y(n18765));
  NAND2X1 g15336(.A(n18765), .B(n18764), .Y(P1_U2931));
  NAND2X1 g15337(.A(n18750), .B(P1_EAX_REG_6__SCAN_IN), .Y(n18767));
  AOI22X1 g15338(.A0(n18749), .A1(P1_DATAO_REG_6__SCAN_IN), .B0(P1_LWORD_REG_6__SCAN_IN), .B1(n18752), .Y(n18768));
  NAND2X1 g15339(.A(n18768), .B(n18767), .Y(P1_U2930));
  NAND2X1 g15340(.A(n18750), .B(P1_EAX_REG_7__SCAN_IN), .Y(n18770));
  AOI22X1 g15341(.A0(n18749), .A1(P1_DATAO_REG_7__SCAN_IN), .B0(P1_LWORD_REG_7__SCAN_IN), .B1(n18752), .Y(n18771));
  NAND2X1 g15342(.A(n18771), .B(n18770), .Y(P1_U2929));
  NAND2X1 g15343(.A(n18750), .B(P1_EAX_REG_8__SCAN_IN), .Y(n18773));
  AOI22X1 g15344(.A0(n18749), .A1(P1_DATAO_REG_8__SCAN_IN), .B0(P1_LWORD_REG_8__SCAN_IN), .B1(n18752), .Y(n18774));
  NAND2X1 g15345(.A(n18774), .B(n18773), .Y(P1_U2928));
  AOI22X1 g15346(.A0(n18749), .A1(P1_DATAO_REG_9__SCAN_IN), .B0(P1_LWORD_REG_9__SCAN_IN), .B1(n18752), .Y(n18776));
  OAI21X1 g15347(.A0(n18751), .A1(n17886), .B0(n18776), .Y(P1_U2927));
  AOI22X1 g15348(.A0(n18749), .A1(P1_DATAO_REG_10__SCAN_IN), .B0(P1_LWORD_REG_10__SCAN_IN), .B1(n18752), .Y(n18778));
  OAI21X1 g15349(.A0(n18751), .A1(n17908), .B0(n18778), .Y(P1_U2926));
  AOI22X1 g15350(.A0(n18749), .A1(P1_DATAO_REG_11__SCAN_IN), .B0(P1_LWORD_REG_11__SCAN_IN), .B1(n18752), .Y(n18780));
  OAI21X1 g15351(.A0(n18751), .A1(n17927), .B0(n18780), .Y(P1_U2925));
  AOI22X1 g15352(.A0(n18749), .A1(P1_DATAO_REG_12__SCAN_IN), .B0(P1_LWORD_REG_12__SCAN_IN), .B1(n18752), .Y(n18782));
  OAI21X1 g15353(.A0(n18751), .A1(n17944), .B0(n18782), .Y(P1_U2924));
  AOI22X1 g15354(.A0(n18749), .A1(P1_DATAO_REG_13__SCAN_IN), .B0(P1_LWORD_REG_13__SCAN_IN), .B1(n18752), .Y(n18784));
  OAI21X1 g15355(.A0(n18751), .A1(n17970), .B0(n18784), .Y(P1_U2923));
  AOI22X1 g15356(.A0(n18749), .A1(P1_DATAO_REG_14__SCAN_IN), .B0(P1_LWORD_REG_14__SCAN_IN), .B1(n18752), .Y(n18786));
  OAI21X1 g15357(.A0(n18751), .A1(n17992), .B0(n18786), .Y(P1_U2922));
  AOI22X1 g15358(.A0(n18749), .A1(P1_DATAO_REG_15__SCAN_IN), .B0(P1_LWORD_REG_15__SCAN_IN), .B1(n18752), .Y(n18788));
  OAI21X1 g15359(.A0(n18751), .A1(n18012), .B0(n18788), .Y(P1_U2921));
  INVX1   g15360(.A(P1_EAX_REG_16__SCAN_IN), .Y(n18790));
  NAND2X1 g15361(.A(n18750), .B(n14806), .Y(n18791));
  AOI22X1 g15362(.A0(n18749), .A1(P1_DATAO_REG_16__SCAN_IN), .B0(P1_UWORD_REG_0__SCAN_IN), .B1(n18752), .Y(n18792));
  OAI21X1 g15363(.A0(n18791), .A1(n18790), .B0(n18792), .Y(P1_U2920));
  INVX1   g15364(.A(P1_EAX_REG_17__SCAN_IN), .Y(n18794));
  AOI22X1 g15365(.A0(n18749), .A1(P1_DATAO_REG_17__SCAN_IN), .B0(P1_UWORD_REG_1__SCAN_IN), .B1(n18752), .Y(n18795));
  OAI21X1 g15366(.A0(n18791), .A1(n18794), .B0(n18795), .Y(P1_U2919));
  INVX1   g15367(.A(P1_EAX_REG_18__SCAN_IN), .Y(n18797));
  AOI22X1 g15368(.A0(n18749), .A1(P1_DATAO_REG_18__SCAN_IN), .B0(P1_UWORD_REG_2__SCAN_IN), .B1(n18752), .Y(n18798));
  OAI21X1 g15369(.A0(n18791), .A1(n18797), .B0(n18798), .Y(P1_U2918));
  INVX1   g15370(.A(P1_EAX_REG_19__SCAN_IN), .Y(n18800));
  AOI22X1 g15371(.A0(n18749), .A1(P1_DATAO_REG_19__SCAN_IN), .B0(P1_UWORD_REG_3__SCAN_IN), .B1(n18752), .Y(n18801));
  OAI21X1 g15372(.A0(n18791), .A1(n18800), .B0(n18801), .Y(P1_U2917));
  INVX1   g15373(.A(P1_EAX_REG_20__SCAN_IN), .Y(n18803));
  AOI22X1 g15374(.A0(n18749), .A1(P1_DATAO_REG_20__SCAN_IN), .B0(P1_UWORD_REG_4__SCAN_IN), .B1(n18752), .Y(n18804));
  OAI21X1 g15375(.A0(n18791), .A1(n18803), .B0(n18804), .Y(P1_U2916));
  AOI22X1 g15376(.A0(n18749), .A1(P1_DATAO_REG_21__SCAN_IN), .B0(P1_UWORD_REG_5__SCAN_IN), .B1(n18752), .Y(n18806));
  OAI21X1 g15377(.A0(n18791), .A1(n18234), .B0(n18806), .Y(P1_U2915));
  AOI22X1 g15378(.A0(n18749), .A1(P1_DATAO_REG_22__SCAN_IN), .B0(P1_UWORD_REG_6__SCAN_IN), .B1(n18752), .Y(n18808));
  OAI21X1 g15379(.A0(n18791), .A1(n18271), .B0(n18808), .Y(P1_U2914));
  AOI22X1 g15380(.A0(n18749), .A1(P1_DATAO_REG_23__SCAN_IN), .B0(P1_UWORD_REG_7__SCAN_IN), .B1(n18752), .Y(n18810));
  OAI21X1 g15381(.A0(n18791), .A1(n18336), .B0(n18810), .Y(P1_U2913));
  AOI22X1 g15382(.A0(n18749), .A1(P1_DATAO_REG_24__SCAN_IN), .B0(P1_UWORD_REG_8__SCAN_IN), .B1(n18752), .Y(n18812));
  OAI21X1 g15383(.A0(n18791), .A1(n18371), .B0(n18812), .Y(P1_U2912));
  INVX1   g15384(.A(P1_EAX_REG_25__SCAN_IN), .Y(n18814));
  AOI22X1 g15385(.A0(n18749), .A1(P1_DATAO_REG_25__SCAN_IN), .B0(P1_UWORD_REG_9__SCAN_IN), .B1(n18752), .Y(n18815));
  OAI21X1 g15386(.A0(n18791), .A1(n18814), .B0(n18815), .Y(P1_U2911));
  INVX1   g15387(.A(P1_EAX_REG_26__SCAN_IN), .Y(n18817));
  AOI22X1 g15388(.A0(n18749), .A1(P1_DATAO_REG_26__SCAN_IN), .B0(P1_UWORD_REG_10__SCAN_IN), .B1(n18752), .Y(n18818));
  OAI21X1 g15389(.A0(n18791), .A1(n18817), .B0(n18818), .Y(P1_U2910));
  INVX1   g15390(.A(P1_EAX_REG_27__SCAN_IN), .Y(n18820));
  AOI22X1 g15391(.A0(n18749), .A1(P1_DATAO_REG_27__SCAN_IN), .B0(P1_UWORD_REG_11__SCAN_IN), .B1(n18752), .Y(n18821));
  OAI21X1 g15392(.A0(n18791), .A1(n18820), .B0(n18821), .Y(P1_U2909));
  INVX1   g15393(.A(P1_EAX_REG_28__SCAN_IN), .Y(n18823));
  AOI22X1 g15394(.A0(n18749), .A1(P1_DATAO_REG_28__SCAN_IN), .B0(P1_UWORD_REG_12__SCAN_IN), .B1(n18752), .Y(n18824));
  OAI21X1 g15395(.A0(n18791), .A1(n18823), .B0(n18824), .Y(P1_U2908));
  INVX1   g15396(.A(P1_EAX_REG_29__SCAN_IN), .Y(n18826));
  AOI22X1 g15397(.A0(n18749), .A1(P1_DATAO_REG_29__SCAN_IN), .B0(P1_UWORD_REG_13__SCAN_IN), .B1(n18752), .Y(n18827));
  OAI21X1 g15398(.A0(n18791), .A1(n18826), .B0(n18827), .Y(P1_U2907));
  AOI22X1 g15399(.A0(n18749), .A1(P1_DATAO_REG_30__SCAN_IN), .B0(P1_UWORD_REG_14__SCAN_IN), .B1(n18752), .Y(n18829));
  OAI21X1 g15400(.A0(n18791), .A1(n18585), .B0(n18829), .Y(P1_U2906));
  INVX1   g15401(.A(n18749), .Y(n18831));
  NOR2X1  g15402(.A(n18831), .B(n2966), .Y(P1_U2905));
  NOR4X1  g15403(.A(n15268), .B(n14807), .C(n14650), .D(n14987), .Y(n18833));
  NOR3X1  g15404(.A(n15286), .B(n15137), .C(n15150), .Y(n18834));
  OAI21X1 g15405(.A0(n18834), .A1(n18833), .B0(n14550), .Y(n18835));
  NOR4X1  g15406(.A(n14985), .B(n14940), .C(n15150), .D(n15000), .Y(n18836));
  NOR4X1  g15407(.A(n15065), .B(n15046), .C(n15150), .D(n15070), .Y(n18837));
  AOI21X1 g15408(.A0(n18836), .A1(n15007), .B0(n18837), .Y(n18838));
  AOI21X1 g15409(.A0(n18838), .A1(n18835), .B0(n15157), .Y(n18839));
  OAI21X1 g15410(.A0(n15022), .A1(n14962), .B0(n18839), .Y(n18840));
  INVX1   g15411(.A(n18839), .Y(n18841));
  NOR3X1  g15412(.A(n18841), .B(n15022), .C(n14962), .Y(n18842));
  AOI22X1 g15413(.A0(n18841), .A1(P1_EAX_REG_0__SCAN_IN), .B0(n18696), .B1(n18842), .Y(n18843));
  OAI21X1 g15414(.A0(n18840), .A1(n17679), .B0(n18843), .Y(P1_U2904));
  AOI22X1 g15415(.A0(n18841), .A1(P1_EAX_REG_1__SCAN_IN), .B0(n18692), .B1(n18842), .Y(n18845));
  OAI21X1 g15416(.A0(n18840), .A1(n17715), .B0(n18845), .Y(P1_U2903));
  AOI22X1 g15417(.A0(n18841), .A1(P1_EAX_REG_2__SCAN_IN), .B0(n18688), .B1(n18842), .Y(n18847));
  OAI21X1 g15418(.A0(n18840), .A1(n17741), .B0(n18847), .Y(P1_U2902));
  INVX1   g15419(.A(n17762), .Y(n18849));
  AOI22X1 g15420(.A0(n18841), .A1(P1_EAX_REG_3__SCAN_IN), .B0(n18684), .B1(n18842), .Y(n18850));
  OAI21X1 g15421(.A0(n18840), .A1(n18849), .B0(n18850), .Y(P1_U2901));
  AOI22X1 g15422(.A0(n18841), .A1(P1_EAX_REG_4__SCAN_IN), .B0(n18680), .B1(n18842), .Y(n18852));
  OAI21X1 g15423(.A0(n18840), .A1(n17786), .B0(n18852), .Y(P1_U2900));
  AOI22X1 g15424(.A0(n18841), .A1(P1_EAX_REG_5__SCAN_IN), .B0(n18676), .B1(n18842), .Y(n18854));
  OAI21X1 g15425(.A0(n18840), .A1(n17809), .B0(n18854), .Y(P1_U2899));
  AOI22X1 g15426(.A0(n18841), .A1(P1_EAX_REG_6__SCAN_IN), .B0(n18672), .B1(n18842), .Y(n18856));
  OAI21X1 g15427(.A0(n18840), .A1(n17831), .B0(n18856), .Y(P1_U2898));
  AOI22X1 g15428(.A0(n18841), .A1(P1_EAX_REG_7__SCAN_IN), .B0(n18668), .B1(n18842), .Y(n18858));
  OAI21X1 g15429(.A0(n18840), .A1(n17849), .B0(n18858), .Y(P1_U2897));
  AOI22X1 g15430(.A0(n18841), .A1(P1_EAX_REG_8__SCAN_IN), .B0(n18664), .B1(n18842), .Y(n18860));
  OAI21X1 g15431(.A0(n18840), .A1(n17876), .B0(n18860), .Y(P1_U2896));
  AOI22X1 g15432(.A0(n18841), .A1(P1_EAX_REG_9__SCAN_IN), .B0(n18659), .B1(n18842), .Y(n18862));
  OAI21X1 g15433(.A0(n18840), .A1(n17896), .B0(n18862), .Y(P1_U2895));
  AOI22X1 g15434(.A0(n18841), .A1(P1_EAX_REG_10__SCAN_IN), .B0(n18654), .B1(n18842), .Y(n18864));
  OAI21X1 g15435(.A0(n18840), .A1(n17918), .B0(n18864), .Y(P1_U2894));
  INVX1   g15436(.A(n17937), .Y(n18866));
  AOI22X1 g15437(.A0(n18841), .A1(P1_EAX_REG_11__SCAN_IN), .B0(n18649), .B1(n18842), .Y(n18867));
  OAI21X1 g15438(.A0(n18840), .A1(n18866), .B0(n18867), .Y(P1_U2893));
  AOI22X1 g15439(.A0(n18841), .A1(P1_EAX_REG_12__SCAN_IN), .B0(n18644), .B1(n18842), .Y(n18869));
  OAI21X1 g15440(.A0(n18840), .A1(n17962), .B0(n18869), .Y(P1_U2892));
  AOI22X1 g15441(.A0(n18841), .A1(P1_EAX_REG_13__SCAN_IN), .B0(n18639), .B1(n18842), .Y(n18871));
  OAI21X1 g15442(.A0(n18840), .A1(n17980), .B0(n18871), .Y(P1_U2891));
  AOI22X1 g15443(.A0(n18841), .A1(P1_EAX_REG_14__SCAN_IN), .B0(n18634), .B1(n18842), .Y(n18873));
  OAI21X1 g15444(.A0(n18840), .A1(n18003), .B0(n18873), .Y(P1_U2890));
  INVX1   g15445(.A(n18025), .Y(n18875));
  AOI22X1 g15446(.A0(n18841), .A1(P1_EAX_REG_15__SCAN_IN), .B0(n18625), .B1(n18842), .Y(n18876));
  OAI21X1 g15447(.A0(n18840), .A1(n18875), .B0(n18876), .Y(P1_U2889));
  NOR3X1  g15448(.A(n18841), .B(n14962), .C(n14801), .Y(n18878));
  NOR2X1  g15449(.A(n18841), .B(n14993), .Y(n18879));
  INVX1   g15450(.A(n18879), .Y(n18880));
  OAI22X1 g15451(.A0(n18839), .A1(n18790), .B0(n15619), .B1(n18880), .Y(n18881));
  AOI21X1 g15452(.A0(n18878), .A1(n18696), .B0(n18881), .Y(n18882));
  OAI21X1 g15453(.A0(n18840), .A1(n18080), .B0(n18882), .Y(P1_U2888));
  OAI22X1 g15454(.A0(n18839), .A1(n18794), .B0(n15603), .B1(n18880), .Y(n18884));
  AOI21X1 g15455(.A0(n18878), .A1(n18692), .B0(n18884), .Y(n18885));
  OAI21X1 g15456(.A0(n18840), .A1(n18108), .B0(n18885), .Y(P1_U2887));
  INVX1   g15457(.A(n18141), .Y(n18887));
  OAI22X1 g15458(.A0(n18839), .A1(n18797), .B0(n15587), .B1(n18880), .Y(n18888));
  AOI21X1 g15459(.A0(n18878), .A1(n18688), .B0(n18888), .Y(n18889));
  OAI21X1 g15460(.A0(n18840), .A1(n18887), .B0(n18889), .Y(P1_U2886));
  OAI22X1 g15461(.A0(n18839), .A1(n18800), .B0(n15571), .B1(n18880), .Y(n18891));
  AOI21X1 g15462(.A0(n18878), .A1(n18684), .B0(n18891), .Y(n18892));
  OAI21X1 g15463(.A0(n18840), .A1(n18173), .B0(n18892), .Y(P1_U2885));
  OAI22X1 g15464(.A0(n18839), .A1(n18803), .B0(n15557), .B1(n18880), .Y(n18894));
  AOI21X1 g15465(.A0(n18878), .A1(n18680), .B0(n18894), .Y(n18895));
  OAI21X1 g15466(.A0(n18840), .A1(n18202), .B0(n18895), .Y(P1_U2884));
  OAI22X1 g15467(.A0(n18839), .A1(n18234), .B0(n15542), .B1(n18880), .Y(n18897));
  AOI21X1 g15468(.A0(n18878), .A1(n18676), .B0(n18897), .Y(n18898));
  OAI21X1 g15469(.A0(n18840), .A1(n18245), .B0(n18898), .Y(P1_U2883));
  OAI22X1 g15470(.A0(n18839), .A1(n18271), .B0(n15527), .B1(n18880), .Y(n18900));
  AOI21X1 g15471(.A0(n18878), .A1(n18672), .B0(n18900), .Y(n18901));
  OAI21X1 g15472(.A0(n18840), .A1(n18283), .B0(n18901), .Y(P1_U2882));
  OAI22X1 g15473(.A0(n18839), .A1(n18336), .B0(n15510), .B1(n18880), .Y(n18903));
  AOI21X1 g15474(.A0(n18878), .A1(n18668), .B0(n18903), .Y(n18904));
  OAI21X1 g15475(.A0(n18840), .A1(n18348), .B0(n18904), .Y(P1_U2881));
  OAI22X1 g15476(.A0(n18839), .A1(n18371), .B0(n15616), .B1(n18880), .Y(n18906));
  AOI21X1 g15477(.A0(n18878), .A1(n18664), .B0(n18906), .Y(n18907));
  OAI21X1 g15478(.A0(n18840), .A1(n18380), .B0(n18907), .Y(P1_U2880));
  OAI22X1 g15479(.A0(n18839), .A1(n18814), .B0(n15600), .B1(n18880), .Y(n18909));
  AOI21X1 g15480(.A0(n18878), .A1(n18659), .B0(n18909), .Y(n18910));
  OAI21X1 g15481(.A0(n18840), .A1(n18412), .B0(n18910), .Y(P1_U2879));
  OAI22X1 g15482(.A0(n18839), .A1(n18817), .B0(n15584), .B1(n18880), .Y(n18912));
  AOI21X1 g15483(.A0(n18878), .A1(n18654), .B0(n18912), .Y(n18913));
  OAI21X1 g15484(.A0(n18840), .A1(n18449), .B0(n18913), .Y(P1_U2878));
  INVX1   g15485(.A(n18485), .Y(n18915));
  OAI22X1 g15486(.A0(n18839), .A1(n18820), .B0(n15568), .B1(n18880), .Y(n18916));
  AOI21X1 g15487(.A0(n18878), .A1(n18649), .B0(n18916), .Y(n18917));
  OAI21X1 g15488(.A0(n18840), .A1(n18915), .B0(n18917), .Y(P1_U2877));
  OAI22X1 g15489(.A0(n18839), .A1(n18823), .B0(n15553), .B1(n18880), .Y(n18919));
  AOI21X1 g15490(.A0(n18878), .A1(n18644), .B0(n18919), .Y(n18920));
  OAI21X1 g15491(.A0(n18840), .A1(n18523), .B0(n18920), .Y(P1_U2876));
  OAI22X1 g15492(.A0(n18839), .A1(n18826), .B0(n15538), .B1(n18880), .Y(n18922));
  AOI21X1 g15493(.A0(n18878), .A1(n18639), .B0(n18922), .Y(n18923));
  OAI21X1 g15494(.A0(n18840), .A1(n18555), .B0(n18923), .Y(P1_U2875));
  OAI22X1 g15495(.A0(n18839), .A1(n18585), .B0(n15523), .B1(n18880), .Y(n18925));
  AOI21X1 g15496(.A0(n18878), .A1(n18634), .B0(n18925), .Y(n18926));
  OAI21X1 g15497(.A0(n18840), .A1(n18591), .B0(n18926), .Y(P1_U2874));
  NAND2X1 g15498(.A(n18839), .B(n14962), .Y(n18928));
  NOR3X1  g15499(.A(n18841), .B(n15506), .C(n14993), .Y(n18929));
  AOI21X1 g15500(.A0(n18841), .A1(P1_EAX_REG_31__SCAN_IN), .B0(n18929), .Y(n18930));
  OAI21X1 g15501(.A0(n18928), .A1(n18618), .B0(n18930), .Y(P1_U2873));
  NAND2X1 g15502(.A(n14984), .B(P1_STATE2_REG_0__SCAN_IN), .Y(n18932));
  NOR4X1  g15503(.A(n15024), .B(n14769), .C(n14707), .D(n18932), .Y(n18933));
  NOR3X1  g15504(.A(n15011), .B(n15007), .C(n14650), .Y(n18934));
  AOI21X1 g15505(.A0(n18933), .A1(n15072), .B0(n18934), .Y(n18935));
  NOR2X1  g15506(.A(n18935), .B(n15157), .Y(n18936));
  NAND2X1 g15507(.A(n18936), .B(n15042), .Y(n18937));
  INVX1   g15508(.A(n18936), .Y(n18938));
  NOR3X1  g15509(.A(n18935), .B(n15157), .C(n15042), .Y(n18939));
  AOI22X1 g15510(.A0(n18938), .A1(P1_EBX_REG_0__SCAN_IN), .B0(n16556), .B1(n18939), .Y(n18940));
  OAI21X1 g15511(.A0(n18937), .A1(n17679), .B0(n18940), .Y(P1_U2872));
  AOI22X1 g15512(.A0(n18938), .A1(P1_EBX_REG_1__SCAN_IN), .B0(n16569), .B1(n18939), .Y(n18942));
  OAI21X1 g15513(.A0(n18937), .A1(n17715), .B0(n18942), .Y(P1_U2871));
  AOI22X1 g15514(.A0(n18938), .A1(P1_EBX_REG_2__SCAN_IN), .B0(n16613), .B1(n18939), .Y(n18944));
  OAI21X1 g15515(.A0(n18937), .A1(n17741), .B0(n18944), .Y(P1_U2870));
  INVX1   g15516(.A(n16634), .Y(n18946));
  AOI22X1 g15517(.A0(n18938), .A1(P1_EBX_REG_3__SCAN_IN), .B0(n18946), .B1(n18939), .Y(n18947));
  OAI21X1 g15518(.A0(n18937), .A1(n18849), .B0(n18947), .Y(P1_U2869));
  INVX1   g15519(.A(n16689), .Y(n18949));
  AOI22X1 g15520(.A0(n18938), .A1(P1_EBX_REG_4__SCAN_IN), .B0(n18949), .B1(n18939), .Y(n18950));
  OAI21X1 g15521(.A0(n18937), .A1(n17786), .B0(n18950), .Y(P1_U2868));
  INVX1   g15522(.A(n16748), .Y(n18952));
  AOI22X1 g15523(.A0(n18938), .A1(P1_EBX_REG_5__SCAN_IN), .B0(n18952), .B1(n18939), .Y(n18953));
  OAI21X1 g15524(.A0(n18937), .A1(n17809), .B0(n18953), .Y(P1_U2867));
  INVX1   g15525(.A(n16802), .Y(n18955));
  AOI22X1 g15526(.A0(n18938), .A1(P1_EBX_REG_6__SCAN_IN), .B0(n18955), .B1(n18939), .Y(n18956));
  OAI21X1 g15527(.A0(n18937), .A1(n17831), .B0(n18956), .Y(P1_U2866));
  INVX1   g15528(.A(n16850), .Y(n18958));
  AOI22X1 g15529(.A0(n18938), .A1(P1_EBX_REG_7__SCAN_IN), .B0(n18958), .B1(n18939), .Y(n18959));
  OAI21X1 g15530(.A0(n18937), .A1(n17849), .B0(n18959), .Y(P1_U2865));
  INVX1   g15531(.A(n16917), .Y(n18961));
  AOI22X1 g15532(.A0(n18938), .A1(P1_EBX_REG_8__SCAN_IN), .B0(n18961), .B1(n18939), .Y(n18962));
  OAI21X1 g15533(.A0(n18937), .A1(n17876), .B0(n18962), .Y(P1_U2864));
  INVX1   g15534(.A(n16956), .Y(n18964));
  AOI22X1 g15535(.A0(n18938), .A1(P1_EBX_REG_9__SCAN_IN), .B0(n18964), .B1(n18939), .Y(n18965));
  OAI21X1 g15536(.A0(n18937), .A1(n17896), .B0(n18965), .Y(P1_U2863));
  INVX1   g15537(.A(n16999), .Y(n18967));
  AOI22X1 g15538(.A0(n18938), .A1(P1_EBX_REG_10__SCAN_IN), .B0(n18967), .B1(n18939), .Y(n18968));
  OAI21X1 g15539(.A0(n18937), .A1(n17918), .B0(n18968), .Y(P1_U2862));
  INVX1   g15540(.A(n17046), .Y(n18970));
  AOI22X1 g15541(.A0(n18938), .A1(P1_EBX_REG_11__SCAN_IN), .B0(n18970), .B1(n18939), .Y(n18971));
  OAI21X1 g15542(.A0(n18937), .A1(n18866), .B0(n18971), .Y(P1_U2861));
  INVX1   g15543(.A(n17090), .Y(n18973));
  AOI22X1 g15544(.A0(n18938), .A1(P1_EBX_REG_12__SCAN_IN), .B0(n18973), .B1(n18939), .Y(n18974));
  OAI21X1 g15545(.A0(n18937), .A1(n17962), .B0(n18974), .Y(P1_U2860));
  INVX1   g15546(.A(n17119), .Y(n18976));
  AOI22X1 g15547(.A0(n18938), .A1(P1_EBX_REG_13__SCAN_IN), .B0(n18976), .B1(n18939), .Y(n18977));
  OAI21X1 g15548(.A0(n18937), .A1(n17980), .B0(n18977), .Y(P1_U2859));
  INVX1   g15549(.A(n17162), .Y(n18979));
  AOI22X1 g15550(.A0(n18938), .A1(P1_EBX_REG_14__SCAN_IN), .B0(n18979), .B1(n18939), .Y(n18980));
  OAI21X1 g15551(.A0(n18937), .A1(n18003), .B0(n18980), .Y(P1_U2858));
  INVX1   g15552(.A(n17204), .Y(n18982));
  AOI22X1 g15553(.A0(n18938), .A1(P1_EBX_REG_15__SCAN_IN), .B0(n18982), .B1(n18939), .Y(n18983));
  OAI21X1 g15554(.A0(n18937), .A1(n18875), .B0(n18983), .Y(P1_U2857));
  INVX1   g15555(.A(n17239), .Y(n18985));
  AOI22X1 g15556(.A0(n18938), .A1(P1_EBX_REG_16__SCAN_IN), .B0(n18985), .B1(n18939), .Y(n18986));
  OAI21X1 g15557(.A0(n18937), .A1(n18080), .B0(n18986), .Y(P1_U2856));
  INVX1   g15558(.A(n17264), .Y(n18988));
  AOI22X1 g15559(.A0(n18938), .A1(P1_EBX_REG_17__SCAN_IN), .B0(n18988), .B1(n18939), .Y(n18989));
  OAI21X1 g15560(.A0(n18937), .A1(n18108), .B0(n18989), .Y(P1_U2855));
  INVX1   g15561(.A(n17289), .Y(n18991));
  AOI22X1 g15562(.A0(n18938), .A1(P1_EBX_REG_18__SCAN_IN), .B0(n18991), .B1(n18939), .Y(n18992));
  OAI21X1 g15563(.A0(n18937), .A1(n18887), .B0(n18992), .Y(P1_U2854));
  INVX1   g15564(.A(n17315), .Y(n18994));
  AOI22X1 g15565(.A0(n18938), .A1(P1_EBX_REG_19__SCAN_IN), .B0(n18994), .B1(n18939), .Y(n18995));
  OAI21X1 g15566(.A0(n18937), .A1(n18173), .B0(n18995), .Y(P1_U2853));
  INVX1   g15567(.A(n17337), .Y(n18997));
  AOI22X1 g15568(.A0(n18938), .A1(P1_EBX_REG_20__SCAN_IN), .B0(n18997), .B1(n18939), .Y(n18998));
  OAI21X1 g15569(.A0(n18937), .A1(n18202), .B0(n18998), .Y(P1_U2852));
  INVX1   g15570(.A(n17359), .Y(n19000));
  AOI22X1 g15571(.A0(n18938), .A1(P1_EBX_REG_21__SCAN_IN), .B0(n19000), .B1(n18939), .Y(n19001));
  OAI21X1 g15572(.A0(n18937), .A1(n18245), .B0(n19001), .Y(P1_U2851));
  INVX1   g15573(.A(n17385), .Y(n19003));
  AOI22X1 g15574(.A0(n18938), .A1(P1_EBX_REG_22__SCAN_IN), .B0(n19003), .B1(n18939), .Y(n19004));
  OAI21X1 g15575(.A0(n18937), .A1(n18283), .B0(n19004), .Y(P1_U2850));
  INVX1   g15576(.A(n17416), .Y(n19006));
  AOI22X1 g15577(.A0(n18938), .A1(P1_EBX_REG_23__SCAN_IN), .B0(n19006), .B1(n18939), .Y(n19007));
  OAI21X1 g15578(.A0(n18937), .A1(n18348), .B0(n19007), .Y(P1_U2849));
  INVX1   g15579(.A(n17437), .Y(n19009));
  AOI22X1 g15580(.A0(n18938), .A1(P1_EBX_REG_24__SCAN_IN), .B0(n19009), .B1(n18939), .Y(n19010));
  OAI21X1 g15581(.A0(n18937), .A1(n18380), .B0(n19010), .Y(P1_U2848));
  INVX1   g15582(.A(n17460), .Y(n19012));
  AOI22X1 g15583(.A0(n18938), .A1(P1_EBX_REG_25__SCAN_IN), .B0(n19012), .B1(n18939), .Y(n19013));
  OAI21X1 g15584(.A0(n18937), .A1(n18412), .B0(n19013), .Y(P1_U2847));
  INVX1   g15585(.A(n17487), .Y(n19015));
  AOI22X1 g15586(.A0(n18938), .A1(P1_EBX_REG_26__SCAN_IN), .B0(n19015), .B1(n18939), .Y(n19016));
  OAI21X1 g15587(.A0(n18937), .A1(n18449), .B0(n19016), .Y(P1_U2846));
  INVX1   g15588(.A(n17511), .Y(n19018));
  AOI22X1 g15589(.A0(n18938), .A1(P1_EBX_REG_27__SCAN_IN), .B0(n19018), .B1(n18939), .Y(n19019));
  OAI21X1 g15590(.A0(n18937), .A1(n18915), .B0(n19019), .Y(P1_U2845));
  INVX1   g15591(.A(n18939), .Y(n19021));
  NOR2X1  g15592(.A(n19021), .B(n17537), .Y(n19022));
  AOI21X1 g15593(.A0(n18938), .A1(P1_EBX_REG_28__SCAN_IN), .B0(n19022), .Y(n19023));
  OAI21X1 g15594(.A0(n18937), .A1(n18523), .B0(n19023), .Y(P1_U2844));
  NOR2X1  g15595(.A(n19021), .B(n17580), .Y(n19025));
  AOI21X1 g15596(.A0(n18938), .A1(P1_EBX_REG_29__SCAN_IN), .B0(n19025), .Y(n19026));
  OAI21X1 g15597(.A0(n18937), .A1(n18555), .B0(n19026), .Y(P1_U2843));
  NOR2X1  g15598(.A(n19021), .B(n17608), .Y(n19028));
  AOI21X1 g15599(.A0(n18938), .A1(P1_EBX_REG_30__SCAN_IN), .B0(n19028), .Y(n19029));
  OAI21X1 g15600(.A0(n18937), .A1(n18591), .B0(n19029), .Y(P1_U2842));
  INVX1   g15601(.A(P1_EBX_REG_31__SCAN_IN), .Y(n19031));
  OAI22X1 g15602(.A0(n18936), .A1(n19031), .B0(n17649), .B1(n19021), .Y(P1_U2841));
  INVX1   g15603(.A(P1_EBX_REG_0__SCAN_IN), .Y(n19033));
  NOR3X1  g15604(.A(n15339), .B(n17680), .C(n14987), .Y(n19034));
  INVX1   g15605(.A(n19034), .Y(n19035));
  AOI22X1 g15606(.A0(n15123), .A1(n15030), .B0(n15007), .B1(n15237), .Y(n19036));
  AOI21X1 g15607(.A0(n19036), .A1(n19035), .B0(n15157), .Y(n19037));
  NOR4X1  g15608(.A(n16527), .B(n15341), .C(n15315), .D(n19037), .Y(n19038));
  NOR4X1  g15609(.A(n15294), .B(n14807), .C(n15155), .D(n19038), .Y(n19039));
  NOR3X1  g15610(.A(n19038), .B(n15021), .C(n15155), .Y(n19040));
  OAI21X1 g15611(.A0(n15295), .A1(n15276), .B0(n19040), .Y(n19041));
  INVX1   g15612(.A(n19041), .Y(n19042));
  AOI21X1 g15613(.A0(n19039), .A1(n19031), .B0(n19042), .Y(n19043));
  NOR3X1  g15614(.A(n19038), .B(n14807), .C(n15155), .Y(n19044));
  NOR4X1  g15615(.A(n15276), .B(n15021), .C(n15155), .D(n19038), .Y(n19045));
  OAI21X1 g15616(.A0(n19045), .A1(n19044), .B0(n15294), .Y(n19046));
  INVX1   g15617(.A(n19046), .Y(n19047));
  NAND3X1 g15618(.A(n19039), .B(n16556), .C(P1_EBX_REG_31__SCAN_IN), .Y(n19048));
  INVX1   g15619(.A(n17679), .Y(n19049));
  AOI22X1 g15620(.A0(n15001), .A1(P1_STATE2_REG_2__SCAN_IN), .B0(P1_STATE2_REG_1__SCAN_IN), .B1(n18601), .Y(n19050));
  NOR2X1  g15621(.A(n19050), .B(n19038), .Y(n19051));
  NAND2X1 g15622(.A(n19051), .B(n19049), .Y(n19052));
  NOR3X1  g15623(.A(n19038), .B(n18601), .C(n15093), .Y(n19053));
  AOI22X1 g15624(.A0(n19038), .A1(P1_REIP_REG_0__SCAN_IN), .B0(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B1(n19053), .Y(n19054));
  NOR2X1  g15625(.A(n19038), .B(n14649), .Y(n19055));
  NOR4X1  g15626(.A(n14769), .B(n14806), .C(n15155), .D(n19038), .Y(n19056));
  AOI22X1 g15627(.A0(n19055), .A1(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B0(n15131), .B1(n19056), .Y(n19057));
  NAND4X1 g15628(.A(n19054), .B(n19052), .C(n19048), .D(n19057), .Y(n19058));
  AOI21X1 g15629(.A0(n19047), .A1(P1_REIP_REG_0__SCAN_IN), .B0(n19058), .Y(n19059));
  OAI21X1 g15630(.A0(n19043), .A1(n19033), .B0(n19059), .Y(P1_U2840));
  INVX1   g15631(.A(n19043), .Y(n19061));
  NAND2X1 g15632(.A(n19061), .B(P1_EBX_REG_1__SCAN_IN), .Y(n19062));
  NAND2X1 g15633(.A(n19047), .B(n14541), .Y(n19063));
  NAND3X1 g15634(.A(n19039), .B(n16569), .C(P1_EBX_REG_31__SCAN_IN), .Y(n19064));
  AOI22X1 g15635(.A0(n19038), .A1(P1_REIP_REG_1__SCAN_IN), .B0(n17701), .B1(n19053), .Y(n19065));
  NAND2X1 g15636(.A(n19055), .B(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .Y(n19066));
  NAND2X1 g15637(.A(n19056), .B(n15168), .Y(n19067));
  NAND3X1 g15638(.A(n19067), .B(n19066), .C(n19065), .Y(n19068));
  AOI21X1 g15639(.A0(n19051), .A1(n17716), .B0(n19068), .Y(n19069));
  NAND4X1 g15640(.A(n19064), .B(n19063), .C(n19062), .D(n19069), .Y(P1_U2839));
  NAND2X1 g15641(.A(n19061), .B(P1_EBX_REG_2__SCAN_IN), .Y(n19071));
  NAND2X1 g15642(.A(n19051), .B(n17740), .Y(n19072));
  XOR2X1  g15643(.A(P1_REIP_REG_1__SCAN_IN), .B(P1_REIP_REG_2__SCAN_IN), .Y(n19073));
  NAND3X1 g15644(.A(n19039), .B(n16613), .C(P1_EBX_REG_31__SCAN_IN), .Y(n19074));
  AOI22X1 g15645(.A0(n19038), .A1(P1_REIP_REG_2__SCAN_IN), .B0(n17729), .B1(n19053), .Y(n19075));
  AOI22X1 g15646(.A0(n19055), .A1(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B0(n15802), .B1(n19056), .Y(n19076));
  NAND3X1 g15647(.A(n19076), .B(n19075), .C(n19074), .Y(n19077));
  AOI21X1 g15648(.A0(n19073), .A1(n19047), .B0(n19077), .Y(n19078));
  NAND3X1 g15649(.A(n19078), .B(n19072), .C(n19071), .Y(P1_U2838));
  INVX1   g15650(.A(n19051), .Y(n19080));
  NAND2X1 g15651(.A(P1_REIP_REG_1__SCAN_IN), .B(P1_REIP_REG_2__SCAN_IN), .Y(n19081));
  XOR2X1  g15652(.A(n19081), .B(P1_REIP_REG_3__SCAN_IN), .Y(n19082));
  NAND2X1 g15653(.A(n19039), .B(P1_EBX_REG_31__SCAN_IN), .Y(n19083));
  INVX1   g15654(.A(n19083), .Y(n19084));
  AOI22X1 g15655(.A0(n19038), .A1(P1_REIP_REG_3__SCAN_IN), .B0(n17752), .B1(n19053), .Y(n19085));
  AOI22X1 g15656(.A0(n19055), .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B0(n15218), .B1(n19056), .Y(n19086));
  NAND2X1 g15657(.A(n19086), .B(n19085), .Y(n19087));
  AOI21X1 g15658(.A0(n19084), .A1(n18946), .B0(n19087), .Y(n19088));
  OAI21X1 g15659(.A0(n19082), .A1(n19046), .B0(n19088), .Y(n19089));
  AOI21X1 g15660(.A0(n19061), .A1(P1_EBX_REG_3__SCAN_IN), .B0(n19089), .Y(n19090));
  OAI21X1 g15661(.A0(n19080), .A1(n18849), .B0(n19090), .Y(P1_U2837));
  NAND3X1 g15662(.A(P1_REIP_REG_1__SCAN_IN), .B(P1_REIP_REG_2__SCAN_IN), .C(P1_REIP_REG_3__SCAN_IN), .Y(n19092));
  XOR2X1  g15663(.A(n19092), .B(n14532), .Y(n19093));
  NAND2X1 g15664(.A(n19093), .B(n19047), .Y(n19094));
  NAND3X1 g15665(.A(n19039), .B(n18949), .C(P1_EBX_REG_31__SCAN_IN), .Y(n19095));
  INVX1   g15666(.A(n19038), .Y(n19096));
  OAI21X1 g15667(.A0(n19096), .A1(n14532), .B0(n16586), .Y(n19098));
  AOI21X1 g15668(.A0(n19055), .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B0(n19098), .Y(n19099));
  AOI22X1 g15669(.A0(n19053), .A1(n17772), .B0(n16460), .B1(n19056), .Y(n19100));
  NAND4X1 g15670(.A(n19099), .B(n19095), .C(n19094), .D(n19100), .Y(n19101));
  AOI21X1 g15671(.A0(n19061), .A1(P1_EBX_REG_4__SCAN_IN), .B0(n19101), .Y(n19102));
  OAI21X1 g15672(.A0(n19080), .A1(n17786), .B0(n19102), .Y(P1_U2836));
  NAND4X1 g15673(.A(P1_REIP_REG_2__SCAN_IN), .B(P1_REIP_REG_3__SCAN_IN), .C(P1_REIP_REG_4__SCAN_IN), .D(P1_REIP_REG_1__SCAN_IN), .Y(n19104));
  XOR2X1  g15674(.A(n19104), .B(n14529), .Y(n19105));
  NAND2X1 g15675(.A(n19105), .B(n19047), .Y(n19106));
  NAND3X1 g15676(.A(n19039), .B(n18952), .C(P1_EBX_REG_31__SCAN_IN), .Y(n19107));
  OAI21X1 g15677(.A0(n19096), .A1(n14529), .B0(n16586), .Y(n19108));
  AOI21X1 g15678(.A0(n19055), .A1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B0(n19108), .Y(n19109));
  AOI22X1 g15679(.A0(n19053), .A1(n17811), .B0(n17792), .B1(n19056), .Y(n19110));
  NAND4X1 g15680(.A(n19109), .B(n19107), .C(n19106), .D(n19110), .Y(n19111));
  AOI21X1 g15681(.A0(n19061), .A1(P1_EBX_REG_5__SCAN_IN), .B0(n19111), .Y(n19112));
  OAI21X1 g15682(.A0(n19080), .A1(n17809), .B0(n19112), .Y(P1_U2835));
  NAND3X1 g15683(.A(n19096), .B(n18601), .C(P1_STATE2_REG_1__SCAN_IN), .Y(n19114));
  NOR2X1  g15684(.A(n19104), .B(n14529), .Y(n19115));
  XOR2X1  g15685(.A(n19115), .B(P1_REIP_REG_6__SCAN_IN), .Y(n19116));
  NAND2X1 g15686(.A(n19116), .B(n19047), .Y(n19117));
  NAND3X1 g15687(.A(n19039), .B(n18955), .C(P1_EBX_REG_31__SCAN_IN), .Y(n19118));
  NAND2X1 g15688(.A(n19055), .B(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .Y(n19119));
  OAI21X1 g15689(.A0(n19096), .A1(n14526), .B0(n16586), .Y(n19120));
  AOI21X1 g15690(.A0(n19053), .A1(n17833), .B0(n19120), .Y(n19121));
  NAND4X1 g15691(.A(n19119), .B(n19118), .C(n19117), .D(n19121), .Y(n19122));
  AOI21X1 g15692(.A0(n19061), .A1(P1_EBX_REG_6__SCAN_IN), .B0(n19122), .Y(n19123));
  OAI21X1 g15693(.A0(n19114), .A1(n17831), .B0(n19123), .Y(P1_U2834));
  NOR3X1  g15694(.A(n19104), .B(n14529), .C(n14526), .Y(n19125));
  XOR2X1  g15695(.A(n19125), .B(P1_REIP_REG_7__SCAN_IN), .Y(n19126));
  NAND2X1 g15696(.A(n19126), .B(n19047), .Y(n19127));
  NAND3X1 g15697(.A(n19039), .B(n18958), .C(P1_EBX_REG_31__SCAN_IN), .Y(n19128));
  NAND2X1 g15698(.A(n19055), .B(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .Y(n19129));
  OAI21X1 g15699(.A0(n19096), .A1(n14523), .B0(n16586), .Y(n19130));
  AOI21X1 g15700(.A0(n19053), .A1(n17853), .B0(n19130), .Y(n19131));
  NAND4X1 g15701(.A(n19129), .B(n19128), .C(n19127), .D(n19131), .Y(n19132));
  AOI21X1 g15702(.A0(n19061), .A1(P1_EBX_REG_7__SCAN_IN), .B0(n19132), .Y(n19133));
  OAI21X1 g15703(.A0(n19114), .A1(n17849), .B0(n19133), .Y(P1_U2833));
  NOR4X1  g15704(.A(n14529), .B(n14526), .C(n14523), .D(n19104), .Y(n19135));
  XOR2X1  g15705(.A(n19135), .B(P1_REIP_REG_8__SCAN_IN), .Y(n19136));
  NAND2X1 g15706(.A(n19136), .B(n19047), .Y(n19137));
  NAND3X1 g15707(.A(n19039), .B(n18961), .C(P1_EBX_REG_31__SCAN_IN), .Y(n19138));
  NAND2X1 g15708(.A(n19055), .B(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .Y(n19139));
  OAI21X1 g15709(.A0(n19096), .A1(n14520), .B0(n16586), .Y(n19140));
  AOI21X1 g15710(.A0(n19053), .A1(n17878), .B0(n19140), .Y(n19141));
  NAND4X1 g15711(.A(n19139), .B(n19138), .C(n19137), .D(n19141), .Y(n19142));
  AOI21X1 g15712(.A0(n19061), .A1(P1_EBX_REG_8__SCAN_IN), .B0(n19142), .Y(n19143));
  OAI21X1 g15713(.A0(n19114), .A1(n17876), .B0(n19143), .Y(P1_U2832));
  NAND2X1 g15714(.A(n19135), .B(P1_REIP_REG_8__SCAN_IN), .Y(n19145));
  XOR2X1  g15715(.A(n19145), .B(n14517), .Y(n19146));
  NAND2X1 g15716(.A(n19146), .B(n19047), .Y(n19147));
  NAND3X1 g15717(.A(n19039), .B(n18964), .C(P1_EBX_REG_31__SCAN_IN), .Y(n19148));
  NAND2X1 g15718(.A(n19055), .B(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .Y(n19149));
  OAI21X1 g15719(.A0(n19096), .A1(n14517), .B0(n16586), .Y(n19150));
  AOI21X1 g15720(.A0(n19053), .A1(n17885), .B0(n19150), .Y(n19151));
  NAND4X1 g15721(.A(n19149), .B(n19148), .C(n19147), .D(n19151), .Y(n19152));
  AOI21X1 g15722(.A0(n19061), .A1(P1_EBX_REG_9__SCAN_IN), .B0(n19152), .Y(n19153));
  OAI21X1 g15723(.A0(n19114), .A1(n17896), .B0(n19153), .Y(P1_U2831));
  NAND3X1 g15724(.A(n19135), .B(P1_REIP_REG_8__SCAN_IN), .C(P1_REIP_REG_9__SCAN_IN), .Y(n19155));
  XOR2X1  g15725(.A(n19155), .B(n14514), .Y(n19156));
  NAND2X1 g15726(.A(n19156), .B(n19047), .Y(n19157));
  NAND3X1 g15727(.A(n19039), .B(n18967), .C(P1_EBX_REG_31__SCAN_IN), .Y(n19158));
  NAND2X1 g15728(.A(n19055), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .Y(n19159));
  OAI21X1 g15729(.A0(n19096), .A1(n14514), .B0(n16586), .Y(n19160));
  AOI21X1 g15730(.A0(n19053), .A1(n17907), .B0(n19160), .Y(n19161));
  NAND4X1 g15731(.A(n19159), .B(n19158), .C(n19157), .D(n19161), .Y(n19162));
  AOI21X1 g15732(.A0(n19061), .A1(P1_EBX_REG_10__SCAN_IN), .B0(n19162), .Y(n19163));
  OAI21X1 g15733(.A0(n19114), .A1(n17918), .B0(n19163), .Y(P1_U2830));
  NAND4X1 g15734(.A(P1_REIP_REG_8__SCAN_IN), .B(P1_REIP_REG_9__SCAN_IN), .C(P1_REIP_REG_10__SCAN_IN), .D(n19135), .Y(n19165));
  XOR2X1  g15735(.A(n19165), .B(n14511), .Y(n19166));
  NAND2X1 g15736(.A(n19166), .B(n19047), .Y(n19167));
  NAND3X1 g15737(.A(n19039), .B(n18970), .C(P1_EBX_REG_31__SCAN_IN), .Y(n19168));
  NAND2X1 g15738(.A(n19055), .B(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .Y(n19169));
  OAI21X1 g15739(.A0(n19096), .A1(n14511), .B0(n16586), .Y(n19170));
  AOI21X1 g15740(.A0(n19053), .A1(n17926), .B0(n19170), .Y(n19171));
  NAND4X1 g15741(.A(n19169), .B(n19168), .C(n19167), .D(n19171), .Y(n19172));
  AOI21X1 g15742(.A0(n19061), .A1(P1_EBX_REG_11__SCAN_IN), .B0(n19172), .Y(n19173));
  OAI21X1 g15743(.A0(n19114), .A1(n18866), .B0(n19173), .Y(P1_U2829));
  NOR2X1  g15744(.A(n19165), .B(n14511), .Y(n19175));
  XOR2X1  g15745(.A(n19175), .B(P1_REIP_REG_12__SCAN_IN), .Y(n19176));
  NAND2X1 g15746(.A(n19176), .B(n19047), .Y(n19177));
  NAND3X1 g15747(.A(n19039), .B(n18973), .C(P1_EBX_REG_31__SCAN_IN), .Y(n19178));
  NAND2X1 g15748(.A(n19055), .B(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .Y(n19179));
  OAI21X1 g15749(.A0(n19096), .A1(n14508), .B0(n16586), .Y(n19180));
  AOI21X1 g15750(.A0(n19053), .A1(n17943), .B0(n19180), .Y(n19181));
  NAND4X1 g15751(.A(n19179), .B(n19178), .C(n19177), .D(n19181), .Y(n19182));
  AOI21X1 g15752(.A0(n19061), .A1(P1_EBX_REG_12__SCAN_IN), .B0(n19182), .Y(n19183));
  OAI21X1 g15753(.A0(n19114), .A1(n17962), .B0(n19183), .Y(P1_U2828));
  NOR3X1  g15754(.A(n19165), .B(n14511), .C(n14508), .Y(n19185));
  XOR2X1  g15755(.A(n19185), .B(P1_REIP_REG_13__SCAN_IN), .Y(n19186));
  NAND2X1 g15756(.A(n19186), .B(n19047), .Y(n19187));
  NAND3X1 g15757(.A(n19039), .B(n18976), .C(P1_EBX_REG_31__SCAN_IN), .Y(n19188));
  NAND2X1 g15758(.A(n19055), .B(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .Y(n19189));
  OAI21X1 g15759(.A0(n19096), .A1(n14505), .B0(n16586), .Y(n19190));
  AOI21X1 g15760(.A0(n19053), .A1(n17969), .B0(n19190), .Y(n19191));
  NAND4X1 g15761(.A(n19189), .B(n19188), .C(n19187), .D(n19191), .Y(n19192));
  AOI21X1 g15762(.A0(n19061), .A1(P1_EBX_REG_13__SCAN_IN), .B0(n19192), .Y(n19193));
  OAI21X1 g15763(.A0(n19114), .A1(n17980), .B0(n19193), .Y(P1_U2827));
  NOR4X1  g15764(.A(n14511), .B(n14508), .C(n14505), .D(n19165), .Y(n19195));
  XOR2X1  g15765(.A(n19195), .B(P1_REIP_REG_14__SCAN_IN), .Y(n19196));
  NAND2X1 g15766(.A(n19196), .B(n19047), .Y(n19197));
  NAND3X1 g15767(.A(n19039), .B(n18979), .C(P1_EBX_REG_31__SCAN_IN), .Y(n19198));
  NAND2X1 g15768(.A(n19055), .B(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .Y(n19199));
  OAI21X1 g15769(.A0(n19096), .A1(n14502), .B0(n16586), .Y(n19200));
  AOI21X1 g15770(.A0(n19053), .A1(n17991), .B0(n19200), .Y(n19201));
  NAND4X1 g15771(.A(n19199), .B(n19198), .C(n19197), .D(n19201), .Y(n19202));
  AOI21X1 g15772(.A0(n19061), .A1(P1_EBX_REG_14__SCAN_IN), .B0(n19202), .Y(n19203));
  OAI21X1 g15773(.A0(n19114), .A1(n18003), .B0(n19203), .Y(P1_U2826));
  NAND2X1 g15774(.A(n19195), .B(P1_REIP_REG_14__SCAN_IN), .Y(n19205));
  XOR2X1  g15775(.A(n19205), .B(n14499), .Y(n19206));
  NAND2X1 g15776(.A(n19206), .B(n19047), .Y(n19207));
  NAND3X1 g15777(.A(n19039), .B(n18982), .C(P1_EBX_REG_31__SCAN_IN), .Y(n19208));
  NAND2X1 g15778(.A(n19055), .B(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .Y(n19209));
  OAI21X1 g15779(.A0(n19096), .A1(n14499), .B0(n16586), .Y(n19210));
  AOI21X1 g15780(.A0(n19053), .A1(n18011), .B0(n19210), .Y(n19211));
  NAND4X1 g15781(.A(n19209), .B(n19208), .C(n19207), .D(n19211), .Y(n19212));
  AOI21X1 g15782(.A0(n19061), .A1(P1_EBX_REG_15__SCAN_IN), .B0(n19212), .Y(n19213));
  OAI21X1 g15783(.A0(n19114), .A1(n18875), .B0(n19213), .Y(P1_U2825));
  NAND3X1 g15784(.A(n19195), .B(P1_REIP_REG_14__SCAN_IN), .C(P1_REIP_REG_15__SCAN_IN), .Y(n19215));
  XOR2X1  g15785(.A(n19215), .B(n14496), .Y(n19216));
  NAND2X1 g15786(.A(n19216), .B(n19047), .Y(n19217));
  NAND3X1 g15787(.A(n19039), .B(n18985), .C(P1_EBX_REG_31__SCAN_IN), .Y(n19218));
  NAND2X1 g15788(.A(n19055), .B(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .Y(n19219));
  OAI21X1 g15789(.A0(n19096), .A1(n14496), .B0(n16586), .Y(n19220));
  AOI21X1 g15790(.A0(n19053), .A1(n18032), .B0(n19220), .Y(n19221));
  NAND4X1 g15791(.A(n19219), .B(n19218), .C(n19217), .D(n19221), .Y(n19222));
  AOI21X1 g15792(.A0(n19061), .A1(P1_EBX_REG_16__SCAN_IN), .B0(n19222), .Y(n19223));
  OAI21X1 g15793(.A0(n19114), .A1(n18080), .B0(n19223), .Y(P1_U2824));
  NAND4X1 g15794(.A(P1_REIP_REG_14__SCAN_IN), .B(P1_REIP_REG_15__SCAN_IN), .C(P1_REIP_REG_16__SCAN_IN), .D(n19195), .Y(n19225));
  XOR2X1  g15795(.A(n19225), .B(n14493), .Y(n19226));
  NAND2X1 g15796(.A(n19226), .B(n19047), .Y(n19227));
  NAND3X1 g15797(.A(n19039), .B(n18988), .C(P1_EBX_REG_31__SCAN_IN), .Y(n19228));
  NAND2X1 g15798(.A(n19055), .B(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .Y(n19229));
  OAI21X1 g15799(.A0(n19096), .A1(n14493), .B0(n16586), .Y(n19230));
  AOI21X1 g15800(.A0(n19053), .A1(n18090), .B0(n19230), .Y(n19231));
  NAND4X1 g15801(.A(n19229), .B(n19228), .C(n19227), .D(n19231), .Y(n19232));
  AOI21X1 g15802(.A0(n19061), .A1(P1_EBX_REG_17__SCAN_IN), .B0(n19232), .Y(n19233));
  OAI21X1 g15803(.A0(n19114), .A1(n18108), .B0(n19233), .Y(P1_U2823));
  NOR2X1  g15804(.A(n19225), .B(n14493), .Y(n19235));
  XOR2X1  g15805(.A(n19235), .B(P1_REIP_REG_18__SCAN_IN), .Y(n19236));
  NAND2X1 g15806(.A(n19236), .B(n19047), .Y(n19237));
  NAND3X1 g15807(.A(n19039), .B(n18991), .C(P1_EBX_REG_31__SCAN_IN), .Y(n19238));
  NAND2X1 g15808(.A(n19055), .B(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .Y(n19239));
  OAI21X1 g15809(.A0(n19096), .A1(n14490), .B0(n16586), .Y(n19240));
  AOI21X1 g15810(.A0(n19053), .A1(n18118), .B0(n19240), .Y(n19241));
  NAND4X1 g15811(.A(n19239), .B(n19238), .C(n19237), .D(n19241), .Y(n19242));
  AOI21X1 g15812(.A0(n19061), .A1(P1_EBX_REG_18__SCAN_IN), .B0(n19242), .Y(n19243));
  OAI21X1 g15813(.A0(n19114), .A1(n18887), .B0(n19243), .Y(P1_U2822));
  NOR3X1  g15814(.A(n19225), .B(n14493), .C(n14490), .Y(n19245));
  XOR2X1  g15815(.A(n19245), .B(P1_REIP_REG_19__SCAN_IN), .Y(n19246));
  NAND2X1 g15816(.A(n19246), .B(n19047), .Y(n19247));
  NAND3X1 g15817(.A(n19039), .B(n18994), .C(P1_EBX_REG_31__SCAN_IN), .Y(n19248));
  NAND2X1 g15818(.A(n19055), .B(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .Y(n19249));
  OAI21X1 g15819(.A0(n19096), .A1(n14487), .B0(n16586), .Y(n19250));
  AOI21X1 g15820(.A0(n19053), .A1(n18149), .B0(n19250), .Y(n19251));
  NAND4X1 g15821(.A(n19249), .B(n19248), .C(n19247), .D(n19251), .Y(n19252));
  AOI21X1 g15822(.A0(n19061), .A1(P1_EBX_REG_19__SCAN_IN), .B0(n19252), .Y(n19253));
  OAI21X1 g15823(.A0(n19114), .A1(n18173), .B0(n19253), .Y(P1_U2821));
  NOR4X1  g15824(.A(n14493), .B(n14490), .C(n14487), .D(n19225), .Y(n19255));
  XOR2X1  g15825(.A(n19255), .B(P1_REIP_REG_20__SCAN_IN), .Y(n19256));
  NAND2X1 g15826(.A(n19256), .B(n19047), .Y(n19257));
  NAND3X1 g15827(.A(n19039), .B(n18997), .C(P1_EBX_REG_31__SCAN_IN), .Y(n19258));
  INVX1   g15828(.A(n19053), .Y(n19259));
  OAI22X1 g15829(.A0(n19096), .A1(n14484), .B0(n18181), .B1(n19259), .Y(n19260));
  AOI21X1 g15830(.A0(n19055), .A1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B0(n19260), .Y(n19261));
  NAND3X1 g15831(.A(n19261), .B(n19258), .C(n19257), .Y(n19262));
  AOI21X1 g15832(.A0(n19061), .A1(P1_EBX_REG_20__SCAN_IN), .B0(n19262), .Y(n19263));
  OAI21X1 g15833(.A0(n19114), .A1(n18202), .B0(n19263), .Y(P1_U2820));
  NAND2X1 g15834(.A(n19255), .B(P1_REIP_REG_20__SCAN_IN), .Y(n19265));
  XOR2X1  g15835(.A(n19265), .B(n14481), .Y(n19266));
  NAND2X1 g15836(.A(n19266), .B(n19047), .Y(n19267));
  NAND3X1 g15837(.A(n19039), .B(n19000), .C(P1_EBX_REG_31__SCAN_IN), .Y(n19268));
  OAI22X1 g15838(.A0(n19096), .A1(n14481), .B0(n18209), .B1(n19259), .Y(n19269));
  AOI21X1 g15839(.A0(n19055), .A1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B0(n19269), .Y(n19270));
  NAND3X1 g15840(.A(n19270), .B(n19268), .C(n19267), .Y(n19271));
  AOI21X1 g15841(.A0(n19061), .A1(P1_EBX_REG_21__SCAN_IN), .B0(n19271), .Y(n19272));
  OAI21X1 g15842(.A0(n19114), .A1(n18245), .B0(n19272), .Y(P1_U2819));
  NAND3X1 g15843(.A(n19255), .B(P1_REIP_REG_20__SCAN_IN), .C(P1_REIP_REG_21__SCAN_IN), .Y(n19274));
  XOR2X1  g15844(.A(n19274), .B(n14478), .Y(n19275));
  NAND2X1 g15845(.A(n19275), .B(n19047), .Y(n19276));
  NAND3X1 g15846(.A(n19039), .B(n19003), .C(P1_EBX_REG_31__SCAN_IN), .Y(n19277));
  OAI22X1 g15847(.A0(n19096), .A1(n14478), .B0(n18253), .B1(n19259), .Y(n19278));
  AOI21X1 g15848(.A0(n19055), .A1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B0(n19278), .Y(n19279));
  NAND3X1 g15849(.A(n19279), .B(n19277), .C(n19276), .Y(n19280));
  AOI21X1 g15850(.A0(n19061), .A1(P1_EBX_REG_22__SCAN_IN), .B0(n19280), .Y(n19281));
  OAI21X1 g15851(.A0(n19114), .A1(n18283), .B0(n19281), .Y(P1_U2818));
  NAND4X1 g15852(.A(P1_REIP_REG_20__SCAN_IN), .B(P1_REIP_REG_21__SCAN_IN), .C(P1_REIP_REG_22__SCAN_IN), .D(n19255), .Y(n19283));
  XOR2X1  g15853(.A(n19283), .B(P1_REIP_REG_23__SCAN_IN), .Y(n19284));
  NAND2X1 g15854(.A(n19055), .B(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .Y(n19285));
  AOI22X1 g15855(.A0(n19038), .A1(P1_REIP_REG_23__SCAN_IN), .B0(n18292), .B1(n19053), .Y(n19286));
  NAND2X1 g15856(.A(n19286), .B(n19285), .Y(n19287));
  AOI21X1 g15857(.A0(n19084), .A1(n19006), .B0(n19287), .Y(n19288));
  OAI21X1 g15858(.A0(n19284), .A1(n19046), .B0(n19288), .Y(n19289));
  AOI21X1 g15859(.A0(n19061), .A1(P1_EBX_REG_23__SCAN_IN), .B0(n19289), .Y(n19290));
  OAI21X1 g15860(.A0(n19114), .A1(n18348), .B0(n19290), .Y(P1_U2817));
  NOR2X1  g15861(.A(n19283), .B(n14475), .Y(n19292));
  XOR2X1  g15862(.A(n19292), .B(P1_REIP_REG_24__SCAN_IN), .Y(n19293));
  NAND2X1 g15863(.A(n19293), .B(n19047), .Y(n19294));
  NAND2X1 g15864(.A(n19084), .B(n19009), .Y(n19295));
  OAI22X1 g15865(.A0(n19096), .A1(n14472), .B0(n18356), .B1(n19259), .Y(n19296));
  AOI21X1 g15866(.A0(n19055), .A1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B0(n19296), .Y(n19297));
  NAND3X1 g15867(.A(n19297), .B(n19295), .C(n19294), .Y(n19298));
  AOI21X1 g15868(.A0(n19061), .A1(P1_EBX_REG_24__SCAN_IN), .B0(n19298), .Y(n19299));
  OAI21X1 g15869(.A0(n19114), .A1(n18380), .B0(n19299), .Y(P1_U2816));
  NOR3X1  g15870(.A(n19283), .B(n14475), .C(n14472), .Y(n19301));
  XOR2X1  g15871(.A(n19301), .B(n14469), .Y(n19302));
  NAND2X1 g15872(.A(n19055), .B(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .Y(n19303));
  AOI22X1 g15873(.A0(n19038), .A1(P1_REIP_REG_25__SCAN_IN), .B0(n18388), .B1(n19053), .Y(n19304));
  NAND2X1 g15874(.A(n19304), .B(n19303), .Y(n19305));
  AOI21X1 g15875(.A0(n19084), .A1(n19012), .B0(n19305), .Y(n19306));
  OAI21X1 g15876(.A0(n19302), .A1(n19046), .B0(n19306), .Y(n19307));
  AOI21X1 g15877(.A0(n19061), .A1(P1_EBX_REG_25__SCAN_IN), .B0(n19307), .Y(n19308));
  OAI21X1 g15878(.A0(n19114), .A1(n18412), .B0(n19308), .Y(P1_U2815));
  NOR4X1  g15879(.A(n14475), .B(n14472), .C(n14469), .D(n19283), .Y(n19310));
  XOR2X1  g15880(.A(n19310), .B(P1_REIP_REG_26__SCAN_IN), .Y(n19311));
  NAND2X1 g15881(.A(n19311), .B(n19047), .Y(n19312));
  NAND2X1 g15882(.A(n19084), .B(n19015), .Y(n19313));
  NAND2X1 g15883(.A(n19055), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .Y(n19314));
  AOI22X1 g15884(.A0(n19038), .A1(P1_REIP_REG_26__SCAN_IN), .B0(n18421), .B1(n19053), .Y(n19315));
  NAND4X1 g15885(.A(n19314), .B(n19313), .C(n19312), .D(n19315), .Y(n19316));
  AOI21X1 g15886(.A0(n19061), .A1(P1_EBX_REG_26__SCAN_IN), .B0(n19316), .Y(n19317));
  OAI21X1 g15887(.A0(n19114), .A1(n18449), .B0(n19317), .Y(P1_U2814));
  NAND2X1 g15888(.A(n19310), .B(P1_REIP_REG_26__SCAN_IN), .Y(n19319));
  XOR2X1  g15889(.A(n19319), .B(n14463), .Y(n19320));
  NAND2X1 g15890(.A(n19320), .B(n19047), .Y(n19321));
  NAND2X1 g15891(.A(n19084), .B(n19018), .Y(n19322));
  OAI22X1 g15892(.A0(n19096), .A1(n14463), .B0(n18457), .B1(n19259), .Y(n19323));
  AOI21X1 g15893(.A0(n19055), .A1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B0(n19323), .Y(n19324));
  NAND3X1 g15894(.A(n19324), .B(n19322), .C(n19321), .Y(n19325));
  AOI21X1 g15895(.A0(n19061), .A1(P1_EBX_REG_27__SCAN_IN), .B0(n19325), .Y(n19326));
  OAI21X1 g15896(.A0(n19114), .A1(n18915), .B0(n19326), .Y(P1_U2813));
  INVX1   g15897(.A(P1_EBX_REG_28__SCAN_IN), .Y(n19328));
  NOR2X1  g15898(.A(n19043), .B(n19328), .Y(n19329));
  NOR2X1  g15899(.A(n19083), .B(n17537), .Y(n19330));
  NAND3X1 g15900(.A(n19310), .B(P1_REIP_REG_26__SCAN_IN), .C(P1_REIP_REG_27__SCAN_IN), .Y(n19331));
  XOR2X1  g15901(.A(n19331), .B(P1_REIP_REG_28__SCAN_IN), .Y(n19332));
  OAI22X1 g15902(.A0(n19096), .A1(n14460), .B0(n18491), .B1(n19259), .Y(n19333));
  AOI21X1 g15903(.A0(n19055), .A1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B0(n19333), .Y(n19334));
  OAI21X1 g15904(.A0(n19332), .A1(n19046), .B0(n19334), .Y(n19335));
  NOR3X1  g15905(.A(n19335), .B(n19330), .C(n19329), .Y(n19336));
  OAI21X1 g15906(.A0(n19114), .A1(n18523), .B0(n19336), .Y(P1_U2812));
  NOR2X1  g15907(.A(n19083), .B(n17580), .Y(n19338));
  INVX1   g15908(.A(P1_EBX_REG_29__SCAN_IN), .Y(n19339));
  NOR2X1  g15909(.A(n19043), .B(n19339), .Y(n19340));
  NAND4X1 g15910(.A(P1_REIP_REG_26__SCAN_IN), .B(P1_REIP_REG_27__SCAN_IN), .C(P1_REIP_REG_28__SCAN_IN), .D(n19310), .Y(n19341));
  XOR2X1  g15911(.A(n19341), .B(P1_REIP_REG_29__SCAN_IN), .Y(n19342));
  OAI22X1 g15912(.A0(n19096), .A1(n14457), .B0(n18530), .B1(n19259), .Y(n19343));
  AOI21X1 g15913(.A0(n19055), .A1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B0(n19343), .Y(n19344));
  OAI21X1 g15914(.A0(n19342), .A1(n19046), .B0(n19344), .Y(n19345));
  NOR3X1  g15915(.A(n19345), .B(n19340), .C(n19338), .Y(n19346));
  OAI21X1 g15916(.A0(n19114), .A1(n18555), .B0(n19346), .Y(P1_U2811));
  NOR2X1  g15917(.A(n19083), .B(n17608), .Y(n19348));
  INVX1   g15918(.A(P1_EBX_REG_30__SCAN_IN), .Y(n19349));
  NOR2X1  g15919(.A(n19043), .B(n19349), .Y(n19350));
  NOR2X1  g15920(.A(n19341), .B(n14457), .Y(n19351));
  XOR2X1  g15921(.A(n19351), .B(n14452), .Y(n19352));
  OAI22X1 g15922(.A0(n19096), .A1(n14452), .B0(n18567), .B1(n19259), .Y(n19353));
  AOI21X1 g15923(.A0(n19055), .A1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B0(n19353), .Y(n19354));
  OAI21X1 g15924(.A0(n19352), .A1(n19046), .B0(n19354), .Y(n19355));
  NOR3X1  g15925(.A(n19355), .B(n19350), .C(n19348), .Y(n19356));
  OAI21X1 g15926(.A0(n19114), .A1(n18591), .B0(n19356), .Y(P1_U2810));
  NOR2X1  g15927(.A(n19083), .B(n17649), .Y(n19358));
  NOR2X1  g15928(.A(n19043), .B(n19031), .Y(n19359));
  NOR3X1  g15929(.A(n19341), .B(n14457), .C(n14452), .Y(n19360));
  XOR2X1  g15930(.A(n19360), .B(n18619), .Y(n19361));
  OAI22X1 g15931(.A0(n19096), .A1(n18619), .B0(n18600), .B1(n19259), .Y(n19362));
  AOI21X1 g15932(.A0(n19055), .A1(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B0(n19362), .Y(n19363));
  OAI21X1 g15933(.A0(n19361), .A1(n19046), .B0(n19363), .Y(n19364));
  NOR3X1  g15934(.A(n19364), .B(n19359), .C(n19358), .Y(n19365));
  OAI21X1 g15935(.A0(n19114), .A1(n18618), .B0(n19365), .Y(P1_U2809));
  NOR4X1  g15936(.A(P1_DATAWIDTH_REG_15__SCAN_IN), .B(P1_DATAWIDTH_REG_14__SCAN_IN), .C(P1_DATAWIDTH_REG_13__SCAN_IN), .D(P1_DATAWIDTH_REG_16__SCAN_IN), .Y(n19367));
  NOR4X1  g15937(.A(P1_DATAWIDTH_REG_12__SCAN_IN), .B(P1_DATAWIDTH_REG_11__SCAN_IN), .C(P1_DATAWIDTH_REG_10__SCAN_IN), .D(P1_DATAWIDTH_REG_26__SCAN_IN), .Y(n19368));
  NOR4X1  g15938(.A(P1_DATAWIDTH_REG_7__SCAN_IN), .B(P1_DATAWIDTH_REG_6__SCAN_IN), .C(P1_DATAWIDTH_REG_5__SCAN_IN), .D(P1_DATAWIDTH_REG_8__SCAN_IN), .Y(n19369));
  NOR4X1  g15939(.A(P1_DATAWIDTH_REG_4__SCAN_IN), .B(P1_DATAWIDTH_REG_3__SCAN_IN), .C(P1_DATAWIDTH_REG_2__SCAN_IN), .D(P1_DATAWIDTH_REG_17__SCAN_IN), .Y(n19370));
  NAND4X1 g15940(.A(n19369), .B(n19368), .C(n19367), .D(n19370), .Y(n19371));
  NOR4X1  g15941(.A(P1_DATAWIDTH_REG_22__SCAN_IN), .B(P1_DATAWIDTH_REG_21__SCAN_IN), .C(P1_DATAWIDTH_REG_20__SCAN_IN), .D(P1_DATAWIDTH_REG_23__SCAN_IN), .Y(n19372));
  INVX1   g15942(.A(P1_DATAWIDTH_REG_0__SCAN_IN), .Y(n19373));
  NOR2X1  g15943(.A(n14585), .B(n19373), .Y(n19374));
  NOR3X1  g15944(.A(n19374), .B(P1_DATAWIDTH_REG_19__SCAN_IN), .C(P1_DATAWIDTH_REG_18__SCAN_IN), .Y(n19375));
  NOR4X1  g15945(.A(P1_DATAWIDTH_REG_29__SCAN_IN), .B(P1_DATAWIDTH_REG_28__SCAN_IN), .C(P1_DATAWIDTH_REG_27__SCAN_IN), .D(P1_DATAWIDTH_REG_30__SCAN_IN), .Y(n19376));
  NOR4X1  g15946(.A(P1_DATAWIDTH_REG_25__SCAN_IN), .B(P1_DATAWIDTH_REG_24__SCAN_IN), .C(P1_DATAWIDTH_REG_9__SCAN_IN), .D(P1_DATAWIDTH_REG_31__SCAN_IN), .Y(n19377));
  NAND4X1 g15947(.A(n19376), .B(n19375), .C(n19372), .D(n19377), .Y(n19378));
  NOR2X1  g15948(.A(n19378), .B(n19371), .Y(n19379));
  NAND3X1 g15949(.A(n19379), .B(n14585), .C(n14541), .Y(n19380));
  NOR2X1  g15950(.A(P1_DATAWIDTH_REG_1__SCAN_IN), .B(P1_DATAWIDTH_REG_0__SCAN_IN), .Y(n19381));
  NAND3X1 g15951(.A(n19381), .B(n19379), .C(n17690), .Y(n19382));
  OAI21X1 g15952(.A0(n19378), .A1(n19371), .B0(P1_BYTEENABLE_REG_3__SCAN_IN), .Y(n19383));
  NAND3X1 g15953(.A(n19383), .B(n19382), .C(n19380), .Y(P1_U2808));
  NAND2X1 g15954(.A(P1_REIP_REG_0__SCAN_IN), .B(P1_REIP_REG_1__SCAN_IN), .Y(n19385));
  AOI21X1 g15955(.A0(P1_DATAWIDTH_REG_0__SCAN_IN), .A1(n17690), .B0(n19381), .Y(n19386));
  OAI21X1 g15956(.A0(n19386), .A1(P1_REIP_REG_1__SCAN_IN), .B0(n19385), .Y(n19387));
  NAND2X1 g15957(.A(n19387), .B(n19379), .Y(n19388));
  OAI21X1 g15958(.A0(n19379), .A1(n14441), .B0(n19388), .Y(P1_U3481));
  NAND2X1 g15959(.A(n19379), .B(P1_REIP_REG_1__SCAN_IN), .Y(n19390));
  OAI21X1 g15960(.A0(n19378), .A1(n19371), .B0(P1_BYTEENABLE_REG_1__SCAN_IN), .Y(n19391));
  NAND3X1 g15961(.A(n19391), .B(n19390), .C(n19382), .Y(P1_U2807));
  OAI21X1 g15962(.A0(P1_REIP_REG_0__SCAN_IN), .A1(P1_REIP_REG_1__SCAN_IN), .B0(n19379), .Y(n19393));
  OAI21X1 g15963(.A0(n19379), .A1(n14449), .B0(n19393), .Y(P1_U3482));
  OAI21X1 g15964(.A0(P1_STATE_REG_0__SCAN_IN), .A1(n14438), .B0(P1_W_R_N_REG_SCAN_IN), .Y(n19395));
  OAI21X1 g15965(.A0(n14443), .A1(P1_READREQUEST_REG_SCAN_IN), .B0(n19395), .Y(P1_U3483));
  NOR2X1  g15966(.A(n15339), .B(n15278), .Y(n19397));
  OAI21X1 g15967(.A0(n19397), .A1(n15322), .B0(n17683), .Y(P1_U2806));
  NAND2X1 g15968(.A(n19397), .B(n15288), .Y(n19399));
  OAI21X1 g15969(.A0(n15339), .A1(n15278), .B0(P1_MORE_REG_SCAN_IN), .Y(n19400));
  NAND2X1 g15970(.A(n19400), .B(n19399), .Y(P1_U3484));
  AOI22X1 g15971(.A0(n14559), .A1(n14436), .B0(P1_STATEBS16_REG_SCAN_IN), .B1(n14582), .Y(n19402));
  OAI21X1 g15972(.A0(n14582), .A1(n3439), .B0(n19402), .Y(P1_U2805));
  OAI21X1 g15973(.A0(n15276), .A1(n15305), .B0(n15020), .Y(n19404));
  NAND3X1 g15974(.A(n19404), .B(n14550), .C(P1_STATE2_REG_2__SCAN_IN), .Y(n19405));
  OAI22X1 g15975(.A0(n15106), .A1(n15275), .B0(P1_STATE2_REG_1__SCAN_IN), .B1(P1_STATE2_REG_2__SCAN_IN), .Y(n19406));
  AOI21X1 g15976(.A0(n19405), .A1(P1_STATE2_REG_0__SCAN_IN), .B0(n19406), .Y(n19407));
  NOR4X1  g15977(.A(P1_STATE2_REG_0__SCAN_IN), .B(n15093), .C(n15155), .D(n14549), .Y(n19408));
  NOR4X1  g15978(.A(n19037), .B(n16508), .C(n15095), .D(n19408), .Y(n19409));
  NAND2X1 g15979(.A(n19409), .B(P1_REQUESTPENDING_REG_SCAN_IN), .Y(n19410));
  OAI21X1 g15980(.A0(n19409), .A1(n19407), .B0(n19410), .Y(P1_U3485));
  OAI21X1 g15981(.A0(P1_STATE_REG_0__SCAN_IN), .A1(n14438), .B0(P1_D_C_N_REG_SCAN_IN), .Y(n19412));
  NOR3X1  g15982(.A(P1_STATE_REG_0__SCAN_IN), .B(n14438), .C(P1_CODEFETCH_REG_SCAN_IN), .Y(n19413));
  AOI21X1 g15983(.A0(n14559), .A1(n14436), .B0(n19413), .Y(n19414));
  NAND2X1 g15984(.A(n19414), .B(n19412), .Y(P1_U2804));
  NAND3X1 g15985(.A(n14436), .B(P1_STATE_REG_1__SCAN_IN), .C(P1_MEMORYFETCH_REG_SCAN_IN), .Y(n19416));
  OAI21X1 g15986(.A0(P1_STATE_REG_0__SCAN_IN), .A1(n14438), .B0(P1_M_IO_N_REG_SCAN_IN), .Y(n19417));
  NAND2X1 g15987(.A(n19417), .B(n19416), .Y(P1_U3486));
  NAND2X1 g15988(.A(n16508), .B(n15093), .Y(n19419));
  OAI21X1 g15989(.A0(n15339), .A1(n15274), .B0(P1_CODEFETCH_REG_SCAN_IN), .Y(n19420));
  OAI21X1 g15990(.A0(n19419), .A1(n14650), .B0(n19420), .Y(P1_U2803));
  NAND2X1 g15991(.A(P1_STATE_REG_0__SCAN_IN), .B(P1_ADS_N_REG_SCAN_IN), .Y(n19422));
  NAND2X1 g15992(.A(n19422), .B(n14582), .Y(P1_U2802));
  NOR3X1  g15993(.A(n15008), .B(n15001), .C(n15155), .Y(n19424));
  AOI21X1 g15994(.A0(n16508), .A1(n15093), .B0(n19037), .Y(n19425));
  NAND2X1 g15995(.A(n19425), .B(P1_READREQUEST_REG_SCAN_IN), .Y(n19426));
  OAI21X1 g15996(.A0(n19425), .A1(n19424), .B0(n19426), .Y(P1_U3487));
  NOR2X1  g15997(.A(n15272), .B(n15137), .Y(n19428));
  NAND3X1 g15998(.A(n19428), .B(n15156), .C(n14824), .Y(n19429));
  OAI21X1 g15999(.A0(n19429), .A1(n15270), .B0(P1_MEMORYFETCH_REG_SCAN_IN), .Y(n19430));
  NAND3X1 g16000(.A(n19430), .B(n19419), .C(n19035), .Y(P1_U2801));
endmodule


