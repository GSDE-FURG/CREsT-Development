// Benchmark "top" written by ABC on Wed Sep 29 17:25:37 2021

module top ( 
    \A[0] , \A[1] , \A[2] , \A[3] , \A[4] , \A[5] , \A[6] , \A[7] , \A[8] ,
    \A[9] , \A[10] , \A[11] , \A[12] , \A[13] , \A[14] , \A[15] , \A[16] ,
    \A[17] , \A[18] , \A[19] , \A[20] , \A[21] , \A[22] , \A[23] , \A[24] ,
    \A[25] , \A[26] , \A[27] , \A[28] , \A[29] , \A[30] , \A[31] , \A[32] ,
    \A[33] , \A[34] , \A[35] , \A[36] , \A[37] , \A[38] , \A[39] , \A[40] ,
    \A[41] , \A[42] , \A[43] , \A[44] , \A[45] , \A[46] , \A[47] , \A[48] ,
    \A[49] , \A[50] , \A[51] , \A[52] , \A[53] , \A[54] , \A[55] , \A[56] ,
    \A[57] , \A[58] , \A[59] , \A[60] , \A[61] , \A[62] , \A[63] , \A[64] ,
    \A[65] , \A[66] , \A[67] , \A[68] , \A[69] , \A[70] , \A[71] , \A[72] ,
    \A[73] , \A[74] , \A[75] , \A[76] , \A[77] , \A[78] , \A[79] , \A[80] ,
    \A[81] , \A[82] , \A[83] , \A[84] , \A[85] , \A[86] , \A[87] , \A[88] ,
    \A[89] , \A[90] , \A[91] , \A[92] , \A[93] , \A[94] , \A[95] , \A[96] ,
    \A[97] , \A[98] , \A[99] , \A[100] , \A[101] , \A[102] , \A[103] ,
    \A[104] , \A[105] , \A[106] , \A[107] , \A[108] , \A[109] , \A[110] ,
    \A[111] , \A[112] , \A[113] , \A[114] , \A[115] , \A[116] , \A[117] ,
    \A[118] , \A[119] , \A[120] , \A[121] , \A[122] , \A[123] , \A[124] ,
    \A[125] , \A[126] , \A[127] , \A[128] , \A[129] , \A[130] , \A[131] ,
    \A[132] , \A[133] , \A[134] , \A[135] , \A[136] , \A[137] , \A[138] ,
    \A[139] , \A[140] , \A[141] , \A[142] , \A[143] , \A[144] , \A[145] ,
    \A[146] , \A[147] , \A[148] , \A[149] , \A[150] , \A[151] , \A[152] ,
    \A[153] , \A[154] , \A[155] , \A[156] , \A[157] , \A[158] , \A[159] ,
    \A[160] , \A[161] , \A[162] , \A[163] , \A[164] , \A[165] , \A[166] ,
    \A[167] , \A[168] , \A[169] , \A[170] , \A[171] , \A[172] , \A[173] ,
    \A[174] , \A[175] , \A[176] , \A[177] , \A[178] , \A[179] , \A[180] ,
    \A[181] , \A[182] , \A[183] , \A[184] , \A[185] , \A[186] , \A[187] ,
    \A[188] , \A[189] , \A[190] , \A[191] , \A[192] , \A[193] , \A[194] ,
    \A[195] , \A[196] , \A[197] , \A[198] , \A[199] , \A[200] , \A[201] ,
    \A[202] , \A[203] , \A[204] , \A[205] , \A[206] , \A[207] , \A[208] ,
    \A[209] , \A[210] , \A[211] , \A[212] , \A[213] , \A[214] , \A[215] ,
    \A[216] , \A[217] , \A[218] , \A[219] , \A[220] , \A[221] , \A[222] ,
    \A[223] , \A[224] , \A[225] , \A[226] , \A[227] , \A[228] , \A[229] ,
    \A[230] , \A[231] , \A[232] , \A[233] , \A[234] , \A[235] , \A[236] ,
    \A[237] , \A[238] , \A[239] , \A[240] , \A[241] , \A[242] , \A[243] ,
    \A[244] , \A[245] , \A[246] , \A[247] , \A[248] , \A[249] , \A[250] ,
    \A[251] , \A[252] , \A[253] , \A[254] , \A[255] , \A[256] , \A[257] ,
    \A[258] , \A[259] , \A[260] , \A[261] , \A[262] , \A[263] , \A[264] ,
    \A[265] , \A[266] , \A[267] , \A[268] , \A[269] , \A[270] , \A[271] ,
    \A[272] , \A[273] , \A[274] , \A[275] , \A[276] , \A[277] , \A[278] ,
    \A[279] , \A[280] , \A[281] , \A[282] , \A[283] , \A[284] , \A[285] ,
    \A[286] , \A[287] , \A[288] , \A[289] , \A[290] , \A[291] , \A[292] ,
    \A[293] , \A[294] , \A[295] , \A[296] , \A[297] , \A[298] , \A[299] ,
    \A[300] , \A[301] , \A[302] , \A[303] , \A[304] , \A[305] , \A[306] ,
    \A[307] , \A[308] , \A[309] , \A[310] , \A[311] , \A[312] , \A[313] ,
    \A[314] , \A[315] , \A[316] , \A[317] , \A[318] , \A[319] , \A[320] ,
    \A[321] , \A[322] , \A[323] , \A[324] , \A[325] , \A[326] , \A[327] ,
    \A[328] , \A[329] , \A[330] , \A[331] , \A[332] , \A[333] , \A[334] ,
    \A[335] , \A[336] , \A[337] , \A[338] , \A[339] , \A[340] , \A[341] ,
    \A[342] , \A[343] , \A[344] , \A[345] , \A[346] , \A[347] , \A[348] ,
    \A[349] , \A[350] , \A[351] , \A[352] , \A[353] , \A[354] , \A[355] ,
    \A[356] , \A[357] , \A[358] , \A[359] , \A[360] , \A[361] , \A[362] ,
    \A[363] , \A[364] , \A[365] , \A[366] , \A[367] , \A[368] , \A[369] ,
    \A[370] , \A[371] , \A[372] , \A[373] , \A[374] , \A[375] , \A[376] ,
    \A[377] , \A[378] , \A[379] , \A[380] , \A[381] , \A[382] , \A[383] ,
    \A[384] , \A[385] , \A[386] , \A[387] , \A[388] , \A[389] , \A[390] ,
    \A[391] , \A[392] , \A[393] , \A[394] , \A[395] , \A[396] , \A[397] ,
    \A[398] , \A[399] , \A[400] , \A[401] , \A[402] , \A[403] , \A[404] ,
    \A[405] , \A[406] , \A[407] , \A[408] , \A[409] , \A[410] , \A[411] ,
    \A[412] , \A[413] , \A[414] , \A[415] , \A[416] , \A[417] , \A[418] ,
    \A[419] , \A[420] , \A[421] , \A[422] , \A[423] , \A[424] , \A[425] ,
    \A[426] , \A[427] , \A[428] , \A[429] , \A[430] , \A[431] , \A[432] ,
    \A[433] , \A[434] , \A[435] , \A[436] , \A[437] , \A[438] , \A[439] ,
    \A[440] , \A[441] , \A[442] , \A[443] , \A[444] , \A[445] , \A[446] ,
    \A[447] , \A[448] , \A[449] , \A[450] , \A[451] , \A[452] , \A[453] ,
    \A[454] , \A[455] , \A[456] , \A[457] , \A[458] , \A[459] , \A[460] ,
    \A[461] , \A[462] , \A[463] , \A[464] , \A[465] , \A[466] , \A[467] ,
    \A[468] , \A[469] , \A[470] , \A[471] , \A[472] , \A[473] , \A[474] ,
    \A[475] , \A[476] , \A[477] , \A[478] , \A[479] , \A[480] , \A[481] ,
    \A[482] , \A[483] , \A[484] , \A[485] , \A[486] , \A[487] , \A[488] ,
    \A[489] , \A[490] , \A[491] , \A[492] , \A[493] , \A[494] , \A[495] ,
    \A[496] , \A[497] , \A[498] , \A[499] , \A[500] , \A[501] , \A[502] ,
    \A[503] , \A[504] , \A[505] , \A[506] , \A[507] , \A[508] , \A[509] ,
    \A[510] , \A[511] , \A[512] , \A[513] , \A[514] , \A[515] , \A[516] ,
    \A[517] , \A[518] , \A[519] , \A[520] , \A[521] , \A[522] , \A[523] ,
    \A[524] , \A[525] , \A[526] , \A[527] , \A[528] , \A[529] , \A[530] ,
    \A[531] , \A[532] , \A[533] , \A[534] , \A[535] , \A[536] , \A[537] ,
    \A[538] , \A[539] , \A[540] , \A[541] , \A[542] , \A[543] , \A[544] ,
    \A[545] , \A[546] , \A[547] , \A[548] , \A[549] , \A[550] , \A[551] ,
    \A[552] , \A[553] , \A[554] , \A[555] , \A[556] , \A[557] , \A[558] ,
    \A[559] , \A[560] , \A[561] , \A[562] , \A[563] , \A[564] , \A[565] ,
    \A[566] , \A[567] , \A[568] , \A[569] , \A[570] , \A[571] , \A[572] ,
    \A[573] , \A[574] , \A[575] , \A[576] , \A[577] , \A[578] , \A[579] ,
    \A[580] , \A[581] , \A[582] , \A[583] , \A[584] , \A[585] , \A[586] ,
    \A[587] , \A[588] , \A[589] , \A[590] , \A[591] , \A[592] , \A[593] ,
    \A[594] , \A[595] , \A[596] , \A[597] , \A[598] , \A[599] , \A[600] ,
    \A[601] , \A[602] , \A[603] , \A[604] , \A[605] , \A[606] , \A[607] ,
    \A[608] , \A[609] , \A[610] , \A[611] , \A[612] , \A[613] , \A[614] ,
    \A[615] , \A[616] , \A[617] , \A[618] , \A[619] , \A[620] , \A[621] ,
    \A[622] , \A[623] , \A[624] , \A[625] , \A[626] , \A[627] , \A[628] ,
    \A[629] , \A[630] , \A[631] , \A[632] , \A[633] , \A[634] , \A[635] ,
    \A[636] , \A[637] , \A[638] , \A[639] , \A[640] , \A[641] , \A[642] ,
    \A[643] , \A[644] , \A[645] , \A[646] , \A[647] , \A[648] , \A[649] ,
    \A[650] , \A[651] , \A[652] , \A[653] , \A[654] , \A[655] , \A[656] ,
    \A[657] , \A[658] , \A[659] , \A[660] , \A[661] , \A[662] , \A[663] ,
    \A[664] , \A[665] , \A[666] , \A[667] , \A[668] , \A[669] , \A[670] ,
    \A[671] , \A[672] , \A[673] , \A[674] , \A[675] , \A[676] , \A[677] ,
    \A[678] , \A[679] , \A[680] , \A[681] , \A[682] , \A[683] , \A[684] ,
    \A[685] , \A[686] , \A[687] , \A[688] , \A[689] , \A[690] , \A[691] ,
    \A[692] , \A[693] , \A[694] , \A[695] , \A[696] , \A[697] , \A[698] ,
    \A[699] , \A[700] , \A[701] , \A[702] , \A[703] , \A[704] , \A[705] ,
    \A[706] , \A[707] , \A[708] , \A[709] , \A[710] , \A[711] , \A[712] ,
    \A[713] , \A[714] , \A[715] , \A[716] , \A[717] , \A[718] , \A[719] ,
    \A[720] , \A[721] , \A[722] , \A[723] , \A[724] , \A[725] , \A[726] ,
    \A[727] , \A[728] , \A[729] , \A[730] , \A[731] , \A[732] , \A[733] ,
    \A[734] , \A[735] , \A[736] , \A[737] , \A[738] , \A[739] , \A[740] ,
    \A[741] , \A[742] , \A[743] , \A[744] , \A[745] , \A[746] , \A[747] ,
    \A[748] , \A[749] , \A[750] , \A[751] , \A[752] , \A[753] , \A[754] ,
    \A[755] , \A[756] , \A[757] , \A[758] , \A[759] , \A[760] , \A[761] ,
    \A[762] , \A[763] , \A[764] , \A[765] , \A[766] , \A[767] , \A[768] ,
    \A[769] , \A[770] , \A[771] , \A[772] , \A[773] , \A[774] , \A[775] ,
    \A[776] , \A[777] , \A[778] , \A[779] , \A[780] , \A[781] , \A[782] ,
    \A[783] , \A[784] , \A[785] , \A[786] , \A[787] , \A[788] , \A[789] ,
    \A[790] , \A[791] , \A[792] , \A[793] , \A[794] , \A[795] , \A[796] ,
    \A[797] , \A[798] , \A[799] , \A[800] , \A[801] , \A[802] , \A[803] ,
    \A[804] , \A[805] , \A[806] , \A[807] , \A[808] , \A[809] , \A[810] ,
    \A[811] , \A[812] , \A[813] , \A[814] , \A[815] , \A[816] , \A[817] ,
    \A[818] , \A[819] , \A[820] , \A[821] , \A[822] , \A[823] , \A[824] ,
    \A[825] , \A[826] , \A[827] , \A[828] , \A[829] , \A[830] , \A[831] ,
    \A[832] , \A[833] , \A[834] , \A[835] , \A[836] , \A[837] , \A[838] ,
    \A[839] , \A[840] , \A[841] , \A[842] , \A[843] , \A[844] , \A[845] ,
    \A[846] , \A[847] , \A[848] , \A[849] , \A[850] , \A[851] , \A[852] ,
    \A[853] , \A[854] , \A[855] , \A[856] , \A[857] , \A[858] , \A[859] ,
    \A[860] , \A[861] , \A[862] , \A[863] , \A[864] , \A[865] , \A[866] ,
    \A[867] , \A[868] , \A[869] , \A[870] , \A[871] , \A[872] , \A[873] ,
    \A[874] , \A[875] , \A[876] , \A[877] , \A[878] , \A[879] , \A[880] ,
    \A[881] , \A[882] , \A[883] , \A[884] , \A[885] , \A[886] , \A[887] ,
    \A[888] , \A[889] , \A[890] , \A[891] , \A[892] , \A[893] , \A[894] ,
    \A[895] , \A[896] , \A[897] , \A[898] , \A[899] , \A[900] , \A[901] ,
    \A[902] , \A[903] , \A[904] , \A[905] , \A[906] , \A[907] , \A[908] ,
    \A[909] , \A[910] , \A[911] , \A[912] , \A[913] , \A[914] , \A[915] ,
    \A[916] , \A[917] , \A[918] , \A[919] , \A[920] , \A[921] , \A[922] ,
    \A[923] , \A[924] , \A[925] , \A[926] , \A[927] , \A[928] , \A[929] ,
    \A[930] , \A[931] , \A[932] , \A[933] , \A[934] , \A[935] , \A[936] ,
    \A[937] , \A[938] , \A[939] , \A[940] , \A[941] , \A[942] , \A[943] ,
    \A[944] , \A[945] , \A[946] , \A[947] , \A[948] , \A[949] , \A[950] ,
    \A[951] , \A[952] , \A[953] , \A[954] , \A[955] , \A[956] , \A[957] ,
    \A[958] , \A[959] , \A[960] , \A[961] , \A[962] , \A[963] , \A[964] ,
    \A[965] , \A[966] , \A[967] , \A[968] , \A[969] , \A[970] , \A[971] ,
    \A[972] , \A[973] , \A[974] , \A[975] , \A[976] , \A[977] , \A[978] ,
    \A[979] , \A[980] , \A[981] , \A[982] , \A[983] , \A[984] , \A[985] ,
    \A[986] , \A[987] , \A[988] , \A[989] , \A[990] , \A[991] , \A[992] ,
    \A[993] , \A[994] , \A[995] , \A[996] , \A[997] , \A[998] , \A[999] ,
    \A[1000] ,
    maj  );
  input  \A[0] , \A[1] , \A[2] , \A[3] , \A[4] , \A[5] , \A[6] , \A[7] ,
    \A[8] , \A[9] , \A[10] , \A[11] , \A[12] , \A[13] , \A[14] , \A[15] ,
    \A[16] , \A[17] , \A[18] , \A[19] , \A[20] , \A[21] , \A[22] , \A[23] ,
    \A[24] , \A[25] , \A[26] , \A[27] , \A[28] , \A[29] , \A[30] , \A[31] ,
    \A[32] , \A[33] , \A[34] , \A[35] , \A[36] , \A[37] , \A[38] , \A[39] ,
    \A[40] , \A[41] , \A[42] , \A[43] , \A[44] , \A[45] , \A[46] , \A[47] ,
    \A[48] , \A[49] , \A[50] , \A[51] , \A[52] , \A[53] , \A[54] , \A[55] ,
    \A[56] , \A[57] , \A[58] , \A[59] , \A[60] , \A[61] , \A[62] , \A[63] ,
    \A[64] , \A[65] , \A[66] , \A[67] , \A[68] , \A[69] , \A[70] , \A[71] ,
    \A[72] , \A[73] , \A[74] , \A[75] , \A[76] , \A[77] , \A[78] , \A[79] ,
    \A[80] , \A[81] , \A[82] , \A[83] , \A[84] , \A[85] , \A[86] , \A[87] ,
    \A[88] , \A[89] , \A[90] , \A[91] , \A[92] , \A[93] , \A[94] , \A[95] ,
    \A[96] , \A[97] , \A[98] , \A[99] , \A[100] , \A[101] , \A[102] ,
    \A[103] , \A[104] , \A[105] , \A[106] , \A[107] , \A[108] , \A[109] ,
    \A[110] , \A[111] , \A[112] , \A[113] , \A[114] , \A[115] , \A[116] ,
    \A[117] , \A[118] , \A[119] , \A[120] , \A[121] , \A[122] , \A[123] ,
    \A[124] , \A[125] , \A[126] , \A[127] , \A[128] , \A[129] , \A[130] ,
    \A[131] , \A[132] , \A[133] , \A[134] , \A[135] , \A[136] , \A[137] ,
    \A[138] , \A[139] , \A[140] , \A[141] , \A[142] , \A[143] , \A[144] ,
    \A[145] , \A[146] , \A[147] , \A[148] , \A[149] , \A[150] , \A[151] ,
    \A[152] , \A[153] , \A[154] , \A[155] , \A[156] , \A[157] , \A[158] ,
    \A[159] , \A[160] , \A[161] , \A[162] , \A[163] , \A[164] , \A[165] ,
    \A[166] , \A[167] , \A[168] , \A[169] , \A[170] , \A[171] , \A[172] ,
    \A[173] , \A[174] , \A[175] , \A[176] , \A[177] , \A[178] , \A[179] ,
    \A[180] , \A[181] , \A[182] , \A[183] , \A[184] , \A[185] , \A[186] ,
    \A[187] , \A[188] , \A[189] , \A[190] , \A[191] , \A[192] , \A[193] ,
    \A[194] , \A[195] , \A[196] , \A[197] , \A[198] , \A[199] , \A[200] ,
    \A[201] , \A[202] , \A[203] , \A[204] , \A[205] , \A[206] , \A[207] ,
    \A[208] , \A[209] , \A[210] , \A[211] , \A[212] , \A[213] , \A[214] ,
    \A[215] , \A[216] , \A[217] , \A[218] , \A[219] , \A[220] , \A[221] ,
    \A[222] , \A[223] , \A[224] , \A[225] , \A[226] , \A[227] , \A[228] ,
    \A[229] , \A[230] , \A[231] , \A[232] , \A[233] , \A[234] , \A[235] ,
    \A[236] , \A[237] , \A[238] , \A[239] , \A[240] , \A[241] , \A[242] ,
    \A[243] , \A[244] , \A[245] , \A[246] , \A[247] , \A[248] , \A[249] ,
    \A[250] , \A[251] , \A[252] , \A[253] , \A[254] , \A[255] , \A[256] ,
    \A[257] , \A[258] , \A[259] , \A[260] , \A[261] , \A[262] , \A[263] ,
    \A[264] , \A[265] , \A[266] , \A[267] , \A[268] , \A[269] , \A[270] ,
    \A[271] , \A[272] , \A[273] , \A[274] , \A[275] , \A[276] , \A[277] ,
    \A[278] , \A[279] , \A[280] , \A[281] , \A[282] , \A[283] , \A[284] ,
    \A[285] , \A[286] , \A[287] , \A[288] , \A[289] , \A[290] , \A[291] ,
    \A[292] , \A[293] , \A[294] , \A[295] , \A[296] , \A[297] , \A[298] ,
    \A[299] , \A[300] , \A[301] , \A[302] , \A[303] , \A[304] , \A[305] ,
    \A[306] , \A[307] , \A[308] , \A[309] , \A[310] , \A[311] , \A[312] ,
    \A[313] , \A[314] , \A[315] , \A[316] , \A[317] , \A[318] , \A[319] ,
    \A[320] , \A[321] , \A[322] , \A[323] , \A[324] , \A[325] , \A[326] ,
    \A[327] , \A[328] , \A[329] , \A[330] , \A[331] , \A[332] , \A[333] ,
    \A[334] , \A[335] , \A[336] , \A[337] , \A[338] , \A[339] , \A[340] ,
    \A[341] , \A[342] , \A[343] , \A[344] , \A[345] , \A[346] , \A[347] ,
    \A[348] , \A[349] , \A[350] , \A[351] , \A[352] , \A[353] , \A[354] ,
    \A[355] , \A[356] , \A[357] , \A[358] , \A[359] , \A[360] , \A[361] ,
    \A[362] , \A[363] , \A[364] , \A[365] , \A[366] , \A[367] , \A[368] ,
    \A[369] , \A[370] , \A[371] , \A[372] , \A[373] , \A[374] , \A[375] ,
    \A[376] , \A[377] , \A[378] , \A[379] , \A[380] , \A[381] , \A[382] ,
    \A[383] , \A[384] , \A[385] , \A[386] , \A[387] , \A[388] , \A[389] ,
    \A[390] , \A[391] , \A[392] , \A[393] , \A[394] , \A[395] , \A[396] ,
    \A[397] , \A[398] , \A[399] , \A[400] , \A[401] , \A[402] , \A[403] ,
    \A[404] , \A[405] , \A[406] , \A[407] , \A[408] , \A[409] , \A[410] ,
    \A[411] , \A[412] , \A[413] , \A[414] , \A[415] , \A[416] , \A[417] ,
    \A[418] , \A[419] , \A[420] , \A[421] , \A[422] , \A[423] , \A[424] ,
    \A[425] , \A[426] , \A[427] , \A[428] , \A[429] , \A[430] , \A[431] ,
    \A[432] , \A[433] , \A[434] , \A[435] , \A[436] , \A[437] , \A[438] ,
    \A[439] , \A[440] , \A[441] , \A[442] , \A[443] , \A[444] , \A[445] ,
    \A[446] , \A[447] , \A[448] , \A[449] , \A[450] , \A[451] , \A[452] ,
    \A[453] , \A[454] , \A[455] , \A[456] , \A[457] , \A[458] , \A[459] ,
    \A[460] , \A[461] , \A[462] , \A[463] , \A[464] , \A[465] , \A[466] ,
    \A[467] , \A[468] , \A[469] , \A[470] , \A[471] , \A[472] , \A[473] ,
    \A[474] , \A[475] , \A[476] , \A[477] , \A[478] , \A[479] , \A[480] ,
    \A[481] , \A[482] , \A[483] , \A[484] , \A[485] , \A[486] , \A[487] ,
    \A[488] , \A[489] , \A[490] , \A[491] , \A[492] , \A[493] , \A[494] ,
    \A[495] , \A[496] , \A[497] , \A[498] , \A[499] , \A[500] , \A[501] ,
    \A[502] , \A[503] , \A[504] , \A[505] , \A[506] , \A[507] , \A[508] ,
    \A[509] , \A[510] , \A[511] , \A[512] , \A[513] , \A[514] , \A[515] ,
    \A[516] , \A[517] , \A[518] , \A[519] , \A[520] , \A[521] , \A[522] ,
    \A[523] , \A[524] , \A[525] , \A[526] , \A[527] , \A[528] , \A[529] ,
    \A[530] , \A[531] , \A[532] , \A[533] , \A[534] , \A[535] , \A[536] ,
    \A[537] , \A[538] , \A[539] , \A[540] , \A[541] , \A[542] , \A[543] ,
    \A[544] , \A[545] , \A[546] , \A[547] , \A[548] , \A[549] , \A[550] ,
    \A[551] , \A[552] , \A[553] , \A[554] , \A[555] , \A[556] , \A[557] ,
    \A[558] , \A[559] , \A[560] , \A[561] , \A[562] , \A[563] , \A[564] ,
    \A[565] , \A[566] , \A[567] , \A[568] , \A[569] , \A[570] , \A[571] ,
    \A[572] , \A[573] , \A[574] , \A[575] , \A[576] , \A[577] , \A[578] ,
    \A[579] , \A[580] , \A[581] , \A[582] , \A[583] , \A[584] , \A[585] ,
    \A[586] , \A[587] , \A[588] , \A[589] , \A[590] , \A[591] , \A[592] ,
    \A[593] , \A[594] , \A[595] , \A[596] , \A[597] , \A[598] , \A[599] ,
    \A[600] , \A[601] , \A[602] , \A[603] , \A[604] , \A[605] , \A[606] ,
    \A[607] , \A[608] , \A[609] , \A[610] , \A[611] , \A[612] , \A[613] ,
    \A[614] , \A[615] , \A[616] , \A[617] , \A[618] , \A[619] , \A[620] ,
    \A[621] , \A[622] , \A[623] , \A[624] , \A[625] , \A[626] , \A[627] ,
    \A[628] , \A[629] , \A[630] , \A[631] , \A[632] , \A[633] , \A[634] ,
    \A[635] , \A[636] , \A[637] , \A[638] , \A[639] , \A[640] , \A[641] ,
    \A[642] , \A[643] , \A[644] , \A[645] , \A[646] , \A[647] , \A[648] ,
    \A[649] , \A[650] , \A[651] , \A[652] , \A[653] , \A[654] , \A[655] ,
    \A[656] , \A[657] , \A[658] , \A[659] , \A[660] , \A[661] , \A[662] ,
    \A[663] , \A[664] , \A[665] , \A[666] , \A[667] , \A[668] , \A[669] ,
    \A[670] , \A[671] , \A[672] , \A[673] , \A[674] , \A[675] , \A[676] ,
    \A[677] , \A[678] , \A[679] , \A[680] , \A[681] , \A[682] , \A[683] ,
    \A[684] , \A[685] , \A[686] , \A[687] , \A[688] , \A[689] , \A[690] ,
    \A[691] , \A[692] , \A[693] , \A[694] , \A[695] , \A[696] , \A[697] ,
    \A[698] , \A[699] , \A[700] , \A[701] , \A[702] , \A[703] , \A[704] ,
    \A[705] , \A[706] , \A[707] , \A[708] , \A[709] , \A[710] , \A[711] ,
    \A[712] , \A[713] , \A[714] , \A[715] , \A[716] , \A[717] , \A[718] ,
    \A[719] , \A[720] , \A[721] , \A[722] , \A[723] , \A[724] , \A[725] ,
    \A[726] , \A[727] , \A[728] , \A[729] , \A[730] , \A[731] , \A[732] ,
    \A[733] , \A[734] , \A[735] , \A[736] , \A[737] , \A[738] , \A[739] ,
    \A[740] , \A[741] , \A[742] , \A[743] , \A[744] , \A[745] , \A[746] ,
    \A[747] , \A[748] , \A[749] , \A[750] , \A[751] , \A[752] , \A[753] ,
    \A[754] , \A[755] , \A[756] , \A[757] , \A[758] , \A[759] , \A[760] ,
    \A[761] , \A[762] , \A[763] , \A[764] , \A[765] , \A[766] , \A[767] ,
    \A[768] , \A[769] , \A[770] , \A[771] , \A[772] , \A[773] , \A[774] ,
    \A[775] , \A[776] , \A[777] , \A[778] , \A[779] , \A[780] , \A[781] ,
    \A[782] , \A[783] , \A[784] , \A[785] , \A[786] , \A[787] , \A[788] ,
    \A[789] , \A[790] , \A[791] , \A[792] , \A[793] , \A[794] , \A[795] ,
    \A[796] , \A[797] , \A[798] , \A[799] , \A[800] , \A[801] , \A[802] ,
    \A[803] , \A[804] , \A[805] , \A[806] , \A[807] , \A[808] , \A[809] ,
    \A[810] , \A[811] , \A[812] , \A[813] , \A[814] , \A[815] , \A[816] ,
    \A[817] , \A[818] , \A[819] , \A[820] , \A[821] , \A[822] , \A[823] ,
    \A[824] , \A[825] , \A[826] , \A[827] , \A[828] , \A[829] , \A[830] ,
    \A[831] , \A[832] , \A[833] , \A[834] , \A[835] , \A[836] , \A[837] ,
    \A[838] , \A[839] , \A[840] , \A[841] , \A[842] , \A[843] , \A[844] ,
    \A[845] , \A[846] , \A[847] , \A[848] , \A[849] , \A[850] , \A[851] ,
    \A[852] , \A[853] , \A[854] , \A[855] , \A[856] , \A[857] , \A[858] ,
    \A[859] , \A[860] , \A[861] , \A[862] , \A[863] , \A[864] , \A[865] ,
    \A[866] , \A[867] , \A[868] , \A[869] , \A[870] , \A[871] , \A[872] ,
    \A[873] , \A[874] , \A[875] , \A[876] , \A[877] , \A[878] , \A[879] ,
    \A[880] , \A[881] , \A[882] , \A[883] , \A[884] , \A[885] , \A[886] ,
    \A[887] , \A[888] , \A[889] , \A[890] , \A[891] , \A[892] , \A[893] ,
    \A[894] , \A[895] , \A[896] , \A[897] , \A[898] , \A[899] , \A[900] ,
    \A[901] , \A[902] , \A[903] , \A[904] , \A[905] , \A[906] , \A[907] ,
    \A[908] , \A[909] , \A[910] , \A[911] , \A[912] , \A[913] , \A[914] ,
    \A[915] , \A[916] , \A[917] , \A[918] , \A[919] , \A[920] , \A[921] ,
    \A[922] , \A[923] , \A[924] , \A[925] , \A[926] , \A[927] , \A[928] ,
    \A[929] , \A[930] , \A[931] , \A[932] , \A[933] , \A[934] , \A[935] ,
    \A[936] , \A[937] , \A[938] , \A[939] , \A[940] , \A[941] , \A[942] ,
    \A[943] , \A[944] , \A[945] , \A[946] , \A[947] , \A[948] , \A[949] ,
    \A[950] , \A[951] , \A[952] , \A[953] , \A[954] , \A[955] , \A[956] ,
    \A[957] , \A[958] , \A[959] , \A[960] , \A[961] , \A[962] , \A[963] ,
    \A[964] , \A[965] , \A[966] , \A[967] , \A[968] , \A[969] , \A[970] ,
    \A[971] , \A[972] , \A[973] , \A[974] , \A[975] , \A[976] , \A[977] ,
    \A[978] , \A[979] , \A[980] , \A[981] , \A[982] , \A[983] , \A[984] ,
    \A[985] , \A[986] , \A[987] , \A[988] , \A[989] , \A[990] , \A[991] ,
    \A[992] , \A[993] , \A[994] , \A[995] , \A[996] , \A[997] , \A[998] ,
    \A[999] , \A[1000] ;
  output maj;
  wire new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_,
    new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_,
    new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_,
    new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_,
    new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_,
    new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_,
    new_n1038_, new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_,
    new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_,
    new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_,
    new_n1056_, new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_,
    new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_,
    new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1072_, new_n1073_,
    new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1078_, new_n1079_,
    new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1085_,
    new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_, new_n1091_,
    new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_,
    new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_,
    new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_,
    new_n1110_, new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1115_,
    new_n1116_, new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1121_,
    new_n1122_, new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_,
    new_n1128_, new_n1129_, new_n1130_, new_n1131_, new_n1132_, new_n1133_,
    new_n1134_, new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1139_,
    new_n1140_, new_n1141_, new_n1142_, new_n1143_, new_n1144_, new_n1145_,
    new_n1146_, new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_,
    new_n1152_, new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_,
    new_n1158_, new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_,
    new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_,
    new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_,
    new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_,
    new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1187_,
    new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1193_,
    new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1199_,
    new_n1200_, new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_,
    new_n1206_, new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_,
    new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_,
    new_n1218_, new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_,
    new_n1224_, new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_,
    new_n1230_, new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_,
    new_n1236_, new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_,
    new_n1242_, new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_,
    new_n1248_, new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_,
    new_n1254_, new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_,
    new_n1260_, new_n1261_, new_n1262_, new_n1263_, new_n1264_, new_n1265_,
    new_n1266_, new_n1267_, new_n1268_, new_n1269_, new_n1270_, new_n1271_,
    new_n1272_, new_n1273_, new_n1274_, new_n1275_, new_n1276_, new_n1277_,
    new_n1278_, new_n1279_, new_n1280_, new_n1281_, new_n1282_, new_n1283_,
    new_n1284_, new_n1285_, new_n1286_, new_n1287_, new_n1288_, new_n1289_,
    new_n1290_, new_n1291_, new_n1292_, new_n1293_, new_n1294_, new_n1295_,
    new_n1296_, new_n1297_, new_n1298_, new_n1299_, new_n1300_, new_n1301_,
    new_n1302_, new_n1303_, new_n1304_, new_n1305_, new_n1306_, new_n1307_,
    new_n1308_, new_n1309_, new_n1310_, new_n1311_, new_n1312_, new_n1313_,
    new_n1314_, new_n1315_, new_n1316_, new_n1317_, new_n1318_, new_n1319_,
    new_n1320_, new_n1321_, new_n1322_, new_n1323_, new_n1324_, new_n1325_,
    new_n1326_, new_n1327_, new_n1328_, new_n1329_, new_n1330_, new_n1331_,
    new_n1332_, new_n1333_, new_n1334_, new_n1335_, new_n1336_, new_n1337_,
    new_n1338_, new_n1339_, new_n1340_, new_n1341_, new_n1342_, new_n1343_,
    new_n1344_, new_n1345_, new_n1346_, new_n1347_, new_n1348_, new_n1349_,
    new_n1350_, new_n1351_, new_n1352_, new_n1353_, new_n1354_, new_n1355_,
    new_n1356_, new_n1357_, new_n1358_, new_n1359_, new_n1360_, new_n1361_,
    new_n1362_, new_n1363_, new_n1364_, new_n1365_, new_n1366_, new_n1367_,
    new_n1368_, new_n1369_, new_n1370_, new_n1371_, new_n1372_, new_n1373_,
    new_n1374_, new_n1375_, new_n1376_, new_n1377_, new_n1378_, new_n1379_,
    new_n1380_, new_n1381_, new_n1382_, new_n1383_, new_n1384_, new_n1385_,
    new_n1386_, new_n1387_, new_n1388_, new_n1389_, new_n1390_, new_n1391_,
    new_n1392_, new_n1393_, new_n1394_, new_n1395_, new_n1396_, new_n1397_,
    new_n1398_, new_n1399_, new_n1400_, new_n1401_, new_n1402_, new_n1403_,
    new_n1404_, new_n1405_, new_n1406_, new_n1407_, new_n1408_, new_n1409_,
    new_n1410_, new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_,
    new_n1416_, new_n1417_, new_n1418_, new_n1419_, new_n1420_, new_n1421_,
    new_n1422_, new_n1423_, new_n1424_, new_n1425_, new_n1426_, new_n1427_,
    new_n1428_, new_n1429_, new_n1430_, new_n1431_, new_n1432_, new_n1433_,
    new_n1434_, new_n1435_, new_n1436_, new_n1437_, new_n1438_, new_n1439_,
    new_n1440_, new_n1441_, new_n1442_, new_n1443_, new_n1444_, new_n1445_,
    new_n1446_, new_n1447_, new_n1448_, new_n1449_, new_n1450_, new_n1451_,
    new_n1452_, new_n1453_, new_n1454_, new_n1455_, new_n1456_, new_n1457_,
    new_n1458_, new_n1459_, new_n1460_, new_n1461_, new_n1462_, new_n1463_,
    new_n1464_, new_n1465_, new_n1466_, new_n1467_, new_n1468_, new_n1469_,
    new_n1470_, new_n1471_, new_n1472_, new_n1473_, new_n1474_, new_n1475_,
    new_n1476_, new_n1477_, new_n1478_, new_n1479_, new_n1480_, new_n1481_,
    new_n1482_, new_n1483_, new_n1484_, new_n1485_, new_n1486_, new_n1487_,
    new_n1488_, new_n1489_, new_n1490_, new_n1491_, new_n1492_, new_n1493_,
    new_n1494_, new_n1495_, new_n1496_, new_n1497_, new_n1498_, new_n1499_,
    new_n1500_, new_n1501_, new_n1502_, new_n1503_, new_n1504_, new_n1505_,
    new_n1506_, new_n1507_, new_n1508_, new_n1509_, new_n1510_, new_n1511_,
    new_n1512_, new_n1513_, new_n1514_, new_n1515_, new_n1516_, new_n1517_,
    new_n1518_, new_n1519_, new_n1520_, new_n1521_, new_n1522_, new_n1523_,
    new_n1524_, new_n1525_, new_n1526_, new_n1527_, new_n1528_, new_n1529_,
    new_n1530_, new_n1531_, new_n1532_, new_n1533_, new_n1534_, new_n1535_,
    new_n1536_, new_n1537_, new_n1538_, new_n1539_, new_n1540_, new_n1541_,
    new_n1542_, new_n1543_, new_n1544_, new_n1545_, new_n1546_, new_n1547_,
    new_n1548_, new_n1549_, new_n1550_, new_n1551_, new_n1552_, new_n1553_,
    new_n1554_, new_n1555_, new_n1556_, new_n1557_, new_n1558_, new_n1559_,
    new_n1560_, new_n1561_, new_n1562_, new_n1563_, new_n1564_, new_n1565_,
    new_n1566_, new_n1567_, new_n1568_, new_n1569_, new_n1570_, new_n1571_,
    new_n1572_, new_n1573_, new_n1574_, new_n1575_, new_n1576_, new_n1577_,
    new_n1578_, new_n1579_, new_n1580_, new_n1581_, new_n1582_, new_n1583_,
    new_n1584_, new_n1585_, new_n1586_, new_n1587_, new_n1588_, new_n1589_,
    new_n1590_, new_n1591_, new_n1592_, new_n1593_, new_n1594_, new_n1595_,
    new_n1596_, new_n1597_, new_n1598_, new_n1599_, new_n1600_, new_n1601_,
    new_n1602_, new_n1603_, new_n1604_, new_n1605_, new_n1606_, new_n1607_,
    new_n1608_, new_n1609_, new_n1610_, new_n1611_, new_n1612_, new_n1613_,
    new_n1614_, new_n1615_, new_n1616_, new_n1617_, new_n1618_, new_n1619_,
    new_n1620_, new_n1621_, new_n1622_, new_n1623_, new_n1624_, new_n1625_,
    new_n1626_, new_n1627_, new_n1628_, new_n1629_, new_n1630_, new_n1631_,
    new_n1632_, new_n1633_, new_n1634_, new_n1635_, new_n1636_, new_n1637_,
    new_n1638_, new_n1639_, new_n1640_, new_n1641_, new_n1642_, new_n1643_,
    new_n1644_, new_n1645_, new_n1646_, new_n1647_, new_n1648_, new_n1649_,
    new_n1650_, new_n1651_, new_n1652_, new_n1653_, new_n1654_, new_n1655_,
    new_n1656_, new_n1657_, new_n1658_, new_n1659_, new_n1660_, new_n1661_,
    new_n1662_, new_n1663_, new_n1664_, new_n1665_, new_n1666_, new_n1667_,
    new_n1668_, new_n1669_, new_n1670_, new_n1671_, new_n1672_, new_n1673_,
    new_n1674_, new_n1675_, new_n1676_, new_n1677_, new_n1678_, new_n1679_,
    new_n1680_, new_n1681_, new_n1682_, new_n1683_, new_n1684_, new_n1685_,
    new_n1686_, new_n1687_, new_n1688_, new_n1689_, new_n1690_, new_n1691_,
    new_n1692_, new_n1693_, new_n1694_, new_n1695_, new_n1696_, new_n1697_,
    new_n1698_, new_n1699_, new_n1700_, new_n1701_, new_n1702_, new_n1703_,
    new_n1704_, new_n1705_, new_n1706_, new_n1707_, new_n1708_, new_n1709_,
    new_n1710_, new_n1711_, new_n1712_, new_n1713_, new_n1714_, new_n1715_,
    new_n1716_, new_n1717_, new_n1718_, new_n1719_, new_n1720_, new_n1721_,
    new_n1722_, new_n1723_, new_n1724_, new_n1725_, new_n1726_, new_n1727_,
    new_n1728_, new_n1729_, new_n1730_, new_n1731_, new_n1732_, new_n1733_,
    new_n1734_, new_n1735_, new_n1736_, new_n1737_, new_n1738_, new_n1739_,
    new_n1740_, new_n1741_, new_n1742_, new_n1743_, new_n1744_, new_n1745_,
    new_n1746_, new_n1747_, new_n1748_, new_n1749_, new_n1750_, new_n1751_,
    new_n1752_, new_n1753_, new_n1754_, new_n1755_, new_n1756_, new_n1757_,
    new_n1758_, new_n1759_, new_n1760_, new_n1761_, new_n1762_, new_n1763_,
    new_n1764_, new_n1765_, new_n1766_, new_n1767_, new_n1768_, new_n1769_,
    new_n1770_, new_n1771_, new_n1772_, new_n1773_, new_n1774_, new_n1775_,
    new_n1776_, new_n1777_, new_n1778_, new_n1779_, new_n1780_, new_n1781_,
    new_n1782_, new_n1783_, new_n1784_, new_n1785_, new_n1786_, new_n1787_,
    new_n1788_, new_n1789_, new_n1790_, new_n1791_, new_n1792_, new_n1793_,
    new_n1794_, new_n1795_, new_n1796_, new_n1797_, new_n1798_, new_n1799_,
    new_n1800_, new_n1801_, new_n1802_, new_n1803_, new_n1804_, new_n1805_,
    new_n1806_, new_n1807_, new_n1808_, new_n1809_, new_n1810_, new_n1811_,
    new_n1812_, new_n1813_, new_n1814_, new_n1815_, new_n1816_, new_n1817_,
    new_n1818_, new_n1819_, new_n1820_, new_n1821_, new_n1822_, new_n1823_,
    new_n1824_, new_n1825_, new_n1826_, new_n1827_, new_n1828_, new_n1829_,
    new_n1830_, new_n1831_, new_n1832_, new_n1833_, new_n1834_, new_n1835_,
    new_n1836_, new_n1837_, new_n1838_, new_n1839_, new_n1840_, new_n1841_,
    new_n1842_, new_n1843_, new_n1844_, new_n1845_, new_n1846_, new_n1847_,
    new_n1848_, new_n1849_, new_n1850_, new_n1851_, new_n1852_, new_n1853_,
    new_n1854_, new_n1855_, new_n1856_, new_n1857_, new_n1858_, new_n1859_,
    new_n1860_, new_n1861_, new_n1862_, new_n1863_, new_n1864_, new_n1865_,
    new_n1866_, new_n1867_, new_n1868_, new_n1869_, new_n1870_, new_n1871_,
    new_n1872_, new_n1873_, new_n1874_, new_n1875_, new_n1876_, new_n1877_,
    new_n1878_, new_n1879_, new_n1880_, new_n1881_, new_n1882_, new_n1883_,
    new_n1884_, new_n1885_, new_n1886_, new_n1887_, new_n1888_, new_n1889_,
    new_n1890_, new_n1891_, new_n1892_, new_n1893_, new_n1894_, new_n1895_,
    new_n1896_, new_n1897_, new_n1898_, new_n1899_, new_n1900_, new_n1901_,
    new_n1902_, new_n1903_, new_n1904_, new_n1905_, new_n1906_, new_n1907_,
    new_n1908_, new_n1909_, new_n1910_, new_n1911_, new_n1912_, new_n1913_,
    new_n1914_, new_n1915_, new_n1916_, new_n1917_, new_n1918_, new_n1919_,
    new_n1920_, new_n1921_, new_n1922_, new_n1923_, new_n1924_, new_n1925_,
    new_n1926_, new_n1927_, new_n1928_, new_n1929_, new_n1930_, new_n1931_,
    new_n1932_, new_n1933_, new_n1934_, new_n1935_, new_n1936_, new_n1937_,
    new_n1938_, new_n1939_, new_n1940_, new_n1941_, new_n1942_, new_n1943_,
    new_n1944_, new_n1945_, new_n1946_, new_n1947_, new_n1948_, new_n1949_,
    new_n1950_, new_n1951_, new_n1952_, new_n1953_, new_n1954_, new_n1955_,
    new_n1956_, new_n1957_, new_n1958_, new_n1959_, new_n1960_, new_n1961_,
    new_n1962_, new_n1963_, new_n1964_, new_n1965_, new_n1966_, new_n1967_,
    new_n1968_, new_n1969_, new_n1970_, new_n1971_, new_n1972_, new_n1973_,
    new_n1974_, new_n1975_, new_n1976_, new_n1977_, new_n1978_, new_n1979_,
    new_n1980_, new_n1981_, new_n1982_, new_n1983_, new_n1984_, new_n1985_,
    new_n1986_, new_n1987_, new_n1988_, new_n1989_, new_n1990_, new_n1991_,
    new_n1992_, new_n1993_, new_n1994_, new_n1995_, new_n1996_, new_n1997_,
    new_n1998_, new_n1999_, new_n2000_, new_n2001_, new_n2002_, new_n2003_,
    new_n2004_, new_n2005_, new_n2006_, new_n2007_, new_n2008_, new_n2009_,
    new_n2010_, new_n2011_, new_n2012_, new_n2013_, new_n2014_, new_n2015_,
    new_n2016_, new_n2017_, new_n2018_, new_n2019_, new_n2020_, new_n2021_,
    new_n2022_, new_n2023_, new_n2024_, new_n2025_, new_n2026_, new_n2027_,
    new_n2028_, new_n2029_, new_n2030_, new_n2031_, new_n2032_, new_n2033_,
    new_n2034_, new_n2035_, new_n2036_, new_n2037_, new_n2038_, new_n2039_,
    new_n2040_, new_n2041_, new_n2042_, new_n2043_, new_n2044_, new_n2045_,
    new_n2046_, new_n2047_, new_n2048_, new_n2049_, new_n2050_, new_n2051_,
    new_n2052_, new_n2053_, new_n2054_, new_n2055_, new_n2056_, new_n2057_,
    new_n2058_, new_n2059_, new_n2060_, new_n2061_, new_n2062_, new_n2063_,
    new_n2064_, new_n2065_, new_n2066_, new_n2067_, new_n2068_, new_n2069_,
    new_n2070_, new_n2071_, new_n2072_, new_n2073_, new_n2074_, new_n2075_,
    new_n2076_, new_n2077_, new_n2078_, new_n2079_, new_n2080_, new_n2081_,
    new_n2082_, new_n2083_, new_n2084_, new_n2085_, new_n2086_, new_n2087_,
    new_n2088_, new_n2089_, new_n2090_, new_n2091_, new_n2092_, new_n2093_,
    new_n2094_, new_n2095_, new_n2096_, new_n2097_, new_n2098_, new_n2099_,
    new_n2100_, new_n2101_, new_n2102_, new_n2103_, new_n2104_, new_n2105_,
    new_n2106_, new_n2107_, new_n2108_, new_n2109_, new_n2110_, new_n2111_,
    new_n2112_, new_n2113_, new_n2114_, new_n2115_, new_n2116_, new_n2117_,
    new_n2118_, new_n2119_, new_n2120_, new_n2121_, new_n2122_, new_n2123_,
    new_n2124_, new_n2125_, new_n2126_, new_n2127_, new_n2128_, new_n2129_,
    new_n2130_, new_n2131_, new_n2132_, new_n2133_, new_n2134_, new_n2135_,
    new_n2136_, new_n2137_, new_n2138_, new_n2139_, new_n2140_, new_n2141_,
    new_n2142_, new_n2143_, new_n2144_, new_n2145_, new_n2146_, new_n2147_,
    new_n2148_, new_n2149_, new_n2150_, new_n2151_, new_n2152_, new_n2153_,
    new_n2154_, new_n2155_, new_n2156_, new_n2157_, new_n2158_, new_n2159_,
    new_n2160_, new_n2161_, new_n2162_, new_n2163_, new_n2164_, new_n2165_,
    new_n2166_, new_n2167_, new_n2168_, new_n2169_, new_n2170_, new_n2171_,
    new_n2172_, new_n2173_, new_n2174_, new_n2175_, new_n2176_, new_n2177_,
    new_n2178_, new_n2179_, new_n2180_, new_n2181_, new_n2182_, new_n2183_,
    new_n2184_, new_n2185_, new_n2186_, new_n2187_, new_n2188_, new_n2189_,
    new_n2190_, new_n2191_, new_n2192_, new_n2193_, new_n2194_, new_n2195_,
    new_n2196_, new_n2197_, new_n2198_, new_n2199_, new_n2200_, new_n2201_,
    new_n2202_, new_n2203_, new_n2204_, new_n2205_, new_n2206_, new_n2207_,
    new_n2208_, new_n2209_, new_n2210_, new_n2211_, new_n2212_, new_n2213_,
    new_n2214_, new_n2215_, new_n2216_, new_n2217_, new_n2218_, new_n2219_,
    new_n2220_, new_n2221_, new_n2222_, new_n2223_, new_n2224_, new_n2225_,
    new_n2226_, new_n2227_, new_n2228_, new_n2229_, new_n2230_, new_n2231_,
    new_n2232_, new_n2233_, new_n2234_, new_n2235_, new_n2236_, new_n2237_,
    new_n2238_, new_n2239_, new_n2240_, new_n2241_, new_n2242_, new_n2243_,
    new_n2244_, new_n2245_, new_n2246_, new_n2247_, new_n2248_, new_n2249_,
    new_n2250_, new_n2251_, new_n2252_, new_n2253_, new_n2254_, new_n2255_,
    new_n2256_, new_n2257_, new_n2258_, new_n2259_, new_n2260_, new_n2261_,
    new_n2262_, new_n2263_, new_n2264_, new_n2265_, new_n2266_, new_n2267_,
    new_n2268_, new_n2269_, new_n2270_, new_n2271_, new_n2272_, new_n2273_,
    new_n2274_, new_n2275_, new_n2276_, new_n2277_, new_n2278_, new_n2279_,
    new_n2280_, new_n2281_, new_n2282_, new_n2283_, new_n2284_, new_n2285_,
    new_n2286_, new_n2287_, new_n2288_, new_n2289_, new_n2290_, new_n2291_,
    new_n2292_, new_n2293_, new_n2294_, new_n2295_, new_n2296_, new_n2297_,
    new_n2298_, new_n2299_, new_n2300_, new_n2301_, new_n2302_, new_n2303_,
    new_n2304_, new_n2305_, new_n2306_, new_n2307_, new_n2308_, new_n2309_,
    new_n2310_, new_n2311_, new_n2312_, new_n2313_, new_n2314_, new_n2315_,
    new_n2316_, new_n2317_, new_n2318_, new_n2319_, new_n2320_, new_n2321_,
    new_n2322_, new_n2323_, new_n2324_, new_n2325_, new_n2326_, new_n2327_,
    new_n2328_, new_n2329_, new_n2330_, new_n2331_, new_n2332_, new_n2333_,
    new_n2334_, new_n2335_, new_n2336_, new_n2337_, new_n2338_, new_n2339_,
    new_n2340_, new_n2341_, new_n2342_, new_n2343_, new_n2344_, new_n2345_,
    new_n2346_, new_n2347_, new_n2348_, new_n2349_, new_n2350_, new_n2351_,
    new_n2352_, new_n2353_, new_n2354_, new_n2355_, new_n2356_, new_n2357_,
    new_n2358_, new_n2359_, new_n2360_, new_n2361_, new_n2362_, new_n2363_,
    new_n2364_, new_n2365_, new_n2366_, new_n2367_, new_n2368_, new_n2369_,
    new_n2370_, new_n2371_, new_n2372_, new_n2373_, new_n2374_, new_n2375_,
    new_n2376_, new_n2377_, new_n2378_, new_n2379_, new_n2380_, new_n2381_,
    new_n2382_, new_n2383_, new_n2384_, new_n2385_, new_n2386_, new_n2387_,
    new_n2388_, new_n2389_, new_n2390_, new_n2391_, new_n2392_, new_n2393_,
    new_n2394_, new_n2395_, new_n2396_, new_n2397_, new_n2398_, new_n2399_,
    new_n2400_, new_n2401_, new_n2402_, new_n2403_, new_n2404_, new_n2405_,
    new_n2406_, new_n2407_, new_n2408_, new_n2409_, new_n2410_, new_n2411_,
    new_n2412_, new_n2413_, new_n2414_, new_n2415_, new_n2416_, new_n2417_,
    new_n2418_, new_n2419_, new_n2420_, new_n2421_, new_n2422_, new_n2423_,
    new_n2424_, new_n2425_, new_n2426_, new_n2427_, new_n2428_, new_n2429_,
    new_n2430_, new_n2431_, new_n2432_, new_n2433_, new_n2434_, new_n2435_,
    new_n2436_, new_n2437_, new_n2438_, new_n2439_, new_n2440_, new_n2441_,
    new_n2442_, new_n2443_, new_n2444_, new_n2445_, new_n2446_, new_n2447_,
    new_n2448_, new_n2449_, new_n2450_, new_n2451_, new_n2452_, new_n2453_,
    new_n2454_, new_n2455_, new_n2456_, new_n2457_, new_n2458_, new_n2459_,
    new_n2460_, new_n2461_, new_n2462_, new_n2463_, new_n2464_, new_n2465_,
    new_n2466_, new_n2467_, new_n2468_, new_n2469_, new_n2470_, new_n2471_,
    new_n2472_, new_n2473_, new_n2474_, new_n2475_, new_n2476_, new_n2477_,
    new_n2478_, new_n2479_, new_n2480_, new_n2481_, new_n2482_, new_n2483_,
    new_n2484_, new_n2485_, new_n2486_, new_n2487_, new_n2488_, new_n2489_,
    new_n2490_, new_n2491_, new_n2492_, new_n2493_, new_n2494_, new_n2495_,
    new_n2496_, new_n2497_, new_n2498_, new_n2499_, new_n2500_, new_n2501_,
    new_n2502_, new_n2503_, new_n2504_, new_n2505_, new_n2506_, new_n2507_,
    new_n2508_, new_n2509_, new_n2510_, new_n2511_, new_n2512_, new_n2513_,
    new_n2514_, new_n2515_, new_n2516_, new_n2517_, new_n2518_, new_n2519_,
    new_n2520_, new_n2521_, new_n2522_, new_n2523_, new_n2524_, new_n2525_,
    new_n2526_, new_n2527_, new_n2528_, new_n2529_, new_n2530_, new_n2531_,
    new_n2532_, new_n2533_, new_n2534_, new_n2535_, new_n2536_, new_n2537_,
    new_n2538_, new_n2539_, new_n2540_, new_n2541_, new_n2542_, new_n2543_,
    new_n2544_, new_n2545_, new_n2546_, new_n2547_, new_n2548_, new_n2549_,
    new_n2550_, new_n2551_, new_n2552_, new_n2553_, new_n2554_, new_n2555_,
    new_n2556_, new_n2557_, new_n2558_, new_n2559_, new_n2560_, new_n2561_,
    new_n2562_, new_n2563_, new_n2564_, new_n2565_, new_n2566_, new_n2567_,
    new_n2568_, new_n2569_, new_n2570_, new_n2571_, new_n2572_, new_n2573_,
    new_n2574_, new_n2575_, new_n2576_, new_n2577_, new_n2578_, new_n2579_,
    new_n2580_, new_n2581_, new_n2582_, new_n2583_, new_n2584_, new_n2585_,
    new_n2586_, new_n2587_, new_n2588_, new_n2589_, new_n2590_, new_n2591_,
    new_n2592_, new_n2593_, new_n2594_, new_n2595_, new_n2596_, new_n2597_,
    new_n2598_, new_n2599_, new_n2600_, new_n2601_, new_n2602_, new_n2603_,
    new_n2604_, new_n2605_, new_n2606_, new_n2607_, new_n2608_, new_n2609_,
    new_n2610_, new_n2611_, new_n2612_, new_n2613_, new_n2614_, new_n2615_,
    new_n2616_, new_n2617_, new_n2618_, new_n2619_, new_n2620_, new_n2621_,
    new_n2622_, new_n2623_, new_n2624_, new_n2625_, new_n2626_, new_n2627_,
    new_n2628_, new_n2629_, new_n2630_, new_n2631_, new_n2632_, new_n2633_,
    new_n2634_, new_n2635_, new_n2636_, new_n2637_, new_n2638_, new_n2639_,
    new_n2640_, new_n2641_, new_n2642_, new_n2643_, new_n2644_, new_n2645_,
    new_n2646_, new_n2647_, new_n2648_, new_n2649_, new_n2650_, new_n2651_,
    new_n2652_, new_n2653_, new_n2654_, new_n2655_, new_n2656_, new_n2657_,
    new_n2658_, new_n2659_, new_n2660_, new_n2661_, new_n2662_, new_n2663_,
    new_n2664_, new_n2665_, new_n2666_, new_n2667_, new_n2668_, new_n2669_,
    new_n2670_, new_n2671_, new_n2672_, new_n2673_, new_n2674_, new_n2675_,
    new_n2676_, new_n2677_, new_n2678_, new_n2679_, new_n2680_, new_n2681_,
    new_n2682_, new_n2683_, new_n2684_, new_n2685_, new_n2686_, new_n2687_,
    new_n2688_, new_n2689_, new_n2690_, new_n2691_, new_n2692_, new_n2693_,
    new_n2694_, new_n2695_, new_n2696_, new_n2697_, new_n2698_, new_n2699_,
    new_n2700_, new_n2701_, new_n2702_, new_n2703_, new_n2704_, new_n2705_,
    new_n2706_, new_n2707_, new_n2708_, new_n2709_, new_n2710_, new_n2711_,
    new_n2712_, new_n2713_, new_n2714_, new_n2715_, new_n2716_, new_n2717_,
    new_n2718_, new_n2719_, new_n2720_, new_n2721_, new_n2722_, new_n2723_,
    new_n2724_, new_n2725_, new_n2726_, new_n2727_, new_n2728_, new_n2729_,
    new_n2730_, new_n2731_, new_n2732_, new_n2733_, new_n2734_, new_n2735_,
    new_n2736_, new_n2737_, new_n2738_, new_n2739_, new_n2740_, new_n2741_,
    new_n2742_, new_n2743_, new_n2744_, new_n2745_, new_n2746_, new_n2747_,
    new_n2748_, new_n2749_, new_n2750_, new_n2751_, new_n2752_, new_n2753_,
    new_n2754_, new_n2755_, new_n2756_, new_n2757_, new_n2758_, new_n2759_,
    new_n2760_, new_n2761_, new_n2762_, new_n2763_, new_n2764_, new_n2765_,
    new_n2766_, new_n2767_, new_n2768_, new_n2769_, new_n2770_, new_n2771_,
    new_n2772_, new_n2773_, new_n2774_, new_n2775_, new_n2776_, new_n2777_,
    new_n2778_, new_n2779_, new_n2780_, new_n2781_, new_n2782_, new_n2783_,
    new_n2784_, new_n2785_, new_n2786_, new_n2787_, new_n2788_, new_n2789_,
    new_n2790_, new_n2791_, new_n2792_, new_n2793_, new_n2794_, new_n2795_,
    new_n2796_, new_n2797_, new_n2798_, new_n2799_, new_n2800_, new_n2801_,
    new_n2802_, new_n2803_, new_n2804_, new_n2805_, new_n2806_, new_n2807_,
    new_n2808_, new_n2809_, new_n2810_, new_n2811_, new_n2812_, new_n2813_,
    new_n2814_, new_n2815_, new_n2816_, new_n2817_, new_n2818_, new_n2819_,
    new_n2820_, new_n2821_, new_n2822_, new_n2823_, new_n2824_, new_n2825_,
    new_n2826_, new_n2827_, new_n2828_, new_n2829_, new_n2830_, new_n2831_,
    new_n2832_, new_n2833_, new_n2834_, new_n2835_, new_n2836_, new_n2837_,
    new_n2838_, new_n2839_, new_n2840_, new_n2841_, new_n2842_, new_n2843_,
    new_n2844_, new_n2845_, new_n2846_, new_n2847_, new_n2848_, new_n2849_,
    new_n2850_, new_n2851_, new_n2852_, new_n2853_, new_n2854_, new_n2855_,
    new_n2856_, new_n2857_, new_n2858_, new_n2859_, new_n2860_, new_n2861_,
    new_n2862_, new_n2863_, new_n2864_, new_n2865_, new_n2866_, new_n2867_,
    new_n2868_, new_n2869_, new_n2870_, new_n2871_, new_n2872_, new_n2873_,
    new_n2874_, new_n2875_, new_n2876_, new_n2877_, new_n2878_, new_n2879_,
    new_n2880_, new_n2881_, new_n2882_, new_n2883_, new_n2884_, new_n2885_,
    new_n2886_, new_n2887_, new_n2888_, new_n2889_, new_n2890_, new_n2891_,
    new_n2892_, new_n2893_, new_n2894_, new_n2895_, new_n2896_, new_n2897_,
    new_n2898_, new_n2899_, new_n2900_, new_n2901_, new_n2902_, new_n2903_,
    new_n2904_, new_n2905_, new_n2906_, new_n2907_, new_n2908_, new_n2909_,
    new_n2910_, new_n2911_, new_n2912_, new_n2913_, new_n2914_, new_n2915_,
    new_n2916_, new_n2917_, new_n2918_, new_n2919_, new_n2920_, new_n2921_,
    new_n2922_, new_n2923_, new_n2924_, new_n2925_, new_n2926_, new_n2927_,
    new_n2928_, new_n2929_, new_n2930_, new_n2931_, new_n2932_, new_n2933_,
    new_n2934_, new_n2935_, new_n2936_, new_n2937_, new_n2938_, new_n2939_,
    new_n2940_, new_n2941_, new_n2942_, new_n2943_, new_n2944_, new_n2945_,
    new_n2946_, new_n2947_, new_n2948_, new_n2949_, new_n2950_, new_n2951_,
    new_n2952_, new_n2953_, new_n2954_, new_n2955_, new_n2956_, new_n2957_,
    new_n2958_, new_n2959_, new_n2960_, new_n2961_, new_n2962_, new_n2963_,
    new_n2964_, new_n2965_, new_n2966_, new_n2967_, new_n2968_, new_n2969_,
    new_n2970_, new_n2971_, new_n2972_, new_n2973_, new_n2974_, new_n2975_,
    new_n2976_, new_n2977_, new_n2978_, new_n2979_, new_n2980_, new_n2981_,
    new_n2982_, new_n2983_, new_n2984_, new_n2985_, new_n2986_, new_n2987_,
    new_n2988_, new_n2989_, new_n2990_, new_n2991_, new_n2992_, new_n2993_,
    new_n2994_, new_n2995_, new_n2996_, new_n2997_, new_n2998_, new_n2999_,
    new_n3000_, new_n3001_, new_n3002_, new_n3003_, new_n3004_, new_n3005_,
    new_n3006_, new_n3007_, new_n3008_, new_n3009_, new_n3010_, new_n3011_,
    new_n3012_, new_n3013_, new_n3014_, new_n3015_, new_n3016_, new_n3017_,
    new_n3018_, new_n3019_, new_n3020_, new_n3021_, new_n3022_, new_n3023_,
    new_n3024_, new_n3025_, new_n3026_, new_n3027_, new_n3028_, new_n3029_,
    new_n3030_, new_n3031_, new_n3032_, new_n3033_, new_n3034_, new_n3035_,
    new_n3036_, new_n3037_, new_n3038_, new_n3039_, new_n3040_, new_n3041_,
    new_n3042_, new_n3043_, new_n3044_, new_n3045_, new_n3046_, new_n3047_,
    new_n3048_, new_n3049_, new_n3050_, new_n3051_, new_n3052_, new_n3053_,
    new_n3054_, new_n3055_, new_n3056_, new_n3057_, new_n3058_, new_n3059_,
    new_n3060_, new_n3061_, new_n3062_, new_n3063_, new_n3064_, new_n3065_,
    new_n3066_, new_n3067_, new_n3068_, new_n3069_, new_n3070_, new_n3071_,
    new_n3072_, new_n3073_, new_n3074_, new_n3075_, new_n3076_, new_n3077_,
    new_n3078_, new_n3079_, new_n3080_, new_n3081_, new_n3082_, new_n3083_,
    new_n3084_, new_n3085_, new_n3086_, new_n3087_, new_n3088_, new_n3089_,
    new_n3090_, new_n3091_, new_n3092_, new_n3093_, new_n3094_, new_n3095_,
    new_n3096_, new_n3097_, new_n3098_, new_n3099_, new_n3100_, new_n3101_,
    new_n3102_, new_n3103_, new_n3104_, new_n3105_, new_n3106_, new_n3107_,
    new_n3108_, new_n3109_, new_n3110_, new_n3111_, new_n3112_, new_n3113_,
    new_n3114_, new_n3115_, new_n3116_, new_n3117_, new_n3118_, new_n3119_,
    new_n3120_, new_n3121_, new_n3122_, new_n3123_, new_n3124_, new_n3125_,
    new_n3126_, new_n3127_, new_n3128_, new_n3129_, new_n3130_, new_n3131_,
    new_n3132_, new_n3133_, new_n3134_, new_n3135_, new_n3136_, new_n3137_,
    new_n3138_, new_n3139_, new_n3140_, new_n3141_, new_n3142_, new_n3143_,
    new_n3144_, new_n3145_, new_n3146_, new_n3147_, new_n3148_, new_n3149_,
    new_n3150_, new_n3151_, new_n3152_, new_n3153_, new_n3154_, new_n3155_,
    new_n3156_, new_n3157_, new_n3158_, new_n3159_, new_n3160_, new_n3161_,
    new_n3162_, new_n3163_, new_n3164_, new_n3165_, new_n3166_, new_n3167_,
    new_n3168_, new_n3169_, new_n3170_, new_n3171_, new_n3172_, new_n3173_,
    new_n3174_, new_n3175_, new_n3176_, new_n3177_, new_n3178_, new_n3179_,
    new_n3180_, new_n3181_, new_n3182_, new_n3183_, new_n3184_, new_n3185_,
    new_n3186_, new_n3187_, new_n3188_, new_n3189_, new_n3190_, new_n3191_,
    new_n3192_, new_n3193_, new_n3194_, new_n3195_, new_n3196_, new_n3197_,
    new_n3198_, new_n3199_, new_n3200_, new_n3201_, new_n3202_, new_n3203_,
    new_n3204_, new_n3205_, new_n3206_, new_n3207_, new_n3208_, new_n3209_,
    new_n3210_, new_n3211_, new_n3212_, new_n3213_, new_n3214_, new_n3215_,
    new_n3216_, new_n3217_, new_n3218_, new_n3219_, new_n3220_, new_n3221_,
    new_n3222_, new_n3223_, new_n3224_, new_n3225_, new_n3226_, new_n3227_,
    new_n3228_, new_n3229_, new_n3230_, new_n3231_, new_n3232_, new_n3233_,
    new_n3234_, new_n3235_, new_n3236_, new_n3237_, new_n3238_, new_n3239_,
    new_n3240_, new_n3241_, new_n3242_, new_n3243_, new_n3244_, new_n3245_,
    new_n3246_, new_n3247_, new_n3248_, new_n3249_, new_n3250_, new_n3251_,
    new_n3252_, new_n3253_, new_n3254_, new_n3255_, new_n3256_, new_n3257_,
    new_n3258_, new_n3259_, new_n3260_, new_n3261_, new_n3262_, new_n3263_,
    new_n3264_, new_n3265_, new_n3266_, new_n3267_, new_n3268_, new_n3269_,
    new_n3270_, new_n3271_, new_n3272_, new_n3273_, new_n3274_, new_n3275_,
    new_n3276_, new_n3277_, new_n3278_, new_n3279_, new_n3280_, new_n3281_,
    new_n3282_, new_n3283_, new_n3284_, new_n3285_, new_n3286_, new_n3287_,
    new_n3288_, new_n3289_, new_n3290_, new_n3291_, new_n3292_, new_n3293_,
    new_n3294_, new_n3295_, new_n3296_, new_n3297_, new_n3298_, new_n3299_,
    new_n3300_, new_n3301_, new_n3302_, new_n3303_, new_n3304_, new_n3305_,
    new_n3306_, new_n3307_, new_n3308_, new_n3309_, new_n3310_, new_n3311_,
    new_n3312_, new_n3313_, new_n3314_, new_n3315_, new_n3316_, new_n3317_,
    new_n3318_, new_n3319_, new_n3320_, new_n3321_, new_n3322_, new_n3323_,
    new_n3324_, new_n3325_, new_n3326_, new_n3327_, new_n3328_, new_n3329_,
    new_n3330_, new_n3331_, new_n3332_, new_n3333_, new_n3334_, new_n3335_,
    new_n3336_, new_n3337_, new_n3338_, new_n3339_, new_n3340_, new_n3341_,
    new_n3342_, new_n3343_, new_n3344_, new_n3345_, new_n3346_, new_n3347_,
    new_n3348_, new_n3349_, new_n3350_, new_n3351_, new_n3352_, new_n3353_,
    new_n3354_, new_n3355_, new_n3356_, new_n3357_, new_n3358_, new_n3359_,
    new_n3360_, new_n3361_, new_n3362_, new_n3363_, new_n3364_, new_n3365_,
    new_n3366_, new_n3367_, new_n3368_, new_n3369_, new_n3370_, new_n3371_,
    new_n3372_, new_n3373_, new_n3374_, new_n3375_, new_n3376_, new_n3377_,
    new_n3378_, new_n3379_, new_n3380_, new_n3381_, new_n3382_, new_n3383_,
    new_n3384_, new_n3385_, new_n3386_, new_n3387_, new_n3388_, new_n3389_,
    new_n3390_, new_n3391_, new_n3392_, new_n3393_, new_n3394_, new_n3395_,
    new_n3396_, new_n3397_, new_n3398_, new_n3399_, new_n3400_, new_n3401_,
    new_n3402_, new_n3403_, new_n3404_, new_n3405_, new_n3406_, new_n3407_,
    new_n3408_, new_n3409_, new_n3410_, new_n3411_, new_n3412_, new_n3413_,
    new_n3414_, new_n3415_, new_n3416_, new_n3417_, new_n3418_, new_n3419_,
    new_n3420_, new_n3421_, new_n3422_, new_n3423_, new_n3424_, new_n3425_,
    new_n3426_, new_n3427_, new_n3428_, new_n3429_, new_n3430_, new_n3431_,
    new_n3432_, new_n3433_, new_n3434_, new_n3435_, new_n3436_, new_n3437_,
    new_n3438_, new_n3439_, new_n3440_, new_n3441_, new_n3442_, new_n3443_,
    new_n3444_, new_n3445_, new_n3446_, new_n3447_, new_n3448_, new_n3449_,
    new_n3450_, new_n3451_, new_n3452_, new_n3453_, new_n3454_, new_n3455_,
    new_n3456_, new_n3457_, new_n3458_, new_n3459_, new_n3460_, new_n3461_,
    new_n3462_, new_n3463_, new_n3464_, new_n3465_, new_n3466_, new_n3467_,
    new_n3468_, new_n3469_, new_n3470_, new_n3471_, new_n3472_, new_n3473_,
    new_n3474_, new_n3475_, new_n3476_, new_n3477_, new_n3478_, new_n3479_,
    new_n3480_, new_n3481_, new_n3482_, new_n3483_, new_n3484_, new_n3485_,
    new_n3486_, new_n3487_, new_n3488_, new_n3489_, new_n3490_, new_n3491_,
    new_n3492_, new_n3493_, new_n3494_, new_n3495_, new_n3496_, new_n3497_,
    new_n3498_, new_n3499_, new_n3500_, new_n3501_, new_n3502_, new_n3503_,
    new_n3504_, new_n3505_, new_n3506_, new_n3507_, new_n3508_, new_n3509_,
    new_n3510_, new_n3511_, new_n3512_, new_n3513_, new_n3514_, new_n3515_,
    new_n3516_, new_n3517_, new_n3518_, new_n3519_, new_n3520_, new_n3521_,
    new_n3522_, new_n3523_, new_n3524_, new_n3525_, new_n3526_, new_n3527_,
    new_n3528_, new_n3529_, new_n3530_, new_n3531_, new_n3532_, new_n3533_,
    new_n3534_, new_n3535_, new_n3536_, new_n3537_, new_n3538_, new_n3539_,
    new_n3540_, new_n3541_, new_n3542_, new_n3543_, new_n3544_, new_n3545_,
    new_n3546_, new_n3547_, new_n3548_, new_n3549_, new_n3550_, new_n3551_,
    new_n3552_, new_n3553_, new_n3554_, new_n3555_, new_n3556_, new_n3557_,
    new_n3558_, new_n3559_, new_n3560_, new_n3561_, new_n3562_, new_n3563_,
    new_n3564_, new_n3565_, new_n3566_, new_n3567_, new_n3568_, new_n3569_,
    new_n3570_, new_n3571_, new_n3572_, new_n3573_, new_n3574_, new_n3575_,
    new_n3576_, new_n3577_, new_n3578_, new_n3579_, new_n3580_, new_n3581_,
    new_n3582_, new_n3583_, new_n3584_, new_n3585_, new_n3586_, new_n3587_,
    new_n3588_, new_n3589_, new_n3590_, new_n3591_, new_n3592_, new_n3593_,
    new_n3594_, new_n3595_, new_n3596_, new_n3597_, new_n3598_, new_n3599_,
    new_n3600_, new_n3601_, new_n3602_, new_n3603_, new_n3604_, new_n3605_,
    new_n3606_, new_n3607_, new_n3608_, new_n3609_, new_n3610_, new_n3611_,
    new_n3612_, new_n3613_, new_n3614_, new_n3615_, new_n3616_, new_n3617_,
    new_n3618_, new_n3619_, new_n3620_, new_n3621_, new_n3622_, new_n3623_,
    new_n3624_, new_n3625_, new_n3626_, new_n3627_, new_n3628_, new_n3629_,
    new_n3630_, new_n3631_, new_n3632_, new_n3633_, new_n3634_, new_n3635_,
    new_n3636_, new_n3637_, new_n3638_, new_n3639_, new_n3640_, new_n3641_,
    new_n3642_, new_n3643_, new_n3644_, new_n3645_, new_n3646_, new_n3647_,
    new_n3648_, new_n3649_, new_n3650_, new_n3651_, new_n3652_, new_n3653_,
    new_n3654_, new_n3655_, new_n3656_, new_n3657_, new_n3658_, new_n3659_,
    new_n3660_, new_n3661_, new_n3662_, new_n3663_, new_n3664_, new_n3665_,
    new_n3666_, new_n3667_, new_n3668_, new_n3669_, new_n3670_, new_n3671_,
    new_n3672_, new_n3673_, new_n3674_, new_n3675_, new_n3676_, new_n3677_,
    new_n3678_, new_n3679_, new_n3680_, new_n3681_, new_n3682_, new_n3683_,
    new_n3684_, new_n3685_, new_n3686_, new_n3687_, new_n3688_, new_n3689_,
    new_n3690_, new_n3691_, new_n3692_, new_n3693_, new_n3694_, new_n3695_,
    new_n3696_, new_n3697_, new_n3698_, new_n3699_, new_n3700_, new_n3701_,
    new_n3702_, new_n3703_, new_n3704_, new_n3705_, new_n3706_, new_n3707_,
    new_n3708_, new_n3709_, new_n3710_, new_n3711_, new_n3712_, new_n3713_,
    new_n3714_, new_n3715_, new_n3716_, new_n3717_, new_n3718_, new_n3719_,
    new_n3720_, new_n3721_, new_n3722_, new_n3723_, new_n3724_, new_n3725_,
    new_n3726_, new_n3727_, new_n3728_, new_n3729_, new_n3730_, new_n3731_,
    new_n3732_, new_n3733_, new_n3734_, new_n3735_, new_n3736_, new_n3737_,
    new_n3738_, new_n3739_, new_n3740_, new_n3741_, new_n3742_, new_n3743_,
    new_n3744_, new_n3745_, new_n3746_, new_n3747_, new_n3748_, new_n3749_,
    new_n3750_, new_n3751_, new_n3752_, new_n3753_, new_n3754_, new_n3755_,
    new_n3756_, new_n3757_, new_n3758_, new_n3759_, new_n3760_, new_n3761_,
    new_n3762_, new_n3763_, new_n3764_, new_n3765_, new_n3766_, new_n3767_,
    new_n3768_, new_n3769_, new_n3770_, new_n3771_, new_n3772_, new_n3773_,
    new_n3774_, new_n3775_, new_n3776_, new_n3777_, new_n3778_, new_n3779_,
    new_n3780_, new_n3781_, new_n3782_, new_n3783_, new_n3784_, new_n3785_,
    new_n3786_, new_n3787_, new_n3788_, new_n3789_, new_n3790_, new_n3791_,
    new_n3792_, new_n3793_, new_n3794_, new_n3795_, new_n3796_, new_n3797_,
    new_n3798_, new_n3799_, new_n3800_, new_n3801_, new_n3802_, new_n3803_,
    new_n3804_, new_n3805_, new_n3806_, new_n3807_, new_n3808_, new_n3809_,
    new_n3810_, new_n3811_, new_n3812_, new_n3813_, new_n3814_, new_n3815_,
    new_n3816_, new_n3817_, new_n3818_, new_n3819_, new_n3820_, new_n3821_,
    new_n3822_, new_n3823_, new_n3824_, new_n3825_, new_n3826_, new_n3827_,
    new_n3828_, new_n3829_, new_n3830_, new_n3831_, new_n3832_, new_n3833_,
    new_n3834_, new_n3835_, new_n3836_, new_n3837_, new_n3838_, new_n3839_,
    new_n3840_, new_n3841_, new_n3842_, new_n3843_, new_n3844_, new_n3845_,
    new_n3846_, new_n3847_, new_n3848_, new_n3849_, new_n3850_, new_n3851_,
    new_n3852_, new_n3853_, new_n3854_, new_n3855_, new_n3856_, new_n3857_,
    new_n3858_, new_n3859_, new_n3860_, new_n3861_, new_n3862_, new_n3863_,
    new_n3864_, new_n3865_, new_n3866_, new_n3867_, new_n3868_, new_n3869_,
    new_n3870_, new_n3871_, new_n3872_, new_n3873_, new_n3874_, new_n3875_,
    new_n3876_, new_n3877_, new_n3878_, new_n3879_, new_n3880_, new_n3881_,
    new_n3882_, new_n3883_, new_n3884_, new_n3885_, new_n3886_, new_n3887_,
    new_n3888_, new_n3889_, new_n3890_, new_n3891_, new_n3892_, new_n3893_,
    new_n3894_, new_n3895_, new_n3896_, new_n3897_, new_n3898_, new_n3899_,
    new_n3900_, new_n3901_, new_n3902_, new_n3903_, new_n3904_, new_n3905_,
    new_n3906_, new_n3907_, new_n3908_, new_n3909_, new_n3910_, new_n3911_,
    new_n3912_, new_n3913_, new_n3914_, new_n3915_, new_n3916_, new_n3917_,
    new_n3918_, new_n3919_, new_n3920_, new_n3921_, new_n3922_, new_n3923_,
    new_n3924_, new_n3925_, new_n3926_, new_n3927_, new_n3928_, new_n3929_,
    new_n3930_, new_n3931_, new_n3932_, new_n3933_, new_n3934_, new_n3935_,
    new_n3936_, new_n3937_, new_n3938_, new_n3939_, new_n3940_, new_n3941_,
    new_n3942_, new_n3943_, new_n3944_, new_n3945_, new_n3946_, new_n3947_,
    new_n3948_, new_n3949_, new_n3950_, new_n3951_, new_n3952_, new_n3953_,
    new_n3954_, new_n3955_, new_n3956_, new_n3957_, new_n3958_, new_n3959_,
    new_n3960_, new_n3961_, new_n3962_, new_n3963_, new_n3964_, new_n3965_,
    new_n3966_, new_n3967_, new_n3968_, new_n3969_, new_n3970_, new_n3971_,
    new_n3972_, new_n3973_, new_n3974_, new_n3975_, new_n3976_, new_n3977_,
    new_n3978_, new_n3979_, new_n3980_, new_n3981_, new_n3982_, new_n3983_,
    new_n3984_, new_n3985_, new_n3986_, new_n3987_, new_n3988_, new_n3989_,
    new_n3990_, new_n3991_, new_n3992_, new_n3993_, new_n3994_, new_n3995_,
    new_n3996_, new_n3997_, new_n3998_, new_n3999_, new_n4000_, new_n4001_,
    new_n4002_, new_n4003_, new_n4004_, new_n4005_, new_n4006_, new_n4007_,
    new_n4008_, new_n4009_, new_n4010_, new_n4011_, new_n4012_, new_n4013_,
    new_n4014_, new_n4015_, new_n4016_, new_n4017_, new_n4018_, new_n4019_,
    new_n4020_, new_n4021_, new_n4022_, new_n4023_, new_n4024_, new_n4025_,
    new_n4026_, new_n4027_, new_n4028_, new_n4029_, new_n4030_, new_n4031_,
    new_n4032_, new_n4033_, new_n4034_, new_n4035_, new_n4036_, new_n4037_,
    new_n4038_, new_n4039_, new_n4040_, new_n4041_, new_n4042_, new_n4043_,
    new_n4044_, new_n4045_, new_n4046_, new_n4047_, new_n4048_, new_n4049_,
    new_n4050_, new_n4051_, new_n4052_, new_n4053_, new_n4054_, new_n4055_,
    new_n4056_, new_n4057_, new_n4058_, new_n4059_, new_n4060_, new_n4061_,
    new_n4062_, new_n4063_, new_n4064_, new_n4065_, new_n4066_, new_n4067_,
    new_n4068_, new_n4069_, new_n4070_, new_n4071_, new_n4072_, new_n4073_,
    new_n4074_, new_n4075_, new_n4076_, new_n4077_, new_n4078_, new_n4079_,
    new_n4080_, new_n4081_, new_n4082_, new_n4083_, new_n4084_, new_n4085_,
    new_n4086_, new_n4087_, new_n4088_, new_n4089_, new_n4090_, new_n4091_,
    new_n4092_, new_n4093_, new_n4094_, new_n4095_, new_n4096_, new_n4097_,
    new_n4098_, new_n4099_, new_n4100_, new_n4101_, new_n4102_, new_n4103_,
    new_n4104_, new_n4105_, new_n4106_, new_n4107_, new_n4108_, new_n4109_,
    new_n4110_, new_n4111_, new_n4112_, new_n4113_, new_n4114_, new_n4115_,
    new_n4116_, new_n4117_, new_n4118_, new_n4119_, new_n4120_, new_n4121_,
    new_n4122_, new_n4123_, new_n4124_, new_n4125_, new_n4126_, new_n4127_,
    new_n4128_, new_n4129_, new_n4130_, new_n4131_, new_n4132_, new_n4133_,
    new_n4134_, new_n4135_, new_n4136_, new_n4137_, new_n4138_, new_n4139_,
    new_n4140_, new_n4141_, new_n4142_, new_n4143_, new_n4144_, new_n4145_,
    new_n4146_, new_n4147_, new_n4148_, new_n4149_, new_n4150_, new_n4151_,
    new_n4152_, new_n4153_, new_n4154_, new_n4155_, new_n4156_, new_n4157_,
    new_n4158_, new_n4159_, new_n4160_, new_n4161_, new_n4162_, new_n4163_,
    new_n4164_, new_n4165_, new_n4166_, new_n4167_, new_n4168_, new_n4169_,
    new_n4170_, new_n4171_, new_n4172_, new_n4173_, new_n4174_, new_n4175_,
    new_n4176_, new_n4177_, new_n4178_, new_n4179_, new_n4180_, new_n4181_,
    new_n4182_, new_n4183_, new_n4184_, new_n4185_, new_n4186_, new_n4187_,
    new_n4188_, new_n4189_, new_n4190_, new_n4191_, new_n4192_, new_n4193_,
    new_n4194_, new_n4195_, new_n4196_, new_n4197_, new_n4198_, new_n4199_,
    new_n4200_, new_n4201_, new_n4202_, new_n4203_, new_n4204_, new_n4205_,
    new_n4206_, new_n4207_, new_n4208_, new_n4209_, new_n4210_, new_n4211_,
    new_n4212_, new_n4213_, new_n4214_, new_n4215_, new_n4216_, new_n4217_,
    new_n4218_, new_n4219_, new_n4220_, new_n4221_, new_n4222_, new_n4223_,
    new_n4224_, new_n4225_, new_n4226_, new_n4227_, new_n4228_, new_n4229_,
    new_n4230_, new_n4231_, new_n4232_, new_n4233_, new_n4234_, new_n4235_,
    new_n4236_, new_n4237_, new_n4238_, new_n4239_, new_n4240_, new_n4241_,
    new_n4242_, new_n4243_, new_n4244_, new_n4245_, new_n4246_, new_n4247_,
    new_n4248_, new_n4249_, new_n4250_, new_n4251_, new_n4252_, new_n4253_,
    new_n4254_, new_n4255_, new_n4256_, new_n4257_, new_n4258_, new_n4259_,
    new_n4260_, new_n4261_, new_n4262_, new_n4263_, new_n4264_, new_n4265_,
    new_n4266_, new_n4267_, new_n4268_, new_n4269_, new_n4270_, new_n4271_,
    new_n4272_, new_n4273_, new_n4274_, new_n4275_, new_n4276_, new_n4277_,
    new_n4278_, new_n4279_, new_n4280_, new_n4281_, new_n4282_, new_n4283_,
    new_n4284_, new_n4285_, new_n4286_, new_n4287_, new_n4288_, new_n4289_,
    new_n4290_, new_n4291_, new_n4292_, new_n4293_, new_n4294_, new_n4295_,
    new_n4296_, new_n4297_, new_n4298_, new_n4299_, new_n4300_, new_n4301_,
    new_n4302_, new_n4303_, new_n4304_, new_n4305_, new_n4306_, new_n4307_,
    new_n4308_, new_n4309_, new_n4310_, new_n4311_, new_n4312_, new_n4313_,
    new_n4314_, new_n4315_, new_n4316_, new_n4317_, new_n4318_, new_n4319_,
    new_n4320_, new_n4321_, new_n4322_, new_n4323_, new_n4324_, new_n4325_,
    new_n4326_, new_n4327_, new_n4328_, new_n4329_, new_n4330_, new_n4331_,
    new_n4332_, new_n4333_, new_n4334_, new_n4335_, new_n4336_, new_n4337_,
    new_n4338_, new_n4339_, new_n4340_, new_n4341_, new_n4342_, new_n4343_,
    new_n4344_, new_n4345_, new_n4346_, new_n4347_, new_n4348_, new_n4349_,
    new_n4350_, new_n4351_, new_n4352_, new_n4353_, new_n4354_, new_n4355_,
    new_n4356_, new_n4357_, new_n4358_, new_n4359_, new_n4360_, new_n4361_,
    new_n4362_, new_n4363_, new_n4364_, new_n4365_, new_n4366_, new_n4367_,
    new_n4368_, new_n4369_, new_n4370_, new_n4371_, new_n4372_, new_n4373_,
    new_n4374_, new_n4375_, new_n4376_, new_n4377_, new_n4378_, new_n4379_,
    new_n4380_, new_n4381_, new_n4382_, new_n4383_, new_n4384_, new_n4385_,
    new_n4386_, new_n4387_, new_n4388_, new_n4389_, new_n4390_, new_n4391_,
    new_n4392_, new_n4393_, new_n4394_, new_n4395_, new_n4396_, new_n4397_,
    new_n4398_, new_n4399_, new_n4400_, new_n4401_, new_n4402_, new_n4403_,
    new_n4404_, new_n4405_, new_n4406_, new_n4407_, new_n4408_, new_n4409_,
    new_n4410_, new_n4411_, new_n4412_, new_n4413_, new_n4414_, new_n4415_,
    new_n4416_, new_n4417_, new_n4418_, new_n4419_, new_n4420_, new_n4421_,
    new_n4422_, new_n4423_, new_n4424_, new_n4425_, new_n4426_, new_n4427_,
    new_n4428_, new_n4429_, new_n4430_, new_n4431_, new_n4432_, new_n4433_,
    new_n4434_, new_n4435_, new_n4436_, new_n4437_, new_n4438_, new_n4439_,
    new_n4440_, new_n4441_, new_n4442_, new_n4443_, new_n4444_, new_n4445_,
    new_n4446_, new_n4447_, new_n4448_, new_n4449_, new_n4450_, new_n4451_,
    new_n4452_, new_n4453_, new_n4454_, new_n4455_, new_n4456_, new_n4457_,
    new_n4458_, new_n4459_, new_n4460_, new_n4461_, new_n4462_, new_n4463_,
    new_n4464_, new_n4465_, new_n4466_, new_n4467_, new_n4468_, new_n4469_,
    new_n4470_, new_n4471_, new_n4472_, new_n4473_, new_n4474_, new_n4475_,
    new_n4476_, new_n4477_, new_n4478_, new_n4479_, new_n4480_, new_n4481_,
    new_n4482_, new_n4483_, new_n4484_, new_n4485_, new_n4486_, new_n4487_,
    new_n4488_, new_n4489_, new_n4490_, new_n4491_, new_n4492_, new_n4493_,
    new_n4494_, new_n4495_, new_n4496_, new_n4497_, new_n4498_, new_n4499_,
    new_n4500_, new_n4501_, new_n4502_, new_n4503_, new_n4504_, new_n4505_,
    new_n4506_, new_n4507_, new_n4508_, new_n4509_, new_n4510_, new_n4511_,
    new_n4512_, new_n4513_, new_n4514_, new_n4515_, new_n4516_, new_n4517_,
    new_n4518_, new_n4519_, new_n4520_, new_n4521_, new_n4522_, new_n4523_,
    new_n4524_, new_n4525_, new_n4526_, new_n4527_, new_n4528_, new_n4529_,
    new_n4530_, new_n4531_, new_n4532_, new_n4533_, new_n4534_, new_n4535_,
    new_n4536_, new_n4537_, new_n4538_, new_n4539_, new_n4540_, new_n4541_,
    new_n4542_, new_n4543_, new_n4544_, new_n4545_, new_n4546_, new_n4547_,
    new_n4548_, new_n4549_, new_n4550_, new_n4551_, new_n4552_, new_n4553_,
    new_n4554_, new_n4555_, new_n4556_, new_n4557_, new_n4558_, new_n4559_,
    new_n4560_, new_n4561_, new_n4562_, new_n4563_, new_n4564_, new_n4565_,
    new_n4566_, new_n4567_, new_n4568_, new_n4569_, new_n4570_, new_n4571_,
    new_n4572_, new_n4573_, new_n4574_, new_n4575_, new_n4576_, new_n4577_,
    new_n4578_, new_n4579_, new_n4580_, new_n4581_, new_n4582_, new_n4583_,
    new_n4584_, new_n4585_, new_n4586_, new_n4587_, new_n4588_, new_n4589_,
    new_n4590_, new_n4591_, new_n4592_, new_n4593_, new_n4594_, new_n4595_,
    new_n4596_, new_n4597_, new_n4598_, new_n4599_, new_n4600_, new_n4601_,
    new_n4602_, new_n4603_, new_n4604_, new_n4605_, new_n4606_, new_n4607_,
    new_n4608_, new_n4609_, new_n4610_, new_n4611_, new_n4612_, new_n4613_,
    new_n4614_, new_n4615_, new_n4616_, new_n4617_, new_n4618_, new_n4619_,
    new_n4620_, new_n4621_, new_n4622_, new_n4623_, new_n4624_, new_n4625_,
    new_n4626_, new_n4627_, new_n4628_, new_n4629_, new_n4630_, new_n4631_,
    new_n4632_, new_n4633_, new_n4634_, new_n4635_, new_n4636_, new_n4637_,
    new_n4638_, new_n4639_, new_n4640_, new_n4641_, new_n4642_, new_n4643_,
    new_n4644_, new_n4645_, new_n4646_, new_n4647_, new_n4648_, new_n4649_,
    new_n4650_, new_n4651_, new_n4652_, new_n4653_, new_n4654_, new_n4655_,
    new_n4656_, new_n4657_, new_n4658_, new_n4659_, new_n4660_, new_n4661_,
    new_n4662_, new_n4663_, new_n4664_, new_n4665_, new_n4666_, new_n4667_,
    new_n4668_, new_n4669_, new_n4670_, new_n4671_, new_n4672_, new_n4673_,
    new_n4674_, new_n4675_, new_n4676_, new_n4677_, new_n4678_, new_n4679_,
    new_n4680_, new_n4681_, new_n4682_, new_n4683_, new_n4684_, new_n4685_,
    new_n4686_, new_n4687_, new_n4688_, new_n4689_, new_n4690_, new_n4691_,
    new_n4692_, new_n4693_, new_n4694_, new_n4695_, new_n4696_, new_n4697_,
    new_n4698_, new_n4699_, new_n4700_, new_n4701_, new_n4702_, new_n4703_,
    new_n4704_, new_n4705_, new_n4706_, new_n4707_, new_n4708_, new_n4709_,
    new_n4710_, new_n4711_, new_n4712_, new_n4713_, new_n4714_, new_n4715_,
    new_n4716_, new_n4717_, new_n4718_, new_n4719_, new_n4720_, new_n4721_,
    new_n4722_, new_n4723_, new_n4724_, new_n4725_, new_n4726_, new_n4727_,
    new_n4728_, new_n4729_, new_n4730_, new_n4731_, new_n4732_, new_n4733_,
    new_n4734_, new_n4735_, new_n4736_, new_n4737_, new_n4738_, new_n4739_,
    new_n4740_, new_n4741_, new_n4742_, new_n4743_, new_n4744_, new_n4745_,
    new_n4746_, new_n4747_, new_n4748_, new_n4749_, new_n4750_, new_n4751_,
    new_n4752_, new_n4753_, new_n4754_, new_n4755_, new_n4756_, new_n4757_,
    new_n4758_, new_n4759_, new_n4760_, new_n4761_, new_n4762_, new_n4763_,
    new_n4764_, new_n4765_, new_n4766_, new_n4767_, new_n4768_, new_n4769_,
    new_n4770_, new_n4771_, new_n4772_, new_n4773_, new_n4774_, new_n4775_,
    new_n4776_, new_n4777_, new_n4778_, new_n4779_, new_n4780_, new_n4781_,
    new_n4782_, new_n4783_, new_n4784_, new_n4785_, new_n4786_, new_n4787_,
    new_n4788_, new_n4789_, new_n4790_, new_n4791_, new_n4792_, new_n4793_,
    new_n4794_, new_n4795_, new_n4796_, new_n4797_, new_n4798_, new_n4799_,
    new_n4800_, new_n4801_, new_n4802_, new_n4803_, new_n4804_, new_n4805_,
    new_n4806_, new_n4807_, new_n4808_, new_n4809_, new_n4810_, new_n4811_,
    new_n4812_, new_n4813_, new_n4814_, new_n4815_, new_n4816_, new_n4817_,
    new_n4818_, new_n4819_, new_n4820_, new_n4821_, new_n4822_, new_n4823_,
    new_n4824_, new_n4825_, new_n4826_, new_n4827_, new_n4828_, new_n4829_,
    new_n4830_, new_n4831_, new_n4832_, new_n4833_, new_n4834_, new_n4835_,
    new_n4836_, new_n4837_, new_n4838_, new_n4839_, new_n4840_, new_n4841_,
    new_n4842_, new_n4843_, new_n4844_, new_n4845_, new_n4846_, new_n4847_,
    new_n4848_, new_n4849_, new_n4850_, new_n4851_, new_n4852_, new_n4853_,
    new_n4854_, new_n4855_, new_n4856_, new_n4857_, new_n4858_, new_n4859_,
    new_n4860_, new_n4861_, new_n4862_, new_n4863_, new_n4864_, new_n4865_,
    new_n4866_, new_n4867_, new_n4868_, new_n4869_, new_n4870_, new_n4871_,
    new_n4872_, new_n4873_, new_n4874_, new_n4875_, new_n4876_, new_n4877_,
    new_n4878_, new_n4879_, new_n4880_, new_n4881_, new_n4882_, new_n4883_,
    new_n4884_, new_n4885_, new_n4886_, new_n4887_, new_n4888_, new_n4889_,
    new_n4890_, new_n4891_, new_n4892_, new_n4893_, new_n4894_, new_n4895_,
    new_n4896_, new_n4897_, new_n4898_, new_n4899_, new_n4900_, new_n4901_,
    new_n4902_, new_n4903_, new_n4904_, new_n4905_, new_n4906_, new_n4907_,
    new_n4908_, new_n4909_, new_n4910_, new_n4911_, new_n4912_, new_n4913_,
    new_n4914_, new_n4915_, new_n4916_, new_n4917_, new_n4918_, new_n4919_,
    new_n4920_, new_n4921_, new_n4922_, new_n4923_, new_n4924_, new_n4925_,
    new_n4926_, new_n4927_, new_n4928_, new_n4929_, new_n4930_, new_n4931_,
    new_n4932_, new_n4933_, new_n4934_, new_n4935_, new_n4936_, new_n4937_,
    new_n4938_, new_n4939_, new_n4940_, new_n4941_, new_n4942_, new_n4943_,
    new_n4944_, new_n4945_, new_n4946_, new_n4947_, new_n4948_, new_n4949_,
    new_n4950_, new_n4951_, new_n4952_, new_n4953_, new_n4954_, new_n4955_,
    new_n4956_, new_n4957_, new_n4958_, new_n4959_, new_n4960_, new_n4961_,
    new_n4962_, new_n4963_, new_n4964_, new_n4965_, new_n4966_, new_n4967_,
    new_n4968_, new_n4969_, new_n4970_, new_n4971_, new_n4972_, new_n4973_,
    new_n4974_, new_n4975_, new_n4976_, new_n4977_, new_n4978_, new_n4979_,
    new_n4980_, new_n4981_, new_n4982_, new_n4983_, new_n4984_, new_n4985_,
    new_n4986_, new_n4987_, new_n4988_, new_n4989_, new_n4990_, new_n4991_,
    new_n4992_, new_n4993_, new_n4994_, new_n4995_, new_n4996_, new_n4997_,
    new_n4998_, new_n4999_, new_n5000_, new_n5001_, new_n5002_, new_n5003_,
    new_n5004_, new_n5005_, new_n5006_, new_n5007_, new_n5008_, new_n5009_,
    new_n5010_, new_n5011_, new_n5012_, new_n5013_, new_n5014_, new_n5015_,
    new_n5016_, new_n5017_, new_n5018_, new_n5019_, new_n5020_, new_n5021_,
    new_n5022_, new_n5023_, new_n5024_, new_n5025_, new_n5026_, new_n5027_,
    new_n5028_, new_n5029_, new_n5030_, new_n5031_, new_n5032_, new_n5033_,
    new_n5034_, new_n5035_, new_n5036_, new_n5037_, new_n5038_, new_n5039_,
    new_n5040_, new_n5041_, new_n5042_, new_n5043_, new_n5044_, new_n5045_,
    new_n5046_, new_n5047_, new_n5048_, new_n5049_, new_n5050_, new_n5051_,
    new_n5052_, new_n5053_, new_n5054_, new_n5055_, new_n5056_, new_n5057_,
    new_n5058_, new_n5059_, new_n5060_, new_n5061_, new_n5062_, new_n5063_,
    new_n5064_, new_n5065_, new_n5066_, new_n5067_, new_n5068_, new_n5069_,
    new_n5070_, new_n5071_, new_n5072_, new_n5073_, new_n5074_, new_n5075_,
    new_n5076_, new_n5077_, new_n5078_, new_n5079_, new_n5080_, new_n5081_,
    new_n5082_, new_n5083_, new_n5084_, new_n5085_, new_n5086_, new_n5087_,
    new_n5088_, new_n5089_, new_n5090_, new_n5091_, new_n5092_, new_n5093_,
    new_n5094_, new_n5095_, new_n5096_, new_n5097_, new_n5098_, new_n5099_,
    new_n5100_, new_n5101_, new_n5102_, new_n5103_, new_n5104_, new_n5105_,
    new_n5106_, new_n5107_, new_n5108_, new_n5109_, new_n5110_, new_n5111_,
    new_n5112_, new_n5113_, new_n5114_, new_n5115_, new_n5116_, new_n5117_,
    new_n5118_, new_n5119_, new_n5120_, new_n5121_, new_n5122_, new_n5123_,
    new_n5124_, new_n5125_, new_n5126_, new_n5127_, new_n5128_, new_n5129_,
    new_n5130_, new_n5131_, new_n5132_, new_n5133_, new_n5134_, new_n5135_,
    new_n5136_, new_n5137_, new_n5138_, new_n5139_, new_n5140_, new_n5141_,
    new_n5142_, new_n5143_, new_n5144_, new_n5145_, new_n5146_, new_n5147_,
    new_n5148_, new_n5149_, new_n5150_, new_n5151_, new_n5152_, new_n5153_,
    new_n5154_, new_n5155_, new_n5156_, new_n5157_, new_n5158_, new_n5159_,
    new_n5160_, new_n5161_, new_n5162_, new_n5163_, new_n5164_, new_n5165_,
    new_n5166_, new_n5167_, new_n5168_, new_n5169_, new_n5170_, new_n5171_,
    new_n5172_, new_n5173_, new_n5174_, new_n5175_, new_n5176_, new_n5177_,
    new_n5178_, new_n5179_, new_n5180_, new_n5181_, new_n5182_, new_n5183_,
    new_n5184_, new_n5185_, new_n5186_, new_n5187_, new_n5188_, new_n5189_,
    new_n5190_, new_n5191_, new_n5192_, new_n5193_, new_n5194_, new_n5195_,
    new_n5196_, new_n5197_, new_n5198_, new_n5199_, new_n5200_, new_n5201_,
    new_n5202_, new_n5203_, new_n5204_, new_n5205_, new_n5206_, new_n5207_,
    new_n5208_, new_n5209_, new_n5210_, new_n5211_, new_n5212_, new_n5213_,
    new_n5214_, new_n5215_, new_n5216_, new_n5217_, new_n5218_, new_n5219_,
    new_n5220_, new_n5221_, new_n5222_, new_n5223_, new_n5224_, new_n5225_,
    new_n5226_, new_n5227_, new_n5228_, new_n5229_, new_n5230_, new_n5231_,
    new_n5232_, new_n5233_, new_n5234_, new_n5235_, new_n5236_, new_n5237_,
    new_n5238_, new_n5239_, new_n5240_, new_n5241_, new_n5242_, new_n5243_,
    new_n5244_, new_n5245_, new_n5246_, new_n5247_, new_n5248_, new_n5249_,
    new_n5250_, new_n5251_, new_n5252_, new_n5253_, new_n5254_, new_n5255_,
    new_n5256_, new_n5257_, new_n5258_, new_n5259_, new_n5260_, new_n5261_,
    new_n5262_, new_n5263_, new_n5264_, new_n5265_, new_n5266_, new_n5267_,
    new_n5268_, new_n5269_, new_n5270_, new_n5271_, new_n5272_, new_n5273_,
    new_n5274_, new_n5275_, new_n5276_, new_n5277_, new_n5278_, new_n5279_,
    new_n5280_, new_n5281_, new_n5282_, new_n5283_, new_n5284_, new_n5285_,
    new_n5286_, new_n5287_, new_n5288_, new_n5289_, new_n5290_, new_n5291_,
    new_n5292_, new_n5293_, new_n5294_, new_n5295_, new_n5296_, new_n5297_,
    new_n5298_, new_n5299_, new_n5300_, new_n5301_, new_n5302_, new_n5303_,
    new_n5304_, new_n5305_, new_n5306_, new_n5307_, new_n5308_, new_n5309_,
    new_n5310_, new_n5311_, new_n5312_, new_n5313_, new_n5314_, new_n5315_,
    new_n5316_, new_n5317_, new_n5318_, new_n5319_, new_n5320_, new_n5321_,
    new_n5322_, new_n5323_, new_n5324_, new_n5325_, new_n5326_, new_n5327_,
    new_n5328_, new_n5329_, new_n5330_, new_n5331_, new_n5332_, new_n5333_,
    new_n5334_, new_n5335_, new_n5336_, new_n5337_, new_n5338_, new_n5339_,
    new_n5340_, new_n5341_, new_n5342_, new_n5343_, new_n5344_, new_n5345_,
    new_n5346_, new_n5347_, new_n5348_, new_n5349_, new_n5350_, new_n5351_,
    new_n5352_, new_n5353_, new_n5354_, new_n5355_, new_n5356_, new_n5357_,
    new_n5358_, new_n5359_, new_n5360_, new_n5361_, new_n5362_, new_n5363_,
    new_n5364_, new_n5365_, new_n5366_, new_n5367_, new_n5368_, new_n5369_,
    new_n5370_, new_n5371_, new_n5372_, new_n5373_, new_n5374_, new_n5375_,
    new_n5376_, new_n5377_, new_n5378_, new_n5379_, new_n5380_, new_n5381_,
    new_n5382_, new_n5383_, new_n5384_, new_n5385_, new_n5386_, new_n5387_,
    new_n5388_, new_n5389_, new_n5390_, new_n5391_, new_n5392_, new_n5393_,
    new_n5394_, new_n5395_, new_n5396_, new_n5397_, new_n5398_, new_n5399_,
    new_n5400_, new_n5401_, new_n5402_, new_n5403_, new_n5404_, new_n5405_,
    new_n5406_, new_n5407_, new_n5408_, new_n5409_, new_n5410_, new_n5411_,
    new_n5412_, new_n5413_, new_n5414_, new_n5415_, new_n5416_, new_n5417_,
    new_n5418_, new_n5419_, new_n5420_, new_n5421_, new_n5422_, new_n5423_,
    new_n5424_, new_n5425_, new_n5426_, new_n5427_, new_n5428_, new_n5429_,
    new_n5430_, new_n5431_, new_n5432_, new_n5433_, new_n5434_, new_n5435_,
    new_n5436_, new_n5437_, new_n5438_, new_n5439_, new_n5440_, new_n5441_,
    new_n5442_, new_n5443_, new_n5444_, new_n5445_, new_n5446_, new_n5447_,
    new_n5448_, new_n5449_, new_n5450_, new_n5451_, new_n5452_, new_n5453_,
    new_n5454_, new_n5455_, new_n5456_, new_n5457_, new_n5458_, new_n5459_,
    new_n5460_, new_n5461_, new_n5462_, new_n5463_, new_n5464_, new_n5465_,
    new_n5466_, new_n5467_, new_n5468_, new_n5469_, new_n5470_, new_n5471_,
    new_n5472_, new_n5473_, new_n5474_, new_n5475_, new_n5476_, new_n5477_,
    new_n5478_, new_n5479_, new_n5480_, new_n5481_, new_n5482_, new_n5483_,
    new_n5484_, new_n5485_, new_n5486_, new_n5487_, new_n5488_, new_n5489_,
    new_n5490_, new_n5491_, new_n5492_, new_n5493_, new_n5494_, new_n5495_,
    new_n5496_, new_n5497_, new_n5498_, new_n5499_, new_n5500_, new_n5501_,
    new_n5502_, new_n5503_, new_n5504_, new_n5505_, new_n5506_, new_n5507_,
    new_n5508_, new_n5509_, new_n5510_, new_n5511_, new_n5512_, new_n5513_,
    new_n5514_, new_n5515_, new_n5516_, new_n5517_, new_n5518_, new_n5519_,
    new_n5520_, new_n5521_, new_n5522_, new_n5523_, new_n5524_, new_n5525_,
    new_n5526_, new_n5527_, new_n5528_, new_n5529_, new_n5530_, new_n5531_,
    new_n5532_, new_n5533_, new_n5534_, new_n5535_, new_n5536_, new_n5537_,
    new_n5538_, new_n5539_, new_n5540_, new_n5541_, new_n5542_, new_n5543_,
    new_n5544_, new_n5545_, new_n5546_, new_n5547_, new_n5548_, new_n5549_,
    new_n5550_, new_n5551_, new_n5552_, new_n5553_, new_n5554_, new_n5555_,
    new_n5556_, new_n5557_, new_n5558_, new_n5559_, new_n5560_, new_n5561_,
    new_n5562_, new_n5563_, new_n5564_, new_n5565_, new_n5566_, new_n5567_,
    new_n5568_, new_n5569_, new_n5570_, new_n5571_, new_n5572_, new_n5573_,
    new_n5574_, new_n5575_, new_n5576_, new_n5577_, new_n5578_, new_n5579_,
    new_n5580_, new_n5581_, new_n5582_, new_n5583_, new_n5584_, new_n5585_,
    new_n5586_, new_n5587_, new_n5588_, new_n5589_, new_n5590_, new_n5591_,
    new_n5592_, new_n5593_, new_n5594_, new_n5595_, new_n5596_, new_n5597_,
    new_n5598_, new_n5599_, new_n5600_, new_n5601_, new_n5602_, new_n5603_,
    new_n5604_, new_n5605_, new_n5606_, new_n5607_, new_n5608_, new_n5609_,
    new_n5610_, new_n5611_, new_n5612_, new_n5613_, new_n5614_, new_n5615_,
    new_n5616_, new_n5617_, new_n5618_, new_n5619_, new_n5620_, new_n5621_,
    new_n5622_, new_n5623_, new_n5624_, new_n5625_, new_n5626_, new_n5627_,
    new_n5628_, new_n5629_, new_n5630_, new_n5631_, new_n5632_, new_n5633_,
    new_n5634_, new_n5635_, new_n5636_, new_n5637_, new_n5638_, new_n5639_,
    new_n5640_, new_n5641_, new_n5642_, new_n5643_, new_n5644_, new_n5645_,
    new_n5646_, new_n5647_, new_n5648_, new_n5649_, new_n5650_, new_n5651_,
    new_n5652_, new_n5653_, new_n5654_, new_n5655_, new_n5656_, new_n5657_,
    new_n5658_, new_n5659_, new_n5660_, new_n5661_, new_n5662_, new_n5663_,
    new_n5664_, new_n5665_, new_n5666_, new_n5667_, new_n5668_, new_n5669_,
    new_n5670_, new_n5671_, new_n5672_, new_n5673_, new_n5674_, new_n5675_,
    new_n5676_, new_n5677_, new_n5678_, new_n5679_, new_n5680_, new_n5681_,
    new_n5682_, new_n5683_, new_n5684_, new_n5685_, new_n5686_, new_n5687_,
    new_n5688_, new_n5689_, new_n5690_, new_n5691_, new_n5692_, new_n5693_,
    new_n5694_, new_n5695_, new_n5696_, new_n5697_, new_n5698_, new_n5699_,
    new_n5700_, new_n5701_, new_n5702_, new_n5703_, new_n5704_, new_n5705_,
    new_n5706_, new_n5707_, new_n5708_, new_n5709_, new_n5710_, new_n5711_,
    new_n5712_, new_n5713_, new_n5714_, new_n5715_, new_n5716_, new_n5717_,
    new_n5718_, new_n5719_, new_n5720_, new_n5721_, new_n5722_, new_n5723_,
    new_n5724_, new_n5725_, new_n5726_, new_n5727_, new_n5728_, new_n5729_,
    new_n5730_, new_n5731_, new_n5732_, new_n5733_, new_n5734_, new_n5735_,
    new_n5736_, new_n5737_, new_n5738_, new_n5739_, new_n5740_, new_n5741_,
    new_n5742_, new_n5743_, new_n5744_, new_n5745_, new_n5746_, new_n5747_,
    new_n5748_, new_n5749_, new_n5750_, new_n5751_, new_n5752_, new_n5753_,
    new_n5754_, new_n5755_, new_n5756_, new_n5757_, new_n5758_, new_n5759_,
    new_n5760_, new_n5761_, new_n5762_, new_n5763_, new_n5764_, new_n5765_,
    new_n5766_, new_n5767_, new_n5768_, new_n5769_, new_n5770_, new_n5771_,
    new_n5772_, new_n5773_, new_n5774_, new_n5775_, new_n5776_, new_n5777_,
    new_n5778_, new_n5779_, new_n5780_, new_n5781_, new_n5782_, new_n5783_,
    new_n5784_, new_n5785_, new_n5786_, new_n5787_, new_n5788_, new_n5789_,
    new_n5790_, new_n5791_, new_n5792_, new_n5793_, new_n5794_, new_n5795_,
    new_n5796_, new_n5797_, new_n5798_, new_n5799_, new_n5800_, new_n5801_,
    new_n5802_, new_n5803_, new_n5804_, new_n5805_, new_n5806_, new_n5807_,
    new_n5808_, new_n5809_, new_n5810_, new_n5811_, new_n5812_, new_n5813_,
    new_n5814_, new_n5815_, new_n5816_, new_n5817_, new_n5818_, new_n5819_,
    new_n5820_, new_n5821_, new_n5822_, new_n5823_, new_n5824_, new_n5825_,
    new_n5826_, new_n5827_, new_n5828_, new_n5829_, new_n5830_, new_n5831_,
    new_n5832_, new_n5833_, new_n5834_, new_n5835_, new_n5836_, new_n5837_,
    new_n5838_, new_n5839_, new_n5840_, new_n5841_, new_n5842_, new_n5843_,
    new_n5844_, new_n5845_, new_n5846_, new_n5847_, new_n5848_, new_n5849_,
    new_n5850_, new_n5851_, new_n5852_, new_n5853_, new_n5854_, new_n5855_,
    new_n5856_, new_n5857_, new_n5858_, new_n5859_, new_n5860_, new_n5861_,
    new_n5862_, new_n5863_, new_n5864_, new_n5865_, new_n5866_, new_n5867_,
    new_n5868_, new_n5869_, new_n5870_, new_n5871_, new_n5872_, new_n5873_,
    new_n5874_, new_n5875_, new_n5876_, new_n5877_, new_n5878_, new_n5879_,
    new_n5880_, new_n5881_, new_n5882_, new_n5883_, new_n5884_, new_n5885_,
    new_n5886_, new_n5887_, new_n5888_, new_n5889_, new_n5890_, new_n5891_,
    new_n5892_, new_n5893_, new_n5894_, new_n5895_, new_n5896_, new_n5897_,
    new_n5898_, new_n5899_, new_n5900_, new_n5901_, new_n5902_, new_n5903_,
    new_n5904_, new_n5905_, new_n5906_, new_n5907_, new_n5908_, new_n5909_,
    new_n5910_, new_n5911_, new_n5912_, new_n5913_, new_n5914_, new_n5915_,
    new_n5916_, new_n5917_, new_n5918_, new_n5919_, new_n5920_, new_n5921_,
    new_n5922_, new_n5923_, new_n5924_, new_n5925_, new_n5926_, new_n5927_,
    new_n5928_, new_n5929_, new_n5930_, new_n5931_, new_n5932_, new_n5933_,
    new_n5934_, new_n5935_, new_n5936_, new_n5937_, new_n5938_, new_n5939_,
    new_n5940_, new_n5941_, new_n5942_, new_n5943_, new_n5944_, new_n5945_,
    new_n5946_, new_n5947_, new_n5948_, new_n5949_, new_n5950_, new_n5951_,
    new_n5952_, new_n5953_, new_n5954_, new_n5955_, new_n5956_, new_n5957_,
    new_n5958_, new_n5959_, new_n5960_, new_n5961_, new_n5962_, new_n5963_,
    new_n5964_, new_n5965_, new_n5966_, new_n5967_, new_n5968_, new_n5969_,
    new_n5970_, new_n5971_, new_n5972_, new_n5973_, new_n5974_, new_n5975_,
    new_n5976_, new_n5977_, new_n5978_, new_n5979_, new_n5980_, new_n5981_,
    new_n5982_, new_n5983_, new_n5984_, new_n5985_, new_n5986_, new_n5987_,
    new_n5988_, new_n5989_, new_n5990_, new_n5991_, new_n5992_, new_n5993_,
    new_n5994_, new_n5995_, new_n5996_, new_n5997_, new_n5998_, new_n5999_,
    new_n6000_, new_n6001_, new_n6002_, new_n6003_, new_n6004_, new_n6005_,
    new_n6006_, new_n6007_, new_n6008_, new_n6009_, new_n6010_, new_n6011_,
    new_n6012_, new_n6013_, new_n6014_, new_n6015_, new_n6016_, new_n6017_,
    new_n6018_, new_n6019_, new_n6020_, new_n6021_, new_n6022_, new_n6023_,
    new_n6024_, new_n6025_, new_n6026_, new_n6027_, new_n6028_, new_n6029_,
    new_n6030_, new_n6031_, new_n6032_, new_n6033_, new_n6034_, new_n6035_,
    new_n6036_, new_n6037_, new_n6038_, new_n6039_, new_n6040_, new_n6041_,
    new_n6042_, new_n6043_, new_n6044_, new_n6045_, new_n6046_, new_n6047_,
    new_n6048_, new_n6049_, new_n6050_, new_n6051_, new_n6052_, new_n6053_,
    new_n6054_, new_n6055_, new_n6056_, new_n6057_, new_n6058_, new_n6059_,
    new_n6060_, new_n6061_, new_n6062_, new_n6063_, new_n6064_, new_n6065_,
    new_n6066_, new_n6067_, new_n6068_, new_n6069_, new_n6070_, new_n6071_,
    new_n6072_, new_n6073_, new_n6074_, new_n6075_, new_n6076_, new_n6077_,
    new_n6078_, new_n6079_, new_n6080_, new_n6081_, new_n6082_, new_n6083_,
    new_n6084_, new_n6085_, new_n6086_, new_n6087_, new_n6088_, new_n6089_,
    new_n6090_, new_n6091_, new_n6092_, new_n6093_, new_n6094_, new_n6095_,
    new_n6096_, new_n6097_, new_n6098_, new_n6099_, new_n6100_, new_n6101_,
    new_n6102_, new_n6103_, new_n6104_, new_n6105_, new_n6106_, new_n6107_,
    new_n6108_, new_n6109_, new_n6110_, new_n6111_, new_n6112_, new_n6113_,
    new_n6114_, new_n6115_, new_n6116_, new_n6117_, new_n6118_, new_n6119_,
    new_n6120_, new_n6121_, new_n6122_, new_n6123_, new_n6124_, new_n6125_,
    new_n6126_, new_n6127_, new_n6128_, new_n6129_, new_n6130_, new_n6131_,
    new_n6132_, new_n6133_, new_n6134_, new_n6135_, new_n6136_, new_n6137_,
    new_n6138_, new_n6139_, new_n6140_, new_n6141_, new_n6142_, new_n6143_,
    new_n6144_, new_n6145_, new_n6146_, new_n6147_, new_n6148_, new_n6149_,
    new_n6150_, new_n6151_, new_n6152_, new_n6153_, new_n6154_, new_n6155_,
    new_n6156_, new_n6157_, new_n6158_, new_n6159_, new_n6160_, new_n6161_,
    new_n6162_, new_n6163_, new_n6164_, new_n6165_, new_n6166_, new_n6167_,
    new_n6168_, new_n6169_, new_n6170_, new_n6171_, new_n6172_, new_n6173_,
    new_n6174_, new_n6175_, new_n6176_, new_n6177_, new_n6178_, new_n6179_,
    new_n6180_, new_n6181_, new_n6182_, new_n6183_, new_n6184_, new_n6185_,
    new_n6186_, new_n6187_, new_n6188_, new_n6189_, new_n6190_, new_n6191_,
    new_n6192_, new_n6193_, new_n6194_, new_n6195_, new_n6196_, new_n6197_,
    new_n6198_, new_n6199_, new_n6200_, new_n6201_, new_n6202_, new_n6203_,
    new_n6204_, new_n6205_, new_n6206_, new_n6207_, new_n6208_, new_n6209_,
    new_n6210_, new_n6211_, new_n6212_, new_n6213_, new_n6214_, new_n6215_,
    new_n6216_, new_n6217_, new_n6218_, new_n6219_, new_n6220_, new_n6221_,
    new_n6222_, new_n6223_, new_n6224_, new_n6225_, new_n6226_, new_n6227_,
    new_n6228_, new_n6229_, new_n6230_, new_n6231_, new_n6232_, new_n6233_,
    new_n6234_, new_n6235_, new_n6236_, new_n6237_, new_n6238_, new_n6239_,
    new_n6240_, new_n6241_, new_n6242_, new_n6243_, new_n6244_, new_n6245_,
    new_n6246_, new_n6247_, new_n6248_, new_n6249_, new_n6250_, new_n6251_,
    new_n6252_, new_n6253_, new_n6254_, new_n6255_, new_n6256_, new_n6257_,
    new_n6258_, new_n6259_, new_n6260_, new_n6261_, new_n6262_, new_n6263_,
    new_n6264_, new_n6265_, new_n6266_, new_n6267_, new_n6268_, new_n6269_,
    new_n6270_, new_n6271_, new_n6272_, new_n6273_, new_n6274_, new_n6275_,
    new_n6276_, new_n6277_, new_n6278_, new_n6279_, new_n6280_, new_n6281_,
    new_n6282_, new_n6283_, new_n6284_, new_n6285_, new_n6286_, new_n6287_,
    new_n6288_, new_n6289_, new_n6290_, new_n6291_, new_n6292_, new_n6293_,
    new_n6294_, new_n6295_, new_n6296_, new_n6297_, new_n6298_, new_n6299_,
    new_n6300_, new_n6301_, new_n6302_, new_n6303_, new_n6304_, new_n6305_,
    new_n6306_, new_n6307_, new_n6308_, new_n6309_, new_n6310_, new_n6311_,
    new_n6312_, new_n6313_, new_n6314_, new_n6315_, new_n6316_, new_n6317_,
    new_n6318_, new_n6319_, new_n6320_, new_n6321_, new_n6322_, new_n6323_,
    new_n6324_, new_n6325_, new_n6326_, new_n6327_, new_n6328_, new_n6329_,
    new_n6330_, new_n6331_, new_n6332_, new_n6333_, new_n6334_, new_n6335_,
    new_n6336_, new_n6337_, new_n6338_, new_n6339_, new_n6340_, new_n6341_,
    new_n6342_, new_n6343_, new_n6344_, new_n6345_, new_n6346_, new_n6347_,
    new_n6348_, new_n6349_, new_n6350_, new_n6351_, new_n6352_, new_n6353_,
    new_n6354_, new_n6355_, new_n6356_, new_n6357_, new_n6358_, new_n6359_,
    new_n6360_, new_n6361_, new_n6362_, new_n6363_, new_n6364_, new_n6365_,
    new_n6366_, new_n6367_, new_n6368_, new_n6369_, new_n6370_, new_n6371_,
    new_n6372_, new_n6373_, new_n6374_, new_n6375_, new_n6376_, new_n6377_,
    new_n6378_, new_n6379_, new_n6380_, new_n6381_, new_n6382_, new_n6383_,
    new_n6384_, new_n6385_, new_n6386_, new_n6387_, new_n6388_, new_n6389_,
    new_n6390_, new_n6391_, new_n6392_, new_n6393_, new_n6394_, new_n6395_,
    new_n6396_, new_n6397_, new_n6398_, new_n6399_, new_n6400_, new_n6401_,
    new_n6402_, new_n6403_, new_n6404_, new_n6405_, new_n6406_, new_n6407_,
    new_n6408_, new_n6409_, new_n6410_, new_n6411_, new_n6412_, new_n6413_,
    new_n6414_, new_n6415_, new_n6416_, new_n6417_, new_n6418_, new_n6419_,
    new_n6420_, new_n6421_, new_n6422_, new_n6423_, new_n6424_, new_n6425_,
    new_n6426_, new_n6427_, new_n6428_, new_n6429_, new_n6430_, new_n6431_,
    new_n6432_, new_n6433_, new_n6434_, new_n6435_, new_n6436_, new_n6437_,
    new_n6438_, new_n6439_, new_n6440_, new_n6441_, new_n6442_, new_n6443_,
    new_n6444_, new_n6445_, new_n6446_, new_n6447_, new_n6448_, new_n6449_,
    new_n6450_, new_n6451_, new_n6452_, new_n6453_, new_n6454_, new_n6455_,
    new_n6456_, new_n6457_, new_n6458_, new_n6459_, new_n6460_, new_n6461_,
    new_n6462_, new_n6463_, new_n6464_, new_n6465_, new_n6466_, new_n6467_,
    new_n6468_, new_n6469_, new_n6470_, new_n6471_, new_n6472_, new_n6473_,
    new_n6474_, new_n6475_, new_n6476_, new_n6477_, new_n6478_, new_n6479_,
    new_n6480_, new_n6481_, new_n6482_, new_n6483_, new_n6484_, new_n6485_,
    new_n6486_, new_n6487_, new_n6488_, new_n6489_, new_n6490_, new_n6491_,
    new_n6492_, new_n6493_, new_n6494_, new_n6495_, new_n6496_, new_n6497_,
    new_n6498_, new_n6499_, new_n6500_, new_n6501_, new_n6502_, new_n6503_,
    new_n6504_, new_n6505_, new_n6506_, new_n6507_, new_n6508_, new_n6509_,
    new_n6510_, new_n6511_, new_n6512_, new_n6513_, new_n6514_, new_n6515_,
    new_n6516_, new_n6517_, new_n6518_, new_n6519_, new_n6520_, new_n6521_,
    new_n6522_, new_n6523_, new_n6524_, new_n6525_, new_n6526_, new_n6527_,
    new_n6528_, new_n6529_, new_n6530_, new_n6531_, new_n6532_, new_n6533_,
    new_n6534_, new_n6535_, new_n6536_, new_n6537_, new_n6538_, new_n6539_,
    new_n6540_, new_n6541_, new_n6542_, new_n6543_, new_n6544_, new_n6545_,
    new_n6546_, new_n6547_, new_n6548_, new_n6549_, new_n6550_, new_n6551_,
    new_n6552_, new_n6553_, new_n6554_, new_n6555_, new_n6556_, new_n6557_,
    new_n6558_, new_n6559_, new_n6560_, new_n6561_, new_n6562_, new_n6563_,
    new_n6564_, new_n6565_, new_n6566_, new_n6567_, new_n6568_, new_n6569_,
    new_n6570_, new_n6571_, new_n6572_, new_n6573_, new_n6574_, new_n6575_,
    new_n6576_, new_n6577_, new_n6578_, new_n6579_, new_n6580_, new_n6581_,
    new_n6582_, new_n6583_, new_n6584_, new_n6585_, new_n6586_, new_n6587_,
    new_n6588_, new_n6589_, new_n6590_, new_n6591_, new_n6592_, new_n6593_,
    new_n6594_, new_n6595_, new_n6596_, new_n6597_, new_n6598_, new_n6599_,
    new_n6600_, new_n6601_, new_n6602_, new_n6603_, new_n6604_, new_n6605_,
    new_n6606_, new_n6607_, new_n6608_, new_n6609_, new_n6610_, new_n6611_,
    new_n6612_, new_n6613_, new_n6614_, new_n6615_, new_n6616_, new_n6617_,
    new_n6618_, new_n6619_, new_n6620_, new_n6621_, new_n6622_, new_n6623_,
    new_n6624_, new_n6625_, new_n6626_, new_n6627_, new_n6628_, new_n6629_,
    new_n6630_, new_n6631_, new_n6632_, new_n6633_, new_n6634_, new_n6635_,
    new_n6636_, new_n6637_, new_n6638_, new_n6639_, new_n6640_, new_n6641_,
    new_n6642_, new_n6643_, new_n6644_, new_n6645_, new_n6646_, new_n6647_,
    new_n6648_, new_n6649_, new_n6650_, new_n6651_, new_n6652_, new_n6653_,
    new_n6654_, new_n6655_, new_n6656_, new_n6657_, new_n6658_, new_n6659_,
    new_n6660_, new_n6661_, new_n6662_, new_n6663_, new_n6664_, new_n6665_,
    new_n6666_, new_n6667_, new_n6668_, new_n6669_, new_n6670_, new_n6671_,
    new_n6672_, new_n6673_, new_n6674_, new_n6675_, new_n6676_, new_n6677_,
    new_n6678_, new_n6679_, new_n6680_, new_n6681_, new_n6682_, new_n6683_,
    new_n6684_, new_n6685_, new_n6686_, new_n6687_, new_n6688_, new_n6689_,
    new_n6690_, new_n6691_, new_n6692_, new_n6693_, new_n6694_, new_n6695_,
    new_n6696_, new_n6697_, new_n6698_, new_n6699_, new_n6700_, new_n6701_,
    new_n6702_, new_n6703_, new_n6704_, new_n6705_, new_n6706_, new_n6707_,
    new_n6708_, new_n6709_, new_n6710_, new_n6711_, new_n6712_, new_n6713_,
    new_n6714_, new_n6715_, new_n6716_, new_n6717_, new_n6718_, new_n6719_,
    new_n6720_, new_n6721_, new_n6722_, new_n6723_, new_n6724_, new_n6725_,
    new_n6726_, new_n6727_, new_n6728_, new_n6729_, new_n6730_, new_n6731_,
    new_n6732_, new_n6733_, new_n6734_, new_n6735_, new_n6736_, new_n6737_,
    new_n6738_, new_n6739_, new_n6740_, new_n6741_, new_n6742_, new_n6743_,
    new_n6744_, new_n6745_, new_n6746_, new_n6747_, new_n6748_, new_n6749_,
    new_n6750_, new_n6751_, new_n6752_, new_n6753_, new_n6754_, new_n6755_,
    new_n6756_, new_n6757_, new_n6758_, new_n6759_, new_n6760_, new_n6761_,
    new_n6762_, new_n6763_, new_n6764_, new_n6765_, new_n6766_, new_n6767_,
    new_n6768_, new_n6769_, new_n6770_, new_n6771_, new_n6772_, new_n6773_,
    new_n6774_, new_n6775_, new_n6776_, new_n6777_, new_n6778_, new_n6779_,
    new_n6780_, new_n6781_, new_n6782_, new_n6783_, new_n6784_, new_n6785_,
    new_n6786_, new_n6787_, new_n6788_, new_n6789_, new_n6790_, new_n6791_,
    new_n6792_, new_n6793_, new_n6794_, new_n6795_, new_n6796_, new_n6797_,
    new_n6798_, new_n6799_, new_n6800_, new_n6801_, new_n6802_, new_n6803_,
    new_n6804_, new_n6805_, new_n6806_, new_n6807_, new_n6808_, new_n6809_,
    new_n6810_, new_n6811_, new_n6812_, new_n6813_, new_n6814_, new_n6815_,
    new_n6816_, new_n6817_, new_n6818_, new_n6819_, new_n6820_, new_n6821_,
    new_n6822_, new_n6823_, new_n6824_, new_n6825_, new_n6826_, new_n6827_,
    new_n6828_, new_n6829_, new_n6830_, new_n6831_, new_n6832_, new_n6833_,
    new_n6834_, new_n6835_, new_n6836_, new_n6837_, new_n6838_, new_n6839_,
    new_n6840_, new_n6841_, new_n6842_, new_n6843_, new_n6844_, new_n6845_,
    new_n6846_, new_n6847_, new_n6848_, new_n6849_, new_n6850_, new_n6851_,
    new_n6852_, new_n6853_, new_n6854_, new_n6855_, new_n6856_, new_n6857_,
    new_n6858_, new_n6859_, new_n6860_, new_n6861_, new_n6862_, new_n6863_,
    new_n6864_, new_n6865_, new_n6866_, new_n6867_, new_n6868_, new_n6869_,
    new_n6870_, new_n6871_, new_n6872_, new_n6873_, new_n6874_, new_n6875_,
    new_n6876_, new_n6877_, new_n6878_, new_n6879_, new_n6880_, new_n6881_,
    new_n6882_, new_n6883_, new_n6884_, new_n6885_, new_n6886_, new_n6887_,
    new_n6888_, new_n6889_, new_n6890_, new_n6891_, new_n6892_, new_n6893_,
    new_n6894_, new_n6895_, new_n6896_, new_n6897_, new_n6898_, new_n6899_,
    new_n6900_, new_n6901_, new_n6902_, new_n6903_, new_n6904_, new_n6905_,
    new_n6906_, new_n6907_, new_n6908_, new_n6909_, new_n6910_, new_n6911_,
    new_n6912_, new_n6913_, new_n6914_, new_n6915_, new_n6916_, new_n6917_,
    new_n6918_, new_n6919_, new_n6920_, new_n6921_, new_n6922_, new_n6923_,
    new_n6924_, new_n6925_, new_n6926_, new_n6927_, new_n6928_, new_n6929_,
    new_n6930_, new_n6931_, new_n6932_, new_n6933_, new_n6934_, new_n6935_,
    new_n6936_, new_n6937_, new_n6938_, new_n6939_, new_n6940_, new_n6941_,
    new_n6942_, new_n6943_, new_n6944_, new_n6945_, new_n6946_, new_n6947_,
    new_n6948_, new_n6949_, new_n6950_, new_n6951_, new_n6952_, new_n6953_,
    new_n6954_, new_n6955_, new_n6956_, new_n6957_, new_n6958_, new_n6959_,
    new_n6960_, new_n6961_, new_n6962_, new_n6963_, new_n6964_, new_n6965_,
    new_n6966_, new_n6967_, new_n6968_, new_n6969_, new_n6970_, new_n6971_,
    new_n6972_, new_n6973_, new_n6974_, new_n6975_, new_n6976_, new_n6977_,
    new_n6978_, new_n6979_, new_n6980_, new_n6981_, new_n6982_, new_n6983_,
    new_n6984_, new_n6985_, new_n6986_, new_n6987_, new_n6988_, new_n6989_,
    new_n6990_, new_n6991_, new_n6992_, new_n6993_, new_n6994_, new_n6995_,
    new_n6996_, new_n6997_, new_n6998_, new_n6999_, new_n7000_, new_n7001_,
    new_n7002_, new_n7003_, new_n7004_, new_n7005_, new_n7006_, new_n7007_,
    new_n7008_, new_n7009_, new_n7010_, new_n7011_, new_n7012_, new_n7013_,
    new_n7014_, new_n7015_, new_n7016_, new_n7017_, new_n7018_, new_n7019_,
    new_n7020_, new_n7021_, new_n7022_, new_n7023_, new_n7024_, new_n7025_,
    new_n7026_, new_n7027_, new_n7028_, new_n7029_, new_n7030_, new_n7031_,
    new_n7032_, new_n7033_, new_n7034_, new_n7035_, new_n7036_, new_n7037_,
    new_n7038_, new_n7039_, new_n7040_, new_n7041_, new_n7042_, new_n7043_,
    new_n7044_, new_n7045_, new_n7046_, new_n7047_, new_n7048_, new_n7049_,
    new_n7050_, new_n7051_, new_n7052_, new_n7053_, new_n7054_, new_n7055_,
    new_n7056_, new_n7057_, new_n7058_, new_n7059_, new_n7060_, new_n7061_,
    new_n7062_, new_n7063_, new_n7064_, new_n7065_, new_n7066_, new_n7067_,
    new_n7068_, new_n7069_, new_n7070_, new_n7071_, new_n7072_, new_n7073_,
    new_n7074_, new_n7075_, new_n7076_, new_n7077_, new_n7078_, new_n7079_,
    new_n7080_, new_n7081_, new_n7082_, new_n7083_, new_n7084_, new_n7085_,
    new_n7086_, new_n7087_, new_n7088_, new_n7089_, new_n7090_, new_n7091_,
    new_n7092_, new_n7093_, new_n7094_, new_n7095_, new_n7096_, new_n7097_,
    new_n7098_, new_n7099_, new_n7100_, new_n7101_, new_n7102_, new_n7103_,
    new_n7104_, new_n7105_, new_n7106_, new_n7107_, new_n7108_, new_n7109_,
    new_n7110_, new_n7111_, new_n7112_, new_n7113_, new_n7114_, new_n7115_,
    new_n7116_, new_n7117_, new_n7118_, new_n7119_, new_n7120_, new_n7121_,
    new_n7122_, new_n7123_, new_n7124_, new_n7125_, new_n7126_, new_n7127_,
    new_n7128_, new_n7129_, new_n7130_, new_n7131_, new_n7132_, new_n7133_,
    new_n7134_, new_n7135_, new_n7136_, new_n7137_, new_n7138_, new_n7139_,
    new_n7140_, new_n7141_, new_n7142_, new_n7143_, new_n7144_, new_n7145_,
    new_n7146_, new_n7147_, new_n7148_, new_n7149_, new_n7150_, new_n7151_,
    new_n7152_, new_n7153_, new_n7154_, new_n7155_, new_n7156_, new_n7157_,
    new_n7158_, new_n7159_, new_n7160_, new_n7161_, new_n7162_, new_n7163_,
    new_n7164_, new_n7165_, new_n7166_, new_n7167_, new_n7168_, new_n7169_,
    new_n7170_, new_n7171_, new_n7172_, new_n7173_, new_n7174_, new_n7175_,
    new_n7176_, new_n7177_, new_n7178_, new_n7179_, new_n7180_, new_n7181_,
    new_n7182_, new_n7183_, new_n7184_, new_n7185_, new_n7186_, new_n7187_,
    new_n7188_, new_n7189_, new_n7190_, new_n7191_, new_n7192_, new_n7193_,
    new_n7194_, new_n7195_, new_n7196_, new_n7197_, new_n7198_, new_n7199_,
    new_n7200_, new_n7201_, new_n7202_, new_n7203_, new_n7204_, new_n7205_,
    new_n7206_, new_n7207_, new_n7208_, new_n7209_, new_n7210_, new_n7211_,
    new_n7212_, new_n7213_, new_n7214_, new_n7215_, new_n7216_, new_n7217_,
    new_n7218_, new_n7219_, new_n7220_, new_n7221_, new_n7222_, new_n7223_,
    new_n7224_, new_n7225_, new_n7226_, new_n7227_, new_n7228_, new_n7229_,
    new_n7230_, new_n7231_, new_n7232_, new_n7233_, new_n7234_, new_n7235_,
    new_n7236_, new_n7237_, new_n7238_, new_n7239_, new_n7240_, new_n7241_,
    new_n7242_, new_n7243_, new_n7244_, new_n7245_, new_n7246_, new_n7247_,
    new_n7248_, new_n7249_, new_n7250_, new_n7251_, new_n7252_, new_n7253_,
    new_n7254_, new_n7255_, new_n7256_, new_n7257_, new_n7258_, new_n7259_,
    new_n7260_, new_n7261_, new_n7262_, new_n7263_, new_n7264_, new_n7265_,
    new_n7266_, new_n7267_, new_n7268_, new_n7269_, new_n7270_, new_n7271_,
    new_n7272_, new_n7273_, new_n7274_, new_n7275_, new_n7276_, new_n7277_,
    new_n7278_, new_n7279_, new_n7280_, new_n7281_, new_n7282_, new_n7283_,
    new_n7284_, new_n7285_, new_n7286_, new_n7287_, new_n7288_, new_n7289_,
    new_n7290_, new_n7291_, new_n7292_, new_n7293_, new_n7294_, new_n7295_,
    new_n7296_, new_n7297_, new_n7298_, new_n7299_, new_n7300_, new_n7301_,
    new_n7302_, new_n7303_, new_n7304_, new_n7305_, new_n7306_, new_n7307_,
    new_n7308_, new_n7309_, new_n7310_, new_n7311_, new_n7312_, new_n7313_,
    new_n7314_, new_n7315_, new_n7316_, new_n7317_, new_n7318_, new_n7319_,
    new_n7320_, new_n7321_, new_n7322_, new_n7323_, new_n7324_, new_n7325_,
    new_n7326_, new_n7327_, new_n7328_, new_n7329_, new_n7330_, new_n7331_,
    new_n7332_, new_n7333_, new_n7334_, new_n7335_, new_n7336_, new_n7337_,
    new_n7338_, new_n7339_, new_n7340_, new_n7341_, new_n7342_, new_n7343_,
    new_n7344_, new_n7345_, new_n7346_, new_n7347_, new_n7348_, new_n7349_,
    new_n7350_, new_n7351_, new_n7352_, new_n7353_, new_n7354_, new_n7355_,
    new_n7356_, new_n7357_, new_n7358_, new_n7359_, new_n7360_, new_n7361_,
    new_n7362_, new_n7363_, new_n7364_, new_n7365_, new_n7366_, new_n7367_,
    new_n7368_, new_n7369_, new_n7370_, new_n7371_, new_n7372_, new_n7373_,
    new_n7374_, new_n7375_, new_n7376_, new_n7377_, new_n7378_, new_n7379_,
    new_n7380_, new_n7381_, new_n7382_, new_n7383_, new_n7384_, new_n7385_,
    new_n7386_, new_n7387_, new_n7388_, new_n7389_, new_n7390_, new_n7391_,
    new_n7392_, new_n7393_, new_n7394_, new_n7395_, new_n7396_, new_n7397_,
    new_n7398_, new_n7399_, new_n7400_, new_n7401_, new_n7402_, new_n7403_,
    new_n7404_, new_n7405_, new_n7406_, new_n7407_, new_n7408_, new_n7409_,
    new_n7410_, new_n7411_, new_n7412_, new_n7413_, new_n7414_, new_n7415_,
    new_n7416_, new_n7417_, new_n7418_, new_n7419_, new_n7420_, new_n7421_,
    new_n7422_, new_n7423_, new_n7424_, new_n7425_, new_n7426_, new_n7427_,
    new_n7428_, new_n7429_, new_n7430_, new_n7431_, new_n7432_, new_n7433_,
    new_n7434_, new_n7435_, new_n7436_, new_n7437_, new_n7438_, new_n7439_,
    new_n7440_, new_n7441_, new_n7442_, new_n7443_, new_n7444_, new_n7445_,
    new_n7446_, new_n7447_, new_n7448_, new_n7449_, new_n7450_, new_n7451_,
    new_n7452_, new_n7453_, new_n7454_, new_n7455_, new_n7456_, new_n7457_,
    new_n7458_, new_n7459_, new_n7460_, new_n7461_, new_n7462_, new_n7463_,
    new_n7464_, new_n7465_, new_n7466_, new_n7467_, new_n7468_, new_n7469_,
    new_n7470_, new_n7471_, new_n7472_, new_n7473_, new_n7474_, new_n7475_,
    new_n7476_, new_n7477_, new_n7478_, new_n7479_, new_n7480_, new_n7481_,
    new_n7482_, new_n7483_, new_n7484_, new_n7485_, new_n7486_, new_n7487_,
    new_n7488_, new_n7489_, new_n7490_, new_n7491_, new_n7492_, new_n7493_,
    new_n7494_, new_n7495_, new_n7496_, new_n7497_, new_n7498_, new_n7499_,
    new_n7500_, new_n7501_, new_n7502_, new_n7503_, new_n7504_, new_n7505_,
    new_n7506_, new_n7507_, new_n7508_, new_n7509_, new_n7510_, new_n7511_,
    new_n7512_, new_n7513_, new_n7514_, new_n7515_, new_n7516_, new_n7517_,
    new_n7518_, new_n7519_, new_n7520_, new_n7521_, new_n7522_, new_n7523_,
    new_n7524_, new_n7525_, new_n7526_, new_n7527_, new_n7528_, new_n7529_,
    new_n7530_, new_n7531_, new_n7532_, new_n7533_, new_n7534_, new_n7535_,
    new_n7536_, new_n7537_, new_n7538_, new_n7539_, new_n7540_, new_n7541_,
    new_n7542_, new_n7543_, new_n7544_, new_n7545_, new_n7546_, new_n7547_,
    new_n7548_, new_n7549_, new_n7550_, new_n7551_, new_n7552_, new_n7553_,
    new_n7554_, new_n7555_, new_n7556_, new_n7557_, new_n7558_, new_n7559_,
    new_n7560_, new_n7561_, new_n7562_, new_n7563_, new_n7564_, new_n7565_,
    new_n7566_, new_n7567_, new_n7568_, new_n7569_, new_n7570_, new_n7571_,
    new_n7572_, new_n7573_, new_n7574_, new_n7575_, new_n7576_, new_n7577_,
    new_n7578_, new_n7579_, new_n7580_, new_n7581_, new_n7582_, new_n7583_,
    new_n7584_, new_n7585_, new_n7586_, new_n7587_, new_n7588_, new_n7589_,
    new_n7590_, new_n7591_, new_n7592_, new_n7593_, new_n7594_, new_n7595_,
    new_n7596_, new_n7597_, new_n7598_, new_n7599_, new_n7600_, new_n7601_,
    new_n7602_, new_n7603_, new_n7604_, new_n7605_, new_n7606_, new_n7607_,
    new_n7608_, new_n7609_, new_n7610_, new_n7611_, new_n7612_, new_n7613_,
    new_n7614_, new_n7615_, new_n7616_, new_n7617_, new_n7618_, new_n7619_,
    new_n7620_, new_n7621_, new_n7622_, new_n7623_, new_n7624_, new_n7625_,
    new_n7626_, new_n7627_, new_n7628_, new_n7629_, new_n7630_, new_n7631_,
    new_n7632_, new_n7633_, new_n7634_, new_n7635_, new_n7636_, new_n7637_,
    new_n7638_, new_n7639_, new_n7640_, new_n7641_, new_n7642_, new_n7643_,
    new_n7644_, new_n7645_, new_n7646_, new_n7647_, new_n7648_, new_n7649_,
    new_n7650_, new_n7651_, new_n7652_, new_n7653_, new_n7654_, new_n7655_,
    new_n7656_, new_n7657_, new_n7658_, new_n7659_, new_n7660_, new_n7661_,
    new_n7662_, new_n7663_, new_n7664_, new_n7665_, new_n7666_, new_n7667_,
    new_n7668_, new_n7669_, new_n7670_, new_n7671_, new_n7672_, new_n7673_,
    new_n7674_, new_n7675_, new_n7676_, new_n7677_, new_n7678_, new_n7679_,
    new_n7680_, new_n7681_, new_n7682_, new_n7683_, new_n7684_, new_n7685_,
    new_n7686_, new_n7687_, new_n7688_, new_n7689_, new_n7690_, new_n7691_,
    new_n7692_, new_n7693_, new_n7694_, new_n7695_, new_n7696_, new_n7697_,
    new_n7698_, new_n7699_, new_n7700_, new_n7701_, new_n7702_, new_n7703_,
    new_n7704_, new_n7705_, new_n7706_, new_n7707_, new_n7708_, new_n7709_,
    new_n7710_, new_n7711_, new_n7712_, new_n7713_, new_n7714_, new_n7715_,
    new_n7716_, new_n7717_, new_n7718_, new_n7719_, new_n7720_, new_n7721_,
    new_n7722_, new_n7723_, new_n7724_, new_n7725_, new_n7726_, new_n7727_,
    new_n7728_, new_n7729_, new_n7730_, new_n7731_, new_n7732_, new_n7733_,
    new_n7734_, new_n7735_, new_n7736_, new_n7737_, new_n7738_, new_n7739_,
    new_n7740_, new_n7741_, new_n7742_, new_n7743_, new_n7744_, new_n7745_,
    new_n7746_, new_n7747_, new_n7748_, new_n7749_, new_n7750_, new_n7751_,
    new_n7752_, new_n7753_, new_n7754_, new_n7755_, new_n7756_, new_n7757_,
    new_n7758_, new_n7759_, new_n7760_, new_n7761_, new_n7762_, new_n7763_,
    new_n7764_, new_n7765_, new_n7766_, new_n7767_, new_n7768_, new_n7769_,
    new_n7770_, new_n7771_, new_n7772_, new_n7773_, new_n7774_, new_n7775_,
    new_n7776_, new_n7777_, new_n7778_, new_n7779_, new_n7780_, new_n7781_,
    new_n7782_, new_n7783_, new_n7784_, new_n7785_, new_n7786_, new_n7787_,
    new_n7788_, new_n7789_, new_n7790_, new_n7791_, new_n7792_, new_n7793_,
    new_n7794_, new_n7795_, new_n7796_, new_n7797_, new_n7798_, new_n7799_,
    new_n7800_, new_n7801_, new_n7802_, new_n7803_, new_n7804_, new_n7805_,
    new_n7806_, new_n7807_, new_n7808_, new_n7809_, new_n7810_, new_n7811_,
    new_n7812_, new_n7813_, new_n7814_, new_n7815_, new_n7816_, new_n7817_,
    new_n7818_, new_n7819_, new_n7820_, new_n7821_, new_n7822_, new_n7823_,
    new_n7824_, new_n7825_, new_n7826_, new_n7827_, new_n7828_, new_n7829_,
    new_n7830_, new_n7831_, new_n7832_, new_n7833_, new_n7834_, new_n7835_,
    new_n7836_, new_n7837_, new_n7838_, new_n7839_, new_n7840_, new_n7841_,
    new_n7842_, new_n7843_, new_n7844_, new_n7845_, new_n7846_, new_n7847_,
    new_n7848_, new_n7849_, new_n7850_, new_n7851_, new_n7852_, new_n7853_,
    new_n7854_, new_n7855_, new_n7856_, new_n7857_, new_n7858_, new_n7859_,
    new_n7860_, new_n7861_, new_n7862_, new_n7863_, new_n7864_, new_n7865_,
    new_n7866_, new_n7867_, new_n7868_, new_n7869_, new_n7870_, new_n7871_,
    new_n7872_, new_n7873_, new_n7874_, new_n7875_, new_n7876_, new_n7877_,
    new_n7878_, new_n7879_, new_n7880_, new_n7881_, new_n7882_, new_n7883_,
    new_n7884_, new_n7885_, new_n7886_, new_n7887_, new_n7888_, new_n7889_,
    new_n7890_, new_n7891_, new_n7892_, new_n7893_, new_n7894_, new_n7895_,
    new_n7896_, new_n7897_, new_n7898_, new_n7899_, new_n7900_, new_n7901_,
    new_n7902_, new_n7903_, new_n7904_, new_n7905_, new_n7906_, new_n7907_,
    new_n7908_, new_n7909_, new_n7910_, new_n7911_, new_n7912_, new_n7913_,
    new_n7914_, new_n7915_, new_n7916_, new_n7917_, new_n7918_, new_n7919_,
    new_n7920_, new_n7921_, new_n7922_, new_n7923_, new_n7924_, new_n7925_,
    new_n7926_, new_n7927_, new_n7928_, new_n7929_, new_n7930_, new_n7931_,
    new_n7932_, new_n7933_, new_n7934_, new_n7935_, new_n7936_, new_n7937_,
    new_n7938_, new_n7939_, new_n7940_, new_n7941_, new_n7942_, new_n7943_,
    new_n7944_, new_n7945_, new_n7946_, new_n7947_, new_n7948_, new_n7949_,
    new_n7950_, new_n7951_, new_n7952_, new_n7953_, new_n7954_, new_n7955_,
    new_n7956_, new_n7957_, new_n7958_, new_n7959_, new_n7960_, new_n7961_,
    new_n7962_, new_n7963_, new_n7964_, new_n7965_, new_n7966_, new_n7967_,
    new_n7968_, new_n7969_, new_n7970_, new_n7971_, new_n7972_, new_n7973_,
    new_n7974_, new_n7975_, new_n7976_, new_n7977_, new_n7978_, new_n7979_,
    new_n7980_, new_n7981_, new_n7982_, new_n7983_, new_n7984_, new_n7985_,
    new_n7986_, new_n7987_, new_n7988_, new_n7989_, new_n7990_, new_n7991_,
    new_n7992_, new_n7993_, new_n7994_, new_n7995_, new_n7996_, new_n7997_,
    new_n7998_, new_n7999_, new_n8000_, new_n8001_, new_n8002_, new_n8003_,
    new_n8004_, new_n8005_, new_n8006_, new_n8007_, new_n8008_, new_n8009_,
    new_n8010_, new_n8011_, new_n8012_, new_n8013_, new_n8014_, new_n8015_,
    new_n8016_, new_n8017_, new_n8018_, new_n8019_, new_n8020_, new_n8021_,
    new_n8022_, new_n8023_, new_n8024_, new_n8025_, new_n8026_, new_n8027_,
    new_n8028_, new_n8029_, new_n8030_, new_n8031_, new_n8032_, new_n8033_,
    new_n8034_, new_n8035_, new_n8036_, new_n8037_, new_n8038_, new_n8039_,
    new_n8040_, new_n8041_, new_n8042_, new_n8043_, new_n8044_, new_n8045_,
    new_n8046_, new_n8047_, new_n8048_, new_n8049_, new_n8050_, new_n8051_,
    new_n8052_, new_n8053_, new_n8054_, new_n8055_, new_n8056_, new_n8057_,
    new_n8058_, new_n8059_, new_n8060_, new_n8061_, new_n8062_, new_n8063_,
    new_n8064_, new_n8065_, new_n8066_, new_n8067_, new_n8068_, new_n8069_,
    new_n8070_, new_n8071_, new_n8072_, new_n8073_, new_n8074_, new_n8075_,
    new_n8076_, new_n8077_, new_n8078_, new_n8079_, new_n8080_, new_n8081_,
    new_n8082_, new_n8083_, new_n8084_, new_n8085_, new_n8086_, new_n8087_,
    new_n8088_, new_n8089_, new_n8090_, new_n8091_, new_n8092_, new_n8093_,
    new_n8094_, new_n8095_, new_n8096_, new_n8097_, new_n8098_, new_n8099_,
    new_n8100_, new_n8101_, new_n8102_, new_n8103_, new_n8104_, new_n8105_,
    new_n8106_, new_n8107_, new_n8108_, new_n8109_, new_n8110_, new_n8111_,
    new_n8112_, new_n8113_, new_n8114_, new_n8115_, new_n8116_, new_n8117_,
    new_n8118_, new_n8119_, new_n8120_, new_n8121_, new_n8122_, new_n8123_,
    new_n8124_, new_n8125_, new_n8126_, new_n8127_, new_n8128_, new_n8129_,
    new_n8130_, new_n8131_, new_n8132_, new_n8133_, new_n8134_, new_n8135_,
    new_n8136_, new_n8137_, new_n8138_, new_n8139_, new_n8140_, new_n8141_,
    new_n8142_, new_n8143_, new_n8144_, new_n8145_, new_n8146_, new_n8147_,
    new_n8148_, new_n8149_, new_n8150_, new_n8151_, new_n8152_, new_n8153_,
    new_n8154_, new_n8155_, new_n8156_, new_n8157_, new_n8158_, new_n8159_,
    new_n8160_, new_n8161_, new_n8162_, new_n8163_, new_n8164_, new_n8165_,
    new_n8166_, new_n8167_, new_n8168_, new_n8169_, new_n8170_, new_n8171_,
    new_n8172_, new_n8173_, new_n8174_, new_n8175_, new_n8176_, new_n8177_,
    new_n8178_, new_n8179_, new_n8180_, new_n8181_, new_n8182_, new_n8183_,
    new_n8184_, new_n8185_, new_n8186_, new_n8187_, new_n8188_, new_n8189_,
    new_n8190_, new_n8191_, new_n8192_, new_n8193_, new_n8194_, new_n8195_,
    new_n8196_, new_n8197_, new_n8198_, new_n8199_, new_n8200_, new_n8201_,
    new_n8202_, new_n8203_, new_n8204_, new_n8205_, new_n8206_, new_n8207_,
    new_n8208_, new_n8209_, new_n8210_, new_n8211_, new_n8212_, new_n8213_,
    new_n8214_, new_n8215_, new_n8216_, new_n8217_, new_n8218_, new_n8219_,
    new_n8220_, new_n8221_, new_n8222_, new_n8223_, new_n8224_, new_n8225_,
    new_n8226_, new_n8227_, new_n8228_, new_n8229_, new_n8230_, new_n8231_,
    new_n8232_, new_n8233_, new_n8234_, new_n8235_, new_n8236_, new_n8237_,
    new_n8238_, new_n8239_, new_n8240_, new_n8241_, new_n8242_, new_n8243_,
    new_n8244_, new_n8245_, new_n8246_, new_n8247_, new_n8248_, new_n8249_,
    new_n8250_, new_n8251_, new_n8252_, new_n8253_, new_n8254_, new_n8255_,
    new_n8256_, new_n8257_, new_n8258_, new_n8259_, new_n8260_, new_n8261_,
    new_n8262_, new_n8263_, new_n8264_, new_n8265_, new_n8266_, new_n8267_,
    new_n8268_, new_n8269_, new_n8270_, new_n8271_, new_n8272_, new_n8273_,
    new_n8274_, new_n8275_, new_n8276_, new_n8277_, new_n8278_, new_n8279_,
    new_n8280_, new_n8281_, new_n8282_, new_n8283_, new_n8284_, new_n8285_,
    new_n8286_, new_n8287_, new_n8288_, new_n8289_, new_n8290_, new_n8291_,
    new_n8292_, new_n8293_, new_n8294_, new_n8295_, new_n8296_, new_n8297_,
    new_n8298_, new_n8299_, new_n8300_, new_n8301_, new_n8302_, new_n8303_,
    new_n8304_, new_n8305_, new_n8306_, new_n8307_, new_n8308_, new_n8309_,
    new_n8310_, new_n8311_, new_n8312_, new_n8313_, new_n8314_, new_n8315_,
    new_n8316_, new_n8317_, new_n8318_, new_n8319_, new_n8320_, new_n8321_,
    new_n8322_, new_n8323_, new_n8324_, new_n8325_, new_n8326_, new_n8327_,
    new_n8328_, new_n8329_, new_n8330_, new_n8331_, new_n8332_, new_n8333_,
    new_n8334_, new_n8335_, new_n8336_, new_n8337_, new_n8338_, new_n8339_,
    new_n8340_, new_n8341_, new_n8342_, new_n8343_, new_n8344_, new_n8345_,
    new_n8346_, new_n8347_, new_n8348_, new_n8349_, new_n8350_, new_n8351_,
    new_n8352_, new_n8353_, new_n8354_, new_n8355_, new_n8356_, new_n8357_,
    new_n8358_, new_n8359_, new_n8360_, new_n8361_, new_n8362_, new_n8363_,
    new_n8364_, new_n8365_, new_n8366_, new_n8367_, new_n8368_, new_n8369_,
    new_n8370_, new_n8371_, new_n8372_, new_n8373_, new_n8374_, new_n8375_,
    new_n8376_, new_n8377_, new_n8378_, new_n8379_, new_n8380_, new_n8381_,
    new_n8382_, new_n8383_, new_n8384_, new_n8385_, new_n8386_, new_n8387_,
    new_n8388_, new_n8389_, new_n8390_, new_n8391_, new_n8392_, new_n8393_,
    new_n8394_, new_n8395_, new_n8396_, new_n8397_, new_n8398_, new_n8399_,
    new_n8400_, new_n8401_, new_n8402_, new_n8403_, new_n8404_, new_n8405_,
    new_n8406_, new_n8407_, new_n8408_, new_n8409_, new_n8410_, new_n8411_,
    new_n8412_, new_n8413_, new_n8414_, new_n8415_, new_n8416_, new_n8417_,
    new_n8418_, new_n8419_, new_n8420_, new_n8421_, new_n8422_, new_n8423_,
    new_n8424_, new_n8425_, new_n8426_, new_n8427_, new_n8428_, new_n8429_,
    new_n8430_, new_n8431_, new_n8432_, new_n8433_, new_n8434_, new_n8435_,
    new_n8436_, new_n8437_, new_n8438_, new_n8439_, new_n8440_, new_n8441_,
    new_n8442_, new_n8443_, new_n8444_, new_n8445_, new_n8446_, new_n8447_,
    new_n8448_, new_n8449_, new_n8450_, new_n8451_, new_n8452_, new_n8453_,
    new_n8454_, new_n8455_, new_n8456_, new_n8457_, new_n8458_, new_n8459_,
    new_n8460_, new_n8461_, new_n8462_, new_n8463_, new_n8464_, new_n8465_,
    new_n8466_, new_n8467_, new_n8468_, new_n8469_, new_n8470_, new_n8471_,
    new_n8472_, new_n8473_, new_n8474_, new_n8475_, new_n8476_, new_n8477_,
    new_n8478_, new_n8479_, new_n8480_, new_n8481_, new_n8482_, new_n8483_,
    new_n8484_, new_n8485_, new_n8486_, new_n8487_, new_n8488_, new_n8489_,
    new_n8490_, new_n8491_, new_n8492_, new_n8493_, new_n8494_, new_n8495_,
    new_n8496_, new_n8497_, new_n8498_, new_n8499_, new_n8500_, new_n8501_,
    new_n8502_, new_n8503_, new_n8504_, new_n8505_, new_n8506_, new_n8507_,
    new_n8508_, new_n8509_, new_n8510_, new_n8511_, new_n8512_, new_n8513_,
    new_n8514_, new_n8515_, new_n8516_, new_n8517_, new_n8518_, new_n8519_,
    new_n8520_, new_n8521_, new_n8522_, new_n8523_, new_n8524_, new_n8525_,
    new_n8526_, new_n8527_, new_n8528_, new_n8529_, new_n8530_, new_n8531_,
    new_n8532_, new_n8533_, new_n8534_, new_n8535_, new_n8536_, new_n8537_,
    new_n8538_, new_n8539_, new_n8540_, new_n8541_, new_n8542_, new_n8543_,
    new_n8544_, new_n8545_, new_n8546_, new_n8547_, new_n8548_, new_n8549_,
    new_n8550_, new_n8551_, new_n8552_, new_n8553_, new_n8554_, new_n8555_,
    new_n8556_, new_n8557_, new_n8558_, new_n8559_, new_n8560_, new_n8561_,
    new_n8562_, new_n8563_, new_n8564_, new_n8565_, new_n8566_, new_n8567_,
    new_n8568_, new_n8569_, new_n8570_, new_n8571_, new_n8572_, new_n8573_,
    new_n8574_, new_n8575_, new_n8576_, new_n8577_, new_n8578_, new_n8579_,
    new_n8580_, new_n8581_, new_n8582_, new_n8583_, new_n8584_, new_n8585_,
    new_n8586_, new_n8587_, new_n8588_, new_n8589_, new_n8590_, new_n8591_,
    new_n8592_, new_n8593_, new_n8594_, new_n8595_, new_n8596_, new_n8597_,
    new_n8598_, new_n8599_, new_n8600_, new_n8601_, new_n8602_, new_n8603_,
    new_n8604_, new_n8605_, new_n8606_, new_n8607_, new_n8608_, new_n8609_,
    new_n8610_, new_n8611_, new_n8612_, new_n8613_, new_n8614_, new_n8615_,
    new_n8616_, new_n8617_, new_n8618_, new_n8619_, new_n8620_, new_n8621_,
    new_n8622_, new_n8623_, new_n8624_, new_n8625_, new_n8626_, new_n8627_,
    new_n8628_, new_n8629_, new_n8630_, new_n8631_, new_n8632_, new_n8633_,
    new_n8634_, new_n8635_, new_n8636_, new_n8637_, new_n8638_, new_n8639_,
    new_n8640_, new_n8641_, new_n8642_, new_n8643_, new_n8644_, new_n8645_,
    new_n8646_, new_n8647_, new_n8648_, new_n8649_, new_n8650_, new_n8651_,
    new_n8652_, new_n8653_, new_n8654_, new_n8655_, new_n8656_, new_n8657_,
    new_n8658_, new_n8659_, new_n8660_, new_n8661_, new_n8662_, new_n8663_,
    new_n8664_, new_n8665_, new_n8666_, new_n8667_, new_n8668_, new_n8669_,
    new_n8670_, new_n8671_, new_n8672_, new_n8673_, new_n8674_, new_n8675_,
    new_n8676_, new_n8677_, new_n8678_, new_n8679_, new_n8680_, new_n8681_,
    new_n8682_, new_n8683_, new_n8684_, new_n8685_, new_n8686_, new_n8687_,
    new_n8688_, new_n8689_, new_n8690_, new_n8691_, new_n8692_, new_n8693_,
    new_n8694_, new_n8695_, new_n8696_, new_n8697_, new_n8698_, new_n8699_,
    new_n8700_, new_n8701_, new_n8702_, new_n8703_, new_n8704_, new_n8705_,
    new_n8706_, new_n8707_, new_n8708_, new_n8709_, new_n8710_, new_n8711_,
    new_n8712_, new_n8713_, new_n8714_, new_n8715_, new_n8716_, new_n8717_,
    new_n8718_, new_n8719_, new_n8720_, new_n8721_, new_n8722_, new_n8723_,
    new_n8724_, new_n8725_, new_n8726_, new_n8727_, new_n8728_, new_n8729_,
    new_n8730_, new_n8731_, new_n8732_, new_n8733_, new_n8734_, new_n8735_,
    new_n8736_, new_n8737_, new_n8738_, new_n8739_, new_n8740_, new_n8741_,
    new_n8742_, new_n8743_, new_n8744_, new_n8745_, new_n8746_, new_n8747_,
    new_n8748_, new_n8749_, new_n8750_, new_n8751_, new_n8752_, new_n8753_,
    new_n8754_, new_n8755_, new_n8756_, new_n8757_, new_n8758_, new_n8759_,
    new_n8760_, new_n8761_, new_n8762_, new_n8763_, new_n8764_, new_n8765_,
    new_n8766_, new_n8767_, new_n8768_, new_n8769_, new_n8770_, new_n8771_,
    new_n8772_, new_n8773_, new_n8774_, new_n8775_, new_n8776_, new_n8777_,
    new_n8778_, new_n8779_, new_n8780_, new_n8781_, new_n8782_, new_n8783_,
    new_n8784_, new_n8785_, new_n8786_, new_n8787_, new_n8788_, new_n8789_,
    new_n8790_, new_n8791_, new_n8792_, new_n8793_, new_n8794_, new_n8795_,
    new_n8796_, new_n8797_, new_n8798_, new_n8799_, new_n8800_, new_n8801_,
    new_n8802_, new_n8803_, new_n8804_, new_n8805_, new_n8806_, new_n8807_,
    new_n8808_, new_n8809_, new_n8810_, new_n8811_, new_n8812_, new_n8813_,
    new_n8814_, new_n8815_, new_n8816_, new_n8817_, new_n8818_, new_n8819_,
    new_n8820_, new_n8821_, new_n8822_, new_n8823_, new_n8824_, new_n8825_,
    new_n8826_, new_n8827_, new_n8828_, new_n8829_, new_n8830_, new_n8831_,
    new_n8832_, new_n8833_, new_n8834_, new_n8835_, new_n8836_, new_n8837_,
    new_n8838_, new_n8839_, new_n8840_, new_n8841_, new_n8842_, new_n8843_,
    new_n8844_, new_n8845_, new_n8846_, new_n8847_, new_n8848_, new_n8849_,
    new_n8850_, new_n8851_, new_n8852_, new_n8853_, new_n8854_, new_n8855_,
    new_n8856_, new_n8857_, new_n8858_, new_n8859_, new_n8860_, new_n8861_,
    new_n8862_, new_n8863_, new_n8864_, new_n8865_, new_n8866_, new_n8867_,
    new_n8868_, new_n8869_, new_n8870_, new_n8871_, new_n8872_, new_n8873_,
    new_n8874_, new_n8875_, new_n8876_, new_n8877_, new_n8878_, new_n8879_,
    new_n8880_, new_n8881_, new_n8882_, new_n8883_, new_n8884_, new_n8885_,
    new_n8886_, new_n8887_, new_n8888_, new_n8889_, new_n8890_, new_n8891_,
    new_n8892_, new_n8893_, new_n8894_, new_n8895_, new_n8896_, new_n8897_,
    new_n8898_, new_n8899_, new_n8900_, new_n8901_, new_n8902_, new_n8903_,
    new_n8904_, new_n8905_, new_n8906_, new_n8907_, new_n8908_, new_n8909_,
    new_n8910_, new_n8911_, new_n8912_, new_n8913_, new_n8914_, new_n8915_,
    new_n8916_, new_n8917_, new_n8918_, new_n8919_, new_n8920_, new_n8921_,
    new_n8922_, new_n8923_, new_n8924_, new_n8925_, new_n8926_, new_n8927_,
    new_n8928_, new_n8929_, new_n8930_, new_n8931_, new_n8932_, new_n8933_,
    new_n8934_, new_n8935_, new_n8936_, new_n8937_, new_n8938_, new_n8939_,
    new_n8940_, new_n8941_, new_n8942_, new_n8943_, new_n8944_, new_n8945_,
    new_n8946_, new_n8947_, new_n8948_, new_n8949_, new_n8950_, new_n8951_,
    new_n8952_, new_n8953_, new_n8954_, new_n8955_, new_n8956_, new_n8957_,
    new_n8958_, new_n8959_, new_n8960_, new_n8961_, new_n8962_, new_n8963_,
    new_n8964_, new_n8965_, new_n8966_, new_n8967_, new_n8968_, new_n8969_,
    new_n8970_, new_n8971_, new_n8972_, new_n8973_, new_n8974_, new_n8975_,
    new_n8976_, new_n8977_, new_n8978_, new_n8979_, new_n8980_, new_n8981_,
    new_n8982_, new_n8983_, new_n8984_, new_n8985_, new_n8986_, new_n8987_,
    new_n8988_, new_n8989_, new_n8990_, new_n8991_, new_n8992_, new_n8993_,
    new_n8994_, new_n8995_, new_n8996_, new_n8997_, new_n8998_, new_n8999_,
    new_n9000_, new_n9001_, new_n9002_, new_n9003_, new_n9004_, new_n9005_,
    new_n9006_, new_n9007_, new_n9008_, new_n9009_, new_n9010_, new_n9011_,
    new_n9012_, new_n9013_, new_n9014_, new_n9015_, new_n9016_, new_n9017_,
    new_n9018_, new_n9019_, new_n9020_, new_n9021_, new_n9022_, new_n9023_,
    new_n9024_, new_n9025_, new_n9026_, new_n9027_, new_n9028_, new_n9029_,
    new_n9030_, new_n9031_, new_n9032_, new_n9033_, new_n9034_, new_n9035_,
    new_n9036_, new_n9037_, new_n9038_, new_n9039_, new_n9040_, new_n9041_,
    new_n9042_, new_n9043_, new_n9044_, new_n9045_, new_n9046_, new_n9047_,
    new_n9048_, new_n9049_, new_n9050_, new_n9051_, new_n9052_, new_n9053_,
    new_n9054_, new_n9055_, new_n9056_, new_n9057_, new_n9058_, new_n9059_,
    new_n9060_, new_n9061_, new_n9062_, new_n9063_, new_n9064_, new_n9065_,
    new_n9066_, new_n9067_, new_n9068_, new_n9069_, new_n9070_, new_n9071_,
    new_n9072_, new_n9073_, new_n9074_, new_n9075_, new_n9076_, new_n9077_,
    new_n9078_, new_n9079_, new_n9080_, new_n9081_, new_n9082_, new_n9083_,
    new_n9084_, new_n9085_, new_n9086_, new_n9087_, new_n9088_, new_n9089_,
    new_n9090_, new_n9091_, new_n9092_, new_n9093_, new_n9094_, new_n9095_,
    new_n9096_, new_n9097_, new_n9098_, new_n9099_, new_n9100_, new_n9101_,
    new_n9102_, new_n9103_, new_n9104_, new_n9105_, new_n9106_, new_n9107_,
    new_n9108_, new_n9109_, new_n9110_, new_n9111_, new_n9112_, new_n9113_,
    new_n9114_, new_n9115_, new_n9116_, new_n9117_, new_n9118_, new_n9119_,
    new_n9120_, new_n9121_, new_n9122_, new_n9123_, new_n9124_, new_n9125_,
    new_n9126_, new_n9127_, new_n9128_, new_n9129_, new_n9130_, new_n9131_,
    new_n9132_, new_n9133_, new_n9134_, new_n9135_, new_n9136_, new_n9137_,
    new_n9138_, new_n9139_, new_n9140_, new_n9141_, new_n9142_, new_n9143_,
    new_n9144_, new_n9145_, new_n9146_, new_n9147_, new_n9148_, new_n9149_,
    new_n9150_, new_n9151_, new_n9152_, new_n9153_, new_n9154_, new_n9155_,
    new_n9156_, new_n9157_, new_n9158_, new_n9159_, new_n9160_, new_n9161_,
    new_n9162_, new_n9163_, new_n9164_, new_n9165_, new_n9166_, new_n9167_,
    new_n9168_, new_n9169_, new_n9170_, new_n9171_, new_n9172_, new_n9173_,
    new_n9174_, new_n9175_, new_n9176_, new_n9177_, new_n9178_, new_n9179_,
    new_n9180_, new_n9181_, new_n9182_, new_n9183_, new_n9184_, new_n9185_,
    new_n9186_, new_n9187_, new_n9188_, new_n9189_, new_n9190_, new_n9191_,
    new_n9192_, new_n9193_, new_n9194_, new_n9195_, new_n9196_, new_n9197_,
    new_n9198_, new_n9199_, new_n9200_, new_n9201_, new_n9202_, new_n9203_,
    new_n9204_, new_n9205_, new_n9206_, new_n9207_, new_n9208_, new_n9209_,
    new_n9210_, new_n9211_, new_n9212_, new_n9213_, new_n9214_, new_n9215_,
    new_n9216_, new_n9217_, new_n9218_, new_n9219_, new_n9220_, new_n9221_,
    new_n9222_, new_n9223_, new_n9224_, new_n9225_, new_n9226_, new_n9227_,
    new_n9228_, new_n9229_, new_n9230_, new_n9231_, new_n9232_, new_n9233_,
    new_n9234_, new_n9235_, new_n9236_, new_n9237_, new_n9238_, new_n9239_,
    new_n9240_, new_n9241_, new_n9242_, new_n9243_, new_n9244_, new_n9245_,
    new_n9246_, new_n9247_, new_n9248_, new_n9249_, new_n9250_, new_n9251_,
    new_n9252_, new_n9253_, new_n9254_, new_n9255_, new_n9256_, new_n9257_,
    new_n9258_, new_n9259_, new_n9260_, new_n9261_, new_n9262_, new_n9263_,
    new_n9264_, new_n9265_, new_n9266_, new_n9267_, new_n9268_, new_n9269_,
    new_n9270_, new_n9271_, new_n9272_, new_n9273_, new_n9274_, new_n9275_,
    new_n9276_, new_n9277_, new_n9278_, new_n9279_, new_n9280_, new_n9281_,
    new_n9282_, new_n9283_, new_n9284_, new_n9285_, new_n9286_, new_n9287_,
    new_n9288_, new_n9289_, new_n9290_, new_n9291_, new_n9292_, new_n9293_,
    new_n9294_, new_n9295_, new_n9296_, new_n9297_, new_n9298_, new_n9299_,
    new_n9300_, new_n9301_, new_n9302_, new_n9303_, new_n9304_, new_n9305_,
    new_n9306_, new_n9307_, new_n9308_, new_n9309_, new_n9310_, new_n9311_,
    new_n9312_, new_n9313_, new_n9314_, new_n9315_, new_n9316_, new_n9317_,
    new_n9318_, new_n9319_, new_n9320_, new_n9321_, new_n9322_, new_n9323_,
    new_n9324_, new_n9325_, new_n9326_, new_n9327_, new_n9328_, new_n9329_,
    new_n9330_, new_n9331_, new_n9332_, new_n9333_, new_n9334_, new_n9335_,
    new_n9336_, new_n9337_, new_n9338_, new_n9339_, new_n9340_, new_n9341_,
    new_n9342_, new_n9343_, new_n9344_, new_n9345_, new_n9346_, new_n9347_,
    new_n9348_, new_n9349_, new_n9350_, new_n9351_, new_n9352_, new_n9353_,
    new_n9354_, new_n9355_, new_n9356_, new_n9357_, new_n9358_, new_n9359_,
    new_n9360_, new_n9361_, new_n9362_, new_n9363_, new_n9364_, new_n9365_,
    new_n9366_, new_n9367_, new_n9368_, new_n9369_, new_n9370_, new_n9371_,
    new_n9372_, new_n9373_, new_n9374_, new_n9375_, new_n9376_, new_n9377_,
    new_n9378_, new_n9379_, new_n9380_, new_n9381_, new_n9382_, new_n9383_,
    new_n9384_, new_n9385_, new_n9386_, new_n9387_, new_n9388_, new_n9389_,
    new_n9390_, new_n9391_, new_n9392_, new_n9393_, new_n9394_, new_n9395_,
    new_n9396_, new_n9397_, new_n9398_, new_n9399_, new_n9400_, new_n9401_,
    new_n9402_, new_n9403_, new_n9404_, new_n9405_, new_n9406_, new_n9407_,
    new_n9408_, new_n9409_, new_n9410_, new_n9411_, new_n9412_, new_n9413_,
    new_n9414_, new_n9415_, new_n9416_, new_n9417_, new_n9418_, new_n9419_,
    new_n9420_, new_n9421_, new_n9422_, new_n9423_, new_n9424_, new_n9425_,
    new_n9426_, new_n9427_, new_n9428_, new_n9429_, new_n9430_, new_n9431_,
    new_n9432_, new_n9433_, new_n9434_, new_n9435_, new_n9436_, new_n9437_,
    new_n9438_, new_n9439_, new_n9440_, new_n9441_, new_n9442_, new_n9443_,
    new_n9444_, new_n9445_, new_n9446_, new_n9447_, new_n9448_, new_n9449_,
    new_n9450_, new_n9451_, new_n9452_, new_n9453_, new_n9454_, new_n9455_,
    new_n9456_, new_n9457_, new_n9458_, new_n9459_, new_n9460_, new_n9461_,
    new_n9462_, new_n9463_, new_n9464_, new_n9465_, new_n9466_, new_n9467_,
    new_n9468_, new_n9469_, new_n9470_, new_n9471_, new_n9472_, new_n9473_,
    new_n9474_, new_n9475_, new_n9476_, new_n9477_, new_n9478_, new_n9479_,
    new_n9480_, new_n9481_, new_n9482_, new_n9483_, new_n9484_, new_n9485_,
    new_n9486_, new_n9487_, new_n9488_, new_n9489_, new_n9490_, new_n9491_,
    new_n9492_, new_n9493_, new_n9494_, new_n9495_, new_n9496_, new_n9497_,
    new_n9498_, new_n9499_, new_n9500_, new_n9501_, new_n9502_, new_n9503_,
    new_n9504_, new_n9505_, new_n9506_, new_n9507_, new_n9508_, new_n9509_,
    new_n9510_, new_n9511_, new_n9512_, new_n9513_, new_n9514_, new_n9515_,
    new_n9516_, new_n9517_, new_n9518_, new_n9519_, new_n9520_, new_n9521_,
    new_n9522_, new_n9523_, new_n9524_, new_n9525_, new_n9526_, new_n9527_,
    new_n9528_, new_n9529_, new_n9530_, new_n9531_, new_n9532_, new_n9533_,
    new_n9534_, new_n9535_, new_n9536_, new_n9537_, new_n9538_, new_n9539_,
    new_n9540_, new_n9541_, new_n9542_, new_n9543_, new_n9544_, new_n9545_,
    new_n9546_, new_n9547_, new_n9548_, new_n9549_, new_n9550_, new_n9551_,
    new_n9552_, new_n9553_, new_n9554_, new_n9555_, new_n9556_, new_n9557_,
    new_n9558_, new_n9559_, new_n9560_, new_n9561_, new_n9562_, new_n9563_,
    new_n9564_, new_n9565_, new_n9566_, new_n9567_, new_n9568_, new_n9569_,
    new_n9570_, new_n9571_, new_n9572_, new_n9573_, new_n9574_, new_n9575_,
    new_n9576_, new_n9577_, new_n9578_, new_n9579_, new_n9580_, new_n9581_,
    new_n9582_, new_n9583_, new_n9584_, new_n9585_, new_n9586_, new_n9587_,
    new_n9588_, new_n9589_, new_n9590_, new_n9591_, new_n9592_, new_n9593_,
    new_n9594_, new_n9595_, new_n9596_, new_n9597_, new_n9598_, new_n9599_,
    new_n9600_, new_n9601_, new_n9602_, new_n9603_, new_n9604_, new_n9605_,
    new_n9606_, new_n9607_, new_n9608_, new_n9609_, new_n9610_, new_n9611_,
    new_n9612_, new_n9613_, new_n9614_, new_n9615_, new_n9616_, new_n9617_,
    new_n9618_, new_n9619_, new_n9620_, new_n9621_, new_n9622_, new_n9623_,
    new_n9624_, new_n9625_, new_n9626_, new_n9627_, new_n9628_, new_n9629_,
    new_n9630_, new_n9631_, new_n9632_, new_n9633_, new_n9634_, new_n9635_,
    new_n9636_, new_n9637_, new_n9638_, new_n9639_, new_n9640_, new_n9641_,
    new_n9642_, new_n9643_, new_n9644_, new_n9645_, new_n9646_, new_n9647_,
    new_n9648_, new_n9649_, new_n9650_, new_n9651_, new_n9652_, new_n9653_,
    new_n9654_, new_n9655_, new_n9656_, new_n9657_, new_n9658_, new_n9659_,
    new_n9660_, new_n9661_, new_n9662_, new_n9663_, new_n9664_, new_n9665_,
    new_n9666_, new_n9667_, new_n9668_, new_n9669_, new_n9670_, new_n9671_,
    new_n9672_, new_n9673_, new_n9674_, new_n9675_, new_n9676_, new_n9677_,
    new_n9678_, new_n9679_, new_n9680_, new_n9681_, new_n9682_, new_n9683_,
    new_n9684_, new_n9685_, new_n9686_, new_n9687_, new_n9688_, new_n9689_,
    new_n9690_, new_n9691_, new_n9692_, new_n9693_, new_n9694_, new_n9695_,
    new_n9696_, new_n9697_, new_n9698_, new_n9699_, new_n9700_, new_n9701_,
    new_n9702_, new_n9703_, new_n9704_, new_n9705_, new_n9706_, new_n9707_,
    new_n9708_, new_n9709_, new_n9710_, new_n9711_, new_n9712_, new_n9713_,
    new_n9714_, new_n9715_, new_n9716_, new_n9717_, new_n9718_, new_n9719_,
    new_n9720_, new_n9721_, new_n9722_, new_n9723_, new_n9724_, new_n9725_,
    new_n9726_, new_n9727_, new_n9728_, new_n9729_, new_n9730_, new_n9731_,
    new_n9732_, new_n9733_, new_n9734_, new_n9735_, new_n9736_, new_n9737_,
    new_n9738_, new_n9739_, new_n9740_, new_n9741_, new_n9742_, new_n9743_,
    new_n9744_, new_n9745_, new_n9746_, new_n9747_, new_n9748_, new_n9749_,
    new_n9750_, new_n9751_, new_n9752_, new_n9753_, new_n9754_, new_n9755_,
    new_n9756_, new_n9757_, new_n9758_, new_n9759_, new_n9760_, new_n9761_,
    new_n9762_, new_n9763_, new_n9764_, new_n9765_, new_n9766_, new_n9767_,
    new_n9768_, new_n9769_, new_n9770_, new_n9771_, new_n9772_, new_n9773_,
    new_n9774_, new_n9775_, new_n9776_, new_n9777_, new_n9778_, new_n9779_,
    new_n9780_, new_n9781_, new_n9782_, new_n9783_, new_n9784_, new_n9785_,
    new_n9786_, new_n9787_, new_n9788_, new_n9789_, new_n9790_, new_n9791_,
    new_n9792_, new_n9793_, new_n9794_, new_n9795_, new_n9796_, new_n9797_,
    new_n9798_, new_n9799_, new_n9800_, new_n9801_, new_n9802_, new_n9803_,
    new_n9804_, new_n9805_, new_n9806_, new_n9807_, new_n9808_, new_n9809_,
    new_n9810_, new_n9811_, new_n9812_, new_n9813_, new_n9814_, new_n9815_,
    new_n9816_, new_n9817_, new_n9818_, new_n9819_, new_n9820_, new_n9821_,
    new_n9822_, new_n9823_, new_n9824_, new_n9825_, new_n9826_, new_n9827_,
    new_n9828_, new_n9829_, new_n9830_, new_n9831_, new_n9832_, new_n9833_,
    new_n9834_, new_n9835_, new_n9836_, new_n9837_, new_n9838_, new_n9839_,
    new_n9840_, new_n9841_, new_n9842_, new_n9843_, new_n9844_, new_n9845_,
    new_n9846_, new_n9847_, new_n9848_, new_n9849_, new_n9850_, new_n9851_,
    new_n9852_, new_n9853_, new_n9854_, new_n9855_, new_n9856_, new_n9857_,
    new_n9858_, new_n9859_, new_n9860_, new_n9861_, new_n9862_, new_n9863_,
    new_n9864_, new_n9865_, new_n9866_, new_n9867_, new_n9868_, new_n9869_,
    new_n9870_, new_n9871_, new_n9872_, new_n9873_, new_n9874_, new_n9875_,
    new_n9876_, new_n9877_, new_n9878_, new_n9879_, new_n9880_, new_n9881_,
    new_n9882_, new_n9883_, new_n9884_, new_n9885_, new_n9886_, new_n9887_,
    new_n9888_, new_n9889_, new_n9890_, new_n9891_, new_n9892_, new_n9893_,
    new_n9894_, new_n9895_, new_n9896_, new_n9897_, new_n9898_, new_n9899_,
    new_n9900_, new_n9901_, new_n9902_, new_n9903_, new_n9904_, new_n9905_,
    new_n9906_, new_n9907_, new_n9908_, new_n9909_, new_n9910_, new_n9911_,
    new_n9912_, new_n9913_, new_n9914_, new_n9915_, new_n9916_, new_n9917_,
    new_n9918_, new_n9919_, new_n9920_, new_n9921_, new_n9922_, new_n9923_,
    new_n9924_, new_n9925_, new_n9926_, new_n9927_, new_n9928_, new_n9929_,
    new_n9930_, new_n9931_, new_n9932_, new_n9933_, new_n9934_, new_n9935_,
    new_n9936_, new_n9937_, new_n9938_, new_n9939_, new_n9940_, new_n9941_,
    new_n9942_, new_n9943_, new_n9944_, new_n9945_, new_n9946_, new_n9947_,
    new_n9948_, new_n9949_, new_n9950_, new_n9951_, new_n9952_, new_n9953_,
    new_n9954_, new_n9955_, new_n9956_, new_n9957_, new_n9958_, new_n9959_,
    new_n9960_, new_n9961_, new_n9962_, new_n9963_, new_n9964_, new_n9965_,
    new_n9966_, new_n9967_, new_n9968_, new_n9969_, new_n9970_, new_n9971_,
    new_n9972_, new_n9973_, new_n9974_, new_n9975_, new_n9976_, new_n9977_,
    new_n9978_, new_n9979_, new_n9980_, new_n9981_, new_n9982_, new_n9983_,
    new_n9984_, new_n9985_, new_n9986_, new_n9987_, new_n9988_, new_n9989_,
    new_n9990_, new_n9991_, new_n9992_, new_n9993_, new_n9994_, new_n9995_,
    new_n9996_, new_n9997_, new_n9998_, new_n9999_, new_n10000_,
    new_n10001_, new_n10002_, new_n10003_, new_n10004_, new_n10005_,
    new_n10006_, new_n10007_, new_n10008_, new_n10009_, new_n10010_,
    new_n10011_, new_n10012_, new_n10013_, new_n10014_, new_n10015_,
    new_n10016_, new_n10017_, new_n10018_, new_n10019_, new_n10020_,
    new_n10021_, new_n10022_, new_n10023_, new_n10024_, new_n10025_,
    new_n10026_, new_n10027_, new_n10028_, new_n10029_, new_n10030_,
    new_n10031_, new_n10032_, new_n10033_, new_n10034_, new_n10035_,
    new_n10036_, new_n10037_, new_n10038_, new_n10039_, new_n10040_,
    new_n10041_, new_n10042_, new_n10043_, new_n10044_, new_n10045_,
    new_n10046_, new_n10047_, new_n10048_, new_n10049_, new_n10050_,
    new_n10051_, new_n10052_, new_n10053_, new_n10054_, new_n10055_,
    new_n10056_, new_n10057_, new_n10058_, new_n10059_, new_n10060_,
    new_n10061_, new_n10062_, new_n10063_, new_n10064_, new_n10065_,
    new_n10066_, new_n10067_, new_n10068_, new_n10069_, new_n10070_,
    new_n10071_, new_n10072_, new_n10073_, new_n10074_, new_n10075_,
    new_n10076_, new_n10077_, new_n10078_, new_n10079_, new_n10080_,
    new_n10081_, new_n10082_, new_n10083_, new_n10084_, new_n10085_,
    new_n10086_, new_n10087_, new_n10088_, new_n10089_, new_n10090_,
    new_n10091_, new_n10092_, new_n10093_, new_n10094_, new_n10095_,
    new_n10096_, new_n10097_, new_n10098_, new_n10099_, new_n10100_,
    new_n10101_, new_n10102_, new_n10103_, new_n10104_, new_n10105_,
    new_n10106_, new_n10107_, new_n10108_, new_n10109_, new_n10110_,
    new_n10111_, new_n10112_, new_n10113_, new_n10114_, new_n10115_,
    new_n10116_, new_n10117_, new_n10118_, new_n10119_, new_n10120_,
    new_n10121_, new_n10122_, new_n10123_, new_n10124_, new_n10125_,
    new_n10126_, new_n10127_, new_n10128_, new_n10129_, new_n10130_,
    new_n10131_, new_n10132_, new_n10133_, new_n10134_, new_n10135_,
    new_n10136_, new_n10137_, new_n10138_, new_n10139_, new_n10140_,
    new_n10141_, new_n10142_, new_n10143_, new_n10144_, new_n10145_,
    new_n10146_, new_n10147_, new_n10148_, new_n10149_, new_n10150_,
    new_n10151_, new_n10152_, new_n10153_, new_n10154_, new_n10155_,
    new_n10156_, new_n10157_, new_n10158_, new_n10159_, new_n10160_,
    new_n10161_, new_n10162_, new_n10163_, new_n10164_, new_n10165_,
    new_n10166_, new_n10167_, new_n10168_, new_n10169_, new_n10170_,
    new_n10171_, new_n10172_, new_n10173_, new_n10174_, new_n10175_,
    new_n10176_, new_n10177_, new_n10178_, new_n10179_, new_n10180_,
    new_n10181_, new_n10182_, new_n10183_, new_n10184_, new_n10185_,
    new_n10186_, new_n10187_, new_n10188_, new_n10189_, new_n10190_,
    new_n10191_, new_n10192_, new_n10193_, new_n10194_, new_n10195_,
    new_n10196_, new_n10197_, new_n10198_, new_n10199_, new_n10200_,
    new_n10201_, new_n10202_, new_n10203_, new_n10204_, new_n10205_,
    new_n10206_, new_n10207_, new_n10208_, new_n10209_, new_n10210_,
    new_n10211_, new_n10212_, new_n10213_, new_n10214_, new_n10215_,
    new_n10216_, new_n10217_, new_n10218_, new_n10219_, new_n10220_,
    new_n10221_, new_n10222_, new_n10223_, new_n10224_, new_n10225_,
    new_n10226_, new_n10227_, new_n10228_, new_n10229_, new_n10230_,
    new_n10231_, new_n10232_, new_n10233_, new_n10234_, new_n10235_,
    new_n10236_, new_n10237_, new_n10238_, new_n10239_, new_n10240_,
    new_n10241_, new_n10242_, new_n10243_, new_n10244_, new_n10245_,
    new_n10246_, new_n10247_, new_n10248_, new_n10249_, new_n10250_,
    new_n10251_, new_n10252_, new_n10253_, new_n10254_, new_n10255_,
    new_n10256_, new_n10257_, new_n10258_, new_n10259_, new_n10260_,
    new_n10261_, new_n10262_, new_n10263_, new_n10264_, new_n10265_,
    new_n10266_, new_n10267_, new_n10268_, new_n10269_, new_n10270_,
    new_n10271_, new_n10272_, new_n10273_, new_n10274_, new_n10275_,
    new_n10276_, new_n10277_, new_n10278_, new_n10279_, new_n10280_,
    new_n10281_, new_n10282_, new_n10283_, new_n10284_, new_n10285_,
    new_n10286_, new_n10287_, new_n10288_, new_n10289_, new_n10290_,
    new_n10291_, new_n10292_, new_n10293_, new_n10294_, new_n10295_,
    new_n10296_, new_n10297_, new_n10298_, new_n10299_, new_n10300_,
    new_n10301_, new_n10302_, new_n10303_, new_n10304_, new_n10305_,
    new_n10306_, new_n10307_, new_n10308_, new_n10309_, new_n10310_,
    new_n10311_, new_n10312_, new_n10313_, new_n10314_, new_n10315_,
    new_n10316_, new_n10317_, new_n10318_, new_n10319_, new_n10320_,
    new_n10321_, new_n10322_, new_n10323_, new_n10324_, new_n10325_,
    new_n10326_, new_n10327_, new_n10328_, new_n10329_, new_n10330_,
    new_n10331_, new_n10332_, new_n10333_, new_n10334_, new_n10335_,
    new_n10336_, new_n10337_, new_n10338_, new_n10339_, new_n10340_,
    new_n10341_, new_n10342_, new_n10343_, new_n10344_, new_n10345_,
    new_n10346_, new_n10347_, new_n10348_, new_n10349_, new_n10350_,
    new_n10351_, new_n10352_, new_n10353_, new_n10354_, new_n10355_,
    new_n10356_, new_n10357_, new_n10358_, new_n10359_, new_n10360_,
    new_n10361_, new_n10362_, new_n10363_, new_n10364_, new_n10365_,
    new_n10366_, new_n10367_, new_n10368_, new_n10369_, new_n10370_,
    new_n10371_, new_n10372_, new_n10373_, new_n10374_, new_n10375_,
    new_n10376_, new_n10377_, new_n10378_, new_n10379_, new_n10380_,
    new_n10381_, new_n10382_, new_n10383_, new_n10384_, new_n10385_,
    new_n10386_, new_n10387_, new_n10388_, new_n10389_, new_n10390_,
    new_n10391_, new_n10392_, new_n10393_, new_n10394_, new_n10395_,
    new_n10396_, new_n10397_, new_n10398_, new_n10399_, new_n10400_,
    new_n10401_, new_n10402_, new_n10403_, new_n10404_, new_n10405_,
    new_n10406_, new_n10407_, new_n10408_, new_n10409_, new_n10410_,
    new_n10411_, new_n10412_, new_n10413_, new_n10414_, new_n10415_,
    new_n10416_, new_n10417_, new_n10418_, new_n10419_, new_n10420_,
    new_n10421_, new_n10422_, new_n10423_, new_n10424_, new_n10425_,
    new_n10426_, new_n10427_, new_n10428_, new_n10429_, new_n10430_,
    new_n10431_, new_n10432_, new_n10433_, new_n10434_, new_n10435_,
    new_n10436_, new_n10437_, new_n10438_, new_n10439_, new_n10440_,
    new_n10441_, new_n10442_, new_n10443_, new_n10444_, new_n10445_,
    new_n10446_, new_n10447_, new_n10448_, new_n10449_, new_n10450_,
    new_n10451_, new_n10452_, new_n10453_, new_n10454_, new_n10455_,
    new_n10456_, new_n10457_, new_n10458_, new_n10459_, new_n10460_,
    new_n10461_, new_n10462_, new_n10463_, new_n10464_, new_n10465_,
    new_n10466_, new_n10467_, new_n10468_, new_n10469_, new_n10470_,
    new_n10471_, new_n10472_, new_n10473_, new_n10474_, new_n10475_,
    new_n10476_, new_n10477_, new_n10478_, new_n10479_, new_n10480_,
    new_n10481_, new_n10482_, new_n10483_, new_n10484_, new_n10485_,
    new_n10486_, new_n10487_, new_n10488_, new_n10489_, new_n10490_,
    new_n10491_, new_n10492_, new_n10493_, new_n10494_, new_n10495_,
    new_n10496_, new_n10497_, new_n10498_, new_n10499_, new_n10500_,
    new_n10501_, new_n10502_, new_n10503_, new_n10504_, new_n10505_,
    new_n10506_, new_n10507_, new_n10508_, new_n10509_, new_n10510_,
    new_n10511_, new_n10512_, new_n10513_, new_n10514_, new_n10515_,
    new_n10516_, new_n10517_, new_n10518_, new_n10519_, new_n10520_,
    new_n10521_, new_n10522_, new_n10523_, new_n10524_, new_n10525_,
    new_n10526_, new_n10527_, new_n10528_, new_n10529_, new_n10530_,
    new_n10531_, new_n10532_, new_n10533_, new_n10534_, new_n10535_,
    new_n10536_, new_n10537_, new_n10538_, new_n10539_, new_n10540_,
    new_n10541_, new_n10542_, new_n10543_, new_n10544_, new_n10545_,
    new_n10546_, new_n10547_, new_n10548_, new_n10549_, new_n10550_,
    new_n10551_, new_n10552_, new_n10553_, new_n10554_, new_n10555_,
    new_n10556_, new_n10557_, new_n10558_, new_n10559_, new_n10560_,
    new_n10561_, new_n10562_, new_n10563_, new_n10564_, new_n10565_,
    new_n10566_, new_n10567_, new_n10568_, new_n10569_, new_n10570_,
    new_n10571_, new_n10572_, new_n10573_, new_n10574_, new_n10575_,
    new_n10576_, new_n10577_, new_n10578_, new_n10579_, new_n10580_,
    new_n10581_, new_n10582_, new_n10583_, new_n10584_, new_n10585_,
    new_n10586_, new_n10587_, new_n10588_, new_n10589_, new_n10590_,
    new_n10591_, new_n10592_, new_n10593_, new_n10594_, new_n10595_,
    new_n10596_, new_n10597_, new_n10598_, new_n10599_, new_n10600_,
    new_n10601_, new_n10602_, new_n10603_, new_n10604_, new_n10605_,
    new_n10606_, new_n10607_, new_n10608_, new_n10609_, new_n10610_,
    new_n10611_, new_n10612_, new_n10613_, new_n10614_, new_n10615_,
    new_n10616_, new_n10617_, new_n10618_, new_n10619_, new_n10620_,
    new_n10621_, new_n10622_, new_n10623_, new_n10624_, new_n10625_,
    new_n10626_, new_n10627_, new_n10628_, new_n10629_, new_n10630_,
    new_n10631_, new_n10632_, new_n10633_, new_n10634_, new_n10635_,
    new_n10636_, new_n10637_, new_n10638_, new_n10639_, new_n10640_,
    new_n10641_, new_n10642_, new_n10643_, new_n10644_, new_n10645_,
    new_n10646_, new_n10647_, new_n10648_, new_n10649_, new_n10650_,
    new_n10651_, new_n10652_, new_n10653_, new_n10654_, new_n10655_,
    new_n10656_, new_n10657_, new_n10658_, new_n10659_, new_n10660_,
    new_n10661_, new_n10662_, new_n10663_, new_n10664_, new_n10665_,
    new_n10666_, new_n10667_, new_n10668_, new_n10669_, new_n10670_,
    new_n10671_, new_n10672_, new_n10673_, new_n10674_, new_n10675_,
    new_n10676_, new_n10677_, new_n10678_, new_n10679_, new_n10680_,
    new_n10681_, new_n10682_, new_n10683_, new_n10684_, new_n10685_,
    new_n10686_, new_n10687_, new_n10688_, new_n10689_, new_n10690_,
    new_n10691_, new_n10692_, new_n10693_, new_n10694_, new_n10695_,
    new_n10696_, new_n10697_, new_n10698_, new_n10699_, new_n10700_,
    new_n10701_, new_n10702_, new_n10703_, new_n10704_, new_n10705_,
    new_n10706_, new_n10707_, new_n10708_, new_n10709_, new_n10710_,
    new_n10711_, new_n10712_, new_n10713_, new_n10714_, new_n10715_,
    new_n10716_, new_n10717_, new_n10718_, new_n10719_, new_n10720_,
    new_n10721_, new_n10722_, new_n10723_, new_n10724_, new_n10725_,
    new_n10726_, new_n10727_, new_n10728_, new_n10729_, new_n10730_,
    new_n10731_, new_n10732_, new_n10733_, new_n10734_, new_n10735_,
    new_n10736_, new_n10737_, new_n10738_, new_n10739_, new_n10740_,
    new_n10741_, new_n10742_, new_n10743_, new_n10744_, new_n10745_,
    new_n10746_, new_n10747_, new_n10748_, new_n10749_, new_n10750_,
    new_n10751_, new_n10752_, new_n10753_, new_n10754_, new_n10755_,
    new_n10756_, new_n10757_, new_n10758_, new_n10759_, new_n10760_,
    new_n10761_, new_n10762_, new_n10763_, new_n10764_, new_n10765_,
    new_n10766_, new_n10767_, new_n10768_, new_n10769_, new_n10770_,
    new_n10771_, new_n10772_, new_n10773_, new_n10774_, new_n10775_,
    new_n10776_, new_n10777_, new_n10778_, new_n10779_, new_n10780_,
    new_n10781_, new_n10782_, new_n10783_, new_n10784_, new_n10785_,
    new_n10786_, new_n10787_, new_n10788_, new_n10789_, new_n10790_,
    new_n10791_, new_n10792_, new_n10793_, new_n10794_, new_n10795_,
    new_n10796_, new_n10797_, new_n10798_, new_n10799_, new_n10800_,
    new_n10801_, new_n10802_, new_n10803_, new_n10804_, new_n10805_,
    new_n10806_, new_n10807_, new_n10808_, new_n10809_, new_n10810_,
    new_n10811_, new_n10812_, new_n10813_, new_n10814_, new_n10815_,
    new_n10816_, new_n10817_, new_n10818_, new_n10819_, new_n10820_,
    new_n10821_, new_n10822_, new_n10823_, new_n10824_, new_n10825_,
    new_n10826_, new_n10827_, new_n10828_, new_n10829_, new_n10830_,
    new_n10831_, new_n10832_, new_n10833_, new_n10834_, new_n10835_,
    new_n10836_, new_n10837_, new_n10838_, new_n10839_, new_n10840_,
    new_n10841_, new_n10842_, new_n10843_, new_n10844_, new_n10845_,
    new_n10846_, new_n10847_, new_n10848_, new_n10849_, new_n10850_,
    new_n10851_, new_n10852_, new_n10853_, new_n10854_, new_n10855_,
    new_n10856_, new_n10857_, new_n10858_, new_n10859_, new_n10860_,
    new_n10861_, new_n10862_, new_n10863_, new_n10864_, new_n10865_,
    new_n10866_, new_n10867_, new_n10868_, new_n10869_, new_n10870_,
    new_n10871_, new_n10872_, new_n10873_, new_n10874_, new_n10875_,
    new_n10876_, new_n10877_, new_n10878_, new_n10879_, new_n10880_,
    new_n10881_, new_n10882_, new_n10883_, new_n10884_, new_n10885_,
    new_n10886_, new_n10887_, new_n10888_, new_n10889_, new_n10890_,
    new_n10891_, new_n10892_, new_n10893_, new_n10894_, new_n10895_,
    new_n10896_, new_n10897_, new_n10898_, new_n10899_, new_n10900_,
    new_n10901_, new_n10902_, new_n10903_, new_n10904_, new_n10905_,
    new_n10906_, new_n10907_, new_n10908_, new_n10909_, new_n10910_,
    new_n10911_, new_n10912_, new_n10913_, new_n10914_, new_n10915_,
    new_n10916_, new_n10917_, new_n10918_, new_n10919_, new_n10920_,
    new_n10921_, new_n10922_, new_n10923_, new_n10924_, new_n10925_,
    new_n10926_, new_n10927_, new_n10928_, new_n10929_, new_n10930_,
    new_n10931_, new_n10932_, new_n10933_, new_n10934_, new_n10935_,
    new_n10936_, new_n10937_, new_n10938_, new_n10939_, new_n10940_,
    new_n10941_, new_n10942_, new_n10943_, new_n10944_, new_n10945_,
    new_n10946_, new_n10947_, new_n10948_, new_n10949_, new_n10950_,
    new_n10951_, new_n10952_, new_n10953_, new_n10954_, new_n10955_,
    new_n10956_, new_n10957_, new_n10958_, new_n10959_, new_n10960_,
    new_n10961_, new_n10962_, new_n10963_, new_n10964_, new_n10965_,
    new_n10966_, new_n10967_, new_n10968_, new_n10969_, new_n10970_,
    new_n10971_, new_n10972_, new_n10973_, new_n10974_, new_n10975_,
    new_n10976_, new_n10977_, new_n10978_, new_n10979_, new_n10980_,
    new_n10981_, new_n10982_, new_n10983_, new_n10984_, new_n10985_,
    new_n10986_, new_n10987_, new_n10988_, new_n10989_, new_n10990_,
    new_n10991_, new_n10992_, new_n10993_, new_n10994_, new_n10995_,
    new_n10996_, new_n10997_, new_n10998_, new_n10999_, new_n11000_,
    new_n11001_, new_n11002_, new_n11003_, new_n11004_, new_n11005_,
    new_n11006_, new_n11007_, new_n11008_, new_n11009_, new_n11010_,
    new_n11011_, new_n11012_, new_n11013_, new_n11014_, new_n11015_,
    new_n11016_, new_n11017_, new_n11018_, new_n11019_, new_n11020_,
    new_n11021_, new_n11022_, new_n11023_, new_n11024_, new_n11025_,
    new_n11026_, new_n11027_, new_n11028_, new_n11029_, new_n11030_,
    new_n11031_, new_n11032_, new_n11033_, new_n11034_, new_n11035_,
    new_n11036_, new_n11037_, new_n11038_, new_n11039_, new_n11040_,
    new_n11041_, new_n11042_, new_n11043_, new_n11044_, new_n11045_,
    new_n11046_, new_n11047_, new_n11048_, new_n11049_, new_n11050_,
    new_n11051_, new_n11052_, new_n11053_, new_n11054_, new_n11055_,
    new_n11056_, new_n11057_, new_n11058_, new_n11059_, new_n11060_,
    new_n11061_, new_n11062_, new_n11063_, new_n11064_, new_n11065_,
    new_n11066_, new_n11067_, new_n11068_, new_n11069_, new_n11070_,
    new_n11071_, new_n11072_, new_n11073_, new_n11074_, new_n11075_,
    new_n11076_, new_n11077_, new_n11078_, new_n11079_, new_n11080_,
    new_n11081_, new_n11082_, new_n11083_, new_n11084_, new_n11085_,
    new_n11086_, new_n11087_, new_n11088_, new_n11089_, new_n11090_,
    new_n11091_, new_n11092_, new_n11093_, new_n11094_, new_n11095_,
    new_n11096_, new_n11097_, new_n11098_, new_n11099_, new_n11100_,
    new_n11101_, new_n11102_, new_n11103_, new_n11104_, new_n11105_,
    new_n11106_, new_n11107_, new_n11108_, new_n11109_, new_n11110_,
    new_n11111_, new_n11112_, new_n11113_, new_n11114_, new_n11115_,
    new_n11116_, new_n11117_, new_n11118_, new_n11119_, new_n11120_,
    new_n11121_, new_n11122_, new_n11123_, new_n11124_, new_n11125_,
    new_n11126_, new_n11127_, new_n11128_, new_n11129_, new_n11130_,
    new_n11131_, new_n11132_, new_n11133_, new_n11134_, new_n11135_,
    new_n11136_, new_n11137_, new_n11138_, new_n11139_, new_n11140_,
    new_n11141_, new_n11142_, new_n11143_, new_n11144_, new_n11145_,
    new_n11146_, new_n11147_, new_n11148_, new_n11149_, new_n11150_,
    new_n11151_, new_n11152_, new_n11153_, new_n11154_, new_n11155_,
    new_n11156_, new_n11157_, new_n11158_, new_n11159_, new_n11160_,
    new_n11161_, new_n11162_, new_n11163_, new_n11164_, new_n11165_,
    new_n11166_, new_n11167_, new_n11168_, new_n11169_, new_n11170_,
    new_n11171_, new_n11172_, new_n11173_, new_n11174_, new_n11175_,
    new_n11176_, new_n11177_, new_n11178_, new_n11179_, new_n11180_,
    new_n11181_, new_n11182_, new_n11183_, new_n11184_, new_n11185_,
    new_n11186_, new_n11187_, new_n11188_, new_n11189_, new_n11190_,
    new_n11191_, new_n11192_, new_n11193_, new_n11194_, new_n11195_,
    new_n11196_, new_n11197_, new_n11198_, new_n11199_, new_n11200_,
    new_n11201_, new_n11202_, new_n11203_, new_n11204_, new_n11205_,
    new_n11206_, new_n11207_, new_n11208_, new_n11209_, new_n11210_,
    new_n11211_, new_n11212_, new_n11213_, new_n11214_, new_n11215_,
    new_n11216_, new_n11217_, new_n11218_, new_n11219_, new_n11220_,
    new_n11221_, new_n11222_, new_n11223_, new_n11224_, new_n11225_,
    new_n11226_, new_n11227_, new_n11228_, new_n11229_, new_n11230_,
    new_n11231_, new_n11232_, new_n11233_, new_n11234_, new_n11235_,
    new_n11236_, new_n11237_, new_n11238_, new_n11239_, new_n11240_,
    new_n11241_, new_n11242_, new_n11243_, new_n11244_, new_n11245_,
    new_n11246_, new_n11247_, new_n11248_, new_n11249_, new_n11250_,
    new_n11251_, new_n11252_, new_n11253_, new_n11254_, new_n11255_,
    new_n11256_, new_n11257_, new_n11258_, new_n11259_, new_n11260_,
    new_n11261_, new_n11262_, new_n11263_, new_n11264_, new_n11265_,
    new_n11266_, new_n11267_, new_n11268_, new_n11269_, new_n11270_,
    new_n11271_, new_n11272_, new_n11273_, new_n11274_, new_n11275_,
    new_n11276_, new_n11277_, new_n11278_, new_n11279_, new_n11280_,
    new_n11281_, new_n11282_, new_n11283_, new_n11284_, new_n11285_,
    new_n11286_, new_n11287_, new_n11288_, new_n11289_, new_n11290_,
    new_n11291_, new_n11292_, new_n11293_, new_n11294_, new_n11295_,
    new_n11296_, new_n11297_, new_n11298_, new_n11299_, new_n11300_,
    new_n11301_, new_n11302_, new_n11303_, new_n11304_, new_n11305_,
    new_n11306_, new_n11307_, new_n11308_, new_n11309_, new_n11310_,
    new_n11311_, new_n11312_, new_n11313_, new_n11314_, new_n11315_,
    new_n11316_, new_n11317_, new_n11318_, new_n11319_, new_n11320_,
    new_n11321_, new_n11322_, new_n11323_, new_n11324_, new_n11325_,
    new_n11326_, new_n11327_, new_n11328_, new_n11329_, new_n11330_,
    new_n11331_, new_n11332_, new_n11333_, new_n11334_, new_n11335_,
    new_n11336_, new_n11337_, new_n11338_, new_n11339_, new_n11340_,
    new_n11341_, new_n11342_, new_n11343_, new_n11344_, new_n11345_,
    new_n11346_, new_n11347_, new_n11348_, new_n11349_, new_n11350_,
    new_n11351_, new_n11352_, new_n11353_, new_n11354_, new_n11355_,
    new_n11356_, new_n11357_, new_n11358_, new_n11359_, new_n11360_,
    new_n11361_, new_n11362_, new_n11363_, new_n11364_, new_n11365_,
    new_n11366_, new_n11367_, new_n11368_, new_n11369_, new_n11370_,
    new_n11371_, new_n11372_, new_n11373_, new_n11374_, new_n11375_,
    new_n11376_, new_n11377_, new_n11378_, new_n11379_, new_n11380_,
    new_n11381_, new_n11382_, new_n11383_, new_n11384_, new_n11385_,
    new_n11386_, new_n11387_, new_n11388_, new_n11389_, new_n11390_,
    new_n11391_, new_n11392_, new_n11393_, new_n11394_, new_n11395_,
    new_n11396_, new_n11397_, new_n11398_, new_n11399_, new_n11400_,
    new_n11401_, new_n11402_, new_n11403_, new_n11404_, new_n11405_,
    new_n11406_, new_n11407_, new_n11408_, new_n11409_, new_n11410_,
    new_n11411_, new_n11412_, new_n11413_, new_n11414_, new_n11415_,
    new_n11416_, new_n11417_, new_n11418_, new_n11419_, new_n11420_,
    new_n11421_, new_n11422_, new_n11423_, new_n11424_, new_n11425_,
    new_n11426_, new_n11427_, new_n11428_, new_n11429_, new_n11430_,
    new_n11431_, new_n11432_, new_n11433_, new_n11434_, new_n11435_,
    new_n11436_, new_n11437_, new_n11438_, new_n11439_, new_n11440_,
    new_n11441_, new_n11442_, new_n11443_, new_n11444_, new_n11445_,
    new_n11446_, new_n11447_, new_n11448_, new_n11449_, new_n11450_,
    new_n11451_, new_n11452_, new_n11453_, new_n11454_, new_n11455_,
    new_n11456_, new_n11457_, new_n11458_, new_n11459_, new_n11460_,
    new_n11461_, new_n11462_, new_n11463_, new_n11464_, new_n11465_,
    new_n11466_, new_n11467_, new_n11468_, new_n11469_, new_n11470_,
    new_n11471_, new_n11472_, new_n11473_, new_n11474_, new_n11475_,
    new_n11476_, new_n11477_, new_n11478_, new_n11479_, new_n11480_,
    new_n11481_, new_n11482_, new_n11483_, new_n11484_, new_n11485_,
    new_n11486_, new_n11487_, new_n11488_, new_n11489_, new_n11490_,
    new_n11491_, new_n11492_, new_n11493_, new_n11494_, new_n11495_,
    new_n11496_, new_n11497_, new_n11498_, new_n11499_, new_n11500_,
    new_n11501_, new_n11502_, new_n11503_, new_n11504_, new_n11505_,
    new_n11506_, new_n11507_, new_n11508_, new_n11509_, new_n11510_,
    new_n11511_, new_n11512_, new_n11513_, new_n11514_, new_n11515_,
    new_n11516_, new_n11517_, new_n11518_, new_n11519_, new_n11520_,
    new_n11521_, new_n11522_, new_n11523_, new_n11524_, new_n11525_,
    new_n11526_, new_n11527_, new_n11528_, new_n11529_, new_n11530_,
    new_n11531_, new_n11532_, new_n11533_, new_n11534_, new_n11535_,
    new_n11536_, new_n11537_, new_n11538_, new_n11539_, new_n11540_,
    new_n11541_, new_n11542_, new_n11543_, new_n11544_, new_n11545_,
    new_n11546_, new_n11547_, new_n11548_, new_n11549_, new_n11550_,
    new_n11551_, new_n11552_, new_n11553_, new_n11554_, new_n11555_,
    new_n11556_, new_n11557_, new_n11558_, new_n11559_, new_n11560_,
    new_n11561_, new_n11562_, new_n11563_, new_n11564_, new_n11565_,
    new_n11566_, new_n11567_, new_n11568_, new_n11569_, new_n11570_,
    new_n11571_, new_n11572_, new_n11573_, new_n11574_, new_n11575_,
    new_n11576_, new_n11577_, new_n11578_, new_n11579_, new_n11580_,
    new_n11581_, new_n11582_, new_n11583_, new_n11584_, new_n11585_,
    new_n11586_, new_n11587_, new_n11588_, new_n11589_, new_n11590_,
    new_n11591_, new_n11592_, new_n11593_, new_n11594_, new_n11595_,
    new_n11596_, new_n11597_, new_n11598_, new_n11599_, new_n11600_,
    new_n11601_, new_n11602_, new_n11603_, new_n11604_, new_n11605_,
    new_n11606_, new_n11607_, new_n11608_, new_n11609_, new_n11610_,
    new_n11611_, new_n11612_, new_n11613_, new_n11614_, new_n11615_,
    new_n11616_, new_n11617_, new_n11618_, new_n11619_, new_n11620_,
    new_n11621_, new_n11622_, new_n11623_, new_n11624_, new_n11625_,
    new_n11626_, new_n11627_, new_n11628_, new_n11629_, new_n11630_,
    new_n11631_, new_n11632_, new_n11633_, new_n11634_, new_n11635_,
    new_n11636_, new_n11637_, new_n11638_, new_n11639_, new_n11640_,
    new_n11641_, new_n11642_, new_n11643_, new_n11644_, new_n11645_,
    new_n11646_, new_n11647_, new_n11648_, new_n11649_, new_n11650_,
    new_n11651_, new_n11652_, new_n11653_, new_n11654_, new_n11655_,
    new_n11656_, new_n11657_, new_n11658_, new_n11659_, new_n11660_,
    new_n11661_, new_n11662_, new_n11663_, new_n11664_, new_n11665_,
    new_n11666_, new_n11667_, new_n11668_, new_n11669_, new_n11670_,
    new_n11671_, new_n11672_, new_n11673_, new_n11674_, new_n11675_,
    new_n11676_, new_n11677_, new_n11678_, new_n11679_, new_n11680_,
    new_n11681_, new_n11682_, new_n11683_, new_n11684_, new_n11685_,
    new_n11686_, new_n11687_, new_n11688_, new_n11689_, new_n11690_,
    new_n11691_, new_n11692_, new_n11693_, new_n11694_, new_n11695_,
    new_n11696_, new_n11697_, new_n11698_, new_n11699_, new_n11700_,
    new_n11701_, new_n11702_, new_n11703_, new_n11704_, new_n11705_,
    new_n11706_, new_n11707_, new_n11708_, new_n11709_, new_n11710_,
    new_n11711_, new_n11712_, new_n11713_, new_n11714_, new_n11715_,
    new_n11716_, new_n11717_, new_n11718_, new_n11719_, new_n11720_,
    new_n11721_, new_n11722_, new_n11723_, new_n11724_, new_n11725_,
    new_n11726_, new_n11727_, new_n11728_, new_n11729_, new_n11730_,
    new_n11731_, new_n11732_, new_n11733_, new_n11734_, new_n11735_,
    new_n11736_, new_n11737_, new_n11738_, new_n11739_, new_n11740_,
    new_n11741_, new_n11742_, new_n11743_, new_n11744_, new_n11745_,
    new_n11746_, new_n11747_, new_n11748_, new_n11749_, new_n11750_,
    new_n11751_, new_n11752_, new_n11753_, new_n11754_, new_n11755_,
    new_n11756_, new_n11757_, new_n11758_, new_n11759_, new_n11760_,
    new_n11761_, new_n11762_, new_n11763_, new_n11764_, new_n11765_,
    new_n11766_, new_n11767_, new_n11768_, new_n11769_, new_n11770_,
    new_n11771_, new_n11772_, new_n11773_, new_n11774_, new_n11775_,
    new_n11776_, new_n11777_, new_n11778_, new_n11779_, new_n11780_,
    new_n11781_, new_n11782_, new_n11783_, new_n11784_, new_n11785_,
    new_n11786_, new_n11787_, new_n11788_, new_n11789_, new_n11790_,
    new_n11791_, new_n11792_, new_n11793_, new_n11794_, new_n11795_,
    new_n11796_, new_n11797_, new_n11798_, new_n11799_, new_n11800_,
    new_n11801_, new_n11802_, new_n11803_, new_n11804_, new_n11805_,
    new_n11806_, new_n11807_, new_n11808_, new_n11809_, new_n11810_,
    new_n11811_, new_n11812_, new_n11813_, new_n11814_, new_n11815_,
    new_n11816_, new_n11817_, new_n11818_, new_n11819_, new_n11820_,
    new_n11821_, new_n11822_, new_n11823_, new_n11824_, new_n11825_,
    new_n11826_, new_n11827_, new_n11828_, new_n11829_, new_n11830_,
    new_n11831_, new_n11832_, new_n11833_, new_n11834_, new_n11835_,
    new_n11836_, new_n11837_, new_n11838_, new_n11839_, new_n11840_,
    new_n11841_, new_n11842_, new_n11843_, new_n11844_, new_n11845_,
    new_n11846_, new_n11847_, new_n11848_, new_n11849_, new_n11850_,
    new_n11851_, new_n11852_, new_n11853_, new_n11854_, new_n11855_,
    new_n11856_, new_n11857_, new_n11858_, new_n11859_, new_n11860_,
    new_n11861_, new_n11862_, new_n11863_, new_n11864_, new_n11865_,
    new_n11866_, new_n11867_, new_n11868_, new_n11869_, new_n11870_,
    new_n11871_, new_n11872_, new_n11873_, new_n11874_, new_n11875_,
    new_n11876_, new_n11877_, new_n11878_, new_n11879_, new_n11880_,
    new_n11881_, new_n11882_, new_n11883_, new_n11884_, new_n11885_,
    new_n11886_, new_n11887_, new_n11888_, new_n11889_, new_n11890_,
    new_n11891_, new_n11892_, new_n11893_, new_n11894_, new_n11895_,
    new_n11896_, new_n11897_, new_n11898_, new_n11899_, new_n11900_,
    new_n11901_, new_n11902_, new_n11903_, new_n11904_, new_n11905_,
    new_n11906_, new_n11907_, new_n11908_, new_n11909_, new_n11910_,
    new_n11911_, new_n11912_, new_n11913_, new_n11914_, new_n11915_,
    new_n11916_, new_n11917_, new_n11918_, new_n11919_, new_n11920_,
    new_n11921_, new_n11922_, new_n11923_, new_n11924_, new_n11925_,
    new_n11926_, new_n11927_, new_n11928_, new_n11929_, new_n11930_,
    new_n11931_, new_n11932_, new_n11933_, new_n11934_, new_n11935_,
    new_n11936_, new_n11937_, new_n11938_, new_n11939_, new_n11940_,
    new_n11941_, new_n11942_, new_n11943_, new_n11944_, new_n11945_,
    new_n11946_, new_n11947_, new_n11948_, new_n11949_, new_n11950_,
    new_n11951_, new_n11952_, new_n11953_, new_n11954_, new_n11955_,
    new_n11956_, new_n11957_, new_n11958_, new_n11959_, new_n11960_,
    new_n11961_, new_n11962_, new_n11963_, new_n11964_, new_n11965_,
    new_n11966_, new_n11967_, new_n11968_, new_n11969_, new_n11970_,
    new_n11971_, new_n11972_, new_n11973_, new_n11974_, new_n11975_,
    new_n11976_, new_n11977_, new_n11978_, new_n11979_, new_n11980_,
    new_n11981_, new_n11982_, new_n11983_, new_n11984_, new_n11985_,
    new_n11986_, new_n11987_, new_n11988_, new_n11989_, new_n11990_,
    new_n11991_, new_n11992_, new_n11993_, new_n11994_, new_n11995_,
    new_n11996_, new_n11997_, new_n11998_, new_n11999_, new_n12000_,
    new_n12001_, new_n12002_, new_n12003_, new_n12004_, new_n12005_,
    new_n12006_, new_n12007_, new_n12008_, new_n12009_, new_n12010_,
    new_n12011_, new_n12012_, new_n12013_, new_n12014_, new_n12015_,
    new_n12016_, new_n12017_, new_n12018_, new_n12019_, new_n12020_,
    new_n12021_, new_n12022_, new_n12023_, new_n12024_, new_n12025_,
    new_n12026_, new_n12027_, new_n12028_, new_n12029_, new_n12030_,
    new_n12031_, new_n12032_, new_n12033_, new_n12034_, new_n12035_,
    new_n12036_, new_n12037_, new_n12038_, new_n12039_, new_n12040_,
    new_n12041_, new_n12042_, new_n12043_, new_n12044_, new_n12045_,
    new_n12046_, new_n12047_, new_n12048_, new_n12049_, new_n12050_,
    new_n12051_, new_n12052_, new_n12053_, new_n12054_, new_n12055_,
    new_n12056_, new_n12057_, new_n12058_, new_n12059_, new_n12060_,
    new_n12061_, new_n12062_, new_n12063_, new_n12064_, new_n12065_,
    new_n12066_, new_n12067_, new_n12068_, new_n12069_, new_n12070_,
    new_n12071_, new_n12072_, new_n12073_, new_n12074_, new_n12075_,
    new_n12076_, new_n12077_, new_n12078_, new_n12079_, new_n12080_,
    new_n12081_, new_n12082_, new_n12083_, new_n12084_, new_n12085_,
    new_n12086_, new_n12087_, new_n12088_, new_n12089_, new_n12090_,
    new_n12091_, new_n12092_, new_n12093_, new_n12094_, new_n12095_,
    new_n12096_, new_n12097_, new_n12098_, new_n12099_, new_n12100_,
    new_n12101_, new_n12102_, new_n12103_, new_n12104_, new_n12105_,
    new_n12106_, new_n12107_, new_n12108_, new_n12109_, new_n12110_,
    new_n12111_, new_n12112_, new_n12113_, new_n12114_, new_n12115_,
    new_n12116_, new_n12117_, new_n12118_, new_n12119_, new_n12120_,
    new_n12121_, new_n12122_, new_n12123_, new_n12124_, new_n12125_,
    new_n12126_, new_n12127_, new_n12128_, new_n12129_, new_n12130_,
    new_n12131_, new_n12132_, new_n12133_, new_n12134_, new_n12135_,
    new_n12136_, new_n12137_, new_n12138_, new_n12139_, new_n12140_,
    new_n12141_, new_n12142_, new_n12143_, new_n12144_, new_n12145_,
    new_n12146_, new_n12147_, new_n12148_, new_n12149_, new_n12150_,
    new_n12151_, new_n12152_, new_n12153_, new_n12154_, new_n12155_,
    new_n12156_, new_n12157_, new_n12158_, new_n12159_, new_n12160_,
    new_n12161_, new_n12162_, new_n12163_, new_n12164_, new_n12165_,
    new_n12166_, new_n12167_, new_n12168_, new_n12169_, new_n12170_,
    new_n12171_, new_n12172_, new_n12173_, new_n12174_, new_n12175_,
    new_n12176_, new_n12177_, new_n12178_, new_n12179_, new_n12180_,
    new_n12181_, new_n12182_, new_n12183_, new_n12184_, new_n12185_,
    new_n12186_, new_n12187_, new_n12188_, new_n12189_, new_n12190_,
    new_n12191_, new_n12192_, new_n12193_, new_n12194_, new_n12195_,
    new_n12196_, new_n12197_, new_n12198_, new_n12199_, new_n12200_,
    new_n12201_, new_n12202_, new_n12203_, new_n12204_, new_n12205_,
    new_n12206_, new_n12207_, new_n12208_, new_n12209_, new_n12210_,
    new_n12211_, new_n12212_, new_n12213_, new_n12214_, new_n12215_,
    new_n12216_, new_n12217_, new_n12218_, new_n12219_, new_n12220_,
    new_n12221_, new_n12222_, new_n12223_, new_n12224_, new_n12225_,
    new_n12226_, new_n12227_, new_n12228_, new_n12229_, new_n12230_,
    new_n12231_, new_n12232_, new_n12233_, new_n12234_, new_n12235_,
    new_n12236_, new_n12237_, new_n12238_, new_n12239_, new_n12240_,
    new_n12241_, new_n12242_, new_n12243_, new_n12244_, new_n12245_,
    new_n12246_, new_n12247_, new_n12248_, new_n12249_, new_n12250_,
    new_n12251_, new_n12252_, new_n12253_, new_n12254_, new_n12255_,
    new_n12256_, new_n12257_, new_n12258_, new_n12259_, new_n12260_,
    new_n12261_, new_n12262_, new_n12263_, new_n12264_, new_n12265_,
    new_n12266_, new_n12267_, new_n12268_, new_n12269_, new_n12270_,
    new_n12271_, new_n12272_, new_n12273_, new_n12274_, new_n12275_,
    new_n12276_, new_n12277_, new_n12278_, new_n12279_, new_n12280_,
    new_n12281_, new_n12282_, new_n12283_, new_n12284_, new_n12285_,
    new_n12286_, new_n12287_, new_n12288_, new_n12289_, new_n12290_,
    new_n12291_, new_n12292_, new_n12293_, new_n12294_, new_n12295_,
    new_n12296_, new_n12297_, new_n12298_, new_n12299_, new_n12300_,
    new_n12301_, new_n12302_, new_n12303_, new_n12304_, new_n12305_,
    new_n12306_, new_n12307_, new_n12308_, new_n12309_, new_n12310_,
    new_n12311_, new_n12312_, new_n12313_, new_n12314_, new_n12315_,
    new_n12316_, new_n12317_, new_n12318_, new_n12319_, new_n12320_,
    new_n12321_, new_n12322_, new_n12323_, new_n12324_, new_n12325_,
    new_n12326_, new_n12327_, new_n12328_, new_n12329_, new_n12330_,
    new_n12331_, new_n12332_, new_n12333_, new_n12334_, new_n12335_,
    new_n12336_, new_n12337_, new_n12338_, new_n12339_, new_n12340_,
    new_n12341_, new_n12342_, new_n12343_, new_n12344_, new_n12345_,
    new_n12346_, new_n12347_, new_n12348_, new_n12349_, new_n12350_,
    new_n12351_, new_n12352_, new_n12353_, new_n12354_, new_n12355_,
    new_n12356_, new_n12357_, new_n12358_, new_n12359_, new_n12360_,
    new_n12361_, new_n12362_, new_n12363_, new_n12364_, new_n12365_,
    new_n12366_, new_n12367_, new_n12368_, new_n12369_, new_n12370_,
    new_n12371_, new_n12372_, new_n12373_, new_n12374_, new_n12375_,
    new_n12376_, new_n12377_, new_n12378_, new_n12379_, new_n12380_,
    new_n12381_, new_n12382_, new_n12383_, new_n12384_, new_n12385_,
    new_n12386_, new_n12387_, new_n12388_, new_n12389_, new_n12390_,
    new_n12391_, new_n12392_, new_n12393_, new_n12394_, new_n12395_,
    new_n12396_, new_n12397_, new_n12398_, new_n12399_, new_n12400_,
    new_n12401_, new_n12402_, new_n12403_, new_n12404_, new_n12405_,
    new_n12406_, new_n12407_, new_n12408_, new_n12409_, new_n12410_,
    new_n12411_, new_n12412_, new_n12413_, new_n12414_, new_n12415_,
    new_n12416_, new_n12417_, new_n12418_, new_n12419_, new_n12420_,
    new_n12421_, new_n12422_, new_n12423_, new_n12424_, new_n12425_,
    new_n12426_, new_n12427_, new_n12428_, new_n12429_, new_n12430_,
    new_n12431_, new_n12432_, new_n12433_, new_n12434_, new_n12435_,
    new_n12436_, new_n12437_, new_n12438_, new_n12439_, new_n12440_,
    new_n12441_, new_n12442_, new_n12443_, new_n12444_, new_n12445_,
    new_n12446_, new_n12447_, new_n12448_, new_n12449_, new_n12450_,
    new_n12451_, new_n12452_, new_n12453_, new_n12454_, new_n12455_,
    new_n12456_, new_n12457_, new_n12458_, new_n12459_, new_n12460_,
    new_n12461_, new_n12462_, new_n12463_, new_n12464_, new_n12465_,
    new_n12466_, new_n12467_, new_n12468_, new_n12469_, new_n12470_,
    new_n12471_, new_n12472_, new_n12473_, new_n12474_, new_n12475_,
    new_n12476_, new_n12477_, new_n12478_, new_n12479_, new_n12480_,
    new_n12481_, new_n12482_, new_n12483_, new_n12484_, new_n12485_,
    new_n12486_, new_n12487_, new_n12488_, new_n12489_, new_n12490_,
    new_n12491_, new_n12492_, new_n12493_, new_n12494_, new_n12495_,
    new_n12496_, new_n12497_, new_n12498_, new_n12499_, new_n12500_,
    new_n12501_, new_n12502_, new_n12503_, new_n12504_, new_n12505_,
    new_n12506_, new_n12507_, new_n12508_, new_n12509_, new_n12510_,
    new_n12511_, new_n12512_, new_n12513_, new_n12514_, new_n12515_,
    new_n12516_, new_n12517_, new_n12518_, new_n12519_, new_n12520_,
    new_n12521_, new_n12522_, new_n12523_, new_n12524_, new_n12525_,
    new_n12526_, new_n12527_, new_n12528_, new_n12529_, new_n12530_,
    new_n12531_, new_n12532_, new_n12533_, new_n12534_, new_n12535_,
    new_n12536_, new_n12537_, new_n12538_, new_n12539_, new_n12540_,
    new_n12541_, new_n12542_, new_n12543_, new_n12544_, new_n12545_,
    new_n12546_, new_n12547_, new_n12548_, new_n12549_, new_n12550_,
    new_n12551_, new_n12552_, new_n12553_, new_n12554_, new_n12555_,
    new_n12556_, new_n12557_, new_n12558_, new_n12559_, new_n12560_,
    new_n12561_, new_n12562_, new_n12563_, new_n12564_, new_n12565_,
    new_n12566_, new_n12567_, new_n12568_, new_n12569_, new_n12570_,
    new_n12571_, new_n12572_, new_n12573_, new_n12574_, new_n12575_,
    new_n12576_, new_n12577_, new_n12578_, new_n12579_, new_n12580_,
    new_n12581_, new_n12582_, new_n12583_, new_n12584_, new_n12585_,
    new_n12586_, new_n12587_, new_n12588_, new_n12589_, new_n12590_,
    new_n12591_, new_n12592_, new_n12593_, new_n12594_, new_n12595_,
    new_n12596_, new_n12597_, new_n12598_, new_n12599_, new_n12600_,
    new_n12601_, new_n12602_, new_n12603_, new_n12604_, new_n12605_,
    new_n12606_, new_n12607_, new_n12608_, new_n12609_, new_n12610_,
    new_n12611_, new_n12612_, new_n12613_, new_n12614_, new_n12615_,
    new_n12616_, new_n12617_, new_n12618_, new_n12619_, new_n12620_,
    new_n12621_, new_n12622_, new_n12623_, new_n12624_, new_n12625_,
    new_n12626_, new_n12627_, new_n12628_, new_n12629_, new_n12630_,
    new_n12631_, new_n12632_, new_n12633_, new_n12634_, new_n12635_,
    new_n12636_, new_n12637_, new_n12638_, new_n12639_, new_n12640_,
    new_n12641_, new_n12642_, new_n12643_, new_n12644_, new_n12645_,
    new_n12646_, new_n12647_, new_n12648_, new_n12649_, new_n12650_,
    new_n12651_, new_n12652_, new_n12653_, new_n12654_, new_n12655_,
    new_n12656_, new_n12657_, new_n12658_, new_n12659_, new_n12660_,
    new_n12661_, new_n12662_, new_n12663_, new_n12664_, new_n12665_,
    new_n12666_, new_n12667_, new_n12668_, new_n12669_, new_n12670_,
    new_n12671_, new_n12672_, new_n12673_, new_n12674_, new_n12675_,
    new_n12676_, new_n12677_, new_n12678_, new_n12679_, new_n12680_,
    new_n12681_, new_n12682_, new_n12683_, new_n12684_, new_n12685_,
    new_n12686_, new_n12687_, new_n12688_, new_n12689_, new_n12690_,
    new_n12691_, new_n12692_, new_n12693_, new_n12694_, new_n12695_,
    new_n12696_, new_n12697_, new_n12698_, new_n12699_, new_n12700_,
    new_n12701_, new_n12702_, new_n12703_, new_n12704_, new_n12705_,
    new_n12706_, new_n12707_, new_n12708_, new_n12709_, new_n12710_,
    new_n12711_, new_n12712_, new_n12713_, new_n12714_, new_n12715_,
    new_n12716_, new_n12717_, new_n12718_, new_n12719_, new_n12720_,
    new_n12721_, new_n12722_, new_n12723_, new_n12724_, new_n12725_,
    new_n12726_, new_n12727_, new_n12728_, new_n12729_, new_n12730_,
    new_n12731_, new_n12732_, new_n12733_, new_n12734_, new_n12735_,
    new_n12736_, new_n12737_, new_n12738_, new_n12739_, new_n12740_,
    new_n12741_, new_n12742_, new_n12743_, new_n12744_, new_n12745_,
    new_n12746_, new_n12747_, new_n12748_, new_n12749_, new_n12750_,
    new_n12751_, new_n12752_, new_n12753_, new_n12754_, new_n12755_,
    new_n12756_, new_n12757_, new_n12758_, new_n12759_, new_n12760_,
    new_n12761_, new_n12762_, new_n12763_, new_n12764_, new_n12765_,
    new_n12766_, new_n12767_, new_n12768_, new_n12769_, new_n12770_,
    new_n12771_, new_n12772_, new_n12773_, new_n12774_, new_n12775_,
    new_n12776_, new_n12777_, new_n12778_, new_n12779_, new_n12780_,
    new_n12781_, new_n12782_, new_n12783_, new_n12784_, new_n12785_,
    new_n12786_, new_n12787_, new_n12788_, new_n12789_, new_n12790_,
    new_n12791_, new_n12792_, new_n12793_, new_n12794_, new_n12795_,
    new_n12796_, new_n12797_, new_n12798_, new_n12799_, new_n12800_,
    new_n12801_, new_n12802_, new_n12803_, new_n12804_, new_n12805_,
    new_n12806_, new_n12807_, new_n12808_, new_n12809_, new_n12810_,
    new_n12811_, new_n12812_, new_n12813_, new_n12814_, new_n12815_,
    new_n12816_, new_n12817_, new_n12818_, new_n12819_, new_n12820_,
    new_n12821_, new_n12822_, new_n12823_, new_n12824_, new_n12825_,
    new_n12826_, new_n12827_, new_n12828_, new_n12829_, new_n12830_,
    new_n12831_, new_n12832_, new_n12833_, new_n12834_, new_n12835_,
    new_n12836_, new_n12837_, new_n12838_, new_n12839_, new_n12840_,
    new_n12841_, new_n12842_, new_n12843_, new_n12844_, new_n12845_,
    new_n12846_, new_n12847_, new_n12848_, new_n12849_, new_n12850_,
    new_n12851_, new_n12852_, new_n12853_, new_n12854_, new_n12855_,
    new_n12856_, new_n12857_, new_n12858_, new_n12859_, new_n12860_,
    new_n12861_, new_n12862_, new_n12863_, new_n12864_, new_n12865_,
    new_n12866_, new_n12867_, new_n12868_, new_n12869_, new_n12870_,
    new_n12871_, new_n12872_, new_n12873_, new_n12874_, new_n12875_,
    new_n12876_, new_n12877_, new_n12878_, new_n12879_, new_n12880_,
    new_n12881_, new_n12882_, new_n12883_, new_n12884_, new_n12885_,
    new_n12886_, new_n12887_, new_n12888_, new_n12889_, new_n12890_,
    new_n12891_, new_n12892_, new_n12893_, new_n12894_, new_n12895_,
    new_n12896_, new_n12897_, new_n12898_, new_n12899_, new_n12900_,
    new_n12901_, new_n12902_, new_n12903_, new_n12904_, new_n12905_,
    new_n12906_, new_n12907_, new_n12908_, new_n12909_, new_n12910_,
    new_n12911_, new_n12912_, new_n12913_, new_n12914_, new_n12915_,
    new_n12916_, new_n12917_, new_n12918_, new_n12919_, new_n12920_,
    new_n12921_, new_n12922_, new_n12923_, new_n12924_, new_n12925_,
    new_n12926_, new_n12927_, new_n12928_, new_n12929_, new_n12930_,
    new_n12931_, new_n12932_, new_n12933_, new_n12934_, new_n12935_,
    new_n12936_, new_n12937_, new_n12938_, new_n12939_, new_n12940_,
    new_n12941_, new_n12942_, new_n12943_, new_n12944_, new_n12945_,
    new_n12946_, new_n12947_, new_n12948_, new_n12949_, new_n12950_,
    new_n12951_, new_n12952_, new_n12953_, new_n12954_, new_n12955_,
    new_n12956_, new_n12957_, new_n12958_, new_n12959_, new_n12960_,
    new_n12961_, new_n12962_, new_n12963_, new_n12964_, new_n12965_,
    new_n12966_, new_n12967_, new_n12968_, new_n12969_, new_n12970_,
    new_n12971_, new_n12972_, new_n12973_, new_n12974_, new_n12975_,
    new_n12976_, new_n12977_, new_n12978_, new_n12979_, new_n12980_,
    new_n12981_, new_n12982_, new_n12983_, new_n12984_, new_n12985_,
    new_n12986_, new_n12987_, new_n12988_, new_n12989_, new_n12990_,
    new_n12991_, new_n12992_, new_n12993_, new_n12994_, new_n12995_,
    new_n12996_, new_n12997_, new_n12998_, new_n12999_, new_n13000_,
    new_n13001_, new_n13002_, new_n13003_, new_n13004_, new_n13005_,
    new_n13006_, new_n13007_, new_n13008_, new_n13009_, new_n13010_,
    new_n13011_, new_n13012_, new_n13013_, new_n13014_, new_n13015_,
    new_n13016_, new_n13017_, new_n13018_, new_n13019_, new_n13020_,
    new_n13021_, new_n13022_, new_n13023_, new_n13024_, new_n13025_,
    new_n13026_, new_n13027_, new_n13028_, new_n13029_, new_n13030_,
    new_n13031_, new_n13032_, new_n13033_, new_n13034_, new_n13035_,
    new_n13036_, new_n13037_, new_n13038_, new_n13039_, new_n13040_,
    new_n13041_, new_n13042_, new_n13043_, new_n13044_, new_n13045_,
    new_n13046_, new_n13047_, new_n13048_, new_n13049_, new_n13050_,
    new_n13051_, new_n13052_, new_n13053_, new_n13054_, new_n13055_,
    new_n13056_, new_n13057_, new_n13058_, new_n13059_, new_n13060_,
    new_n13061_, new_n13062_, new_n13063_, new_n13064_, new_n13065_,
    new_n13066_, new_n13067_, new_n13068_, new_n13069_, new_n13070_,
    new_n13071_, new_n13072_, new_n13073_, new_n13074_, new_n13075_,
    new_n13076_, new_n13077_, new_n13078_, new_n13079_, new_n13080_,
    new_n13081_, new_n13082_, new_n13083_, new_n13084_, new_n13085_,
    new_n13086_, new_n13087_, new_n13088_, new_n13089_, new_n13090_,
    new_n13091_, new_n13092_, new_n13093_, new_n13094_, new_n13095_,
    new_n13096_, new_n13097_, new_n13098_, new_n13099_, new_n13100_,
    new_n13101_, new_n13102_, new_n13103_, new_n13104_, new_n13105_,
    new_n13106_, new_n13107_, new_n13108_, new_n13109_, new_n13110_,
    new_n13111_, new_n13112_, new_n13113_, new_n13114_, new_n13115_,
    new_n13116_, new_n13117_, new_n13118_, new_n13119_, new_n13120_,
    new_n13121_, new_n13122_, new_n13123_, new_n13124_, new_n13125_,
    new_n13126_, new_n13127_, new_n13128_, new_n13129_, new_n13130_,
    new_n13131_, new_n13132_, new_n13133_, new_n13134_, new_n13135_,
    new_n13136_, new_n13137_, new_n13138_, new_n13139_, new_n13140_,
    new_n13141_, new_n13142_, new_n13143_, new_n13144_, new_n13145_,
    new_n13146_, new_n13147_, new_n13148_, new_n13149_, new_n13150_,
    new_n13151_, new_n13152_, new_n13153_, new_n13154_, new_n13155_,
    new_n13156_, new_n13157_, new_n13158_, new_n13159_, new_n13160_,
    new_n13161_, new_n13162_, new_n13163_, new_n13164_, new_n13165_,
    new_n13166_, new_n13167_, new_n13168_, new_n13169_, new_n13170_,
    new_n13171_, new_n13172_, new_n13173_, new_n13174_, new_n13175_,
    new_n13176_, new_n13177_, new_n13178_, new_n13179_, new_n13180_,
    new_n13181_, new_n13182_, new_n13183_, new_n13184_, new_n13185_,
    new_n13186_, new_n13187_, new_n13188_, new_n13189_, new_n13190_,
    new_n13191_, new_n13192_, new_n13193_, new_n13194_, new_n13195_,
    new_n13196_, new_n13197_, new_n13198_, new_n13199_, new_n13200_,
    new_n13201_, new_n13202_, new_n13203_, new_n13204_, new_n13205_,
    new_n13206_, new_n13207_, new_n13208_, new_n13209_, new_n13210_,
    new_n13211_, new_n13212_, new_n13213_, new_n13214_, new_n13215_,
    new_n13216_, new_n13217_, new_n13218_, new_n13219_, new_n13220_,
    new_n13221_, new_n13222_, new_n13223_, new_n13224_, new_n13225_,
    new_n13226_, new_n13227_, new_n13228_, new_n13229_, new_n13230_,
    new_n13231_, new_n13232_, new_n13233_, new_n13234_, new_n13235_,
    new_n13236_, new_n13237_, new_n13238_, new_n13239_, new_n13240_,
    new_n13241_, new_n13242_, new_n13243_, new_n13244_, new_n13245_,
    new_n13246_, new_n13247_, new_n13248_, new_n13249_, new_n13250_,
    new_n13251_, new_n13252_, new_n13253_, new_n13254_, new_n13255_,
    new_n13256_, new_n13257_, new_n13258_, new_n13259_, new_n13260_,
    new_n13261_, new_n13262_, new_n13263_, new_n13264_, new_n13265_,
    new_n13266_, new_n13267_, new_n13268_, new_n13269_, new_n13270_,
    new_n13271_, new_n13272_, new_n13273_, new_n13274_, new_n13275_,
    new_n13276_, new_n13277_, new_n13278_, new_n13279_, new_n13280_,
    new_n13281_, new_n13282_, new_n13283_, new_n13284_, new_n13285_,
    new_n13286_, new_n13287_, new_n13288_, new_n13289_, new_n13290_,
    new_n13291_, new_n13292_, new_n13293_, new_n13294_, new_n13295_,
    new_n13296_, new_n13297_, new_n13298_, new_n13299_, new_n13300_,
    new_n13301_, new_n13302_, new_n13303_, new_n13304_, new_n13305_,
    new_n13306_, new_n13307_, new_n13308_, new_n13309_, new_n13310_,
    new_n13311_, new_n13312_, new_n13313_, new_n13314_, new_n13315_,
    new_n13316_, new_n13317_, new_n13318_, new_n13319_, new_n13320_,
    new_n13321_, new_n13322_, new_n13323_, new_n13324_, new_n13325_,
    new_n13326_, new_n13327_, new_n13328_, new_n13329_, new_n13330_,
    new_n13331_, new_n13332_, new_n13333_, new_n13334_, new_n13335_,
    new_n13336_, new_n13337_, new_n13338_, new_n13339_, new_n13340_,
    new_n13341_, new_n13342_, new_n13343_, new_n13344_, new_n13345_,
    new_n13346_, new_n13347_, new_n13348_, new_n13349_, new_n13350_,
    new_n13351_, new_n13352_, new_n13353_, new_n13354_, new_n13355_,
    new_n13356_, new_n13357_, new_n13358_, new_n13359_, new_n13360_,
    new_n13361_, new_n13362_, new_n13363_, new_n13364_, new_n13365_,
    new_n13366_, new_n13367_, new_n13368_, new_n13369_, new_n13370_,
    new_n13371_, new_n13372_, new_n13373_, new_n13374_, new_n13375_,
    new_n13376_, new_n13377_, new_n13378_, new_n13379_, new_n13380_,
    new_n13381_, new_n13382_, new_n13383_, new_n13384_, new_n13385_,
    new_n13386_, new_n13387_, new_n13388_, new_n13389_, new_n13390_,
    new_n13391_, new_n13392_, new_n13393_, new_n13394_, new_n13395_,
    new_n13396_, new_n13397_, new_n13398_, new_n13399_, new_n13400_,
    new_n13401_, new_n13402_, new_n13403_, new_n13404_, new_n13405_,
    new_n13406_, new_n13407_, new_n13408_, new_n13409_, new_n13410_,
    new_n13411_, new_n13412_, new_n13413_, new_n13414_, new_n13415_,
    new_n13416_, new_n13417_, new_n13418_, new_n13419_, new_n13420_,
    new_n13421_, new_n13422_, new_n13423_, new_n13424_, new_n13425_,
    new_n13426_, new_n13427_, new_n13428_, new_n13429_, new_n13430_,
    new_n13431_, new_n13432_, new_n13433_, new_n13434_, new_n13435_,
    new_n13436_, new_n13437_, new_n13438_, new_n13439_, new_n13440_,
    new_n13441_, new_n13442_, new_n13443_, new_n13444_, new_n13445_,
    new_n13446_, new_n13447_, new_n13448_, new_n13449_, new_n13450_,
    new_n13451_, new_n13452_, new_n13453_, new_n13454_, new_n13455_,
    new_n13456_, new_n13457_, new_n13458_, new_n13459_, new_n13460_,
    new_n13461_, new_n13462_, new_n13463_, new_n13464_, new_n13465_,
    new_n13466_, new_n13467_, new_n13468_, new_n13469_, new_n13470_,
    new_n13471_, new_n13472_, new_n13473_, new_n13474_, new_n13475_,
    new_n13476_, new_n13477_, new_n13478_, new_n13479_, new_n13480_,
    new_n13481_, new_n13482_, new_n13483_, new_n13484_, new_n13485_,
    new_n13486_, new_n13487_, new_n13488_, new_n13489_, new_n13490_,
    new_n13491_, new_n13492_, new_n13493_, new_n13494_, new_n13495_,
    new_n13496_, new_n13497_, new_n13498_, new_n13499_, new_n13500_,
    new_n13501_, new_n13502_, new_n13503_, new_n13504_, new_n13505_,
    new_n13506_, new_n13507_, new_n13508_, new_n13509_, new_n13510_,
    new_n13511_, new_n13512_, new_n13513_, new_n13514_, new_n13515_,
    new_n13516_, new_n13517_, new_n13518_, new_n13519_, new_n13520_,
    new_n13521_, new_n13522_, new_n13523_, new_n13524_, new_n13525_,
    new_n13526_, new_n13527_, new_n13528_, new_n13529_, new_n13530_,
    new_n13531_, new_n13532_, new_n13533_, new_n13534_, new_n13535_,
    new_n13536_, new_n13537_, new_n13538_, new_n13539_, new_n13540_,
    new_n13541_, new_n13542_, new_n13543_, new_n13544_, new_n13545_,
    new_n13546_, new_n13547_, new_n13548_, new_n13549_, new_n13550_,
    new_n13551_, new_n13552_, new_n13553_, new_n13554_, new_n13555_,
    new_n13556_, new_n13557_, new_n13558_, new_n13559_, new_n13560_,
    new_n13561_, new_n13562_, new_n13563_, new_n13564_, new_n13565_,
    new_n13566_, new_n13567_, new_n13568_, new_n13569_, new_n13570_,
    new_n13571_, new_n13572_, new_n13573_, new_n13574_, new_n13575_,
    new_n13576_, new_n13577_, new_n13578_, new_n13579_, new_n13580_,
    new_n13581_, new_n13582_, new_n13583_, new_n13584_, new_n13585_,
    new_n13586_, new_n13587_, new_n13588_, new_n13589_, new_n13590_,
    new_n13591_, new_n13592_, new_n13593_, new_n13594_, new_n13595_,
    new_n13596_, new_n13597_, new_n13598_, new_n13599_, new_n13600_,
    new_n13601_, new_n13602_, new_n13603_, new_n13604_, new_n13605_,
    new_n13606_, new_n13607_, new_n13608_, new_n13609_, new_n13610_,
    new_n13611_, new_n13612_, new_n13613_, new_n13614_, new_n13615_,
    new_n13616_, new_n13617_, new_n13618_, new_n13619_, new_n13620_,
    new_n13621_, new_n13622_, new_n13623_, new_n13624_, new_n13625_,
    new_n13626_, new_n13627_, new_n13628_, new_n13629_, new_n13630_,
    new_n13631_, new_n13632_, new_n13633_, new_n13634_, new_n13635_,
    new_n13636_, new_n13637_, new_n13638_, new_n13639_, new_n13640_,
    new_n13641_, new_n13642_, new_n13643_, new_n13644_, new_n13645_,
    new_n13646_, new_n13647_, new_n13648_, new_n13649_, new_n13650_,
    new_n13651_, new_n13652_, new_n13653_, new_n13654_, new_n13655_,
    new_n13656_, new_n13657_, new_n13658_, new_n13659_, new_n13660_,
    new_n13661_, new_n13662_, new_n13663_, new_n13664_, new_n13665_,
    new_n13666_, new_n13667_, new_n13668_, new_n13669_, new_n13670_,
    new_n13671_, new_n13672_, new_n13673_, new_n13674_, new_n13675_,
    new_n13676_, new_n13677_, new_n13678_, new_n13679_, new_n13680_,
    new_n13681_, new_n13682_, new_n13683_, new_n13684_, new_n13685_,
    new_n13686_, new_n13687_, new_n13688_, new_n13689_, new_n13690_,
    new_n13691_, new_n13692_, new_n13693_, new_n13694_, new_n13695_,
    new_n13696_, new_n13697_, new_n13698_, new_n13699_, new_n13700_,
    new_n13701_, new_n13702_, new_n13703_, new_n13704_, new_n13705_,
    new_n13706_, new_n13707_, new_n13708_, new_n13709_, new_n13710_,
    new_n13711_, new_n13712_, new_n13713_, new_n13714_, new_n13715_,
    new_n13716_, new_n13717_, new_n13718_, new_n13719_, new_n13720_,
    new_n13721_, new_n13722_, new_n13723_, new_n13724_, new_n13725_,
    new_n13726_, new_n13727_, new_n13728_, new_n13729_, new_n13730_,
    new_n13731_, new_n13732_, new_n13733_, new_n13734_, new_n13735_,
    new_n13736_, new_n13737_, new_n13738_, new_n13739_, new_n13740_,
    new_n13741_, new_n13742_, new_n13743_, new_n13744_, new_n13745_,
    new_n13746_, new_n13747_, new_n13748_, new_n13749_, new_n13750_,
    new_n13751_, new_n13752_, new_n13753_, new_n13754_, new_n13755_,
    new_n13756_, new_n13757_, new_n13758_, new_n13759_, new_n13760_,
    new_n13761_, new_n13762_, new_n13763_, new_n13764_, new_n13765_,
    new_n13766_, new_n13767_, new_n13768_, new_n13769_, new_n13770_,
    new_n13771_, new_n13772_, new_n13773_, new_n13774_, new_n13775_,
    new_n13776_, new_n13777_, new_n13778_, new_n13779_, new_n13780_,
    new_n13781_, new_n13782_, new_n13783_, new_n13784_, new_n13785_,
    new_n13786_, new_n13787_, new_n13788_, new_n13789_, new_n13790_,
    new_n13791_, new_n13792_, new_n13793_, new_n13794_, new_n13795_,
    new_n13796_, new_n13797_, new_n13798_, new_n13799_, new_n13800_,
    new_n13801_, new_n13802_, new_n13803_, new_n13804_, new_n13805_,
    new_n13806_, new_n13807_, new_n13808_, new_n13809_, new_n13810_,
    new_n13811_, new_n13812_, new_n13813_, new_n13814_, new_n13815_,
    new_n13816_, new_n13817_, new_n13818_, new_n13819_, new_n13820_,
    new_n13821_, new_n13822_, new_n13823_, new_n13824_, new_n13825_,
    new_n13826_, new_n13827_, new_n13828_, new_n13829_, new_n13830_,
    new_n13831_, new_n13832_, new_n13833_, new_n13834_, new_n13835_,
    new_n13836_, new_n13837_, new_n13838_, new_n13839_, new_n13840_,
    new_n13841_, new_n13842_, new_n13843_, new_n13844_, new_n13845_,
    new_n13846_, new_n13847_, new_n13848_, new_n13849_, new_n13850_,
    new_n13851_, new_n13852_, new_n13853_, new_n13854_, new_n13855_,
    new_n13856_, new_n13857_, new_n13858_, new_n13859_, new_n13860_,
    new_n13861_, new_n13862_, new_n13863_, new_n13864_, new_n13865_,
    new_n13866_, new_n13867_, new_n13868_, new_n13869_, new_n13870_,
    new_n13871_, new_n13872_, new_n13873_, new_n13874_, new_n13875_,
    new_n13876_, new_n13877_, new_n13878_, new_n13879_, new_n13880_,
    new_n13881_, new_n13882_, new_n13883_, new_n13884_, new_n13885_,
    new_n13886_, new_n13887_, new_n13888_, new_n13889_, new_n13890_,
    new_n13891_, new_n13892_, new_n13893_, new_n13894_, new_n13895_,
    new_n13896_, new_n13897_, new_n13898_, new_n13899_, new_n13900_,
    new_n13901_, new_n13902_, new_n13903_, new_n13904_, new_n13905_,
    new_n13906_, new_n13907_, new_n13908_, new_n13909_, new_n13910_,
    new_n13911_, new_n13912_, new_n13913_, new_n13914_, new_n13915_,
    new_n13916_, new_n13917_, new_n13918_, new_n13919_, new_n13920_,
    new_n13921_, new_n13922_, new_n13923_, new_n13924_, new_n13925_,
    new_n13926_, new_n13927_, new_n13928_, new_n13929_, new_n13930_,
    new_n13931_, new_n13932_, new_n13933_, new_n13934_, new_n13935_,
    new_n13936_, new_n13937_, new_n13938_, new_n13939_, new_n13940_,
    new_n13941_, new_n13942_, new_n13943_, new_n13944_, new_n13945_,
    new_n13946_, new_n13947_, new_n13948_, new_n13949_, new_n13950_,
    new_n13951_, new_n13952_, new_n13953_, new_n13954_, new_n13955_,
    new_n13956_, new_n13957_, new_n13958_, new_n13959_, new_n13960_,
    new_n13961_, new_n13962_, new_n13963_, new_n13964_, new_n13965_,
    new_n13966_, new_n13967_, new_n13968_, new_n13969_, new_n13970_,
    new_n13971_, new_n13972_, new_n13973_, new_n13974_, new_n13975_,
    new_n13976_, new_n13977_, new_n13978_, new_n13979_, new_n13980_,
    new_n13981_, new_n13982_, new_n13983_, new_n13984_, new_n13985_,
    new_n13986_, new_n13987_, new_n13988_, new_n13989_, new_n13990_,
    new_n13991_, new_n13992_, new_n13993_, new_n13994_, new_n13995_,
    new_n13996_, new_n13997_, new_n13998_, new_n13999_, new_n14000_,
    new_n14001_, new_n14002_, new_n14003_, new_n14004_, new_n14005_,
    new_n14006_, new_n14007_, new_n14008_, new_n14009_, new_n14010_,
    new_n14011_, new_n14012_, new_n14013_, new_n14014_, new_n14015_,
    new_n14016_, new_n14017_, new_n14018_, new_n14019_, new_n14020_,
    new_n14021_, new_n14022_, new_n14023_, new_n14024_, new_n14025_,
    new_n14026_, new_n14027_, new_n14028_, new_n14029_, new_n14030_,
    new_n14031_, new_n14032_, new_n14033_, new_n14034_, new_n14035_,
    new_n14036_, new_n14037_, new_n14038_, new_n14039_, new_n14040_,
    new_n14041_, new_n14042_, new_n14043_, new_n14044_, new_n14045_,
    new_n14046_, new_n14047_, new_n14048_, new_n14049_, new_n14050_,
    new_n14051_, new_n14052_, new_n14053_, new_n14054_, new_n14055_,
    new_n14056_, new_n14057_, new_n14058_, new_n14059_, new_n14060_,
    new_n14061_, new_n14062_, new_n14063_, new_n14064_, new_n14065_,
    new_n14066_, new_n14067_, new_n14068_, new_n14069_, new_n14070_,
    new_n14071_, new_n14072_, new_n14073_, new_n14074_, new_n14075_,
    new_n14076_, new_n14077_, new_n14078_, new_n14079_, new_n14080_,
    new_n14081_, new_n14082_, new_n14083_, new_n14084_, new_n14085_,
    new_n14086_, new_n14087_, new_n14088_, new_n14089_, new_n14090_,
    new_n14091_, new_n14092_, new_n14093_, new_n14094_, new_n14095_,
    new_n14096_, new_n14097_, new_n14098_, new_n14099_, new_n14100_,
    new_n14101_, new_n14102_, new_n14103_, new_n14104_, new_n14105_,
    new_n14106_, new_n14107_, new_n14108_, new_n14109_, new_n14110_,
    new_n14111_, new_n14112_, new_n14113_, new_n14114_, new_n14115_,
    new_n14116_, new_n14117_, new_n14118_, new_n14119_, new_n14120_,
    new_n14121_, new_n14122_, new_n14123_, new_n14124_, new_n14125_,
    new_n14126_, new_n14127_, new_n14128_, new_n14129_, new_n14130_,
    new_n14131_, new_n14132_, new_n14133_, new_n14134_, new_n14135_,
    new_n14136_, new_n14137_, new_n14138_, new_n14139_, new_n14140_,
    new_n14141_, new_n14142_, new_n14143_, new_n14144_, new_n14145_,
    new_n14146_, new_n14147_, new_n14148_, new_n14149_, new_n14150_,
    new_n14151_, new_n14152_, new_n14153_, new_n14154_, new_n14155_,
    new_n14156_, new_n14157_, new_n14158_, new_n14159_, new_n14160_,
    new_n14161_, new_n14162_, new_n14163_, new_n14164_, new_n14165_,
    new_n14166_, new_n14167_, new_n14168_, new_n14169_, new_n14170_,
    new_n14171_, new_n14172_, new_n14173_, new_n14174_, new_n14175_,
    new_n14176_, new_n14177_, new_n14178_, new_n14179_, new_n14180_,
    new_n14181_, new_n14182_, new_n14183_, new_n14184_, new_n14185_,
    new_n14186_, new_n14187_, new_n14188_, new_n14189_, new_n14190_,
    new_n14191_, new_n14192_, new_n14193_, new_n14194_, new_n14195_,
    new_n14196_, new_n14197_, new_n14198_, new_n14199_, new_n14200_,
    new_n14201_, new_n14202_, new_n14203_, new_n14204_, new_n14205_,
    new_n14206_, new_n14207_, new_n14208_, new_n14209_, new_n14210_,
    new_n14211_, new_n14212_, new_n14213_, new_n14214_, new_n14215_,
    new_n14216_, new_n14217_, new_n14218_, new_n14219_, new_n14220_,
    new_n14221_, new_n14222_, new_n14223_, new_n14224_, new_n14225_,
    new_n14226_, new_n14227_, new_n14228_, new_n14229_, new_n14230_,
    new_n14231_, new_n14232_, new_n14233_, new_n14234_, new_n14235_,
    new_n14236_, new_n14237_, new_n14238_, new_n14239_, new_n14240_,
    new_n14241_, new_n14242_, new_n14243_, new_n14244_, new_n14245_,
    new_n14246_, new_n14247_, new_n14248_, new_n14249_, new_n14250_,
    new_n14251_, new_n14252_, new_n14253_, new_n14254_, new_n14255_,
    new_n14256_, new_n14257_, new_n14258_, new_n14259_, new_n14260_,
    new_n14261_, new_n14262_, new_n14263_, new_n14264_, new_n14265_,
    new_n14266_, new_n14267_, new_n14268_, new_n14269_, new_n14270_,
    new_n14271_, new_n14272_, new_n14273_, new_n14274_, new_n14275_,
    new_n14276_, new_n14277_, new_n14278_, new_n14279_, new_n14280_,
    new_n14281_, new_n14282_, new_n14283_, new_n14284_, new_n14285_,
    new_n14286_, new_n14287_, new_n14288_, new_n14289_, new_n14290_,
    new_n14291_, new_n14292_, new_n14293_, new_n14294_, new_n14295_,
    new_n14296_, new_n14297_, new_n14298_, new_n14299_, new_n14300_,
    new_n14301_, new_n14302_, new_n14303_, new_n14304_, new_n14305_,
    new_n14306_, new_n14307_, new_n14308_, new_n14309_, new_n14310_,
    new_n14311_, new_n14312_, new_n14313_, new_n14314_, new_n14315_,
    new_n14316_, new_n14317_, new_n14318_, new_n14319_, new_n14320_,
    new_n14321_, new_n14322_, new_n14323_, new_n14324_, new_n14325_,
    new_n14326_, new_n14327_, new_n14328_, new_n14329_, new_n14330_,
    new_n14331_, new_n14332_, new_n14333_, new_n14334_, new_n14335_,
    new_n14336_, new_n14337_, new_n14338_, new_n14339_, new_n14340_,
    new_n14341_, new_n14342_, new_n14343_, new_n14344_, new_n14345_,
    new_n14346_, new_n14347_, new_n14348_, new_n14349_, new_n14350_,
    new_n14351_, new_n14352_, new_n14353_, new_n14354_, new_n14355_,
    new_n14356_, new_n14357_, new_n14358_, new_n14359_, new_n14360_,
    new_n14361_, new_n14362_, new_n14363_, new_n14364_, new_n14365_,
    new_n14366_, new_n14367_, new_n14368_, new_n14369_, new_n14370_,
    new_n14371_, new_n14372_, new_n14373_, new_n14374_, new_n14375_,
    new_n14376_, new_n14377_, new_n14378_, new_n14379_, new_n14380_,
    new_n14381_, new_n14382_, new_n14383_, new_n14384_, new_n14385_,
    new_n14386_, new_n14387_, new_n14388_, new_n14389_, new_n14390_,
    new_n14391_, new_n14392_, new_n14393_, new_n14394_, new_n14395_,
    new_n14396_, new_n14397_, new_n14398_, new_n14399_, new_n14400_,
    new_n14401_, new_n14402_, new_n14403_, new_n14404_, new_n14405_,
    new_n14406_, new_n14407_, new_n14408_, new_n14409_, new_n14410_,
    new_n14411_, new_n14412_, new_n14413_, new_n14414_, new_n14415_,
    new_n14416_, new_n14417_, new_n14418_, new_n14419_, new_n14420_,
    new_n14421_, new_n14422_, new_n14423_, new_n14424_, new_n14425_,
    new_n14426_, new_n14427_, new_n14428_, new_n14429_, new_n14430_,
    new_n14431_, new_n14432_, new_n14433_, new_n14434_, new_n14435_,
    new_n14436_, new_n14437_, new_n14438_, new_n14439_, new_n14440_,
    new_n14441_, new_n14442_, new_n14443_, new_n14444_, new_n14445_,
    new_n14446_, new_n14447_, new_n14448_, new_n14449_, new_n14450_,
    new_n14451_, new_n14452_, new_n14453_, new_n14454_, new_n14455_,
    new_n14456_, new_n14457_, new_n14458_, new_n14459_, new_n14460_,
    new_n14461_, new_n14462_, new_n14463_, new_n14464_, new_n14465_,
    new_n14466_, new_n14467_, new_n14468_, new_n14469_, new_n14470_,
    new_n14471_, new_n14472_, new_n14473_, new_n14474_, new_n14475_,
    new_n14476_, new_n14477_, new_n14478_, new_n14479_, new_n14480_,
    new_n14481_, new_n14482_, new_n14483_, new_n14484_, new_n14485_,
    new_n14486_, new_n14487_, new_n14488_, new_n14489_, new_n14490_,
    new_n14491_, new_n14492_, new_n14493_, new_n14494_, new_n14495_,
    new_n14496_, new_n14497_, new_n14498_, new_n14499_, new_n14500_,
    new_n14501_, new_n14502_, new_n14503_, new_n14504_, new_n14505_,
    new_n14506_, new_n14507_, new_n14508_, new_n14509_, new_n14510_,
    new_n14511_, new_n14512_, new_n14513_, new_n14514_, new_n14515_,
    new_n14516_, new_n14517_, new_n14518_, new_n14519_, new_n14520_,
    new_n14521_, new_n14522_, new_n14523_, new_n14524_, new_n14525_,
    new_n14526_, new_n14527_, new_n14528_, new_n14529_, new_n14530_,
    new_n14531_, new_n14532_, new_n14533_, new_n14534_, new_n14535_,
    new_n14536_, new_n14537_, new_n14538_, new_n14539_, new_n14540_,
    new_n14541_, new_n14542_, new_n14543_, new_n14544_, new_n14545_,
    new_n14546_, new_n14547_, new_n14548_, new_n14549_, new_n14550_,
    new_n14551_, new_n14552_, new_n14553_, new_n14554_, new_n14555_,
    new_n14556_, new_n14557_, new_n14558_, new_n14559_, new_n14560_,
    new_n14561_, new_n14562_, new_n14563_, new_n14564_, new_n14565_,
    new_n14566_, new_n14567_, new_n14568_, new_n14569_, new_n14570_,
    new_n14571_, new_n14572_, new_n14573_, new_n14574_, new_n14575_,
    new_n14576_, new_n14577_, new_n14578_, new_n14579_, new_n14580_,
    new_n14581_, new_n14582_, new_n14583_, new_n14584_, new_n14585_,
    new_n14586_, new_n14587_, new_n14588_, new_n14589_, new_n14590_,
    new_n14591_, new_n14592_, new_n14593_, new_n14594_, new_n14595_,
    new_n14596_, new_n14597_, new_n14598_, new_n14599_, new_n14600_,
    new_n14601_, new_n14602_, new_n14603_, new_n14604_, new_n14605_,
    new_n14606_, new_n14607_, new_n14608_, new_n14609_, new_n14610_,
    new_n14611_, new_n14612_, new_n14613_, new_n14614_, new_n14615_,
    new_n14616_, new_n14617_, new_n14618_, new_n14619_, new_n14620_,
    new_n14621_, new_n14622_, new_n14623_, new_n14624_, new_n14625_,
    new_n14626_, new_n14627_, new_n14628_, new_n14629_, new_n14630_,
    new_n14631_, new_n14632_, new_n14633_, new_n14634_, new_n14635_,
    new_n14636_, new_n14637_, new_n14638_, new_n14639_, new_n14640_,
    new_n14641_, new_n14642_, new_n14643_, new_n14644_, new_n14645_,
    new_n14646_, new_n14647_, new_n14648_, new_n14649_, new_n14650_,
    new_n14651_, new_n14652_, new_n14653_, new_n14654_, new_n14655_,
    new_n14656_, new_n14657_, new_n14658_, new_n14659_, new_n14660_,
    new_n14661_, new_n14662_, new_n14663_, new_n14664_, new_n14665_,
    new_n14666_, new_n14667_, new_n14668_, new_n14669_, new_n14670_,
    new_n14671_, new_n14672_, new_n14673_, new_n14674_, new_n14675_,
    new_n14676_, new_n14677_, new_n14678_, new_n14679_, new_n14680_,
    new_n14681_, new_n14682_, new_n14683_, new_n14684_, new_n14685_,
    new_n14686_, new_n14687_, new_n14688_, new_n14689_, new_n14690_,
    new_n14691_, new_n14692_, new_n14693_, new_n14694_, new_n14695_,
    new_n14696_, new_n14697_, new_n14698_, new_n14699_, new_n14700_,
    new_n14701_, new_n14702_, new_n14703_, new_n14704_, new_n14705_,
    new_n14706_, new_n14707_, new_n14708_, new_n14709_, new_n14710_,
    new_n14711_, new_n14712_, new_n14713_, new_n14714_, new_n14715_,
    new_n14716_, new_n14717_, new_n14718_, new_n14719_, new_n14720_,
    new_n14721_, new_n14722_, new_n14723_, new_n14724_, new_n14725_,
    new_n14726_, new_n14727_, new_n14728_, new_n14729_, new_n14730_,
    new_n14731_, new_n14732_, new_n14733_, new_n14734_, new_n14735_,
    new_n14736_, new_n14737_, new_n14738_, new_n14739_, new_n14740_,
    new_n14741_, new_n14742_, new_n14743_, new_n14744_, new_n14745_,
    new_n14746_, new_n14747_, new_n14748_, new_n14749_, new_n14750_,
    new_n14751_, new_n14752_, new_n14753_, new_n14754_, new_n14755_,
    new_n14756_, new_n14757_, new_n14758_, new_n14759_, new_n14760_,
    new_n14761_, new_n14762_, new_n14763_, new_n14764_, new_n14765_,
    new_n14766_, new_n14767_, new_n14768_, new_n14769_, new_n14770_,
    new_n14771_, new_n14772_, new_n14773_, new_n14774_, new_n14775_,
    new_n14776_, new_n14777_, new_n14778_, new_n14779_, new_n14780_,
    new_n14781_, new_n14782_, new_n14783_, new_n14784_, new_n14785_,
    new_n14786_, new_n14787_, new_n14788_, new_n14789_, new_n14790_,
    new_n14791_, new_n14792_, new_n14793_, new_n14794_, new_n14795_,
    new_n14796_, new_n14797_, new_n14798_, new_n14799_, new_n14800_,
    new_n14801_, new_n14802_, new_n14803_, new_n14804_, new_n14805_,
    new_n14806_, new_n14807_, new_n14808_, new_n14809_, new_n14810_,
    new_n14811_, new_n14812_, new_n14813_, new_n14814_, new_n14815_,
    new_n14816_, new_n14817_, new_n14818_, new_n14819_, new_n14820_,
    new_n14821_, new_n14822_, new_n14823_, new_n14824_, new_n14825_,
    new_n14826_, new_n14827_, new_n14828_, new_n14829_, new_n14830_,
    new_n14831_, new_n14832_, new_n14833_, new_n14834_, new_n14835_,
    new_n14836_, new_n14837_, new_n14838_, new_n14839_, new_n14840_,
    new_n14841_, new_n14842_, new_n14843_, new_n14844_, new_n14845_,
    new_n14846_, new_n14847_, new_n14848_, new_n14849_, new_n14850_,
    new_n14851_, new_n14852_, new_n14853_, new_n14854_, new_n14855_,
    new_n14856_, new_n14857_, new_n14858_, new_n14859_, new_n14860_,
    new_n14861_, new_n14862_, new_n14863_, new_n14864_, new_n14865_,
    new_n14866_, new_n14867_, new_n14868_, new_n14869_, new_n14870_,
    new_n14871_, new_n14872_, new_n14873_, new_n14874_, new_n14875_,
    new_n14876_, new_n14877_, new_n14878_, new_n14879_, new_n14880_,
    new_n14881_, new_n14882_, new_n14883_, new_n14884_, new_n14885_,
    new_n14886_, new_n14887_, new_n14888_, new_n14889_, new_n14890_,
    new_n14891_, new_n14892_, new_n14893_, new_n14894_, new_n14895_,
    new_n14896_, new_n14897_, new_n14898_, new_n14899_, new_n14900_,
    new_n14901_, new_n14902_, new_n14903_, new_n14904_, new_n14905_,
    new_n14906_, new_n14907_, new_n14908_, new_n14909_, new_n14910_,
    new_n14911_, new_n14912_, new_n14913_, new_n14914_, new_n14915_,
    new_n14916_, new_n14917_, new_n14918_, new_n14919_, new_n14920_,
    new_n14921_, new_n14922_, new_n14923_, new_n14924_, new_n14925_,
    new_n14926_, new_n14927_, new_n14928_, new_n14929_, new_n14930_,
    new_n14931_, new_n14932_, new_n14933_, new_n14934_, new_n14935_,
    new_n14936_, new_n14937_, new_n14938_, new_n14939_, new_n14940_,
    new_n14941_, new_n14942_, new_n14943_, new_n14944_, new_n14945_,
    new_n14946_, new_n14947_, new_n14948_, new_n14949_, new_n14950_,
    new_n14951_, new_n14952_, new_n14953_, new_n14954_, new_n14955_,
    new_n14956_, new_n14957_, new_n14958_, new_n14959_, new_n14960_,
    new_n14961_, new_n14962_, new_n14963_, new_n14964_, new_n14965_,
    new_n14966_, new_n14967_, new_n14968_, new_n14969_, new_n14970_,
    new_n14971_, new_n14972_, new_n14973_, new_n14974_, new_n14975_,
    new_n14976_, new_n14977_, new_n14978_, new_n14979_, new_n14980_,
    new_n14981_, new_n14982_, new_n14983_, new_n14984_, new_n14985_,
    new_n14986_, new_n14987_, new_n14988_, new_n14989_, new_n14990_,
    new_n14991_, new_n14992_, new_n14993_, new_n14994_, new_n14995_,
    new_n14996_, new_n14997_, new_n14998_, new_n14999_, new_n15000_,
    new_n15001_, new_n15002_, new_n15003_, new_n15004_, new_n15005_,
    new_n15006_, new_n15007_, new_n15008_, new_n15009_, new_n15010_,
    new_n15011_, new_n15012_, new_n15013_, new_n15014_, new_n15015_,
    new_n15016_, new_n15017_, new_n15018_, new_n15019_, new_n15020_,
    new_n15021_, new_n15022_, new_n15023_, new_n15024_, new_n15025_,
    new_n15026_, new_n15027_, new_n15028_, new_n15029_, new_n15030_,
    new_n15031_, new_n15032_, new_n15033_, new_n15034_, new_n15035_,
    new_n15036_, new_n15037_, new_n15038_, new_n15039_, new_n15040_,
    new_n15041_, new_n15042_, new_n15043_, new_n15044_, new_n15045_,
    new_n15046_, new_n15047_, new_n15048_, new_n15049_, new_n15050_,
    new_n15051_, new_n15052_, new_n15053_, new_n15054_, new_n15055_,
    new_n15056_, new_n15057_, new_n15058_, new_n15059_, new_n15060_,
    new_n15061_, new_n15062_, new_n15063_, new_n15064_, new_n15065_,
    new_n15066_, new_n15067_, new_n15068_, new_n15069_, new_n15070_,
    new_n15071_, new_n15072_, new_n15073_, new_n15074_, new_n15075_,
    new_n15076_, new_n15077_, new_n15078_, new_n15079_, new_n15080_,
    new_n15081_, new_n15082_, new_n15083_, new_n15084_, new_n15085_,
    new_n15086_, new_n15087_, new_n15088_, new_n15089_, new_n15090_,
    new_n15091_, new_n15092_, new_n15093_, new_n15094_, new_n15095_,
    new_n15096_, new_n15097_, new_n15098_, new_n15099_, new_n15100_,
    new_n15101_, new_n15102_, new_n15103_, new_n15104_, new_n15105_,
    new_n15106_, new_n15107_, new_n15108_, new_n15109_, new_n15110_,
    new_n15111_, new_n15112_, new_n15113_, new_n15114_, new_n15115_,
    new_n15116_, new_n15117_, new_n15118_, new_n15119_, new_n15120_,
    new_n15121_, new_n15122_, new_n15123_, new_n15124_, new_n15125_,
    new_n15126_, new_n15127_, new_n15128_, new_n15129_, new_n15130_,
    new_n15131_, new_n15132_, new_n15133_, new_n15134_, new_n15135_,
    new_n15136_, new_n15137_, new_n15138_, new_n15139_, new_n15140_,
    new_n15141_, new_n15142_, new_n15143_, new_n15144_, new_n15145_,
    new_n15146_, new_n15147_, new_n15148_, new_n15149_, new_n15150_,
    new_n15151_, new_n15152_, new_n15153_, new_n15154_, new_n15155_,
    new_n15156_, new_n15157_, new_n15158_, new_n15159_, new_n15160_,
    new_n15161_, new_n15162_, new_n15163_, new_n15164_, new_n15165_,
    new_n15166_, new_n15167_, new_n15168_, new_n15169_, new_n15170_,
    new_n15171_, new_n15172_, new_n15173_, new_n15174_, new_n15175_,
    new_n15176_, new_n15177_, new_n15178_, new_n15179_, new_n15180_,
    new_n15181_, new_n15182_, new_n15183_, new_n15184_, new_n15185_,
    new_n15186_, new_n15187_, new_n15188_, new_n15189_, new_n15190_,
    new_n15191_, new_n15192_, new_n15193_, new_n15194_, new_n15195_,
    new_n15196_, new_n15197_, new_n15198_, new_n15199_, new_n15200_,
    new_n15201_, new_n15202_, new_n15203_, new_n15204_, new_n15205_,
    new_n15206_, new_n15207_, new_n15208_, new_n15209_, new_n15210_,
    new_n15211_, new_n15212_, new_n15213_, new_n15214_, new_n15215_,
    new_n15216_, new_n15217_, new_n15218_, new_n15219_, new_n15220_,
    new_n15221_, new_n15222_, new_n15223_, new_n15224_, new_n15225_,
    new_n15226_, new_n15227_, new_n15228_, new_n15229_, new_n15230_,
    new_n15231_, new_n15232_, new_n15233_, new_n15234_, new_n15235_,
    new_n15236_, new_n15237_, new_n15238_, new_n15239_, new_n15240_,
    new_n15241_, new_n15242_, new_n15243_, new_n15244_, new_n15245_,
    new_n15246_, new_n15247_, new_n15248_, new_n15249_, new_n15250_,
    new_n15251_, new_n15252_, new_n15253_, new_n15254_, new_n15255_,
    new_n15256_, new_n15257_, new_n15258_, new_n15259_, new_n15260_,
    new_n15261_, new_n15262_, new_n15263_, new_n15264_, new_n15265_,
    new_n15266_, new_n15267_, new_n15268_, new_n15269_, new_n15270_,
    new_n15271_, new_n15272_, new_n15273_, new_n15274_, new_n15275_,
    new_n15276_, new_n15277_, new_n15278_, new_n15279_, new_n15280_,
    new_n15281_, new_n15282_, new_n15283_, new_n15284_, new_n15285_,
    new_n15286_, new_n15287_, new_n15288_, new_n15289_, new_n15290_,
    new_n15291_, new_n15292_, new_n15293_, new_n15294_, new_n15295_,
    new_n15296_, new_n15297_, new_n15298_, new_n15299_, new_n15300_,
    new_n15301_, new_n15302_, new_n15303_, new_n15304_, new_n15305_,
    new_n15306_, new_n15307_, new_n15308_, new_n15309_, new_n15310_,
    new_n15311_, new_n15312_, new_n15313_, new_n15314_, new_n15315_,
    new_n15316_, new_n15317_, new_n15318_, new_n15319_, new_n15320_,
    new_n15321_, new_n15322_, new_n15323_, new_n15324_, new_n15325_,
    new_n15326_, new_n15327_, new_n15328_, new_n15329_, new_n15330_,
    new_n15331_, new_n15332_, new_n15333_, new_n15334_, new_n15335_,
    new_n15336_, new_n15337_, new_n15338_, new_n15339_, new_n15340_,
    new_n15341_, new_n15342_, new_n15343_, new_n15344_, new_n15345_,
    new_n15346_, new_n15347_, new_n15348_, new_n15349_, new_n15350_,
    new_n15351_, new_n15352_, new_n15353_, new_n15354_, new_n15355_,
    new_n15356_, new_n15357_, new_n15358_, new_n15359_, new_n15360_,
    new_n15361_, new_n15362_, new_n15363_, new_n15364_, new_n15365_,
    new_n15366_, new_n15367_, new_n15368_, new_n15369_, new_n15370_,
    new_n15371_, new_n15372_, new_n15373_, new_n15374_, new_n15375_,
    new_n15376_, new_n15377_, new_n15378_, new_n15379_, new_n15380_,
    new_n15381_, new_n15382_, new_n15383_, new_n15384_, new_n15385_,
    new_n15386_, new_n15387_, new_n15388_, new_n15389_, new_n15390_,
    new_n15391_, new_n15392_, new_n15393_, new_n15394_, new_n15395_,
    new_n15396_, new_n15397_, new_n15398_, new_n15399_, new_n15400_,
    new_n15401_, new_n15402_, new_n15403_, new_n15404_, new_n15405_,
    new_n15406_, new_n15407_, new_n15408_, new_n15409_, new_n15410_,
    new_n15411_, new_n15412_, new_n15413_, new_n15414_, new_n15415_,
    new_n15416_, new_n15417_, new_n15418_, new_n15419_, new_n15420_,
    new_n15421_, new_n15422_, new_n15423_, new_n15424_, new_n15425_,
    new_n15426_, new_n15427_, new_n15428_, new_n15429_, new_n15430_,
    new_n15431_, new_n15432_, new_n15433_, new_n15434_, new_n15435_,
    new_n15436_, new_n15437_, new_n15438_, new_n15439_, new_n15440_,
    new_n15441_, new_n15442_, new_n15443_, new_n15444_, new_n15445_,
    new_n15446_, new_n15447_, new_n15448_, new_n15449_, new_n15450_,
    new_n15451_, new_n15452_, new_n15453_, new_n15454_, new_n15455_,
    new_n15456_, new_n15457_, new_n15458_, new_n15459_, new_n15460_,
    new_n15461_, new_n15462_, new_n15463_, new_n15464_, new_n15465_,
    new_n15466_, new_n15467_, new_n15468_, new_n15469_, new_n15470_,
    new_n15471_, new_n15472_, new_n15473_, new_n15474_, new_n15475_,
    new_n15476_, new_n15477_, new_n15478_, new_n15479_, new_n15480_,
    new_n15481_, new_n15482_, new_n15483_, new_n15484_, new_n15485_,
    new_n15486_, new_n15487_, new_n15488_, new_n15489_, new_n15490_,
    new_n15491_, new_n15492_, new_n15493_, new_n15494_, new_n15495_,
    new_n15496_, new_n15497_, new_n15498_, new_n15499_, new_n15500_,
    new_n15501_, new_n15502_, new_n15503_, new_n15504_, new_n15505_,
    new_n15506_, new_n15507_, new_n15508_, new_n15509_, new_n15510_,
    new_n15511_, new_n15512_, new_n15513_, new_n15514_, new_n15515_,
    new_n15516_, new_n15517_, new_n15518_, new_n15519_, new_n15520_,
    new_n15521_, new_n15522_, new_n15523_, new_n15524_, new_n15525_,
    new_n15526_, new_n15527_, new_n15528_, new_n15529_, new_n15530_,
    new_n15531_, new_n15532_, new_n15533_, new_n15534_, new_n15535_,
    new_n15536_, new_n15537_, new_n15538_, new_n15539_, new_n15540_,
    new_n15541_, new_n15542_, new_n15543_, new_n15544_, new_n15545_,
    new_n15546_, new_n15547_, new_n15548_, new_n15549_, new_n15550_,
    new_n15551_, new_n15552_, new_n15553_, new_n15554_, new_n15555_,
    new_n15556_, new_n15557_, new_n15558_, new_n15559_, new_n15560_,
    new_n15561_, new_n15562_, new_n15563_, new_n15564_, new_n15565_,
    new_n15566_, new_n15567_, new_n15568_, new_n15569_, new_n15570_,
    new_n15571_, new_n15572_, new_n15573_, new_n15574_, new_n15575_,
    new_n15576_, new_n15577_, new_n15578_, new_n15579_, new_n15580_,
    new_n15581_, new_n15582_, new_n15583_, new_n15584_, new_n15585_,
    new_n15586_, new_n15587_, new_n15588_, new_n15589_, new_n15590_,
    new_n15591_, new_n15592_, new_n15593_, new_n15594_, new_n15595_,
    new_n15596_, new_n15597_, new_n15598_, new_n15599_, new_n15600_,
    new_n15601_, new_n15602_, new_n15603_, new_n15604_, new_n15605_,
    new_n15606_, new_n15607_, new_n15608_, new_n15609_, new_n15610_,
    new_n15611_, new_n15612_, new_n15613_, new_n15614_, new_n15615_,
    new_n15616_, new_n15617_, new_n15618_, new_n15619_, new_n15620_,
    new_n15621_, new_n15622_, new_n15623_, new_n15624_, new_n15625_,
    new_n15626_, new_n15627_, new_n15628_, new_n15629_, new_n15630_,
    new_n15631_, new_n15632_, new_n15633_, new_n15634_, new_n15635_,
    new_n15636_, new_n15637_, new_n15638_, new_n15639_, new_n15640_,
    new_n15641_, new_n15642_, new_n15643_, new_n15644_, new_n15645_,
    new_n15646_, new_n15647_, new_n15648_, new_n15649_, new_n15650_,
    new_n15651_, new_n15652_, new_n15653_, new_n15654_, new_n15655_,
    new_n15656_, new_n15657_, new_n15658_, new_n15659_, new_n15660_,
    new_n15661_, new_n15662_, new_n15663_, new_n15664_, new_n15665_,
    new_n15666_, new_n15667_, new_n15668_, new_n15669_, new_n15670_,
    new_n15671_, new_n15672_, new_n15673_, new_n15674_, new_n15675_,
    new_n15676_, new_n15677_, new_n15678_, new_n15679_, new_n15680_,
    new_n15681_, new_n15682_, new_n15683_, new_n15684_, new_n15685_,
    new_n15686_, new_n15687_, new_n15688_, new_n15689_, new_n15690_,
    new_n15691_, new_n15692_, new_n15693_, new_n15694_, new_n15695_,
    new_n15696_, new_n15697_, new_n15698_, new_n15699_, new_n15700_,
    new_n15701_, new_n15702_, new_n15703_, new_n15704_, new_n15705_,
    new_n15706_, new_n15707_, new_n15708_, new_n15709_, new_n15710_,
    new_n15711_, new_n15712_, new_n15713_, new_n15714_, new_n15715_,
    new_n15716_, new_n15717_, new_n15718_, new_n15719_, new_n15720_,
    new_n15721_, new_n15722_, new_n15723_, new_n15724_, new_n15725_,
    new_n15726_, new_n15727_, new_n15728_, new_n15729_, new_n15730_,
    new_n15731_, new_n15732_, new_n15733_, new_n15734_, new_n15735_,
    new_n15736_, new_n15737_, new_n15738_, new_n15739_, new_n15740_,
    new_n15741_, new_n15742_, new_n15743_, new_n15744_, new_n15745_,
    new_n15746_, new_n15747_, new_n15748_, new_n15749_, new_n15750_,
    new_n15751_, new_n15752_, new_n15753_, new_n15754_, new_n15755_,
    new_n15756_, new_n15757_, new_n15758_, new_n15759_, new_n15760_,
    new_n15761_, new_n15762_, new_n15763_, new_n15764_, new_n15765_,
    new_n15766_, new_n15767_, new_n15768_, new_n15769_, new_n15770_,
    new_n15771_, new_n15772_, new_n15773_, new_n15774_, new_n15775_,
    new_n15776_, new_n15777_, new_n15778_, new_n15779_, new_n15780_,
    new_n15781_, new_n15782_, new_n15783_, new_n15784_, new_n15785_,
    new_n15786_, new_n15787_, new_n15788_, new_n15789_, new_n15790_,
    new_n15791_, new_n15792_, new_n15793_, new_n15794_, new_n15795_,
    new_n15796_, new_n15797_, new_n15798_, new_n15799_, new_n15800_,
    new_n15801_, new_n15802_, new_n15803_, new_n15804_, new_n15805_,
    new_n15806_, new_n15807_, new_n15808_, new_n15809_, new_n15810_,
    new_n15811_, new_n15812_, new_n15813_, new_n15814_, new_n15815_,
    new_n15816_, new_n15817_, new_n15818_, new_n15819_, new_n15820_,
    new_n15821_, new_n15822_, new_n15823_, new_n15824_, new_n15825_,
    new_n15826_, new_n15827_, new_n15828_, new_n15829_, new_n15830_,
    new_n15831_, new_n15832_, new_n15833_, new_n15834_, new_n15835_,
    new_n15836_, new_n15837_, new_n15838_, new_n15839_, new_n15840_,
    new_n15841_, new_n15842_, new_n15843_, new_n15844_, new_n15845_,
    new_n15846_, new_n15847_, new_n15848_, new_n15849_, new_n15850_,
    new_n15851_, new_n15852_, new_n15853_, new_n15854_, new_n15855_,
    new_n15856_, new_n15857_, new_n15858_, new_n15859_, new_n15860_,
    new_n15861_, new_n15862_, new_n15863_, new_n15864_, new_n15865_,
    new_n15866_, new_n15867_, new_n15868_, new_n15869_, new_n15870_,
    new_n15871_, new_n15872_, new_n15873_, new_n15874_, new_n15875_,
    new_n15876_, new_n15877_, new_n15878_, new_n15879_, new_n15880_,
    new_n15881_, new_n15882_, new_n15883_, new_n15884_, new_n15885_,
    new_n15886_, new_n15887_, new_n15888_, new_n15889_, new_n15890_,
    new_n15891_, new_n15892_, new_n15893_, new_n15894_, new_n15895_,
    new_n15896_, new_n15897_, new_n15898_, new_n15899_, new_n15900_,
    new_n15901_, new_n15902_, new_n15903_, new_n15904_, new_n15905_,
    new_n15906_, new_n15907_, new_n15908_, new_n15909_, new_n15910_,
    new_n15911_, new_n15912_, new_n15913_, new_n15914_, new_n15915_,
    new_n15916_, new_n15917_, new_n15918_, new_n15919_, new_n15920_,
    new_n15921_, new_n15922_, new_n15923_, new_n15924_, new_n15925_,
    new_n15926_, new_n15927_, new_n15928_, new_n15929_, new_n15930_,
    new_n15931_, new_n15932_, new_n15933_, new_n15934_, new_n15935_,
    new_n15936_, new_n15937_, new_n15938_, new_n15939_, new_n15940_,
    new_n15941_, new_n15942_, new_n15943_, new_n15944_, new_n15945_,
    new_n15946_, new_n15947_, new_n15948_, new_n15949_, new_n15950_,
    new_n15951_, new_n15952_, new_n15953_, new_n15954_, new_n15955_,
    new_n15956_, new_n15957_, new_n15958_, new_n15959_, new_n15960_,
    new_n15961_, new_n15962_, new_n15963_, new_n15964_, new_n15965_,
    new_n15966_, new_n15967_, new_n15968_, new_n15969_, new_n15970_,
    new_n15971_, new_n15972_, new_n15973_, new_n15974_, new_n15975_,
    new_n15976_, new_n15977_, new_n15978_, new_n15979_, new_n15980_,
    new_n15981_, new_n15982_, new_n15983_, new_n15984_, new_n15985_,
    new_n15986_, new_n15987_, new_n15988_, new_n15989_, new_n15990_,
    new_n15991_, new_n15992_, new_n15993_, new_n15994_, new_n15995_,
    new_n15996_, new_n15997_, new_n15998_, new_n15999_, new_n16000_,
    new_n16001_, new_n16002_, new_n16003_, new_n16004_, new_n16005_,
    new_n16006_, new_n16007_, new_n16008_, new_n16009_, new_n16010_,
    new_n16011_, new_n16012_, new_n16013_, new_n16014_, new_n16015_,
    new_n16016_, new_n16017_, new_n16018_, new_n16019_, new_n16020_,
    new_n16021_, new_n16022_, new_n16023_, new_n16024_, new_n16025_,
    new_n16026_, new_n16027_, new_n16028_, new_n16029_, new_n16030_,
    new_n16031_, new_n16032_, new_n16033_, new_n16034_, new_n16035_,
    new_n16036_, new_n16037_, new_n16038_, new_n16039_, new_n16040_,
    new_n16041_, new_n16042_, new_n16043_, new_n16044_, new_n16045_,
    new_n16046_, new_n16047_, new_n16048_, new_n16049_, new_n16050_,
    new_n16051_, new_n16052_, new_n16053_, new_n16054_, new_n16055_,
    new_n16056_, new_n16057_, new_n16058_, new_n16059_, new_n16060_,
    new_n16061_, new_n16062_, new_n16063_, new_n16064_, new_n16065_,
    new_n16066_, new_n16067_, new_n16068_, new_n16069_, new_n16070_,
    new_n16071_, new_n16073_, new_n16074_, new_n16075_, new_n16076_,
    new_n16077_;
  INV    g00000(.A(\A[717] ), .Y(new_n1003_));
  INV    g00001(.A(\A[715] ), .Y(new_n1004_));
  NAND2  g00002(.A(\A[716] ), .B(new_n1004_), .Y(new_n1005_));
  INV    g00003(.A(\A[716] ), .Y(new_n1006_));
  AOI21  g00004(.A0(new_n1006_), .A1(\A[715] ), .B0(new_n1003_), .Y(new_n1007_));
  XOR2   g00005(.A(\A[716] ), .B(\A[715] ), .Y(new_n1008_));
  AOI22  g00006(.A0(new_n1008_), .A1(new_n1003_), .B0(new_n1007_), .B1(new_n1005_), .Y(new_n1009_));
  INV    g00007(.A(\A[720] ), .Y(new_n1010_));
  INV    g00008(.A(\A[718] ), .Y(new_n1011_));
  NAND2  g00009(.A(\A[719] ), .B(new_n1011_), .Y(new_n1012_));
  INV    g00010(.A(\A[719] ), .Y(new_n1013_));
  AOI21  g00011(.A0(new_n1013_), .A1(\A[718] ), .B0(new_n1010_), .Y(new_n1014_));
  XOR2   g00012(.A(\A[719] ), .B(\A[718] ), .Y(new_n1015_));
  AOI22  g00013(.A0(new_n1015_), .A1(new_n1010_), .B0(new_n1014_), .B1(new_n1012_), .Y(new_n1016_));
  NOR2   g00014(.A(new_n1016_), .B(new_n1009_), .Y(new_n1017_));
  NAND2  g00015(.A(\A[719] ), .B(\A[718] ), .Y(new_n1018_));
  NAND2  g00016(.A(new_n1015_), .B(\A[720] ), .Y(new_n1019_));
  NAND2  g00017(.A(new_n1019_), .B(new_n1018_), .Y(new_n1020_));
  NOR2   g00018(.A(new_n1006_), .B(new_n1004_), .Y(new_n1021_));
  AOI21  g00019(.A0(new_n1008_), .A1(\A[717] ), .B0(new_n1021_), .Y(new_n1022_));
  XOR2   g00020(.A(new_n1022_), .B(new_n1020_), .Y(new_n1023_));
  XOR2   g00021(.A(new_n1023_), .B(new_n1017_), .Y(new_n1024_));
  XOR2   g00022(.A(new_n1016_), .B(new_n1009_), .Y(new_n1025_));
  NOR2   g00023(.A(new_n1006_), .B(\A[715] ), .Y(new_n1026_));
  OAI21  g00024(.A0(\A[716] ), .A1(new_n1004_), .B0(\A[717] ), .Y(new_n1027_));
  XOR2   g00025(.A(\A[716] ), .B(new_n1004_), .Y(new_n1028_));
  OAI22  g00026(.A0(new_n1028_), .A1(\A[717] ), .B0(new_n1027_), .B1(new_n1026_), .Y(new_n1029_));
  NOR2   g00027(.A(new_n1013_), .B(\A[718] ), .Y(new_n1030_));
  OAI21  g00028(.A0(\A[719] ), .A1(new_n1011_), .B0(\A[720] ), .Y(new_n1031_));
  XOR2   g00029(.A(\A[719] ), .B(new_n1011_), .Y(new_n1032_));
  OAI22  g00030(.A0(new_n1032_), .A1(\A[720] ), .B0(new_n1031_), .B1(new_n1030_), .Y(new_n1033_));
  NAND2  g00031(.A(new_n1033_), .B(new_n1029_), .Y(new_n1034_));
  NAND2  g00032(.A(\A[716] ), .B(\A[715] ), .Y(new_n1035_));
  OAI21  g00033(.A0(new_n1028_), .A1(new_n1003_), .B0(new_n1035_), .Y(new_n1036_));
  NAND2  g00034(.A(new_n1036_), .B(new_n1020_), .Y(new_n1037_));
  OAI21  g00035(.A0(new_n1023_), .A1(new_n1034_), .B0(new_n1037_), .Y(new_n1038_));
  AOI21  g00036(.A0(new_n1038_), .A1(new_n1025_), .B0(new_n1024_), .Y(new_n1039_));
  INV    g00037(.A(\A[724] ), .Y(new_n1040_));
  INV    g00038(.A(\A[725] ), .Y(new_n1041_));
  XOR2   g00039(.A(\A[725] ), .B(\A[724] ), .Y(new_n1042_));
  NAND2  g00040(.A(new_n1042_), .B(\A[726] ), .Y(new_n1043_));
  OAI21  g00041(.A0(new_n1041_), .A1(new_n1040_), .B0(new_n1043_), .Y(new_n1044_));
  INV    g00042(.A(\A[721] ), .Y(new_n1045_));
  INV    g00043(.A(\A[722] ), .Y(new_n1046_));
  XOR2   g00044(.A(\A[722] ), .B(\A[721] ), .Y(new_n1047_));
  NAND2  g00045(.A(new_n1047_), .B(\A[723] ), .Y(new_n1048_));
  OAI21  g00046(.A0(new_n1046_), .A1(new_n1045_), .B0(new_n1048_), .Y(new_n1049_));
  NOR2   g00047(.A(new_n1046_), .B(\A[721] ), .Y(new_n1050_));
  OAI21  g00048(.A0(\A[722] ), .A1(new_n1045_), .B0(\A[723] ), .Y(new_n1051_));
  INV    g00049(.A(\A[723] ), .Y(new_n1052_));
  NAND2  g00050(.A(new_n1047_), .B(new_n1052_), .Y(new_n1053_));
  OAI21  g00051(.A0(new_n1051_), .A1(new_n1050_), .B0(new_n1053_), .Y(new_n1054_));
  NOR2   g00052(.A(new_n1041_), .B(\A[724] ), .Y(new_n1055_));
  OAI21  g00053(.A0(\A[725] ), .A1(new_n1040_), .B0(\A[726] ), .Y(new_n1056_));
  INV    g00054(.A(\A[726] ), .Y(new_n1057_));
  NAND2  g00055(.A(new_n1042_), .B(new_n1057_), .Y(new_n1058_));
  OAI21  g00056(.A0(new_n1056_), .A1(new_n1055_), .B0(new_n1058_), .Y(new_n1059_));
  NAND4  g00057(.A(new_n1059_), .B(new_n1054_), .C(new_n1049_), .D(new_n1044_), .Y(new_n1060_));
  NAND4  g00058(.A(new_n1036_), .B(new_n1020_), .C(new_n1033_), .D(new_n1029_), .Y(new_n1061_));
  NAND2  g00059(.A(\A[722] ), .B(new_n1045_), .Y(new_n1062_));
  AOI21  g00060(.A0(new_n1046_), .A1(\A[721] ), .B0(new_n1052_), .Y(new_n1063_));
  AOI22  g00061(.A0(new_n1063_), .A1(new_n1062_), .B0(new_n1047_), .B1(new_n1052_), .Y(new_n1064_));
  NAND2  g00062(.A(\A[725] ), .B(new_n1040_), .Y(new_n1065_));
  AOI21  g00063(.A0(new_n1041_), .A1(\A[724] ), .B0(new_n1057_), .Y(new_n1066_));
  AOI22  g00064(.A0(new_n1066_), .A1(new_n1065_), .B0(new_n1042_), .B1(new_n1057_), .Y(new_n1067_));
  XOR2   g00065(.A(new_n1067_), .B(new_n1064_), .Y(new_n1068_));
  NAND4  g00066(.A(new_n1068_), .B(new_n1061_), .C(new_n1060_), .D(new_n1025_), .Y(new_n1069_));
  NOR2   g00067(.A(new_n1046_), .B(new_n1045_), .Y(new_n1070_));
  AOI21  g00068(.A0(new_n1047_), .A1(\A[723] ), .B0(new_n1070_), .Y(new_n1071_));
  XOR2   g00069(.A(new_n1071_), .B(new_n1044_), .Y(new_n1072_));
  NAND2  g00070(.A(new_n1059_), .B(new_n1054_), .Y(new_n1073_));
  NAND2  g00071(.A(new_n1049_), .B(new_n1044_), .Y(new_n1074_));
  OAI21  g00072(.A0(new_n1073_), .A1(new_n1072_), .B0(new_n1074_), .Y(new_n1075_));
  NOR2   g00073(.A(new_n1067_), .B(new_n1064_), .Y(new_n1076_));
  XOR2   g00074(.A(new_n1076_), .B(new_n1072_), .Y(new_n1077_));
  AOI21  g00075(.A0(new_n1068_), .A1(new_n1075_), .B0(new_n1077_), .Y(new_n1078_));
  XOR2   g00076(.A(new_n1078_), .B(new_n1069_), .Y(new_n1079_));
  NOR2   g00077(.A(new_n1079_), .B(new_n1039_), .Y(new_n1080_));
  XOR2   g00078(.A(new_n1023_), .B(new_n1034_), .Y(new_n1081_));
  INV    g00079(.A(new_n1025_), .Y(new_n1082_));
  NOR2   g00080(.A(new_n1023_), .B(new_n1034_), .Y(new_n1083_));
  AOI21  g00081(.A0(new_n1036_), .A1(new_n1020_), .B0(new_n1083_), .Y(new_n1084_));
  OAI21  g00082(.A0(new_n1084_), .A1(new_n1082_), .B0(new_n1081_), .Y(new_n1085_));
  XOR2   g00083(.A(new_n1049_), .B(new_n1044_), .Y(new_n1086_));
  NOR2   g00084(.A(new_n1041_), .B(new_n1040_), .Y(new_n1087_));
  AOI21  g00085(.A0(new_n1042_), .A1(\A[726] ), .B0(new_n1087_), .Y(new_n1088_));
  NOR2   g00086(.A(new_n1071_), .B(new_n1088_), .Y(new_n1089_));
  AOI21  g00087(.A0(new_n1076_), .A1(new_n1086_), .B0(new_n1089_), .Y(new_n1090_));
  XOR2   g00088(.A(new_n1076_), .B(new_n1086_), .Y(new_n1091_));
  XOR2   g00089(.A(new_n1067_), .B(new_n1054_), .Y(new_n1092_));
  OAI21  g00090(.A0(new_n1092_), .A1(new_n1090_), .B0(new_n1091_), .Y(new_n1093_));
  AOI211 g00091(.A0(new_n1019_), .A1(new_n1018_), .B(new_n1022_), .C(new_n1034_), .Y(new_n1094_));
  NAND2  g00092(.A(new_n1068_), .B(new_n1025_), .Y(new_n1095_));
  AOI211 g00093(.A0(new_n1067_), .A1(new_n1064_), .B(new_n1071_), .C(new_n1088_), .Y(new_n1096_));
  NOR4   g00094(.A(new_n1096_), .B(new_n1095_), .C(new_n1094_), .D(new_n1077_), .Y(new_n1097_));
  AOI21  g00095(.A0(new_n1093_), .A1(new_n1069_), .B0(new_n1097_), .Y(new_n1098_));
  NOR2   g00096(.A(new_n1098_), .B(new_n1085_), .Y(new_n1099_));
  NAND2  g00097(.A(new_n1068_), .B(new_n1060_), .Y(new_n1100_));
  NAND2  g00098(.A(new_n1061_), .B(new_n1025_), .Y(new_n1101_));
  XOR2   g00099(.A(new_n1101_), .B(new_n1100_), .Y(new_n1102_));
  INV    g00100(.A(\A[711] ), .Y(new_n1103_));
  INV    g00101(.A(\A[710] ), .Y(new_n1104_));
  NAND2  g00102(.A(new_n1104_), .B(\A[709] ), .Y(new_n1105_));
  INV    g00103(.A(\A[709] ), .Y(new_n1106_));
  AOI21  g00104(.A0(\A[710] ), .A1(new_n1106_), .B0(new_n1103_), .Y(new_n1107_));
  XOR2   g00105(.A(\A[710] ), .B(\A[709] ), .Y(new_n1108_));
  AOI22  g00106(.A0(new_n1108_), .A1(new_n1103_), .B0(new_n1107_), .B1(new_n1105_), .Y(new_n1109_));
  INV    g00107(.A(\A[714] ), .Y(new_n1110_));
  INV    g00108(.A(\A[713] ), .Y(new_n1111_));
  NAND2  g00109(.A(new_n1111_), .B(\A[712] ), .Y(new_n1112_));
  INV    g00110(.A(\A[712] ), .Y(new_n1113_));
  AOI21  g00111(.A0(\A[713] ), .A1(new_n1113_), .B0(new_n1110_), .Y(new_n1114_));
  XOR2   g00112(.A(\A[713] ), .B(\A[712] ), .Y(new_n1115_));
  AOI22  g00113(.A0(new_n1115_), .A1(new_n1110_), .B0(new_n1114_), .B1(new_n1112_), .Y(new_n1116_));
  NOR2   g00114(.A(new_n1111_), .B(new_n1113_), .Y(new_n1117_));
  AOI21  g00115(.A0(new_n1115_), .A1(\A[714] ), .B0(new_n1117_), .Y(new_n1118_));
  NOR2   g00116(.A(new_n1104_), .B(new_n1106_), .Y(new_n1119_));
  AOI21  g00117(.A0(new_n1108_), .A1(\A[711] ), .B0(new_n1119_), .Y(new_n1120_));
  XOR2   g00118(.A(new_n1116_), .B(new_n1109_), .Y(new_n1121_));
  INV    g00119(.A(\A[705] ), .Y(new_n1122_));
  INV    g00120(.A(\A[704] ), .Y(new_n1123_));
  NAND2  g00121(.A(new_n1123_), .B(\A[703] ), .Y(new_n1124_));
  INV    g00122(.A(\A[703] ), .Y(new_n1125_));
  AOI21  g00123(.A0(\A[704] ), .A1(new_n1125_), .B0(new_n1122_), .Y(new_n1126_));
  XOR2   g00124(.A(\A[704] ), .B(\A[703] ), .Y(new_n1127_));
  AOI22  g00125(.A0(new_n1127_), .A1(new_n1122_), .B0(new_n1126_), .B1(new_n1124_), .Y(new_n1128_));
  INV    g00126(.A(\A[708] ), .Y(new_n1129_));
  INV    g00127(.A(\A[707] ), .Y(new_n1130_));
  NAND2  g00128(.A(new_n1130_), .B(\A[706] ), .Y(new_n1131_));
  INV    g00129(.A(\A[706] ), .Y(new_n1132_));
  AOI21  g00130(.A0(\A[707] ), .A1(new_n1132_), .B0(new_n1129_), .Y(new_n1133_));
  XOR2   g00131(.A(\A[707] ), .B(\A[706] ), .Y(new_n1134_));
  AOI22  g00132(.A0(new_n1134_), .A1(new_n1129_), .B0(new_n1133_), .B1(new_n1131_), .Y(new_n1135_));
  NOR2   g00133(.A(new_n1130_), .B(new_n1132_), .Y(new_n1136_));
  AOI21  g00134(.A0(new_n1134_), .A1(\A[708] ), .B0(new_n1136_), .Y(new_n1137_));
  NOR2   g00135(.A(new_n1123_), .B(new_n1125_), .Y(new_n1138_));
  AOI21  g00136(.A0(new_n1127_), .A1(\A[705] ), .B0(new_n1138_), .Y(new_n1139_));
  XOR2   g00137(.A(new_n1135_), .B(new_n1128_), .Y(new_n1140_));
  XOR2   g00138(.A(new_n1140_), .B(new_n1121_), .Y(new_n1141_));
  NAND2  g00139(.A(new_n1141_), .B(new_n1102_), .Y(new_n1142_));
  NOR3   g00140(.A(new_n1142_), .B(new_n1099_), .C(new_n1080_), .Y(new_n1143_));
  NOR4   g00141(.A(new_n1067_), .B(new_n1064_), .C(new_n1071_), .D(new_n1088_), .Y(new_n1144_));
  NOR3   g00142(.A(new_n1095_), .B(new_n1094_), .C(new_n1144_), .Y(new_n1145_));
  XOR2   g00143(.A(new_n1078_), .B(new_n1145_), .Y(new_n1146_));
  NAND2  g00144(.A(new_n1146_), .B(new_n1085_), .Y(new_n1147_));
  NOR2   g00145(.A(new_n1078_), .B(new_n1145_), .Y(new_n1148_));
  OAI21  g00146(.A0(new_n1097_), .A1(new_n1148_), .B0(new_n1039_), .Y(new_n1149_));
  NOR2   g00147(.A(new_n1092_), .B(new_n1144_), .Y(new_n1150_));
  XOR2   g00148(.A(new_n1101_), .B(new_n1150_), .Y(new_n1151_));
  INV    g00149(.A(new_n1141_), .Y(new_n1152_));
  NOR2   g00150(.A(new_n1152_), .B(new_n1151_), .Y(new_n1153_));
  AOI21  g00151(.A0(new_n1149_), .A1(new_n1147_), .B0(new_n1153_), .Y(new_n1154_));
  NOR2   g00152(.A(new_n1154_), .B(new_n1143_), .Y(new_n1155_));
  XOR2   g00153(.A(new_n1135_), .B(new_n1128_), .Y(new_n1156_));
  XOR2   g00154(.A(new_n1139_), .B(new_n1137_), .Y(new_n1157_));
  NOR2   g00155(.A(new_n1135_), .B(new_n1128_), .Y(new_n1158_));
  NAND2  g00156(.A(new_n1158_), .B(new_n1157_), .Y(new_n1159_));
  OAI21  g00157(.A0(new_n1139_), .A1(new_n1137_), .B0(new_n1159_), .Y(new_n1160_));
  INV    g00158(.A(new_n1134_), .Y(new_n1161_));
  NAND2  g00159(.A(\A[707] ), .B(\A[706] ), .Y(new_n1162_));
  OAI21  g00160(.A0(new_n1161_), .A1(new_n1129_), .B0(new_n1162_), .Y(new_n1163_));
  XOR2   g00161(.A(new_n1139_), .B(new_n1163_), .Y(new_n1164_));
  XOR2   g00162(.A(new_n1158_), .B(new_n1164_), .Y(new_n1165_));
  AOI21  g00163(.A0(new_n1160_), .A1(new_n1156_), .B0(new_n1165_), .Y(new_n1166_));
  XOR2   g00164(.A(new_n1116_), .B(new_n1109_), .Y(new_n1167_));
  NOR2   g00165(.A(\A[710] ), .B(new_n1106_), .Y(new_n1168_));
  OAI21  g00166(.A0(new_n1104_), .A1(\A[709] ), .B0(\A[711] ), .Y(new_n1169_));
  NAND2  g00167(.A(new_n1108_), .B(new_n1103_), .Y(new_n1170_));
  OAI21  g00168(.A0(new_n1169_), .A1(new_n1168_), .B0(new_n1170_), .Y(new_n1171_));
  NOR2   g00169(.A(\A[713] ), .B(new_n1113_), .Y(new_n1172_));
  OAI21  g00170(.A0(new_n1111_), .A1(\A[712] ), .B0(\A[714] ), .Y(new_n1173_));
  NAND2  g00171(.A(new_n1115_), .B(new_n1110_), .Y(new_n1174_));
  OAI21  g00172(.A0(new_n1173_), .A1(new_n1172_), .B0(new_n1174_), .Y(new_n1175_));
  NAND2  g00173(.A(new_n1115_), .B(\A[714] ), .Y(new_n1176_));
  OAI21  g00174(.A0(new_n1111_), .A1(new_n1113_), .B0(new_n1176_), .Y(new_n1177_));
  NAND2  g00175(.A(new_n1108_), .B(\A[711] ), .Y(new_n1178_));
  OAI21  g00176(.A0(new_n1104_), .A1(new_n1106_), .B0(new_n1178_), .Y(new_n1179_));
  NAND4  g00177(.A(new_n1179_), .B(new_n1177_), .C(new_n1175_), .D(new_n1171_), .Y(new_n1180_));
  INV    g00178(.A(new_n1127_), .Y(new_n1181_));
  NOR2   g00179(.A(new_n1181_), .B(new_n1122_), .Y(new_n1182_));
  OAI211 g00180(.A0(new_n1182_), .A1(new_n1138_), .B0(new_n1158_), .B1(new_n1163_), .Y(new_n1183_));
  NAND4  g00181(.A(new_n1183_), .B(new_n1156_), .C(new_n1180_), .D(new_n1167_), .Y(new_n1184_));
  XOR2   g00182(.A(new_n1120_), .B(new_n1177_), .Y(new_n1185_));
  NAND2  g00183(.A(new_n1175_), .B(new_n1171_), .Y(new_n1186_));
  NAND2  g00184(.A(new_n1179_), .B(new_n1177_), .Y(new_n1187_));
  OAI21  g00185(.A0(new_n1186_), .A1(new_n1185_), .B0(new_n1187_), .Y(new_n1188_));
  NOR2   g00186(.A(new_n1116_), .B(new_n1109_), .Y(new_n1189_));
  XOR2   g00187(.A(new_n1189_), .B(new_n1185_), .Y(new_n1190_));
  AOI21  g00188(.A0(new_n1188_), .A1(new_n1167_), .B0(new_n1190_), .Y(new_n1191_));
  XOR2   g00189(.A(new_n1191_), .B(new_n1184_), .Y(new_n1192_));
  XOR2   g00190(.A(new_n1116_), .B(new_n1171_), .Y(new_n1193_));
  XOR2   g00191(.A(new_n1120_), .B(new_n1118_), .Y(new_n1194_));
  NOR2   g00192(.A(new_n1120_), .B(new_n1118_), .Y(new_n1195_));
  AOI21  g00193(.A0(new_n1189_), .A1(new_n1194_), .B0(new_n1195_), .Y(new_n1196_));
  XOR2   g00194(.A(new_n1189_), .B(new_n1194_), .Y(new_n1197_));
  OAI21  g00195(.A0(new_n1196_), .A1(new_n1193_), .B0(new_n1197_), .Y(new_n1198_));
  NAND2  g00196(.A(new_n1198_), .B(new_n1184_), .Y(new_n1199_));
  NAND2  g00197(.A(new_n1126_), .B(new_n1124_), .Y(new_n1200_));
  OAI21  g00198(.A0(new_n1181_), .A1(\A[705] ), .B0(new_n1200_), .Y(new_n1201_));
  XOR2   g00199(.A(new_n1135_), .B(new_n1201_), .Y(new_n1202_));
  NOR4   g00200(.A(new_n1202_), .B(new_n1190_), .C(new_n1188_), .D(new_n1193_), .Y(new_n1203_));
  OAI211 g00201(.A0(new_n1196_), .A1(new_n1193_), .B0(new_n1203_), .B1(new_n1183_), .Y(new_n1204_));
  NAND2  g00202(.A(new_n1204_), .B(new_n1199_), .Y(new_n1205_));
  NAND2  g00203(.A(new_n1205_), .B(new_n1166_), .Y(new_n1206_));
  OAI21  g00204(.A0(new_n1192_), .A1(new_n1166_), .B0(new_n1206_), .Y(new_n1207_));
  NOR2   g00205(.A(new_n1207_), .B(new_n1155_), .Y(new_n1208_));
  NOR2   g00206(.A(new_n1192_), .B(new_n1166_), .Y(new_n1209_));
  NOR2   g00207(.A(new_n1139_), .B(new_n1137_), .Y(new_n1210_));
  AOI21  g00208(.A0(new_n1158_), .A1(new_n1157_), .B0(new_n1210_), .Y(new_n1211_));
  XOR2   g00209(.A(new_n1158_), .B(new_n1157_), .Y(new_n1212_));
  OAI21  g00210(.A0(new_n1211_), .A1(new_n1202_), .B0(new_n1212_), .Y(new_n1213_));
  AOI21  g00211(.A0(new_n1204_), .A1(new_n1199_), .B0(new_n1213_), .Y(new_n1214_));
  NOR2   g00212(.A(new_n1214_), .B(new_n1209_), .Y(new_n1215_));
  NAND3  g00213(.A(new_n1142_), .B(new_n1149_), .C(new_n1147_), .Y(new_n1216_));
  OAI21  g00214(.A0(new_n1099_), .A1(new_n1080_), .B0(new_n1153_), .Y(new_n1217_));
  AOI21  g00215(.A0(new_n1217_), .A1(new_n1216_), .B0(new_n1215_), .Y(new_n1218_));
  NOR2   g00216(.A(new_n1218_), .B(new_n1208_), .Y(new_n1219_));
  INV    g00217(.A(\A[729] ), .Y(new_n1220_));
  INV    g00218(.A(\A[727] ), .Y(new_n1221_));
  NAND2  g00219(.A(\A[728] ), .B(new_n1221_), .Y(new_n1222_));
  INV    g00220(.A(\A[728] ), .Y(new_n1223_));
  AOI21  g00221(.A0(new_n1223_), .A1(\A[727] ), .B0(new_n1220_), .Y(new_n1224_));
  XOR2   g00222(.A(\A[728] ), .B(\A[727] ), .Y(new_n1225_));
  AOI22  g00223(.A0(new_n1225_), .A1(new_n1220_), .B0(new_n1224_), .B1(new_n1222_), .Y(new_n1226_));
  INV    g00224(.A(\A[732] ), .Y(new_n1227_));
  INV    g00225(.A(\A[730] ), .Y(new_n1228_));
  NAND2  g00226(.A(\A[731] ), .B(new_n1228_), .Y(new_n1229_));
  INV    g00227(.A(\A[731] ), .Y(new_n1230_));
  AOI21  g00228(.A0(new_n1230_), .A1(\A[730] ), .B0(new_n1227_), .Y(new_n1231_));
  XOR2   g00229(.A(\A[731] ), .B(\A[730] ), .Y(new_n1232_));
  AOI22  g00230(.A0(new_n1232_), .A1(new_n1227_), .B0(new_n1231_), .B1(new_n1229_), .Y(new_n1233_));
  NOR2   g00231(.A(new_n1233_), .B(new_n1226_), .Y(new_n1234_));
  NAND2  g00232(.A(\A[731] ), .B(\A[730] ), .Y(new_n1235_));
  NAND2  g00233(.A(new_n1232_), .B(\A[732] ), .Y(new_n1236_));
  NAND2  g00234(.A(new_n1236_), .B(new_n1235_), .Y(new_n1237_));
  NOR2   g00235(.A(new_n1223_), .B(new_n1221_), .Y(new_n1238_));
  AOI21  g00236(.A0(new_n1225_), .A1(\A[729] ), .B0(new_n1238_), .Y(new_n1239_));
  XOR2   g00237(.A(new_n1239_), .B(new_n1237_), .Y(new_n1240_));
  XOR2   g00238(.A(new_n1240_), .B(new_n1234_), .Y(new_n1241_));
  XOR2   g00239(.A(new_n1233_), .B(new_n1226_), .Y(new_n1242_));
  NOR2   g00240(.A(new_n1223_), .B(\A[727] ), .Y(new_n1243_));
  OAI21  g00241(.A0(\A[728] ), .A1(new_n1221_), .B0(\A[729] ), .Y(new_n1244_));
  XOR2   g00242(.A(\A[728] ), .B(new_n1221_), .Y(new_n1245_));
  OAI22  g00243(.A0(new_n1245_), .A1(\A[729] ), .B0(new_n1244_), .B1(new_n1243_), .Y(new_n1246_));
  NOR2   g00244(.A(new_n1230_), .B(\A[730] ), .Y(new_n1247_));
  OAI21  g00245(.A0(\A[731] ), .A1(new_n1228_), .B0(\A[732] ), .Y(new_n1248_));
  XOR2   g00246(.A(\A[731] ), .B(new_n1228_), .Y(new_n1249_));
  OAI22  g00247(.A0(new_n1249_), .A1(\A[732] ), .B0(new_n1248_), .B1(new_n1247_), .Y(new_n1250_));
  NAND2  g00248(.A(new_n1250_), .B(new_n1246_), .Y(new_n1251_));
  NAND2  g00249(.A(\A[728] ), .B(\A[727] ), .Y(new_n1252_));
  OAI21  g00250(.A0(new_n1245_), .A1(new_n1220_), .B0(new_n1252_), .Y(new_n1253_));
  NAND2  g00251(.A(new_n1253_), .B(new_n1237_), .Y(new_n1254_));
  OAI21  g00252(.A0(new_n1240_), .A1(new_n1251_), .B0(new_n1254_), .Y(new_n1255_));
  AOI21  g00253(.A0(new_n1255_), .A1(new_n1242_), .B0(new_n1241_), .Y(new_n1256_));
  NAND2  g00254(.A(\A[737] ), .B(\A[736] ), .Y(new_n1257_));
  XOR2   g00255(.A(\A[737] ), .B(\A[736] ), .Y(new_n1258_));
  NAND2  g00256(.A(new_n1258_), .B(\A[738] ), .Y(new_n1259_));
  NAND2  g00257(.A(new_n1259_), .B(new_n1257_), .Y(new_n1260_));
  INV    g00258(.A(\A[733] ), .Y(new_n1261_));
  INV    g00259(.A(\A[734] ), .Y(new_n1262_));
  XOR2   g00260(.A(\A[734] ), .B(\A[733] ), .Y(new_n1263_));
  NAND2  g00261(.A(new_n1263_), .B(\A[735] ), .Y(new_n1264_));
  OAI21  g00262(.A0(new_n1262_), .A1(new_n1261_), .B0(new_n1264_), .Y(new_n1265_));
  NOR2   g00263(.A(new_n1262_), .B(\A[733] ), .Y(new_n1266_));
  OAI21  g00264(.A0(\A[734] ), .A1(new_n1261_), .B0(\A[735] ), .Y(new_n1267_));
  INV    g00265(.A(\A[735] ), .Y(new_n1268_));
  NAND2  g00266(.A(new_n1263_), .B(new_n1268_), .Y(new_n1269_));
  OAI21  g00267(.A0(new_n1267_), .A1(new_n1266_), .B0(new_n1269_), .Y(new_n1270_));
  INV    g00268(.A(\A[737] ), .Y(new_n1271_));
  NOR2   g00269(.A(new_n1271_), .B(\A[736] ), .Y(new_n1272_));
  INV    g00270(.A(\A[736] ), .Y(new_n1273_));
  OAI21  g00271(.A0(\A[737] ), .A1(new_n1273_), .B0(\A[738] ), .Y(new_n1274_));
  INV    g00272(.A(\A[738] ), .Y(new_n1275_));
  NAND2  g00273(.A(new_n1258_), .B(new_n1275_), .Y(new_n1276_));
  OAI21  g00274(.A0(new_n1274_), .A1(new_n1272_), .B0(new_n1276_), .Y(new_n1277_));
  NAND4  g00275(.A(new_n1277_), .B(new_n1270_), .C(new_n1265_), .D(new_n1260_), .Y(new_n1278_));
  NAND4  g00276(.A(new_n1253_), .B(new_n1237_), .C(new_n1250_), .D(new_n1246_), .Y(new_n1279_));
  NAND2  g00277(.A(\A[734] ), .B(new_n1261_), .Y(new_n1280_));
  AOI21  g00278(.A0(new_n1262_), .A1(\A[733] ), .B0(new_n1268_), .Y(new_n1281_));
  AOI22  g00279(.A0(new_n1281_), .A1(new_n1280_), .B0(new_n1263_), .B1(new_n1268_), .Y(new_n1282_));
  NAND2  g00280(.A(\A[737] ), .B(new_n1273_), .Y(new_n1283_));
  AOI21  g00281(.A0(new_n1271_), .A1(\A[736] ), .B0(new_n1275_), .Y(new_n1284_));
  AOI22  g00282(.A0(new_n1284_), .A1(new_n1283_), .B0(new_n1258_), .B1(new_n1275_), .Y(new_n1285_));
  XOR2   g00283(.A(new_n1285_), .B(new_n1282_), .Y(new_n1286_));
  NAND4  g00284(.A(new_n1286_), .B(new_n1279_), .C(new_n1278_), .D(new_n1242_), .Y(new_n1287_));
  NOR2   g00285(.A(new_n1262_), .B(new_n1261_), .Y(new_n1288_));
  AOI21  g00286(.A0(new_n1263_), .A1(\A[735] ), .B0(new_n1288_), .Y(new_n1289_));
  XOR2   g00287(.A(new_n1289_), .B(new_n1260_), .Y(new_n1290_));
  NAND2  g00288(.A(new_n1277_), .B(new_n1270_), .Y(new_n1291_));
  NAND2  g00289(.A(new_n1265_), .B(new_n1260_), .Y(new_n1292_));
  OAI21  g00290(.A0(new_n1291_), .A1(new_n1290_), .B0(new_n1292_), .Y(new_n1293_));
  NOR2   g00291(.A(new_n1285_), .B(new_n1282_), .Y(new_n1294_));
  XOR2   g00292(.A(new_n1294_), .B(new_n1290_), .Y(new_n1295_));
  AOI21  g00293(.A0(new_n1286_), .A1(new_n1293_), .B0(new_n1295_), .Y(new_n1296_));
  XOR2   g00294(.A(new_n1296_), .B(new_n1287_), .Y(new_n1297_));
  XOR2   g00295(.A(new_n1265_), .B(new_n1260_), .Y(new_n1298_));
  XOR2   g00296(.A(new_n1294_), .B(new_n1298_), .Y(new_n1299_));
  AOI211 g00297(.A0(new_n1236_), .A1(new_n1235_), .B(new_n1239_), .C(new_n1251_), .Y(new_n1300_));
  NAND2  g00298(.A(new_n1286_), .B(new_n1242_), .Y(new_n1301_));
  AOI211 g00299(.A0(new_n1299_), .A1(new_n1293_), .B(new_n1301_), .C(new_n1300_), .Y(new_n1302_));
  NOR2   g00300(.A(new_n1296_), .B(new_n1302_), .Y(new_n1303_));
  AOI221 g00301(.A0(new_n1285_), .A1(new_n1282_), .C0(new_n1289_), .B0(new_n1259_), .B1(new_n1257_), .Y(new_n1304_));
  NOR4   g00302(.A(new_n1304_), .B(new_n1301_), .C(new_n1300_), .D(new_n1295_), .Y(new_n1305_));
  OAI21  g00303(.A0(new_n1305_), .A1(new_n1303_), .B0(new_n1256_), .Y(new_n1306_));
  OAI21  g00304(.A0(new_n1297_), .A1(new_n1256_), .B0(new_n1306_), .Y(new_n1307_));
  INV    g00305(.A(\A[740] ), .Y(new_n1308_));
  NOR2   g00306(.A(new_n1308_), .B(\A[739] ), .Y(new_n1309_));
  INV    g00307(.A(\A[739] ), .Y(new_n1310_));
  OAI21  g00308(.A0(\A[740] ), .A1(new_n1310_), .B0(\A[741] ), .Y(new_n1311_));
  XOR2   g00309(.A(\A[740] ), .B(new_n1310_), .Y(new_n1312_));
  OAI22  g00310(.A0(new_n1312_), .A1(\A[741] ), .B0(new_n1311_), .B1(new_n1309_), .Y(new_n1313_));
  INV    g00311(.A(\A[743] ), .Y(new_n1314_));
  NOR2   g00312(.A(new_n1314_), .B(\A[742] ), .Y(new_n1315_));
  INV    g00313(.A(\A[742] ), .Y(new_n1316_));
  OAI21  g00314(.A0(\A[743] ), .A1(new_n1316_), .B0(\A[744] ), .Y(new_n1317_));
  XOR2   g00315(.A(\A[743] ), .B(new_n1316_), .Y(new_n1318_));
  OAI22  g00316(.A0(new_n1318_), .A1(\A[744] ), .B0(new_n1317_), .B1(new_n1315_), .Y(new_n1319_));
  NAND2  g00317(.A(new_n1319_), .B(new_n1313_), .Y(new_n1320_));
  NAND2  g00318(.A(\A[743] ), .B(\A[742] ), .Y(new_n1321_));
  XOR2   g00319(.A(\A[743] ), .B(\A[742] ), .Y(new_n1322_));
  NAND2  g00320(.A(new_n1322_), .B(\A[744] ), .Y(new_n1323_));
  NAND2  g00321(.A(new_n1323_), .B(new_n1321_), .Y(new_n1324_));
  XOR2   g00322(.A(\A[740] ), .B(\A[739] ), .Y(new_n1325_));
  NOR2   g00323(.A(new_n1308_), .B(new_n1310_), .Y(new_n1326_));
  AOI21  g00324(.A0(new_n1325_), .A1(\A[741] ), .B0(new_n1326_), .Y(new_n1327_));
  XOR2   g00325(.A(new_n1327_), .B(new_n1324_), .Y(new_n1328_));
  XOR2   g00326(.A(new_n1328_), .B(new_n1320_), .Y(new_n1329_));
  INV    g00327(.A(\A[741] ), .Y(new_n1330_));
  NAND2  g00328(.A(\A[740] ), .B(new_n1310_), .Y(new_n1331_));
  AOI21  g00329(.A0(new_n1308_), .A1(\A[739] ), .B0(new_n1330_), .Y(new_n1332_));
  AOI22  g00330(.A0(new_n1325_), .A1(new_n1330_), .B0(new_n1332_), .B1(new_n1331_), .Y(new_n1333_));
  INV    g00331(.A(\A[744] ), .Y(new_n1334_));
  NAND2  g00332(.A(\A[743] ), .B(new_n1316_), .Y(new_n1335_));
  AOI21  g00333(.A0(new_n1314_), .A1(\A[742] ), .B0(new_n1334_), .Y(new_n1336_));
  AOI22  g00334(.A0(new_n1322_), .A1(new_n1334_), .B0(new_n1336_), .B1(new_n1335_), .Y(new_n1337_));
  XOR2   g00335(.A(new_n1337_), .B(new_n1333_), .Y(new_n1338_));
  INV    g00336(.A(new_n1338_), .Y(new_n1339_));
  NAND2  g00337(.A(\A[740] ), .B(\A[739] ), .Y(new_n1340_));
  OAI21  g00338(.A0(new_n1312_), .A1(new_n1330_), .B0(new_n1340_), .Y(new_n1341_));
  NOR2   g00339(.A(new_n1328_), .B(new_n1320_), .Y(new_n1342_));
  AOI21  g00340(.A0(new_n1341_), .A1(new_n1324_), .B0(new_n1342_), .Y(new_n1343_));
  OAI21  g00341(.A0(new_n1343_), .A1(new_n1339_), .B0(new_n1329_), .Y(new_n1344_));
  INV    g00342(.A(\A[748] ), .Y(new_n1345_));
  INV    g00343(.A(\A[749] ), .Y(new_n1346_));
  NOR2   g00344(.A(new_n1346_), .B(new_n1345_), .Y(new_n1347_));
  XOR2   g00345(.A(\A[749] ), .B(\A[748] ), .Y(new_n1348_));
  AOI21  g00346(.A0(new_n1348_), .A1(\A[750] ), .B0(new_n1347_), .Y(new_n1349_));
  INV    g00347(.A(\A[745] ), .Y(new_n1350_));
  INV    g00348(.A(\A[746] ), .Y(new_n1351_));
  NOR2   g00349(.A(new_n1351_), .B(new_n1350_), .Y(new_n1352_));
  XOR2   g00350(.A(\A[746] ), .B(\A[745] ), .Y(new_n1353_));
  AOI21  g00351(.A0(new_n1353_), .A1(\A[747] ), .B0(new_n1352_), .Y(new_n1354_));
  INV    g00352(.A(\A[747] ), .Y(new_n1355_));
  NAND2  g00353(.A(\A[746] ), .B(new_n1350_), .Y(new_n1356_));
  AOI21  g00354(.A0(new_n1351_), .A1(\A[745] ), .B0(new_n1355_), .Y(new_n1357_));
  AOI22  g00355(.A0(new_n1357_), .A1(new_n1356_), .B0(new_n1353_), .B1(new_n1355_), .Y(new_n1358_));
  INV    g00356(.A(\A[750] ), .Y(new_n1359_));
  NAND2  g00357(.A(\A[749] ), .B(new_n1345_), .Y(new_n1360_));
  AOI21  g00358(.A0(new_n1346_), .A1(\A[748] ), .B0(new_n1359_), .Y(new_n1361_));
  AOI22  g00359(.A0(new_n1361_), .A1(new_n1360_), .B0(new_n1348_), .B1(new_n1359_), .Y(new_n1362_));
  NOR4   g00360(.A(new_n1362_), .B(new_n1358_), .C(new_n1354_), .D(new_n1349_), .Y(new_n1363_));
  AOI211 g00361(.A0(new_n1323_), .A1(new_n1321_), .B(new_n1327_), .C(new_n1320_), .Y(new_n1364_));
  XOR2   g00362(.A(new_n1362_), .B(new_n1358_), .Y(new_n1365_));
  NAND2  g00363(.A(new_n1365_), .B(new_n1338_), .Y(new_n1366_));
  NOR3   g00364(.A(new_n1366_), .B(new_n1364_), .C(new_n1363_), .Y(new_n1367_));
  NAND2  g00365(.A(new_n1348_), .B(\A[750] ), .Y(new_n1368_));
  OAI21  g00366(.A0(new_n1346_), .A1(new_n1345_), .B0(new_n1368_), .Y(new_n1369_));
  XOR2   g00367(.A(new_n1354_), .B(new_n1369_), .Y(new_n1370_));
  NOR2   g00368(.A(new_n1351_), .B(\A[745] ), .Y(new_n1371_));
  OAI21  g00369(.A0(\A[746] ), .A1(new_n1350_), .B0(\A[747] ), .Y(new_n1372_));
  NAND2  g00370(.A(new_n1353_), .B(new_n1355_), .Y(new_n1373_));
  OAI21  g00371(.A0(new_n1372_), .A1(new_n1371_), .B0(new_n1373_), .Y(new_n1374_));
  NOR2   g00372(.A(new_n1346_), .B(\A[748] ), .Y(new_n1375_));
  OAI21  g00373(.A0(\A[749] ), .A1(new_n1345_), .B0(\A[750] ), .Y(new_n1376_));
  NAND2  g00374(.A(new_n1348_), .B(new_n1359_), .Y(new_n1377_));
  OAI21  g00375(.A0(new_n1376_), .A1(new_n1375_), .B0(new_n1377_), .Y(new_n1378_));
  NAND2  g00376(.A(new_n1378_), .B(new_n1374_), .Y(new_n1379_));
  NAND2  g00377(.A(new_n1353_), .B(\A[747] ), .Y(new_n1380_));
  OAI21  g00378(.A0(new_n1351_), .A1(new_n1350_), .B0(new_n1380_), .Y(new_n1381_));
  NAND2  g00379(.A(new_n1381_), .B(new_n1369_), .Y(new_n1382_));
  OAI21  g00380(.A0(new_n1379_), .A1(new_n1370_), .B0(new_n1382_), .Y(new_n1383_));
  NOR2   g00381(.A(new_n1362_), .B(new_n1358_), .Y(new_n1384_));
  XOR2   g00382(.A(new_n1384_), .B(new_n1370_), .Y(new_n1385_));
  AOI21  g00383(.A0(new_n1365_), .A1(new_n1383_), .B0(new_n1385_), .Y(new_n1386_));
  XOR2   g00384(.A(new_n1386_), .B(new_n1367_), .Y(new_n1387_));
  NAND2  g00385(.A(new_n1387_), .B(new_n1344_), .Y(new_n1388_));
  NOR2   g00386(.A(new_n1337_), .B(new_n1333_), .Y(new_n1389_));
  XOR2   g00387(.A(new_n1328_), .B(new_n1389_), .Y(new_n1390_));
  NAND2  g00388(.A(new_n1341_), .B(new_n1324_), .Y(new_n1391_));
  OAI21  g00389(.A0(new_n1328_), .A1(new_n1320_), .B0(new_n1391_), .Y(new_n1392_));
  AOI21  g00390(.A0(new_n1392_), .A1(new_n1338_), .B0(new_n1390_), .Y(new_n1393_));
  NOR2   g00391(.A(new_n1386_), .B(new_n1367_), .Y(new_n1394_));
  AOI211 g00392(.A0(new_n1362_), .A1(new_n1358_), .B(new_n1354_), .C(new_n1349_), .Y(new_n1395_));
  NOR4   g00393(.A(new_n1395_), .B(new_n1366_), .C(new_n1364_), .D(new_n1385_), .Y(new_n1396_));
  OAI21  g00394(.A0(new_n1396_), .A1(new_n1394_), .B0(new_n1393_), .Y(new_n1397_));
  XOR2   g00395(.A(new_n1362_), .B(new_n1374_), .Y(new_n1398_));
  NOR2   g00396(.A(new_n1398_), .B(new_n1363_), .Y(new_n1399_));
  NAND4  g00397(.A(new_n1341_), .B(new_n1324_), .C(new_n1319_), .D(new_n1313_), .Y(new_n1400_));
  NAND2  g00398(.A(new_n1400_), .B(new_n1338_), .Y(new_n1401_));
  XOR2   g00399(.A(new_n1401_), .B(new_n1399_), .Y(new_n1402_));
  NAND2  g00400(.A(new_n1286_), .B(new_n1278_), .Y(new_n1403_));
  NAND3  g00401(.A(new_n1403_), .B(new_n1279_), .C(new_n1242_), .Y(new_n1404_));
  NAND2  g00402(.A(new_n1279_), .B(new_n1242_), .Y(new_n1405_));
  NAND3  g00403(.A(new_n1405_), .B(new_n1286_), .C(new_n1278_), .Y(new_n1406_));
  AOI21  g00404(.A0(new_n1406_), .A1(new_n1404_), .B0(new_n1402_), .Y(new_n1407_));
  NAND3  g00405(.A(new_n1407_), .B(new_n1397_), .C(new_n1388_), .Y(new_n1408_));
  NAND4  g00406(.A(new_n1378_), .B(new_n1374_), .C(new_n1381_), .D(new_n1369_), .Y(new_n1409_));
  NAND4  g00407(.A(new_n1365_), .B(new_n1400_), .C(new_n1409_), .D(new_n1338_), .Y(new_n1410_));
  XOR2   g00408(.A(new_n1386_), .B(new_n1410_), .Y(new_n1411_));
  NOR2   g00409(.A(new_n1411_), .B(new_n1393_), .Y(new_n1412_));
  XOR2   g00410(.A(new_n1381_), .B(new_n1369_), .Y(new_n1413_));
  NOR2   g00411(.A(new_n1354_), .B(new_n1349_), .Y(new_n1414_));
  AOI21  g00412(.A0(new_n1384_), .A1(new_n1413_), .B0(new_n1414_), .Y(new_n1415_));
  XOR2   g00413(.A(new_n1384_), .B(new_n1413_), .Y(new_n1416_));
  OAI21  g00414(.A0(new_n1398_), .A1(new_n1415_), .B0(new_n1416_), .Y(new_n1417_));
  AOI21  g00415(.A0(new_n1417_), .A1(new_n1410_), .B0(new_n1396_), .Y(new_n1418_));
  NOR2   g00416(.A(new_n1418_), .B(new_n1344_), .Y(new_n1419_));
  NAND2  g00417(.A(new_n1365_), .B(new_n1409_), .Y(new_n1420_));
  XOR2   g00418(.A(new_n1401_), .B(new_n1420_), .Y(new_n1421_));
  XOR2   g00419(.A(new_n1405_), .B(new_n1403_), .Y(new_n1422_));
  NAND2  g00420(.A(new_n1422_), .B(new_n1421_), .Y(new_n1423_));
  OAI21  g00421(.A0(new_n1419_), .A1(new_n1412_), .B0(new_n1423_), .Y(new_n1424_));
  AOI21  g00422(.A0(new_n1424_), .A1(new_n1408_), .B0(new_n1307_), .Y(new_n1425_));
  NOR2   g00423(.A(new_n1297_), .B(new_n1256_), .Y(new_n1426_));
  AOI21  g00424(.A0(new_n1259_), .A1(new_n1257_), .B0(new_n1289_), .Y(new_n1427_));
  AOI21  g00425(.A0(new_n1294_), .A1(new_n1298_), .B0(new_n1427_), .Y(new_n1428_));
  XOR2   g00426(.A(new_n1285_), .B(new_n1270_), .Y(new_n1429_));
  OAI21  g00427(.A0(new_n1429_), .A1(new_n1428_), .B0(new_n1299_), .Y(new_n1430_));
  AOI21  g00428(.A0(new_n1430_), .A1(new_n1287_), .B0(new_n1305_), .Y(new_n1431_));
  AOI211 g00429(.A0(new_n1255_), .A1(new_n1242_), .B(new_n1431_), .C(new_n1241_), .Y(new_n1432_));
  NOR2   g00430(.A(new_n1432_), .B(new_n1426_), .Y(new_n1433_));
  NAND3  g00431(.A(new_n1423_), .B(new_n1397_), .C(new_n1388_), .Y(new_n1434_));
  OAI21  g00432(.A0(new_n1419_), .A1(new_n1412_), .B0(new_n1407_), .Y(new_n1435_));
  AOI21  g00433(.A0(new_n1435_), .A1(new_n1434_), .B0(new_n1433_), .Y(new_n1436_));
  XOR2   g00434(.A(new_n1422_), .B(new_n1402_), .Y(new_n1437_));
  XOR2   g00435(.A(new_n1152_), .B(new_n1102_), .Y(new_n1438_));
  NOR2   g00436(.A(new_n1438_), .B(new_n1437_), .Y(new_n1439_));
  INV    g00437(.A(new_n1439_), .Y(new_n1440_));
  NOR3   g00438(.A(new_n1440_), .B(new_n1436_), .C(new_n1425_), .Y(new_n1441_));
  NAND2  g00439(.A(new_n1424_), .B(new_n1408_), .Y(new_n1442_));
  NAND2  g00440(.A(new_n1442_), .B(new_n1433_), .Y(new_n1443_));
  NAND2  g00441(.A(new_n1435_), .B(new_n1434_), .Y(new_n1444_));
  NAND2  g00442(.A(new_n1444_), .B(new_n1307_), .Y(new_n1445_));
  AOI21  g00443(.A0(new_n1445_), .A1(new_n1443_), .B0(new_n1439_), .Y(new_n1446_));
  OAI21  g00444(.A0(new_n1446_), .A1(new_n1441_), .B0(new_n1219_), .Y(new_n1447_));
  OAI21  g00445(.A0(new_n1154_), .A1(new_n1143_), .B0(new_n1215_), .Y(new_n1448_));
  OAI21  g00446(.A0(new_n1098_), .A1(new_n1085_), .B0(new_n1142_), .Y(new_n1449_));
  NOR2   g00447(.A(new_n1449_), .B(new_n1080_), .Y(new_n1450_));
  AOI21  g00448(.A0(new_n1149_), .A1(new_n1147_), .B0(new_n1142_), .Y(new_n1451_));
  OAI22  g00449(.A0(new_n1451_), .A1(new_n1450_), .B0(new_n1214_), .B1(new_n1209_), .Y(new_n1452_));
  NAND2  g00450(.A(new_n1452_), .B(new_n1448_), .Y(new_n1453_));
  NOR3   g00451(.A(new_n1439_), .B(new_n1436_), .C(new_n1425_), .Y(new_n1454_));
  AOI21  g00452(.A0(new_n1445_), .A1(new_n1443_), .B0(new_n1440_), .Y(new_n1455_));
  OAI21  g00453(.A0(new_n1455_), .A1(new_n1454_), .B0(new_n1453_), .Y(new_n1456_));
  XOR2   g00454(.A(new_n1438_), .B(new_n1437_), .Y(new_n1457_));
  INV    g00455(.A(new_n1457_), .Y(new_n1458_));
  INV    g00456(.A(\A[699] ), .Y(new_n1459_));
  INV    g00457(.A(\A[698] ), .Y(new_n1460_));
  NAND2  g00458(.A(new_n1460_), .B(\A[697] ), .Y(new_n1461_));
  INV    g00459(.A(\A[697] ), .Y(new_n1462_));
  AOI21  g00460(.A0(\A[698] ), .A1(new_n1462_), .B0(new_n1459_), .Y(new_n1463_));
  XOR2   g00461(.A(\A[698] ), .B(\A[697] ), .Y(new_n1464_));
  AOI22  g00462(.A0(new_n1464_), .A1(new_n1459_), .B0(new_n1463_), .B1(new_n1461_), .Y(new_n1465_));
  INV    g00463(.A(\A[702] ), .Y(new_n1466_));
  INV    g00464(.A(\A[701] ), .Y(new_n1467_));
  NAND2  g00465(.A(new_n1467_), .B(\A[700] ), .Y(new_n1468_));
  INV    g00466(.A(\A[700] ), .Y(new_n1469_));
  AOI21  g00467(.A0(\A[701] ), .A1(new_n1469_), .B0(new_n1466_), .Y(new_n1470_));
  XOR2   g00468(.A(\A[701] ), .B(\A[700] ), .Y(new_n1471_));
  AOI22  g00469(.A0(new_n1471_), .A1(new_n1466_), .B0(new_n1470_), .B1(new_n1468_), .Y(new_n1472_));
  NOR2   g00470(.A(new_n1467_), .B(new_n1469_), .Y(new_n1473_));
  AOI21  g00471(.A0(new_n1471_), .A1(\A[702] ), .B0(new_n1473_), .Y(new_n1474_));
  NOR2   g00472(.A(new_n1460_), .B(new_n1462_), .Y(new_n1475_));
  AOI21  g00473(.A0(new_n1464_), .A1(\A[699] ), .B0(new_n1475_), .Y(new_n1476_));
  XOR2   g00474(.A(new_n1472_), .B(new_n1465_), .Y(new_n1477_));
  INV    g00475(.A(\A[693] ), .Y(new_n1478_));
  INV    g00476(.A(\A[692] ), .Y(new_n1479_));
  NAND2  g00477(.A(new_n1479_), .B(\A[691] ), .Y(new_n1480_));
  INV    g00478(.A(\A[691] ), .Y(new_n1481_));
  AOI21  g00479(.A0(\A[692] ), .A1(new_n1481_), .B0(new_n1478_), .Y(new_n1482_));
  XOR2   g00480(.A(\A[692] ), .B(\A[691] ), .Y(new_n1483_));
  AOI22  g00481(.A0(new_n1483_), .A1(new_n1478_), .B0(new_n1482_), .B1(new_n1480_), .Y(new_n1484_));
  INV    g00482(.A(\A[696] ), .Y(new_n1485_));
  INV    g00483(.A(\A[695] ), .Y(new_n1486_));
  NAND2  g00484(.A(new_n1486_), .B(\A[694] ), .Y(new_n1487_));
  INV    g00485(.A(\A[694] ), .Y(new_n1488_));
  AOI21  g00486(.A0(\A[695] ), .A1(new_n1488_), .B0(new_n1485_), .Y(new_n1489_));
  XOR2   g00487(.A(\A[695] ), .B(\A[694] ), .Y(new_n1490_));
  AOI22  g00488(.A0(new_n1490_), .A1(new_n1485_), .B0(new_n1489_), .B1(new_n1487_), .Y(new_n1491_));
  NOR2   g00489(.A(new_n1486_), .B(new_n1488_), .Y(new_n1492_));
  AOI21  g00490(.A0(new_n1490_), .A1(\A[696] ), .B0(new_n1492_), .Y(new_n1493_));
  NOR2   g00491(.A(new_n1479_), .B(new_n1481_), .Y(new_n1494_));
  AOI21  g00492(.A0(new_n1483_), .A1(\A[693] ), .B0(new_n1494_), .Y(new_n1495_));
  XOR2   g00493(.A(new_n1491_), .B(new_n1484_), .Y(new_n1496_));
  XOR2   g00494(.A(new_n1496_), .B(new_n1477_), .Y(new_n1497_));
  INV    g00495(.A(\A[687] ), .Y(new_n1498_));
  INV    g00496(.A(\A[686] ), .Y(new_n1499_));
  NAND2  g00497(.A(new_n1499_), .B(\A[685] ), .Y(new_n1500_));
  INV    g00498(.A(\A[685] ), .Y(new_n1501_));
  AOI21  g00499(.A0(\A[686] ), .A1(new_n1501_), .B0(new_n1498_), .Y(new_n1502_));
  XOR2   g00500(.A(\A[686] ), .B(\A[685] ), .Y(new_n1503_));
  AOI22  g00501(.A0(new_n1503_), .A1(new_n1498_), .B0(new_n1502_), .B1(new_n1500_), .Y(new_n1504_));
  INV    g00502(.A(\A[690] ), .Y(new_n1505_));
  INV    g00503(.A(\A[689] ), .Y(new_n1506_));
  NAND2  g00504(.A(new_n1506_), .B(\A[688] ), .Y(new_n1507_));
  INV    g00505(.A(\A[688] ), .Y(new_n1508_));
  AOI21  g00506(.A0(\A[689] ), .A1(new_n1508_), .B0(new_n1505_), .Y(new_n1509_));
  XOR2   g00507(.A(\A[689] ), .B(\A[688] ), .Y(new_n1510_));
  AOI22  g00508(.A0(new_n1510_), .A1(new_n1505_), .B0(new_n1509_), .B1(new_n1507_), .Y(new_n1511_));
  NOR2   g00509(.A(new_n1506_), .B(new_n1508_), .Y(new_n1512_));
  AOI21  g00510(.A0(new_n1510_), .A1(\A[690] ), .B0(new_n1512_), .Y(new_n1513_));
  NOR2   g00511(.A(new_n1499_), .B(new_n1501_), .Y(new_n1514_));
  AOI21  g00512(.A0(new_n1503_), .A1(\A[687] ), .B0(new_n1514_), .Y(new_n1515_));
  XOR2   g00513(.A(new_n1511_), .B(new_n1504_), .Y(new_n1516_));
  INV    g00514(.A(\A[681] ), .Y(new_n1517_));
  INV    g00515(.A(\A[680] ), .Y(new_n1518_));
  NAND2  g00516(.A(new_n1518_), .B(\A[679] ), .Y(new_n1519_));
  INV    g00517(.A(\A[679] ), .Y(new_n1520_));
  AOI21  g00518(.A0(\A[680] ), .A1(new_n1520_), .B0(new_n1517_), .Y(new_n1521_));
  XOR2   g00519(.A(\A[680] ), .B(\A[679] ), .Y(new_n1522_));
  AOI22  g00520(.A0(new_n1522_), .A1(new_n1517_), .B0(new_n1521_), .B1(new_n1519_), .Y(new_n1523_));
  INV    g00521(.A(\A[684] ), .Y(new_n1524_));
  INV    g00522(.A(\A[683] ), .Y(new_n1525_));
  NAND2  g00523(.A(new_n1525_), .B(\A[682] ), .Y(new_n1526_));
  INV    g00524(.A(\A[682] ), .Y(new_n1527_));
  AOI21  g00525(.A0(\A[683] ), .A1(new_n1527_), .B0(new_n1524_), .Y(new_n1528_));
  XOR2   g00526(.A(\A[683] ), .B(\A[682] ), .Y(new_n1529_));
  AOI22  g00527(.A0(new_n1529_), .A1(new_n1524_), .B0(new_n1528_), .B1(new_n1526_), .Y(new_n1530_));
  NOR2   g00528(.A(new_n1525_), .B(new_n1527_), .Y(new_n1531_));
  AOI21  g00529(.A0(new_n1529_), .A1(\A[684] ), .B0(new_n1531_), .Y(new_n1532_));
  NOR2   g00530(.A(new_n1518_), .B(new_n1520_), .Y(new_n1533_));
  AOI21  g00531(.A0(new_n1522_), .A1(\A[681] ), .B0(new_n1533_), .Y(new_n1534_));
  XOR2   g00532(.A(new_n1530_), .B(new_n1523_), .Y(new_n1535_));
  XOR2   g00533(.A(new_n1535_), .B(new_n1516_), .Y(new_n1536_));
  INV    g00534(.A(new_n1536_), .Y(new_n1537_));
  XOR2   g00535(.A(new_n1537_), .B(new_n1497_), .Y(new_n1538_));
  INV    g00536(.A(new_n1538_), .Y(new_n1539_));
  INV    g00537(.A(\A[675] ), .Y(new_n1540_));
  INV    g00538(.A(\A[674] ), .Y(new_n1541_));
  NAND2  g00539(.A(new_n1541_), .B(\A[673] ), .Y(new_n1542_));
  INV    g00540(.A(\A[673] ), .Y(new_n1543_));
  AOI21  g00541(.A0(\A[674] ), .A1(new_n1543_), .B0(new_n1540_), .Y(new_n1544_));
  XOR2   g00542(.A(\A[674] ), .B(\A[673] ), .Y(new_n1545_));
  AOI22  g00543(.A0(new_n1545_), .A1(new_n1540_), .B0(new_n1544_), .B1(new_n1542_), .Y(new_n1546_));
  INV    g00544(.A(\A[678] ), .Y(new_n1547_));
  INV    g00545(.A(\A[677] ), .Y(new_n1548_));
  NAND2  g00546(.A(new_n1548_), .B(\A[676] ), .Y(new_n1549_));
  INV    g00547(.A(\A[676] ), .Y(new_n1550_));
  AOI21  g00548(.A0(\A[677] ), .A1(new_n1550_), .B0(new_n1547_), .Y(new_n1551_));
  XOR2   g00549(.A(\A[677] ), .B(\A[676] ), .Y(new_n1552_));
  AOI22  g00550(.A0(new_n1552_), .A1(new_n1547_), .B0(new_n1551_), .B1(new_n1549_), .Y(new_n1553_));
  NOR2   g00551(.A(new_n1548_), .B(new_n1550_), .Y(new_n1554_));
  AOI21  g00552(.A0(new_n1552_), .A1(\A[678] ), .B0(new_n1554_), .Y(new_n1555_));
  NOR2   g00553(.A(new_n1541_), .B(new_n1543_), .Y(new_n1556_));
  AOI21  g00554(.A0(new_n1545_), .A1(\A[675] ), .B0(new_n1556_), .Y(new_n1557_));
  XOR2   g00555(.A(new_n1553_), .B(new_n1546_), .Y(new_n1558_));
  INV    g00556(.A(\A[669] ), .Y(new_n1559_));
  INV    g00557(.A(\A[668] ), .Y(new_n1560_));
  NAND2  g00558(.A(new_n1560_), .B(\A[667] ), .Y(new_n1561_));
  INV    g00559(.A(\A[667] ), .Y(new_n1562_));
  AOI21  g00560(.A0(\A[668] ), .A1(new_n1562_), .B0(new_n1559_), .Y(new_n1563_));
  XOR2   g00561(.A(\A[668] ), .B(\A[667] ), .Y(new_n1564_));
  AOI22  g00562(.A0(new_n1564_), .A1(new_n1559_), .B0(new_n1563_), .B1(new_n1561_), .Y(new_n1565_));
  INV    g00563(.A(\A[672] ), .Y(new_n1566_));
  INV    g00564(.A(\A[671] ), .Y(new_n1567_));
  NAND2  g00565(.A(new_n1567_), .B(\A[670] ), .Y(new_n1568_));
  INV    g00566(.A(\A[670] ), .Y(new_n1569_));
  AOI21  g00567(.A0(\A[671] ), .A1(new_n1569_), .B0(new_n1566_), .Y(new_n1570_));
  XOR2   g00568(.A(\A[671] ), .B(\A[670] ), .Y(new_n1571_));
  AOI22  g00569(.A0(new_n1571_), .A1(new_n1566_), .B0(new_n1570_), .B1(new_n1568_), .Y(new_n1572_));
  NOR2   g00570(.A(new_n1567_), .B(new_n1569_), .Y(new_n1573_));
  AOI21  g00571(.A0(new_n1571_), .A1(\A[672] ), .B0(new_n1573_), .Y(new_n1574_));
  NOR2   g00572(.A(new_n1560_), .B(new_n1562_), .Y(new_n1575_));
  AOI21  g00573(.A0(new_n1564_), .A1(\A[669] ), .B0(new_n1575_), .Y(new_n1576_));
  XOR2   g00574(.A(new_n1572_), .B(new_n1565_), .Y(new_n1577_));
  XOR2   g00575(.A(new_n1577_), .B(new_n1558_), .Y(new_n1578_));
  INV    g00576(.A(\A[663] ), .Y(new_n1579_));
  INV    g00577(.A(\A[662] ), .Y(new_n1580_));
  NAND2  g00578(.A(new_n1580_), .B(\A[661] ), .Y(new_n1581_));
  INV    g00579(.A(\A[661] ), .Y(new_n1582_));
  AOI21  g00580(.A0(\A[662] ), .A1(new_n1582_), .B0(new_n1579_), .Y(new_n1583_));
  XOR2   g00581(.A(\A[662] ), .B(\A[661] ), .Y(new_n1584_));
  AOI22  g00582(.A0(new_n1584_), .A1(new_n1579_), .B0(new_n1583_), .B1(new_n1581_), .Y(new_n1585_));
  INV    g00583(.A(\A[666] ), .Y(new_n1586_));
  INV    g00584(.A(\A[665] ), .Y(new_n1587_));
  NAND2  g00585(.A(new_n1587_), .B(\A[664] ), .Y(new_n1588_));
  INV    g00586(.A(\A[664] ), .Y(new_n1589_));
  AOI21  g00587(.A0(\A[665] ), .A1(new_n1589_), .B0(new_n1586_), .Y(new_n1590_));
  XOR2   g00588(.A(\A[665] ), .B(\A[664] ), .Y(new_n1591_));
  AOI22  g00589(.A0(new_n1591_), .A1(new_n1586_), .B0(new_n1590_), .B1(new_n1588_), .Y(new_n1592_));
  NOR2   g00590(.A(new_n1587_), .B(new_n1589_), .Y(new_n1593_));
  AOI21  g00591(.A0(new_n1591_), .A1(\A[666] ), .B0(new_n1593_), .Y(new_n1594_));
  NOR2   g00592(.A(new_n1580_), .B(new_n1582_), .Y(new_n1595_));
  AOI21  g00593(.A0(new_n1584_), .A1(\A[663] ), .B0(new_n1595_), .Y(new_n1596_));
  XOR2   g00594(.A(new_n1592_), .B(new_n1585_), .Y(new_n1597_));
  INV    g00595(.A(\A[657] ), .Y(new_n1598_));
  INV    g00596(.A(\A[656] ), .Y(new_n1599_));
  NAND2  g00597(.A(new_n1599_), .B(\A[655] ), .Y(new_n1600_));
  INV    g00598(.A(\A[655] ), .Y(new_n1601_));
  AOI21  g00599(.A0(\A[656] ), .A1(new_n1601_), .B0(new_n1598_), .Y(new_n1602_));
  XOR2   g00600(.A(\A[656] ), .B(\A[655] ), .Y(new_n1603_));
  AOI22  g00601(.A0(new_n1603_), .A1(new_n1598_), .B0(new_n1602_), .B1(new_n1600_), .Y(new_n1604_));
  INV    g00602(.A(\A[660] ), .Y(new_n1605_));
  INV    g00603(.A(\A[659] ), .Y(new_n1606_));
  NAND2  g00604(.A(new_n1606_), .B(\A[658] ), .Y(new_n1607_));
  INV    g00605(.A(\A[658] ), .Y(new_n1608_));
  AOI21  g00606(.A0(\A[659] ), .A1(new_n1608_), .B0(new_n1605_), .Y(new_n1609_));
  XOR2   g00607(.A(\A[659] ), .B(\A[658] ), .Y(new_n1610_));
  AOI22  g00608(.A0(new_n1610_), .A1(new_n1605_), .B0(new_n1609_), .B1(new_n1607_), .Y(new_n1611_));
  NOR2   g00609(.A(new_n1606_), .B(new_n1608_), .Y(new_n1612_));
  AOI21  g00610(.A0(new_n1610_), .A1(\A[660] ), .B0(new_n1612_), .Y(new_n1613_));
  NOR2   g00611(.A(new_n1599_), .B(new_n1601_), .Y(new_n1614_));
  AOI21  g00612(.A0(new_n1603_), .A1(\A[657] ), .B0(new_n1614_), .Y(new_n1615_));
  XOR2   g00613(.A(new_n1611_), .B(new_n1604_), .Y(new_n1616_));
  XOR2   g00614(.A(new_n1616_), .B(new_n1597_), .Y(new_n1617_));
  INV    g00615(.A(new_n1617_), .Y(new_n1618_));
  XOR2   g00616(.A(new_n1618_), .B(new_n1578_), .Y(new_n1619_));
  XOR2   g00617(.A(new_n1619_), .B(new_n1539_), .Y(new_n1620_));
  NOR2   g00618(.A(new_n1620_), .B(new_n1458_), .Y(new_n1621_));
  NAND3  g00619(.A(new_n1621_), .B(new_n1456_), .C(new_n1447_), .Y(new_n1622_));
  NAND3  g00620(.A(new_n1439_), .B(new_n1445_), .C(new_n1443_), .Y(new_n1623_));
  OAI21  g00621(.A0(new_n1436_), .A1(new_n1425_), .B0(new_n1440_), .Y(new_n1624_));
  AOI21  g00622(.A0(new_n1624_), .A1(new_n1623_), .B0(new_n1453_), .Y(new_n1625_));
  NAND3  g00623(.A(new_n1440_), .B(new_n1445_), .C(new_n1443_), .Y(new_n1626_));
  OAI21  g00624(.A0(new_n1436_), .A1(new_n1425_), .B0(new_n1439_), .Y(new_n1627_));
  AOI21  g00625(.A0(new_n1627_), .A1(new_n1626_), .B0(new_n1219_), .Y(new_n1628_));
  INV    g00626(.A(new_n1621_), .Y(new_n1629_));
  OAI21  g00627(.A0(new_n1628_), .A1(new_n1625_), .B0(new_n1629_), .Y(new_n1630_));
  XOR2   g00628(.A(new_n1611_), .B(new_n1604_), .Y(new_n1631_));
  XOR2   g00629(.A(\A[659] ), .B(new_n1608_), .Y(new_n1632_));
  NAND2  g00630(.A(\A[659] ), .B(\A[658] ), .Y(new_n1633_));
  OAI21  g00631(.A0(new_n1632_), .A1(new_n1605_), .B0(new_n1633_), .Y(new_n1634_));
  XOR2   g00632(.A(new_n1615_), .B(new_n1634_), .Y(new_n1635_));
  NOR2   g00633(.A(\A[656] ), .B(new_n1601_), .Y(new_n1636_));
  OAI21  g00634(.A0(new_n1599_), .A1(\A[655] ), .B0(\A[657] ), .Y(new_n1637_));
  XOR2   g00635(.A(\A[656] ), .B(new_n1601_), .Y(new_n1638_));
  OAI22  g00636(.A0(new_n1638_), .A1(\A[657] ), .B0(new_n1637_), .B1(new_n1636_), .Y(new_n1639_));
  NOR2   g00637(.A(\A[659] ), .B(new_n1608_), .Y(new_n1640_));
  OAI21  g00638(.A0(new_n1606_), .A1(\A[658] ), .B0(\A[660] ), .Y(new_n1641_));
  OAI22  g00639(.A0(new_n1632_), .A1(\A[660] ), .B0(new_n1641_), .B1(new_n1640_), .Y(new_n1642_));
  NAND2  g00640(.A(new_n1642_), .B(new_n1639_), .Y(new_n1643_));
  NAND2  g00641(.A(\A[656] ), .B(\A[655] ), .Y(new_n1644_));
  OAI21  g00642(.A0(new_n1638_), .A1(new_n1598_), .B0(new_n1644_), .Y(new_n1645_));
  NAND2  g00643(.A(new_n1645_), .B(new_n1634_), .Y(new_n1646_));
  OAI21  g00644(.A0(new_n1643_), .A1(new_n1635_), .B0(new_n1646_), .Y(new_n1647_));
  NOR2   g00645(.A(new_n1611_), .B(new_n1604_), .Y(new_n1648_));
  XOR2   g00646(.A(new_n1648_), .B(new_n1635_), .Y(new_n1649_));
  AOI21  g00647(.A0(new_n1647_), .A1(new_n1631_), .B0(new_n1649_), .Y(new_n1650_));
  XOR2   g00648(.A(new_n1592_), .B(new_n1585_), .Y(new_n1651_));
  NOR2   g00649(.A(\A[662] ), .B(new_n1582_), .Y(new_n1652_));
  OAI21  g00650(.A0(new_n1580_), .A1(\A[661] ), .B0(\A[663] ), .Y(new_n1653_));
  NAND2  g00651(.A(new_n1584_), .B(new_n1579_), .Y(new_n1654_));
  OAI21  g00652(.A0(new_n1653_), .A1(new_n1652_), .B0(new_n1654_), .Y(new_n1655_));
  NOR2   g00653(.A(\A[665] ), .B(new_n1589_), .Y(new_n1656_));
  OAI21  g00654(.A0(new_n1587_), .A1(\A[664] ), .B0(\A[666] ), .Y(new_n1657_));
  NAND2  g00655(.A(new_n1591_), .B(new_n1586_), .Y(new_n1658_));
  OAI21  g00656(.A0(new_n1657_), .A1(new_n1656_), .B0(new_n1658_), .Y(new_n1659_));
  NAND2  g00657(.A(new_n1591_), .B(\A[666] ), .Y(new_n1660_));
  OAI21  g00658(.A0(new_n1587_), .A1(new_n1589_), .B0(new_n1660_), .Y(new_n1661_));
  NAND2  g00659(.A(new_n1584_), .B(\A[663] ), .Y(new_n1662_));
  OAI21  g00660(.A0(new_n1580_), .A1(new_n1582_), .B0(new_n1662_), .Y(new_n1663_));
  NAND4  g00661(.A(new_n1663_), .B(new_n1661_), .C(new_n1659_), .D(new_n1655_), .Y(new_n1664_));
  NAND4  g00662(.A(new_n1645_), .B(new_n1634_), .C(new_n1642_), .D(new_n1639_), .Y(new_n1665_));
  NAND4  g00663(.A(new_n1665_), .B(new_n1631_), .C(new_n1664_), .D(new_n1651_), .Y(new_n1666_));
  XOR2   g00664(.A(new_n1596_), .B(new_n1661_), .Y(new_n1667_));
  NAND2  g00665(.A(new_n1659_), .B(new_n1655_), .Y(new_n1668_));
  NAND2  g00666(.A(new_n1663_), .B(new_n1661_), .Y(new_n1669_));
  OAI21  g00667(.A0(new_n1668_), .A1(new_n1667_), .B0(new_n1669_), .Y(new_n1670_));
  NOR2   g00668(.A(new_n1592_), .B(new_n1585_), .Y(new_n1671_));
  XOR2   g00669(.A(new_n1671_), .B(new_n1667_), .Y(new_n1672_));
  AOI21  g00670(.A0(new_n1670_), .A1(new_n1651_), .B0(new_n1672_), .Y(new_n1673_));
  XOR2   g00671(.A(new_n1673_), .B(new_n1666_), .Y(new_n1674_));
  XOR2   g00672(.A(new_n1592_), .B(new_n1655_), .Y(new_n1675_));
  NOR4   g00673(.A(new_n1596_), .B(new_n1594_), .C(new_n1592_), .D(new_n1585_), .Y(new_n1676_));
  XOR2   g00674(.A(new_n1611_), .B(new_n1639_), .Y(new_n1677_));
  NOR4   g00675(.A(new_n1615_), .B(new_n1613_), .C(new_n1611_), .D(new_n1604_), .Y(new_n1678_));
  NOR4   g00676(.A(new_n1678_), .B(new_n1677_), .C(new_n1676_), .D(new_n1675_), .Y(new_n1679_));
  XOR2   g00677(.A(new_n1596_), .B(new_n1594_), .Y(new_n1680_));
  NOR2   g00678(.A(new_n1596_), .B(new_n1594_), .Y(new_n1681_));
  AOI21  g00679(.A0(new_n1671_), .A1(new_n1680_), .B0(new_n1681_), .Y(new_n1682_));
  NOR4   g00680(.A(new_n1677_), .B(new_n1676_), .C(new_n1672_), .D(new_n1675_), .Y(new_n1683_));
  OAI211 g00681(.A0(new_n1682_), .A1(new_n1675_), .B0(new_n1683_), .B1(new_n1665_), .Y(new_n1684_));
  OAI21  g00682(.A0(new_n1673_), .A1(new_n1679_), .B0(new_n1684_), .Y(new_n1685_));
  NAND2  g00683(.A(new_n1685_), .B(new_n1650_), .Y(new_n1686_));
  OAI21  g00684(.A0(new_n1674_), .A1(new_n1650_), .B0(new_n1686_), .Y(new_n1687_));
  XOR2   g00685(.A(new_n1572_), .B(new_n1565_), .Y(new_n1688_));
  XOR2   g00686(.A(\A[671] ), .B(new_n1569_), .Y(new_n1689_));
  NAND2  g00687(.A(\A[671] ), .B(\A[670] ), .Y(new_n1690_));
  OAI21  g00688(.A0(new_n1689_), .A1(new_n1566_), .B0(new_n1690_), .Y(new_n1691_));
  XOR2   g00689(.A(new_n1576_), .B(new_n1691_), .Y(new_n1692_));
  NOR2   g00690(.A(\A[668] ), .B(new_n1562_), .Y(new_n1693_));
  OAI21  g00691(.A0(new_n1560_), .A1(\A[667] ), .B0(\A[669] ), .Y(new_n1694_));
  XOR2   g00692(.A(\A[668] ), .B(new_n1562_), .Y(new_n1695_));
  OAI22  g00693(.A0(new_n1695_), .A1(\A[669] ), .B0(new_n1694_), .B1(new_n1693_), .Y(new_n1696_));
  NOR2   g00694(.A(\A[671] ), .B(new_n1569_), .Y(new_n1697_));
  OAI21  g00695(.A0(new_n1567_), .A1(\A[670] ), .B0(\A[672] ), .Y(new_n1698_));
  OAI22  g00696(.A0(new_n1689_), .A1(\A[672] ), .B0(new_n1698_), .B1(new_n1697_), .Y(new_n1699_));
  NAND2  g00697(.A(new_n1699_), .B(new_n1696_), .Y(new_n1700_));
  NAND2  g00698(.A(\A[668] ), .B(\A[667] ), .Y(new_n1701_));
  OAI21  g00699(.A0(new_n1695_), .A1(new_n1559_), .B0(new_n1701_), .Y(new_n1702_));
  NAND2  g00700(.A(new_n1702_), .B(new_n1691_), .Y(new_n1703_));
  OAI21  g00701(.A0(new_n1700_), .A1(new_n1692_), .B0(new_n1703_), .Y(new_n1704_));
  NOR2   g00702(.A(new_n1572_), .B(new_n1565_), .Y(new_n1705_));
  XOR2   g00703(.A(new_n1705_), .B(new_n1692_), .Y(new_n1706_));
  AOI21  g00704(.A0(new_n1704_), .A1(new_n1688_), .B0(new_n1706_), .Y(new_n1707_));
  XOR2   g00705(.A(new_n1553_), .B(new_n1546_), .Y(new_n1708_));
  NOR2   g00706(.A(\A[674] ), .B(new_n1543_), .Y(new_n1709_));
  OAI21  g00707(.A0(new_n1541_), .A1(\A[673] ), .B0(\A[675] ), .Y(new_n1710_));
  NAND2  g00708(.A(new_n1545_), .B(new_n1540_), .Y(new_n1711_));
  OAI21  g00709(.A0(new_n1710_), .A1(new_n1709_), .B0(new_n1711_), .Y(new_n1712_));
  NOR2   g00710(.A(\A[677] ), .B(new_n1550_), .Y(new_n1713_));
  OAI21  g00711(.A0(new_n1548_), .A1(\A[676] ), .B0(\A[678] ), .Y(new_n1714_));
  NAND2  g00712(.A(new_n1552_), .B(new_n1547_), .Y(new_n1715_));
  OAI21  g00713(.A0(new_n1714_), .A1(new_n1713_), .B0(new_n1715_), .Y(new_n1716_));
  NAND2  g00714(.A(new_n1552_), .B(\A[678] ), .Y(new_n1717_));
  OAI21  g00715(.A0(new_n1548_), .A1(new_n1550_), .B0(new_n1717_), .Y(new_n1718_));
  NAND2  g00716(.A(new_n1545_), .B(\A[675] ), .Y(new_n1719_));
  OAI21  g00717(.A0(new_n1541_), .A1(new_n1543_), .B0(new_n1719_), .Y(new_n1720_));
  NAND4  g00718(.A(new_n1720_), .B(new_n1718_), .C(new_n1716_), .D(new_n1712_), .Y(new_n1721_));
  NAND4  g00719(.A(new_n1702_), .B(new_n1691_), .C(new_n1699_), .D(new_n1696_), .Y(new_n1722_));
  NAND4  g00720(.A(new_n1722_), .B(new_n1688_), .C(new_n1721_), .D(new_n1708_), .Y(new_n1723_));
  XOR2   g00721(.A(new_n1557_), .B(new_n1718_), .Y(new_n1724_));
  NAND2  g00722(.A(new_n1716_), .B(new_n1712_), .Y(new_n1725_));
  NAND2  g00723(.A(new_n1720_), .B(new_n1718_), .Y(new_n1726_));
  OAI21  g00724(.A0(new_n1725_), .A1(new_n1724_), .B0(new_n1726_), .Y(new_n1727_));
  NOR2   g00725(.A(new_n1553_), .B(new_n1546_), .Y(new_n1728_));
  XOR2   g00726(.A(new_n1728_), .B(new_n1724_), .Y(new_n1729_));
  AOI21  g00727(.A0(new_n1727_), .A1(new_n1708_), .B0(new_n1729_), .Y(new_n1730_));
  XOR2   g00728(.A(new_n1730_), .B(new_n1723_), .Y(new_n1731_));
  NOR2   g00729(.A(new_n1731_), .B(new_n1707_), .Y(new_n1732_));
  XOR2   g00730(.A(new_n1572_), .B(new_n1696_), .Y(new_n1733_));
  XOR2   g00731(.A(new_n1576_), .B(new_n1574_), .Y(new_n1734_));
  NOR2   g00732(.A(new_n1576_), .B(new_n1574_), .Y(new_n1735_));
  AOI21  g00733(.A0(new_n1705_), .A1(new_n1734_), .B0(new_n1735_), .Y(new_n1736_));
  XOR2   g00734(.A(new_n1705_), .B(new_n1734_), .Y(new_n1737_));
  OAI21  g00735(.A0(new_n1736_), .A1(new_n1733_), .B0(new_n1737_), .Y(new_n1738_));
  XOR2   g00736(.A(new_n1553_), .B(new_n1712_), .Y(new_n1739_));
  XOR2   g00737(.A(new_n1557_), .B(new_n1555_), .Y(new_n1740_));
  NOR2   g00738(.A(new_n1557_), .B(new_n1555_), .Y(new_n1741_));
  AOI21  g00739(.A0(new_n1728_), .A1(new_n1740_), .B0(new_n1741_), .Y(new_n1742_));
  XOR2   g00740(.A(new_n1728_), .B(new_n1740_), .Y(new_n1743_));
  OAI21  g00741(.A0(new_n1742_), .A1(new_n1739_), .B0(new_n1743_), .Y(new_n1744_));
  NAND2  g00742(.A(new_n1744_), .B(new_n1723_), .Y(new_n1745_));
  NOR4   g00743(.A(new_n1557_), .B(new_n1555_), .C(new_n1553_), .D(new_n1546_), .Y(new_n1746_));
  NOR4   g00744(.A(new_n1733_), .B(new_n1746_), .C(new_n1729_), .D(new_n1739_), .Y(new_n1747_));
  OAI211 g00745(.A0(new_n1742_), .A1(new_n1739_), .B0(new_n1747_), .B1(new_n1722_), .Y(new_n1748_));
  AOI21  g00746(.A0(new_n1748_), .A1(new_n1745_), .B0(new_n1738_), .Y(new_n1749_));
  NAND2  g00747(.A(new_n1617_), .B(new_n1578_), .Y(new_n1750_));
  NOR3   g00748(.A(new_n1750_), .B(new_n1749_), .C(new_n1732_), .Y(new_n1751_));
  NOR4   g00749(.A(new_n1576_), .B(new_n1574_), .C(new_n1572_), .D(new_n1565_), .Y(new_n1752_));
  NOR4   g00750(.A(new_n1752_), .B(new_n1733_), .C(new_n1746_), .D(new_n1739_), .Y(new_n1753_));
  XOR2   g00751(.A(new_n1730_), .B(new_n1753_), .Y(new_n1754_));
  NAND2  g00752(.A(new_n1754_), .B(new_n1738_), .Y(new_n1755_));
  NAND4  g00753(.A(new_n1688_), .B(new_n1721_), .C(new_n1743_), .D(new_n1708_), .Y(new_n1756_));
  OAI21  g00754(.A0(new_n1742_), .A1(new_n1739_), .B0(new_n1722_), .Y(new_n1757_));
  OAI22  g00755(.A0(new_n1757_), .A1(new_n1756_), .B0(new_n1730_), .B1(new_n1753_), .Y(new_n1758_));
  NAND2  g00756(.A(new_n1758_), .B(new_n1707_), .Y(new_n1759_));
  INV    g00757(.A(new_n1750_), .Y(new_n1760_));
  AOI21  g00758(.A0(new_n1759_), .A1(new_n1755_), .B0(new_n1760_), .Y(new_n1761_));
  NOR2   g00759(.A(new_n1761_), .B(new_n1751_), .Y(new_n1762_));
  NOR2   g00760(.A(new_n1687_), .B(new_n1762_), .Y(new_n1763_));
  NOR2   g00761(.A(new_n1749_), .B(new_n1732_), .Y(new_n1764_));
  NAND3  g00762(.A(new_n1750_), .B(new_n1759_), .C(new_n1755_), .Y(new_n1765_));
  OAI21  g00763(.A0(new_n1764_), .A1(new_n1750_), .B0(new_n1765_), .Y(new_n1766_));
  AOI21  g00764(.A0(new_n1766_), .A1(new_n1687_), .B0(new_n1763_), .Y(new_n1767_));
  XOR2   g00765(.A(new_n1530_), .B(new_n1523_), .Y(new_n1768_));
  XOR2   g00766(.A(\A[683] ), .B(new_n1527_), .Y(new_n1769_));
  NAND2  g00767(.A(\A[683] ), .B(\A[682] ), .Y(new_n1770_));
  OAI21  g00768(.A0(new_n1769_), .A1(new_n1524_), .B0(new_n1770_), .Y(new_n1771_));
  XOR2   g00769(.A(new_n1534_), .B(new_n1771_), .Y(new_n1772_));
  NOR2   g00770(.A(\A[680] ), .B(new_n1520_), .Y(new_n1773_));
  OAI21  g00771(.A0(new_n1518_), .A1(\A[679] ), .B0(\A[681] ), .Y(new_n1774_));
  XOR2   g00772(.A(\A[680] ), .B(new_n1520_), .Y(new_n1775_));
  OAI22  g00773(.A0(new_n1775_), .A1(\A[681] ), .B0(new_n1774_), .B1(new_n1773_), .Y(new_n1776_));
  NOR2   g00774(.A(\A[683] ), .B(new_n1527_), .Y(new_n1777_));
  OAI21  g00775(.A0(new_n1525_), .A1(\A[682] ), .B0(\A[684] ), .Y(new_n1778_));
  OAI22  g00776(.A0(new_n1769_), .A1(\A[684] ), .B0(new_n1778_), .B1(new_n1777_), .Y(new_n1779_));
  NAND2  g00777(.A(new_n1779_), .B(new_n1776_), .Y(new_n1780_));
  NAND2  g00778(.A(\A[680] ), .B(\A[679] ), .Y(new_n1781_));
  OAI21  g00779(.A0(new_n1775_), .A1(new_n1517_), .B0(new_n1781_), .Y(new_n1782_));
  NAND2  g00780(.A(new_n1782_), .B(new_n1771_), .Y(new_n1783_));
  OAI21  g00781(.A0(new_n1780_), .A1(new_n1772_), .B0(new_n1783_), .Y(new_n1784_));
  NOR2   g00782(.A(new_n1530_), .B(new_n1523_), .Y(new_n1785_));
  XOR2   g00783(.A(new_n1785_), .B(new_n1772_), .Y(new_n1786_));
  AOI21  g00784(.A0(new_n1784_), .A1(new_n1768_), .B0(new_n1786_), .Y(new_n1787_));
  XOR2   g00785(.A(new_n1511_), .B(new_n1504_), .Y(new_n1788_));
  NOR2   g00786(.A(\A[686] ), .B(new_n1501_), .Y(new_n1789_));
  OAI21  g00787(.A0(new_n1499_), .A1(\A[685] ), .B0(\A[687] ), .Y(new_n1790_));
  NAND2  g00788(.A(new_n1503_), .B(new_n1498_), .Y(new_n1791_));
  OAI21  g00789(.A0(new_n1790_), .A1(new_n1789_), .B0(new_n1791_), .Y(new_n1792_));
  NOR2   g00790(.A(\A[689] ), .B(new_n1508_), .Y(new_n1793_));
  OAI21  g00791(.A0(new_n1506_), .A1(\A[688] ), .B0(\A[690] ), .Y(new_n1794_));
  NAND2  g00792(.A(new_n1510_), .B(new_n1505_), .Y(new_n1795_));
  OAI21  g00793(.A0(new_n1794_), .A1(new_n1793_), .B0(new_n1795_), .Y(new_n1796_));
  NAND2  g00794(.A(new_n1510_), .B(\A[690] ), .Y(new_n1797_));
  OAI21  g00795(.A0(new_n1506_), .A1(new_n1508_), .B0(new_n1797_), .Y(new_n1798_));
  NAND2  g00796(.A(new_n1503_), .B(\A[687] ), .Y(new_n1799_));
  OAI21  g00797(.A0(new_n1499_), .A1(new_n1501_), .B0(new_n1799_), .Y(new_n1800_));
  NAND4  g00798(.A(new_n1800_), .B(new_n1798_), .C(new_n1796_), .D(new_n1792_), .Y(new_n1801_));
  NAND4  g00799(.A(new_n1782_), .B(new_n1771_), .C(new_n1779_), .D(new_n1776_), .Y(new_n1802_));
  NAND4  g00800(.A(new_n1802_), .B(new_n1768_), .C(new_n1801_), .D(new_n1788_), .Y(new_n1803_));
  XOR2   g00801(.A(new_n1515_), .B(new_n1798_), .Y(new_n1804_));
  NAND2  g00802(.A(new_n1796_), .B(new_n1792_), .Y(new_n1805_));
  NAND2  g00803(.A(new_n1800_), .B(new_n1798_), .Y(new_n1806_));
  OAI21  g00804(.A0(new_n1805_), .A1(new_n1804_), .B0(new_n1806_), .Y(new_n1807_));
  NOR2   g00805(.A(new_n1511_), .B(new_n1504_), .Y(new_n1808_));
  XOR2   g00806(.A(new_n1808_), .B(new_n1804_), .Y(new_n1809_));
  AOI21  g00807(.A0(new_n1807_), .A1(new_n1788_), .B0(new_n1809_), .Y(new_n1810_));
  XOR2   g00808(.A(new_n1810_), .B(new_n1803_), .Y(new_n1811_));
  XOR2   g00809(.A(new_n1511_), .B(new_n1792_), .Y(new_n1812_));
  NOR4   g00810(.A(new_n1515_), .B(new_n1513_), .C(new_n1511_), .D(new_n1504_), .Y(new_n1813_));
  XOR2   g00811(.A(new_n1530_), .B(new_n1776_), .Y(new_n1814_));
  NOR4   g00812(.A(new_n1534_), .B(new_n1532_), .C(new_n1530_), .D(new_n1523_), .Y(new_n1815_));
  NOR4   g00813(.A(new_n1815_), .B(new_n1814_), .C(new_n1813_), .D(new_n1812_), .Y(new_n1816_));
  XOR2   g00814(.A(new_n1515_), .B(new_n1513_), .Y(new_n1817_));
  NOR2   g00815(.A(new_n1515_), .B(new_n1513_), .Y(new_n1818_));
  AOI21  g00816(.A0(new_n1808_), .A1(new_n1817_), .B0(new_n1818_), .Y(new_n1819_));
  NOR4   g00817(.A(new_n1814_), .B(new_n1813_), .C(new_n1809_), .D(new_n1812_), .Y(new_n1820_));
  OAI211 g00818(.A0(new_n1819_), .A1(new_n1812_), .B0(new_n1820_), .B1(new_n1802_), .Y(new_n1821_));
  OAI21  g00819(.A0(new_n1810_), .A1(new_n1816_), .B0(new_n1821_), .Y(new_n1822_));
  NAND2  g00820(.A(new_n1822_), .B(new_n1787_), .Y(new_n1823_));
  OAI21  g00821(.A0(new_n1811_), .A1(new_n1787_), .B0(new_n1823_), .Y(new_n1824_));
  NOR2   g00822(.A(\A[692] ), .B(new_n1481_), .Y(new_n1825_));
  OAI21  g00823(.A0(new_n1479_), .A1(\A[691] ), .B0(\A[693] ), .Y(new_n1826_));
  XOR2   g00824(.A(\A[692] ), .B(new_n1481_), .Y(new_n1827_));
  OAI22  g00825(.A0(new_n1827_), .A1(\A[693] ), .B0(new_n1826_), .B1(new_n1825_), .Y(new_n1828_));
  XOR2   g00826(.A(new_n1491_), .B(new_n1828_), .Y(new_n1829_));
  XOR2   g00827(.A(new_n1495_), .B(new_n1493_), .Y(new_n1830_));
  NOR2   g00828(.A(new_n1491_), .B(new_n1484_), .Y(new_n1831_));
  NOR2   g00829(.A(new_n1495_), .B(new_n1493_), .Y(new_n1832_));
  AOI21  g00830(.A0(new_n1831_), .A1(new_n1830_), .B0(new_n1832_), .Y(new_n1833_));
  XOR2   g00831(.A(new_n1831_), .B(new_n1830_), .Y(new_n1834_));
  OAI21  g00832(.A0(new_n1833_), .A1(new_n1829_), .B0(new_n1834_), .Y(new_n1835_));
  NOR2   g00833(.A(\A[698] ), .B(new_n1462_), .Y(new_n1836_));
  OAI21  g00834(.A0(new_n1460_), .A1(\A[697] ), .B0(\A[699] ), .Y(new_n1837_));
  NAND2  g00835(.A(new_n1464_), .B(new_n1459_), .Y(new_n1838_));
  OAI21  g00836(.A0(new_n1837_), .A1(new_n1836_), .B0(new_n1838_), .Y(new_n1839_));
  XOR2   g00837(.A(new_n1472_), .B(new_n1839_), .Y(new_n1840_));
  NOR4   g00838(.A(new_n1476_), .B(new_n1474_), .C(new_n1472_), .D(new_n1465_), .Y(new_n1841_));
  NOR4   g00839(.A(new_n1495_), .B(new_n1493_), .C(new_n1491_), .D(new_n1484_), .Y(new_n1842_));
  NOR4   g00840(.A(new_n1842_), .B(new_n1829_), .C(new_n1841_), .D(new_n1840_), .Y(new_n1843_));
  XOR2   g00841(.A(new_n1472_), .B(new_n1465_), .Y(new_n1844_));
  NAND2  g00842(.A(new_n1471_), .B(\A[702] ), .Y(new_n1845_));
  OAI21  g00843(.A0(new_n1467_), .A1(new_n1469_), .B0(new_n1845_), .Y(new_n1846_));
  XOR2   g00844(.A(new_n1476_), .B(new_n1846_), .Y(new_n1847_));
  NOR2   g00845(.A(\A[701] ), .B(new_n1469_), .Y(new_n1848_));
  OAI21  g00846(.A0(new_n1467_), .A1(\A[700] ), .B0(\A[702] ), .Y(new_n1849_));
  NAND2  g00847(.A(new_n1471_), .B(new_n1466_), .Y(new_n1850_));
  OAI21  g00848(.A0(new_n1849_), .A1(new_n1848_), .B0(new_n1850_), .Y(new_n1851_));
  NAND2  g00849(.A(new_n1851_), .B(new_n1839_), .Y(new_n1852_));
  NAND2  g00850(.A(new_n1464_), .B(\A[699] ), .Y(new_n1853_));
  OAI21  g00851(.A0(new_n1460_), .A1(new_n1462_), .B0(new_n1853_), .Y(new_n1854_));
  NAND2  g00852(.A(new_n1854_), .B(new_n1846_), .Y(new_n1855_));
  OAI21  g00853(.A0(new_n1852_), .A1(new_n1847_), .B0(new_n1855_), .Y(new_n1856_));
  NOR2   g00854(.A(new_n1472_), .B(new_n1465_), .Y(new_n1857_));
  XOR2   g00855(.A(new_n1857_), .B(new_n1847_), .Y(new_n1858_));
  AOI21  g00856(.A0(new_n1856_), .A1(new_n1844_), .B0(new_n1858_), .Y(new_n1859_));
  XOR2   g00857(.A(new_n1859_), .B(new_n1843_), .Y(new_n1860_));
  NAND2  g00858(.A(new_n1860_), .B(new_n1835_), .Y(new_n1861_));
  XOR2   g00859(.A(new_n1491_), .B(new_n1484_), .Y(new_n1862_));
  XOR2   g00860(.A(\A[695] ), .B(new_n1488_), .Y(new_n1863_));
  NAND2  g00861(.A(\A[695] ), .B(\A[694] ), .Y(new_n1864_));
  OAI21  g00862(.A0(new_n1863_), .A1(new_n1485_), .B0(new_n1864_), .Y(new_n1865_));
  XOR2   g00863(.A(new_n1495_), .B(new_n1865_), .Y(new_n1866_));
  NOR2   g00864(.A(\A[695] ), .B(new_n1488_), .Y(new_n1867_));
  OAI21  g00865(.A0(new_n1486_), .A1(\A[694] ), .B0(\A[696] ), .Y(new_n1868_));
  OAI22  g00866(.A0(new_n1863_), .A1(\A[696] ), .B0(new_n1868_), .B1(new_n1867_), .Y(new_n1869_));
  NAND2  g00867(.A(new_n1869_), .B(new_n1828_), .Y(new_n1870_));
  NAND2  g00868(.A(\A[692] ), .B(\A[691] ), .Y(new_n1871_));
  OAI21  g00869(.A0(new_n1827_), .A1(new_n1478_), .B0(new_n1871_), .Y(new_n1872_));
  NAND2  g00870(.A(new_n1872_), .B(new_n1865_), .Y(new_n1873_));
  OAI21  g00871(.A0(new_n1870_), .A1(new_n1866_), .B0(new_n1873_), .Y(new_n1874_));
  XOR2   g00872(.A(new_n1831_), .B(new_n1866_), .Y(new_n1875_));
  AOI21  g00873(.A0(new_n1874_), .A1(new_n1862_), .B0(new_n1875_), .Y(new_n1876_));
  XOR2   g00874(.A(new_n1476_), .B(new_n1474_), .Y(new_n1877_));
  XOR2   g00875(.A(new_n1857_), .B(new_n1877_), .Y(new_n1878_));
  NAND4  g00876(.A(new_n1854_), .B(new_n1846_), .C(new_n1851_), .D(new_n1839_), .Y(new_n1879_));
  NAND4  g00877(.A(new_n1862_), .B(new_n1879_), .C(new_n1878_), .D(new_n1844_), .Y(new_n1880_));
  NOR2   g00878(.A(new_n1476_), .B(new_n1474_), .Y(new_n1881_));
  AOI21  g00879(.A0(new_n1857_), .A1(new_n1877_), .B0(new_n1881_), .Y(new_n1882_));
  NAND4  g00880(.A(new_n1872_), .B(new_n1865_), .C(new_n1869_), .D(new_n1828_), .Y(new_n1883_));
  OAI21  g00881(.A0(new_n1882_), .A1(new_n1840_), .B0(new_n1883_), .Y(new_n1884_));
  OAI22  g00882(.A0(new_n1884_), .A1(new_n1880_), .B0(new_n1859_), .B1(new_n1843_), .Y(new_n1885_));
  NAND2  g00883(.A(new_n1885_), .B(new_n1876_), .Y(new_n1886_));
  NAND2  g00884(.A(new_n1536_), .B(new_n1497_), .Y(new_n1887_));
  INV    g00885(.A(new_n1887_), .Y(new_n1888_));
  NAND3  g00886(.A(new_n1888_), .B(new_n1886_), .C(new_n1861_), .Y(new_n1889_));
  NAND2  g00887(.A(new_n1886_), .B(new_n1861_), .Y(new_n1890_));
  NAND2  g00888(.A(new_n1890_), .B(new_n1887_), .Y(new_n1891_));
  AOI21  g00889(.A0(new_n1891_), .A1(new_n1889_), .B0(new_n1824_), .Y(new_n1892_));
  NOR2   g00890(.A(new_n1811_), .B(new_n1787_), .Y(new_n1893_));
  AOI21  g00891(.A0(new_n1822_), .A1(new_n1787_), .B0(new_n1893_), .Y(new_n1894_));
  NAND4  g00892(.A(new_n1883_), .B(new_n1862_), .C(new_n1879_), .D(new_n1844_), .Y(new_n1895_));
  XOR2   g00893(.A(new_n1859_), .B(new_n1895_), .Y(new_n1896_));
  NOR2   g00894(.A(new_n1896_), .B(new_n1876_), .Y(new_n1897_));
  AOI211 g00895(.A0(new_n1885_), .A1(new_n1876_), .B(new_n1888_), .C(new_n1897_), .Y(new_n1898_));
  AOI21  g00896(.A0(new_n1886_), .A1(new_n1861_), .B0(new_n1887_), .Y(new_n1899_));
  NOR2   g00897(.A(new_n1899_), .B(new_n1898_), .Y(new_n1900_));
  NOR2   g00898(.A(new_n1619_), .B(new_n1538_), .Y(new_n1901_));
  OAI21  g00899(.A0(new_n1900_), .A1(new_n1894_), .B0(new_n1901_), .Y(new_n1902_));
  NOR2   g00900(.A(new_n1902_), .B(new_n1892_), .Y(new_n1903_));
  AOI21  g00901(.A0(new_n1885_), .A1(new_n1876_), .B0(new_n1897_), .Y(new_n1904_));
  OAI21  g00902(.A0(new_n1904_), .A1(new_n1888_), .B0(new_n1889_), .Y(new_n1905_));
  NAND2  g00903(.A(new_n1905_), .B(new_n1894_), .Y(new_n1906_));
  NAND3  g00904(.A(new_n1887_), .B(new_n1886_), .C(new_n1861_), .Y(new_n1907_));
  OAI21  g00905(.A0(new_n1904_), .A1(new_n1887_), .B0(new_n1907_), .Y(new_n1908_));
  NAND2  g00906(.A(new_n1908_), .B(new_n1824_), .Y(new_n1909_));
  AOI21  g00907(.A0(new_n1909_), .A1(new_n1906_), .B0(new_n1901_), .Y(new_n1910_));
  OAI21  g00908(.A0(new_n1910_), .A1(new_n1903_), .B0(new_n1767_), .Y(new_n1911_));
  NOR2   g00909(.A(new_n1900_), .B(new_n1894_), .Y(new_n1912_));
  NOR3   g00910(.A(new_n1901_), .B(new_n1912_), .C(new_n1892_), .Y(new_n1913_));
  INV    g00911(.A(new_n1901_), .Y(new_n1914_));
  AOI21  g00912(.A0(new_n1909_), .A1(new_n1906_), .B0(new_n1914_), .Y(new_n1915_));
  NOR2   g00913(.A(new_n1915_), .B(new_n1913_), .Y(new_n1916_));
  OAI21  g00914(.A0(new_n1916_), .A1(new_n1767_), .B0(new_n1911_), .Y(new_n1917_));
  AOI21  g00915(.A0(new_n1630_), .A1(new_n1622_), .B0(new_n1917_), .Y(new_n1918_));
  OAI21  g00916(.A0(new_n1912_), .A1(new_n1892_), .B0(new_n1914_), .Y(new_n1919_));
  OAI21  g00917(.A0(new_n1902_), .A1(new_n1892_), .B0(new_n1919_), .Y(new_n1920_));
  AOI21  g00918(.A0(new_n1908_), .A1(new_n1824_), .B0(new_n1901_), .Y(new_n1921_));
  NAND2  g00919(.A(new_n1921_), .B(new_n1906_), .Y(new_n1922_));
  OAI21  g00920(.A0(new_n1912_), .A1(new_n1892_), .B0(new_n1901_), .Y(new_n1923_));
  AOI21  g00921(.A0(new_n1923_), .A1(new_n1922_), .B0(new_n1767_), .Y(new_n1924_));
  AOI21  g00922(.A0(new_n1767_), .A1(new_n1920_), .B0(new_n1924_), .Y(new_n1925_));
  NAND3  g00923(.A(new_n1629_), .B(new_n1456_), .C(new_n1447_), .Y(new_n1926_));
  OAI21  g00924(.A0(new_n1628_), .A1(new_n1625_), .B0(new_n1621_), .Y(new_n1927_));
  AOI21  g00925(.A0(new_n1927_), .A1(new_n1926_), .B0(new_n1925_), .Y(new_n1928_));
  NOR2   g00926(.A(new_n1928_), .B(new_n1918_), .Y(new_n1929_));
  INV    g00927(.A(\A[753] ), .Y(new_n1930_));
  INV    g00928(.A(\A[752] ), .Y(new_n1931_));
  NAND2  g00929(.A(new_n1931_), .B(\A[751] ), .Y(new_n1932_));
  INV    g00930(.A(\A[751] ), .Y(new_n1933_));
  AOI21  g00931(.A0(\A[752] ), .A1(new_n1933_), .B0(new_n1930_), .Y(new_n1934_));
  XOR2   g00932(.A(\A[752] ), .B(\A[751] ), .Y(new_n1935_));
  AOI22  g00933(.A0(new_n1935_), .A1(new_n1930_), .B0(new_n1934_), .B1(new_n1932_), .Y(new_n1936_));
  INV    g00934(.A(\A[756] ), .Y(new_n1937_));
  INV    g00935(.A(\A[755] ), .Y(new_n1938_));
  NAND2  g00936(.A(new_n1938_), .B(\A[754] ), .Y(new_n1939_));
  INV    g00937(.A(\A[754] ), .Y(new_n1940_));
  AOI21  g00938(.A0(\A[755] ), .A1(new_n1940_), .B0(new_n1937_), .Y(new_n1941_));
  XOR2   g00939(.A(\A[755] ), .B(\A[754] ), .Y(new_n1942_));
  AOI22  g00940(.A0(new_n1942_), .A1(new_n1937_), .B0(new_n1941_), .B1(new_n1939_), .Y(new_n1943_));
  XOR2   g00941(.A(new_n1943_), .B(new_n1936_), .Y(new_n1944_));
  XOR2   g00942(.A(\A[755] ), .B(new_n1940_), .Y(new_n1945_));
  NAND2  g00943(.A(\A[755] ), .B(\A[754] ), .Y(new_n1946_));
  OAI21  g00944(.A0(new_n1945_), .A1(new_n1937_), .B0(new_n1946_), .Y(new_n1947_));
  NOR2   g00945(.A(new_n1931_), .B(new_n1933_), .Y(new_n1948_));
  AOI21  g00946(.A0(new_n1935_), .A1(\A[753] ), .B0(new_n1948_), .Y(new_n1949_));
  XOR2   g00947(.A(new_n1949_), .B(new_n1947_), .Y(new_n1950_));
  NOR2   g00948(.A(\A[752] ), .B(new_n1933_), .Y(new_n1951_));
  OAI21  g00949(.A0(new_n1931_), .A1(\A[751] ), .B0(\A[753] ), .Y(new_n1952_));
  XOR2   g00950(.A(\A[752] ), .B(new_n1933_), .Y(new_n1953_));
  OAI22  g00951(.A0(new_n1953_), .A1(\A[753] ), .B0(new_n1952_), .B1(new_n1951_), .Y(new_n1954_));
  NOR2   g00952(.A(\A[755] ), .B(new_n1940_), .Y(new_n1955_));
  OAI21  g00953(.A0(new_n1938_), .A1(\A[754] ), .B0(\A[756] ), .Y(new_n1956_));
  OAI22  g00954(.A0(new_n1945_), .A1(\A[756] ), .B0(new_n1956_), .B1(new_n1955_), .Y(new_n1957_));
  NAND2  g00955(.A(new_n1957_), .B(new_n1954_), .Y(new_n1958_));
  NAND2  g00956(.A(\A[752] ), .B(\A[751] ), .Y(new_n1959_));
  OAI21  g00957(.A0(new_n1953_), .A1(new_n1930_), .B0(new_n1959_), .Y(new_n1960_));
  NAND2  g00958(.A(new_n1960_), .B(new_n1947_), .Y(new_n1961_));
  OAI21  g00959(.A0(new_n1958_), .A1(new_n1950_), .B0(new_n1961_), .Y(new_n1962_));
  NOR2   g00960(.A(new_n1943_), .B(new_n1936_), .Y(new_n1963_));
  XOR2   g00961(.A(new_n1963_), .B(new_n1950_), .Y(new_n1964_));
  AOI21  g00962(.A0(new_n1962_), .A1(new_n1944_), .B0(new_n1964_), .Y(new_n1965_));
  INV    g00963(.A(\A[759] ), .Y(new_n1966_));
  INV    g00964(.A(\A[758] ), .Y(new_n1967_));
  NAND2  g00965(.A(new_n1967_), .B(\A[757] ), .Y(new_n1968_));
  INV    g00966(.A(\A[757] ), .Y(new_n1969_));
  AOI21  g00967(.A0(\A[758] ), .A1(new_n1969_), .B0(new_n1966_), .Y(new_n1970_));
  XOR2   g00968(.A(\A[758] ), .B(\A[757] ), .Y(new_n1971_));
  AOI22  g00969(.A0(new_n1971_), .A1(new_n1966_), .B0(new_n1970_), .B1(new_n1968_), .Y(new_n1972_));
  INV    g00970(.A(\A[762] ), .Y(new_n1973_));
  INV    g00971(.A(\A[761] ), .Y(new_n1974_));
  NAND2  g00972(.A(new_n1974_), .B(\A[760] ), .Y(new_n1975_));
  INV    g00973(.A(\A[760] ), .Y(new_n1976_));
  AOI21  g00974(.A0(\A[761] ), .A1(new_n1976_), .B0(new_n1973_), .Y(new_n1977_));
  XOR2   g00975(.A(\A[761] ), .B(\A[760] ), .Y(new_n1978_));
  AOI22  g00976(.A0(new_n1978_), .A1(new_n1973_), .B0(new_n1977_), .B1(new_n1975_), .Y(new_n1979_));
  XOR2   g00977(.A(new_n1979_), .B(new_n1972_), .Y(new_n1980_));
  NOR2   g00978(.A(\A[758] ), .B(new_n1969_), .Y(new_n1981_));
  OAI21  g00979(.A0(new_n1967_), .A1(\A[757] ), .B0(\A[759] ), .Y(new_n1982_));
  NAND2  g00980(.A(new_n1971_), .B(new_n1966_), .Y(new_n1983_));
  OAI21  g00981(.A0(new_n1982_), .A1(new_n1981_), .B0(new_n1983_), .Y(new_n1984_));
  NOR2   g00982(.A(\A[761] ), .B(new_n1976_), .Y(new_n1985_));
  OAI21  g00983(.A0(new_n1974_), .A1(\A[760] ), .B0(\A[762] ), .Y(new_n1986_));
  NAND2  g00984(.A(new_n1978_), .B(new_n1973_), .Y(new_n1987_));
  OAI21  g00985(.A0(new_n1986_), .A1(new_n1985_), .B0(new_n1987_), .Y(new_n1988_));
  NAND2  g00986(.A(new_n1978_), .B(\A[762] ), .Y(new_n1989_));
  OAI21  g00987(.A0(new_n1974_), .A1(new_n1976_), .B0(new_n1989_), .Y(new_n1990_));
  NAND2  g00988(.A(new_n1971_), .B(\A[759] ), .Y(new_n1991_));
  OAI21  g00989(.A0(new_n1967_), .A1(new_n1969_), .B0(new_n1991_), .Y(new_n1992_));
  NAND4  g00990(.A(new_n1992_), .B(new_n1990_), .C(new_n1988_), .D(new_n1984_), .Y(new_n1993_));
  NAND4  g00991(.A(new_n1960_), .B(new_n1947_), .C(new_n1957_), .D(new_n1954_), .Y(new_n1994_));
  NAND4  g00992(.A(new_n1994_), .B(new_n1944_), .C(new_n1993_), .D(new_n1980_), .Y(new_n1995_));
  NOR2   g00993(.A(new_n1967_), .B(new_n1969_), .Y(new_n1996_));
  AOI21  g00994(.A0(new_n1971_), .A1(\A[759] ), .B0(new_n1996_), .Y(new_n1997_));
  XOR2   g00995(.A(new_n1997_), .B(new_n1990_), .Y(new_n1998_));
  NAND2  g00996(.A(new_n1988_), .B(new_n1984_), .Y(new_n1999_));
  NAND2  g00997(.A(new_n1992_), .B(new_n1990_), .Y(new_n2000_));
  OAI21  g00998(.A0(new_n1999_), .A1(new_n1998_), .B0(new_n2000_), .Y(new_n2001_));
  NOR2   g00999(.A(new_n1979_), .B(new_n1972_), .Y(new_n2002_));
  XOR2   g01000(.A(new_n2002_), .B(new_n1998_), .Y(new_n2003_));
  AOI21  g01001(.A0(new_n2001_), .A1(new_n1980_), .B0(new_n2003_), .Y(new_n2004_));
  XOR2   g01002(.A(new_n2004_), .B(new_n1995_), .Y(new_n2005_));
  XOR2   g01003(.A(new_n1979_), .B(new_n1984_), .Y(new_n2006_));
  NOR2   g01004(.A(new_n1974_), .B(new_n1976_), .Y(new_n2007_));
  AOI21  g01005(.A0(new_n1978_), .A1(\A[762] ), .B0(new_n2007_), .Y(new_n2008_));
  NOR4   g01006(.A(new_n1997_), .B(new_n2008_), .C(new_n1979_), .D(new_n1972_), .Y(new_n2009_));
  XOR2   g01007(.A(new_n1943_), .B(new_n1954_), .Y(new_n2010_));
  NOR2   g01008(.A(new_n1938_), .B(new_n1940_), .Y(new_n2011_));
  AOI21  g01009(.A0(new_n1942_), .A1(\A[756] ), .B0(new_n2011_), .Y(new_n2012_));
  NOR4   g01010(.A(new_n1949_), .B(new_n2012_), .C(new_n1943_), .D(new_n1936_), .Y(new_n2013_));
  NOR4   g01011(.A(new_n2013_), .B(new_n2010_), .C(new_n2009_), .D(new_n2006_), .Y(new_n2014_));
  XOR2   g01012(.A(new_n1997_), .B(new_n2008_), .Y(new_n2015_));
  NOR2   g01013(.A(new_n1997_), .B(new_n2008_), .Y(new_n2016_));
  AOI21  g01014(.A0(new_n2002_), .A1(new_n2015_), .B0(new_n2016_), .Y(new_n2017_));
  NOR4   g01015(.A(new_n2010_), .B(new_n2009_), .C(new_n2003_), .D(new_n2006_), .Y(new_n2018_));
  OAI211 g01016(.A0(new_n2017_), .A1(new_n2006_), .B0(new_n2018_), .B1(new_n1994_), .Y(new_n2019_));
  OAI21  g01017(.A0(new_n2004_), .A1(new_n2014_), .B0(new_n2019_), .Y(new_n2020_));
  NAND2  g01018(.A(new_n2020_), .B(new_n1965_), .Y(new_n2021_));
  OAI21  g01019(.A0(new_n2005_), .A1(new_n1965_), .B0(new_n2021_), .Y(new_n2022_));
  INV    g01020(.A(\A[765] ), .Y(new_n2023_));
  INV    g01021(.A(\A[764] ), .Y(new_n2024_));
  NAND2  g01022(.A(new_n2024_), .B(\A[763] ), .Y(new_n2025_));
  INV    g01023(.A(\A[763] ), .Y(new_n2026_));
  AOI21  g01024(.A0(\A[764] ), .A1(new_n2026_), .B0(new_n2023_), .Y(new_n2027_));
  XOR2   g01025(.A(\A[764] ), .B(\A[763] ), .Y(new_n2028_));
  AOI22  g01026(.A0(new_n2028_), .A1(new_n2023_), .B0(new_n2027_), .B1(new_n2025_), .Y(new_n2029_));
  INV    g01027(.A(\A[768] ), .Y(new_n2030_));
  INV    g01028(.A(\A[767] ), .Y(new_n2031_));
  NAND2  g01029(.A(new_n2031_), .B(\A[766] ), .Y(new_n2032_));
  INV    g01030(.A(\A[766] ), .Y(new_n2033_));
  AOI21  g01031(.A0(\A[767] ), .A1(new_n2033_), .B0(new_n2030_), .Y(new_n2034_));
  XOR2   g01032(.A(\A[767] ), .B(\A[766] ), .Y(new_n2035_));
  AOI22  g01033(.A0(new_n2035_), .A1(new_n2030_), .B0(new_n2034_), .B1(new_n2032_), .Y(new_n2036_));
  XOR2   g01034(.A(new_n2036_), .B(new_n2029_), .Y(new_n2037_));
  XOR2   g01035(.A(\A[767] ), .B(new_n2033_), .Y(new_n2038_));
  NAND2  g01036(.A(\A[767] ), .B(\A[766] ), .Y(new_n2039_));
  OAI21  g01037(.A0(new_n2038_), .A1(new_n2030_), .B0(new_n2039_), .Y(new_n2040_));
  NOR2   g01038(.A(new_n2024_), .B(new_n2026_), .Y(new_n2041_));
  AOI21  g01039(.A0(new_n2028_), .A1(\A[765] ), .B0(new_n2041_), .Y(new_n2042_));
  XOR2   g01040(.A(new_n2042_), .B(new_n2040_), .Y(new_n2043_));
  NOR2   g01041(.A(\A[764] ), .B(new_n2026_), .Y(new_n2044_));
  OAI21  g01042(.A0(new_n2024_), .A1(\A[763] ), .B0(\A[765] ), .Y(new_n2045_));
  XOR2   g01043(.A(\A[764] ), .B(new_n2026_), .Y(new_n2046_));
  OAI22  g01044(.A0(new_n2046_), .A1(\A[765] ), .B0(new_n2045_), .B1(new_n2044_), .Y(new_n2047_));
  NOR2   g01045(.A(\A[767] ), .B(new_n2033_), .Y(new_n2048_));
  OAI21  g01046(.A0(new_n2031_), .A1(\A[766] ), .B0(\A[768] ), .Y(new_n2049_));
  OAI22  g01047(.A0(new_n2038_), .A1(\A[768] ), .B0(new_n2049_), .B1(new_n2048_), .Y(new_n2050_));
  NAND2  g01048(.A(new_n2050_), .B(new_n2047_), .Y(new_n2051_));
  NAND2  g01049(.A(\A[764] ), .B(\A[763] ), .Y(new_n2052_));
  OAI21  g01050(.A0(new_n2046_), .A1(new_n2023_), .B0(new_n2052_), .Y(new_n2053_));
  NAND2  g01051(.A(new_n2053_), .B(new_n2040_), .Y(new_n2054_));
  OAI21  g01052(.A0(new_n2051_), .A1(new_n2043_), .B0(new_n2054_), .Y(new_n2055_));
  NOR2   g01053(.A(new_n2036_), .B(new_n2029_), .Y(new_n2056_));
  XOR2   g01054(.A(new_n2056_), .B(new_n2043_), .Y(new_n2057_));
  AOI21  g01055(.A0(new_n2055_), .A1(new_n2037_), .B0(new_n2057_), .Y(new_n2058_));
  INV    g01056(.A(\A[771] ), .Y(new_n2059_));
  INV    g01057(.A(\A[770] ), .Y(new_n2060_));
  NAND2  g01058(.A(new_n2060_), .B(\A[769] ), .Y(new_n2061_));
  INV    g01059(.A(\A[769] ), .Y(new_n2062_));
  AOI21  g01060(.A0(\A[770] ), .A1(new_n2062_), .B0(new_n2059_), .Y(new_n2063_));
  XOR2   g01061(.A(\A[770] ), .B(\A[769] ), .Y(new_n2064_));
  AOI22  g01062(.A0(new_n2064_), .A1(new_n2059_), .B0(new_n2063_), .B1(new_n2061_), .Y(new_n2065_));
  INV    g01063(.A(\A[774] ), .Y(new_n2066_));
  INV    g01064(.A(\A[773] ), .Y(new_n2067_));
  NAND2  g01065(.A(new_n2067_), .B(\A[772] ), .Y(new_n2068_));
  INV    g01066(.A(\A[772] ), .Y(new_n2069_));
  AOI21  g01067(.A0(\A[773] ), .A1(new_n2069_), .B0(new_n2066_), .Y(new_n2070_));
  XOR2   g01068(.A(\A[773] ), .B(\A[772] ), .Y(new_n2071_));
  AOI22  g01069(.A0(new_n2071_), .A1(new_n2066_), .B0(new_n2070_), .B1(new_n2068_), .Y(new_n2072_));
  XOR2   g01070(.A(new_n2072_), .B(new_n2065_), .Y(new_n2073_));
  NOR2   g01071(.A(\A[770] ), .B(new_n2062_), .Y(new_n2074_));
  OAI21  g01072(.A0(new_n2060_), .A1(\A[769] ), .B0(\A[771] ), .Y(new_n2075_));
  NAND2  g01073(.A(new_n2064_), .B(new_n2059_), .Y(new_n2076_));
  OAI21  g01074(.A0(new_n2075_), .A1(new_n2074_), .B0(new_n2076_), .Y(new_n2077_));
  NOR2   g01075(.A(\A[773] ), .B(new_n2069_), .Y(new_n2078_));
  OAI21  g01076(.A0(new_n2067_), .A1(\A[772] ), .B0(\A[774] ), .Y(new_n2079_));
  NAND2  g01077(.A(new_n2071_), .B(new_n2066_), .Y(new_n2080_));
  OAI21  g01078(.A0(new_n2079_), .A1(new_n2078_), .B0(new_n2080_), .Y(new_n2081_));
  NAND2  g01079(.A(new_n2071_), .B(\A[774] ), .Y(new_n2082_));
  OAI21  g01080(.A0(new_n2067_), .A1(new_n2069_), .B0(new_n2082_), .Y(new_n2083_));
  NAND2  g01081(.A(new_n2064_), .B(\A[771] ), .Y(new_n2084_));
  OAI21  g01082(.A0(new_n2060_), .A1(new_n2062_), .B0(new_n2084_), .Y(new_n2085_));
  NAND4  g01083(.A(new_n2085_), .B(new_n2083_), .C(new_n2081_), .D(new_n2077_), .Y(new_n2086_));
  NAND4  g01084(.A(new_n2053_), .B(new_n2040_), .C(new_n2050_), .D(new_n2047_), .Y(new_n2087_));
  NAND4  g01085(.A(new_n2087_), .B(new_n2037_), .C(new_n2086_), .D(new_n2073_), .Y(new_n2088_));
  NOR2   g01086(.A(new_n2060_), .B(new_n2062_), .Y(new_n2089_));
  AOI21  g01087(.A0(new_n2064_), .A1(\A[771] ), .B0(new_n2089_), .Y(new_n2090_));
  XOR2   g01088(.A(new_n2090_), .B(new_n2083_), .Y(new_n2091_));
  NAND2  g01089(.A(new_n2081_), .B(new_n2077_), .Y(new_n2092_));
  NAND2  g01090(.A(new_n2085_), .B(new_n2083_), .Y(new_n2093_));
  OAI21  g01091(.A0(new_n2092_), .A1(new_n2091_), .B0(new_n2093_), .Y(new_n2094_));
  NOR2   g01092(.A(new_n2072_), .B(new_n2065_), .Y(new_n2095_));
  XOR2   g01093(.A(new_n2095_), .B(new_n2091_), .Y(new_n2096_));
  AOI21  g01094(.A0(new_n2094_), .A1(new_n2073_), .B0(new_n2096_), .Y(new_n2097_));
  XOR2   g01095(.A(new_n2097_), .B(new_n2088_), .Y(new_n2098_));
  NOR2   g01096(.A(new_n2098_), .B(new_n2058_), .Y(new_n2099_));
  XOR2   g01097(.A(new_n2036_), .B(new_n2047_), .Y(new_n2100_));
  NOR2   g01098(.A(new_n2031_), .B(new_n2033_), .Y(new_n2101_));
  AOI21  g01099(.A0(new_n2035_), .A1(\A[768] ), .B0(new_n2101_), .Y(new_n2102_));
  XOR2   g01100(.A(new_n2042_), .B(new_n2102_), .Y(new_n2103_));
  NOR2   g01101(.A(new_n2042_), .B(new_n2102_), .Y(new_n2104_));
  AOI21  g01102(.A0(new_n2056_), .A1(new_n2103_), .B0(new_n2104_), .Y(new_n2105_));
  XOR2   g01103(.A(new_n2056_), .B(new_n2103_), .Y(new_n2106_));
  OAI21  g01104(.A0(new_n2105_), .A1(new_n2100_), .B0(new_n2106_), .Y(new_n2107_));
  XOR2   g01105(.A(new_n2072_), .B(new_n2077_), .Y(new_n2108_));
  NOR2   g01106(.A(new_n2067_), .B(new_n2069_), .Y(new_n2109_));
  AOI21  g01107(.A0(new_n2071_), .A1(\A[774] ), .B0(new_n2109_), .Y(new_n2110_));
  XOR2   g01108(.A(new_n2090_), .B(new_n2110_), .Y(new_n2111_));
  NOR2   g01109(.A(new_n2090_), .B(new_n2110_), .Y(new_n2112_));
  AOI21  g01110(.A0(new_n2095_), .A1(new_n2111_), .B0(new_n2112_), .Y(new_n2113_));
  XOR2   g01111(.A(new_n2095_), .B(new_n2111_), .Y(new_n2114_));
  OAI21  g01112(.A0(new_n2113_), .A1(new_n2108_), .B0(new_n2114_), .Y(new_n2115_));
  NAND2  g01113(.A(new_n2115_), .B(new_n2088_), .Y(new_n2116_));
  NOR4   g01114(.A(new_n2090_), .B(new_n2110_), .C(new_n2072_), .D(new_n2065_), .Y(new_n2117_));
  NOR4   g01115(.A(new_n2100_), .B(new_n2117_), .C(new_n2096_), .D(new_n2108_), .Y(new_n2118_));
  OAI211 g01116(.A0(new_n2113_), .A1(new_n2108_), .B0(new_n2118_), .B1(new_n2087_), .Y(new_n2119_));
  AOI21  g01117(.A0(new_n2119_), .A1(new_n2116_), .B0(new_n2107_), .Y(new_n2120_));
  XOR2   g01118(.A(new_n2072_), .B(new_n2065_), .Y(new_n2121_));
  XOR2   g01119(.A(new_n2036_), .B(new_n2029_), .Y(new_n2122_));
  XOR2   g01120(.A(new_n2122_), .B(new_n2121_), .Y(new_n2123_));
  XOR2   g01121(.A(new_n1979_), .B(new_n1972_), .Y(new_n2124_));
  XOR2   g01122(.A(new_n1943_), .B(new_n1936_), .Y(new_n2125_));
  XOR2   g01123(.A(new_n2125_), .B(new_n2124_), .Y(new_n2126_));
  NAND2  g01124(.A(new_n2126_), .B(new_n2123_), .Y(new_n2127_));
  NOR3   g01125(.A(new_n2127_), .B(new_n2120_), .C(new_n2099_), .Y(new_n2128_));
  NOR4   g01126(.A(new_n2042_), .B(new_n2102_), .C(new_n2036_), .D(new_n2029_), .Y(new_n2129_));
  NOR4   g01127(.A(new_n2129_), .B(new_n2100_), .C(new_n2117_), .D(new_n2108_), .Y(new_n2130_));
  XOR2   g01128(.A(new_n2097_), .B(new_n2130_), .Y(new_n2131_));
  NAND2  g01129(.A(new_n2131_), .B(new_n2107_), .Y(new_n2132_));
  NAND4  g01130(.A(new_n2037_), .B(new_n2086_), .C(new_n2114_), .D(new_n2073_), .Y(new_n2133_));
  OAI21  g01131(.A0(new_n2113_), .A1(new_n2108_), .B0(new_n2087_), .Y(new_n2134_));
  OAI22  g01132(.A0(new_n2134_), .A1(new_n2133_), .B0(new_n2097_), .B1(new_n2130_), .Y(new_n2135_));
  NAND2  g01133(.A(new_n2135_), .B(new_n2058_), .Y(new_n2136_));
  INV    g01134(.A(new_n2127_), .Y(new_n2137_));
  AOI21  g01135(.A0(new_n2136_), .A1(new_n2132_), .B0(new_n2137_), .Y(new_n2138_));
  NOR2   g01136(.A(new_n2138_), .B(new_n2128_), .Y(new_n2139_));
  NOR2   g01137(.A(new_n2022_), .B(new_n2139_), .Y(new_n2140_));
  NOR2   g01138(.A(new_n2120_), .B(new_n2099_), .Y(new_n2141_));
  NAND3  g01139(.A(new_n2127_), .B(new_n2136_), .C(new_n2132_), .Y(new_n2142_));
  OAI21  g01140(.A0(new_n2141_), .A1(new_n2127_), .B0(new_n2142_), .Y(new_n2143_));
  AOI21  g01141(.A0(new_n2143_), .A1(new_n2022_), .B0(new_n2140_), .Y(new_n2144_));
  INV    g01142(.A(\A[776] ), .Y(new_n2145_));
  NOR2   g01143(.A(new_n2145_), .B(\A[775] ), .Y(new_n2146_));
  INV    g01144(.A(\A[775] ), .Y(new_n2147_));
  OAI21  g01145(.A0(\A[776] ), .A1(new_n2147_), .B0(\A[777] ), .Y(new_n2148_));
  XOR2   g01146(.A(\A[776] ), .B(new_n2147_), .Y(new_n2149_));
  OAI22  g01147(.A0(new_n2149_), .A1(\A[777] ), .B0(new_n2148_), .B1(new_n2146_), .Y(new_n2150_));
  INV    g01148(.A(\A[779] ), .Y(new_n2151_));
  NOR2   g01149(.A(new_n2151_), .B(\A[778] ), .Y(new_n2152_));
  INV    g01150(.A(\A[778] ), .Y(new_n2153_));
  OAI21  g01151(.A0(\A[779] ), .A1(new_n2153_), .B0(\A[780] ), .Y(new_n2154_));
  XOR2   g01152(.A(\A[779] ), .B(new_n2153_), .Y(new_n2155_));
  OAI22  g01153(.A0(new_n2155_), .A1(\A[780] ), .B0(new_n2154_), .B1(new_n2152_), .Y(new_n2156_));
  NAND2  g01154(.A(new_n2156_), .B(new_n2150_), .Y(new_n2157_));
  NAND2  g01155(.A(\A[779] ), .B(\A[778] ), .Y(new_n2158_));
  XOR2   g01156(.A(\A[779] ), .B(\A[778] ), .Y(new_n2159_));
  NAND2  g01157(.A(new_n2159_), .B(\A[780] ), .Y(new_n2160_));
  NAND2  g01158(.A(new_n2160_), .B(new_n2158_), .Y(new_n2161_));
  XOR2   g01159(.A(\A[776] ), .B(\A[775] ), .Y(new_n2162_));
  NOR2   g01160(.A(new_n2145_), .B(new_n2147_), .Y(new_n2163_));
  AOI21  g01161(.A0(new_n2162_), .A1(\A[777] ), .B0(new_n2163_), .Y(new_n2164_));
  XOR2   g01162(.A(new_n2164_), .B(new_n2161_), .Y(new_n2165_));
  XOR2   g01163(.A(new_n2165_), .B(new_n2157_), .Y(new_n2166_));
  INV    g01164(.A(\A[780] ), .Y(new_n2167_));
  NAND2  g01165(.A(\A[779] ), .B(new_n2153_), .Y(new_n2168_));
  AOI21  g01166(.A0(new_n2151_), .A1(\A[778] ), .B0(new_n2167_), .Y(new_n2169_));
  AOI22  g01167(.A0(new_n2159_), .A1(new_n2167_), .B0(new_n2169_), .B1(new_n2168_), .Y(new_n2170_));
  XOR2   g01168(.A(new_n2170_), .B(new_n2150_), .Y(new_n2171_));
  INV    g01169(.A(\A[777] ), .Y(new_n2172_));
  NAND2  g01170(.A(\A[776] ), .B(\A[775] ), .Y(new_n2173_));
  OAI21  g01171(.A0(new_n2149_), .A1(new_n2172_), .B0(new_n2173_), .Y(new_n2174_));
  NOR2   g01172(.A(new_n2165_), .B(new_n2157_), .Y(new_n2175_));
  AOI21  g01173(.A0(new_n2174_), .A1(new_n2161_), .B0(new_n2175_), .Y(new_n2176_));
  OAI21  g01174(.A0(new_n2176_), .A1(new_n2171_), .B0(new_n2166_), .Y(new_n2177_));
  NAND2  g01175(.A(\A[785] ), .B(\A[784] ), .Y(new_n2178_));
  XOR2   g01176(.A(\A[785] ), .B(\A[784] ), .Y(new_n2179_));
  NAND2  g01177(.A(new_n2179_), .B(\A[786] ), .Y(new_n2180_));
  NAND2  g01178(.A(new_n2180_), .B(new_n2178_), .Y(new_n2181_));
  INV    g01179(.A(\A[781] ), .Y(new_n2182_));
  INV    g01180(.A(\A[782] ), .Y(new_n2183_));
  NOR2   g01181(.A(new_n2183_), .B(new_n2182_), .Y(new_n2184_));
  XOR2   g01182(.A(\A[782] ), .B(\A[781] ), .Y(new_n2185_));
  AOI21  g01183(.A0(new_n2185_), .A1(\A[783] ), .B0(new_n2184_), .Y(new_n2186_));
  XOR2   g01184(.A(new_n2186_), .B(new_n2181_), .Y(new_n2187_));
  NOR2   g01185(.A(new_n2183_), .B(\A[781] ), .Y(new_n2188_));
  OAI21  g01186(.A0(\A[782] ), .A1(new_n2182_), .B0(\A[783] ), .Y(new_n2189_));
  INV    g01187(.A(\A[783] ), .Y(new_n2190_));
  NAND2  g01188(.A(new_n2185_), .B(new_n2190_), .Y(new_n2191_));
  OAI21  g01189(.A0(new_n2189_), .A1(new_n2188_), .B0(new_n2191_), .Y(new_n2192_));
  INV    g01190(.A(\A[785] ), .Y(new_n2193_));
  NOR2   g01191(.A(new_n2193_), .B(\A[784] ), .Y(new_n2194_));
  INV    g01192(.A(\A[784] ), .Y(new_n2195_));
  OAI21  g01193(.A0(\A[785] ), .A1(new_n2195_), .B0(\A[786] ), .Y(new_n2196_));
  INV    g01194(.A(\A[786] ), .Y(new_n2197_));
  NAND2  g01195(.A(new_n2179_), .B(new_n2197_), .Y(new_n2198_));
  OAI21  g01196(.A0(new_n2196_), .A1(new_n2194_), .B0(new_n2198_), .Y(new_n2199_));
  NAND2  g01197(.A(new_n2199_), .B(new_n2192_), .Y(new_n2200_));
  NAND2  g01198(.A(new_n2185_), .B(\A[783] ), .Y(new_n2201_));
  OAI21  g01199(.A0(new_n2183_), .A1(new_n2182_), .B0(new_n2201_), .Y(new_n2202_));
  NAND2  g01200(.A(new_n2202_), .B(new_n2181_), .Y(new_n2203_));
  OAI21  g01201(.A0(new_n2200_), .A1(new_n2187_), .B0(new_n2203_), .Y(new_n2204_));
  XOR2   g01202(.A(new_n2202_), .B(new_n2181_), .Y(new_n2205_));
  NAND2  g01203(.A(\A[782] ), .B(new_n2182_), .Y(new_n2206_));
  AOI21  g01204(.A0(new_n2183_), .A1(\A[781] ), .B0(new_n2190_), .Y(new_n2207_));
  AOI22  g01205(.A0(new_n2207_), .A1(new_n2206_), .B0(new_n2185_), .B1(new_n2190_), .Y(new_n2208_));
  NAND2  g01206(.A(\A[785] ), .B(new_n2195_), .Y(new_n2209_));
  AOI21  g01207(.A0(new_n2193_), .A1(\A[784] ), .B0(new_n2197_), .Y(new_n2210_));
  AOI22  g01208(.A0(new_n2210_), .A1(new_n2209_), .B0(new_n2179_), .B1(new_n2197_), .Y(new_n2211_));
  NOR2   g01209(.A(new_n2211_), .B(new_n2208_), .Y(new_n2212_));
  XOR2   g01210(.A(new_n2212_), .B(new_n2205_), .Y(new_n2213_));
  AOI211 g01211(.A0(new_n2160_), .A1(new_n2158_), .B(new_n2164_), .C(new_n2157_), .Y(new_n2214_));
  NAND2  g01212(.A(\A[776] ), .B(new_n2147_), .Y(new_n2215_));
  AOI21  g01213(.A0(new_n2145_), .A1(\A[775] ), .B0(new_n2172_), .Y(new_n2216_));
  AOI22  g01214(.A0(new_n2162_), .A1(new_n2172_), .B0(new_n2216_), .B1(new_n2215_), .Y(new_n2217_));
  XOR2   g01215(.A(new_n2170_), .B(new_n2217_), .Y(new_n2218_));
  XOR2   g01216(.A(new_n2211_), .B(new_n2208_), .Y(new_n2219_));
  NAND2  g01217(.A(new_n2219_), .B(new_n2218_), .Y(new_n2220_));
  AOI211 g01218(.A0(new_n2213_), .A1(new_n2204_), .B(new_n2220_), .C(new_n2214_), .Y(new_n2221_));
  XOR2   g01219(.A(new_n2212_), .B(new_n2187_), .Y(new_n2222_));
  AOI21  g01220(.A0(new_n2219_), .A1(new_n2204_), .B0(new_n2222_), .Y(new_n2223_));
  XOR2   g01221(.A(new_n2223_), .B(new_n2221_), .Y(new_n2224_));
  NAND2  g01222(.A(new_n2224_), .B(new_n2177_), .Y(new_n2225_));
  NAND4  g01223(.A(new_n2199_), .B(new_n2192_), .C(new_n2202_), .D(new_n2181_), .Y(new_n2226_));
  NAND4  g01224(.A(new_n2174_), .B(new_n2161_), .C(new_n2156_), .D(new_n2150_), .Y(new_n2227_));
  NAND4  g01225(.A(new_n2219_), .B(new_n2227_), .C(new_n2226_), .D(new_n2218_), .Y(new_n2228_));
  AOI21  g01226(.A0(new_n2180_), .A1(new_n2178_), .B0(new_n2186_), .Y(new_n2229_));
  AOI21  g01227(.A0(new_n2212_), .A1(new_n2205_), .B0(new_n2229_), .Y(new_n2230_));
  XOR2   g01228(.A(new_n2211_), .B(new_n2192_), .Y(new_n2231_));
  OAI21  g01229(.A0(new_n2231_), .A1(new_n2230_), .B0(new_n2213_), .Y(new_n2232_));
  AOI221 g01230(.A0(new_n2211_), .A1(new_n2208_), .C0(new_n2186_), .B0(new_n2180_), .B1(new_n2178_), .Y(new_n2233_));
  NOR4   g01231(.A(new_n2233_), .B(new_n2220_), .C(new_n2214_), .D(new_n2222_), .Y(new_n2234_));
  AOI21  g01232(.A0(new_n2232_), .A1(new_n2228_), .B0(new_n2234_), .Y(new_n2235_));
  OAI21  g01233(.A0(new_n2235_), .A1(new_n2177_), .B0(new_n2225_), .Y(new_n2236_));
  INV    g01234(.A(\A[788] ), .Y(new_n2237_));
  NOR2   g01235(.A(new_n2237_), .B(\A[787] ), .Y(new_n2238_));
  INV    g01236(.A(\A[787] ), .Y(new_n2239_));
  OAI21  g01237(.A0(\A[788] ), .A1(new_n2239_), .B0(\A[789] ), .Y(new_n2240_));
  XOR2   g01238(.A(\A[788] ), .B(new_n2239_), .Y(new_n2241_));
  OAI22  g01239(.A0(new_n2241_), .A1(\A[789] ), .B0(new_n2240_), .B1(new_n2238_), .Y(new_n2242_));
  INV    g01240(.A(\A[791] ), .Y(new_n2243_));
  NOR2   g01241(.A(new_n2243_), .B(\A[790] ), .Y(new_n2244_));
  INV    g01242(.A(\A[790] ), .Y(new_n2245_));
  OAI21  g01243(.A0(\A[791] ), .A1(new_n2245_), .B0(\A[792] ), .Y(new_n2246_));
  XOR2   g01244(.A(\A[791] ), .B(new_n2245_), .Y(new_n2247_));
  OAI22  g01245(.A0(new_n2247_), .A1(\A[792] ), .B0(new_n2246_), .B1(new_n2244_), .Y(new_n2248_));
  NAND2  g01246(.A(new_n2248_), .B(new_n2242_), .Y(new_n2249_));
  NAND2  g01247(.A(\A[791] ), .B(\A[790] ), .Y(new_n2250_));
  XOR2   g01248(.A(\A[791] ), .B(\A[790] ), .Y(new_n2251_));
  NAND2  g01249(.A(new_n2251_), .B(\A[792] ), .Y(new_n2252_));
  NAND2  g01250(.A(new_n2252_), .B(new_n2250_), .Y(new_n2253_));
  XOR2   g01251(.A(\A[788] ), .B(\A[787] ), .Y(new_n2254_));
  NOR2   g01252(.A(new_n2237_), .B(new_n2239_), .Y(new_n2255_));
  AOI21  g01253(.A0(new_n2254_), .A1(\A[789] ), .B0(new_n2255_), .Y(new_n2256_));
  XOR2   g01254(.A(new_n2256_), .B(new_n2253_), .Y(new_n2257_));
  XOR2   g01255(.A(new_n2257_), .B(new_n2249_), .Y(new_n2258_));
  INV    g01256(.A(\A[789] ), .Y(new_n2259_));
  NAND2  g01257(.A(\A[788] ), .B(new_n2239_), .Y(new_n2260_));
  AOI21  g01258(.A0(new_n2237_), .A1(\A[787] ), .B0(new_n2259_), .Y(new_n2261_));
  AOI22  g01259(.A0(new_n2254_), .A1(new_n2259_), .B0(new_n2261_), .B1(new_n2260_), .Y(new_n2262_));
  INV    g01260(.A(\A[792] ), .Y(new_n2263_));
  NAND2  g01261(.A(\A[791] ), .B(new_n2245_), .Y(new_n2264_));
  AOI21  g01262(.A0(new_n2243_), .A1(\A[790] ), .B0(new_n2263_), .Y(new_n2265_));
  AOI22  g01263(.A0(new_n2251_), .A1(new_n2263_), .B0(new_n2265_), .B1(new_n2264_), .Y(new_n2266_));
  XOR2   g01264(.A(new_n2266_), .B(new_n2262_), .Y(new_n2267_));
  INV    g01265(.A(new_n2267_), .Y(new_n2268_));
  NAND2  g01266(.A(\A[788] ), .B(\A[787] ), .Y(new_n2269_));
  OAI21  g01267(.A0(new_n2241_), .A1(new_n2259_), .B0(new_n2269_), .Y(new_n2270_));
  NOR2   g01268(.A(new_n2257_), .B(new_n2249_), .Y(new_n2271_));
  AOI21  g01269(.A0(new_n2270_), .A1(new_n2253_), .B0(new_n2271_), .Y(new_n2272_));
  OAI21  g01270(.A0(new_n2272_), .A1(new_n2268_), .B0(new_n2258_), .Y(new_n2273_));
  INV    g01271(.A(\A[796] ), .Y(new_n2274_));
  INV    g01272(.A(\A[797] ), .Y(new_n2275_));
  NOR2   g01273(.A(new_n2275_), .B(new_n2274_), .Y(new_n2276_));
  XOR2   g01274(.A(\A[797] ), .B(\A[796] ), .Y(new_n2277_));
  AOI21  g01275(.A0(new_n2277_), .A1(\A[798] ), .B0(new_n2276_), .Y(new_n2278_));
  INV    g01276(.A(\A[793] ), .Y(new_n2279_));
  INV    g01277(.A(\A[794] ), .Y(new_n2280_));
  NOR2   g01278(.A(new_n2280_), .B(new_n2279_), .Y(new_n2281_));
  XOR2   g01279(.A(\A[794] ), .B(\A[793] ), .Y(new_n2282_));
  AOI21  g01280(.A0(new_n2282_), .A1(\A[795] ), .B0(new_n2281_), .Y(new_n2283_));
  INV    g01281(.A(\A[795] ), .Y(new_n2284_));
  NAND2  g01282(.A(\A[794] ), .B(new_n2279_), .Y(new_n2285_));
  AOI21  g01283(.A0(new_n2280_), .A1(\A[793] ), .B0(new_n2284_), .Y(new_n2286_));
  AOI22  g01284(.A0(new_n2286_), .A1(new_n2285_), .B0(new_n2282_), .B1(new_n2284_), .Y(new_n2287_));
  INV    g01285(.A(\A[798] ), .Y(new_n2288_));
  NAND2  g01286(.A(\A[797] ), .B(new_n2274_), .Y(new_n2289_));
  AOI21  g01287(.A0(new_n2275_), .A1(\A[796] ), .B0(new_n2288_), .Y(new_n2290_));
  AOI22  g01288(.A0(new_n2290_), .A1(new_n2289_), .B0(new_n2277_), .B1(new_n2288_), .Y(new_n2291_));
  NOR4   g01289(.A(new_n2291_), .B(new_n2287_), .C(new_n2283_), .D(new_n2278_), .Y(new_n2292_));
  AOI211 g01290(.A0(new_n2252_), .A1(new_n2250_), .B(new_n2256_), .C(new_n2249_), .Y(new_n2293_));
  XOR2   g01291(.A(new_n2291_), .B(new_n2287_), .Y(new_n2294_));
  NAND2  g01292(.A(new_n2294_), .B(new_n2267_), .Y(new_n2295_));
  NOR3   g01293(.A(new_n2295_), .B(new_n2293_), .C(new_n2292_), .Y(new_n2296_));
  NAND2  g01294(.A(new_n2277_), .B(\A[798] ), .Y(new_n2297_));
  OAI21  g01295(.A0(new_n2275_), .A1(new_n2274_), .B0(new_n2297_), .Y(new_n2298_));
  XOR2   g01296(.A(new_n2283_), .B(new_n2298_), .Y(new_n2299_));
  NOR2   g01297(.A(new_n2280_), .B(\A[793] ), .Y(new_n2300_));
  OAI21  g01298(.A0(\A[794] ), .A1(new_n2279_), .B0(\A[795] ), .Y(new_n2301_));
  NAND2  g01299(.A(new_n2282_), .B(new_n2284_), .Y(new_n2302_));
  OAI21  g01300(.A0(new_n2301_), .A1(new_n2300_), .B0(new_n2302_), .Y(new_n2303_));
  NOR2   g01301(.A(new_n2275_), .B(\A[796] ), .Y(new_n2304_));
  OAI21  g01302(.A0(\A[797] ), .A1(new_n2274_), .B0(\A[798] ), .Y(new_n2305_));
  NAND2  g01303(.A(new_n2277_), .B(new_n2288_), .Y(new_n2306_));
  OAI21  g01304(.A0(new_n2305_), .A1(new_n2304_), .B0(new_n2306_), .Y(new_n2307_));
  NAND2  g01305(.A(new_n2307_), .B(new_n2303_), .Y(new_n2308_));
  NAND2  g01306(.A(new_n2282_), .B(\A[795] ), .Y(new_n2309_));
  OAI21  g01307(.A0(new_n2280_), .A1(new_n2279_), .B0(new_n2309_), .Y(new_n2310_));
  NAND2  g01308(.A(new_n2310_), .B(new_n2298_), .Y(new_n2311_));
  OAI21  g01309(.A0(new_n2308_), .A1(new_n2299_), .B0(new_n2311_), .Y(new_n2312_));
  NOR2   g01310(.A(new_n2291_), .B(new_n2287_), .Y(new_n2313_));
  XOR2   g01311(.A(new_n2313_), .B(new_n2299_), .Y(new_n2314_));
  AOI21  g01312(.A0(new_n2294_), .A1(new_n2312_), .B0(new_n2314_), .Y(new_n2315_));
  XOR2   g01313(.A(new_n2315_), .B(new_n2296_), .Y(new_n2316_));
  NAND2  g01314(.A(new_n2316_), .B(new_n2273_), .Y(new_n2317_));
  NOR2   g01315(.A(new_n2266_), .B(new_n2262_), .Y(new_n2318_));
  XOR2   g01316(.A(new_n2257_), .B(new_n2318_), .Y(new_n2319_));
  NAND2  g01317(.A(new_n2270_), .B(new_n2253_), .Y(new_n2320_));
  OAI21  g01318(.A0(new_n2257_), .A1(new_n2249_), .B0(new_n2320_), .Y(new_n2321_));
  AOI21  g01319(.A0(new_n2321_), .A1(new_n2267_), .B0(new_n2319_), .Y(new_n2322_));
  NOR2   g01320(.A(new_n2315_), .B(new_n2296_), .Y(new_n2323_));
  AOI211 g01321(.A0(new_n2291_), .A1(new_n2287_), .B(new_n2283_), .C(new_n2278_), .Y(new_n2324_));
  NOR4   g01322(.A(new_n2324_), .B(new_n2295_), .C(new_n2293_), .D(new_n2314_), .Y(new_n2325_));
  OAI21  g01323(.A0(new_n2325_), .A1(new_n2323_), .B0(new_n2322_), .Y(new_n2326_));
  XOR2   g01324(.A(new_n2291_), .B(new_n2303_), .Y(new_n2327_));
  NOR2   g01325(.A(new_n2327_), .B(new_n2292_), .Y(new_n2328_));
  NAND4  g01326(.A(new_n2270_), .B(new_n2253_), .C(new_n2248_), .D(new_n2242_), .Y(new_n2329_));
  NAND2  g01327(.A(new_n2329_), .B(new_n2267_), .Y(new_n2330_));
  XOR2   g01328(.A(new_n2330_), .B(new_n2328_), .Y(new_n2331_));
  NAND2  g01329(.A(new_n2219_), .B(new_n2226_), .Y(new_n2332_));
  NAND3  g01330(.A(new_n2332_), .B(new_n2227_), .C(new_n2218_), .Y(new_n2333_));
  NAND2  g01331(.A(new_n2227_), .B(new_n2218_), .Y(new_n2334_));
  NAND3  g01332(.A(new_n2334_), .B(new_n2219_), .C(new_n2226_), .Y(new_n2335_));
  AOI21  g01333(.A0(new_n2335_), .A1(new_n2333_), .B0(new_n2331_), .Y(new_n2336_));
  NAND3  g01334(.A(new_n2336_), .B(new_n2326_), .C(new_n2317_), .Y(new_n2337_));
  NAND4  g01335(.A(new_n2307_), .B(new_n2303_), .C(new_n2310_), .D(new_n2298_), .Y(new_n2338_));
  NAND4  g01336(.A(new_n2294_), .B(new_n2329_), .C(new_n2338_), .D(new_n2267_), .Y(new_n2339_));
  XOR2   g01337(.A(new_n2315_), .B(new_n2339_), .Y(new_n2340_));
  NOR2   g01338(.A(new_n2340_), .B(new_n2322_), .Y(new_n2341_));
  XOR2   g01339(.A(new_n2310_), .B(new_n2298_), .Y(new_n2342_));
  NOR2   g01340(.A(new_n2283_), .B(new_n2278_), .Y(new_n2343_));
  AOI21  g01341(.A0(new_n2313_), .A1(new_n2342_), .B0(new_n2343_), .Y(new_n2344_));
  XOR2   g01342(.A(new_n2313_), .B(new_n2342_), .Y(new_n2345_));
  OAI21  g01343(.A0(new_n2327_), .A1(new_n2344_), .B0(new_n2345_), .Y(new_n2346_));
  AOI21  g01344(.A0(new_n2346_), .A1(new_n2339_), .B0(new_n2325_), .Y(new_n2347_));
  NOR2   g01345(.A(new_n2347_), .B(new_n2273_), .Y(new_n2348_));
  NAND2  g01346(.A(new_n2294_), .B(new_n2338_), .Y(new_n2349_));
  XOR2   g01347(.A(new_n2330_), .B(new_n2349_), .Y(new_n2350_));
  XOR2   g01348(.A(new_n2334_), .B(new_n2332_), .Y(new_n2351_));
  NAND2  g01349(.A(new_n2351_), .B(new_n2350_), .Y(new_n2352_));
  OAI21  g01350(.A0(new_n2348_), .A1(new_n2341_), .B0(new_n2352_), .Y(new_n2353_));
  AOI21  g01351(.A0(new_n2353_), .A1(new_n2337_), .B0(new_n2236_), .Y(new_n2354_));
  NOR2   g01352(.A(new_n2235_), .B(new_n2177_), .Y(new_n2355_));
  AOI21  g01353(.A0(new_n2224_), .A1(new_n2177_), .B0(new_n2355_), .Y(new_n2356_));
  NAND3  g01354(.A(new_n2352_), .B(new_n2326_), .C(new_n2317_), .Y(new_n2357_));
  OAI21  g01355(.A0(new_n2348_), .A1(new_n2341_), .B0(new_n2336_), .Y(new_n2358_));
  AOI21  g01356(.A0(new_n2358_), .A1(new_n2357_), .B0(new_n2356_), .Y(new_n2359_));
  XOR2   g01357(.A(new_n2351_), .B(new_n2331_), .Y(new_n2360_));
  INV    g01358(.A(new_n2126_), .Y(new_n2361_));
  XOR2   g01359(.A(new_n2361_), .B(new_n2123_), .Y(new_n2362_));
  NOR2   g01360(.A(new_n2362_), .B(new_n2360_), .Y(new_n2363_));
  INV    g01361(.A(new_n2363_), .Y(new_n2364_));
  NOR3   g01362(.A(new_n2364_), .B(new_n2359_), .C(new_n2354_), .Y(new_n2365_));
  NOR2   g01363(.A(new_n2359_), .B(new_n2354_), .Y(new_n2366_));
  NOR2   g01364(.A(new_n2366_), .B(new_n2363_), .Y(new_n2367_));
  OAI21  g01365(.A0(new_n2367_), .A1(new_n2365_), .B0(new_n2144_), .Y(new_n2368_));
  NOR3   g01366(.A(new_n2363_), .B(new_n2359_), .C(new_n2354_), .Y(new_n2369_));
  NOR2   g01367(.A(new_n2366_), .B(new_n2364_), .Y(new_n2370_));
  NOR2   g01368(.A(new_n2370_), .B(new_n2369_), .Y(new_n2371_));
  OAI21  g01369(.A0(new_n2371_), .A1(new_n2144_), .B0(new_n2368_), .Y(new_n2372_));
  INV    g01370(.A(\A[813] ), .Y(new_n2373_));
  INV    g01371(.A(\A[811] ), .Y(new_n2374_));
  NAND2  g01372(.A(\A[812] ), .B(new_n2374_), .Y(new_n2375_));
  INV    g01373(.A(\A[812] ), .Y(new_n2376_));
  AOI21  g01374(.A0(new_n2376_), .A1(\A[811] ), .B0(new_n2373_), .Y(new_n2377_));
  XOR2   g01375(.A(\A[812] ), .B(\A[811] ), .Y(new_n2378_));
  AOI22  g01376(.A0(new_n2378_), .A1(new_n2373_), .B0(new_n2377_), .B1(new_n2375_), .Y(new_n2379_));
  INV    g01377(.A(\A[816] ), .Y(new_n2380_));
  INV    g01378(.A(\A[814] ), .Y(new_n2381_));
  NAND2  g01379(.A(\A[815] ), .B(new_n2381_), .Y(new_n2382_));
  INV    g01380(.A(\A[815] ), .Y(new_n2383_));
  AOI21  g01381(.A0(new_n2383_), .A1(\A[814] ), .B0(new_n2380_), .Y(new_n2384_));
  XOR2   g01382(.A(\A[815] ), .B(\A[814] ), .Y(new_n2385_));
  AOI22  g01383(.A0(new_n2385_), .A1(new_n2380_), .B0(new_n2384_), .B1(new_n2382_), .Y(new_n2386_));
  NOR2   g01384(.A(new_n2386_), .B(new_n2379_), .Y(new_n2387_));
  NAND2  g01385(.A(\A[815] ), .B(\A[814] ), .Y(new_n2388_));
  NAND2  g01386(.A(new_n2385_), .B(\A[816] ), .Y(new_n2389_));
  NAND2  g01387(.A(new_n2389_), .B(new_n2388_), .Y(new_n2390_));
  NOR2   g01388(.A(new_n2376_), .B(new_n2374_), .Y(new_n2391_));
  AOI21  g01389(.A0(new_n2378_), .A1(\A[813] ), .B0(new_n2391_), .Y(new_n2392_));
  XOR2   g01390(.A(new_n2392_), .B(new_n2390_), .Y(new_n2393_));
  XOR2   g01391(.A(new_n2393_), .B(new_n2387_), .Y(new_n2394_));
  XOR2   g01392(.A(new_n2386_), .B(new_n2379_), .Y(new_n2395_));
  NOR2   g01393(.A(new_n2376_), .B(\A[811] ), .Y(new_n2396_));
  OAI21  g01394(.A0(\A[812] ), .A1(new_n2374_), .B0(\A[813] ), .Y(new_n2397_));
  XOR2   g01395(.A(\A[812] ), .B(new_n2374_), .Y(new_n2398_));
  OAI22  g01396(.A0(new_n2398_), .A1(\A[813] ), .B0(new_n2397_), .B1(new_n2396_), .Y(new_n2399_));
  NOR2   g01397(.A(new_n2383_), .B(\A[814] ), .Y(new_n2400_));
  OAI21  g01398(.A0(\A[815] ), .A1(new_n2381_), .B0(\A[816] ), .Y(new_n2401_));
  XOR2   g01399(.A(\A[815] ), .B(new_n2381_), .Y(new_n2402_));
  OAI22  g01400(.A0(new_n2402_), .A1(\A[816] ), .B0(new_n2401_), .B1(new_n2400_), .Y(new_n2403_));
  NAND2  g01401(.A(new_n2403_), .B(new_n2399_), .Y(new_n2404_));
  NAND2  g01402(.A(\A[812] ), .B(\A[811] ), .Y(new_n2405_));
  OAI21  g01403(.A0(new_n2398_), .A1(new_n2373_), .B0(new_n2405_), .Y(new_n2406_));
  NAND2  g01404(.A(new_n2406_), .B(new_n2390_), .Y(new_n2407_));
  OAI21  g01405(.A0(new_n2393_), .A1(new_n2404_), .B0(new_n2407_), .Y(new_n2408_));
  AOI21  g01406(.A0(new_n2408_), .A1(new_n2395_), .B0(new_n2394_), .Y(new_n2409_));
  INV    g01407(.A(\A[820] ), .Y(new_n2410_));
  INV    g01408(.A(\A[821] ), .Y(new_n2411_));
  XOR2   g01409(.A(\A[821] ), .B(\A[820] ), .Y(new_n2412_));
  NAND2  g01410(.A(new_n2412_), .B(\A[822] ), .Y(new_n2413_));
  OAI21  g01411(.A0(new_n2411_), .A1(new_n2410_), .B0(new_n2413_), .Y(new_n2414_));
  INV    g01412(.A(\A[817] ), .Y(new_n2415_));
  INV    g01413(.A(\A[818] ), .Y(new_n2416_));
  XOR2   g01414(.A(\A[818] ), .B(\A[817] ), .Y(new_n2417_));
  NAND2  g01415(.A(new_n2417_), .B(\A[819] ), .Y(new_n2418_));
  OAI21  g01416(.A0(new_n2416_), .A1(new_n2415_), .B0(new_n2418_), .Y(new_n2419_));
  NOR2   g01417(.A(new_n2416_), .B(\A[817] ), .Y(new_n2420_));
  OAI21  g01418(.A0(\A[818] ), .A1(new_n2415_), .B0(\A[819] ), .Y(new_n2421_));
  INV    g01419(.A(\A[819] ), .Y(new_n2422_));
  NAND2  g01420(.A(new_n2417_), .B(new_n2422_), .Y(new_n2423_));
  OAI21  g01421(.A0(new_n2421_), .A1(new_n2420_), .B0(new_n2423_), .Y(new_n2424_));
  NOR2   g01422(.A(new_n2411_), .B(\A[820] ), .Y(new_n2425_));
  OAI21  g01423(.A0(\A[821] ), .A1(new_n2410_), .B0(\A[822] ), .Y(new_n2426_));
  INV    g01424(.A(\A[822] ), .Y(new_n2427_));
  NAND2  g01425(.A(new_n2412_), .B(new_n2427_), .Y(new_n2428_));
  OAI21  g01426(.A0(new_n2426_), .A1(new_n2425_), .B0(new_n2428_), .Y(new_n2429_));
  NAND4  g01427(.A(new_n2429_), .B(new_n2424_), .C(new_n2419_), .D(new_n2414_), .Y(new_n2430_));
  NAND4  g01428(.A(new_n2406_), .B(new_n2390_), .C(new_n2403_), .D(new_n2399_), .Y(new_n2431_));
  NAND2  g01429(.A(\A[818] ), .B(new_n2415_), .Y(new_n2432_));
  AOI21  g01430(.A0(new_n2416_), .A1(\A[817] ), .B0(new_n2422_), .Y(new_n2433_));
  AOI22  g01431(.A0(new_n2433_), .A1(new_n2432_), .B0(new_n2417_), .B1(new_n2422_), .Y(new_n2434_));
  NAND2  g01432(.A(\A[821] ), .B(new_n2410_), .Y(new_n2435_));
  AOI21  g01433(.A0(new_n2411_), .A1(\A[820] ), .B0(new_n2427_), .Y(new_n2436_));
  AOI22  g01434(.A0(new_n2436_), .A1(new_n2435_), .B0(new_n2412_), .B1(new_n2427_), .Y(new_n2437_));
  XOR2   g01435(.A(new_n2437_), .B(new_n2434_), .Y(new_n2438_));
  NAND4  g01436(.A(new_n2438_), .B(new_n2431_), .C(new_n2430_), .D(new_n2395_), .Y(new_n2439_));
  NOR2   g01437(.A(new_n2416_), .B(new_n2415_), .Y(new_n2440_));
  AOI21  g01438(.A0(new_n2417_), .A1(\A[819] ), .B0(new_n2440_), .Y(new_n2441_));
  XOR2   g01439(.A(new_n2441_), .B(new_n2414_), .Y(new_n2442_));
  NAND2  g01440(.A(new_n2429_), .B(new_n2424_), .Y(new_n2443_));
  NAND2  g01441(.A(new_n2419_), .B(new_n2414_), .Y(new_n2444_));
  OAI21  g01442(.A0(new_n2443_), .A1(new_n2442_), .B0(new_n2444_), .Y(new_n2445_));
  NOR2   g01443(.A(new_n2437_), .B(new_n2434_), .Y(new_n2446_));
  XOR2   g01444(.A(new_n2446_), .B(new_n2442_), .Y(new_n2447_));
  AOI21  g01445(.A0(new_n2438_), .A1(new_n2445_), .B0(new_n2447_), .Y(new_n2448_));
  XOR2   g01446(.A(new_n2448_), .B(new_n2439_), .Y(new_n2449_));
  NOR2   g01447(.A(new_n2449_), .B(new_n2409_), .Y(new_n2450_));
  XOR2   g01448(.A(new_n2393_), .B(new_n2404_), .Y(new_n2451_));
  INV    g01449(.A(new_n2395_), .Y(new_n2452_));
  NOR2   g01450(.A(new_n2393_), .B(new_n2404_), .Y(new_n2453_));
  AOI21  g01451(.A0(new_n2406_), .A1(new_n2390_), .B0(new_n2453_), .Y(new_n2454_));
  OAI21  g01452(.A0(new_n2454_), .A1(new_n2452_), .B0(new_n2451_), .Y(new_n2455_));
  XOR2   g01453(.A(new_n2419_), .B(new_n2414_), .Y(new_n2456_));
  NOR2   g01454(.A(new_n2411_), .B(new_n2410_), .Y(new_n2457_));
  AOI21  g01455(.A0(new_n2412_), .A1(\A[822] ), .B0(new_n2457_), .Y(new_n2458_));
  NOR2   g01456(.A(new_n2441_), .B(new_n2458_), .Y(new_n2459_));
  AOI21  g01457(.A0(new_n2446_), .A1(new_n2456_), .B0(new_n2459_), .Y(new_n2460_));
  XOR2   g01458(.A(new_n2446_), .B(new_n2456_), .Y(new_n2461_));
  XOR2   g01459(.A(new_n2437_), .B(new_n2424_), .Y(new_n2462_));
  OAI21  g01460(.A0(new_n2462_), .A1(new_n2460_), .B0(new_n2461_), .Y(new_n2463_));
  AOI211 g01461(.A0(new_n2389_), .A1(new_n2388_), .B(new_n2392_), .C(new_n2404_), .Y(new_n2464_));
  NAND2  g01462(.A(new_n2438_), .B(new_n2395_), .Y(new_n2465_));
  AOI211 g01463(.A0(new_n2437_), .A1(new_n2434_), .B(new_n2441_), .C(new_n2458_), .Y(new_n2466_));
  NOR4   g01464(.A(new_n2466_), .B(new_n2465_), .C(new_n2464_), .D(new_n2447_), .Y(new_n2467_));
  AOI21  g01465(.A0(new_n2463_), .A1(new_n2439_), .B0(new_n2467_), .Y(new_n2468_));
  NOR2   g01466(.A(new_n2468_), .B(new_n2455_), .Y(new_n2469_));
  NAND2  g01467(.A(new_n2438_), .B(new_n2430_), .Y(new_n2470_));
  NAND2  g01468(.A(new_n2431_), .B(new_n2395_), .Y(new_n2471_));
  XOR2   g01469(.A(new_n2471_), .B(new_n2470_), .Y(new_n2472_));
  INV    g01470(.A(\A[807] ), .Y(new_n2473_));
  INV    g01471(.A(\A[806] ), .Y(new_n2474_));
  NAND2  g01472(.A(new_n2474_), .B(\A[805] ), .Y(new_n2475_));
  INV    g01473(.A(\A[805] ), .Y(new_n2476_));
  AOI21  g01474(.A0(\A[806] ), .A1(new_n2476_), .B0(new_n2473_), .Y(new_n2477_));
  XOR2   g01475(.A(\A[806] ), .B(\A[805] ), .Y(new_n2478_));
  AOI22  g01476(.A0(new_n2478_), .A1(new_n2473_), .B0(new_n2477_), .B1(new_n2475_), .Y(new_n2479_));
  INV    g01477(.A(\A[810] ), .Y(new_n2480_));
  INV    g01478(.A(\A[809] ), .Y(new_n2481_));
  NAND2  g01479(.A(new_n2481_), .B(\A[808] ), .Y(new_n2482_));
  INV    g01480(.A(\A[808] ), .Y(new_n2483_));
  AOI21  g01481(.A0(\A[809] ), .A1(new_n2483_), .B0(new_n2480_), .Y(new_n2484_));
  XOR2   g01482(.A(\A[809] ), .B(\A[808] ), .Y(new_n2485_));
  AOI22  g01483(.A0(new_n2485_), .A1(new_n2480_), .B0(new_n2484_), .B1(new_n2482_), .Y(new_n2486_));
  NOR2   g01484(.A(new_n2481_), .B(new_n2483_), .Y(new_n2487_));
  AOI21  g01485(.A0(new_n2485_), .A1(\A[810] ), .B0(new_n2487_), .Y(new_n2488_));
  NOR2   g01486(.A(new_n2474_), .B(new_n2476_), .Y(new_n2489_));
  AOI21  g01487(.A0(new_n2478_), .A1(\A[807] ), .B0(new_n2489_), .Y(new_n2490_));
  XOR2   g01488(.A(new_n2486_), .B(new_n2479_), .Y(new_n2491_));
  INV    g01489(.A(\A[801] ), .Y(new_n2492_));
  INV    g01490(.A(\A[800] ), .Y(new_n2493_));
  NAND2  g01491(.A(new_n2493_), .B(\A[799] ), .Y(new_n2494_));
  INV    g01492(.A(\A[799] ), .Y(new_n2495_));
  AOI21  g01493(.A0(\A[800] ), .A1(new_n2495_), .B0(new_n2492_), .Y(new_n2496_));
  XOR2   g01494(.A(\A[800] ), .B(\A[799] ), .Y(new_n2497_));
  AOI22  g01495(.A0(new_n2497_), .A1(new_n2492_), .B0(new_n2496_), .B1(new_n2494_), .Y(new_n2498_));
  INV    g01496(.A(\A[804] ), .Y(new_n2499_));
  INV    g01497(.A(\A[803] ), .Y(new_n2500_));
  NAND2  g01498(.A(new_n2500_), .B(\A[802] ), .Y(new_n2501_));
  INV    g01499(.A(\A[802] ), .Y(new_n2502_));
  AOI21  g01500(.A0(\A[803] ), .A1(new_n2502_), .B0(new_n2499_), .Y(new_n2503_));
  XOR2   g01501(.A(\A[803] ), .B(\A[802] ), .Y(new_n2504_));
  AOI22  g01502(.A0(new_n2504_), .A1(new_n2499_), .B0(new_n2503_), .B1(new_n2501_), .Y(new_n2505_));
  NOR2   g01503(.A(new_n2500_), .B(new_n2502_), .Y(new_n2506_));
  AOI21  g01504(.A0(new_n2504_), .A1(\A[804] ), .B0(new_n2506_), .Y(new_n2507_));
  NOR2   g01505(.A(new_n2493_), .B(new_n2495_), .Y(new_n2508_));
  AOI21  g01506(.A0(new_n2497_), .A1(\A[801] ), .B0(new_n2508_), .Y(new_n2509_));
  XOR2   g01507(.A(new_n2505_), .B(new_n2498_), .Y(new_n2510_));
  XOR2   g01508(.A(new_n2510_), .B(new_n2491_), .Y(new_n2511_));
  NAND2  g01509(.A(new_n2511_), .B(new_n2472_), .Y(new_n2512_));
  NOR3   g01510(.A(new_n2512_), .B(new_n2469_), .C(new_n2450_), .Y(new_n2513_));
  NOR4   g01511(.A(new_n2437_), .B(new_n2434_), .C(new_n2441_), .D(new_n2458_), .Y(new_n2514_));
  NOR3   g01512(.A(new_n2465_), .B(new_n2464_), .C(new_n2514_), .Y(new_n2515_));
  XOR2   g01513(.A(new_n2448_), .B(new_n2515_), .Y(new_n2516_));
  NAND2  g01514(.A(new_n2516_), .B(new_n2455_), .Y(new_n2517_));
  NOR2   g01515(.A(new_n2448_), .B(new_n2515_), .Y(new_n2518_));
  OAI21  g01516(.A0(new_n2467_), .A1(new_n2518_), .B0(new_n2409_), .Y(new_n2519_));
  NOR2   g01517(.A(new_n2462_), .B(new_n2514_), .Y(new_n2520_));
  XOR2   g01518(.A(new_n2471_), .B(new_n2520_), .Y(new_n2521_));
  INV    g01519(.A(new_n2511_), .Y(new_n2522_));
  NOR2   g01520(.A(new_n2522_), .B(new_n2521_), .Y(new_n2523_));
  AOI21  g01521(.A0(new_n2519_), .A1(new_n2517_), .B0(new_n2523_), .Y(new_n2524_));
  NOR2   g01522(.A(new_n2524_), .B(new_n2513_), .Y(new_n2525_));
  XOR2   g01523(.A(new_n2505_), .B(new_n2498_), .Y(new_n2526_));
  XOR2   g01524(.A(new_n2509_), .B(new_n2507_), .Y(new_n2527_));
  NOR2   g01525(.A(new_n2505_), .B(new_n2498_), .Y(new_n2528_));
  NAND2  g01526(.A(new_n2528_), .B(new_n2527_), .Y(new_n2529_));
  OAI21  g01527(.A0(new_n2509_), .A1(new_n2507_), .B0(new_n2529_), .Y(new_n2530_));
  INV    g01528(.A(new_n2504_), .Y(new_n2531_));
  NAND2  g01529(.A(\A[803] ), .B(\A[802] ), .Y(new_n2532_));
  OAI21  g01530(.A0(new_n2531_), .A1(new_n2499_), .B0(new_n2532_), .Y(new_n2533_));
  XOR2   g01531(.A(new_n2509_), .B(new_n2533_), .Y(new_n2534_));
  XOR2   g01532(.A(new_n2528_), .B(new_n2534_), .Y(new_n2535_));
  AOI21  g01533(.A0(new_n2530_), .A1(new_n2526_), .B0(new_n2535_), .Y(new_n2536_));
  XOR2   g01534(.A(new_n2486_), .B(new_n2479_), .Y(new_n2537_));
  NOR2   g01535(.A(\A[806] ), .B(new_n2476_), .Y(new_n2538_));
  OAI21  g01536(.A0(new_n2474_), .A1(\A[805] ), .B0(\A[807] ), .Y(new_n2539_));
  NAND2  g01537(.A(new_n2478_), .B(new_n2473_), .Y(new_n2540_));
  OAI21  g01538(.A0(new_n2539_), .A1(new_n2538_), .B0(new_n2540_), .Y(new_n2541_));
  NOR2   g01539(.A(\A[809] ), .B(new_n2483_), .Y(new_n2542_));
  OAI21  g01540(.A0(new_n2481_), .A1(\A[808] ), .B0(\A[810] ), .Y(new_n2543_));
  NAND2  g01541(.A(new_n2485_), .B(new_n2480_), .Y(new_n2544_));
  OAI21  g01542(.A0(new_n2543_), .A1(new_n2542_), .B0(new_n2544_), .Y(new_n2545_));
  NAND2  g01543(.A(new_n2485_), .B(\A[810] ), .Y(new_n2546_));
  OAI21  g01544(.A0(new_n2481_), .A1(new_n2483_), .B0(new_n2546_), .Y(new_n2547_));
  NAND2  g01545(.A(new_n2478_), .B(\A[807] ), .Y(new_n2548_));
  OAI21  g01546(.A0(new_n2474_), .A1(new_n2476_), .B0(new_n2548_), .Y(new_n2549_));
  NAND4  g01547(.A(new_n2549_), .B(new_n2547_), .C(new_n2545_), .D(new_n2541_), .Y(new_n2550_));
  INV    g01548(.A(new_n2497_), .Y(new_n2551_));
  NOR2   g01549(.A(new_n2551_), .B(new_n2492_), .Y(new_n2552_));
  OAI211 g01550(.A0(new_n2552_), .A1(new_n2508_), .B0(new_n2528_), .B1(new_n2533_), .Y(new_n2553_));
  NAND4  g01551(.A(new_n2553_), .B(new_n2526_), .C(new_n2550_), .D(new_n2537_), .Y(new_n2554_));
  XOR2   g01552(.A(new_n2490_), .B(new_n2547_), .Y(new_n2555_));
  NAND2  g01553(.A(new_n2545_), .B(new_n2541_), .Y(new_n2556_));
  NAND2  g01554(.A(new_n2549_), .B(new_n2547_), .Y(new_n2557_));
  OAI21  g01555(.A0(new_n2556_), .A1(new_n2555_), .B0(new_n2557_), .Y(new_n2558_));
  NOR2   g01556(.A(new_n2486_), .B(new_n2479_), .Y(new_n2559_));
  XOR2   g01557(.A(new_n2559_), .B(new_n2555_), .Y(new_n2560_));
  AOI21  g01558(.A0(new_n2558_), .A1(new_n2537_), .B0(new_n2560_), .Y(new_n2561_));
  XOR2   g01559(.A(new_n2561_), .B(new_n2554_), .Y(new_n2562_));
  XOR2   g01560(.A(new_n2486_), .B(new_n2541_), .Y(new_n2563_));
  XOR2   g01561(.A(new_n2490_), .B(new_n2488_), .Y(new_n2564_));
  NOR2   g01562(.A(new_n2490_), .B(new_n2488_), .Y(new_n2565_));
  AOI21  g01563(.A0(new_n2559_), .A1(new_n2564_), .B0(new_n2565_), .Y(new_n2566_));
  XOR2   g01564(.A(new_n2559_), .B(new_n2564_), .Y(new_n2567_));
  OAI21  g01565(.A0(new_n2566_), .A1(new_n2563_), .B0(new_n2567_), .Y(new_n2568_));
  NAND2  g01566(.A(new_n2568_), .B(new_n2554_), .Y(new_n2569_));
  NAND2  g01567(.A(new_n2496_), .B(new_n2494_), .Y(new_n2570_));
  OAI21  g01568(.A0(new_n2551_), .A1(\A[801] ), .B0(new_n2570_), .Y(new_n2571_));
  XOR2   g01569(.A(new_n2505_), .B(new_n2571_), .Y(new_n2572_));
  NOR4   g01570(.A(new_n2572_), .B(new_n2560_), .C(new_n2558_), .D(new_n2563_), .Y(new_n2573_));
  OAI211 g01571(.A0(new_n2566_), .A1(new_n2563_), .B0(new_n2573_), .B1(new_n2553_), .Y(new_n2574_));
  NAND2  g01572(.A(new_n2574_), .B(new_n2569_), .Y(new_n2575_));
  NAND2  g01573(.A(new_n2575_), .B(new_n2536_), .Y(new_n2576_));
  OAI21  g01574(.A0(new_n2562_), .A1(new_n2536_), .B0(new_n2576_), .Y(new_n2577_));
  NOR2   g01575(.A(new_n2577_), .B(new_n2525_), .Y(new_n2578_));
  NOR2   g01576(.A(new_n2562_), .B(new_n2536_), .Y(new_n2579_));
  NOR2   g01577(.A(new_n2509_), .B(new_n2507_), .Y(new_n2580_));
  AOI21  g01578(.A0(new_n2528_), .A1(new_n2527_), .B0(new_n2580_), .Y(new_n2581_));
  XOR2   g01579(.A(new_n2528_), .B(new_n2527_), .Y(new_n2582_));
  OAI21  g01580(.A0(new_n2581_), .A1(new_n2572_), .B0(new_n2582_), .Y(new_n2583_));
  AOI21  g01581(.A0(new_n2574_), .A1(new_n2569_), .B0(new_n2583_), .Y(new_n2584_));
  NOR2   g01582(.A(new_n2584_), .B(new_n2579_), .Y(new_n2585_));
  NAND3  g01583(.A(new_n2512_), .B(new_n2519_), .C(new_n2517_), .Y(new_n2586_));
  OAI21  g01584(.A0(new_n2469_), .A1(new_n2450_), .B0(new_n2523_), .Y(new_n2587_));
  AOI21  g01585(.A0(new_n2587_), .A1(new_n2586_), .B0(new_n2585_), .Y(new_n2588_));
  NOR2   g01586(.A(new_n2588_), .B(new_n2578_), .Y(new_n2589_));
  INV    g01587(.A(\A[825] ), .Y(new_n2590_));
  INV    g01588(.A(\A[823] ), .Y(new_n2591_));
  NAND2  g01589(.A(\A[824] ), .B(new_n2591_), .Y(new_n2592_));
  INV    g01590(.A(\A[824] ), .Y(new_n2593_));
  AOI21  g01591(.A0(new_n2593_), .A1(\A[823] ), .B0(new_n2590_), .Y(new_n2594_));
  XOR2   g01592(.A(\A[824] ), .B(\A[823] ), .Y(new_n2595_));
  AOI22  g01593(.A0(new_n2595_), .A1(new_n2590_), .B0(new_n2594_), .B1(new_n2592_), .Y(new_n2596_));
  INV    g01594(.A(\A[828] ), .Y(new_n2597_));
  INV    g01595(.A(\A[826] ), .Y(new_n2598_));
  NAND2  g01596(.A(\A[827] ), .B(new_n2598_), .Y(new_n2599_));
  INV    g01597(.A(\A[827] ), .Y(new_n2600_));
  AOI21  g01598(.A0(new_n2600_), .A1(\A[826] ), .B0(new_n2597_), .Y(new_n2601_));
  XOR2   g01599(.A(\A[827] ), .B(\A[826] ), .Y(new_n2602_));
  AOI22  g01600(.A0(new_n2602_), .A1(new_n2597_), .B0(new_n2601_), .B1(new_n2599_), .Y(new_n2603_));
  NOR2   g01601(.A(new_n2603_), .B(new_n2596_), .Y(new_n2604_));
  NAND2  g01602(.A(\A[827] ), .B(\A[826] ), .Y(new_n2605_));
  NAND2  g01603(.A(new_n2602_), .B(\A[828] ), .Y(new_n2606_));
  NAND2  g01604(.A(new_n2606_), .B(new_n2605_), .Y(new_n2607_));
  NOR2   g01605(.A(new_n2593_), .B(new_n2591_), .Y(new_n2608_));
  AOI21  g01606(.A0(new_n2595_), .A1(\A[825] ), .B0(new_n2608_), .Y(new_n2609_));
  XOR2   g01607(.A(new_n2609_), .B(new_n2607_), .Y(new_n2610_));
  XOR2   g01608(.A(new_n2610_), .B(new_n2604_), .Y(new_n2611_));
  XOR2   g01609(.A(new_n2603_), .B(new_n2596_), .Y(new_n2612_));
  NOR2   g01610(.A(new_n2593_), .B(\A[823] ), .Y(new_n2613_));
  OAI21  g01611(.A0(\A[824] ), .A1(new_n2591_), .B0(\A[825] ), .Y(new_n2614_));
  XOR2   g01612(.A(\A[824] ), .B(new_n2591_), .Y(new_n2615_));
  OAI22  g01613(.A0(new_n2615_), .A1(\A[825] ), .B0(new_n2614_), .B1(new_n2613_), .Y(new_n2616_));
  NOR2   g01614(.A(new_n2600_), .B(\A[826] ), .Y(new_n2617_));
  OAI21  g01615(.A0(\A[827] ), .A1(new_n2598_), .B0(\A[828] ), .Y(new_n2618_));
  XOR2   g01616(.A(\A[827] ), .B(new_n2598_), .Y(new_n2619_));
  OAI22  g01617(.A0(new_n2619_), .A1(\A[828] ), .B0(new_n2618_), .B1(new_n2617_), .Y(new_n2620_));
  NAND2  g01618(.A(new_n2620_), .B(new_n2616_), .Y(new_n2621_));
  NAND2  g01619(.A(\A[824] ), .B(\A[823] ), .Y(new_n2622_));
  OAI21  g01620(.A0(new_n2615_), .A1(new_n2590_), .B0(new_n2622_), .Y(new_n2623_));
  NAND2  g01621(.A(new_n2623_), .B(new_n2607_), .Y(new_n2624_));
  OAI21  g01622(.A0(new_n2610_), .A1(new_n2621_), .B0(new_n2624_), .Y(new_n2625_));
  AOI21  g01623(.A0(new_n2625_), .A1(new_n2612_), .B0(new_n2611_), .Y(new_n2626_));
  NAND2  g01624(.A(\A[833] ), .B(\A[832] ), .Y(new_n2627_));
  XOR2   g01625(.A(\A[833] ), .B(\A[832] ), .Y(new_n2628_));
  NAND2  g01626(.A(new_n2628_), .B(\A[834] ), .Y(new_n2629_));
  NAND2  g01627(.A(new_n2629_), .B(new_n2627_), .Y(new_n2630_));
  INV    g01628(.A(\A[829] ), .Y(new_n2631_));
  INV    g01629(.A(\A[830] ), .Y(new_n2632_));
  XOR2   g01630(.A(\A[830] ), .B(\A[829] ), .Y(new_n2633_));
  NAND2  g01631(.A(new_n2633_), .B(\A[831] ), .Y(new_n2634_));
  OAI21  g01632(.A0(new_n2632_), .A1(new_n2631_), .B0(new_n2634_), .Y(new_n2635_));
  NOR2   g01633(.A(new_n2632_), .B(\A[829] ), .Y(new_n2636_));
  OAI21  g01634(.A0(\A[830] ), .A1(new_n2631_), .B0(\A[831] ), .Y(new_n2637_));
  INV    g01635(.A(\A[831] ), .Y(new_n2638_));
  NAND2  g01636(.A(new_n2633_), .B(new_n2638_), .Y(new_n2639_));
  OAI21  g01637(.A0(new_n2637_), .A1(new_n2636_), .B0(new_n2639_), .Y(new_n2640_));
  INV    g01638(.A(\A[833] ), .Y(new_n2641_));
  NOR2   g01639(.A(new_n2641_), .B(\A[832] ), .Y(new_n2642_));
  INV    g01640(.A(\A[832] ), .Y(new_n2643_));
  OAI21  g01641(.A0(\A[833] ), .A1(new_n2643_), .B0(\A[834] ), .Y(new_n2644_));
  INV    g01642(.A(\A[834] ), .Y(new_n2645_));
  NAND2  g01643(.A(new_n2628_), .B(new_n2645_), .Y(new_n2646_));
  OAI21  g01644(.A0(new_n2644_), .A1(new_n2642_), .B0(new_n2646_), .Y(new_n2647_));
  NAND4  g01645(.A(new_n2647_), .B(new_n2640_), .C(new_n2635_), .D(new_n2630_), .Y(new_n2648_));
  NAND4  g01646(.A(new_n2623_), .B(new_n2607_), .C(new_n2620_), .D(new_n2616_), .Y(new_n2649_));
  NAND2  g01647(.A(\A[830] ), .B(new_n2631_), .Y(new_n2650_));
  AOI21  g01648(.A0(new_n2632_), .A1(\A[829] ), .B0(new_n2638_), .Y(new_n2651_));
  AOI22  g01649(.A0(new_n2651_), .A1(new_n2650_), .B0(new_n2633_), .B1(new_n2638_), .Y(new_n2652_));
  NAND2  g01650(.A(\A[833] ), .B(new_n2643_), .Y(new_n2653_));
  AOI21  g01651(.A0(new_n2641_), .A1(\A[832] ), .B0(new_n2645_), .Y(new_n2654_));
  AOI22  g01652(.A0(new_n2654_), .A1(new_n2653_), .B0(new_n2628_), .B1(new_n2645_), .Y(new_n2655_));
  XOR2   g01653(.A(new_n2655_), .B(new_n2652_), .Y(new_n2656_));
  NAND4  g01654(.A(new_n2656_), .B(new_n2649_), .C(new_n2648_), .D(new_n2612_), .Y(new_n2657_));
  NOR2   g01655(.A(new_n2632_), .B(new_n2631_), .Y(new_n2658_));
  AOI21  g01656(.A0(new_n2633_), .A1(\A[831] ), .B0(new_n2658_), .Y(new_n2659_));
  XOR2   g01657(.A(new_n2659_), .B(new_n2630_), .Y(new_n2660_));
  NAND2  g01658(.A(new_n2647_), .B(new_n2640_), .Y(new_n2661_));
  NAND2  g01659(.A(new_n2635_), .B(new_n2630_), .Y(new_n2662_));
  OAI21  g01660(.A0(new_n2661_), .A1(new_n2660_), .B0(new_n2662_), .Y(new_n2663_));
  NOR2   g01661(.A(new_n2655_), .B(new_n2652_), .Y(new_n2664_));
  XOR2   g01662(.A(new_n2664_), .B(new_n2660_), .Y(new_n2665_));
  AOI21  g01663(.A0(new_n2656_), .A1(new_n2663_), .B0(new_n2665_), .Y(new_n2666_));
  XOR2   g01664(.A(new_n2666_), .B(new_n2657_), .Y(new_n2667_));
  XOR2   g01665(.A(new_n2635_), .B(new_n2630_), .Y(new_n2668_));
  XOR2   g01666(.A(new_n2664_), .B(new_n2668_), .Y(new_n2669_));
  AOI211 g01667(.A0(new_n2606_), .A1(new_n2605_), .B(new_n2609_), .C(new_n2621_), .Y(new_n2670_));
  NAND2  g01668(.A(new_n2656_), .B(new_n2612_), .Y(new_n2671_));
  AOI211 g01669(.A0(new_n2669_), .A1(new_n2663_), .B(new_n2671_), .C(new_n2670_), .Y(new_n2672_));
  NOR2   g01670(.A(new_n2666_), .B(new_n2672_), .Y(new_n2673_));
  AOI221 g01671(.A0(new_n2655_), .A1(new_n2652_), .C0(new_n2659_), .B0(new_n2629_), .B1(new_n2627_), .Y(new_n2674_));
  NOR4   g01672(.A(new_n2674_), .B(new_n2671_), .C(new_n2670_), .D(new_n2665_), .Y(new_n2675_));
  OAI21  g01673(.A0(new_n2675_), .A1(new_n2673_), .B0(new_n2626_), .Y(new_n2676_));
  OAI21  g01674(.A0(new_n2667_), .A1(new_n2626_), .B0(new_n2676_), .Y(new_n2677_));
  INV    g01675(.A(\A[836] ), .Y(new_n2678_));
  NOR2   g01676(.A(new_n2678_), .B(\A[835] ), .Y(new_n2679_));
  INV    g01677(.A(\A[835] ), .Y(new_n2680_));
  OAI21  g01678(.A0(\A[836] ), .A1(new_n2680_), .B0(\A[837] ), .Y(new_n2681_));
  XOR2   g01679(.A(\A[836] ), .B(new_n2680_), .Y(new_n2682_));
  OAI22  g01680(.A0(new_n2682_), .A1(\A[837] ), .B0(new_n2681_), .B1(new_n2679_), .Y(new_n2683_));
  INV    g01681(.A(\A[839] ), .Y(new_n2684_));
  NOR2   g01682(.A(new_n2684_), .B(\A[838] ), .Y(new_n2685_));
  INV    g01683(.A(\A[838] ), .Y(new_n2686_));
  OAI21  g01684(.A0(\A[839] ), .A1(new_n2686_), .B0(\A[840] ), .Y(new_n2687_));
  XOR2   g01685(.A(\A[839] ), .B(new_n2686_), .Y(new_n2688_));
  OAI22  g01686(.A0(new_n2688_), .A1(\A[840] ), .B0(new_n2687_), .B1(new_n2685_), .Y(new_n2689_));
  NAND2  g01687(.A(new_n2689_), .B(new_n2683_), .Y(new_n2690_));
  NAND2  g01688(.A(\A[839] ), .B(\A[838] ), .Y(new_n2691_));
  XOR2   g01689(.A(\A[839] ), .B(\A[838] ), .Y(new_n2692_));
  NAND2  g01690(.A(new_n2692_), .B(\A[840] ), .Y(new_n2693_));
  NAND2  g01691(.A(new_n2693_), .B(new_n2691_), .Y(new_n2694_));
  XOR2   g01692(.A(\A[836] ), .B(\A[835] ), .Y(new_n2695_));
  NOR2   g01693(.A(new_n2678_), .B(new_n2680_), .Y(new_n2696_));
  AOI21  g01694(.A0(new_n2695_), .A1(\A[837] ), .B0(new_n2696_), .Y(new_n2697_));
  XOR2   g01695(.A(new_n2697_), .B(new_n2694_), .Y(new_n2698_));
  XOR2   g01696(.A(new_n2698_), .B(new_n2690_), .Y(new_n2699_));
  INV    g01697(.A(\A[837] ), .Y(new_n2700_));
  NAND2  g01698(.A(\A[836] ), .B(new_n2680_), .Y(new_n2701_));
  AOI21  g01699(.A0(new_n2678_), .A1(\A[835] ), .B0(new_n2700_), .Y(new_n2702_));
  AOI22  g01700(.A0(new_n2695_), .A1(new_n2700_), .B0(new_n2702_), .B1(new_n2701_), .Y(new_n2703_));
  INV    g01701(.A(\A[840] ), .Y(new_n2704_));
  NAND2  g01702(.A(\A[839] ), .B(new_n2686_), .Y(new_n2705_));
  AOI21  g01703(.A0(new_n2684_), .A1(\A[838] ), .B0(new_n2704_), .Y(new_n2706_));
  AOI22  g01704(.A0(new_n2692_), .A1(new_n2704_), .B0(new_n2706_), .B1(new_n2705_), .Y(new_n2707_));
  XOR2   g01705(.A(new_n2707_), .B(new_n2703_), .Y(new_n2708_));
  INV    g01706(.A(new_n2708_), .Y(new_n2709_));
  NAND2  g01707(.A(\A[836] ), .B(\A[835] ), .Y(new_n2710_));
  OAI21  g01708(.A0(new_n2682_), .A1(new_n2700_), .B0(new_n2710_), .Y(new_n2711_));
  NOR2   g01709(.A(new_n2698_), .B(new_n2690_), .Y(new_n2712_));
  AOI21  g01710(.A0(new_n2711_), .A1(new_n2694_), .B0(new_n2712_), .Y(new_n2713_));
  OAI21  g01711(.A0(new_n2713_), .A1(new_n2709_), .B0(new_n2699_), .Y(new_n2714_));
  INV    g01712(.A(\A[844] ), .Y(new_n2715_));
  INV    g01713(.A(\A[845] ), .Y(new_n2716_));
  NOR2   g01714(.A(new_n2716_), .B(new_n2715_), .Y(new_n2717_));
  XOR2   g01715(.A(\A[845] ), .B(\A[844] ), .Y(new_n2718_));
  AOI21  g01716(.A0(new_n2718_), .A1(\A[846] ), .B0(new_n2717_), .Y(new_n2719_));
  INV    g01717(.A(\A[841] ), .Y(new_n2720_));
  INV    g01718(.A(\A[842] ), .Y(new_n2721_));
  NOR2   g01719(.A(new_n2721_), .B(new_n2720_), .Y(new_n2722_));
  XOR2   g01720(.A(\A[842] ), .B(\A[841] ), .Y(new_n2723_));
  AOI21  g01721(.A0(new_n2723_), .A1(\A[843] ), .B0(new_n2722_), .Y(new_n2724_));
  INV    g01722(.A(\A[843] ), .Y(new_n2725_));
  NAND2  g01723(.A(\A[842] ), .B(new_n2720_), .Y(new_n2726_));
  AOI21  g01724(.A0(new_n2721_), .A1(\A[841] ), .B0(new_n2725_), .Y(new_n2727_));
  AOI22  g01725(.A0(new_n2727_), .A1(new_n2726_), .B0(new_n2723_), .B1(new_n2725_), .Y(new_n2728_));
  INV    g01726(.A(\A[846] ), .Y(new_n2729_));
  NAND2  g01727(.A(\A[845] ), .B(new_n2715_), .Y(new_n2730_));
  AOI21  g01728(.A0(new_n2716_), .A1(\A[844] ), .B0(new_n2729_), .Y(new_n2731_));
  AOI22  g01729(.A0(new_n2731_), .A1(new_n2730_), .B0(new_n2718_), .B1(new_n2729_), .Y(new_n2732_));
  NOR4   g01730(.A(new_n2732_), .B(new_n2728_), .C(new_n2724_), .D(new_n2719_), .Y(new_n2733_));
  AOI211 g01731(.A0(new_n2693_), .A1(new_n2691_), .B(new_n2697_), .C(new_n2690_), .Y(new_n2734_));
  XOR2   g01732(.A(new_n2732_), .B(new_n2728_), .Y(new_n2735_));
  NAND2  g01733(.A(new_n2735_), .B(new_n2708_), .Y(new_n2736_));
  NOR3   g01734(.A(new_n2736_), .B(new_n2734_), .C(new_n2733_), .Y(new_n2737_));
  NAND2  g01735(.A(new_n2718_), .B(\A[846] ), .Y(new_n2738_));
  OAI21  g01736(.A0(new_n2716_), .A1(new_n2715_), .B0(new_n2738_), .Y(new_n2739_));
  XOR2   g01737(.A(new_n2724_), .B(new_n2739_), .Y(new_n2740_));
  NOR2   g01738(.A(new_n2721_), .B(\A[841] ), .Y(new_n2741_));
  OAI21  g01739(.A0(\A[842] ), .A1(new_n2720_), .B0(\A[843] ), .Y(new_n2742_));
  NAND2  g01740(.A(new_n2723_), .B(new_n2725_), .Y(new_n2743_));
  OAI21  g01741(.A0(new_n2742_), .A1(new_n2741_), .B0(new_n2743_), .Y(new_n2744_));
  NOR2   g01742(.A(new_n2716_), .B(\A[844] ), .Y(new_n2745_));
  OAI21  g01743(.A0(\A[845] ), .A1(new_n2715_), .B0(\A[846] ), .Y(new_n2746_));
  NAND2  g01744(.A(new_n2718_), .B(new_n2729_), .Y(new_n2747_));
  OAI21  g01745(.A0(new_n2746_), .A1(new_n2745_), .B0(new_n2747_), .Y(new_n2748_));
  NAND2  g01746(.A(new_n2748_), .B(new_n2744_), .Y(new_n2749_));
  NAND2  g01747(.A(new_n2723_), .B(\A[843] ), .Y(new_n2750_));
  OAI21  g01748(.A0(new_n2721_), .A1(new_n2720_), .B0(new_n2750_), .Y(new_n2751_));
  NAND2  g01749(.A(new_n2751_), .B(new_n2739_), .Y(new_n2752_));
  OAI21  g01750(.A0(new_n2749_), .A1(new_n2740_), .B0(new_n2752_), .Y(new_n2753_));
  NOR2   g01751(.A(new_n2732_), .B(new_n2728_), .Y(new_n2754_));
  XOR2   g01752(.A(new_n2754_), .B(new_n2740_), .Y(new_n2755_));
  AOI21  g01753(.A0(new_n2735_), .A1(new_n2753_), .B0(new_n2755_), .Y(new_n2756_));
  XOR2   g01754(.A(new_n2756_), .B(new_n2737_), .Y(new_n2757_));
  NAND2  g01755(.A(new_n2757_), .B(new_n2714_), .Y(new_n2758_));
  NOR2   g01756(.A(new_n2707_), .B(new_n2703_), .Y(new_n2759_));
  XOR2   g01757(.A(new_n2698_), .B(new_n2759_), .Y(new_n2760_));
  NAND2  g01758(.A(new_n2711_), .B(new_n2694_), .Y(new_n2761_));
  OAI21  g01759(.A0(new_n2698_), .A1(new_n2690_), .B0(new_n2761_), .Y(new_n2762_));
  AOI21  g01760(.A0(new_n2762_), .A1(new_n2708_), .B0(new_n2760_), .Y(new_n2763_));
  NOR2   g01761(.A(new_n2756_), .B(new_n2737_), .Y(new_n2764_));
  AOI211 g01762(.A0(new_n2732_), .A1(new_n2728_), .B(new_n2724_), .C(new_n2719_), .Y(new_n2765_));
  NOR4   g01763(.A(new_n2765_), .B(new_n2736_), .C(new_n2734_), .D(new_n2755_), .Y(new_n2766_));
  OAI21  g01764(.A0(new_n2766_), .A1(new_n2764_), .B0(new_n2763_), .Y(new_n2767_));
  XOR2   g01765(.A(new_n2732_), .B(new_n2744_), .Y(new_n2768_));
  NOR2   g01766(.A(new_n2768_), .B(new_n2733_), .Y(new_n2769_));
  NAND4  g01767(.A(new_n2711_), .B(new_n2694_), .C(new_n2689_), .D(new_n2683_), .Y(new_n2770_));
  NAND2  g01768(.A(new_n2770_), .B(new_n2708_), .Y(new_n2771_));
  XOR2   g01769(.A(new_n2771_), .B(new_n2769_), .Y(new_n2772_));
  NAND2  g01770(.A(new_n2656_), .B(new_n2648_), .Y(new_n2773_));
  NAND3  g01771(.A(new_n2773_), .B(new_n2649_), .C(new_n2612_), .Y(new_n2774_));
  NAND2  g01772(.A(new_n2649_), .B(new_n2612_), .Y(new_n2775_));
  NAND3  g01773(.A(new_n2775_), .B(new_n2656_), .C(new_n2648_), .Y(new_n2776_));
  AOI21  g01774(.A0(new_n2776_), .A1(new_n2774_), .B0(new_n2772_), .Y(new_n2777_));
  NAND3  g01775(.A(new_n2777_), .B(new_n2767_), .C(new_n2758_), .Y(new_n2778_));
  NAND4  g01776(.A(new_n2748_), .B(new_n2744_), .C(new_n2751_), .D(new_n2739_), .Y(new_n2779_));
  NAND4  g01777(.A(new_n2735_), .B(new_n2770_), .C(new_n2779_), .D(new_n2708_), .Y(new_n2780_));
  XOR2   g01778(.A(new_n2756_), .B(new_n2780_), .Y(new_n2781_));
  NOR2   g01779(.A(new_n2781_), .B(new_n2763_), .Y(new_n2782_));
  XOR2   g01780(.A(new_n2751_), .B(new_n2739_), .Y(new_n2783_));
  NOR2   g01781(.A(new_n2724_), .B(new_n2719_), .Y(new_n2784_));
  AOI21  g01782(.A0(new_n2754_), .A1(new_n2783_), .B0(new_n2784_), .Y(new_n2785_));
  XOR2   g01783(.A(new_n2754_), .B(new_n2783_), .Y(new_n2786_));
  OAI21  g01784(.A0(new_n2768_), .A1(new_n2785_), .B0(new_n2786_), .Y(new_n2787_));
  AOI21  g01785(.A0(new_n2787_), .A1(new_n2780_), .B0(new_n2766_), .Y(new_n2788_));
  NOR2   g01786(.A(new_n2788_), .B(new_n2714_), .Y(new_n2789_));
  NAND2  g01787(.A(new_n2735_), .B(new_n2779_), .Y(new_n2790_));
  XOR2   g01788(.A(new_n2771_), .B(new_n2790_), .Y(new_n2791_));
  XOR2   g01789(.A(new_n2775_), .B(new_n2773_), .Y(new_n2792_));
  NAND2  g01790(.A(new_n2792_), .B(new_n2791_), .Y(new_n2793_));
  OAI21  g01791(.A0(new_n2789_), .A1(new_n2782_), .B0(new_n2793_), .Y(new_n2794_));
  AOI21  g01792(.A0(new_n2794_), .A1(new_n2778_), .B0(new_n2677_), .Y(new_n2795_));
  NOR2   g01793(.A(new_n2667_), .B(new_n2626_), .Y(new_n2796_));
  AOI21  g01794(.A0(new_n2629_), .A1(new_n2627_), .B0(new_n2659_), .Y(new_n2797_));
  AOI21  g01795(.A0(new_n2664_), .A1(new_n2668_), .B0(new_n2797_), .Y(new_n2798_));
  XOR2   g01796(.A(new_n2655_), .B(new_n2640_), .Y(new_n2799_));
  OAI21  g01797(.A0(new_n2799_), .A1(new_n2798_), .B0(new_n2669_), .Y(new_n2800_));
  AOI21  g01798(.A0(new_n2800_), .A1(new_n2657_), .B0(new_n2675_), .Y(new_n2801_));
  AOI211 g01799(.A0(new_n2625_), .A1(new_n2612_), .B(new_n2801_), .C(new_n2611_), .Y(new_n2802_));
  NOR2   g01800(.A(new_n2802_), .B(new_n2796_), .Y(new_n2803_));
  NAND3  g01801(.A(new_n2793_), .B(new_n2767_), .C(new_n2758_), .Y(new_n2804_));
  OAI21  g01802(.A0(new_n2789_), .A1(new_n2782_), .B0(new_n2777_), .Y(new_n2805_));
  AOI21  g01803(.A0(new_n2805_), .A1(new_n2804_), .B0(new_n2803_), .Y(new_n2806_));
  XOR2   g01804(.A(new_n2792_), .B(new_n2772_), .Y(new_n2807_));
  XOR2   g01805(.A(new_n2522_), .B(new_n2472_), .Y(new_n2808_));
  NOR2   g01806(.A(new_n2808_), .B(new_n2807_), .Y(new_n2809_));
  INV    g01807(.A(new_n2809_), .Y(new_n2810_));
  NOR3   g01808(.A(new_n2810_), .B(new_n2806_), .C(new_n2795_), .Y(new_n2811_));
  NAND2  g01809(.A(new_n2794_), .B(new_n2778_), .Y(new_n2812_));
  NAND2  g01810(.A(new_n2812_), .B(new_n2803_), .Y(new_n2813_));
  NAND2  g01811(.A(new_n2805_), .B(new_n2804_), .Y(new_n2814_));
  NAND2  g01812(.A(new_n2814_), .B(new_n2677_), .Y(new_n2815_));
  AOI21  g01813(.A0(new_n2815_), .A1(new_n2813_), .B0(new_n2809_), .Y(new_n2816_));
  OAI21  g01814(.A0(new_n2816_), .A1(new_n2811_), .B0(new_n2589_), .Y(new_n2817_));
  OAI21  g01815(.A0(new_n2524_), .A1(new_n2513_), .B0(new_n2585_), .Y(new_n2818_));
  OAI21  g01816(.A0(new_n2468_), .A1(new_n2455_), .B0(new_n2512_), .Y(new_n2819_));
  NOR2   g01817(.A(new_n2819_), .B(new_n2450_), .Y(new_n2820_));
  AOI21  g01818(.A0(new_n2519_), .A1(new_n2517_), .B0(new_n2512_), .Y(new_n2821_));
  OAI22  g01819(.A0(new_n2821_), .A1(new_n2820_), .B0(new_n2584_), .B1(new_n2579_), .Y(new_n2822_));
  NAND2  g01820(.A(new_n2822_), .B(new_n2818_), .Y(new_n2823_));
  NOR3   g01821(.A(new_n2809_), .B(new_n2806_), .C(new_n2795_), .Y(new_n2824_));
  AOI21  g01822(.A0(new_n2815_), .A1(new_n2813_), .B0(new_n2810_), .Y(new_n2825_));
  OAI21  g01823(.A0(new_n2825_), .A1(new_n2824_), .B0(new_n2823_), .Y(new_n2826_));
  XOR2   g01824(.A(new_n2808_), .B(new_n2807_), .Y(new_n2827_));
  XOR2   g01825(.A(new_n2362_), .B(new_n2360_), .Y(new_n2828_));
  NAND2  g01826(.A(new_n2828_), .B(new_n2827_), .Y(new_n2829_));
  INV    g01827(.A(new_n2829_), .Y(new_n2830_));
  NAND3  g01828(.A(new_n2830_), .B(new_n2826_), .C(new_n2817_), .Y(new_n2831_));
  NAND3  g01829(.A(new_n2809_), .B(new_n2815_), .C(new_n2813_), .Y(new_n2832_));
  OAI21  g01830(.A0(new_n2806_), .A1(new_n2795_), .B0(new_n2810_), .Y(new_n2833_));
  AOI21  g01831(.A0(new_n2833_), .A1(new_n2832_), .B0(new_n2823_), .Y(new_n2834_));
  NAND3  g01832(.A(new_n2810_), .B(new_n2815_), .C(new_n2813_), .Y(new_n2835_));
  OAI21  g01833(.A0(new_n2806_), .A1(new_n2795_), .B0(new_n2809_), .Y(new_n2836_));
  AOI21  g01834(.A0(new_n2836_), .A1(new_n2835_), .B0(new_n2589_), .Y(new_n2837_));
  OAI21  g01835(.A0(new_n2837_), .A1(new_n2834_), .B0(new_n2829_), .Y(new_n2838_));
  AOI21  g01836(.A0(new_n2838_), .A1(new_n2831_), .B0(new_n2372_), .Y(new_n2839_));
  NAND2  g01837(.A(new_n2353_), .B(new_n2337_), .Y(new_n2840_));
  NAND2  g01838(.A(new_n2840_), .B(new_n2356_), .Y(new_n2841_));
  NOR2   g01839(.A(new_n2364_), .B(new_n2359_), .Y(new_n2842_));
  NAND2  g01840(.A(new_n2842_), .B(new_n2841_), .Y(new_n2843_));
  OAI21  g01841(.A0(new_n2366_), .A1(new_n2363_), .B0(new_n2843_), .Y(new_n2844_));
  NOR2   g01842(.A(new_n2363_), .B(new_n2359_), .Y(new_n2845_));
  NAND2  g01843(.A(new_n2845_), .B(new_n2841_), .Y(new_n2846_));
  OAI21  g01844(.A0(new_n2359_), .A1(new_n2354_), .B0(new_n2363_), .Y(new_n2847_));
  AOI21  g01845(.A0(new_n2847_), .A1(new_n2846_), .B0(new_n2144_), .Y(new_n2848_));
  AOI21  g01846(.A0(new_n2144_), .A1(new_n2844_), .B0(new_n2848_), .Y(new_n2849_));
  NAND3  g01847(.A(new_n2829_), .B(new_n2826_), .C(new_n2817_), .Y(new_n2850_));
  OAI21  g01848(.A0(new_n2837_), .A1(new_n2834_), .B0(new_n2830_), .Y(new_n2851_));
  AOI21  g01849(.A0(new_n2851_), .A1(new_n2850_), .B0(new_n2849_), .Y(new_n2852_));
  INV    g01850(.A(new_n2828_), .Y(new_n2853_));
  XOR2   g01851(.A(new_n2853_), .B(new_n2827_), .Y(new_n2854_));
  XOR2   g01852(.A(new_n1620_), .B(new_n1457_), .Y(new_n2855_));
  NOR2   g01853(.A(new_n2855_), .B(new_n2854_), .Y(new_n2856_));
  INV    g01854(.A(new_n2856_), .Y(new_n2857_));
  NOR3   g01855(.A(new_n2857_), .B(new_n2852_), .C(new_n2839_), .Y(new_n2858_));
  NOR3   g01856(.A(new_n2829_), .B(new_n2837_), .C(new_n2834_), .Y(new_n2859_));
  AOI21  g01857(.A0(new_n2826_), .A1(new_n2817_), .B0(new_n2830_), .Y(new_n2860_));
  OAI21  g01858(.A0(new_n2860_), .A1(new_n2859_), .B0(new_n2849_), .Y(new_n2861_));
  NOR3   g01859(.A(new_n2830_), .B(new_n2837_), .C(new_n2834_), .Y(new_n2862_));
  AOI21  g01860(.A0(new_n2826_), .A1(new_n2817_), .B0(new_n2829_), .Y(new_n2863_));
  OAI21  g01861(.A0(new_n2863_), .A1(new_n2862_), .B0(new_n2372_), .Y(new_n2864_));
  AOI21  g01862(.A0(new_n2864_), .A1(new_n2861_), .B0(new_n2856_), .Y(new_n2865_));
  OAI21  g01863(.A0(new_n2865_), .A1(new_n2858_), .B0(new_n1929_), .Y(new_n2866_));
  NOR3   g01864(.A(new_n1629_), .B(new_n1628_), .C(new_n1625_), .Y(new_n2867_));
  AOI21  g01865(.A0(new_n1456_), .A1(new_n1447_), .B0(new_n1621_), .Y(new_n2868_));
  OAI21  g01866(.A0(new_n2868_), .A1(new_n2867_), .B0(new_n1925_), .Y(new_n2869_));
  NOR3   g01867(.A(new_n1621_), .B(new_n1628_), .C(new_n1625_), .Y(new_n2870_));
  AOI21  g01868(.A0(new_n1456_), .A1(new_n1447_), .B0(new_n1629_), .Y(new_n2871_));
  OAI21  g01869(.A0(new_n2871_), .A1(new_n2870_), .B0(new_n1917_), .Y(new_n2872_));
  NAND2  g01870(.A(new_n2872_), .B(new_n2869_), .Y(new_n2873_));
  NOR3   g01871(.A(new_n2856_), .B(new_n2852_), .C(new_n2839_), .Y(new_n2874_));
  AOI21  g01872(.A0(new_n2864_), .A1(new_n2861_), .B0(new_n2857_), .Y(new_n2875_));
  OAI21  g01873(.A0(new_n2875_), .A1(new_n2874_), .B0(new_n2873_), .Y(new_n2876_));
  INV    g01874(.A(\A[471] ), .Y(new_n2877_));
  INV    g01875(.A(\A[470] ), .Y(new_n2878_));
  NAND2  g01876(.A(new_n2878_), .B(\A[469] ), .Y(new_n2879_));
  INV    g01877(.A(\A[469] ), .Y(new_n2880_));
  AOI21  g01878(.A0(\A[470] ), .A1(new_n2880_), .B0(new_n2877_), .Y(new_n2881_));
  XOR2   g01879(.A(\A[470] ), .B(\A[469] ), .Y(new_n2882_));
  AOI22  g01880(.A0(new_n2882_), .A1(new_n2877_), .B0(new_n2881_), .B1(new_n2879_), .Y(new_n2883_));
  INV    g01881(.A(\A[474] ), .Y(new_n2884_));
  INV    g01882(.A(\A[473] ), .Y(new_n2885_));
  NAND2  g01883(.A(new_n2885_), .B(\A[472] ), .Y(new_n2886_));
  INV    g01884(.A(\A[472] ), .Y(new_n2887_));
  AOI21  g01885(.A0(\A[473] ), .A1(new_n2887_), .B0(new_n2884_), .Y(new_n2888_));
  XOR2   g01886(.A(\A[473] ), .B(\A[472] ), .Y(new_n2889_));
  AOI22  g01887(.A0(new_n2889_), .A1(new_n2884_), .B0(new_n2888_), .B1(new_n2886_), .Y(new_n2890_));
  NOR2   g01888(.A(new_n2885_), .B(new_n2887_), .Y(new_n2891_));
  AOI21  g01889(.A0(new_n2889_), .A1(\A[474] ), .B0(new_n2891_), .Y(new_n2892_));
  NOR2   g01890(.A(new_n2878_), .B(new_n2880_), .Y(new_n2893_));
  AOI21  g01891(.A0(new_n2882_), .A1(\A[471] ), .B0(new_n2893_), .Y(new_n2894_));
  XOR2   g01892(.A(new_n2890_), .B(new_n2883_), .Y(new_n2895_));
  INV    g01893(.A(new_n2895_), .Y(new_n2896_));
  INV    g01894(.A(\A[468] ), .Y(new_n2897_));
  INV    g01895(.A(\A[467] ), .Y(new_n2898_));
  NAND2  g01896(.A(new_n2898_), .B(\A[466] ), .Y(new_n2899_));
  INV    g01897(.A(\A[466] ), .Y(new_n2900_));
  AOI21  g01898(.A0(\A[467] ), .A1(new_n2900_), .B0(new_n2897_), .Y(new_n2901_));
  XOR2   g01899(.A(\A[467] ), .B(\A[466] ), .Y(new_n2902_));
  AOI22  g01900(.A0(new_n2902_), .A1(new_n2897_), .B0(new_n2901_), .B1(new_n2899_), .Y(new_n2903_));
  INV    g01901(.A(\A[465] ), .Y(new_n2904_));
  INV    g01902(.A(\A[464] ), .Y(new_n2905_));
  NAND2  g01903(.A(new_n2905_), .B(\A[463] ), .Y(new_n2906_));
  INV    g01904(.A(\A[463] ), .Y(new_n2907_));
  AOI21  g01905(.A0(\A[464] ), .A1(new_n2907_), .B0(new_n2904_), .Y(new_n2908_));
  XOR2   g01906(.A(\A[464] ), .B(\A[463] ), .Y(new_n2909_));
  AOI22  g01907(.A0(new_n2909_), .A1(new_n2904_), .B0(new_n2908_), .B1(new_n2906_), .Y(new_n2910_));
  XOR2   g01908(.A(new_n2910_), .B(new_n2903_), .Y(new_n2911_));
  NOR2   g01909(.A(\A[467] ), .B(new_n2900_), .Y(new_n2912_));
  OAI21  g01910(.A0(new_n2898_), .A1(\A[466] ), .B0(\A[468] ), .Y(new_n2913_));
  XOR2   g01911(.A(\A[467] ), .B(new_n2900_), .Y(new_n2914_));
  OAI22  g01912(.A0(new_n2914_), .A1(\A[468] ), .B0(new_n2913_), .B1(new_n2912_), .Y(new_n2915_));
  NOR2   g01913(.A(\A[464] ), .B(new_n2907_), .Y(new_n2916_));
  OAI21  g01914(.A0(new_n2905_), .A1(\A[463] ), .B0(\A[465] ), .Y(new_n2917_));
  XOR2   g01915(.A(\A[464] ), .B(new_n2907_), .Y(new_n2918_));
  OAI22  g01916(.A0(new_n2918_), .A1(\A[465] ), .B0(new_n2917_), .B1(new_n2916_), .Y(new_n2919_));
  NAND2  g01917(.A(\A[467] ), .B(\A[466] ), .Y(new_n2920_));
  NAND2  g01918(.A(new_n2902_), .B(\A[468] ), .Y(new_n2921_));
  NAND2  g01919(.A(new_n2921_), .B(new_n2920_), .Y(new_n2922_));
  NAND2  g01920(.A(\A[464] ), .B(\A[463] ), .Y(new_n2923_));
  OAI21  g01921(.A0(new_n2918_), .A1(new_n2904_), .B0(new_n2923_), .Y(new_n2924_));
  NAND4  g01922(.A(new_n2924_), .B(new_n2922_), .C(new_n2919_), .D(new_n2915_), .Y(new_n2925_));
  NAND2  g01923(.A(new_n2925_), .B(new_n2911_), .Y(new_n2926_));
  XOR2   g01924(.A(new_n2926_), .B(new_n2896_), .Y(new_n2927_));
  INV    g01925(.A(\A[483] ), .Y(new_n2928_));
  INV    g01926(.A(\A[482] ), .Y(new_n2929_));
  NAND2  g01927(.A(new_n2929_), .B(\A[481] ), .Y(new_n2930_));
  INV    g01928(.A(\A[481] ), .Y(new_n2931_));
  AOI21  g01929(.A0(\A[482] ), .A1(new_n2931_), .B0(new_n2928_), .Y(new_n2932_));
  XOR2   g01930(.A(\A[482] ), .B(\A[481] ), .Y(new_n2933_));
  AOI22  g01931(.A0(new_n2933_), .A1(new_n2928_), .B0(new_n2932_), .B1(new_n2930_), .Y(new_n2934_));
  INV    g01932(.A(\A[486] ), .Y(new_n2935_));
  INV    g01933(.A(\A[485] ), .Y(new_n2936_));
  NAND2  g01934(.A(new_n2936_), .B(\A[484] ), .Y(new_n2937_));
  INV    g01935(.A(\A[484] ), .Y(new_n2938_));
  AOI21  g01936(.A0(\A[485] ), .A1(new_n2938_), .B0(new_n2935_), .Y(new_n2939_));
  XOR2   g01937(.A(\A[485] ), .B(\A[484] ), .Y(new_n2940_));
  AOI22  g01938(.A0(new_n2940_), .A1(new_n2935_), .B0(new_n2939_), .B1(new_n2937_), .Y(new_n2941_));
  NOR2   g01939(.A(new_n2936_), .B(new_n2938_), .Y(new_n2942_));
  AOI21  g01940(.A0(new_n2940_), .A1(\A[486] ), .B0(new_n2942_), .Y(new_n2943_));
  NOR2   g01941(.A(new_n2929_), .B(new_n2931_), .Y(new_n2944_));
  AOI21  g01942(.A0(new_n2933_), .A1(\A[483] ), .B0(new_n2944_), .Y(new_n2945_));
  XOR2   g01943(.A(new_n2941_), .B(new_n2934_), .Y(new_n2946_));
  INV    g01944(.A(\A[477] ), .Y(new_n2947_));
  INV    g01945(.A(\A[476] ), .Y(new_n2948_));
  NAND2  g01946(.A(new_n2948_), .B(\A[475] ), .Y(new_n2949_));
  INV    g01947(.A(\A[475] ), .Y(new_n2950_));
  AOI21  g01948(.A0(\A[476] ), .A1(new_n2950_), .B0(new_n2947_), .Y(new_n2951_));
  XOR2   g01949(.A(\A[476] ), .B(\A[475] ), .Y(new_n2952_));
  AOI22  g01950(.A0(new_n2952_), .A1(new_n2947_), .B0(new_n2951_), .B1(new_n2949_), .Y(new_n2953_));
  INV    g01951(.A(\A[480] ), .Y(new_n2954_));
  INV    g01952(.A(\A[479] ), .Y(new_n2955_));
  NAND2  g01953(.A(new_n2955_), .B(\A[478] ), .Y(new_n2956_));
  INV    g01954(.A(\A[478] ), .Y(new_n2957_));
  AOI21  g01955(.A0(\A[479] ), .A1(new_n2957_), .B0(new_n2954_), .Y(new_n2958_));
  XOR2   g01956(.A(\A[479] ), .B(\A[478] ), .Y(new_n2959_));
  AOI22  g01957(.A0(new_n2959_), .A1(new_n2954_), .B0(new_n2958_), .B1(new_n2956_), .Y(new_n2960_));
  NOR2   g01958(.A(new_n2955_), .B(new_n2957_), .Y(new_n2961_));
  AOI21  g01959(.A0(new_n2959_), .A1(\A[480] ), .B0(new_n2961_), .Y(new_n2962_));
  NOR2   g01960(.A(new_n2948_), .B(new_n2950_), .Y(new_n2963_));
  AOI21  g01961(.A0(new_n2952_), .A1(\A[477] ), .B0(new_n2963_), .Y(new_n2964_));
  XOR2   g01962(.A(new_n2960_), .B(new_n2953_), .Y(new_n2965_));
  XOR2   g01963(.A(new_n2965_), .B(new_n2946_), .Y(new_n2966_));
  INV    g01964(.A(new_n2966_), .Y(new_n2967_));
  XOR2   g01965(.A(new_n2967_), .B(new_n2927_), .Y(new_n2968_));
  INV    g01966(.A(new_n2968_), .Y(new_n2969_));
  INV    g01967(.A(\A[507] ), .Y(new_n2970_));
  INV    g01968(.A(\A[506] ), .Y(new_n2971_));
  NAND2  g01969(.A(new_n2971_), .B(\A[505] ), .Y(new_n2972_));
  INV    g01970(.A(\A[505] ), .Y(new_n2973_));
  AOI21  g01971(.A0(\A[506] ), .A1(new_n2973_), .B0(new_n2970_), .Y(new_n2974_));
  XOR2   g01972(.A(\A[506] ), .B(\A[505] ), .Y(new_n2975_));
  AOI22  g01973(.A0(new_n2975_), .A1(new_n2970_), .B0(new_n2974_), .B1(new_n2972_), .Y(new_n2976_));
  INV    g01974(.A(\A[510] ), .Y(new_n2977_));
  INV    g01975(.A(\A[509] ), .Y(new_n2978_));
  NAND2  g01976(.A(new_n2978_), .B(\A[508] ), .Y(new_n2979_));
  INV    g01977(.A(\A[508] ), .Y(new_n2980_));
  AOI21  g01978(.A0(\A[509] ), .A1(new_n2980_), .B0(new_n2977_), .Y(new_n2981_));
  XOR2   g01979(.A(\A[509] ), .B(\A[508] ), .Y(new_n2982_));
  AOI22  g01980(.A0(new_n2982_), .A1(new_n2977_), .B0(new_n2981_), .B1(new_n2979_), .Y(new_n2983_));
  NOR2   g01981(.A(new_n2978_), .B(new_n2980_), .Y(new_n2984_));
  AOI21  g01982(.A0(new_n2982_), .A1(\A[510] ), .B0(new_n2984_), .Y(new_n2985_));
  NOR2   g01983(.A(new_n2971_), .B(new_n2973_), .Y(new_n2986_));
  AOI21  g01984(.A0(new_n2975_), .A1(\A[507] ), .B0(new_n2986_), .Y(new_n2987_));
  XOR2   g01985(.A(new_n2983_), .B(new_n2976_), .Y(new_n2988_));
  INV    g01986(.A(\A[501] ), .Y(new_n2989_));
  INV    g01987(.A(\A[500] ), .Y(new_n2990_));
  NAND2  g01988(.A(new_n2990_), .B(\A[499] ), .Y(new_n2991_));
  INV    g01989(.A(\A[499] ), .Y(new_n2992_));
  AOI21  g01990(.A0(\A[500] ), .A1(new_n2992_), .B0(new_n2989_), .Y(new_n2993_));
  XOR2   g01991(.A(\A[500] ), .B(\A[499] ), .Y(new_n2994_));
  AOI22  g01992(.A0(new_n2994_), .A1(new_n2989_), .B0(new_n2993_), .B1(new_n2991_), .Y(new_n2995_));
  INV    g01993(.A(\A[504] ), .Y(new_n2996_));
  INV    g01994(.A(\A[503] ), .Y(new_n2997_));
  NAND2  g01995(.A(new_n2997_), .B(\A[502] ), .Y(new_n2998_));
  INV    g01996(.A(\A[502] ), .Y(new_n2999_));
  AOI21  g01997(.A0(\A[503] ), .A1(new_n2999_), .B0(new_n2996_), .Y(new_n3000_));
  XOR2   g01998(.A(\A[503] ), .B(\A[502] ), .Y(new_n3001_));
  AOI22  g01999(.A0(new_n3001_), .A1(new_n2996_), .B0(new_n3000_), .B1(new_n2998_), .Y(new_n3002_));
  NOR2   g02000(.A(new_n2997_), .B(new_n2999_), .Y(new_n3003_));
  AOI21  g02001(.A0(new_n3001_), .A1(\A[504] ), .B0(new_n3003_), .Y(new_n3004_));
  NOR2   g02002(.A(new_n2990_), .B(new_n2992_), .Y(new_n3005_));
  AOI21  g02003(.A0(new_n2994_), .A1(\A[501] ), .B0(new_n3005_), .Y(new_n3006_));
  XOR2   g02004(.A(new_n3002_), .B(new_n2995_), .Y(new_n3007_));
  XOR2   g02005(.A(new_n3007_), .B(new_n2988_), .Y(new_n3008_));
  INV    g02006(.A(\A[495] ), .Y(new_n3009_));
  INV    g02007(.A(\A[494] ), .Y(new_n3010_));
  NAND2  g02008(.A(new_n3010_), .B(\A[493] ), .Y(new_n3011_));
  INV    g02009(.A(\A[493] ), .Y(new_n3012_));
  AOI21  g02010(.A0(\A[494] ), .A1(new_n3012_), .B0(new_n3009_), .Y(new_n3013_));
  XOR2   g02011(.A(\A[494] ), .B(\A[493] ), .Y(new_n3014_));
  AOI22  g02012(.A0(new_n3014_), .A1(new_n3009_), .B0(new_n3013_), .B1(new_n3011_), .Y(new_n3015_));
  INV    g02013(.A(\A[498] ), .Y(new_n3016_));
  INV    g02014(.A(\A[497] ), .Y(new_n3017_));
  NAND2  g02015(.A(new_n3017_), .B(\A[496] ), .Y(new_n3018_));
  INV    g02016(.A(\A[496] ), .Y(new_n3019_));
  AOI21  g02017(.A0(\A[497] ), .A1(new_n3019_), .B0(new_n3016_), .Y(new_n3020_));
  XOR2   g02018(.A(\A[497] ), .B(\A[496] ), .Y(new_n3021_));
  AOI22  g02019(.A0(new_n3021_), .A1(new_n3016_), .B0(new_n3020_), .B1(new_n3018_), .Y(new_n3022_));
  NOR2   g02020(.A(new_n3017_), .B(new_n3019_), .Y(new_n3023_));
  AOI21  g02021(.A0(new_n3021_), .A1(\A[498] ), .B0(new_n3023_), .Y(new_n3024_));
  NOR2   g02022(.A(new_n3010_), .B(new_n3012_), .Y(new_n3025_));
  AOI21  g02023(.A0(new_n3014_), .A1(\A[495] ), .B0(new_n3025_), .Y(new_n3026_));
  XOR2   g02024(.A(new_n3022_), .B(new_n3015_), .Y(new_n3027_));
  INV    g02025(.A(\A[489] ), .Y(new_n3028_));
  INV    g02026(.A(\A[488] ), .Y(new_n3029_));
  NAND2  g02027(.A(new_n3029_), .B(\A[487] ), .Y(new_n3030_));
  INV    g02028(.A(\A[487] ), .Y(new_n3031_));
  AOI21  g02029(.A0(\A[488] ), .A1(new_n3031_), .B0(new_n3028_), .Y(new_n3032_));
  XOR2   g02030(.A(\A[488] ), .B(\A[487] ), .Y(new_n3033_));
  AOI22  g02031(.A0(new_n3033_), .A1(new_n3028_), .B0(new_n3032_), .B1(new_n3030_), .Y(new_n3034_));
  INV    g02032(.A(\A[492] ), .Y(new_n3035_));
  INV    g02033(.A(\A[491] ), .Y(new_n3036_));
  NAND2  g02034(.A(new_n3036_), .B(\A[490] ), .Y(new_n3037_));
  INV    g02035(.A(\A[490] ), .Y(new_n3038_));
  AOI21  g02036(.A0(\A[491] ), .A1(new_n3038_), .B0(new_n3035_), .Y(new_n3039_));
  XOR2   g02037(.A(\A[491] ), .B(\A[490] ), .Y(new_n3040_));
  AOI22  g02038(.A0(new_n3040_), .A1(new_n3035_), .B0(new_n3039_), .B1(new_n3037_), .Y(new_n3041_));
  NOR2   g02039(.A(new_n3036_), .B(new_n3038_), .Y(new_n3042_));
  AOI21  g02040(.A0(new_n3040_), .A1(\A[492] ), .B0(new_n3042_), .Y(new_n3043_));
  NOR2   g02041(.A(new_n3029_), .B(new_n3031_), .Y(new_n3044_));
  AOI21  g02042(.A0(new_n3033_), .A1(\A[489] ), .B0(new_n3044_), .Y(new_n3045_));
  XOR2   g02043(.A(new_n3041_), .B(new_n3034_), .Y(new_n3046_));
  XOR2   g02044(.A(new_n3046_), .B(new_n3027_), .Y(new_n3047_));
  INV    g02045(.A(new_n3047_), .Y(new_n3048_));
  XOR2   g02046(.A(new_n3048_), .B(new_n3008_), .Y(new_n3049_));
  XOR2   g02047(.A(new_n3049_), .B(new_n2969_), .Y(new_n3050_));
  INV    g02048(.A(new_n3050_), .Y(new_n3051_));
  INV    g02049(.A(\A[555] ), .Y(new_n3052_));
  INV    g02050(.A(\A[554] ), .Y(new_n3053_));
  NAND2  g02051(.A(new_n3053_), .B(\A[553] ), .Y(new_n3054_));
  INV    g02052(.A(\A[553] ), .Y(new_n3055_));
  AOI21  g02053(.A0(\A[554] ), .A1(new_n3055_), .B0(new_n3052_), .Y(new_n3056_));
  XOR2   g02054(.A(\A[554] ), .B(\A[553] ), .Y(new_n3057_));
  AOI22  g02055(.A0(new_n3057_), .A1(new_n3052_), .B0(new_n3056_), .B1(new_n3054_), .Y(new_n3058_));
  INV    g02056(.A(\A[558] ), .Y(new_n3059_));
  INV    g02057(.A(\A[557] ), .Y(new_n3060_));
  NAND2  g02058(.A(new_n3060_), .B(\A[556] ), .Y(new_n3061_));
  INV    g02059(.A(\A[556] ), .Y(new_n3062_));
  AOI21  g02060(.A0(\A[557] ), .A1(new_n3062_), .B0(new_n3059_), .Y(new_n3063_));
  XOR2   g02061(.A(\A[557] ), .B(\A[556] ), .Y(new_n3064_));
  AOI22  g02062(.A0(new_n3064_), .A1(new_n3059_), .B0(new_n3063_), .B1(new_n3061_), .Y(new_n3065_));
  NOR2   g02063(.A(new_n3060_), .B(new_n3062_), .Y(new_n3066_));
  AOI21  g02064(.A0(new_n3064_), .A1(\A[558] ), .B0(new_n3066_), .Y(new_n3067_));
  NOR2   g02065(.A(new_n3053_), .B(new_n3055_), .Y(new_n3068_));
  AOI21  g02066(.A0(new_n3057_), .A1(\A[555] ), .B0(new_n3068_), .Y(new_n3069_));
  XOR2   g02067(.A(new_n3065_), .B(new_n3058_), .Y(new_n3070_));
  INV    g02068(.A(\A[549] ), .Y(new_n3071_));
  INV    g02069(.A(\A[548] ), .Y(new_n3072_));
  NAND2  g02070(.A(new_n3072_), .B(\A[547] ), .Y(new_n3073_));
  INV    g02071(.A(\A[547] ), .Y(new_n3074_));
  AOI21  g02072(.A0(\A[548] ), .A1(new_n3074_), .B0(new_n3071_), .Y(new_n3075_));
  XOR2   g02073(.A(\A[548] ), .B(\A[547] ), .Y(new_n3076_));
  AOI22  g02074(.A0(new_n3076_), .A1(new_n3071_), .B0(new_n3075_), .B1(new_n3073_), .Y(new_n3077_));
  INV    g02075(.A(\A[552] ), .Y(new_n3078_));
  INV    g02076(.A(\A[551] ), .Y(new_n3079_));
  NAND2  g02077(.A(new_n3079_), .B(\A[550] ), .Y(new_n3080_));
  INV    g02078(.A(\A[550] ), .Y(new_n3081_));
  AOI21  g02079(.A0(\A[551] ), .A1(new_n3081_), .B0(new_n3078_), .Y(new_n3082_));
  XOR2   g02080(.A(\A[551] ), .B(\A[550] ), .Y(new_n3083_));
  AOI22  g02081(.A0(new_n3083_), .A1(new_n3078_), .B0(new_n3082_), .B1(new_n3080_), .Y(new_n3084_));
  NAND2  g02082(.A(\A[551] ), .B(\A[550] ), .Y(new_n3085_));
  INV    g02083(.A(new_n3085_), .Y(new_n3086_));
  AOI21  g02084(.A0(new_n3083_), .A1(\A[552] ), .B0(new_n3086_), .Y(new_n3087_));
  NOR2   g02085(.A(new_n3072_), .B(new_n3074_), .Y(new_n3088_));
  AOI21  g02086(.A0(new_n3076_), .A1(\A[549] ), .B0(new_n3088_), .Y(new_n3089_));
  XOR2   g02087(.A(new_n3084_), .B(new_n3077_), .Y(new_n3090_));
  XOR2   g02088(.A(new_n3090_), .B(new_n3070_), .Y(new_n3091_));
  INV    g02089(.A(\A[543] ), .Y(new_n3092_));
  INV    g02090(.A(\A[542] ), .Y(new_n3093_));
  NAND2  g02091(.A(new_n3093_), .B(\A[541] ), .Y(new_n3094_));
  INV    g02092(.A(\A[541] ), .Y(new_n3095_));
  AOI21  g02093(.A0(\A[542] ), .A1(new_n3095_), .B0(new_n3092_), .Y(new_n3096_));
  XOR2   g02094(.A(\A[542] ), .B(\A[541] ), .Y(new_n3097_));
  AOI22  g02095(.A0(new_n3097_), .A1(new_n3092_), .B0(new_n3096_), .B1(new_n3094_), .Y(new_n3098_));
  INV    g02096(.A(\A[546] ), .Y(new_n3099_));
  INV    g02097(.A(\A[545] ), .Y(new_n3100_));
  NAND2  g02098(.A(new_n3100_), .B(\A[544] ), .Y(new_n3101_));
  INV    g02099(.A(\A[544] ), .Y(new_n3102_));
  AOI21  g02100(.A0(\A[545] ), .A1(new_n3102_), .B0(new_n3099_), .Y(new_n3103_));
  XOR2   g02101(.A(\A[545] ), .B(\A[544] ), .Y(new_n3104_));
  AOI22  g02102(.A0(new_n3104_), .A1(new_n3099_), .B0(new_n3103_), .B1(new_n3101_), .Y(new_n3105_));
  NOR2   g02103(.A(new_n3100_), .B(new_n3102_), .Y(new_n3106_));
  AOI21  g02104(.A0(new_n3104_), .A1(\A[546] ), .B0(new_n3106_), .Y(new_n3107_));
  NOR2   g02105(.A(new_n3093_), .B(new_n3095_), .Y(new_n3108_));
  AOI21  g02106(.A0(new_n3097_), .A1(\A[543] ), .B0(new_n3108_), .Y(new_n3109_));
  XOR2   g02107(.A(new_n3105_), .B(new_n3098_), .Y(new_n3110_));
  INV    g02108(.A(\A[537] ), .Y(new_n3111_));
  INV    g02109(.A(\A[536] ), .Y(new_n3112_));
  NAND2  g02110(.A(new_n3112_), .B(\A[535] ), .Y(new_n3113_));
  INV    g02111(.A(\A[535] ), .Y(new_n3114_));
  AOI21  g02112(.A0(\A[536] ), .A1(new_n3114_), .B0(new_n3111_), .Y(new_n3115_));
  XOR2   g02113(.A(\A[536] ), .B(\A[535] ), .Y(new_n3116_));
  AOI22  g02114(.A0(new_n3116_), .A1(new_n3111_), .B0(new_n3115_), .B1(new_n3113_), .Y(new_n3117_));
  INV    g02115(.A(\A[540] ), .Y(new_n3118_));
  INV    g02116(.A(\A[539] ), .Y(new_n3119_));
  NAND2  g02117(.A(new_n3119_), .B(\A[538] ), .Y(new_n3120_));
  INV    g02118(.A(\A[538] ), .Y(new_n3121_));
  AOI21  g02119(.A0(\A[539] ), .A1(new_n3121_), .B0(new_n3118_), .Y(new_n3122_));
  XOR2   g02120(.A(\A[539] ), .B(\A[538] ), .Y(new_n3123_));
  AOI22  g02121(.A0(new_n3123_), .A1(new_n3118_), .B0(new_n3122_), .B1(new_n3120_), .Y(new_n3124_));
  NOR2   g02122(.A(new_n3119_), .B(new_n3121_), .Y(new_n3125_));
  AOI21  g02123(.A0(new_n3123_), .A1(\A[540] ), .B0(new_n3125_), .Y(new_n3126_));
  NOR2   g02124(.A(new_n3112_), .B(new_n3114_), .Y(new_n3127_));
  AOI21  g02125(.A0(new_n3116_), .A1(\A[537] ), .B0(new_n3127_), .Y(new_n3128_));
  XOR2   g02126(.A(new_n3124_), .B(new_n3117_), .Y(new_n3129_));
  XOR2   g02127(.A(new_n3129_), .B(new_n3110_), .Y(new_n3130_));
  INV    g02128(.A(new_n3130_), .Y(new_n3131_));
  XOR2   g02129(.A(new_n3131_), .B(new_n3091_), .Y(new_n3132_));
  INV    g02130(.A(new_n3132_), .Y(new_n3133_));
  INV    g02131(.A(\A[531] ), .Y(new_n3134_));
  INV    g02132(.A(\A[530] ), .Y(new_n3135_));
  NAND2  g02133(.A(new_n3135_), .B(\A[529] ), .Y(new_n3136_));
  INV    g02134(.A(\A[529] ), .Y(new_n3137_));
  AOI21  g02135(.A0(\A[530] ), .A1(new_n3137_), .B0(new_n3134_), .Y(new_n3138_));
  XOR2   g02136(.A(\A[530] ), .B(\A[529] ), .Y(new_n3139_));
  AOI22  g02137(.A0(new_n3139_), .A1(new_n3134_), .B0(new_n3138_), .B1(new_n3136_), .Y(new_n3140_));
  INV    g02138(.A(\A[534] ), .Y(new_n3141_));
  INV    g02139(.A(\A[533] ), .Y(new_n3142_));
  NAND2  g02140(.A(new_n3142_), .B(\A[532] ), .Y(new_n3143_));
  INV    g02141(.A(\A[532] ), .Y(new_n3144_));
  AOI21  g02142(.A0(\A[533] ), .A1(new_n3144_), .B0(new_n3141_), .Y(new_n3145_));
  XOR2   g02143(.A(\A[533] ), .B(\A[532] ), .Y(new_n3146_));
  AOI22  g02144(.A0(new_n3146_), .A1(new_n3141_), .B0(new_n3145_), .B1(new_n3143_), .Y(new_n3147_));
  NOR2   g02145(.A(new_n3142_), .B(new_n3144_), .Y(new_n3148_));
  AOI21  g02146(.A0(new_n3146_), .A1(\A[534] ), .B0(new_n3148_), .Y(new_n3149_));
  NOR2   g02147(.A(new_n3135_), .B(new_n3137_), .Y(new_n3150_));
  AOI21  g02148(.A0(new_n3139_), .A1(\A[531] ), .B0(new_n3150_), .Y(new_n3151_));
  XOR2   g02149(.A(new_n3147_), .B(new_n3140_), .Y(new_n3152_));
  INV    g02150(.A(\A[525] ), .Y(new_n3153_));
  INV    g02151(.A(\A[524] ), .Y(new_n3154_));
  NAND2  g02152(.A(new_n3154_), .B(\A[523] ), .Y(new_n3155_));
  INV    g02153(.A(\A[523] ), .Y(new_n3156_));
  AOI21  g02154(.A0(\A[524] ), .A1(new_n3156_), .B0(new_n3153_), .Y(new_n3157_));
  XOR2   g02155(.A(\A[524] ), .B(\A[523] ), .Y(new_n3158_));
  AOI22  g02156(.A0(new_n3158_), .A1(new_n3153_), .B0(new_n3157_), .B1(new_n3155_), .Y(new_n3159_));
  INV    g02157(.A(\A[528] ), .Y(new_n3160_));
  INV    g02158(.A(\A[527] ), .Y(new_n3161_));
  NAND2  g02159(.A(new_n3161_), .B(\A[526] ), .Y(new_n3162_));
  INV    g02160(.A(\A[526] ), .Y(new_n3163_));
  AOI21  g02161(.A0(\A[527] ), .A1(new_n3163_), .B0(new_n3160_), .Y(new_n3164_));
  XOR2   g02162(.A(\A[527] ), .B(\A[526] ), .Y(new_n3165_));
  AOI22  g02163(.A0(new_n3165_), .A1(new_n3160_), .B0(new_n3164_), .B1(new_n3162_), .Y(new_n3166_));
  NOR2   g02164(.A(new_n3161_), .B(new_n3163_), .Y(new_n3167_));
  AOI21  g02165(.A0(new_n3165_), .A1(\A[528] ), .B0(new_n3167_), .Y(new_n3168_));
  NOR2   g02166(.A(new_n3154_), .B(new_n3156_), .Y(new_n3169_));
  AOI21  g02167(.A0(new_n3158_), .A1(\A[525] ), .B0(new_n3169_), .Y(new_n3170_));
  XOR2   g02168(.A(new_n3166_), .B(new_n3159_), .Y(new_n3171_));
  XOR2   g02169(.A(new_n3171_), .B(new_n3152_), .Y(new_n3172_));
  INV    g02170(.A(\A[519] ), .Y(new_n3173_));
  INV    g02171(.A(\A[518] ), .Y(new_n3174_));
  NAND2  g02172(.A(new_n3174_), .B(\A[517] ), .Y(new_n3175_));
  INV    g02173(.A(\A[517] ), .Y(new_n3176_));
  AOI21  g02174(.A0(\A[518] ), .A1(new_n3176_), .B0(new_n3173_), .Y(new_n3177_));
  XOR2   g02175(.A(\A[518] ), .B(\A[517] ), .Y(new_n3178_));
  AOI22  g02176(.A0(new_n3178_), .A1(new_n3173_), .B0(new_n3177_), .B1(new_n3175_), .Y(new_n3179_));
  INV    g02177(.A(\A[522] ), .Y(new_n3180_));
  INV    g02178(.A(\A[521] ), .Y(new_n3181_));
  NAND2  g02179(.A(new_n3181_), .B(\A[520] ), .Y(new_n3182_));
  INV    g02180(.A(\A[520] ), .Y(new_n3183_));
  AOI21  g02181(.A0(\A[521] ), .A1(new_n3183_), .B0(new_n3180_), .Y(new_n3184_));
  XOR2   g02182(.A(\A[521] ), .B(\A[520] ), .Y(new_n3185_));
  AOI22  g02183(.A0(new_n3185_), .A1(new_n3180_), .B0(new_n3184_), .B1(new_n3182_), .Y(new_n3186_));
  NOR2   g02184(.A(new_n3181_), .B(new_n3183_), .Y(new_n3187_));
  AOI21  g02185(.A0(new_n3185_), .A1(\A[522] ), .B0(new_n3187_), .Y(new_n3188_));
  NOR2   g02186(.A(new_n3174_), .B(new_n3176_), .Y(new_n3189_));
  AOI21  g02187(.A0(new_n3178_), .A1(\A[519] ), .B0(new_n3189_), .Y(new_n3190_));
  XOR2   g02188(.A(new_n3186_), .B(new_n3179_), .Y(new_n3191_));
  INV    g02189(.A(\A[513] ), .Y(new_n3192_));
  INV    g02190(.A(\A[512] ), .Y(new_n3193_));
  NAND2  g02191(.A(new_n3193_), .B(\A[511] ), .Y(new_n3194_));
  INV    g02192(.A(\A[511] ), .Y(new_n3195_));
  AOI21  g02193(.A0(\A[512] ), .A1(new_n3195_), .B0(new_n3192_), .Y(new_n3196_));
  XOR2   g02194(.A(\A[512] ), .B(\A[511] ), .Y(new_n3197_));
  AOI22  g02195(.A0(new_n3197_), .A1(new_n3192_), .B0(new_n3196_), .B1(new_n3194_), .Y(new_n3198_));
  INV    g02196(.A(\A[516] ), .Y(new_n3199_));
  INV    g02197(.A(\A[515] ), .Y(new_n3200_));
  NAND2  g02198(.A(new_n3200_), .B(\A[514] ), .Y(new_n3201_));
  INV    g02199(.A(\A[514] ), .Y(new_n3202_));
  AOI21  g02200(.A0(\A[515] ), .A1(new_n3202_), .B0(new_n3199_), .Y(new_n3203_));
  XOR2   g02201(.A(\A[515] ), .B(\A[514] ), .Y(new_n3204_));
  AOI22  g02202(.A0(new_n3204_), .A1(new_n3199_), .B0(new_n3203_), .B1(new_n3201_), .Y(new_n3205_));
  NOR2   g02203(.A(new_n3200_), .B(new_n3202_), .Y(new_n3206_));
  AOI21  g02204(.A0(new_n3204_), .A1(\A[516] ), .B0(new_n3206_), .Y(new_n3207_));
  NOR2   g02205(.A(new_n3193_), .B(new_n3195_), .Y(new_n3208_));
  AOI21  g02206(.A0(new_n3197_), .A1(\A[513] ), .B0(new_n3208_), .Y(new_n3209_));
  XOR2   g02207(.A(new_n3205_), .B(new_n3198_), .Y(new_n3210_));
  XOR2   g02208(.A(new_n3210_), .B(new_n3191_), .Y(new_n3211_));
  INV    g02209(.A(new_n3211_), .Y(new_n3212_));
  XOR2   g02210(.A(new_n3212_), .B(new_n3172_), .Y(new_n3213_));
  XOR2   g02211(.A(new_n3213_), .B(new_n3133_), .Y(new_n3214_));
  XOR2   g02212(.A(new_n3214_), .B(new_n3051_), .Y(new_n3215_));
  INV    g02213(.A(new_n3215_), .Y(new_n3216_));
  INV    g02214(.A(\A[651] ), .Y(new_n3217_));
  INV    g02215(.A(\A[650] ), .Y(new_n3218_));
  NAND2  g02216(.A(new_n3218_), .B(\A[649] ), .Y(new_n3219_));
  INV    g02217(.A(\A[649] ), .Y(new_n3220_));
  AOI21  g02218(.A0(\A[650] ), .A1(new_n3220_), .B0(new_n3217_), .Y(new_n3221_));
  XOR2   g02219(.A(\A[650] ), .B(\A[649] ), .Y(new_n3222_));
  AOI22  g02220(.A0(new_n3222_), .A1(new_n3217_), .B0(new_n3221_), .B1(new_n3219_), .Y(new_n3223_));
  INV    g02221(.A(\A[654] ), .Y(new_n3224_));
  INV    g02222(.A(\A[653] ), .Y(new_n3225_));
  NAND2  g02223(.A(new_n3225_), .B(\A[652] ), .Y(new_n3226_));
  INV    g02224(.A(\A[652] ), .Y(new_n3227_));
  AOI21  g02225(.A0(\A[653] ), .A1(new_n3227_), .B0(new_n3224_), .Y(new_n3228_));
  XOR2   g02226(.A(\A[653] ), .B(\A[652] ), .Y(new_n3229_));
  AOI22  g02227(.A0(new_n3229_), .A1(new_n3224_), .B0(new_n3228_), .B1(new_n3226_), .Y(new_n3230_));
  NOR2   g02228(.A(new_n3225_), .B(new_n3227_), .Y(new_n3231_));
  AOI21  g02229(.A0(new_n3229_), .A1(\A[654] ), .B0(new_n3231_), .Y(new_n3232_));
  NOR2   g02230(.A(new_n3218_), .B(new_n3220_), .Y(new_n3233_));
  AOI21  g02231(.A0(new_n3222_), .A1(\A[651] ), .B0(new_n3233_), .Y(new_n3234_));
  XOR2   g02232(.A(new_n3230_), .B(new_n3223_), .Y(new_n3235_));
  INV    g02233(.A(\A[645] ), .Y(new_n3236_));
  INV    g02234(.A(\A[644] ), .Y(new_n3237_));
  NAND2  g02235(.A(new_n3237_), .B(\A[643] ), .Y(new_n3238_));
  INV    g02236(.A(\A[643] ), .Y(new_n3239_));
  AOI21  g02237(.A0(\A[644] ), .A1(new_n3239_), .B0(new_n3236_), .Y(new_n3240_));
  XOR2   g02238(.A(\A[644] ), .B(\A[643] ), .Y(new_n3241_));
  AOI22  g02239(.A0(new_n3241_), .A1(new_n3236_), .B0(new_n3240_), .B1(new_n3238_), .Y(new_n3242_));
  INV    g02240(.A(\A[648] ), .Y(new_n3243_));
  INV    g02241(.A(\A[647] ), .Y(new_n3244_));
  NAND2  g02242(.A(new_n3244_), .B(\A[646] ), .Y(new_n3245_));
  INV    g02243(.A(\A[646] ), .Y(new_n3246_));
  AOI21  g02244(.A0(\A[647] ), .A1(new_n3246_), .B0(new_n3243_), .Y(new_n3247_));
  XOR2   g02245(.A(\A[647] ), .B(\A[646] ), .Y(new_n3248_));
  AOI22  g02246(.A0(new_n3248_), .A1(new_n3243_), .B0(new_n3247_), .B1(new_n3245_), .Y(new_n3249_));
  NAND2  g02247(.A(\A[647] ), .B(\A[646] ), .Y(new_n3250_));
  INV    g02248(.A(new_n3250_), .Y(new_n3251_));
  AOI21  g02249(.A0(new_n3248_), .A1(\A[648] ), .B0(new_n3251_), .Y(new_n3252_));
  NOR2   g02250(.A(new_n3237_), .B(new_n3239_), .Y(new_n3253_));
  AOI21  g02251(.A0(new_n3241_), .A1(\A[645] ), .B0(new_n3253_), .Y(new_n3254_));
  XOR2   g02252(.A(new_n3249_), .B(new_n3242_), .Y(new_n3255_));
  XOR2   g02253(.A(new_n3255_), .B(new_n3235_), .Y(new_n3256_));
  INV    g02254(.A(\A[639] ), .Y(new_n3257_));
  INV    g02255(.A(\A[638] ), .Y(new_n3258_));
  NAND2  g02256(.A(new_n3258_), .B(\A[637] ), .Y(new_n3259_));
  INV    g02257(.A(\A[637] ), .Y(new_n3260_));
  AOI21  g02258(.A0(\A[638] ), .A1(new_n3260_), .B0(new_n3257_), .Y(new_n3261_));
  XOR2   g02259(.A(\A[638] ), .B(\A[637] ), .Y(new_n3262_));
  AOI22  g02260(.A0(new_n3262_), .A1(new_n3257_), .B0(new_n3261_), .B1(new_n3259_), .Y(new_n3263_));
  INV    g02261(.A(\A[642] ), .Y(new_n3264_));
  INV    g02262(.A(\A[641] ), .Y(new_n3265_));
  NAND2  g02263(.A(new_n3265_), .B(\A[640] ), .Y(new_n3266_));
  INV    g02264(.A(\A[640] ), .Y(new_n3267_));
  AOI21  g02265(.A0(\A[641] ), .A1(new_n3267_), .B0(new_n3264_), .Y(new_n3268_));
  XOR2   g02266(.A(\A[641] ), .B(\A[640] ), .Y(new_n3269_));
  AOI22  g02267(.A0(new_n3269_), .A1(new_n3264_), .B0(new_n3268_), .B1(new_n3266_), .Y(new_n3270_));
  NOR2   g02268(.A(new_n3265_), .B(new_n3267_), .Y(new_n3271_));
  AOI21  g02269(.A0(new_n3269_), .A1(\A[642] ), .B0(new_n3271_), .Y(new_n3272_));
  NOR2   g02270(.A(new_n3258_), .B(new_n3260_), .Y(new_n3273_));
  AOI21  g02271(.A0(new_n3262_), .A1(\A[639] ), .B0(new_n3273_), .Y(new_n3274_));
  XOR2   g02272(.A(new_n3270_), .B(new_n3263_), .Y(new_n3275_));
  INV    g02273(.A(\A[633] ), .Y(new_n3276_));
  INV    g02274(.A(\A[632] ), .Y(new_n3277_));
  NAND2  g02275(.A(new_n3277_), .B(\A[631] ), .Y(new_n3278_));
  INV    g02276(.A(\A[631] ), .Y(new_n3279_));
  AOI21  g02277(.A0(\A[632] ), .A1(new_n3279_), .B0(new_n3276_), .Y(new_n3280_));
  XOR2   g02278(.A(\A[632] ), .B(\A[631] ), .Y(new_n3281_));
  AOI22  g02279(.A0(new_n3281_), .A1(new_n3276_), .B0(new_n3280_), .B1(new_n3278_), .Y(new_n3282_));
  INV    g02280(.A(\A[636] ), .Y(new_n3283_));
  INV    g02281(.A(\A[635] ), .Y(new_n3284_));
  NAND2  g02282(.A(new_n3284_), .B(\A[634] ), .Y(new_n3285_));
  INV    g02283(.A(\A[634] ), .Y(new_n3286_));
  AOI21  g02284(.A0(\A[635] ), .A1(new_n3286_), .B0(new_n3283_), .Y(new_n3287_));
  XOR2   g02285(.A(\A[635] ), .B(\A[634] ), .Y(new_n3288_));
  AOI22  g02286(.A0(new_n3288_), .A1(new_n3283_), .B0(new_n3287_), .B1(new_n3285_), .Y(new_n3289_));
  NOR2   g02287(.A(new_n3284_), .B(new_n3286_), .Y(new_n3290_));
  AOI21  g02288(.A0(new_n3288_), .A1(\A[636] ), .B0(new_n3290_), .Y(new_n3291_));
  NOR2   g02289(.A(new_n3277_), .B(new_n3279_), .Y(new_n3292_));
  AOI21  g02290(.A0(new_n3281_), .A1(\A[633] ), .B0(new_n3292_), .Y(new_n3293_));
  XOR2   g02291(.A(new_n3289_), .B(new_n3282_), .Y(new_n3294_));
  XOR2   g02292(.A(new_n3294_), .B(new_n3275_), .Y(new_n3295_));
  INV    g02293(.A(new_n3295_), .Y(new_n3296_));
  XOR2   g02294(.A(new_n3296_), .B(new_n3256_), .Y(new_n3297_));
  INV    g02295(.A(new_n3297_), .Y(new_n3298_));
  INV    g02296(.A(\A[627] ), .Y(new_n3299_));
  INV    g02297(.A(\A[626] ), .Y(new_n3300_));
  NAND2  g02298(.A(new_n3300_), .B(\A[625] ), .Y(new_n3301_));
  INV    g02299(.A(\A[625] ), .Y(new_n3302_));
  AOI21  g02300(.A0(\A[626] ), .A1(new_n3302_), .B0(new_n3299_), .Y(new_n3303_));
  XOR2   g02301(.A(\A[626] ), .B(\A[625] ), .Y(new_n3304_));
  AOI22  g02302(.A0(new_n3304_), .A1(new_n3299_), .B0(new_n3303_), .B1(new_n3301_), .Y(new_n3305_));
  INV    g02303(.A(\A[630] ), .Y(new_n3306_));
  INV    g02304(.A(\A[629] ), .Y(new_n3307_));
  NAND2  g02305(.A(new_n3307_), .B(\A[628] ), .Y(new_n3308_));
  INV    g02306(.A(\A[628] ), .Y(new_n3309_));
  AOI21  g02307(.A0(\A[629] ), .A1(new_n3309_), .B0(new_n3306_), .Y(new_n3310_));
  XOR2   g02308(.A(\A[629] ), .B(\A[628] ), .Y(new_n3311_));
  AOI22  g02309(.A0(new_n3311_), .A1(new_n3306_), .B0(new_n3310_), .B1(new_n3308_), .Y(new_n3312_));
  NOR2   g02310(.A(new_n3307_), .B(new_n3309_), .Y(new_n3313_));
  AOI21  g02311(.A0(new_n3311_), .A1(\A[630] ), .B0(new_n3313_), .Y(new_n3314_));
  NOR2   g02312(.A(new_n3300_), .B(new_n3302_), .Y(new_n3315_));
  AOI21  g02313(.A0(new_n3304_), .A1(\A[627] ), .B0(new_n3315_), .Y(new_n3316_));
  XOR2   g02314(.A(new_n3312_), .B(new_n3305_), .Y(new_n3317_));
  INV    g02315(.A(\A[621] ), .Y(new_n3318_));
  INV    g02316(.A(\A[620] ), .Y(new_n3319_));
  NAND2  g02317(.A(new_n3319_), .B(\A[619] ), .Y(new_n3320_));
  INV    g02318(.A(\A[619] ), .Y(new_n3321_));
  AOI21  g02319(.A0(\A[620] ), .A1(new_n3321_), .B0(new_n3318_), .Y(new_n3322_));
  XOR2   g02320(.A(\A[620] ), .B(\A[619] ), .Y(new_n3323_));
  AOI22  g02321(.A0(new_n3323_), .A1(new_n3318_), .B0(new_n3322_), .B1(new_n3320_), .Y(new_n3324_));
  INV    g02322(.A(\A[624] ), .Y(new_n3325_));
  INV    g02323(.A(\A[623] ), .Y(new_n3326_));
  NAND2  g02324(.A(new_n3326_), .B(\A[622] ), .Y(new_n3327_));
  INV    g02325(.A(\A[622] ), .Y(new_n3328_));
  AOI21  g02326(.A0(\A[623] ), .A1(new_n3328_), .B0(new_n3325_), .Y(new_n3329_));
  XOR2   g02327(.A(\A[623] ), .B(\A[622] ), .Y(new_n3330_));
  AOI22  g02328(.A0(new_n3330_), .A1(new_n3325_), .B0(new_n3329_), .B1(new_n3327_), .Y(new_n3331_));
  NOR2   g02329(.A(new_n3326_), .B(new_n3328_), .Y(new_n3332_));
  AOI21  g02330(.A0(new_n3330_), .A1(\A[624] ), .B0(new_n3332_), .Y(new_n3333_));
  NOR2   g02331(.A(new_n3319_), .B(new_n3321_), .Y(new_n3334_));
  AOI21  g02332(.A0(new_n3323_), .A1(\A[621] ), .B0(new_n3334_), .Y(new_n3335_));
  XOR2   g02333(.A(new_n3331_), .B(new_n3324_), .Y(new_n3336_));
  XOR2   g02334(.A(new_n3336_), .B(new_n3317_), .Y(new_n3337_));
  INV    g02335(.A(\A[615] ), .Y(new_n3338_));
  INV    g02336(.A(\A[614] ), .Y(new_n3339_));
  NAND2  g02337(.A(new_n3339_), .B(\A[613] ), .Y(new_n3340_));
  INV    g02338(.A(\A[613] ), .Y(new_n3341_));
  AOI21  g02339(.A0(\A[614] ), .A1(new_n3341_), .B0(new_n3338_), .Y(new_n3342_));
  XOR2   g02340(.A(\A[614] ), .B(\A[613] ), .Y(new_n3343_));
  AOI22  g02341(.A0(new_n3343_), .A1(new_n3338_), .B0(new_n3342_), .B1(new_n3340_), .Y(new_n3344_));
  INV    g02342(.A(\A[618] ), .Y(new_n3345_));
  INV    g02343(.A(\A[617] ), .Y(new_n3346_));
  NAND2  g02344(.A(new_n3346_), .B(\A[616] ), .Y(new_n3347_));
  INV    g02345(.A(\A[616] ), .Y(new_n3348_));
  AOI21  g02346(.A0(\A[617] ), .A1(new_n3348_), .B0(new_n3345_), .Y(new_n3349_));
  XOR2   g02347(.A(\A[617] ), .B(\A[616] ), .Y(new_n3350_));
  AOI22  g02348(.A0(new_n3350_), .A1(new_n3345_), .B0(new_n3349_), .B1(new_n3347_), .Y(new_n3351_));
  NOR2   g02349(.A(new_n3346_), .B(new_n3348_), .Y(new_n3352_));
  AOI21  g02350(.A0(new_n3350_), .A1(\A[618] ), .B0(new_n3352_), .Y(new_n3353_));
  NOR2   g02351(.A(new_n3339_), .B(new_n3341_), .Y(new_n3354_));
  AOI21  g02352(.A0(new_n3343_), .A1(\A[615] ), .B0(new_n3354_), .Y(new_n3355_));
  XOR2   g02353(.A(new_n3351_), .B(new_n3344_), .Y(new_n3356_));
  INV    g02354(.A(\A[609] ), .Y(new_n3357_));
  INV    g02355(.A(\A[608] ), .Y(new_n3358_));
  NAND2  g02356(.A(new_n3358_), .B(\A[607] ), .Y(new_n3359_));
  INV    g02357(.A(\A[607] ), .Y(new_n3360_));
  AOI21  g02358(.A0(\A[608] ), .A1(new_n3360_), .B0(new_n3357_), .Y(new_n3361_));
  XOR2   g02359(.A(\A[608] ), .B(\A[607] ), .Y(new_n3362_));
  AOI22  g02360(.A0(new_n3362_), .A1(new_n3357_), .B0(new_n3361_), .B1(new_n3359_), .Y(new_n3363_));
  INV    g02361(.A(\A[612] ), .Y(new_n3364_));
  INV    g02362(.A(\A[611] ), .Y(new_n3365_));
  NAND2  g02363(.A(new_n3365_), .B(\A[610] ), .Y(new_n3366_));
  INV    g02364(.A(\A[610] ), .Y(new_n3367_));
  AOI21  g02365(.A0(\A[611] ), .A1(new_n3367_), .B0(new_n3364_), .Y(new_n3368_));
  XOR2   g02366(.A(\A[611] ), .B(\A[610] ), .Y(new_n3369_));
  AOI22  g02367(.A0(new_n3369_), .A1(new_n3364_), .B0(new_n3368_), .B1(new_n3366_), .Y(new_n3370_));
  NOR2   g02368(.A(new_n3365_), .B(new_n3367_), .Y(new_n3371_));
  AOI21  g02369(.A0(new_n3369_), .A1(\A[612] ), .B0(new_n3371_), .Y(new_n3372_));
  NOR2   g02370(.A(new_n3358_), .B(new_n3360_), .Y(new_n3373_));
  AOI21  g02371(.A0(new_n3362_), .A1(\A[609] ), .B0(new_n3373_), .Y(new_n3374_));
  XOR2   g02372(.A(new_n3370_), .B(new_n3363_), .Y(new_n3375_));
  XOR2   g02373(.A(new_n3375_), .B(new_n3356_), .Y(new_n3376_));
  INV    g02374(.A(new_n3376_), .Y(new_n3377_));
  XOR2   g02375(.A(new_n3377_), .B(new_n3337_), .Y(new_n3378_));
  XOR2   g02376(.A(new_n3378_), .B(new_n3298_), .Y(new_n3379_));
  INV    g02377(.A(new_n3379_), .Y(new_n3380_));
  INV    g02378(.A(\A[603] ), .Y(new_n3381_));
  INV    g02379(.A(\A[602] ), .Y(new_n3382_));
  NAND2  g02380(.A(new_n3382_), .B(\A[601] ), .Y(new_n3383_));
  INV    g02381(.A(\A[601] ), .Y(new_n3384_));
  AOI21  g02382(.A0(\A[602] ), .A1(new_n3384_), .B0(new_n3381_), .Y(new_n3385_));
  XOR2   g02383(.A(\A[602] ), .B(\A[601] ), .Y(new_n3386_));
  AOI22  g02384(.A0(new_n3386_), .A1(new_n3381_), .B0(new_n3385_), .B1(new_n3383_), .Y(new_n3387_));
  INV    g02385(.A(\A[606] ), .Y(new_n3388_));
  INV    g02386(.A(\A[605] ), .Y(new_n3389_));
  NAND2  g02387(.A(new_n3389_), .B(\A[604] ), .Y(new_n3390_));
  INV    g02388(.A(\A[604] ), .Y(new_n3391_));
  AOI21  g02389(.A0(\A[605] ), .A1(new_n3391_), .B0(new_n3388_), .Y(new_n3392_));
  XOR2   g02390(.A(\A[605] ), .B(\A[604] ), .Y(new_n3393_));
  AOI22  g02391(.A0(new_n3393_), .A1(new_n3388_), .B0(new_n3392_), .B1(new_n3390_), .Y(new_n3394_));
  NOR2   g02392(.A(new_n3389_), .B(new_n3391_), .Y(new_n3395_));
  AOI21  g02393(.A0(new_n3393_), .A1(\A[606] ), .B0(new_n3395_), .Y(new_n3396_));
  NOR2   g02394(.A(new_n3382_), .B(new_n3384_), .Y(new_n3397_));
  AOI21  g02395(.A0(new_n3386_), .A1(\A[603] ), .B0(new_n3397_), .Y(new_n3398_));
  XOR2   g02396(.A(new_n3394_), .B(new_n3387_), .Y(new_n3399_));
  INV    g02397(.A(\A[597] ), .Y(new_n3400_));
  INV    g02398(.A(\A[596] ), .Y(new_n3401_));
  NAND2  g02399(.A(new_n3401_), .B(\A[595] ), .Y(new_n3402_));
  INV    g02400(.A(\A[595] ), .Y(new_n3403_));
  AOI21  g02401(.A0(\A[596] ), .A1(new_n3403_), .B0(new_n3400_), .Y(new_n3404_));
  XOR2   g02402(.A(\A[596] ), .B(\A[595] ), .Y(new_n3405_));
  AOI22  g02403(.A0(new_n3405_), .A1(new_n3400_), .B0(new_n3404_), .B1(new_n3402_), .Y(new_n3406_));
  INV    g02404(.A(\A[600] ), .Y(new_n3407_));
  INV    g02405(.A(\A[599] ), .Y(new_n3408_));
  NAND2  g02406(.A(new_n3408_), .B(\A[598] ), .Y(new_n3409_));
  INV    g02407(.A(\A[598] ), .Y(new_n3410_));
  AOI21  g02408(.A0(\A[599] ), .A1(new_n3410_), .B0(new_n3407_), .Y(new_n3411_));
  XOR2   g02409(.A(\A[599] ), .B(\A[598] ), .Y(new_n3412_));
  AOI22  g02410(.A0(new_n3412_), .A1(new_n3407_), .B0(new_n3411_), .B1(new_n3409_), .Y(new_n3413_));
  NOR2   g02411(.A(new_n3408_), .B(new_n3410_), .Y(new_n3414_));
  AOI21  g02412(.A0(new_n3412_), .A1(\A[600] ), .B0(new_n3414_), .Y(new_n3415_));
  NOR2   g02413(.A(new_n3401_), .B(new_n3403_), .Y(new_n3416_));
  AOI21  g02414(.A0(new_n3405_), .A1(\A[597] ), .B0(new_n3416_), .Y(new_n3417_));
  XOR2   g02415(.A(new_n3413_), .B(new_n3406_), .Y(new_n3418_));
  XOR2   g02416(.A(new_n3418_), .B(new_n3399_), .Y(new_n3419_));
  INV    g02417(.A(\A[591] ), .Y(new_n3420_));
  INV    g02418(.A(\A[590] ), .Y(new_n3421_));
  NAND2  g02419(.A(new_n3421_), .B(\A[589] ), .Y(new_n3422_));
  INV    g02420(.A(\A[589] ), .Y(new_n3423_));
  AOI21  g02421(.A0(\A[590] ), .A1(new_n3423_), .B0(new_n3420_), .Y(new_n3424_));
  XOR2   g02422(.A(\A[590] ), .B(\A[589] ), .Y(new_n3425_));
  AOI22  g02423(.A0(new_n3425_), .A1(new_n3420_), .B0(new_n3424_), .B1(new_n3422_), .Y(new_n3426_));
  INV    g02424(.A(\A[594] ), .Y(new_n3427_));
  INV    g02425(.A(\A[593] ), .Y(new_n3428_));
  NAND2  g02426(.A(new_n3428_), .B(\A[592] ), .Y(new_n3429_));
  INV    g02427(.A(\A[592] ), .Y(new_n3430_));
  AOI21  g02428(.A0(\A[593] ), .A1(new_n3430_), .B0(new_n3427_), .Y(new_n3431_));
  XOR2   g02429(.A(\A[593] ), .B(\A[592] ), .Y(new_n3432_));
  AOI22  g02430(.A0(new_n3432_), .A1(new_n3427_), .B0(new_n3431_), .B1(new_n3429_), .Y(new_n3433_));
  NOR2   g02431(.A(new_n3428_), .B(new_n3430_), .Y(new_n3434_));
  AOI21  g02432(.A0(new_n3432_), .A1(\A[594] ), .B0(new_n3434_), .Y(new_n3435_));
  NOR2   g02433(.A(new_n3421_), .B(new_n3423_), .Y(new_n3436_));
  AOI21  g02434(.A0(new_n3425_), .A1(\A[591] ), .B0(new_n3436_), .Y(new_n3437_));
  XOR2   g02435(.A(new_n3433_), .B(new_n3426_), .Y(new_n3438_));
  INV    g02436(.A(\A[585] ), .Y(new_n3439_));
  INV    g02437(.A(\A[584] ), .Y(new_n3440_));
  NAND2  g02438(.A(new_n3440_), .B(\A[583] ), .Y(new_n3441_));
  INV    g02439(.A(\A[583] ), .Y(new_n3442_));
  AOI21  g02440(.A0(\A[584] ), .A1(new_n3442_), .B0(new_n3439_), .Y(new_n3443_));
  XOR2   g02441(.A(\A[584] ), .B(\A[583] ), .Y(new_n3444_));
  AOI22  g02442(.A0(new_n3444_), .A1(new_n3439_), .B0(new_n3443_), .B1(new_n3441_), .Y(new_n3445_));
  INV    g02443(.A(\A[588] ), .Y(new_n3446_));
  INV    g02444(.A(\A[587] ), .Y(new_n3447_));
  NAND2  g02445(.A(new_n3447_), .B(\A[586] ), .Y(new_n3448_));
  INV    g02446(.A(\A[586] ), .Y(new_n3449_));
  AOI21  g02447(.A0(\A[587] ), .A1(new_n3449_), .B0(new_n3446_), .Y(new_n3450_));
  XOR2   g02448(.A(\A[587] ), .B(\A[586] ), .Y(new_n3451_));
  AOI22  g02449(.A0(new_n3451_), .A1(new_n3446_), .B0(new_n3450_), .B1(new_n3448_), .Y(new_n3452_));
  NOR2   g02450(.A(new_n3447_), .B(new_n3449_), .Y(new_n3453_));
  AOI21  g02451(.A0(new_n3451_), .A1(\A[588] ), .B0(new_n3453_), .Y(new_n3454_));
  NOR2   g02452(.A(new_n3440_), .B(new_n3442_), .Y(new_n3455_));
  AOI21  g02453(.A0(new_n3444_), .A1(\A[585] ), .B0(new_n3455_), .Y(new_n3456_));
  XOR2   g02454(.A(new_n3452_), .B(new_n3445_), .Y(new_n3457_));
  XOR2   g02455(.A(new_n3457_), .B(new_n3438_), .Y(new_n3458_));
  INV    g02456(.A(new_n3458_), .Y(new_n3459_));
  XOR2   g02457(.A(new_n3459_), .B(new_n3419_), .Y(new_n3460_));
  INV    g02458(.A(new_n3460_), .Y(new_n3461_));
  INV    g02459(.A(\A[579] ), .Y(new_n3462_));
  INV    g02460(.A(\A[578] ), .Y(new_n3463_));
  NAND2  g02461(.A(new_n3463_), .B(\A[577] ), .Y(new_n3464_));
  INV    g02462(.A(\A[577] ), .Y(new_n3465_));
  AOI21  g02463(.A0(\A[578] ), .A1(new_n3465_), .B0(new_n3462_), .Y(new_n3466_));
  XOR2   g02464(.A(\A[578] ), .B(\A[577] ), .Y(new_n3467_));
  AOI22  g02465(.A0(new_n3467_), .A1(new_n3462_), .B0(new_n3466_), .B1(new_n3464_), .Y(new_n3468_));
  INV    g02466(.A(\A[582] ), .Y(new_n3469_));
  INV    g02467(.A(\A[581] ), .Y(new_n3470_));
  NAND2  g02468(.A(new_n3470_), .B(\A[580] ), .Y(new_n3471_));
  INV    g02469(.A(\A[580] ), .Y(new_n3472_));
  AOI21  g02470(.A0(\A[581] ), .A1(new_n3472_), .B0(new_n3469_), .Y(new_n3473_));
  XOR2   g02471(.A(\A[581] ), .B(\A[580] ), .Y(new_n3474_));
  AOI22  g02472(.A0(new_n3474_), .A1(new_n3469_), .B0(new_n3473_), .B1(new_n3471_), .Y(new_n3475_));
  NOR2   g02473(.A(new_n3470_), .B(new_n3472_), .Y(new_n3476_));
  AOI21  g02474(.A0(new_n3474_), .A1(\A[582] ), .B0(new_n3476_), .Y(new_n3477_));
  NOR2   g02475(.A(new_n3463_), .B(new_n3465_), .Y(new_n3478_));
  AOI21  g02476(.A0(new_n3467_), .A1(\A[579] ), .B0(new_n3478_), .Y(new_n3479_));
  XOR2   g02477(.A(new_n3475_), .B(new_n3468_), .Y(new_n3480_));
  INV    g02478(.A(\A[573] ), .Y(new_n3481_));
  INV    g02479(.A(\A[572] ), .Y(new_n3482_));
  NAND2  g02480(.A(new_n3482_), .B(\A[571] ), .Y(new_n3483_));
  INV    g02481(.A(\A[571] ), .Y(new_n3484_));
  AOI21  g02482(.A0(\A[572] ), .A1(new_n3484_), .B0(new_n3481_), .Y(new_n3485_));
  XOR2   g02483(.A(\A[572] ), .B(\A[571] ), .Y(new_n3486_));
  AOI22  g02484(.A0(new_n3486_), .A1(new_n3481_), .B0(new_n3485_), .B1(new_n3483_), .Y(new_n3487_));
  INV    g02485(.A(\A[576] ), .Y(new_n3488_));
  INV    g02486(.A(\A[575] ), .Y(new_n3489_));
  NAND2  g02487(.A(new_n3489_), .B(\A[574] ), .Y(new_n3490_));
  INV    g02488(.A(\A[574] ), .Y(new_n3491_));
  AOI21  g02489(.A0(\A[575] ), .A1(new_n3491_), .B0(new_n3488_), .Y(new_n3492_));
  XOR2   g02490(.A(\A[575] ), .B(\A[574] ), .Y(new_n3493_));
  AOI22  g02491(.A0(new_n3493_), .A1(new_n3488_), .B0(new_n3492_), .B1(new_n3490_), .Y(new_n3494_));
  NOR2   g02492(.A(new_n3489_), .B(new_n3491_), .Y(new_n3495_));
  AOI21  g02493(.A0(new_n3493_), .A1(\A[576] ), .B0(new_n3495_), .Y(new_n3496_));
  NOR2   g02494(.A(new_n3482_), .B(new_n3484_), .Y(new_n3497_));
  AOI21  g02495(.A0(new_n3486_), .A1(\A[573] ), .B0(new_n3497_), .Y(new_n3498_));
  XOR2   g02496(.A(new_n3494_), .B(new_n3487_), .Y(new_n3499_));
  XOR2   g02497(.A(new_n3499_), .B(new_n3480_), .Y(new_n3500_));
  INV    g02498(.A(\A[567] ), .Y(new_n3501_));
  INV    g02499(.A(\A[566] ), .Y(new_n3502_));
  NAND2  g02500(.A(new_n3502_), .B(\A[565] ), .Y(new_n3503_));
  INV    g02501(.A(\A[565] ), .Y(new_n3504_));
  AOI21  g02502(.A0(\A[566] ), .A1(new_n3504_), .B0(new_n3501_), .Y(new_n3505_));
  XOR2   g02503(.A(\A[566] ), .B(\A[565] ), .Y(new_n3506_));
  AOI22  g02504(.A0(new_n3506_), .A1(new_n3501_), .B0(new_n3505_), .B1(new_n3503_), .Y(new_n3507_));
  INV    g02505(.A(\A[570] ), .Y(new_n3508_));
  INV    g02506(.A(\A[569] ), .Y(new_n3509_));
  NAND2  g02507(.A(new_n3509_), .B(\A[568] ), .Y(new_n3510_));
  INV    g02508(.A(\A[568] ), .Y(new_n3511_));
  AOI21  g02509(.A0(\A[569] ), .A1(new_n3511_), .B0(new_n3508_), .Y(new_n3512_));
  XOR2   g02510(.A(\A[569] ), .B(\A[568] ), .Y(new_n3513_));
  AOI22  g02511(.A0(new_n3513_), .A1(new_n3508_), .B0(new_n3512_), .B1(new_n3510_), .Y(new_n3514_));
  NOR2   g02512(.A(new_n3509_), .B(new_n3511_), .Y(new_n3515_));
  AOI21  g02513(.A0(new_n3513_), .A1(\A[570] ), .B0(new_n3515_), .Y(new_n3516_));
  NOR2   g02514(.A(new_n3502_), .B(new_n3504_), .Y(new_n3517_));
  AOI21  g02515(.A0(new_n3506_), .A1(\A[567] ), .B0(new_n3517_), .Y(new_n3518_));
  XOR2   g02516(.A(new_n3514_), .B(new_n3507_), .Y(new_n3519_));
  INV    g02517(.A(\A[561] ), .Y(new_n3520_));
  INV    g02518(.A(\A[560] ), .Y(new_n3521_));
  NAND2  g02519(.A(new_n3521_), .B(\A[559] ), .Y(new_n3522_));
  INV    g02520(.A(\A[559] ), .Y(new_n3523_));
  AOI21  g02521(.A0(\A[560] ), .A1(new_n3523_), .B0(new_n3520_), .Y(new_n3524_));
  XOR2   g02522(.A(\A[560] ), .B(\A[559] ), .Y(new_n3525_));
  AOI22  g02523(.A0(new_n3525_), .A1(new_n3520_), .B0(new_n3524_), .B1(new_n3522_), .Y(new_n3526_));
  INV    g02524(.A(\A[564] ), .Y(new_n3527_));
  INV    g02525(.A(\A[563] ), .Y(new_n3528_));
  NAND2  g02526(.A(new_n3528_), .B(\A[562] ), .Y(new_n3529_));
  INV    g02527(.A(\A[562] ), .Y(new_n3530_));
  AOI21  g02528(.A0(\A[563] ), .A1(new_n3530_), .B0(new_n3527_), .Y(new_n3531_));
  XOR2   g02529(.A(\A[563] ), .B(\A[562] ), .Y(new_n3532_));
  AOI22  g02530(.A0(new_n3532_), .A1(new_n3527_), .B0(new_n3531_), .B1(new_n3529_), .Y(new_n3533_));
  NOR2   g02531(.A(new_n3528_), .B(new_n3530_), .Y(new_n3534_));
  AOI21  g02532(.A0(new_n3532_), .A1(\A[564] ), .B0(new_n3534_), .Y(new_n3535_));
  NOR2   g02533(.A(new_n3521_), .B(new_n3523_), .Y(new_n3536_));
  AOI21  g02534(.A0(new_n3525_), .A1(\A[561] ), .B0(new_n3536_), .Y(new_n3537_));
  XOR2   g02535(.A(new_n3533_), .B(new_n3526_), .Y(new_n3538_));
  XOR2   g02536(.A(new_n3538_), .B(new_n3519_), .Y(new_n3539_));
  INV    g02537(.A(new_n3539_), .Y(new_n3540_));
  XOR2   g02538(.A(new_n3540_), .B(new_n3500_), .Y(new_n3541_));
  XOR2   g02539(.A(new_n3541_), .B(new_n3461_), .Y(new_n3542_));
  XOR2   g02540(.A(new_n3542_), .B(new_n3380_), .Y(new_n3543_));
  XOR2   g02541(.A(new_n3543_), .B(new_n3216_), .Y(new_n3544_));
  XOR2   g02542(.A(new_n2855_), .B(new_n2854_), .Y(new_n3545_));
  INV    g02543(.A(new_n3545_), .Y(new_n3546_));
  NOR2   g02544(.A(new_n3546_), .B(new_n3544_), .Y(new_n3547_));
  NAND3  g02545(.A(new_n3547_), .B(new_n2876_), .C(new_n2866_), .Y(new_n3548_));
  NAND3  g02546(.A(new_n2856_), .B(new_n2864_), .C(new_n2861_), .Y(new_n3549_));
  OAI21  g02547(.A0(new_n2852_), .A1(new_n2839_), .B0(new_n2857_), .Y(new_n3550_));
  AOI21  g02548(.A0(new_n3550_), .A1(new_n3549_), .B0(new_n2873_), .Y(new_n3551_));
  NAND3  g02549(.A(new_n2857_), .B(new_n2864_), .C(new_n2861_), .Y(new_n3552_));
  OAI21  g02550(.A0(new_n2852_), .A1(new_n2839_), .B0(new_n2856_), .Y(new_n3553_));
  AOI21  g02551(.A0(new_n3553_), .A1(new_n3552_), .B0(new_n1929_), .Y(new_n3554_));
  INV    g02552(.A(new_n3547_), .Y(new_n3555_));
  OAI21  g02553(.A0(new_n3554_), .A1(new_n3551_), .B0(new_n3555_), .Y(new_n3556_));
  NAND2  g02554(.A(new_n3556_), .B(new_n3548_), .Y(new_n3557_));
  XOR2   g02555(.A(new_n3452_), .B(new_n3445_), .Y(new_n3558_));
  XOR2   g02556(.A(\A[587] ), .B(new_n3449_), .Y(new_n3559_));
  NAND2  g02557(.A(\A[587] ), .B(\A[586] ), .Y(new_n3560_));
  OAI21  g02558(.A0(new_n3559_), .A1(new_n3446_), .B0(new_n3560_), .Y(new_n3561_));
  XOR2   g02559(.A(new_n3456_), .B(new_n3561_), .Y(new_n3562_));
  NOR2   g02560(.A(\A[584] ), .B(new_n3442_), .Y(new_n3563_));
  OAI21  g02561(.A0(new_n3440_), .A1(\A[583] ), .B0(\A[585] ), .Y(new_n3564_));
  XOR2   g02562(.A(\A[584] ), .B(new_n3442_), .Y(new_n3565_));
  OAI22  g02563(.A0(new_n3565_), .A1(\A[585] ), .B0(new_n3564_), .B1(new_n3563_), .Y(new_n3566_));
  NOR2   g02564(.A(\A[587] ), .B(new_n3449_), .Y(new_n3567_));
  OAI21  g02565(.A0(new_n3447_), .A1(\A[586] ), .B0(\A[588] ), .Y(new_n3568_));
  OAI22  g02566(.A0(new_n3559_), .A1(\A[588] ), .B0(new_n3568_), .B1(new_n3567_), .Y(new_n3569_));
  NAND2  g02567(.A(new_n3569_), .B(new_n3566_), .Y(new_n3570_));
  NAND2  g02568(.A(\A[584] ), .B(\A[583] ), .Y(new_n3571_));
  OAI21  g02569(.A0(new_n3565_), .A1(new_n3439_), .B0(new_n3571_), .Y(new_n3572_));
  NAND2  g02570(.A(new_n3572_), .B(new_n3561_), .Y(new_n3573_));
  OAI21  g02571(.A0(new_n3570_), .A1(new_n3562_), .B0(new_n3573_), .Y(new_n3574_));
  NOR2   g02572(.A(new_n3452_), .B(new_n3445_), .Y(new_n3575_));
  XOR2   g02573(.A(new_n3575_), .B(new_n3562_), .Y(new_n3576_));
  AOI21  g02574(.A0(new_n3574_), .A1(new_n3558_), .B0(new_n3576_), .Y(new_n3577_));
  XOR2   g02575(.A(new_n3433_), .B(new_n3426_), .Y(new_n3578_));
  NOR2   g02576(.A(\A[590] ), .B(new_n3423_), .Y(new_n3579_));
  OAI21  g02577(.A0(new_n3421_), .A1(\A[589] ), .B0(\A[591] ), .Y(new_n3580_));
  NAND2  g02578(.A(new_n3425_), .B(new_n3420_), .Y(new_n3581_));
  OAI21  g02579(.A0(new_n3580_), .A1(new_n3579_), .B0(new_n3581_), .Y(new_n3582_));
  NOR2   g02580(.A(\A[593] ), .B(new_n3430_), .Y(new_n3583_));
  OAI21  g02581(.A0(new_n3428_), .A1(\A[592] ), .B0(\A[594] ), .Y(new_n3584_));
  NAND2  g02582(.A(new_n3432_), .B(new_n3427_), .Y(new_n3585_));
  OAI21  g02583(.A0(new_n3584_), .A1(new_n3583_), .B0(new_n3585_), .Y(new_n3586_));
  NAND2  g02584(.A(new_n3432_), .B(\A[594] ), .Y(new_n3587_));
  OAI21  g02585(.A0(new_n3428_), .A1(new_n3430_), .B0(new_n3587_), .Y(new_n3588_));
  NAND2  g02586(.A(new_n3425_), .B(\A[591] ), .Y(new_n3589_));
  OAI21  g02587(.A0(new_n3421_), .A1(new_n3423_), .B0(new_n3589_), .Y(new_n3590_));
  NAND4  g02588(.A(new_n3590_), .B(new_n3588_), .C(new_n3586_), .D(new_n3582_), .Y(new_n3591_));
  NAND4  g02589(.A(new_n3572_), .B(new_n3561_), .C(new_n3569_), .D(new_n3566_), .Y(new_n3592_));
  NAND4  g02590(.A(new_n3592_), .B(new_n3558_), .C(new_n3591_), .D(new_n3578_), .Y(new_n3593_));
  XOR2   g02591(.A(new_n3437_), .B(new_n3588_), .Y(new_n3594_));
  NAND2  g02592(.A(new_n3586_), .B(new_n3582_), .Y(new_n3595_));
  NAND2  g02593(.A(new_n3590_), .B(new_n3588_), .Y(new_n3596_));
  OAI21  g02594(.A0(new_n3595_), .A1(new_n3594_), .B0(new_n3596_), .Y(new_n3597_));
  NOR2   g02595(.A(new_n3433_), .B(new_n3426_), .Y(new_n3598_));
  XOR2   g02596(.A(new_n3598_), .B(new_n3594_), .Y(new_n3599_));
  AOI21  g02597(.A0(new_n3597_), .A1(new_n3578_), .B0(new_n3599_), .Y(new_n3600_));
  XOR2   g02598(.A(new_n3600_), .B(new_n3593_), .Y(new_n3601_));
  XOR2   g02599(.A(new_n3433_), .B(new_n3582_), .Y(new_n3602_));
  NOR4   g02600(.A(new_n3437_), .B(new_n3435_), .C(new_n3433_), .D(new_n3426_), .Y(new_n3603_));
  XOR2   g02601(.A(new_n3452_), .B(new_n3566_), .Y(new_n3604_));
  NOR4   g02602(.A(new_n3456_), .B(new_n3454_), .C(new_n3452_), .D(new_n3445_), .Y(new_n3605_));
  NOR4   g02603(.A(new_n3605_), .B(new_n3604_), .C(new_n3603_), .D(new_n3602_), .Y(new_n3606_));
  XOR2   g02604(.A(new_n3437_), .B(new_n3435_), .Y(new_n3607_));
  NOR2   g02605(.A(new_n3437_), .B(new_n3435_), .Y(new_n3608_));
  AOI21  g02606(.A0(new_n3598_), .A1(new_n3607_), .B0(new_n3608_), .Y(new_n3609_));
  NOR4   g02607(.A(new_n3604_), .B(new_n3603_), .C(new_n3599_), .D(new_n3602_), .Y(new_n3610_));
  OAI211 g02608(.A0(new_n3609_), .A1(new_n3602_), .B0(new_n3610_), .B1(new_n3592_), .Y(new_n3611_));
  OAI21  g02609(.A0(new_n3600_), .A1(new_n3606_), .B0(new_n3611_), .Y(new_n3612_));
  NAND2  g02610(.A(new_n3612_), .B(new_n3577_), .Y(new_n3613_));
  OAI21  g02611(.A0(new_n3601_), .A1(new_n3577_), .B0(new_n3613_), .Y(new_n3614_));
  NOR2   g02612(.A(\A[596] ), .B(new_n3403_), .Y(new_n3615_));
  OAI21  g02613(.A0(new_n3401_), .A1(\A[595] ), .B0(\A[597] ), .Y(new_n3616_));
  XOR2   g02614(.A(\A[596] ), .B(new_n3403_), .Y(new_n3617_));
  OAI22  g02615(.A0(new_n3617_), .A1(\A[597] ), .B0(new_n3616_), .B1(new_n3615_), .Y(new_n3618_));
  XOR2   g02616(.A(new_n3413_), .B(new_n3618_), .Y(new_n3619_));
  XOR2   g02617(.A(new_n3417_), .B(new_n3415_), .Y(new_n3620_));
  NOR2   g02618(.A(new_n3413_), .B(new_n3406_), .Y(new_n3621_));
  NOR2   g02619(.A(new_n3417_), .B(new_n3415_), .Y(new_n3622_));
  AOI21  g02620(.A0(new_n3621_), .A1(new_n3620_), .B0(new_n3622_), .Y(new_n3623_));
  XOR2   g02621(.A(new_n3621_), .B(new_n3620_), .Y(new_n3624_));
  OAI21  g02622(.A0(new_n3623_), .A1(new_n3619_), .B0(new_n3624_), .Y(new_n3625_));
  NOR2   g02623(.A(\A[602] ), .B(new_n3384_), .Y(new_n3626_));
  OAI21  g02624(.A0(new_n3382_), .A1(\A[601] ), .B0(\A[603] ), .Y(new_n3627_));
  NAND2  g02625(.A(new_n3386_), .B(new_n3381_), .Y(new_n3628_));
  OAI21  g02626(.A0(new_n3627_), .A1(new_n3626_), .B0(new_n3628_), .Y(new_n3629_));
  XOR2   g02627(.A(new_n3394_), .B(new_n3629_), .Y(new_n3630_));
  NOR4   g02628(.A(new_n3398_), .B(new_n3396_), .C(new_n3394_), .D(new_n3387_), .Y(new_n3631_));
  NOR4   g02629(.A(new_n3417_), .B(new_n3415_), .C(new_n3413_), .D(new_n3406_), .Y(new_n3632_));
  NOR4   g02630(.A(new_n3632_), .B(new_n3619_), .C(new_n3631_), .D(new_n3630_), .Y(new_n3633_));
  XOR2   g02631(.A(new_n3394_), .B(new_n3387_), .Y(new_n3634_));
  NAND2  g02632(.A(new_n3393_), .B(\A[606] ), .Y(new_n3635_));
  OAI21  g02633(.A0(new_n3389_), .A1(new_n3391_), .B0(new_n3635_), .Y(new_n3636_));
  XOR2   g02634(.A(new_n3398_), .B(new_n3636_), .Y(new_n3637_));
  NOR2   g02635(.A(\A[605] ), .B(new_n3391_), .Y(new_n3638_));
  OAI21  g02636(.A0(new_n3389_), .A1(\A[604] ), .B0(\A[606] ), .Y(new_n3639_));
  NAND2  g02637(.A(new_n3393_), .B(new_n3388_), .Y(new_n3640_));
  OAI21  g02638(.A0(new_n3639_), .A1(new_n3638_), .B0(new_n3640_), .Y(new_n3641_));
  NAND2  g02639(.A(new_n3641_), .B(new_n3629_), .Y(new_n3642_));
  NAND2  g02640(.A(new_n3386_), .B(\A[603] ), .Y(new_n3643_));
  OAI21  g02641(.A0(new_n3382_), .A1(new_n3384_), .B0(new_n3643_), .Y(new_n3644_));
  NAND2  g02642(.A(new_n3644_), .B(new_n3636_), .Y(new_n3645_));
  OAI21  g02643(.A0(new_n3642_), .A1(new_n3637_), .B0(new_n3645_), .Y(new_n3646_));
  NOR2   g02644(.A(new_n3394_), .B(new_n3387_), .Y(new_n3647_));
  XOR2   g02645(.A(new_n3647_), .B(new_n3637_), .Y(new_n3648_));
  AOI21  g02646(.A0(new_n3646_), .A1(new_n3634_), .B0(new_n3648_), .Y(new_n3649_));
  XOR2   g02647(.A(new_n3649_), .B(new_n3633_), .Y(new_n3650_));
  NAND2  g02648(.A(new_n3650_), .B(new_n3625_), .Y(new_n3651_));
  XOR2   g02649(.A(new_n3413_), .B(new_n3406_), .Y(new_n3652_));
  XOR2   g02650(.A(\A[599] ), .B(new_n3410_), .Y(new_n3653_));
  NAND2  g02651(.A(\A[599] ), .B(\A[598] ), .Y(new_n3654_));
  OAI21  g02652(.A0(new_n3653_), .A1(new_n3407_), .B0(new_n3654_), .Y(new_n3655_));
  XOR2   g02653(.A(new_n3417_), .B(new_n3655_), .Y(new_n3656_));
  NOR2   g02654(.A(\A[599] ), .B(new_n3410_), .Y(new_n3657_));
  OAI21  g02655(.A0(new_n3408_), .A1(\A[598] ), .B0(\A[600] ), .Y(new_n3658_));
  OAI22  g02656(.A0(new_n3653_), .A1(\A[600] ), .B0(new_n3658_), .B1(new_n3657_), .Y(new_n3659_));
  NAND2  g02657(.A(new_n3659_), .B(new_n3618_), .Y(new_n3660_));
  NAND2  g02658(.A(\A[596] ), .B(\A[595] ), .Y(new_n3661_));
  OAI21  g02659(.A0(new_n3617_), .A1(new_n3400_), .B0(new_n3661_), .Y(new_n3662_));
  NAND2  g02660(.A(new_n3662_), .B(new_n3655_), .Y(new_n3663_));
  OAI21  g02661(.A0(new_n3660_), .A1(new_n3656_), .B0(new_n3663_), .Y(new_n3664_));
  XOR2   g02662(.A(new_n3621_), .B(new_n3656_), .Y(new_n3665_));
  AOI21  g02663(.A0(new_n3664_), .A1(new_n3652_), .B0(new_n3665_), .Y(new_n3666_));
  XOR2   g02664(.A(new_n3398_), .B(new_n3396_), .Y(new_n3667_));
  XOR2   g02665(.A(new_n3647_), .B(new_n3667_), .Y(new_n3668_));
  NAND4  g02666(.A(new_n3644_), .B(new_n3636_), .C(new_n3641_), .D(new_n3629_), .Y(new_n3669_));
  NAND4  g02667(.A(new_n3652_), .B(new_n3669_), .C(new_n3668_), .D(new_n3634_), .Y(new_n3670_));
  NOR2   g02668(.A(new_n3398_), .B(new_n3396_), .Y(new_n3671_));
  AOI21  g02669(.A0(new_n3647_), .A1(new_n3667_), .B0(new_n3671_), .Y(new_n3672_));
  NAND4  g02670(.A(new_n3662_), .B(new_n3655_), .C(new_n3659_), .D(new_n3618_), .Y(new_n3673_));
  OAI21  g02671(.A0(new_n3672_), .A1(new_n3630_), .B0(new_n3673_), .Y(new_n3674_));
  OAI22  g02672(.A0(new_n3674_), .A1(new_n3670_), .B0(new_n3649_), .B1(new_n3633_), .Y(new_n3675_));
  NAND2  g02673(.A(new_n3675_), .B(new_n3666_), .Y(new_n3676_));
  NAND2  g02674(.A(new_n3458_), .B(new_n3419_), .Y(new_n3677_));
  INV    g02675(.A(new_n3677_), .Y(new_n3678_));
  NAND3  g02676(.A(new_n3678_), .B(new_n3676_), .C(new_n3651_), .Y(new_n3679_));
  NAND2  g02677(.A(new_n3676_), .B(new_n3651_), .Y(new_n3680_));
  NAND2  g02678(.A(new_n3680_), .B(new_n3677_), .Y(new_n3681_));
  AOI21  g02679(.A0(new_n3681_), .A1(new_n3679_), .B0(new_n3614_), .Y(new_n3682_));
  NOR2   g02680(.A(new_n3601_), .B(new_n3577_), .Y(new_n3683_));
  AOI21  g02681(.A0(new_n3612_), .A1(new_n3577_), .B0(new_n3683_), .Y(new_n3684_));
  NAND4  g02682(.A(new_n3673_), .B(new_n3652_), .C(new_n3669_), .D(new_n3634_), .Y(new_n3685_));
  XOR2   g02683(.A(new_n3649_), .B(new_n3685_), .Y(new_n3686_));
  NOR2   g02684(.A(new_n3686_), .B(new_n3666_), .Y(new_n3687_));
  AOI211 g02685(.A0(new_n3675_), .A1(new_n3666_), .B(new_n3678_), .C(new_n3687_), .Y(new_n3688_));
  AOI21  g02686(.A0(new_n3676_), .A1(new_n3651_), .B0(new_n3677_), .Y(new_n3689_));
  NOR2   g02687(.A(new_n3689_), .B(new_n3688_), .Y(new_n3690_));
  NOR2   g02688(.A(new_n3541_), .B(new_n3460_), .Y(new_n3691_));
  OAI21  g02689(.A0(new_n3690_), .A1(new_n3684_), .B0(new_n3691_), .Y(new_n3692_));
  NOR2   g02690(.A(new_n3690_), .B(new_n3684_), .Y(new_n3693_));
  INV    g02691(.A(new_n3691_), .Y(new_n3694_));
  OAI21  g02692(.A0(new_n3693_), .A1(new_n3682_), .B0(new_n3694_), .Y(new_n3695_));
  OAI21  g02693(.A0(new_n3692_), .A1(new_n3682_), .B0(new_n3695_), .Y(new_n3696_));
  XOR2   g02694(.A(new_n3533_), .B(new_n3526_), .Y(new_n3697_));
  XOR2   g02695(.A(\A[563] ), .B(new_n3530_), .Y(new_n3698_));
  NAND2  g02696(.A(\A[563] ), .B(\A[562] ), .Y(new_n3699_));
  OAI21  g02697(.A0(new_n3698_), .A1(new_n3527_), .B0(new_n3699_), .Y(new_n3700_));
  XOR2   g02698(.A(new_n3537_), .B(new_n3700_), .Y(new_n3701_));
  NOR2   g02699(.A(\A[560] ), .B(new_n3523_), .Y(new_n3702_));
  OAI21  g02700(.A0(new_n3521_), .A1(\A[559] ), .B0(\A[561] ), .Y(new_n3703_));
  XOR2   g02701(.A(\A[560] ), .B(new_n3523_), .Y(new_n3704_));
  OAI22  g02702(.A0(new_n3704_), .A1(\A[561] ), .B0(new_n3703_), .B1(new_n3702_), .Y(new_n3705_));
  NOR2   g02703(.A(\A[563] ), .B(new_n3530_), .Y(new_n3706_));
  OAI21  g02704(.A0(new_n3528_), .A1(\A[562] ), .B0(\A[564] ), .Y(new_n3707_));
  OAI22  g02705(.A0(new_n3698_), .A1(\A[564] ), .B0(new_n3707_), .B1(new_n3706_), .Y(new_n3708_));
  NAND2  g02706(.A(new_n3708_), .B(new_n3705_), .Y(new_n3709_));
  NAND2  g02707(.A(\A[560] ), .B(\A[559] ), .Y(new_n3710_));
  OAI21  g02708(.A0(new_n3704_), .A1(new_n3520_), .B0(new_n3710_), .Y(new_n3711_));
  NAND2  g02709(.A(new_n3711_), .B(new_n3700_), .Y(new_n3712_));
  OAI21  g02710(.A0(new_n3709_), .A1(new_n3701_), .B0(new_n3712_), .Y(new_n3713_));
  NOR2   g02711(.A(new_n3533_), .B(new_n3526_), .Y(new_n3714_));
  XOR2   g02712(.A(new_n3714_), .B(new_n3701_), .Y(new_n3715_));
  AOI21  g02713(.A0(new_n3713_), .A1(new_n3697_), .B0(new_n3715_), .Y(new_n3716_));
  XOR2   g02714(.A(new_n3514_), .B(new_n3507_), .Y(new_n3717_));
  NOR2   g02715(.A(\A[566] ), .B(new_n3504_), .Y(new_n3718_));
  OAI21  g02716(.A0(new_n3502_), .A1(\A[565] ), .B0(\A[567] ), .Y(new_n3719_));
  NAND2  g02717(.A(new_n3506_), .B(new_n3501_), .Y(new_n3720_));
  OAI21  g02718(.A0(new_n3719_), .A1(new_n3718_), .B0(new_n3720_), .Y(new_n3721_));
  NOR2   g02719(.A(\A[569] ), .B(new_n3511_), .Y(new_n3722_));
  OAI21  g02720(.A0(new_n3509_), .A1(\A[568] ), .B0(\A[570] ), .Y(new_n3723_));
  NAND2  g02721(.A(new_n3513_), .B(new_n3508_), .Y(new_n3724_));
  OAI21  g02722(.A0(new_n3723_), .A1(new_n3722_), .B0(new_n3724_), .Y(new_n3725_));
  NAND2  g02723(.A(new_n3513_), .B(\A[570] ), .Y(new_n3726_));
  OAI21  g02724(.A0(new_n3509_), .A1(new_n3511_), .B0(new_n3726_), .Y(new_n3727_));
  NAND2  g02725(.A(new_n3506_), .B(\A[567] ), .Y(new_n3728_));
  OAI21  g02726(.A0(new_n3502_), .A1(new_n3504_), .B0(new_n3728_), .Y(new_n3729_));
  NAND4  g02727(.A(new_n3729_), .B(new_n3727_), .C(new_n3725_), .D(new_n3721_), .Y(new_n3730_));
  NAND4  g02728(.A(new_n3711_), .B(new_n3700_), .C(new_n3708_), .D(new_n3705_), .Y(new_n3731_));
  NAND4  g02729(.A(new_n3731_), .B(new_n3697_), .C(new_n3730_), .D(new_n3717_), .Y(new_n3732_));
  XOR2   g02730(.A(new_n3518_), .B(new_n3727_), .Y(new_n3733_));
  NAND2  g02731(.A(new_n3725_), .B(new_n3721_), .Y(new_n3734_));
  NAND2  g02732(.A(new_n3729_), .B(new_n3727_), .Y(new_n3735_));
  OAI21  g02733(.A0(new_n3734_), .A1(new_n3733_), .B0(new_n3735_), .Y(new_n3736_));
  NOR2   g02734(.A(new_n3514_), .B(new_n3507_), .Y(new_n3737_));
  XOR2   g02735(.A(new_n3737_), .B(new_n3733_), .Y(new_n3738_));
  AOI21  g02736(.A0(new_n3736_), .A1(new_n3717_), .B0(new_n3738_), .Y(new_n3739_));
  XOR2   g02737(.A(new_n3739_), .B(new_n3732_), .Y(new_n3740_));
  XOR2   g02738(.A(new_n3514_), .B(new_n3721_), .Y(new_n3741_));
  NOR4   g02739(.A(new_n3518_), .B(new_n3516_), .C(new_n3514_), .D(new_n3507_), .Y(new_n3742_));
  XOR2   g02740(.A(new_n3533_), .B(new_n3705_), .Y(new_n3743_));
  NOR4   g02741(.A(new_n3537_), .B(new_n3535_), .C(new_n3533_), .D(new_n3526_), .Y(new_n3744_));
  NOR4   g02742(.A(new_n3744_), .B(new_n3743_), .C(new_n3742_), .D(new_n3741_), .Y(new_n3745_));
  XOR2   g02743(.A(new_n3518_), .B(new_n3516_), .Y(new_n3746_));
  NOR2   g02744(.A(new_n3518_), .B(new_n3516_), .Y(new_n3747_));
  AOI21  g02745(.A0(new_n3737_), .A1(new_n3746_), .B0(new_n3747_), .Y(new_n3748_));
  NOR4   g02746(.A(new_n3743_), .B(new_n3742_), .C(new_n3738_), .D(new_n3741_), .Y(new_n3749_));
  OAI211 g02747(.A0(new_n3748_), .A1(new_n3741_), .B0(new_n3749_), .B1(new_n3731_), .Y(new_n3750_));
  OAI21  g02748(.A0(new_n3739_), .A1(new_n3745_), .B0(new_n3750_), .Y(new_n3751_));
  NAND2  g02749(.A(new_n3751_), .B(new_n3716_), .Y(new_n3752_));
  OAI21  g02750(.A0(new_n3740_), .A1(new_n3716_), .B0(new_n3752_), .Y(new_n3753_));
  XOR2   g02751(.A(new_n3494_), .B(new_n3487_), .Y(new_n3754_));
  XOR2   g02752(.A(\A[575] ), .B(new_n3491_), .Y(new_n3755_));
  NAND2  g02753(.A(\A[575] ), .B(\A[574] ), .Y(new_n3756_));
  OAI21  g02754(.A0(new_n3755_), .A1(new_n3488_), .B0(new_n3756_), .Y(new_n3757_));
  XOR2   g02755(.A(new_n3498_), .B(new_n3757_), .Y(new_n3758_));
  NOR2   g02756(.A(\A[572] ), .B(new_n3484_), .Y(new_n3759_));
  OAI21  g02757(.A0(new_n3482_), .A1(\A[571] ), .B0(\A[573] ), .Y(new_n3760_));
  XOR2   g02758(.A(\A[572] ), .B(new_n3484_), .Y(new_n3761_));
  OAI22  g02759(.A0(new_n3761_), .A1(\A[573] ), .B0(new_n3760_), .B1(new_n3759_), .Y(new_n3762_));
  NOR2   g02760(.A(\A[575] ), .B(new_n3491_), .Y(new_n3763_));
  OAI21  g02761(.A0(new_n3489_), .A1(\A[574] ), .B0(\A[576] ), .Y(new_n3764_));
  OAI22  g02762(.A0(new_n3755_), .A1(\A[576] ), .B0(new_n3764_), .B1(new_n3763_), .Y(new_n3765_));
  NAND2  g02763(.A(new_n3765_), .B(new_n3762_), .Y(new_n3766_));
  NAND2  g02764(.A(\A[572] ), .B(\A[571] ), .Y(new_n3767_));
  OAI21  g02765(.A0(new_n3761_), .A1(new_n3481_), .B0(new_n3767_), .Y(new_n3768_));
  NAND2  g02766(.A(new_n3768_), .B(new_n3757_), .Y(new_n3769_));
  OAI21  g02767(.A0(new_n3766_), .A1(new_n3758_), .B0(new_n3769_), .Y(new_n3770_));
  NOR2   g02768(.A(new_n3494_), .B(new_n3487_), .Y(new_n3771_));
  XOR2   g02769(.A(new_n3771_), .B(new_n3758_), .Y(new_n3772_));
  AOI21  g02770(.A0(new_n3770_), .A1(new_n3754_), .B0(new_n3772_), .Y(new_n3773_));
  XOR2   g02771(.A(new_n3475_), .B(new_n3468_), .Y(new_n3774_));
  NOR2   g02772(.A(\A[578] ), .B(new_n3465_), .Y(new_n3775_));
  OAI21  g02773(.A0(new_n3463_), .A1(\A[577] ), .B0(\A[579] ), .Y(new_n3776_));
  NAND2  g02774(.A(new_n3467_), .B(new_n3462_), .Y(new_n3777_));
  OAI21  g02775(.A0(new_n3776_), .A1(new_n3775_), .B0(new_n3777_), .Y(new_n3778_));
  NOR2   g02776(.A(\A[581] ), .B(new_n3472_), .Y(new_n3779_));
  OAI21  g02777(.A0(new_n3470_), .A1(\A[580] ), .B0(\A[582] ), .Y(new_n3780_));
  NAND2  g02778(.A(new_n3474_), .B(new_n3469_), .Y(new_n3781_));
  OAI21  g02779(.A0(new_n3780_), .A1(new_n3779_), .B0(new_n3781_), .Y(new_n3782_));
  NAND2  g02780(.A(new_n3474_), .B(\A[582] ), .Y(new_n3783_));
  OAI21  g02781(.A0(new_n3470_), .A1(new_n3472_), .B0(new_n3783_), .Y(new_n3784_));
  NAND2  g02782(.A(new_n3467_), .B(\A[579] ), .Y(new_n3785_));
  OAI21  g02783(.A0(new_n3463_), .A1(new_n3465_), .B0(new_n3785_), .Y(new_n3786_));
  NAND4  g02784(.A(new_n3786_), .B(new_n3784_), .C(new_n3782_), .D(new_n3778_), .Y(new_n3787_));
  NAND4  g02785(.A(new_n3768_), .B(new_n3757_), .C(new_n3765_), .D(new_n3762_), .Y(new_n3788_));
  NAND4  g02786(.A(new_n3788_), .B(new_n3754_), .C(new_n3787_), .D(new_n3774_), .Y(new_n3789_));
  XOR2   g02787(.A(new_n3479_), .B(new_n3784_), .Y(new_n3790_));
  NAND2  g02788(.A(new_n3782_), .B(new_n3778_), .Y(new_n3791_));
  NAND2  g02789(.A(new_n3786_), .B(new_n3784_), .Y(new_n3792_));
  OAI21  g02790(.A0(new_n3791_), .A1(new_n3790_), .B0(new_n3792_), .Y(new_n3793_));
  NOR2   g02791(.A(new_n3475_), .B(new_n3468_), .Y(new_n3794_));
  XOR2   g02792(.A(new_n3794_), .B(new_n3790_), .Y(new_n3795_));
  AOI21  g02793(.A0(new_n3793_), .A1(new_n3774_), .B0(new_n3795_), .Y(new_n3796_));
  XOR2   g02794(.A(new_n3796_), .B(new_n3789_), .Y(new_n3797_));
  NOR2   g02795(.A(new_n3797_), .B(new_n3773_), .Y(new_n3798_));
  XOR2   g02796(.A(new_n3494_), .B(new_n3762_), .Y(new_n3799_));
  XOR2   g02797(.A(new_n3498_), .B(new_n3496_), .Y(new_n3800_));
  NOR2   g02798(.A(new_n3498_), .B(new_n3496_), .Y(new_n3801_));
  AOI21  g02799(.A0(new_n3771_), .A1(new_n3800_), .B0(new_n3801_), .Y(new_n3802_));
  XOR2   g02800(.A(new_n3771_), .B(new_n3800_), .Y(new_n3803_));
  OAI21  g02801(.A0(new_n3802_), .A1(new_n3799_), .B0(new_n3803_), .Y(new_n3804_));
  XOR2   g02802(.A(new_n3475_), .B(new_n3778_), .Y(new_n3805_));
  XOR2   g02803(.A(new_n3479_), .B(new_n3477_), .Y(new_n3806_));
  NOR2   g02804(.A(new_n3479_), .B(new_n3477_), .Y(new_n3807_));
  AOI21  g02805(.A0(new_n3794_), .A1(new_n3806_), .B0(new_n3807_), .Y(new_n3808_));
  XOR2   g02806(.A(new_n3794_), .B(new_n3806_), .Y(new_n3809_));
  OAI21  g02807(.A0(new_n3808_), .A1(new_n3805_), .B0(new_n3809_), .Y(new_n3810_));
  NAND2  g02808(.A(new_n3810_), .B(new_n3789_), .Y(new_n3811_));
  NOR4   g02809(.A(new_n3479_), .B(new_n3477_), .C(new_n3475_), .D(new_n3468_), .Y(new_n3812_));
  NOR4   g02810(.A(new_n3799_), .B(new_n3812_), .C(new_n3795_), .D(new_n3805_), .Y(new_n3813_));
  OAI211 g02811(.A0(new_n3808_), .A1(new_n3805_), .B0(new_n3813_), .B1(new_n3788_), .Y(new_n3814_));
  AOI21  g02812(.A0(new_n3814_), .A1(new_n3811_), .B0(new_n3804_), .Y(new_n3815_));
  NAND2  g02813(.A(new_n3539_), .B(new_n3500_), .Y(new_n3816_));
  NOR3   g02814(.A(new_n3816_), .B(new_n3815_), .C(new_n3798_), .Y(new_n3817_));
  NOR4   g02815(.A(new_n3498_), .B(new_n3496_), .C(new_n3494_), .D(new_n3487_), .Y(new_n3818_));
  NOR4   g02816(.A(new_n3818_), .B(new_n3799_), .C(new_n3812_), .D(new_n3805_), .Y(new_n3819_));
  XOR2   g02817(.A(new_n3796_), .B(new_n3819_), .Y(new_n3820_));
  NAND2  g02818(.A(new_n3820_), .B(new_n3804_), .Y(new_n3821_));
  NAND4  g02819(.A(new_n3754_), .B(new_n3787_), .C(new_n3809_), .D(new_n3774_), .Y(new_n3822_));
  OAI21  g02820(.A0(new_n3808_), .A1(new_n3805_), .B0(new_n3788_), .Y(new_n3823_));
  OAI22  g02821(.A0(new_n3823_), .A1(new_n3822_), .B0(new_n3796_), .B1(new_n3819_), .Y(new_n3824_));
  NAND2  g02822(.A(new_n3824_), .B(new_n3773_), .Y(new_n3825_));
  INV    g02823(.A(new_n3816_), .Y(new_n3826_));
  AOI21  g02824(.A0(new_n3825_), .A1(new_n3821_), .B0(new_n3826_), .Y(new_n3827_));
  NOR2   g02825(.A(new_n3827_), .B(new_n3817_), .Y(new_n3828_));
  NOR2   g02826(.A(new_n3753_), .B(new_n3828_), .Y(new_n3829_));
  NOR2   g02827(.A(new_n3815_), .B(new_n3798_), .Y(new_n3830_));
  NAND3  g02828(.A(new_n3816_), .B(new_n3825_), .C(new_n3821_), .Y(new_n3831_));
  OAI21  g02829(.A0(new_n3830_), .A1(new_n3816_), .B0(new_n3831_), .Y(new_n3832_));
  AOI21  g02830(.A0(new_n3832_), .A1(new_n3753_), .B0(new_n3829_), .Y(new_n3833_));
  AOI21  g02831(.A0(new_n3675_), .A1(new_n3666_), .B0(new_n3687_), .Y(new_n3834_));
  OAI21  g02832(.A0(new_n3834_), .A1(new_n3678_), .B0(new_n3679_), .Y(new_n3835_));
  NAND2  g02833(.A(new_n3835_), .B(new_n3684_), .Y(new_n3836_));
  NAND3  g02834(.A(new_n3677_), .B(new_n3676_), .C(new_n3651_), .Y(new_n3837_));
  OAI21  g02835(.A0(new_n3834_), .A1(new_n3677_), .B0(new_n3837_), .Y(new_n3838_));
  AOI21  g02836(.A0(new_n3838_), .A1(new_n3614_), .B0(new_n3691_), .Y(new_n3839_));
  NAND2  g02837(.A(new_n3839_), .B(new_n3836_), .Y(new_n3840_));
  OAI21  g02838(.A0(new_n3693_), .A1(new_n3682_), .B0(new_n3691_), .Y(new_n3841_));
  AOI21  g02839(.A0(new_n3841_), .A1(new_n3840_), .B0(new_n3833_), .Y(new_n3842_));
  AOI21  g02840(.A0(new_n3833_), .A1(new_n3696_), .B0(new_n3842_), .Y(new_n3843_));
  XOR2   g02841(.A(new_n3331_), .B(new_n3324_), .Y(new_n3844_));
  XOR2   g02842(.A(\A[623] ), .B(new_n3328_), .Y(new_n3845_));
  NAND2  g02843(.A(\A[623] ), .B(\A[622] ), .Y(new_n3846_));
  OAI21  g02844(.A0(new_n3845_), .A1(new_n3325_), .B0(new_n3846_), .Y(new_n3847_));
  XOR2   g02845(.A(new_n3335_), .B(new_n3847_), .Y(new_n3848_));
  NOR2   g02846(.A(\A[620] ), .B(new_n3321_), .Y(new_n3849_));
  OAI21  g02847(.A0(new_n3319_), .A1(\A[619] ), .B0(\A[621] ), .Y(new_n3850_));
  XOR2   g02848(.A(\A[620] ), .B(new_n3321_), .Y(new_n3851_));
  OAI22  g02849(.A0(new_n3851_), .A1(\A[621] ), .B0(new_n3850_), .B1(new_n3849_), .Y(new_n3852_));
  NOR2   g02850(.A(\A[623] ), .B(new_n3328_), .Y(new_n3853_));
  OAI21  g02851(.A0(new_n3326_), .A1(\A[622] ), .B0(\A[624] ), .Y(new_n3854_));
  OAI22  g02852(.A0(new_n3845_), .A1(\A[624] ), .B0(new_n3854_), .B1(new_n3853_), .Y(new_n3855_));
  NAND2  g02853(.A(new_n3855_), .B(new_n3852_), .Y(new_n3856_));
  NAND2  g02854(.A(\A[620] ), .B(\A[619] ), .Y(new_n3857_));
  OAI21  g02855(.A0(new_n3851_), .A1(new_n3318_), .B0(new_n3857_), .Y(new_n3858_));
  NAND2  g02856(.A(new_n3858_), .B(new_n3847_), .Y(new_n3859_));
  OAI21  g02857(.A0(new_n3856_), .A1(new_n3848_), .B0(new_n3859_), .Y(new_n3860_));
  NOR2   g02858(.A(new_n3331_), .B(new_n3324_), .Y(new_n3861_));
  XOR2   g02859(.A(new_n3861_), .B(new_n3848_), .Y(new_n3862_));
  AOI21  g02860(.A0(new_n3860_), .A1(new_n3844_), .B0(new_n3862_), .Y(new_n3863_));
  XOR2   g02861(.A(new_n3312_), .B(new_n3305_), .Y(new_n3864_));
  NOR2   g02862(.A(\A[626] ), .B(new_n3302_), .Y(new_n3865_));
  OAI21  g02863(.A0(new_n3300_), .A1(\A[625] ), .B0(\A[627] ), .Y(new_n3866_));
  NAND2  g02864(.A(new_n3304_), .B(new_n3299_), .Y(new_n3867_));
  OAI21  g02865(.A0(new_n3866_), .A1(new_n3865_), .B0(new_n3867_), .Y(new_n3868_));
  NOR2   g02866(.A(\A[629] ), .B(new_n3309_), .Y(new_n3869_));
  OAI21  g02867(.A0(new_n3307_), .A1(\A[628] ), .B0(\A[630] ), .Y(new_n3870_));
  NAND2  g02868(.A(new_n3311_), .B(new_n3306_), .Y(new_n3871_));
  OAI21  g02869(.A0(new_n3870_), .A1(new_n3869_), .B0(new_n3871_), .Y(new_n3872_));
  NAND2  g02870(.A(new_n3311_), .B(\A[630] ), .Y(new_n3873_));
  OAI21  g02871(.A0(new_n3307_), .A1(new_n3309_), .B0(new_n3873_), .Y(new_n3874_));
  NAND2  g02872(.A(new_n3304_), .B(\A[627] ), .Y(new_n3875_));
  OAI21  g02873(.A0(new_n3300_), .A1(new_n3302_), .B0(new_n3875_), .Y(new_n3876_));
  NAND4  g02874(.A(new_n3876_), .B(new_n3874_), .C(new_n3872_), .D(new_n3868_), .Y(new_n3877_));
  NAND4  g02875(.A(new_n3858_), .B(new_n3847_), .C(new_n3855_), .D(new_n3852_), .Y(new_n3878_));
  NAND4  g02876(.A(new_n3878_), .B(new_n3844_), .C(new_n3877_), .D(new_n3864_), .Y(new_n3879_));
  XOR2   g02877(.A(new_n3316_), .B(new_n3874_), .Y(new_n3880_));
  NAND2  g02878(.A(new_n3872_), .B(new_n3868_), .Y(new_n3881_));
  NAND2  g02879(.A(new_n3876_), .B(new_n3874_), .Y(new_n3882_));
  OAI21  g02880(.A0(new_n3881_), .A1(new_n3880_), .B0(new_n3882_), .Y(new_n3883_));
  NOR2   g02881(.A(new_n3312_), .B(new_n3305_), .Y(new_n3884_));
  XOR2   g02882(.A(new_n3884_), .B(new_n3880_), .Y(new_n3885_));
  AOI21  g02883(.A0(new_n3883_), .A1(new_n3864_), .B0(new_n3885_), .Y(new_n3886_));
  XOR2   g02884(.A(new_n3886_), .B(new_n3879_), .Y(new_n3887_));
  NOR2   g02885(.A(new_n3887_), .B(new_n3863_), .Y(new_n3888_));
  XOR2   g02886(.A(new_n3312_), .B(new_n3868_), .Y(new_n3889_));
  NOR4   g02887(.A(new_n3316_), .B(new_n3314_), .C(new_n3312_), .D(new_n3305_), .Y(new_n3890_));
  XOR2   g02888(.A(new_n3331_), .B(new_n3852_), .Y(new_n3891_));
  NOR4   g02889(.A(new_n3335_), .B(new_n3333_), .C(new_n3331_), .D(new_n3324_), .Y(new_n3892_));
  NOR4   g02890(.A(new_n3892_), .B(new_n3891_), .C(new_n3890_), .D(new_n3889_), .Y(new_n3893_));
  XOR2   g02891(.A(new_n3316_), .B(new_n3314_), .Y(new_n3894_));
  XOR2   g02892(.A(new_n3884_), .B(new_n3894_), .Y(new_n3895_));
  NAND4  g02893(.A(new_n3844_), .B(new_n3877_), .C(new_n3895_), .D(new_n3864_), .Y(new_n3896_));
  NOR2   g02894(.A(new_n3316_), .B(new_n3314_), .Y(new_n3897_));
  AOI21  g02895(.A0(new_n3884_), .A1(new_n3894_), .B0(new_n3897_), .Y(new_n3898_));
  OAI21  g02896(.A0(new_n3898_), .A1(new_n3889_), .B0(new_n3878_), .Y(new_n3899_));
  OAI22  g02897(.A0(new_n3899_), .A1(new_n3896_), .B0(new_n3886_), .B1(new_n3893_), .Y(new_n3900_));
  NAND2  g02898(.A(new_n3376_), .B(new_n3337_), .Y(new_n3901_));
  AOI211 g02899(.A0(new_n3900_), .A1(new_n3863_), .B(new_n3901_), .C(new_n3888_), .Y(new_n3902_));
  XOR2   g02900(.A(new_n3335_), .B(new_n3333_), .Y(new_n3903_));
  NOR2   g02901(.A(new_n3335_), .B(new_n3333_), .Y(new_n3904_));
  AOI21  g02902(.A0(new_n3861_), .A1(new_n3903_), .B0(new_n3904_), .Y(new_n3905_));
  XOR2   g02903(.A(new_n3861_), .B(new_n3903_), .Y(new_n3906_));
  OAI21  g02904(.A0(new_n3905_), .A1(new_n3891_), .B0(new_n3906_), .Y(new_n3907_));
  XOR2   g02905(.A(new_n3886_), .B(new_n3893_), .Y(new_n3908_));
  NAND2  g02906(.A(new_n3908_), .B(new_n3907_), .Y(new_n3909_));
  NAND2  g02907(.A(new_n3900_), .B(new_n3863_), .Y(new_n3910_));
  INV    g02908(.A(new_n3901_), .Y(new_n3911_));
  AOI21  g02909(.A0(new_n3910_), .A1(new_n3909_), .B0(new_n3911_), .Y(new_n3912_));
  XOR2   g02910(.A(new_n3370_), .B(new_n3363_), .Y(new_n3913_));
  XOR2   g02911(.A(new_n3374_), .B(new_n3372_), .Y(new_n3914_));
  NOR2   g02912(.A(new_n3370_), .B(new_n3363_), .Y(new_n3915_));
  NAND2  g02913(.A(new_n3915_), .B(new_n3914_), .Y(new_n3916_));
  OAI21  g02914(.A0(new_n3374_), .A1(new_n3372_), .B0(new_n3916_), .Y(new_n3917_));
  INV    g02915(.A(new_n3369_), .Y(new_n3918_));
  NAND2  g02916(.A(\A[611] ), .B(\A[610] ), .Y(new_n3919_));
  OAI21  g02917(.A0(new_n3918_), .A1(new_n3364_), .B0(new_n3919_), .Y(new_n3920_));
  XOR2   g02918(.A(new_n3374_), .B(new_n3920_), .Y(new_n3921_));
  XOR2   g02919(.A(new_n3915_), .B(new_n3921_), .Y(new_n3922_));
  AOI21  g02920(.A0(new_n3917_), .A1(new_n3913_), .B0(new_n3922_), .Y(new_n3923_));
  XOR2   g02921(.A(new_n3351_), .B(new_n3344_), .Y(new_n3924_));
  NOR2   g02922(.A(\A[614] ), .B(new_n3341_), .Y(new_n3925_));
  OAI21  g02923(.A0(new_n3339_), .A1(\A[613] ), .B0(\A[615] ), .Y(new_n3926_));
  NAND2  g02924(.A(new_n3343_), .B(new_n3338_), .Y(new_n3927_));
  OAI21  g02925(.A0(new_n3926_), .A1(new_n3925_), .B0(new_n3927_), .Y(new_n3928_));
  NOR2   g02926(.A(\A[617] ), .B(new_n3348_), .Y(new_n3929_));
  OAI21  g02927(.A0(new_n3346_), .A1(\A[616] ), .B0(\A[618] ), .Y(new_n3930_));
  NAND2  g02928(.A(new_n3350_), .B(new_n3345_), .Y(new_n3931_));
  OAI21  g02929(.A0(new_n3930_), .A1(new_n3929_), .B0(new_n3931_), .Y(new_n3932_));
  NAND2  g02930(.A(new_n3350_), .B(\A[618] ), .Y(new_n3933_));
  OAI21  g02931(.A0(new_n3346_), .A1(new_n3348_), .B0(new_n3933_), .Y(new_n3934_));
  NAND2  g02932(.A(new_n3343_), .B(\A[615] ), .Y(new_n3935_));
  OAI21  g02933(.A0(new_n3339_), .A1(new_n3341_), .B0(new_n3935_), .Y(new_n3936_));
  NAND4  g02934(.A(new_n3936_), .B(new_n3934_), .C(new_n3932_), .D(new_n3928_), .Y(new_n3937_));
  INV    g02935(.A(new_n3362_), .Y(new_n3938_));
  NOR2   g02936(.A(new_n3938_), .B(new_n3357_), .Y(new_n3939_));
  OAI211 g02937(.A0(new_n3939_), .A1(new_n3373_), .B0(new_n3915_), .B1(new_n3920_), .Y(new_n3940_));
  NAND4  g02938(.A(new_n3940_), .B(new_n3913_), .C(new_n3937_), .D(new_n3924_), .Y(new_n3941_));
  XOR2   g02939(.A(new_n3355_), .B(new_n3934_), .Y(new_n3942_));
  NAND2  g02940(.A(new_n3932_), .B(new_n3928_), .Y(new_n3943_));
  NAND2  g02941(.A(new_n3936_), .B(new_n3934_), .Y(new_n3944_));
  OAI21  g02942(.A0(new_n3943_), .A1(new_n3942_), .B0(new_n3944_), .Y(new_n3945_));
  NOR2   g02943(.A(new_n3351_), .B(new_n3344_), .Y(new_n3946_));
  XOR2   g02944(.A(new_n3946_), .B(new_n3942_), .Y(new_n3947_));
  AOI21  g02945(.A0(new_n3945_), .A1(new_n3924_), .B0(new_n3947_), .Y(new_n3948_));
  XOR2   g02946(.A(new_n3948_), .B(new_n3941_), .Y(new_n3949_));
  NOR2   g02947(.A(new_n3949_), .B(new_n3923_), .Y(new_n3950_));
  NAND2  g02948(.A(new_n3361_), .B(new_n3359_), .Y(new_n3951_));
  OAI21  g02949(.A0(new_n3938_), .A1(\A[609] ), .B0(new_n3951_), .Y(new_n3952_));
  XOR2   g02950(.A(new_n3370_), .B(new_n3952_), .Y(new_n3953_));
  NOR2   g02951(.A(new_n3374_), .B(new_n3372_), .Y(new_n3954_));
  AOI21  g02952(.A0(new_n3915_), .A1(new_n3914_), .B0(new_n3954_), .Y(new_n3955_));
  XOR2   g02953(.A(new_n3915_), .B(new_n3914_), .Y(new_n3956_));
  OAI21  g02954(.A0(new_n3955_), .A1(new_n3953_), .B0(new_n3956_), .Y(new_n3957_));
  XOR2   g02955(.A(new_n3351_), .B(new_n3928_), .Y(new_n3958_));
  XOR2   g02956(.A(new_n3355_), .B(new_n3353_), .Y(new_n3959_));
  NOR2   g02957(.A(new_n3355_), .B(new_n3353_), .Y(new_n3960_));
  AOI21  g02958(.A0(new_n3946_), .A1(new_n3959_), .B0(new_n3960_), .Y(new_n3961_));
  XOR2   g02959(.A(new_n3946_), .B(new_n3959_), .Y(new_n3962_));
  OAI21  g02960(.A0(new_n3961_), .A1(new_n3958_), .B0(new_n3962_), .Y(new_n3963_));
  NAND2  g02961(.A(new_n3963_), .B(new_n3941_), .Y(new_n3964_));
  NOR4   g02962(.A(new_n3953_), .B(new_n3947_), .C(new_n3945_), .D(new_n3958_), .Y(new_n3965_));
  OAI211 g02963(.A0(new_n3961_), .A1(new_n3958_), .B0(new_n3965_), .B1(new_n3940_), .Y(new_n3966_));
  AOI21  g02964(.A0(new_n3966_), .A1(new_n3964_), .B0(new_n3957_), .Y(new_n3967_));
  NOR2   g02965(.A(new_n3967_), .B(new_n3950_), .Y(new_n3968_));
  OAI21  g02966(.A0(new_n3912_), .A1(new_n3902_), .B0(new_n3968_), .Y(new_n3969_));
  AOI211 g02967(.A0(new_n3900_), .A1(new_n3863_), .B(new_n3911_), .C(new_n3888_), .Y(new_n3970_));
  AOI21  g02968(.A0(new_n3910_), .A1(new_n3909_), .B0(new_n3901_), .Y(new_n3971_));
  OAI22  g02969(.A0(new_n3971_), .A1(new_n3970_), .B0(new_n3967_), .B1(new_n3950_), .Y(new_n3972_));
  NAND2  g02970(.A(new_n3972_), .B(new_n3969_), .Y(new_n3973_));
  XOR2   g02971(.A(new_n3289_), .B(new_n3282_), .Y(new_n3974_));
  XOR2   g02972(.A(new_n3293_), .B(new_n3291_), .Y(new_n3975_));
  NOR2   g02973(.A(new_n3289_), .B(new_n3282_), .Y(new_n3976_));
  NAND2  g02974(.A(new_n3976_), .B(new_n3975_), .Y(new_n3977_));
  OAI21  g02975(.A0(new_n3293_), .A1(new_n3291_), .B0(new_n3977_), .Y(new_n3978_));
  INV    g02976(.A(new_n3288_), .Y(new_n3979_));
  NAND2  g02977(.A(\A[635] ), .B(\A[634] ), .Y(new_n3980_));
  OAI21  g02978(.A0(new_n3979_), .A1(new_n3283_), .B0(new_n3980_), .Y(new_n3981_));
  XOR2   g02979(.A(new_n3293_), .B(new_n3981_), .Y(new_n3982_));
  XOR2   g02980(.A(new_n3976_), .B(new_n3982_), .Y(new_n3983_));
  AOI21  g02981(.A0(new_n3978_), .A1(new_n3974_), .B0(new_n3983_), .Y(new_n3984_));
  XOR2   g02982(.A(new_n3270_), .B(new_n3263_), .Y(new_n3985_));
  NOR2   g02983(.A(\A[638] ), .B(new_n3260_), .Y(new_n3986_));
  OAI21  g02984(.A0(new_n3258_), .A1(\A[637] ), .B0(\A[639] ), .Y(new_n3987_));
  NAND2  g02985(.A(new_n3262_), .B(new_n3257_), .Y(new_n3988_));
  OAI21  g02986(.A0(new_n3987_), .A1(new_n3986_), .B0(new_n3988_), .Y(new_n3989_));
  NOR2   g02987(.A(\A[641] ), .B(new_n3267_), .Y(new_n3990_));
  OAI21  g02988(.A0(new_n3265_), .A1(\A[640] ), .B0(\A[642] ), .Y(new_n3991_));
  NAND2  g02989(.A(new_n3269_), .B(new_n3264_), .Y(new_n3992_));
  OAI21  g02990(.A0(new_n3991_), .A1(new_n3990_), .B0(new_n3992_), .Y(new_n3993_));
  NAND2  g02991(.A(new_n3269_), .B(\A[642] ), .Y(new_n3994_));
  OAI21  g02992(.A0(new_n3265_), .A1(new_n3267_), .B0(new_n3994_), .Y(new_n3995_));
  NAND2  g02993(.A(new_n3262_), .B(\A[639] ), .Y(new_n3996_));
  OAI21  g02994(.A0(new_n3258_), .A1(new_n3260_), .B0(new_n3996_), .Y(new_n3997_));
  NAND4  g02995(.A(new_n3997_), .B(new_n3995_), .C(new_n3993_), .D(new_n3989_), .Y(new_n3998_));
  INV    g02996(.A(new_n3281_), .Y(new_n3999_));
  NOR2   g02997(.A(new_n3999_), .B(new_n3276_), .Y(new_n4000_));
  OAI211 g02998(.A0(new_n4000_), .A1(new_n3292_), .B0(new_n3976_), .B1(new_n3981_), .Y(new_n4001_));
  NAND4  g02999(.A(new_n4001_), .B(new_n3974_), .C(new_n3998_), .D(new_n3985_), .Y(new_n4002_));
  XOR2   g03000(.A(new_n3274_), .B(new_n3995_), .Y(new_n4003_));
  NAND2  g03001(.A(new_n3993_), .B(new_n3989_), .Y(new_n4004_));
  NAND2  g03002(.A(new_n3997_), .B(new_n3995_), .Y(new_n4005_));
  OAI21  g03003(.A0(new_n4004_), .A1(new_n4003_), .B0(new_n4005_), .Y(new_n4006_));
  NOR2   g03004(.A(new_n3270_), .B(new_n3263_), .Y(new_n4007_));
  XOR2   g03005(.A(new_n4007_), .B(new_n4003_), .Y(new_n4008_));
  AOI21  g03006(.A0(new_n4006_), .A1(new_n3985_), .B0(new_n4008_), .Y(new_n4009_));
  XOR2   g03007(.A(new_n4009_), .B(new_n4002_), .Y(new_n4010_));
  NOR2   g03008(.A(new_n4010_), .B(new_n3984_), .Y(new_n4011_));
  NAND2  g03009(.A(new_n3280_), .B(new_n3278_), .Y(new_n4012_));
  OAI21  g03010(.A0(new_n3999_), .A1(\A[633] ), .B0(new_n4012_), .Y(new_n4013_));
  XOR2   g03011(.A(new_n3289_), .B(new_n4013_), .Y(new_n4014_));
  NOR2   g03012(.A(new_n3293_), .B(new_n3291_), .Y(new_n4015_));
  AOI21  g03013(.A0(new_n3976_), .A1(new_n3975_), .B0(new_n4015_), .Y(new_n4016_));
  XOR2   g03014(.A(new_n3976_), .B(new_n3975_), .Y(new_n4017_));
  OAI21  g03015(.A0(new_n4016_), .A1(new_n4014_), .B0(new_n4017_), .Y(new_n4018_));
  XOR2   g03016(.A(new_n3270_), .B(new_n3989_), .Y(new_n4019_));
  XOR2   g03017(.A(new_n3274_), .B(new_n3272_), .Y(new_n4020_));
  NOR2   g03018(.A(new_n3274_), .B(new_n3272_), .Y(new_n4021_));
  AOI21  g03019(.A0(new_n4007_), .A1(new_n4020_), .B0(new_n4021_), .Y(new_n4022_));
  XOR2   g03020(.A(new_n4007_), .B(new_n4020_), .Y(new_n4023_));
  OAI21  g03021(.A0(new_n4022_), .A1(new_n4019_), .B0(new_n4023_), .Y(new_n4024_));
  NAND2  g03022(.A(new_n4024_), .B(new_n4002_), .Y(new_n4025_));
  NOR4   g03023(.A(new_n4014_), .B(new_n4008_), .C(new_n4006_), .D(new_n4019_), .Y(new_n4026_));
  OAI211 g03024(.A0(new_n4022_), .A1(new_n4019_), .B0(new_n4026_), .B1(new_n4001_), .Y(new_n4027_));
  AOI21  g03025(.A0(new_n4027_), .A1(new_n4025_), .B0(new_n4018_), .Y(new_n4028_));
  NOR2   g03026(.A(new_n4028_), .B(new_n4011_), .Y(new_n4029_));
  NAND2  g03027(.A(new_n3295_), .B(new_n3256_), .Y(new_n4030_));
  INV    g03028(.A(new_n4030_), .Y(new_n4031_));
  NOR2   g03029(.A(\A[644] ), .B(new_n3239_), .Y(new_n4032_));
  OAI21  g03030(.A0(new_n3237_), .A1(\A[643] ), .B0(\A[645] ), .Y(new_n4033_));
  XOR2   g03031(.A(\A[644] ), .B(new_n3239_), .Y(new_n4034_));
  OAI22  g03032(.A0(new_n4034_), .A1(\A[645] ), .B0(new_n4033_), .B1(new_n4032_), .Y(new_n4035_));
  XOR2   g03033(.A(new_n3249_), .B(new_n4035_), .Y(new_n4036_));
  XOR2   g03034(.A(new_n3254_), .B(new_n3252_), .Y(new_n4037_));
  NOR2   g03035(.A(new_n3249_), .B(new_n3242_), .Y(new_n4038_));
  NOR2   g03036(.A(new_n3254_), .B(new_n3252_), .Y(new_n4039_));
  AOI21  g03037(.A0(new_n4038_), .A1(new_n4037_), .B0(new_n4039_), .Y(new_n4040_));
  XOR2   g03038(.A(new_n4038_), .B(new_n4037_), .Y(new_n4041_));
  OAI21  g03039(.A0(new_n4040_), .A1(new_n4036_), .B0(new_n4041_), .Y(new_n4042_));
  NOR2   g03040(.A(\A[650] ), .B(new_n3220_), .Y(new_n4043_));
  OAI21  g03041(.A0(new_n3218_), .A1(\A[649] ), .B0(\A[651] ), .Y(new_n4044_));
  NAND2  g03042(.A(new_n3222_), .B(new_n3217_), .Y(new_n4045_));
  OAI21  g03043(.A0(new_n4044_), .A1(new_n4043_), .B0(new_n4045_), .Y(new_n4046_));
  XOR2   g03044(.A(new_n3230_), .B(new_n4046_), .Y(new_n4047_));
  NOR4   g03045(.A(new_n3234_), .B(new_n3232_), .C(new_n3230_), .D(new_n3223_), .Y(new_n4048_));
  NOR4   g03046(.A(new_n3254_), .B(new_n3252_), .C(new_n3249_), .D(new_n3242_), .Y(new_n4049_));
  NOR4   g03047(.A(new_n4049_), .B(new_n4036_), .C(new_n4048_), .D(new_n4047_), .Y(new_n4050_));
  XOR2   g03048(.A(new_n3230_), .B(new_n3223_), .Y(new_n4051_));
  NAND2  g03049(.A(new_n3229_), .B(\A[654] ), .Y(new_n4052_));
  OAI21  g03050(.A0(new_n3225_), .A1(new_n3227_), .B0(new_n4052_), .Y(new_n4053_));
  XOR2   g03051(.A(new_n3234_), .B(new_n4053_), .Y(new_n4054_));
  NOR2   g03052(.A(\A[653] ), .B(new_n3227_), .Y(new_n4055_));
  OAI21  g03053(.A0(new_n3225_), .A1(\A[652] ), .B0(\A[654] ), .Y(new_n4056_));
  NAND2  g03054(.A(new_n3229_), .B(new_n3224_), .Y(new_n4057_));
  OAI21  g03055(.A0(new_n4056_), .A1(new_n4055_), .B0(new_n4057_), .Y(new_n4058_));
  NAND2  g03056(.A(new_n4058_), .B(new_n4046_), .Y(new_n4059_));
  NAND2  g03057(.A(new_n3222_), .B(\A[651] ), .Y(new_n4060_));
  OAI21  g03058(.A0(new_n3218_), .A1(new_n3220_), .B0(new_n4060_), .Y(new_n4061_));
  NAND2  g03059(.A(new_n4061_), .B(new_n4053_), .Y(new_n4062_));
  OAI21  g03060(.A0(new_n4059_), .A1(new_n4054_), .B0(new_n4062_), .Y(new_n4063_));
  NOR2   g03061(.A(new_n3230_), .B(new_n3223_), .Y(new_n4064_));
  XOR2   g03062(.A(new_n4064_), .B(new_n4054_), .Y(new_n4065_));
  AOI21  g03063(.A0(new_n4063_), .A1(new_n4051_), .B0(new_n4065_), .Y(new_n4066_));
  XOR2   g03064(.A(new_n4066_), .B(new_n4050_), .Y(new_n4067_));
  NAND2  g03065(.A(new_n4067_), .B(new_n4042_), .Y(new_n4068_));
  XOR2   g03066(.A(new_n3249_), .B(new_n3242_), .Y(new_n4069_));
  XOR2   g03067(.A(\A[647] ), .B(new_n3246_), .Y(new_n4070_));
  OAI21  g03068(.A0(new_n4070_), .A1(new_n3243_), .B0(new_n3250_), .Y(new_n4071_));
  XOR2   g03069(.A(new_n3254_), .B(new_n4071_), .Y(new_n4072_));
  NOR2   g03070(.A(\A[647] ), .B(new_n3246_), .Y(new_n4073_));
  OAI21  g03071(.A0(new_n3244_), .A1(\A[646] ), .B0(\A[648] ), .Y(new_n4074_));
  OAI22  g03072(.A0(new_n4070_), .A1(\A[648] ), .B0(new_n4074_), .B1(new_n4073_), .Y(new_n4075_));
  NAND2  g03073(.A(new_n4075_), .B(new_n4035_), .Y(new_n4076_));
  NAND2  g03074(.A(\A[644] ), .B(\A[643] ), .Y(new_n4077_));
  OAI21  g03075(.A0(new_n4034_), .A1(new_n3236_), .B0(new_n4077_), .Y(new_n4078_));
  NAND2  g03076(.A(new_n4078_), .B(new_n4071_), .Y(new_n4079_));
  OAI21  g03077(.A0(new_n4076_), .A1(new_n4072_), .B0(new_n4079_), .Y(new_n4080_));
  XOR2   g03078(.A(new_n4038_), .B(new_n4072_), .Y(new_n4081_));
  AOI21  g03079(.A0(new_n4080_), .A1(new_n4069_), .B0(new_n4081_), .Y(new_n4082_));
  XOR2   g03080(.A(new_n3234_), .B(new_n3232_), .Y(new_n4083_));
  XOR2   g03081(.A(new_n4064_), .B(new_n4083_), .Y(new_n4084_));
  NAND4  g03082(.A(new_n4061_), .B(new_n4053_), .C(new_n4058_), .D(new_n4046_), .Y(new_n4085_));
  NAND4  g03083(.A(new_n4069_), .B(new_n4085_), .C(new_n4084_), .D(new_n4051_), .Y(new_n4086_));
  NOR2   g03084(.A(new_n3234_), .B(new_n3232_), .Y(new_n4087_));
  AOI21  g03085(.A0(new_n4064_), .A1(new_n4083_), .B0(new_n4087_), .Y(new_n4088_));
  NAND4  g03086(.A(new_n4078_), .B(new_n4071_), .C(new_n4075_), .D(new_n4035_), .Y(new_n4089_));
  OAI21  g03087(.A0(new_n4088_), .A1(new_n4047_), .B0(new_n4089_), .Y(new_n4090_));
  OAI22  g03088(.A0(new_n4090_), .A1(new_n4086_), .B0(new_n4066_), .B1(new_n4050_), .Y(new_n4091_));
  NAND2  g03089(.A(new_n4091_), .B(new_n4082_), .Y(new_n4092_));
  NAND3  g03090(.A(new_n4031_), .B(new_n4092_), .C(new_n4068_), .Y(new_n4093_));
  NAND4  g03091(.A(new_n4089_), .B(new_n4069_), .C(new_n4085_), .D(new_n4051_), .Y(new_n4094_));
  XOR2   g03092(.A(new_n4066_), .B(new_n4094_), .Y(new_n4095_));
  NOR2   g03093(.A(new_n4095_), .B(new_n4082_), .Y(new_n4096_));
  AOI21  g03094(.A0(new_n4091_), .A1(new_n4082_), .B0(new_n4096_), .Y(new_n4097_));
  OAI21  g03095(.A0(new_n4097_), .A1(new_n4031_), .B0(new_n4093_), .Y(new_n4098_));
  NAND2  g03096(.A(new_n4098_), .B(new_n4029_), .Y(new_n4099_));
  AOI211 g03097(.A0(new_n4091_), .A1(new_n4082_), .B(new_n4031_), .C(new_n4096_), .Y(new_n4100_));
  AOI21  g03098(.A0(new_n4092_), .A1(new_n4068_), .B0(new_n4030_), .Y(new_n4101_));
  OAI22  g03099(.A0(new_n4101_), .A1(new_n4100_), .B0(new_n4028_), .B1(new_n4011_), .Y(new_n4102_));
  NOR2   g03100(.A(new_n3378_), .B(new_n3297_), .Y(new_n4103_));
  NAND3  g03101(.A(new_n4103_), .B(new_n4102_), .C(new_n4099_), .Y(new_n4104_));
  NAND2  g03102(.A(new_n4027_), .B(new_n4025_), .Y(new_n4105_));
  NAND2  g03103(.A(new_n4105_), .B(new_n3984_), .Y(new_n4106_));
  OAI21  g03104(.A0(new_n4010_), .A1(new_n3984_), .B0(new_n4106_), .Y(new_n4107_));
  NOR2   g03105(.A(new_n4066_), .B(new_n4050_), .Y(new_n4108_));
  NOR2   g03106(.A(new_n4090_), .B(new_n4086_), .Y(new_n4109_));
  NOR2   g03107(.A(new_n4109_), .B(new_n4108_), .Y(new_n4110_));
  NOR2   g03108(.A(new_n4110_), .B(new_n4042_), .Y(new_n4111_));
  OAI21  g03109(.A0(new_n4111_), .A1(new_n4096_), .B0(new_n4030_), .Y(new_n4112_));
  AOI21  g03110(.A0(new_n4112_), .A1(new_n4093_), .B0(new_n4107_), .Y(new_n4113_));
  NAND3  g03111(.A(new_n4030_), .B(new_n4092_), .C(new_n4068_), .Y(new_n4114_));
  OAI21  g03112(.A0(new_n4111_), .A1(new_n4096_), .B0(new_n4031_), .Y(new_n4115_));
  AOI21  g03113(.A0(new_n4115_), .A1(new_n4114_), .B0(new_n4029_), .Y(new_n4116_));
  INV    g03114(.A(new_n4103_), .Y(new_n4117_));
  OAI21  g03115(.A0(new_n4116_), .A1(new_n4113_), .B0(new_n4117_), .Y(new_n4118_));
  AOI21  g03116(.A0(new_n4118_), .A1(new_n4104_), .B0(new_n3973_), .Y(new_n4119_));
  NOR2   g03117(.A(new_n3912_), .B(new_n3902_), .Y(new_n4120_));
  NAND2  g03118(.A(new_n3966_), .B(new_n3964_), .Y(new_n4121_));
  NAND2  g03119(.A(new_n4121_), .B(new_n3923_), .Y(new_n4122_));
  OAI21  g03120(.A0(new_n3949_), .A1(new_n3923_), .B0(new_n4122_), .Y(new_n4123_));
  NOR2   g03121(.A(new_n4123_), .B(new_n4120_), .Y(new_n4124_));
  NAND3  g03122(.A(new_n3901_), .B(new_n3910_), .C(new_n3909_), .Y(new_n4125_));
  NAND2  g03123(.A(new_n3910_), .B(new_n3909_), .Y(new_n4126_));
  NAND2  g03124(.A(new_n4126_), .B(new_n3911_), .Y(new_n4127_));
  AOI21  g03125(.A0(new_n4127_), .A1(new_n4125_), .B0(new_n3968_), .Y(new_n4128_));
  NOR2   g03126(.A(new_n4128_), .B(new_n4124_), .Y(new_n4129_));
  OAI21  g03127(.A0(new_n4097_), .A1(new_n4030_), .B0(new_n4114_), .Y(new_n4130_));
  AOI21  g03128(.A0(new_n4130_), .A1(new_n4107_), .B0(new_n4103_), .Y(new_n4131_));
  NAND2  g03129(.A(new_n4131_), .B(new_n4099_), .Y(new_n4132_));
  OAI21  g03130(.A0(new_n4116_), .A1(new_n4113_), .B0(new_n4103_), .Y(new_n4133_));
  AOI21  g03131(.A0(new_n4133_), .A1(new_n4132_), .B0(new_n4129_), .Y(new_n4134_));
  NOR2   g03132(.A(new_n3542_), .B(new_n3379_), .Y(new_n4135_));
  INV    g03133(.A(new_n4135_), .Y(new_n4136_));
  NOR3   g03134(.A(new_n4136_), .B(new_n4134_), .C(new_n4119_), .Y(new_n4137_));
  NOR3   g03135(.A(new_n4117_), .B(new_n4116_), .C(new_n4113_), .Y(new_n4138_));
  AOI21  g03136(.A0(new_n4102_), .A1(new_n4099_), .B0(new_n4103_), .Y(new_n4139_));
  OAI21  g03137(.A0(new_n4139_), .A1(new_n4138_), .B0(new_n4129_), .Y(new_n4140_));
  NOR3   g03138(.A(new_n4103_), .B(new_n4116_), .C(new_n4113_), .Y(new_n4141_));
  AOI21  g03139(.A0(new_n4102_), .A1(new_n4099_), .B0(new_n4117_), .Y(new_n4142_));
  OAI21  g03140(.A0(new_n4142_), .A1(new_n4141_), .B0(new_n3973_), .Y(new_n4143_));
  AOI21  g03141(.A0(new_n4143_), .A1(new_n4140_), .B0(new_n4135_), .Y(new_n4144_));
  OAI21  g03142(.A0(new_n4144_), .A1(new_n4137_), .B0(new_n3843_), .Y(new_n4145_));
  NOR2   g03143(.A(new_n3692_), .B(new_n3682_), .Y(new_n4146_));
  NAND2  g03144(.A(new_n3838_), .B(new_n3614_), .Y(new_n4147_));
  AOI21  g03145(.A0(new_n4147_), .A1(new_n3836_), .B0(new_n3691_), .Y(new_n4148_));
  OAI21  g03146(.A0(new_n4148_), .A1(new_n4146_), .B0(new_n3833_), .Y(new_n4149_));
  NOR3   g03147(.A(new_n3691_), .B(new_n3693_), .C(new_n3682_), .Y(new_n4150_));
  AOI21  g03148(.A0(new_n4147_), .A1(new_n3836_), .B0(new_n3694_), .Y(new_n4151_));
  NOR2   g03149(.A(new_n4151_), .B(new_n4150_), .Y(new_n4152_));
  OAI21  g03150(.A0(new_n4152_), .A1(new_n3833_), .B0(new_n4149_), .Y(new_n4153_));
  NOR3   g03151(.A(new_n4135_), .B(new_n4134_), .C(new_n4119_), .Y(new_n4154_));
  AOI21  g03152(.A0(new_n4143_), .A1(new_n4140_), .B0(new_n4136_), .Y(new_n4155_));
  OAI21  g03153(.A0(new_n4155_), .A1(new_n4154_), .B0(new_n4153_), .Y(new_n4156_));
  NOR2   g03154(.A(new_n3543_), .B(new_n3215_), .Y(new_n4157_));
  NAND3  g03155(.A(new_n4157_), .B(new_n4156_), .C(new_n4145_), .Y(new_n4158_));
  NAND3  g03156(.A(new_n4135_), .B(new_n4143_), .C(new_n4140_), .Y(new_n4159_));
  OAI21  g03157(.A0(new_n4134_), .A1(new_n4119_), .B0(new_n4136_), .Y(new_n4160_));
  AOI21  g03158(.A0(new_n4160_), .A1(new_n4159_), .B0(new_n4153_), .Y(new_n4161_));
  NAND3  g03159(.A(new_n4136_), .B(new_n4143_), .C(new_n4140_), .Y(new_n4162_));
  OAI21  g03160(.A0(new_n4134_), .A1(new_n4119_), .B0(new_n4135_), .Y(new_n4163_));
  AOI21  g03161(.A0(new_n4163_), .A1(new_n4162_), .B0(new_n3843_), .Y(new_n4164_));
  INV    g03162(.A(new_n4157_), .Y(new_n4165_));
  OAI21  g03163(.A0(new_n4164_), .A1(new_n4161_), .B0(new_n4165_), .Y(new_n4166_));
  XOR2   g03164(.A(new_n3166_), .B(new_n3159_), .Y(new_n4167_));
  XOR2   g03165(.A(\A[527] ), .B(new_n3163_), .Y(new_n4168_));
  NAND2  g03166(.A(\A[527] ), .B(\A[526] ), .Y(new_n4169_));
  OAI21  g03167(.A0(new_n4168_), .A1(new_n3160_), .B0(new_n4169_), .Y(new_n4170_));
  XOR2   g03168(.A(new_n3170_), .B(new_n4170_), .Y(new_n4171_));
  NOR2   g03169(.A(\A[524] ), .B(new_n3156_), .Y(new_n4172_));
  OAI21  g03170(.A0(new_n3154_), .A1(\A[523] ), .B0(\A[525] ), .Y(new_n4173_));
  XOR2   g03171(.A(\A[524] ), .B(new_n3156_), .Y(new_n4174_));
  OAI22  g03172(.A0(new_n4174_), .A1(\A[525] ), .B0(new_n4173_), .B1(new_n4172_), .Y(new_n4175_));
  NOR2   g03173(.A(\A[527] ), .B(new_n3163_), .Y(new_n4176_));
  OAI21  g03174(.A0(new_n3161_), .A1(\A[526] ), .B0(\A[528] ), .Y(new_n4177_));
  OAI22  g03175(.A0(new_n4168_), .A1(\A[528] ), .B0(new_n4177_), .B1(new_n4176_), .Y(new_n4178_));
  NAND2  g03176(.A(new_n4178_), .B(new_n4175_), .Y(new_n4179_));
  NAND2  g03177(.A(\A[524] ), .B(\A[523] ), .Y(new_n4180_));
  OAI21  g03178(.A0(new_n4174_), .A1(new_n3153_), .B0(new_n4180_), .Y(new_n4181_));
  NAND2  g03179(.A(new_n4181_), .B(new_n4170_), .Y(new_n4182_));
  OAI21  g03180(.A0(new_n4179_), .A1(new_n4171_), .B0(new_n4182_), .Y(new_n4183_));
  NOR2   g03181(.A(new_n3166_), .B(new_n3159_), .Y(new_n4184_));
  XOR2   g03182(.A(new_n4184_), .B(new_n4171_), .Y(new_n4185_));
  AOI21  g03183(.A0(new_n4183_), .A1(new_n4167_), .B0(new_n4185_), .Y(new_n4186_));
  XOR2   g03184(.A(new_n3147_), .B(new_n3140_), .Y(new_n4187_));
  NOR2   g03185(.A(\A[530] ), .B(new_n3137_), .Y(new_n4188_));
  OAI21  g03186(.A0(new_n3135_), .A1(\A[529] ), .B0(\A[531] ), .Y(new_n4189_));
  NAND2  g03187(.A(new_n3139_), .B(new_n3134_), .Y(new_n4190_));
  OAI21  g03188(.A0(new_n4189_), .A1(new_n4188_), .B0(new_n4190_), .Y(new_n4191_));
  NOR2   g03189(.A(\A[533] ), .B(new_n3144_), .Y(new_n4192_));
  OAI21  g03190(.A0(new_n3142_), .A1(\A[532] ), .B0(\A[534] ), .Y(new_n4193_));
  NAND2  g03191(.A(new_n3146_), .B(new_n3141_), .Y(new_n4194_));
  OAI21  g03192(.A0(new_n4193_), .A1(new_n4192_), .B0(new_n4194_), .Y(new_n4195_));
  NAND2  g03193(.A(new_n3146_), .B(\A[534] ), .Y(new_n4196_));
  OAI21  g03194(.A0(new_n3142_), .A1(new_n3144_), .B0(new_n4196_), .Y(new_n4197_));
  NAND2  g03195(.A(new_n3139_), .B(\A[531] ), .Y(new_n4198_));
  OAI21  g03196(.A0(new_n3135_), .A1(new_n3137_), .B0(new_n4198_), .Y(new_n4199_));
  NAND4  g03197(.A(new_n4199_), .B(new_n4197_), .C(new_n4195_), .D(new_n4191_), .Y(new_n4200_));
  NAND4  g03198(.A(new_n4181_), .B(new_n4170_), .C(new_n4178_), .D(new_n4175_), .Y(new_n4201_));
  NAND4  g03199(.A(new_n4201_), .B(new_n4167_), .C(new_n4200_), .D(new_n4187_), .Y(new_n4202_));
  XOR2   g03200(.A(new_n3151_), .B(new_n4197_), .Y(new_n4203_));
  NAND2  g03201(.A(new_n4195_), .B(new_n4191_), .Y(new_n4204_));
  NAND2  g03202(.A(new_n4199_), .B(new_n4197_), .Y(new_n4205_));
  OAI21  g03203(.A0(new_n4204_), .A1(new_n4203_), .B0(new_n4205_), .Y(new_n4206_));
  NOR2   g03204(.A(new_n3147_), .B(new_n3140_), .Y(new_n4207_));
  XOR2   g03205(.A(new_n4207_), .B(new_n4203_), .Y(new_n4208_));
  AOI21  g03206(.A0(new_n4206_), .A1(new_n4187_), .B0(new_n4208_), .Y(new_n4209_));
  XOR2   g03207(.A(new_n4209_), .B(new_n4202_), .Y(new_n4210_));
  NOR2   g03208(.A(new_n4210_), .B(new_n4186_), .Y(new_n4211_));
  XOR2   g03209(.A(new_n3147_), .B(new_n4191_), .Y(new_n4212_));
  NOR4   g03210(.A(new_n3151_), .B(new_n3149_), .C(new_n3147_), .D(new_n3140_), .Y(new_n4213_));
  XOR2   g03211(.A(new_n3166_), .B(new_n4175_), .Y(new_n4214_));
  NOR4   g03212(.A(new_n3170_), .B(new_n3168_), .C(new_n3166_), .D(new_n3159_), .Y(new_n4215_));
  NOR4   g03213(.A(new_n4215_), .B(new_n4214_), .C(new_n4213_), .D(new_n4212_), .Y(new_n4216_));
  XOR2   g03214(.A(new_n3151_), .B(new_n3149_), .Y(new_n4217_));
  XOR2   g03215(.A(new_n4207_), .B(new_n4217_), .Y(new_n4218_));
  NAND4  g03216(.A(new_n4167_), .B(new_n4200_), .C(new_n4218_), .D(new_n4187_), .Y(new_n4219_));
  NOR2   g03217(.A(new_n3151_), .B(new_n3149_), .Y(new_n4220_));
  AOI21  g03218(.A0(new_n4207_), .A1(new_n4217_), .B0(new_n4220_), .Y(new_n4221_));
  OAI21  g03219(.A0(new_n4221_), .A1(new_n4212_), .B0(new_n4201_), .Y(new_n4222_));
  OAI22  g03220(.A0(new_n4222_), .A1(new_n4219_), .B0(new_n4209_), .B1(new_n4216_), .Y(new_n4223_));
  NAND2  g03221(.A(new_n3211_), .B(new_n3172_), .Y(new_n4224_));
  AOI211 g03222(.A0(new_n4223_), .A1(new_n4186_), .B(new_n4224_), .C(new_n4211_), .Y(new_n4225_));
  XOR2   g03223(.A(new_n3170_), .B(new_n3168_), .Y(new_n4226_));
  NOR2   g03224(.A(new_n3170_), .B(new_n3168_), .Y(new_n4227_));
  AOI21  g03225(.A0(new_n4184_), .A1(new_n4226_), .B0(new_n4227_), .Y(new_n4228_));
  XOR2   g03226(.A(new_n4184_), .B(new_n4226_), .Y(new_n4229_));
  OAI21  g03227(.A0(new_n4228_), .A1(new_n4214_), .B0(new_n4229_), .Y(new_n4230_));
  XOR2   g03228(.A(new_n4209_), .B(new_n4216_), .Y(new_n4231_));
  NAND2  g03229(.A(new_n4231_), .B(new_n4230_), .Y(new_n4232_));
  NAND2  g03230(.A(new_n4223_), .B(new_n4186_), .Y(new_n4233_));
  INV    g03231(.A(new_n4224_), .Y(new_n4234_));
  AOI21  g03232(.A0(new_n4233_), .A1(new_n4232_), .B0(new_n4234_), .Y(new_n4235_));
  XOR2   g03233(.A(new_n3205_), .B(new_n3198_), .Y(new_n4236_));
  XOR2   g03234(.A(new_n3209_), .B(new_n3207_), .Y(new_n4237_));
  NOR2   g03235(.A(new_n3205_), .B(new_n3198_), .Y(new_n4238_));
  NAND2  g03236(.A(new_n4238_), .B(new_n4237_), .Y(new_n4239_));
  OAI21  g03237(.A0(new_n3209_), .A1(new_n3207_), .B0(new_n4239_), .Y(new_n4240_));
  INV    g03238(.A(new_n3204_), .Y(new_n4241_));
  NAND2  g03239(.A(\A[515] ), .B(\A[514] ), .Y(new_n4242_));
  OAI21  g03240(.A0(new_n4241_), .A1(new_n3199_), .B0(new_n4242_), .Y(new_n4243_));
  XOR2   g03241(.A(new_n3209_), .B(new_n4243_), .Y(new_n4244_));
  XOR2   g03242(.A(new_n4238_), .B(new_n4244_), .Y(new_n4245_));
  AOI21  g03243(.A0(new_n4240_), .A1(new_n4236_), .B0(new_n4245_), .Y(new_n4246_));
  XOR2   g03244(.A(new_n3186_), .B(new_n3179_), .Y(new_n4247_));
  NOR2   g03245(.A(\A[518] ), .B(new_n3176_), .Y(new_n4248_));
  OAI21  g03246(.A0(new_n3174_), .A1(\A[517] ), .B0(\A[519] ), .Y(new_n4249_));
  NAND2  g03247(.A(new_n3178_), .B(new_n3173_), .Y(new_n4250_));
  OAI21  g03248(.A0(new_n4249_), .A1(new_n4248_), .B0(new_n4250_), .Y(new_n4251_));
  NOR2   g03249(.A(\A[521] ), .B(new_n3183_), .Y(new_n4252_));
  OAI21  g03250(.A0(new_n3181_), .A1(\A[520] ), .B0(\A[522] ), .Y(new_n4253_));
  NAND2  g03251(.A(new_n3185_), .B(new_n3180_), .Y(new_n4254_));
  OAI21  g03252(.A0(new_n4253_), .A1(new_n4252_), .B0(new_n4254_), .Y(new_n4255_));
  NAND2  g03253(.A(new_n3185_), .B(\A[522] ), .Y(new_n4256_));
  OAI21  g03254(.A0(new_n3181_), .A1(new_n3183_), .B0(new_n4256_), .Y(new_n4257_));
  NAND2  g03255(.A(new_n3178_), .B(\A[519] ), .Y(new_n4258_));
  OAI21  g03256(.A0(new_n3174_), .A1(new_n3176_), .B0(new_n4258_), .Y(new_n4259_));
  NAND4  g03257(.A(new_n4259_), .B(new_n4257_), .C(new_n4255_), .D(new_n4251_), .Y(new_n4260_));
  INV    g03258(.A(new_n3197_), .Y(new_n4261_));
  NOR2   g03259(.A(new_n4261_), .B(new_n3192_), .Y(new_n4262_));
  OAI211 g03260(.A0(new_n4262_), .A1(new_n3208_), .B0(new_n4238_), .B1(new_n4243_), .Y(new_n4263_));
  NAND4  g03261(.A(new_n4263_), .B(new_n4236_), .C(new_n4260_), .D(new_n4247_), .Y(new_n4264_));
  XOR2   g03262(.A(new_n3190_), .B(new_n4257_), .Y(new_n4265_));
  NAND2  g03263(.A(new_n4255_), .B(new_n4251_), .Y(new_n4266_));
  NAND2  g03264(.A(new_n4259_), .B(new_n4257_), .Y(new_n4267_));
  OAI21  g03265(.A0(new_n4266_), .A1(new_n4265_), .B0(new_n4267_), .Y(new_n4268_));
  NOR2   g03266(.A(new_n3186_), .B(new_n3179_), .Y(new_n4269_));
  XOR2   g03267(.A(new_n4269_), .B(new_n4265_), .Y(new_n4270_));
  AOI21  g03268(.A0(new_n4268_), .A1(new_n4247_), .B0(new_n4270_), .Y(new_n4271_));
  XOR2   g03269(.A(new_n4271_), .B(new_n4264_), .Y(new_n4272_));
  NOR2   g03270(.A(new_n4272_), .B(new_n4246_), .Y(new_n4273_));
  NAND2  g03271(.A(new_n3196_), .B(new_n3194_), .Y(new_n4274_));
  OAI21  g03272(.A0(new_n4261_), .A1(\A[513] ), .B0(new_n4274_), .Y(new_n4275_));
  XOR2   g03273(.A(new_n3205_), .B(new_n4275_), .Y(new_n4276_));
  NOR2   g03274(.A(new_n3209_), .B(new_n3207_), .Y(new_n4277_));
  AOI21  g03275(.A0(new_n4238_), .A1(new_n4237_), .B0(new_n4277_), .Y(new_n4278_));
  XOR2   g03276(.A(new_n4238_), .B(new_n4237_), .Y(new_n4279_));
  OAI21  g03277(.A0(new_n4278_), .A1(new_n4276_), .B0(new_n4279_), .Y(new_n4280_));
  XOR2   g03278(.A(new_n3186_), .B(new_n4251_), .Y(new_n4281_));
  XOR2   g03279(.A(new_n3190_), .B(new_n3188_), .Y(new_n4282_));
  NOR2   g03280(.A(new_n3190_), .B(new_n3188_), .Y(new_n4283_));
  AOI21  g03281(.A0(new_n4269_), .A1(new_n4282_), .B0(new_n4283_), .Y(new_n4284_));
  XOR2   g03282(.A(new_n4269_), .B(new_n4282_), .Y(new_n4285_));
  OAI21  g03283(.A0(new_n4284_), .A1(new_n4281_), .B0(new_n4285_), .Y(new_n4286_));
  NAND2  g03284(.A(new_n4286_), .B(new_n4264_), .Y(new_n4287_));
  NOR4   g03285(.A(new_n4276_), .B(new_n4270_), .C(new_n4268_), .D(new_n4281_), .Y(new_n4288_));
  OAI211 g03286(.A0(new_n4284_), .A1(new_n4281_), .B0(new_n4288_), .B1(new_n4263_), .Y(new_n4289_));
  AOI21  g03287(.A0(new_n4289_), .A1(new_n4287_), .B0(new_n4280_), .Y(new_n4290_));
  NOR2   g03288(.A(new_n4290_), .B(new_n4273_), .Y(new_n4291_));
  OAI21  g03289(.A0(new_n4235_), .A1(new_n4225_), .B0(new_n4291_), .Y(new_n4292_));
  AOI211 g03290(.A0(new_n4223_), .A1(new_n4186_), .B(new_n4234_), .C(new_n4211_), .Y(new_n4293_));
  AOI21  g03291(.A0(new_n4233_), .A1(new_n4232_), .B0(new_n4224_), .Y(new_n4294_));
  OAI22  g03292(.A0(new_n4294_), .A1(new_n4293_), .B0(new_n4290_), .B1(new_n4273_), .Y(new_n4295_));
  NAND2  g03293(.A(new_n4295_), .B(new_n4292_), .Y(new_n4296_));
  XOR2   g03294(.A(new_n3124_), .B(new_n3117_), .Y(new_n4297_));
  XOR2   g03295(.A(new_n3128_), .B(new_n3126_), .Y(new_n4298_));
  NOR2   g03296(.A(new_n3124_), .B(new_n3117_), .Y(new_n4299_));
  NAND2  g03297(.A(new_n4299_), .B(new_n4298_), .Y(new_n4300_));
  OAI21  g03298(.A0(new_n3128_), .A1(new_n3126_), .B0(new_n4300_), .Y(new_n4301_));
  INV    g03299(.A(new_n3123_), .Y(new_n4302_));
  NAND2  g03300(.A(\A[539] ), .B(\A[538] ), .Y(new_n4303_));
  OAI21  g03301(.A0(new_n4302_), .A1(new_n3118_), .B0(new_n4303_), .Y(new_n4304_));
  XOR2   g03302(.A(new_n3128_), .B(new_n4304_), .Y(new_n4305_));
  XOR2   g03303(.A(new_n4299_), .B(new_n4305_), .Y(new_n4306_));
  AOI21  g03304(.A0(new_n4301_), .A1(new_n4297_), .B0(new_n4306_), .Y(new_n4307_));
  XOR2   g03305(.A(new_n3105_), .B(new_n3098_), .Y(new_n4308_));
  NOR2   g03306(.A(\A[542] ), .B(new_n3095_), .Y(new_n4309_));
  OAI21  g03307(.A0(new_n3093_), .A1(\A[541] ), .B0(\A[543] ), .Y(new_n4310_));
  NAND2  g03308(.A(new_n3097_), .B(new_n3092_), .Y(new_n4311_));
  OAI21  g03309(.A0(new_n4310_), .A1(new_n4309_), .B0(new_n4311_), .Y(new_n4312_));
  NOR2   g03310(.A(\A[545] ), .B(new_n3102_), .Y(new_n4313_));
  OAI21  g03311(.A0(new_n3100_), .A1(\A[544] ), .B0(\A[546] ), .Y(new_n4314_));
  NAND2  g03312(.A(new_n3104_), .B(new_n3099_), .Y(new_n4315_));
  OAI21  g03313(.A0(new_n4314_), .A1(new_n4313_), .B0(new_n4315_), .Y(new_n4316_));
  NAND2  g03314(.A(new_n3104_), .B(\A[546] ), .Y(new_n4317_));
  OAI21  g03315(.A0(new_n3100_), .A1(new_n3102_), .B0(new_n4317_), .Y(new_n4318_));
  NAND2  g03316(.A(new_n3097_), .B(\A[543] ), .Y(new_n4319_));
  OAI21  g03317(.A0(new_n3093_), .A1(new_n3095_), .B0(new_n4319_), .Y(new_n4320_));
  NAND4  g03318(.A(new_n4320_), .B(new_n4318_), .C(new_n4316_), .D(new_n4312_), .Y(new_n4321_));
  INV    g03319(.A(new_n3116_), .Y(new_n4322_));
  NOR2   g03320(.A(new_n4322_), .B(new_n3111_), .Y(new_n4323_));
  OAI211 g03321(.A0(new_n4323_), .A1(new_n3127_), .B0(new_n4299_), .B1(new_n4304_), .Y(new_n4324_));
  NAND4  g03322(.A(new_n4324_), .B(new_n4297_), .C(new_n4321_), .D(new_n4308_), .Y(new_n4325_));
  XOR2   g03323(.A(new_n3109_), .B(new_n4318_), .Y(new_n4326_));
  NAND2  g03324(.A(new_n4316_), .B(new_n4312_), .Y(new_n4327_));
  NAND2  g03325(.A(new_n4320_), .B(new_n4318_), .Y(new_n4328_));
  OAI21  g03326(.A0(new_n4327_), .A1(new_n4326_), .B0(new_n4328_), .Y(new_n4329_));
  NOR2   g03327(.A(new_n3105_), .B(new_n3098_), .Y(new_n4330_));
  XOR2   g03328(.A(new_n4330_), .B(new_n4326_), .Y(new_n4331_));
  AOI21  g03329(.A0(new_n4329_), .A1(new_n4308_), .B0(new_n4331_), .Y(new_n4332_));
  XOR2   g03330(.A(new_n4332_), .B(new_n4325_), .Y(new_n4333_));
  NOR2   g03331(.A(new_n4333_), .B(new_n4307_), .Y(new_n4334_));
  NAND2  g03332(.A(new_n3115_), .B(new_n3113_), .Y(new_n4335_));
  OAI21  g03333(.A0(new_n4322_), .A1(\A[537] ), .B0(new_n4335_), .Y(new_n4336_));
  XOR2   g03334(.A(new_n3124_), .B(new_n4336_), .Y(new_n4337_));
  NOR2   g03335(.A(new_n3128_), .B(new_n3126_), .Y(new_n4338_));
  AOI21  g03336(.A0(new_n4299_), .A1(new_n4298_), .B0(new_n4338_), .Y(new_n4339_));
  XOR2   g03337(.A(new_n4299_), .B(new_n4298_), .Y(new_n4340_));
  OAI21  g03338(.A0(new_n4339_), .A1(new_n4337_), .B0(new_n4340_), .Y(new_n4341_));
  XOR2   g03339(.A(new_n3105_), .B(new_n4312_), .Y(new_n4342_));
  XOR2   g03340(.A(new_n3109_), .B(new_n3107_), .Y(new_n4343_));
  NOR2   g03341(.A(new_n3109_), .B(new_n3107_), .Y(new_n4344_));
  AOI21  g03342(.A0(new_n4330_), .A1(new_n4343_), .B0(new_n4344_), .Y(new_n4345_));
  XOR2   g03343(.A(new_n4330_), .B(new_n4343_), .Y(new_n4346_));
  OAI21  g03344(.A0(new_n4345_), .A1(new_n4342_), .B0(new_n4346_), .Y(new_n4347_));
  NAND2  g03345(.A(new_n4347_), .B(new_n4325_), .Y(new_n4348_));
  NOR4   g03346(.A(new_n4337_), .B(new_n4331_), .C(new_n4329_), .D(new_n4342_), .Y(new_n4349_));
  OAI211 g03347(.A0(new_n4345_), .A1(new_n4342_), .B0(new_n4349_), .B1(new_n4324_), .Y(new_n4350_));
  AOI21  g03348(.A0(new_n4350_), .A1(new_n4348_), .B0(new_n4341_), .Y(new_n4351_));
  NOR2   g03349(.A(new_n4351_), .B(new_n4334_), .Y(new_n4352_));
  NAND2  g03350(.A(new_n3130_), .B(new_n3091_), .Y(new_n4353_));
  INV    g03351(.A(new_n4353_), .Y(new_n4354_));
  NOR2   g03352(.A(\A[548] ), .B(new_n3074_), .Y(new_n4355_));
  OAI21  g03353(.A0(new_n3072_), .A1(\A[547] ), .B0(\A[549] ), .Y(new_n4356_));
  XOR2   g03354(.A(\A[548] ), .B(new_n3074_), .Y(new_n4357_));
  OAI22  g03355(.A0(new_n4357_), .A1(\A[549] ), .B0(new_n4356_), .B1(new_n4355_), .Y(new_n4358_));
  XOR2   g03356(.A(new_n3084_), .B(new_n4358_), .Y(new_n4359_));
  XOR2   g03357(.A(new_n3089_), .B(new_n3087_), .Y(new_n4360_));
  NOR2   g03358(.A(new_n3084_), .B(new_n3077_), .Y(new_n4361_));
  NOR2   g03359(.A(new_n3089_), .B(new_n3087_), .Y(new_n4362_));
  AOI21  g03360(.A0(new_n4361_), .A1(new_n4360_), .B0(new_n4362_), .Y(new_n4363_));
  XOR2   g03361(.A(new_n4361_), .B(new_n4360_), .Y(new_n4364_));
  OAI21  g03362(.A0(new_n4363_), .A1(new_n4359_), .B0(new_n4364_), .Y(new_n4365_));
  NOR2   g03363(.A(\A[554] ), .B(new_n3055_), .Y(new_n4366_));
  OAI21  g03364(.A0(new_n3053_), .A1(\A[553] ), .B0(\A[555] ), .Y(new_n4367_));
  NAND2  g03365(.A(new_n3057_), .B(new_n3052_), .Y(new_n4368_));
  OAI21  g03366(.A0(new_n4367_), .A1(new_n4366_), .B0(new_n4368_), .Y(new_n4369_));
  XOR2   g03367(.A(new_n3065_), .B(new_n4369_), .Y(new_n4370_));
  NOR4   g03368(.A(new_n3069_), .B(new_n3067_), .C(new_n3065_), .D(new_n3058_), .Y(new_n4371_));
  NOR4   g03369(.A(new_n3089_), .B(new_n3087_), .C(new_n3084_), .D(new_n3077_), .Y(new_n4372_));
  NOR4   g03370(.A(new_n4372_), .B(new_n4359_), .C(new_n4371_), .D(new_n4370_), .Y(new_n4373_));
  XOR2   g03371(.A(new_n3065_), .B(new_n3058_), .Y(new_n4374_));
  NAND2  g03372(.A(new_n3064_), .B(\A[558] ), .Y(new_n4375_));
  OAI21  g03373(.A0(new_n3060_), .A1(new_n3062_), .B0(new_n4375_), .Y(new_n4376_));
  XOR2   g03374(.A(new_n3069_), .B(new_n4376_), .Y(new_n4377_));
  NOR2   g03375(.A(\A[557] ), .B(new_n3062_), .Y(new_n4378_));
  OAI21  g03376(.A0(new_n3060_), .A1(\A[556] ), .B0(\A[558] ), .Y(new_n4379_));
  NAND2  g03377(.A(new_n3064_), .B(new_n3059_), .Y(new_n4380_));
  OAI21  g03378(.A0(new_n4379_), .A1(new_n4378_), .B0(new_n4380_), .Y(new_n4381_));
  NAND2  g03379(.A(new_n4381_), .B(new_n4369_), .Y(new_n4382_));
  NAND2  g03380(.A(new_n3057_), .B(\A[555] ), .Y(new_n4383_));
  OAI21  g03381(.A0(new_n3053_), .A1(new_n3055_), .B0(new_n4383_), .Y(new_n4384_));
  NAND2  g03382(.A(new_n4384_), .B(new_n4376_), .Y(new_n4385_));
  OAI21  g03383(.A0(new_n4382_), .A1(new_n4377_), .B0(new_n4385_), .Y(new_n4386_));
  NOR2   g03384(.A(new_n3065_), .B(new_n3058_), .Y(new_n4387_));
  XOR2   g03385(.A(new_n4387_), .B(new_n4377_), .Y(new_n4388_));
  AOI21  g03386(.A0(new_n4386_), .A1(new_n4374_), .B0(new_n4388_), .Y(new_n4389_));
  XOR2   g03387(.A(new_n4389_), .B(new_n4373_), .Y(new_n4390_));
  NAND2  g03388(.A(new_n4390_), .B(new_n4365_), .Y(new_n4391_));
  XOR2   g03389(.A(new_n3084_), .B(new_n3077_), .Y(new_n4392_));
  XOR2   g03390(.A(\A[551] ), .B(new_n3081_), .Y(new_n4393_));
  OAI21  g03391(.A0(new_n4393_), .A1(new_n3078_), .B0(new_n3085_), .Y(new_n4394_));
  XOR2   g03392(.A(new_n3089_), .B(new_n4394_), .Y(new_n4395_));
  NOR2   g03393(.A(\A[551] ), .B(new_n3081_), .Y(new_n4396_));
  OAI21  g03394(.A0(new_n3079_), .A1(\A[550] ), .B0(\A[552] ), .Y(new_n4397_));
  OAI22  g03395(.A0(new_n4393_), .A1(\A[552] ), .B0(new_n4397_), .B1(new_n4396_), .Y(new_n4398_));
  NAND2  g03396(.A(new_n4398_), .B(new_n4358_), .Y(new_n4399_));
  NAND2  g03397(.A(\A[548] ), .B(\A[547] ), .Y(new_n4400_));
  OAI21  g03398(.A0(new_n4357_), .A1(new_n3071_), .B0(new_n4400_), .Y(new_n4401_));
  NAND2  g03399(.A(new_n4401_), .B(new_n4394_), .Y(new_n4402_));
  OAI21  g03400(.A0(new_n4399_), .A1(new_n4395_), .B0(new_n4402_), .Y(new_n4403_));
  XOR2   g03401(.A(new_n4361_), .B(new_n4395_), .Y(new_n4404_));
  AOI21  g03402(.A0(new_n4403_), .A1(new_n4392_), .B0(new_n4404_), .Y(new_n4405_));
  XOR2   g03403(.A(new_n3069_), .B(new_n3067_), .Y(new_n4406_));
  XOR2   g03404(.A(new_n4387_), .B(new_n4406_), .Y(new_n4407_));
  NAND4  g03405(.A(new_n4384_), .B(new_n4376_), .C(new_n4381_), .D(new_n4369_), .Y(new_n4408_));
  NAND4  g03406(.A(new_n4392_), .B(new_n4408_), .C(new_n4407_), .D(new_n4374_), .Y(new_n4409_));
  NOR2   g03407(.A(new_n3069_), .B(new_n3067_), .Y(new_n4410_));
  AOI21  g03408(.A0(new_n4387_), .A1(new_n4406_), .B0(new_n4410_), .Y(new_n4411_));
  NAND4  g03409(.A(new_n4401_), .B(new_n4394_), .C(new_n4398_), .D(new_n4358_), .Y(new_n4412_));
  OAI21  g03410(.A0(new_n4411_), .A1(new_n4370_), .B0(new_n4412_), .Y(new_n4413_));
  OAI22  g03411(.A0(new_n4413_), .A1(new_n4409_), .B0(new_n4389_), .B1(new_n4373_), .Y(new_n4414_));
  NAND2  g03412(.A(new_n4414_), .B(new_n4405_), .Y(new_n4415_));
  NAND3  g03413(.A(new_n4354_), .B(new_n4415_), .C(new_n4391_), .Y(new_n4416_));
  NAND4  g03414(.A(new_n4412_), .B(new_n4392_), .C(new_n4408_), .D(new_n4374_), .Y(new_n4417_));
  XOR2   g03415(.A(new_n4389_), .B(new_n4417_), .Y(new_n4418_));
  NOR2   g03416(.A(new_n4418_), .B(new_n4405_), .Y(new_n4419_));
  AOI21  g03417(.A0(new_n4414_), .A1(new_n4405_), .B0(new_n4419_), .Y(new_n4420_));
  OAI21  g03418(.A0(new_n4420_), .A1(new_n4354_), .B0(new_n4416_), .Y(new_n4421_));
  NAND2  g03419(.A(new_n4421_), .B(new_n4352_), .Y(new_n4422_));
  AOI211 g03420(.A0(new_n4414_), .A1(new_n4405_), .B(new_n4354_), .C(new_n4419_), .Y(new_n4423_));
  AOI21  g03421(.A0(new_n4415_), .A1(new_n4391_), .B0(new_n4353_), .Y(new_n4424_));
  OAI22  g03422(.A0(new_n4424_), .A1(new_n4423_), .B0(new_n4351_), .B1(new_n4334_), .Y(new_n4425_));
  NOR2   g03423(.A(new_n3213_), .B(new_n3132_), .Y(new_n4426_));
  NAND3  g03424(.A(new_n4426_), .B(new_n4425_), .C(new_n4422_), .Y(new_n4427_));
  NAND2  g03425(.A(new_n4350_), .B(new_n4348_), .Y(new_n4428_));
  NAND2  g03426(.A(new_n4428_), .B(new_n4307_), .Y(new_n4429_));
  OAI21  g03427(.A0(new_n4333_), .A1(new_n4307_), .B0(new_n4429_), .Y(new_n4430_));
  NOR2   g03428(.A(new_n4389_), .B(new_n4373_), .Y(new_n4431_));
  NOR2   g03429(.A(new_n4413_), .B(new_n4409_), .Y(new_n4432_));
  NOR2   g03430(.A(new_n4432_), .B(new_n4431_), .Y(new_n4433_));
  NOR2   g03431(.A(new_n4433_), .B(new_n4365_), .Y(new_n4434_));
  OAI21  g03432(.A0(new_n4434_), .A1(new_n4419_), .B0(new_n4353_), .Y(new_n4435_));
  AOI21  g03433(.A0(new_n4435_), .A1(new_n4416_), .B0(new_n4430_), .Y(new_n4436_));
  NAND3  g03434(.A(new_n4353_), .B(new_n4415_), .C(new_n4391_), .Y(new_n4437_));
  OAI21  g03435(.A0(new_n4434_), .A1(new_n4419_), .B0(new_n4354_), .Y(new_n4438_));
  AOI21  g03436(.A0(new_n4438_), .A1(new_n4437_), .B0(new_n4352_), .Y(new_n4439_));
  INV    g03437(.A(new_n4426_), .Y(new_n4440_));
  OAI21  g03438(.A0(new_n4439_), .A1(new_n4436_), .B0(new_n4440_), .Y(new_n4441_));
  AOI21  g03439(.A0(new_n4441_), .A1(new_n4427_), .B0(new_n4296_), .Y(new_n4442_));
  NOR2   g03440(.A(new_n4235_), .B(new_n4225_), .Y(new_n4443_));
  NAND2  g03441(.A(new_n4289_), .B(new_n4287_), .Y(new_n4444_));
  NAND2  g03442(.A(new_n4444_), .B(new_n4246_), .Y(new_n4445_));
  OAI21  g03443(.A0(new_n4272_), .A1(new_n4246_), .B0(new_n4445_), .Y(new_n4446_));
  NOR2   g03444(.A(new_n4446_), .B(new_n4443_), .Y(new_n4447_));
  NAND3  g03445(.A(new_n4224_), .B(new_n4233_), .C(new_n4232_), .Y(new_n4448_));
  NAND2  g03446(.A(new_n4233_), .B(new_n4232_), .Y(new_n4449_));
  NAND2  g03447(.A(new_n4449_), .B(new_n4234_), .Y(new_n4450_));
  AOI21  g03448(.A0(new_n4450_), .A1(new_n4448_), .B0(new_n4291_), .Y(new_n4451_));
  NOR2   g03449(.A(new_n4451_), .B(new_n4447_), .Y(new_n4452_));
  OAI21  g03450(.A0(new_n4420_), .A1(new_n4353_), .B0(new_n4437_), .Y(new_n4453_));
  AOI21  g03451(.A0(new_n4453_), .A1(new_n4430_), .B0(new_n4426_), .Y(new_n4454_));
  NAND2  g03452(.A(new_n4454_), .B(new_n4422_), .Y(new_n4455_));
  OAI21  g03453(.A0(new_n4439_), .A1(new_n4436_), .B0(new_n4426_), .Y(new_n4456_));
  AOI21  g03454(.A0(new_n4456_), .A1(new_n4455_), .B0(new_n4452_), .Y(new_n4457_));
  NOR2   g03455(.A(new_n3214_), .B(new_n3050_), .Y(new_n4458_));
  INV    g03456(.A(new_n4458_), .Y(new_n4459_));
  NOR3   g03457(.A(new_n4459_), .B(new_n4457_), .C(new_n4442_), .Y(new_n4460_));
  NOR3   g03458(.A(new_n4440_), .B(new_n4439_), .C(new_n4436_), .Y(new_n4461_));
  AOI21  g03459(.A0(new_n4425_), .A1(new_n4422_), .B0(new_n4426_), .Y(new_n4462_));
  OAI21  g03460(.A0(new_n4462_), .A1(new_n4461_), .B0(new_n4452_), .Y(new_n4463_));
  NOR3   g03461(.A(new_n4426_), .B(new_n4439_), .C(new_n4436_), .Y(new_n4464_));
  AOI21  g03462(.A0(new_n4425_), .A1(new_n4422_), .B0(new_n4440_), .Y(new_n4465_));
  OAI21  g03463(.A0(new_n4465_), .A1(new_n4464_), .B0(new_n4296_), .Y(new_n4466_));
  AOI21  g03464(.A0(new_n4466_), .A1(new_n4463_), .B0(new_n4458_), .Y(new_n4467_));
  XOR2   g03465(.A(new_n3041_), .B(new_n3034_), .Y(new_n4468_));
  XOR2   g03466(.A(\A[491] ), .B(new_n3038_), .Y(new_n4469_));
  NAND2  g03467(.A(\A[491] ), .B(\A[490] ), .Y(new_n4470_));
  OAI21  g03468(.A0(new_n4469_), .A1(new_n3035_), .B0(new_n4470_), .Y(new_n4471_));
  XOR2   g03469(.A(new_n3045_), .B(new_n4471_), .Y(new_n4472_));
  NOR2   g03470(.A(\A[488] ), .B(new_n3031_), .Y(new_n4473_));
  OAI21  g03471(.A0(new_n3029_), .A1(\A[487] ), .B0(\A[489] ), .Y(new_n4474_));
  XOR2   g03472(.A(\A[488] ), .B(new_n3031_), .Y(new_n4475_));
  OAI22  g03473(.A0(new_n4475_), .A1(\A[489] ), .B0(new_n4474_), .B1(new_n4473_), .Y(new_n4476_));
  NOR2   g03474(.A(\A[491] ), .B(new_n3038_), .Y(new_n4477_));
  OAI21  g03475(.A0(new_n3036_), .A1(\A[490] ), .B0(\A[492] ), .Y(new_n4478_));
  OAI22  g03476(.A0(new_n4469_), .A1(\A[492] ), .B0(new_n4478_), .B1(new_n4477_), .Y(new_n4479_));
  NAND2  g03477(.A(new_n4479_), .B(new_n4476_), .Y(new_n4480_));
  NAND2  g03478(.A(\A[488] ), .B(\A[487] ), .Y(new_n4481_));
  OAI21  g03479(.A0(new_n4475_), .A1(new_n3028_), .B0(new_n4481_), .Y(new_n4482_));
  NAND2  g03480(.A(new_n4482_), .B(new_n4471_), .Y(new_n4483_));
  OAI21  g03481(.A0(new_n4480_), .A1(new_n4472_), .B0(new_n4483_), .Y(new_n4484_));
  NOR2   g03482(.A(new_n3041_), .B(new_n3034_), .Y(new_n4485_));
  XOR2   g03483(.A(new_n4485_), .B(new_n4472_), .Y(new_n4486_));
  AOI21  g03484(.A0(new_n4484_), .A1(new_n4468_), .B0(new_n4486_), .Y(new_n4487_));
  XOR2   g03485(.A(new_n3022_), .B(new_n3015_), .Y(new_n4488_));
  NOR2   g03486(.A(\A[494] ), .B(new_n3012_), .Y(new_n4489_));
  OAI21  g03487(.A0(new_n3010_), .A1(\A[493] ), .B0(\A[495] ), .Y(new_n4490_));
  NAND2  g03488(.A(new_n3014_), .B(new_n3009_), .Y(new_n4491_));
  OAI21  g03489(.A0(new_n4490_), .A1(new_n4489_), .B0(new_n4491_), .Y(new_n4492_));
  NOR2   g03490(.A(\A[497] ), .B(new_n3019_), .Y(new_n4493_));
  OAI21  g03491(.A0(new_n3017_), .A1(\A[496] ), .B0(\A[498] ), .Y(new_n4494_));
  NAND2  g03492(.A(new_n3021_), .B(new_n3016_), .Y(new_n4495_));
  OAI21  g03493(.A0(new_n4494_), .A1(new_n4493_), .B0(new_n4495_), .Y(new_n4496_));
  NAND2  g03494(.A(new_n3021_), .B(\A[498] ), .Y(new_n4497_));
  OAI21  g03495(.A0(new_n3017_), .A1(new_n3019_), .B0(new_n4497_), .Y(new_n4498_));
  NAND2  g03496(.A(new_n3014_), .B(\A[495] ), .Y(new_n4499_));
  OAI21  g03497(.A0(new_n3010_), .A1(new_n3012_), .B0(new_n4499_), .Y(new_n4500_));
  NAND4  g03498(.A(new_n4500_), .B(new_n4498_), .C(new_n4496_), .D(new_n4492_), .Y(new_n4501_));
  NAND4  g03499(.A(new_n4482_), .B(new_n4471_), .C(new_n4479_), .D(new_n4476_), .Y(new_n4502_));
  NAND4  g03500(.A(new_n4502_), .B(new_n4468_), .C(new_n4501_), .D(new_n4488_), .Y(new_n4503_));
  XOR2   g03501(.A(new_n3026_), .B(new_n4498_), .Y(new_n4504_));
  NAND2  g03502(.A(new_n4496_), .B(new_n4492_), .Y(new_n4505_));
  NAND2  g03503(.A(new_n4500_), .B(new_n4498_), .Y(new_n4506_));
  OAI21  g03504(.A0(new_n4505_), .A1(new_n4504_), .B0(new_n4506_), .Y(new_n4507_));
  NOR2   g03505(.A(new_n3022_), .B(new_n3015_), .Y(new_n4508_));
  XOR2   g03506(.A(new_n4508_), .B(new_n4504_), .Y(new_n4509_));
  AOI21  g03507(.A0(new_n4507_), .A1(new_n4488_), .B0(new_n4509_), .Y(new_n4510_));
  XOR2   g03508(.A(new_n4510_), .B(new_n4503_), .Y(new_n4511_));
  XOR2   g03509(.A(new_n3022_), .B(new_n4492_), .Y(new_n4512_));
  NOR4   g03510(.A(new_n3026_), .B(new_n3024_), .C(new_n3022_), .D(new_n3015_), .Y(new_n4513_));
  XOR2   g03511(.A(new_n3041_), .B(new_n4476_), .Y(new_n4514_));
  NOR4   g03512(.A(new_n3045_), .B(new_n3043_), .C(new_n3041_), .D(new_n3034_), .Y(new_n4515_));
  NOR4   g03513(.A(new_n4515_), .B(new_n4514_), .C(new_n4513_), .D(new_n4512_), .Y(new_n4516_));
  XOR2   g03514(.A(new_n3026_), .B(new_n3024_), .Y(new_n4517_));
  NOR2   g03515(.A(new_n3026_), .B(new_n3024_), .Y(new_n4518_));
  AOI21  g03516(.A0(new_n4508_), .A1(new_n4517_), .B0(new_n4518_), .Y(new_n4519_));
  NOR4   g03517(.A(new_n4514_), .B(new_n4513_), .C(new_n4509_), .D(new_n4512_), .Y(new_n4520_));
  OAI211 g03518(.A0(new_n4519_), .A1(new_n4512_), .B0(new_n4520_), .B1(new_n4502_), .Y(new_n4521_));
  OAI21  g03519(.A0(new_n4510_), .A1(new_n4516_), .B0(new_n4521_), .Y(new_n4522_));
  NAND2  g03520(.A(new_n4522_), .B(new_n4487_), .Y(new_n4523_));
  OAI21  g03521(.A0(new_n4511_), .A1(new_n4487_), .B0(new_n4523_), .Y(new_n4524_));
  NOR2   g03522(.A(\A[500] ), .B(new_n2992_), .Y(new_n4525_));
  OAI21  g03523(.A0(new_n2990_), .A1(\A[499] ), .B0(\A[501] ), .Y(new_n4526_));
  XOR2   g03524(.A(\A[500] ), .B(new_n2992_), .Y(new_n4527_));
  OAI22  g03525(.A0(new_n4527_), .A1(\A[501] ), .B0(new_n4526_), .B1(new_n4525_), .Y(new_n4528_));
  XOR2   g03526(.A(new_n3002_), .B(new_n4528_), .Y(new_n4529_));
  XOR2   g03527(.A(new_n3006_), .B(new_n3004_), .Y(new_n4530_));
  NOR2   g03528(.A(new_n3002_), .B(new_n2995_), .Y(new_n4531_));
  NOR2   g03529(.A(new_n3006_), .B(new_n3004_), .Y(new_n4532_));
  AOI21  g03530(.A0(new_n4531_), .A1(new_n4530_), .B0(new_n4532_), .Y(new_n4533_));
  XOR2   g03531(.A(new_n4531_), .B(new_n4530_), .Y(new_n4534_));
  OAI21  g03532(.A0(new_n4533_), .A1(new_n4529_), .B0(new_n4534_), .Y(new_n4535_));
  NOR2   g03533(.A(\A[506] ), .B(new_n2973_), .Y(new_n4536_));
  OAI21  g03534(.A0(new_n2971_), .A1(\A[505] ), .B0(\A[507] ), .Y(new_n4537_));
  NAND2  g03535(.A(new_n2975_), .B(new_n2970_), .Y(new_n4538_));
  OAI21  g03536(.A0(new_n4537_), .A1(new_n4536_), .B0(new_n4538_), .Y(new_n4539_));
  XOR2   g03537(.A(new_n2983_), .B(new_n4539_), .Y(new_n4540_));
  NOR4   g03538(.A(new_n2987_), .B(new_n2985_), .C(new_n2983_), .D(new_n2976_), .Y(new_n4541_));
  NOR4   g03539(.A(new_n3006_), .B(new_n3004_), .C(new_n3002_), .D(new_n2995_), .Y(new_n4542_));
  NOR4   g03540(.A(new_n4542_), .B(new_n4529_), .C(new_n4541_), .D(new_n4540_), .Y(new_n4543_));
  XOR2   g03541(.A(new_n2983_), .B(new_n2976_), .Y(new_n4544_));
  NAND2  g03542(.A(new_n2982_), .B(\A[510] ), .Y(new_n4545_));
  OAI21  g03543(.A0(new_n2978_), .A1(new_n2980_), .B0(new_n4545_), .Y(new_n4546_));
  XOR2   g03544(.A(new_n2987_), .B(new_n4546_), .Y(new_n4547_));
  NOR2   g03545(.A(\A[509] ), .B(new_n2980_), .Y(new_n4548_));
  OAI21  g03546(.A0(new_n2978_), .A1(\A[508] ), .B0(\A[510] ), .Y(new_n4549_));
  NAND2  g03547(.A(new_n2982_), .B(new_n2977_), .Y(new_n4550_));
  OAI21  g03548(.A0(new_n4549_), .A1(new_n4548_), .B0(new_n4550_), .Y(new_n4551_));
  NAND2  g03549(.A(new_n4551_), .B(new_n4539_), .Y(new_n4552_));
  NAND2  g03550(.A(new_n2975_), .B(\A[507] ), .Y(new_n4553_));
  OAI21  g03551(.A0(new_n2971_), .A1(new_n2973_), .B0(new_n4553_), .Y(new_n4554_));
  NAND2  g03552(.A(new_n4554_), .B(new_n4546_), .Y(new_n4555_));
  OAI21  g03553(.A0(new_n4552_), .A1(new_n4547_), .B0(new_n4555_), .Y(new_n4556_));
  NOR2   g03554(.A(new_n2983_), .B(new_n2976_), .Y(new_n4557_));
  XOR2   g03555(.A(new_n4557_), .B(new_n4547_), .Y(new_n4558_));
  AOI21  g03556(.A0(new_n4556_), .A1(new_n4544_), .B0(new_n4558_), .Y(new_n4559_));
  XOR2   g03557(.A(new_n4559_), .B(new_n4543_), .Y(new_n4560_));
  NAND2  g03558(.A(new_n4560_), .B(new_n4535_), .Y(new_n4561_));
  XOR2   g03559(.A(new_n3002_), .B(new_n2995_), .Y(new_n4562_));
  XOR2   g03560(.A(\A[503] ), .B(new_n2999_), .Y(new_n4563_));
  NAND2  g03561(.A(\A[503] ), .B(\A[502] ), .Y(new_n4564_));
  OAI21  g03562(.A0(new_n4563_), .A1(new_n2996_), .B0(new_n4564_), .Y(new_n4565_));
  XOR2   g03563(.A(new_n3006_), .B(new_n4565_), .Y(new_n4566_));
  NOR2   g03564(.A(\A[503] ), .B(new_n2999_), .Y(new_n4567_));
  OAI21  g03565(.A0(new_n2997_), .A1(\A[502] ), .B0(\A[504] ), .Y(new_n4568_));
  OAI22  g03566(.A0(new_n4563_), .A1(\A[504] ), .B0(new_n4568_), .B1(new_n4567_), .Y(new_n4569_));
  NAND2  g03567(.A(new_n4569_), .B(new_n4528_), .Y(new_n4570_));
  NAND2  g03568(.A(\A[500] ), .B(\A[499] ), .Y(new_n4571_));
  OAI21  g03569(.A0(new_n4527_), .A1(new_n2989_), .B0(new_n4571_), .Y(new_n4572_));
  NAND2  g03570(.A(new_n4572_), .B(new_n4565_), .Y(new_n4573_));
  OAI21  g03571(.A0(new_n4570_), .A1(new_n4566_), .B0(new_n4573_), .Y(new_n4574_));
  XOR2   g03572(.A(new_n4531_), .B(new_n4566_), .Y(new_n4575_));
  AOI21  g03573(.A0(new_n4574_), .A1(new_n4562_), .B0(new_n4575_), .Y(new_n4576_));
  XOR2   g03574(.A(new_n2987_), .B(new_n2985_), .Y(new_n4577_));
  XOR2   g03575(.A(new_n4557_), .B(new_n4577_), .Y(new_n4578_));
  NAND4  g03576(.A(new_n4554_), .B(new_n4546_), .C(new_n4551_), .D(new_n4539_), .Y(new_n4579_));
  NAND4  g03577(.A(new_n4562_), .B(new_n4579_), .C(new_n4578_), .D(new_n4544_), .Y(new_n4580_));
  NOR2   g03578(.A(new_n2987_), .B(new_n2985_), .Y(new_n4581_));
  AOI21  g03579(.A0(new_n4557_), .A1(new_n4577_), .B0(new_n4581_), .Y(new_n4582_));
  NAND4  g03580(.A(new_n4572_), .B(new_n4565_), .C(new_n4569_), .D(new_n4528_), .Y(new_n4583_));
  OAI21  g03581(.A0(new_n4582_), .A1(new_n4540_), .B0(new_n4583_), .Y(new_n4584_));
  OAI22  g03582(.A0(new_n4584_), .A1(new_n4580_), .B0(new_n4559_), .B1(new_n4543_), .Y(new_n4585_));
  NAND2  g03583(.A(new_n4585_), .B(new_n4576_), .Y(new_n4586_));
  NAND2  g03584(.A(new_n3047_), .B(new_n3008_), .Y(new_n4587_));
  INV    g03585(.A(new_n4587_), .Y(new_n4588_));
  NAND3  g03586(.A(new_n4588_), .B(new_n4586_), .C(new_n4561_), .Y(new_n4589_));
  NAND2  g03587(.A(new_n4586_), .B(new_n4561_), .Y(new_n4590_));
  NAND2  g03588(.A(new_n4590_), .B(new_n4587_), .Y(new_n4591_));
  AOI21  g03589(.A0(new_n4591_), .A1(new_n4589_), .B0(new_n4524_), .Y(new_n4592_));
  NOR2   g03590(.A(new_n4511_), .B(new_n4487_), .Y(new_n4593_));
  AOI21  g03591(.A0(new_n4522_), .A1(new_n4487_), .B0(new_n4593_), .Y(new_n4594_));
  NAND4  g03592(.A(new_n4583_), .B(new_n4562_), .C(new_n4579_), .D(new_n4544_), .Y(new_n4595_));
  XOR2   g03593(.A(new_n4559_), .B(new_n4595_), .Y(new_n4596_));
  NOR2   g03594(.A(new_n4596_), .B(new_n4576_), .Y(new_n4597_));
  AOI211 g03595(.A0(new_n4585_), .A1(new_n4576_), .B(new_n4588_), .C(new_n4597_), .Y(new_n4598_));
  AOI21  g03596(.A0(new_n4586_), .A1(new_n4561_), .B0(new_n4587_), .Y(new_n4599_));
  NOR2   g03597(.A(new_n4599_), .B(new_n4598_), .Y(new_n4600_));
  NOR2   g03598(.A(new_n3049_), .B(new_n2968_), .Y(new_n4601_));
  OAI21  g03599(.A0(new_n4600_), .A1(new_n4594_), .B0(new_n4601_), .Y(new_n4602_));
  NOR2   g03600(.A(new_n4600_), .B(new_n4594_), .Y(new_n4603_));
  INV    g03601(.A(new_n4601_), .Y(new_n4604_));
  OAI21  g03602(.A0(new_n4603_), .A1(new_n4592_), .B0(new_n4604_), .Y(new_n4605_));
  OAI21  g03603(.A0(new_n4602_), .A1(new_n4592_), .B0(new_n4605_), .Y(new_n4606_));
  NOR2   g03604(.A(new_n2910_), .B(new_n2903_), .Y(new_n4607_));
  NOR2   g03605(.A(new_n2905_), .B(new_n2907_), .Y(new_n4608_));
  AOI21  g03606(.A0(new_n2909_), .A1(\A[465] ), .B0(new_n4608_), .Y(new_n4609_));
  XOR2   g03607(.A(new_n4609_), .B(new_n2922_), .Y(new_n4610_));
  XOR2   g03608(.A(new_n4610_), .B(new_n4607_), .Y(new_n4611_));
  NAND2  g03609(.A(new_n2919_), .B(new_n2915_), .Y(new_n4612_));
  NAND2  g03610(.A(new_n2924_), .B(new_n2922_), .Y(new_n4613_));
  OAI21  g03611(.A0(new_n4610_), .A1(new_n4612_), .B0(new_n4613_), .Y(new_n4614_));
  AOI21  g03612(.A0(new_n4614_), .A1(new_n2911_), .B0(new_n4611_), .Y(new_n4615_));
  XOR2   g03613(.A(new_n2890_), .B(new_n2883_), .Y(new_n4616_));
  NOR2   g03614(.A(\A[470] ), .B(new_n2880_), .Y(new_n4617_));
  OAI21  g03615(.A0(new_n2878_), .A1(\A[469] ), .B0(\A[471] ), .Y(new_n4618_));
  NAND2  g03616(.A(new_n2882_), .B(new_n2877_), .Y(new_n4619_));
  OAI21  g03617(.A0(new_n4618_), .A1(new_n4617_), .B0(new_n4619_), .Y(new_n4620_));
  NOR2   g03618(.A(\A[473] ), .B(new_n2887_), .Y(new_n4621_));
  OAI21  g03619(.A0(new_n2885_), .A1(\A[472] ), .B0(\A[474] ), .Y(new_n4622_));
  NAND2  g03620(.A(new_n2889_), .B(new_n2884_), .Y(new_n4623_));
  OAI21  g03621(.A0(new_n4622_), .A1(new_n4621_), .B0(new_n4623_), .Y(new_n4624_));
  NAND2  g03622(.A(new_n2889_), .B(\A[474] ), .Y(new_n4625_));
  OAI21  g03623(.A0(new_n2885_), .A1(new_n2887_), .B0(new_n4625_), .Y(new_n4626_));
  NAND2  g03624(.A(new_n2882_), .B(\A[471] ), .Y(new_n4627_));
  OAI21  g03625(.A0(new_n2878_), .A1(new_n2880_), .B0(new_n4627_), .Y(new_n4628_));
  NAND4  g03626(.A(new_n4628_), .B(new_n4626_), .C(new_n4624_), .D(new_n4620_), .Y(new_n4629_));
  NAND4  g03627(.A(new_n2925_), .B(new_n2911_), .C(new_n4629_), .D(new_n4616_), .Y(new_n4630_));
  XOR2   g03628(.A(new_n2894_), .B(new_n4626_), .Y(new_n4631_));
  NAND2  g03629(.A(new_n4624_), .B(new_n4620_), .Y(new_n4632_));
  NAND2  g03630(.A(new_n4628_), .B(new_n4626_), .Y(new_n4633_));
  OAI21  g03631(.A0(new_n4632_), .A1(new_n4631_), .B0(new_n4633_), .Y(new_n4634_));
  NOR2   g03632(.A(new_n2890_), .B(new_n2883_), .Y(new_n4635_));
  XOR2   g03633(.A(new_n4635_), .B(new_n4631_), .Y(new_n4636_));
  AOI21  g03634(.A0(new_n4634_), .A1(new_n4616_), .B0(new_n4636_), .Y(new_n4637_));
  XOR2   g03635(.A(new_n4637_), .B(new_n4630_), .Y(new_n4638_));
  XOR2   g03636(.A(new_n2890_), .B(new_n4620_), .Y(new_n4639_));
  NOR4   g03637(.A(new_n2894_), .B(new_n2892_), .C(new_n2890_), .D(new_n2883_), .Y(new_n4640_));
  XOR2   g03638(.A(new_n2910_), .B(new_n2915_), .Y(new_n4641_));
  AOI211 g03639(.A0(new_n2921_), .A1(new_n2920_), .B(new_n4609_), .C(new_n4612_), .Y(new_n4642_));
  NOR4   g03640(.A(new_n4642_), .B(new_n4641_), .C(new_n4640_), .D(new_n4639_), .Y(new_n4643_));
  XOR2   g03641(.A(new_n2894_), .B(new_n2892_), .Y(new_n4644_));
  NOR2   g03642(.A(new_n2894_), .B(new_n2892_), .Y(new_n4645_));
  AOI21  g03643(.A0(new_n4635_), .A1(new_n4644_), .B0(new_n4645_), .Y(new_n4646_));
  NOR4   g03644(.A(new_n4641_), .B(new_n4640_), .C(new_n4636_), .D(new_n4639_), .Y(new_n4647_));
  OAI211 g03645(.A0(new_n4646_), .A1(new_n4639_), .B0(new_n4647_), .B1(new_n2925_), .Y(new_n4648_));
  OAI21  g03646(.A0(new_n4637_), .A1(new_n4643_), .B0(new_n4648_), .Y(new_n4649_));
  NAND2  g03647(.A(new_n4649_), .B(new_n4615_), .Y(new_n4650_));
  OAI21  g03648(.A0(new_n4638_), .A1(new_n4615_), .B0(new_n4650_), .Y(new_n4651_));
  XOR2   g03649(.A(new_n2960_), .B(new_n2953_), .Y(new_n4652_));
  XOR2   g03650(.A(\A[479] ), .B(new_n2957_), .Y(new_n4653_));
  NAND2  g03651(.A(\A[479] ), .B(\A[478] ), .Y(new_n4654_));
  OAI21  g03652(.A0(new_n4653_), .A1(new_n2954_), .B0(new_n4654_), .Y(new_n4655_));
  XOR2   g03653(.A(new_n2964_), .B(new_n4655_), .Y(new_n4656_));
  NOR2   g03654(.A(\A[476] ), .B(new_n2950_), .Y(new_n4657_));
  OAI21  g03655(.A0(new_n2948_), .A1(\A[475] ), .B0(\A[477] ), .Y(new_n4658_));
  XOR2   g03656(.A(\A[476] ), .B(new_n2950_), .Y(new_n4659_));
  OAI22  g03657(.A0(new_n4659_), .A1(\A[477] ), .B0(new_n4658_), .B1(new_n4657_), .Y(new_n4660_));
  NOR2   g03658(.A(\A[479] ), .B(new_n2957_), .Y(new_n4661_));
  OAI21  g03659(.A0(new_n2955_), .A1(\A[478] ), .B0(\A[480] ), .Y(new_n4662_));
  OAI22  g03660(.A0(new_n4653_), .A1(\A[480] ), .B0(new_n4662_), .B1(new_n4661_), .Y(new_n4663_));
  NAND2  g03661(.A(new_n4663_), .B(new_n4660_), .Y(new_n4664_));
  NAND2  g03662(.A(\A[476] ), .B(\A[475] ), .Y(new_n4665_));
  OAI21  g03663(.A0(new_n4659_), .A1(new_n2947_), .B0(new_n4665_), .Y(new_n4666_));
  NAND2  g03664(.A(new_n4666_), .B(new_n4655_), .Y(new_n4667_));
  OAI21  g03665(.A0(new_n4664_), .A1(new_n4656_), .B0(new_n4667_), .Y(new_n4668_));
  NOR2   g03666(.A(new_n2960_), .B(new_n2953_), .Y(new_n4669_));
  XOR2   g03667(.A(new_n4669_), .B(new_n4656_), .Y(new_n4670_));
  AOI21  g03668(.A0(new_n4668_), .A1(new_n4652_), .B0(new_n4670_), .Y(new_n4671_));
  XOR2   g03669(.A(new_n2941_), .B(new_n2934_), .Y(new_n4672_));
  NOR2   g03670(.A(\A[482] ), .B(new_n2931_), .Y(new_n4673_));
  OAI21  g03671(.A0(new_n2929_), .A1(\A[481] ), .B0(\A[483] ), .Y(new_n4674_));
  NAND2  g03672(.A(new_n2933_), .B(new_n2928_), .Y(new_n4675_));
  OAI21  g03673(.A0(new_n4674_), .A1(new_n4673_), .B0(new_n4675_), .Y(new_n4676_));
  NOR2   g03674(.A(\A[485] ), .B(new_n2938_), .Y(new_n4677_));
  OAI21  g03675(.A0(new_n2936_), .A1(\A[484] ), .B0(\A[486] ), .Y(new_n4678_));
  NAND2  g03676(.A(new_n2940_), .B(new_n2935_), .Y(new_n4679_));
  OAI21  g03677(.A0(new_n4678_), .A1(new_n4677_), .B0(new_n4679_), .Y(new_n4680_));
  NAND2  g03678(.A(new_n2940_), .B(\A[486] ), .Y(new_n4681_));
  OAI21  g03679(.A0(new_n2936_), .A1(new_n2938_), .B0(new_n4681_), .Y(new_n4682_));
  NAND2  g03680(.A(new_n2933_), .B(\A[483] ), .Y(new_n4683_));
  OAI21  g03681(.A0(new_n2929_), .A1(new_n2931_), .B0(new_n4683_), .Y(new_n4684_));
  NAND4  g03682(.A(new_n4684_), .B(new_n4682_), .C(new_n4680_), .D(new_n4676_), .Y(new_n4685_));
  NAND4  g03683(.A(new_n4666_), .B(new_n4655_), .C(new_n4663_), .D(new_n4660_), .Y(new_n4686_));
  NAND4  g03684(.A(new_n4686_), .B(new_n4652_), .C(new_n4685_), .D(new_n4672_), .Y(new_n4687_));
  XOR2   g03685(.A(new_n2945_), .B(new_n4682_), .Y(new_n4688_));
  NAND2  g03686(.A(new_n4680_), .B(new_n4676_), .Y(new_n4689_));
  NAND2  g03687(.A(new_n4684_), .B(new_n4682_), .Y(new_n4690_));
  OAI21  g03688(.A0(new_n4689_), .A1(new_n4688_), .B0(new_n4690_), .Y(new_n4691_));
  NOR2   g03689(.A(new_n2941_), .B(new_n2934_), .Y(new_n4692_));
  XOR2   g03690(.A(new_n4692_), .B(new_n4688_), .Y(new_n4693_));
  AOI21  g03691(.A0(new_n4691_), .A1(new_n4672_), .B0(new_n4693_), .Y(new_n4694_));
  XOR2   g03692(.A(new_n4694_), .B(new_n4687_), .Y(new_n4695_));
  NOR2   g03693(.A(new_n4695_), .B(new_n4671_), .Y(new_n4696_));
  XOR2   g03694(.A(new_n2960_), .B(new_n4660_), .Y(new_n4697_));
  XOR2   g03695(.A(new_n2964_), .B(new_n2962_), .Y(new_n4698_));
  NOR2   g03696(.A(new_n2964_), .B(new_n2962_), .Y(new_n4699_));
  AOI21  g03697(.A0(new_n4669_), .A1(new_n4698_), .B0(new_n4699_), .Y(new_n4700_));
  XOR2   g03698(.A(new_n4669_), .B(new_n4698_), .Y(new_n4701_));
  OAI21  g03699(.A0(new_n4700_), .A1(new_n4697_), .B0(new_n4701_), .Y(new_n4702_));
  XOR2   g03700(.A(new_n2941_), .B(new_n4676_), .Y(new_n4703_));
  XOR2   g03701(.A(new_n2945_), .B(new_n2943_), .Y(new_n4704_));
  NOR2   g03702(.A(new_n2945_), .B(new_n2943_), .Y(new_n4705_));
  AOI21  g03703(.A0(new_n4692_), .A1(new_n4704_), .B0(new_n4705_), .Y(new_n4706_));
  XOR2   g03704(.A(new_n4692_), .B(new_n4704_), .Y(new_n4707_));
  OAI21  g03705(.A0(new_n4706_), .A1(new_n4703_), .B0(new_n4707_), .Y(new_n4708_));
  NAND2  g03706(.A(new_n4708_), .B(new_n4687_), .Y(new_n4709_));
  NOR4   g03707(.A(new_n2945_), .B(new_n2943_), .C(new_n2941_), .D(new_n2934_), .Y(new_n4710_));
  NOR4   g03708(.A(new_n4697_), .B(new_n4710_), .C(new_n4693_), .D(new_n4703_), .Y(new_n4711_));
  OAI211 g03709(.A0(new_n4706_), .A1(new_n4703_), .B0(new_n4711_), .B1(new_n4686_), .Y(new_n4712_));
  AOI21  g03710(.A0(new_n4712_), .A1(new_n4709_), .B0(new_n4702_), .Y(new_n4713_));
  NAND2  g03711(.A(new_n2966_), .B(new_n2927_), .Y(new_n4714_));
  NOR3   g03712(.A(new_n4714_), .B(new_n4713_), .C(new_n4696_), .Y(new_n4715_));
  NOR4   g03713(.A(new_n2964_), .B(new_n2962_), .C(new_n2960_), .D(new_n2953_), .Y(new_n4716_));
  NOR4   g03714(.A(new_n4716_), .B(new_n4697_), .C(new_n4710_), .D(new_n4703_), .Y(new_n4717_));
  XOR2   g03715(.A(new_n4694_), .B(new_n4717_), .Y(new_n4718_));
  NAND2  g03716(.A(new_n4718_), .B(new_n4702_), .Y(new_n4719_));
  NAND4  g03717(.A(new_n4652_), .B(new_n4685_), .C(new_n4707_), .D(new_n4672_), .Y(new_n4720_));
  OAI21  g03718(.A0(new_n4706_), .A1(new_n4703_), .B0(new_n4686_), .Y(new_n4721_));
  OAI22  g03719(.A0(new_n4721_), .A1(new_n4720_), .B0(new_n4694_), .B1(new_n4717_), .Y(new_n4722_));
  NAND2  g03720(.A(new_n4722_), .B(new_n4671_), .Y(new_n4723_));
  XOR2   g03721(.A(new_n2926_), .B(new_n2895_), .Y(new_n4724_));
  NOR2   g03722(.A(new_n2967_), .B(new_n4724_), .Y(new_n4725_));
  AOI21  g03723(.A0(new_n4723_), .A1(new_n4719_), .B0(new_n4725_), .Y(new_n4726_));
  NOR2   g03724(.A(new_n4726_), .B(new_n4715_), .Y(new_n4727_));
  NOR2   g03725(.A(new_n4651_), .B(new_n4727_), .Y(new_n4728_));
  NOR2   g03726(.A(new_n4713_), .B(new_n4696_), .Y(new_n4729_));
  NAND3  g03727(.A(new_n4714_), .B(new_n4723_), .C(new_n4719_), .Y(new_n4730_));
  OAI21  g03728(.A0(new_n4729_), .A1(new_n4714_), .B0(new_n4730_), .Y(new_n4731_));
  AOI21  g03729(.A0(new_n4731_), .A1(new_n4651_), .B0(new_n4728_), .Y(new_n4732_));
  AOI21  g03730(.A0(new_n4585_), .A1(new_n4576_), .B0(new_n4597_), .Y(new_n4733_));
  OAI21  g03731(.A0(new_n4733_), .A1(new_n4588_), .B0(new_n4589_), .Y(new_n4734_));
  NAND2  g03732(.A(new_n4734_), .B(new_n4594_), .Y(new_n4735_));
  NAND3  g03733(.A(new_n4587_), .B(new_n4586_), .C(new_n4561_), .Y(new_n4736_));
  OAI21  g03734(.A0(new_n4733_), .A1(new_n4587_), .B0(new_n4736_), .Y(new_n4737_));
  AOI21  g03735(.A0(new_n4737_), .A1(new_n4524_), .B0(new_n4601_), .Y(new_n4738_));
  NAND2  g03736(.A(new_n4738_), .B(new_n4735_), .Y(new_n4739_));
  OAI21  g03737(.A0(new_n4603_), .A1(new_n4592_), .B0(new_n4601_), .Y(new_n4740_));
  AOI21  g03738(.A0(new_n4740_), .A1(new_n4739_), .B0(new_n4732_), .Y(new_n4741_));
  AOI21  g03739(.A0(new_n4732_), .A1(new_n4606_), .B0(new_n4741_), .Y(new_n4742_));
  OAI21  g03740(.A0(new_n4467_), .A1(new_n4460_), .B0(new_n4742_), .Y(new_n4743_));
  NOR2   g03741(.A(new_n4602_), .B(new_n4592_), .Y(new_n4744_));
  NAND2  g03742(.A(new_n4737_), .B(new_n4524_), .Y(new_n4745_));
  AOI21  g03743(.A0(new_n4745_), .A1(new_n4735_), .B0(new_n4601_), .Y(new_n4746_));
  OAI21  g03744(.A0(new_n4746_), .A1(new_n4744_), .B0(new_n4732_), .Y(new_n4747_));
  NOR3   g03745(.A(new_n4601_), .B(new_n4603_), .C(new_n4592_), .Y(new_n4748_));
  AOI21  g03746(.A0(new_n4745_), .A1(new_n4735_), .B0(new_n4604_), .Y(new_n4749_));
  NOR2   g03747(.A(new_n4749_), .B(new_n4748_), .Y(new_n4750_));
  OAI21  g03748(.A0(new_n4750_), .A1(new_n4732_), .B0(new_n4747_), .Y(new_n4751_));
  NOR3   g03749(.A(new_n4458_), .B(new_n4457_), .C(new_n4442_), .Y(new_n4752_));
  AOI21  g03750(.A0(new_n4466_), .A1(new_n4463_), .B0(new_n4459_), .Y(new_n4753_));
  OAI21  g03751(.A0(new_n4753_), .A1(new_n4752_), .B0(new_n4751_), .Y(new_n4754_));
  NAND2  g03752(.A(new_n4754_), .B(new_n4743_), .Y(new_n4755_));
  AOI21  g03753(.A0(new_n4166_), .A1(new_n4158_), .B0(new_n4755_), .Y(new_n4756_));
  NAND3  g03754(.A(new_n4458_), .B(new_n4466_), .C(new_n4463_), .Y(new_n4757_));
  OAI21  g03755(.A0(new_n4457_), .A1(new_n4442_), .B0(new_n4459_), .Y(new_n4758_));
  AOI21  g03756(.A0(new_n4758_), .A1(new_n4757_), .B0(new_n4751_), .Y(new_n4759_));
  NAND3  g03757(.A(new_n4459_), .B(new_n4466_), .C(new_n4463_), .Y(new_n4760_));
  OAI21  g03758(.A0(new_n4457_), .A1(new_n4442_), .B0(new_n4458_), .Y(new_n4761_));
  AOI21  g03759(.A0(new_n4761_), .A1(new_n4760_), .B0(new_n4742_), .Y(new_n4762_));
  NOR2   g03760(.A(new_n4762_), .B(new_n4759_), .Y(new_n4763_));
  NAND3  g03761(.A(new_n4165_), .B(new_n4156_), .C(new_n4145_), .Y(new_n4764_));
  OAI21  g03762(.A0(new_n4164_), .A1(new_n4161_), .B0(new_n4157_), .Y(new_n4765_));
  AOI21  g03763(.A0(new_n4765_), .A1(new_n4764_), .B0(new_n4763_), .Y(new_n4766_));
  NOR2   g03764(.A(new_n4766_), .B(new_n4756_), .Y(new_n4767_));
  NAND3  g03765(.A(new_n3555_), .B(new_n2876_), .C(new_n2866_), .Y(new_n4768_));
  OAI21  g03766(.A0(new_n3554_), .A1(new_n3551_), .B0(new_n3547_), .Y(new_n4769_));
  AOI21  g03767(.A0(new_n4769_), .A1(new_n4768_), .B0(new_n4767_), .Y(new_n4770_));
  AOI21  g03768(.A0(new_n4767_), .A1(new_n3557_), .B0(new_n4770_), .Y(new_n4771_));
  INV    g03769(.A(\A[969] ), .Y(new_n4772_));
  INV    g03770(.A(\A[967] ), .Y(new_n4773_));
  NAND2  g03771(.A(\A[968] ), .B(new_n4773_), .Y(new_n4774_));
  INV    g03772(.A(\A[968] ), .Y(new_n4775_));
  AOI21  g03773(.A0(new_n4775_), .A1(\A[967] ), .B0(new_n4772_), .Y(new_n4776_));
  XOR2   g03774(.A(\A[968] ), .B(\A[967] ), .Y(new_n4777_));
  AOI22  g03775(.A0(new_n4777_), .A1(new_n4772_), .B0(new_n4776_), .B1(new_n4774_), .Y(new_n4778_));
  INV    g03776(.A(\A[972] ), .Y(new_n4779_));
  INV    g03777(.A(\A[970] ), .Y(new_n4780_));
  NAND2  g03778(.A(\A[971] ), .B(new_n4780_), .Y(new_n4781_));
  INV    g03779(.A(\A[971] ), .Y(new_n4782_));
  AOI21  g03780(.A0(new_n4782_), .A1(\A[970] ), .B0(new_n4779_), .Y(new_n4783_));
  XOR2   g03781(.A(\A[971] ), .B(\A[970] ), .Y(new_n4784_));
  AOI22  g03782(.A0(new_n4784_), .A1(new_n4779_), .B0(new_n4783_), .B1(new_n4781_), .Y(new_n4785_));
  NOR2   g03783(.A(new_n4785_), .B(new_n4778_), .Y(new_n4786_));
  NOR2   g03784(.A(new_n4782_), .B(new_n4780_), .Y(new_n4787_));
  AOI21  g03785(.A0(new_n4784_), .A1(\A[972] ), .B0(new_n4787_), .Y(new_n4788_));
  NOR2   g03786(.A(new_n4775_), .B(new_n4773_), .Y(new_n4789_));
  AOI21  g03787(.A0(new_n4777_), .A1(\A[969] ), .B0(new_n4789_), .Y(new_n4790_));
  XOR2   g03788(.A(new_n4790_), .B(new_n4788_), .Y(new_n4791_));
  XOR2   g03789(.A(new_n4791_), .B(new_n4786_), .Y(new_n4792_));
  NAND2  g03790(.A(new_n4776_), .B(new_n4774_), .Y(new_n4793_));
  INV    g03791(.A(new_n4777_), .Y(new_n4794_));
  OAI21  g03792(.A0(new_n4794_), .A1(\A[969] ), .B0(new_n4793_), .Y(new_n4795_));
  XOR2   g03793(.A(new_n4785_), .B(new_n4795_), .Y(new_n4796_));
  NOR2   g03794(.A(new_n4790_), .B(new_n4788_), .Y(new_n4797_));
  AOI21  g03795(.A0(new_n4791_), .A1(new_n4786_), .B0(new_n4797_), .Y(new_n4798_));
  OAI21  g03796(.A0(new_n4798_), .A1(new_n4796_), .B0(new_n4792_), .Y(new_n4799_));
  NAND2  g03797(.A(\A[977] ), .B(\A[976] ), .Y(new_n4800_));
  XOR2   g03798(.A(\A[977] ), .B(\A[976] ), .Y(new_n4801_));
  NAND2  g03799(.A(new_n4801_), .B(\A[978] ), .Y(new_n4802_));
  NAND2  g03800(.A(new_n4802_), .B(new_n4800_), .Y(new_n4803_));
  INV    g03801(.A(\A[973] ), .Y(new_n4804_));
  INV    g03802(.A(\A[974] ), .Y(new_n4805_));
  NOR2   g03803(.A(new_n4805_), .B(new_n4804_), .Y(new_n4806_));
  XOR2   g03804(.A(\A[974] ), .B(\A[973] ), .Y(new_n4807_));
  AOI21  g03805(.A0(new_n4807_), .A1(\A[975] ), .B0(new_n4806_), .Y(new_n4808_));
  XOR2   g03806(.A(new_n4808_), .B(new_n4803_), .Y(new_n4809_));
  NOR2   g03807(.A(new_n4805_), .B(\A[973] ), .Y(new_n4810_));
  OAI21  g03808(.A0(\A[974] ), .A1(new_n4804_), .B0(\A[975] ), .Y(new_n4811_));
  INV    g03809(.A(\A[975] ), .Y(new_n4812_));
  NAND2  g03810(.A(new_n4807_), .B(new_n4812_), .Y(new_n4813_));
  OAI21  g03811(.A0(new_n4811_), .A1(new_n4810_), .B0(new_n4813_), .Y(new_n4814_));
  INV    g03812(.A(\A[977] ), .Y(new_n4815_));
  NOR2   g03813(.A(new_n4815_), .B(\A[976] ), .Y(new_n4816_));
  INV    g03814(.A(\A[976] ), .Y(new_n4817_));
  OAI21  g03815(.A0(\A[977] ), .A1(new_n4817_), .B0(\A[978] ), .Y(new_n4818_));
  INV    g03816(.A(\A[978] ), .Y(new_n4819_));
  NAND2  g03817(.A(new_n4801_), .B(new_n4819_), .Y(new_n4820_));
  OAI21  g03818(.A0(new_n4818_), .A1(new_n4816_), .B0(new_n4820_), .Y(new_n4821_));
  NAND2  g03819(.A(new_n4821_), .B(new_n4814_), .Y(new_n4822_));
  NAND2  g03820(.A(new_n4807_), .B(\A[975] ), .Y(new_n4823_));
  OAI21  g03821(.A0(new_n4805_), .A1(new_n4804_), .B0(new_n4823_), .Y(new_n4824_));
  NAND2  g03822(.A(new_n4824_), .B(new_n4803_), .Y(new_n4825_));
  OAI21  g03823(.A0(new_n4822_), .A1(new_n4809_), .B0(new_n4825_), .Y(new_n4826_));
  XOR2   g03824(.A(new_n4824_), .B(new_n4803_), .Y(new_n4827_));
  NAND2  g03825(.A(\A[974] ), .B(new_n4804_), .Y(new_n4828_));
  AOI21  g03826(.A0(new_n4805_), .A1(\A[973] ), .B0(new_n4812_), .Y(new_n4829_));
  AOI22  g03827(.A0(new_n4829_), .A1(new_n4828_), .B0(new_n4807_), .B1(new_n4812_), .Y(new_n4830_));
  NAND2  g03828(.A(\A[977] ), .B(new_n4817_), .Y(new_n4831_));
  AOI21  g03829(.A0(new_n4815_), .A1(\A[976] ), .B0(new_n4819_), .Y(new_n4832_));
  AOI22  g03830(.A0(new_n4832_), .A1(new_n4831_), .B0(new_n4801_), .B1(new_n4819_), .Y(new_n4833_));
  NOR2   g03831(.A(new_n4833_), .B(new_n4830_), .Y(new_n4834_));
  XOR2   g03832(.A(new_n4834_), .B(new_n4827_), .Y(new_n4835_));
  NOR4   g03833(.A(new_n4790_), .B(new_n4788_), .C(new_n4785_), .D(new_n4778_), .Y(new_n4836_));
  XOR2   g03834(.A(new_n4785_), .B(new_n4778_), .Y(new_n4837_));
  XOR2   g03835(.A(new_n4833_), .B(new_n4830_), .Y(new_n4838_));
  NAND2  g03836(.A(new_n4838_), .B(new_n4837_), .Y(new_n4839_));
  AOI211 g03837(.A0(new_n4835_), .A1(new_n4826_), .B(new_n4839_), .C(new_n4836_), .Y(new_n4840_));
  XOR2   g03838(.A(new_n4834_), .B(new_n4809_), .Y(new_n4841_));
  AOI21  g03839(.A0(new_n4838_), .A1(new_n4826_), .B0(new_n4841_), .Y(new_n4842_));
  XOR2   g03840(.A(new_n4842_), .B(new_n4840_), .Y(new_n4843_));
  NAND2  g03841(.A(new_n4843_), .B(new_n4799_), .Y(new_n4844_));
  NAND4  g03842(.A(new_n4821_), .B(new_n4814_), .C(new_n4824_), .D(new_n4803_), .Y(new_n4845_));
  NAND2  g03843(.A(new_n4784_), .B(\A[972] ), .Y(new_n4846_));
  OAI21  g03844(.A0(new_n4782_), .A1(new_n4780_), .B0(new_n4846_), .Y(new_n4847_));
  NOR2   g03845(.A(new_n4794_), .B(new_n4772_), .Y(new_n4848_));
  OAI211 g03846(.A0(new_n4848_), .A1(new_n4789_), .B0(new_n4847_), .B1(new_n4786_), .Y(new_n4849_));
  NAND4  g03847(.A(new_n4838_), .B(new_n4849_), .C(new_n4845_), .D(new_n4837_), .Y(new_n4850_));
  AOI21  g03848(.A0(new_n4802_), .A1(new_n4800_), .B0(new_n4808_), .Y(new_n4851_));
  AOI21  g03849(.A0(new_n4834_), .A1(new_n4827_), .B0(new_n4851_), .Y(new_n4852_));
  XOR2   g03850(.A(new_n4833_), .B(new_n4814_), .Y(new_n4853_));
  OAI21  g03851(.A0(new_n4853_), .A1(new_n4852_), .B0(new_n4835_), .Y(new_n4854_));
  AOI221 g03852(.A0(new_n4833_), .A1(new_n4830_), .C0(new_n4808_), .B0(new_n4802_), .B1(new_n4800_), .Y(new_n4855_));
  NOR4   g03853(.A(new_n4855_), .B(new_n4839_), .C(new_n4836_), .D(new_n4841_), .Y(new_n4856_));
  AOI21  g03854(.A0(new_n4854_), .A1(new_n4850_), .B0(new_n4856_), .Y(new_n4857_));
  OAI21  g03855(.A0(new_n4857_), .A1(new_n4799_), .B0(new_n4844_), .Y(new_n4858_));
  INV    g03856(.A(\A[981] ), .Y(new_n4859_));
  INV    g03857(.A(\A[979] ), .Y(new_n4860_));
  NAND2  g03858(.A(\A[980] ), .B(new_n4860_), .Y(new_n4861_));
  INV    g03859(.A(\A[980] ), .Y(new_n4862_));
  AOI21  g03860(.A0(new_n4862_), .A1(\A[979] ), .B0(new_n4859_), .Y(new_n4863_));
  XOR2   g03861(.A(\A[980] ), .B(\A[979] ), .Y(new_n4864_));
  AOI22  g03862(.A0(new_n4864_), .A1(new_n4859_), .B0(new_n4863_), .B1(new_n4861_), .Y(new_n4865_));
  INV    g03863(.A(\A[984] ), .Y(new_n4866_));
  INV    g03864(.A(\A[982] ), .Y(new_n4867_));
  NAND2  g03865(.A(\A[983] ), .B(new_n4867_), .Y(new_n4868_));
  INV    g03866(.A(\A[983] ), .Y(new_n4869_));
  AOI21  g03867(.A0(new_n4869_), .A1(\A[982] ), .B0(new_n4866_), .Y(new_n4870_));
  XOR2   g03868(.A(\A[983] ), .B(\A[982] ), .Y(new_n4871_));
  AOI22  g03869(.A0(new_n4871_), .A1(new_n4866_), .B0(new_n4870_), .B1(new_n4868_), .Y(new_n4872_));
  NOR2   g03870(.A(new_n4872_), .B(new_n4865_), .Y(new_n4873_));
  NOR2   g03871(.A(new_n4869_), .B(new_n4867_), .Y(new_n4874_));
  AOI21  g03872(.A0(new_n4871_), .A1(\A[984] ), .B0(new_n4874_), .Y(new_n4875_));
  NOR2   g03873(.A(new_n4862_), .B(new_n4860_), .Y(new_n4876_));
  AOI21  g03874(.A0(new_n4864_), .A1(\A[981] ), .B0(new_n4876_), .Y(new_n4877_));
  XOR2   g03875(.A(new_n4877_), .B(new_n4875_), .Y(new_n4878_));
  XOR2   g03876(.A(new_n4878_), .B(new_n4873_), .Y(new_n4879_));
  NOR2   g03877(.A(new_n4862_), .B(\A[979] ), .Y(new_n4880_));
  OAI21  g03878(.A0(\A[980] ), .A1(new_n4860_), .B0(\A[981] ), .Y(new_n4881_));
  XOR2   g03879(.A(\A[980] ), .B(new_n4860_), .Y(new_n4882_));
  OAI22  g03880(.A0(new_n4882_), .A1(\A[981] ), .B0(new_n4881_), .B1(new_n4880_), .Y(new_n4883_));
  XOR2   g03881(.A(new_n4872_), .B(new_n4883_), .Y(new_n4884_));
  NOR2   g03882(.A(new_n4877_), .B(new_n4875_), .Y(new_n4885_));
  AOI21  g03883(.A0(new_n4878_), .A1(new_n4873_), .B0(new_n4885_), .Y(new_n4886_));
  OAI21  g03884(.A0(new_n4886_), .A1(new_n4884_), .B0(new_n4879_), .Y(new_n4887_));
  INV    g03885(.A(\A[988] ), .Y(new_n4888_));
  INV    g03886(.A(\A[989] ), .Y(new_n4889_));
  NOR2   g03887(.A(new_n4889_), .B(new_n4888_), .Y(new_n4890_));
  XOR2   g03888(.A(\A[989] ), .B(\A[988] ), .Y(new_n4891_));
  AOI21  g03889(.A0(new_n4891_), .A1(\A[990] ), .B0(new_n4890_), .Y(new_n4892_));
  INV    g03890(.A(\A[985] ), .Y(new_n4893_));
  INV    g03891(.A(\A[986] ), .Y(new_n4894_));
  NOR2   g03892(.A(new_n4894_), .B(new_n4893_), .Y(new_n4895_));
  XOR2   g03893(.A(\A[986] ), .B(\A[985] ), .Y(new_n4896_));
  AOI21  g03894(.A0(new_n4896_), .A1(\A[987] ), .B0(new_n4895_), .Y(new_n4897_));
  INV    g03895(.A(\A[987] ), .Y(new_n4898_));
  NAND2  g03896(.A(\A[986] ), .B(new_n4893_), .Y(new_n4899_));
  AOI21  g03897(.A0(new_n4894_), .A1(\A[985] ), .B0(new_n4898_), .Y(new_n4900_));
  AOI22  g03898(.A0(new_n4900_), .A1(new_n4899_), .B0(new_n4896_), .B1(new_n4898_), .Y(new_n4901_));
  INV    g03899(.A(\A[990] ), .Y(new_n4902_));
  NAND2  g03900(.A(\A[989] ), .B(new_n4888_), .Y(new_n4903_));
  AOI21  g03901(.A0(new_n4889_), .A1(\A[988] ), .B0(new_n4902_), .Y(new_n4904_));
  AOI22  g03902(.A0(new_n4904_), .A1(new_n4903_), .B0(new_n4891_), .B1(new_n4902_), .Y(new_n4905_));
  NOR4   g03903(.A(new_n4905_), .B(new_n4901_), .C(new_n4897_), .D(new_n4892_), .Y(new_n4906_));
  NOR4   g03904(.A(new_n4877_), .B(new_n4875_), .C(new_n4872_), .D(new_n4865_), .Y(new_n4907_));
  NOR2   g03905(.A(new_n4894_), .B(\A[985] ), .Y(new_n4908_));
  OAI21  g03906(.A0(\A[986] ), .A1(new_n4893_), .B0(\A[987] ), .Y(new_n4909_));
  NAND2  g03907(.A(new_n4896_), .B(new_n4898_), .Y(new_n4910_));
  OAI21  g03908(.A0(new_n4909_), .A1(new_n4908_), .B0(new_n4910_), .Y(new_n4911_));
  XOR2   g03909(.A(new_n4905_), .B(new_n4911_), .Y(new_n4912_));
  NOR4   g03910(.A(new_n4912_), .B(new_n4907_), .C(new_n4906_), .D(new_n4884_), .Y(new_n4913_));
  NAND2  g03911(.A(new_n4891_), .B(\A[990] ), .Y(new_n4914_));
  OAI21  g03912(.A0(new_n4889_), .A1(new_n4888_), .B0(new_n4914_), .Y(new_n4915_));
  XOR2   g03913(.A(new_n4897_), .B(new_n4915_), .Y(new_n4916_));
  NOR2   g03914(.A(new_n4889_), .B(\A[988] ), .Y(new_n4917_));
  OAI21  g03915(.A0(\A[989] ), .A1(new_n4888_), .B0(\A[990] ), .Y(new_n4918_));
  NAND2  g03916(.A(new_n4891_), .B(new_n4902_), .Y(new_n4919_));
  OAI21  g03917(.A0(new_n4918_), .A1(new_n4917_), .B0(new_n4919_), .Y(new_n4920_));
  NAND2  g03918(.A(new_n4920_), .B(new_n4911_), .Y(new_n4921_));
  NAND2  g03919(.A(new_n4896_), .B(\A[987] ), .Y(new_n4922_));
  OAI21  g03920(.A0(new_n4894_), .A1(new_n4893_), .B0(new_n4922_), .Y(new_n4923_));
  NAND2  g03921(.A(new_n4923_), .B(new_n4915_), .Y(new_n4924_));
  OAI21  g03922(.A0(new_n4921_), .A1(new_n4916_), .B0(new_n4924_), .Y(new_n4925_));
  NOR2   g03923(.A(new_n4905_), .B(new_n4901_), .Y(new_n4926_));
  XOR2   g03924(.A(new_n4926_), .B(new_n4916_), .Y(new_n4927_));
  XOR2   g03925(.A(new_n4905_), .B(new_n4901_), .Y(new_n4928_));
  AOI21  g03926(.A0(new_n4928_), .A1(new_n4925_), .B0(new_n4927_), .Y(new_n4929_));
  XOR2   g03927(.A(new_n4929_), .B(new_n4913_), .Y(new_n4930_));
  NAND2  g03928(.A(new_n4930_), .B(new_n4887_), .Y(new_n4931_));
  INV    g03929(.A(new_n4871_), .Y(new_n4932_));
  NAND2  g03930(.A(\A[983] ), .B(\A[982] ), .Y(new_n4933_));
  OAI21  g03931(.A0(new_n4932_), .A1(new_n4866_), .B0(new_n4933_), .Y(new_n4934_));
  XOR2   g03932(.A(new_n4877_), .B(new_n4934_), .Y(new_n4935_));
  XOR2   g03933(.A(new_n4935_), .B(new_n4873_), .Y(new_n4936_));
  INV    g03934(.A(new_n4884_), .Y(new_n4937_));
  NAND2  g03935(.A(new_n4878_), .B(new_n4873_), .Y(new_n4938_));
  OAI21  g03936(.A0(new_n4877_), .A1(new_n4875_), .B0(new_n4938_), .Y(new_n4939_));
  AOI21  g03937(.A0(new_n4939_), .A1(new_n4937_), .B0(new_n4936_), .Y(new_n4940_));
  XOR2   g03938(.A(new_n4923_), .B(new_n4915_), .Y(new_n4941_));
  XOR2   g03939(.A(new_n4926_), .B(new_n4941_), .Y(new_n4942_));
  NOR2   g03940(.A(new_n4882_), .B(new_n4859_), .Y(new_n4943_));
  OAI211 g03941(.A0(new_n4943_), .A1(new_n4876_), .B0(new_n4934_), .B1(new_n4873_), .Y(new_n4944_));
  NOR2   g03942(.A(new_n4912_), .B(new_n4884_), .Y(new_n4945_));
  OAI211 g03943(.A0(new_n4920_), .A1(new_n4911_), .B0(new_n4923_), .B1(new_n4915_), .Y(new_n4946_));
  NAND4  g03944(.A(new_n4946_), .B(new_n4945_), .C(new_n4944_), .D(new_n4942_), .Y(new_n4947_));
  OAI21  g03945(.A0(new_n4929_), .A1(new_n4913_), .B0(new_n4947_), .Y(new_n4948_));
  NAND2  g03946(.A(new_n4948_), .B(new_n4940_), .Y(new_n4949_));
  NAND4  g03947(.A(new_n4920_), .B(new_n4911_), .C(new_n4923_), .D(new_n4915_), .Y(new_n4950_));
  NAND2  g03948(.A(new_n4928_), .B(new_n4950_), .Y(new_n4951_));
  XOR2   g03949(.A(new_n4872_), .B(new_n4865_), .Y(new_n4952_));
  XOR2   g03950(.A(new_n4952_), .B(new_n4951_), .Y(new_n4953_));
  NAND2  g03951(.A(new_n4838_), .B(new_n4845_), .Y(new_n4954_));
  XOR2   g03952(.A(new_n4785_), .B(new_n4778_), .Y(new_n4955_));
  XOR2   g03953(.A(new_n4955_), .B(new_n4954_), .Y(new_n4956_));
  NOR2   g03954(.A(new_n4956_), .B(new_n4953_), .Y(new_n4957_));
  NAND3  g03955(.A(new_n4957_), .B(new_n4949_), .C(new_n4931_), .Y(new_n4958_));
  NAND3  g03956(.A(new_n4945_), .B(new_n4944_), .C(new_n4950_), .Y(new_n4959_));
  XOR2   g03957(.A(new_n4929_), .B(new_n4959_), .Y(new_n4960_));
  NOR2   g03958(.A(new_n4960_), .B(new_n4940_), .Y(new_n4961_));
  NOR2   g03959(.A(new_n4897_), .B(new_n4892_), .Y(new_n4962_));
  AOI21  g03960(.A0(new_n4926_), .A1(new_n4941_), .B0(new_n4962_), .Y(new_n4963_));
  OAI21  g03961(.A0(new_n4912_), .A1(new_n4963_), .B0(new_n4942_), .Y(new_n4964_));
  NAND2  g03962(.A(new_n4964_), .B(new_n4959_), .Y(new_n4965_));
  AOI21  g03963(.A0(new_n4947_), .A1(new_n4965_), .B0(new_n4887_), .Y(new_n4966_));
  NOR2   g03964(.A(new_n4912_), .B(new_n4906_), .Y(new_n4967_));
  XOR2   g03965(.A(new_n4952_), .B(new_n4967_), .Y(new_n4968_));
  INV    g03966(.A(new_n4955_), .Y(new_n4969_));
  XOR2   g03967(.A(new_n4969_), .B(new_n4954_), .Y(new_n4970_));
  NAND2  g03968(.A(new_n4970_), .B(new_n4968_), .Y(new_n4971_));
  OAI21  g03969(.A0(new_n4966_), .A1(new_n4961_), .B0(new_n4971_), .Y(new_n4972_));
  AOI21  g03970(.A0(new_n4972_), .A1(new_n4958_), .B0(new_n4858_), .Y(new_n4973_));
  XOR2   g03971(.A(new_n4956_), .B(new_n4968_), .Y(new_n4974_));
  INV    g03972(.A(\A[963] ), .Y(new_n4975_));
  INV    g03973(.A(\A[962] ), .Y(new_n4976_));
  NAND2  g03974(.A(new_n4976_), .B(\A[961] ), .Y(new_n4977_));
  INV    g03975(.A(\A[961] ), .Y(new_n4978_));
  AOI21  g03976(.A0(\A[962] ), .A1(new_n4978_), .B0(new_n4975_), .Y(new_n4979_));
  XOR2   g03977(.A(\A[962] ), .B(\A[961] ), .Y(new_n4980_));
  AOI22  g03978(.A0(new_n4980_), .A1(new_n4975_), .B0(new_n4979_), .B1(new_n4977_), .Y(new_n4981_));
  INV    g03979(.A(\A[966] ), .Y(new_n4982_));
  INV    g03980(.A(\A[965] ), .Y(new_n4983_));
  NAND2  g03981(.A(new_n4983_), .B(\A[964] ), .Y(new_n4984_));
  INV    g03982(.A(\A[964] ), .Y(new_n4985_));
  AOI21  g03983(.A0(\A[965] ), .A1(new_n4985_), .B0(new_n4982_), .Y(new_n4986_));
  XOR2   g03984(.A(\A[965] ), .B(\A[964] ), .Y(new_n4987_));
  AOI22  g03985(.A0(new_n4987_), .A1(new_n4982_), .B0(new_n4986_), .B1(new_n4984_), .Y(new_n4988_));
  NOR2   g03986(.A(new_n4983_), .B(new_n4985_), .Y(new_n4989_));
  AOI21  g03987(.A0(new_n4987_), .A1(\A[966] ), .B0(new_n4989_), .Y(new_n4990_));
  NOR2   g03988(.A(new_n4976_), .B(new_n4978_), .Y(new_n4991_));
  AOI21  g03989(.A0(new_n4980_), .A1(\A[963] ), .B0(new_n4991_), .Y(new_n4992_));
  XOR2   g03990(.A(new_n4988_), .B(new_n4981_), .Y(new_n4993_));
  INV    g03991(.A(\A[957] ), .Y(new_n4994_));
  INV    g03992(.A(\A[956] ), .Y(new_n4995_));
  NAND2  g03993(.A(new_n4995_), .B(\A[955] ), .Y(new_n4996_));
  INV    g03994(.A(\A[955] ), .Y(new_n4997_));
  AOI21  g03995(.A0(\A[956] ), .A1(new_n4997_), .B0(new_n4994_), .Y(new_n4998_));
  XOR2   g03996(.A(\A[956] ), .B(\A[955] ), .Y(new_n4999_));
  AOI22  g03997(.A0(new_n4999_), .A1(new_n4994_), .B0(new_n4998_), .B1(new_n4996_), .Y(new_n5000_));
  INV    g03998(.A(\A[960] ), .Y(new_n5001_));
  INV    g03999(.A(\A[959] ), .Y(new_n5002_));
  NAND2  g04000(.A(new_n5002_), .B(\A[958] ), .Y(new_n5003_));
  INV    g04001(.A(\A[958] ), .Y(new_n5004_));
  AOI21  g04002(.A0(\A[959] ), .A1(new_n5004_), .B0(new_n5001_), .Y(new_n5005_));
  XOR2   g04003(.A(\A[959] ), .B(\A[958] ), .Y(new_n5006_));
  AOI22  g04004(.A0(new_n5006_), .A1(new_n5001_), .B0(new_n5005_), .B1(new_n5003_), .Y(new_n5007_));
  NAND2  g04005(.A(\A[959] ), .B(\A[958] ), .Y(new_n5008_));
  INV    g04006(.A(new_n5008_), .Y(new_n5009_));
  AOI21  g04007(.A0(new_n5006_), .A1(\A[960] ), .B0(new_n5009_), .Y(new_n5010_));
  NAND2  g04008(.A(\A[956] ), .B(\A[955] ), .Y(new_n5011_));
  INV    g04009(.A(new_n5011_), .Y(new_n5012_));
  AOI21  g04010(.A0(new_n4999_), .A1(\A[957] ), .B0(new_n5012_), .Y(new_n5013_));
  XOR2   g04011(.A(new_n5007_), .B(new_n5000_), .Y(new_n5014_));
  XOR2   g04012(.A(new_n5014_), .B(new_n4993_), .Y(new_n5015_));
  INV    g04013(.A(\A[951] ), .Y(new_n5016_));
  INV    g04014(.A(\A[950] ), .Y(new_n5017_));
  NAND2  g04015(.A(new_n5017_), .B(\A[949] ), .Y(new_n5018_));
  INV    g04016(.A(\A[949] ), .Y(new_n5019_));
  AOI21  g04017(.A0(\A[950] ), .A1(new_n5019_), .B0(new_n5016_), .Y(new_n5020_));
  XOR2   g04018(.A(\A[950] ), .B(\A[949] ), .Y(new_n5021_));
  AOI22  g04019(.A0(new_n5021_), .A1(new_n5016_), .B0(new_n5020_), .B1(new_n5018_), .Y(new_n5022_));
  INV    g04020(.A(\A[954] ), .Y(new_n5023_));
  INV    g04021(.A(\A[953] ), .Y(new_n5024_));
  NAND2  g04022(.A(new_n5024_), .B(\A[952] ), .Y(new_n5025_));
  INV    g04023(.A(\A[952] ), .Y(new_n5026_));
  AOI21  g04024(.A0(\A[953] ), .A1(new_n5026_), .B0(new_n5023_), .Y(new_n5027_));
  XOR2   g04025(.A(\A[953] ), .B(\A[952] ), .Y(new_n5028_));
  AOI22  g04026(.A0(new_n5028_), .A1(new_n5023_), .B0(new_n5027_), .B1(new_n5025_), .Y(new_n5029_));
  NOR2   g04027(.A(new_n5024_), .B(new_n5026_), .Y(new_n5030_));
  AOI21  g04028(.A0(new_n5028_), .A1(\A[954] ), .B0(new_n5030_), .Y(new_n5031_));
  NOR2   g04029(.A(new_n5017_), .B(new_n5019_), .Y(new_n5032_));
  AOI21  g04030(.A0(new_n5021_), .A1(\A[951] ), .B0(new_n5032_), .Y(new_n5033_));
  XOR2   g04031(.A(new_n5029_), .B(new_n5022_), .Y(new_n5034_));
  INV    g04032(.A(\A[945] ), .Y(new_n5035_));
  INV    g04033(.A(\A[944] ), .Y(new_n5036_));
  NAND2  g04034(.A(new_n5036_), .B(\A[943] ), .Y(new_n5037_));
  INV    g04035(.A(\A[943] ), .Y(new_n5038_));
  AOI21  g04036(.A0(\A[944] ), .A1(new_n5038_), .B0(new_n5035_), .Y(new_n5039_));
  XOR2   g04037(.A(\A[944] ), .B(\A[943] ), .Y(new_n5040_));
  AOI22  g04038(.A0(new_n5040_), .A1(new_n5035_), .B0(new_n5039_), .B1(new_n5037_), .Y(new_n5041_));
  INV    g04039(.A(\A[948] ), .Y(new_n5042_));
  INV    g04040(.A(\A[947] ), .Y(new_n5043_));
  NAND2  g04041(.A(new_n5043_), .B(\A[946] ), .Y(new_n5044_));
  INV    g04042(.A(\A[946] ), .Y(new_n5045_));
  AOI21  g04043(.A0(\A[947] ), .A1(new_n5045_), .B0(new_n5042_), .Y(new_n5046_));
  XOR2   g04044(.A(\A[947] ), .B(\A[946] ), .Y(new_n5047_));
  AOI22  g04045(.A0(new_n5047_), .A1(new_n5042_), .B0(new_n5046_), .B1(new_n5044_), .Y(new_n5048_));
  NAND2  g04046(.A(\A[947] ), .B(\A[946] ), .Y(new_n5049_));
  INV    g04047(.A(new_n5049_), .Y(new_n5050_));
  AOI21  g04048(.A0(new_n5047_), .A1(\A[948] ), .B0(new_n5050_), .Y(new_n5051_));
  NAND2  g04049(.A(\A[944] ), .B(\A[943] ), .Y(new_n5052_));
  INV    g04050(.A(new_n5052_), .Y(new_n5053_));
  AOI21  g04051(.A0(new_n5040_), .A1(\A[945] ), .B0(new_n5053_), .Y(new_n5054_));
  XOR2   g04052(.A(new_n5048_), .B(new_n5041_), .Y(new_n5055_));
  XOR2   g04053(.A(new_n5055_), .B(new_n5034_), .Y(new_n5056_));
  INV    g04054(.A(new_n5056_), .Y(new_n5057_));
  XOR2   g04055(.A(new_n5057_), .B(new_n5015_), .Y(new_n5058_));
  NOR2   g04056(.A(new_n5058_), .B(new_n4974_), .Y(new_n5059_));
  NOR3   g04057(.A(new_n4957_), .B(new_n4966_), .C(new_n4961_), .Y(new_n5060_));
  AOI21  g04058(.A0(new_n4949_), .A1(new_n4931_), .B0(new_n4971_), .Y(new_n5061_));
  OAI21  g04059(.A0(new_n5061_), .A1(new_n5060_), .B0(new_n4858_), .Y(new_n5062_));
  NAND2  g04060(.A(new_n5059_), .B(new_n5062_), .Y(new_n5063_));
  NOR2   g04061(.A(new_n4857_), .B(new_n4799_), .Y(new_n5064_));
  AOI21  g04062(.A0(new_n4843_), .A1(new_n4799_), .B0(new_n5064_), .Y(new_n5065_));
  NAND3  g04063(.A(new_n4971_), .B(new_n4949_), .C(new_n4931_), .Y(new_n5066_));
  OAI21  g04064(.A0(new_n4966_), .A1(new_n4961_), .B0(new_n4957_), .Y(new_n5067_));
  AOI21  g04065(.A0(new_n5067_), .A1(new_n5066_), .B0(new_n5065_), .Y(new_n5068_));
  NOR2   g04066(.A(new_n5068_), .B(new_n4973_), .Y(new_n5069_));
  OAI22  g04067(.A0(new_n5069_), .A1(new_n5059_), .B0(new_n5063_), .B1(new_n4973_), .Y(new_n5070_));
  XOR2   g04068(.A(new_n5048_), .B(new_n5041_), .Y(new_n5071_));
  XOR2   g04069(.A(new_n5054_), .B(new_n5051_), .Y(new_n5072_));
  NOR2   g04070(.A(new_n5048_), .B(new_n5041_), .Y(new_n5073_));
  NAND2  g04071(.A(new_n5073_), .B(new_n5072_), .Y(new_n5074_));
  INV    g04072(.A(new_n5047_), .Y(new_n5075_));
  OAI21  g04073(.A0(new_n5075_), .A1(new_n5042_), .B0(new_n5049_), .Y(new_n5076_));
  INV    g04074(.A(new_n5040_), .Y(new_n5077_));
  OAI21  g04075(.A0(new_n5077_), .A1(new_n5035_), .B0(new_n5052_), .Y(new_n5078_));
  NAND2  g04076(.A(new_n5078_), .B(new_n5076_), .Y(new_n5079_));
  NAND2  g04077(.A(new_n5079_), .B(new_n5074_), .Y(new_n5080_));
  XOR2   g04078(.A(new_n5054_), .B(new_n5076_), .Y(new_n5081_));
  XOR2   g04079(.A(new_n5073_), .B(new_n5081_), .Y(new_n5082_));
  AOI21  g04080(.A0(new_n5080_), .A1(new_n5071_), .B0(new_n5082_), .Y(new_n5083_));
  XOR2   g04081(.A(new_n5029_), .B(new_n5022_), .Y(new_n5084_));
  NOR2   g04082(.A(\A[950] ), .B(new_n5019_), .Y(new_n5085_));
  OAI21  g04083(.A0(new_n5017_), .A1(\A[949] ), .B0(\A[951] ), .Y(new_n5086_));
  NAND2  g04084(.A(new_n5021_), .B(new_n5016_), .Y(new_n5087_));
  OAI21  g04085(.A0(new_n5086_), .A1(new_n5085_), .B0(new_n5087_), .Y(new_n5088_));
  NOR2   g04086(.A(\A[953] ), .B(new_n5026_), .Y(new_n5089_));
  OAI21  g04087(.A0(new_n5024_), .A1(\A[952] ), .B0(\A[954] ), .Y(new_n5090_));
  NAND2  g04088(.A(new_n5028_), .B(new_n5023_), .Y(new_n5091_));
  OAI21  g04089(.A0(new_n5090_), .A1(new_n5089_), .B0(new_n5091_), .Y(new_n5092_));
  NAND2  g04090(.A(new_n5028_), .B(\A[954] ), .Y(new_n5093_));
  OAI21  g04091(.A0(new_n5024_), .A1(new_n5026_), .B0(new_n5093_), .Y(new_n5094_));
  NAND2  g04092(.A(new_n5021_), .B(\A[951] ), .Y(new_n5095_));
  OAI21  g04093(.A0(new_n5017_), .A1(new_n5019_), .B0(new_n5095_), .Y(new_n5096_));
  NAND4  g04094(.A(new_n5096_), .B(new_n5094_), .C(new_n5092_), .D(new_n5088_), .Y(new_n5097_));
  NAND3  g04095(.A(new_n5073_), .B(new_n5078_), .C(new_n5076_), .Y(new_n5098_));
  NAND4  g04096(.A(new_n5098_), .B(new_n5071_), .C(new_n5097_), .D(new_n5084_), .Y(new_n5099_));
  XOR2   g04097(.A(new_n5033_), .B(new_n5094_), .Y(new_n5100_));
  NAND2  g04098(.A(new_n5092_), .B(new_n5088_), .Y(new_n5101_));
  NAND2  g04099(.A(new_n5096_), .B(new_n5094_), .Y(new_n5102_));
  OAI21  g04100(.A0(new_n5101_), .A1(new_n5100_), .B0(new_n5102_), .Y(new_n5103_));
  NOR2   g04101(.A(new_n5029_), .B(new_n5022_), .Y(new_n5104_));
  XOR2   g04102(.A(new_n5104_), .B(new_n5100_), .Y(new_n5105_));
  AOI21  g04103(.A0(new_n5103_), .A1(new_n5084_), .B0(new_n5105_), .Y(new_n5106_));
  XOR2   g04104(.A(new_n5106_), .B(new_n5099_), .Y(new_n5107_));
  XOR2   g04105(.A(new_n5029_), .B(new_n5088_), .Y(new_n5108_));
  NOR4   g04106(.A(new_n5033_), .B(new_n5031_), .C(new_n5029_), .D(new_n5022_), .Y(new_n5109_));
  NAND2  g04107(.A(new_n5039_), .B(new_n5037_), .Y(new_n5110_));
  OAI21  g04108(.A0(new_n5077_), .A1(\A[945] ), .B0(new_n5110_), .Y(new_n5111_));
  XOR2   g04109(.A(new_n5048_), .B(new_n5111_), .Y(new_n5112_));
  NOR4   g04110(.A(new_n5054_), .B(new_n5051_), .C(new_n5048_), .D(new_n5041_), .Y(new_n5113_));
  NOR4   g04111(.A(new_n5113_), .B(new_n5112_), .C(new_n5109_), .D(new_n5108_), .Y(new_n5114_));
  XOR2   g04112(.A(new_n5033_), .B(new_n5031_), .Y(new_n5115_));
  NOR2   g04113(.A(new_n5033_), .B(new_n5031_), .Y(new_n5116_));
  AOI21  g04114(.A0(new_n5104_), .A1(new_n5115_), .B0(new_n5116_), .Y(new_n5117_));
  NOR4   g04115(.A(new_n5112_), .B(new_n5109_), .C(new_n5105_), .D(new_n5108_), .Y(new_n5118_));
  OAI211 g04116(.A0(new_n5117_), .A1(new_n5108_), .B0(new_n5118_), .B1(new_n5098_), .Y(new_n5119_));
  OAI21  g04117(.A0(new_n5106_), .A1(new_n5114_), .B0(new_n5119_), .Y(new_n5120_));
  NAND2  g04118(.A(new_n5120_), .B(new_n5083_), .Y(new_n5121_));
  OAI21  g04119(.A0(new_n5107_), .A1(new_n5083_), .B0(new_n5121_), .Y(new_n5122_));
  XOR2   g04120(.A(new_n5007_), .B(new_n5000_), .Y(new_n5123_));
  XOR2   g04121(.A(new_n5013_), .B(new_n5010_), .Y(new_n5124_));
  NOR2   g04122(.A(new_n5007_), .B(new_n5000_), .Y(new_n5125_));
  NAND2  g04123(.A(new_n5125_), .B(new_n5124_), .Y(new_n5126_));
  OAI21  g04124(.A0(new_n5013_), .A1(new_n5010_), .B0(new_n5126_), .Y(new_n5127_));
  INV    g04125(.A(new_n5006_), .Y(new_n5128_));
  OAI21  g04126(.A0(new_n5128_), .A1(new_n5001_), .B0(new_n5008_), .Y(new_n5129_));
  XOR2   g04127(.A(new_n5013_), .B(new_n5129_), .Y(new_n5130_));
  XOR2   g04128(.A(new_n5125_), .B(new_n5130_), .Y(new_n5131_));
  AOI21  g04129(.A0(new_n5127_), .A1(new_n5123_), .B0(new_n5131_), .Y(new_n5132_));
  XOR2   g04130(.A(new_n4988_), .B(new_n4981_), .Y(new_n5133_));
  NOR2   g04131(.A(\A[962] ), .B(new_n4978_), .Y(new_n5134_));
  OAI21  g04132(.A0(new_n4976_), .A1(\A[961] ), .B0(\A[963] ), .Y(new_n5135_));
  NAND2  g04133(.A(new_n4980_), .B(new_n4975_), .Y(new_n5136_));
  OAI21  g04134(.A0(new_n5135_), .A1(new_n5134_), .B0(new_n5136_), .Y(new_n5137_));
  NOR2   g04135(.A(\A[965] ), .B(new_n4985_), .Y(new_n5138_));
  OAI21  g04136(.A0(new_n4983_), .A1(\A[964] ), .B0(\A[966] ), .Y(new_n5139_));
  NAND2  g04137(.A(new_n4987_), .B(new_n4982_), .Y(new_n5140_));
  OAI21  g04138(.A0(new_n5139_), .A1(new_n5138_), .B0(new_n5140_), .Y(new_n5141_));
  NAND2  g04139(.A(new_n4987_), .B(\A[966] ), .Y(new_n5142_));
  OAI21  g04140(.A0(new_n4983_), .A1(new_n4985_), .B0(new_n5142_), .Y(new_n5143_));
  NAND2  g04141(.A(new_n4980_), .B(\A[963] ), .Y(new_n5144_));
  OAI21  g04142(.A0(new_n4976_), .A1(new_n4978_), .B0(new_n5144_), .Y(new_n5145_));
  NAND4  g04143(.A(new_n5145_), .B(new_n5143_), .C(new_n5141_), .D(new_n5137_), .Y(new_n5146_));
  INV    g04144(.A(new_n4999_), .Y(new_n5147_));
  OAI21  g04145(.A0(new_n5147_), .A1(new_n4994_), .B0(new_n5011_), .Y(new_n5148_));
  NAND3  g04146(.A(new_n5125_), .B(new_n5148_), .C(new_n5129_), .Y(new_n5149_));
  NAND4  g04147(.A(new_n5149_), .B(new_n5123_), .C(new_n5146_), .D(new_n5133_), .Y(new_n5150_));
  XOR2   g04148(.A(new_n4992_), .B(new_n5143_), .Y(new_n5151_));
  NAND2  g04149(.A(new_n5141_), .B(new_n5137_), .Y(new_n5152_));
  NAND2  g04150(.A(new_n5145_), .B(new_n5143_), .Y(new_n5153_));
  OAI21  g04151(.A0(new_n5152_), .A1(new_n5151_), .B0(new_n5153_), .Y(new_n5154_));
  NOR2   g04152(.A(new_n4988_), .B(new_n4981_), .Y(new_n5155_));
  XOR2   g04153(.A(new_n5155_), .B(new_n5151_), .Y(new_n5156_));
  AOI21  g04154(.A0(new_n5154_), .A1(new_n5133_), .B0(new_n5156_), .Y(new_n5157_));
  XOR2   g04155(.A(new_n5157_), .B(new_n5150_), .Y(new_n5158_));
  NOR2   g04156(.A(new_n5158_), .B(new_n5132_), .Y(new_n5159_));
  NAND2  g04157(.A(new_n4998_), .B(new_n4996_), .Y(new_n5160_));
  OAI21  g04158(.A0(new_n5147_), .A1(\A[957] ), .B0(new_n5160_), .Y(new_n5161_));
  XOR2   g04159(.A(new_n5007_), .B(new_n5161_), .Y(new_n5162_));
  NOR2   g04160(.A(new_n5013_), .B(new_n5010_), .Y(new_n5163_));
  AOI21  g04161(.A0(new_n5125_), .A1(new_n5124_), .B0(new_n5163_), .Y(new_n5164_));
  XOR2   g04162(.A(new_n5125_), .B(new_n5124_), .Y(new_n5165_));
  OAI21  g04163(.A0(new_n5164_), .A1(new_n5162_), .B0(new_n5165_), .Y(new_n5166_));
  XOR2   g04164(.A(new_n4988_), .B(new_n5137_), .Y(new_n5167_));
  XOR2   g04165(.A(new_n4992_), .B(new_n4990_), .Y(new_n5168_));
  NOR2   g04166(.A(new_n4992_), .B(new_n4990_), .Y(new_n5169_));
  AOI21  g04167(.A0(new_n5155_), .A1(new_n5168_), .B0(new_n5169_), .Y(new_n5170_));
  XOR2   g04168(.A(new_n5155_), .B(new_n5168_), .Y(new_n5171_));
  OAI21  g04169(.A0(new_n5170_), .A1(new_n5167_), .B0(new_n5171_), .Y(new_n5172_));
  NAND2  g04170(.A(new_n5172_), .B(new_n5150_), .Y(new_n5173_));
  NOR4   g04171(.A(new_n4992_), .B(new_n4990_), .C(new_n4988_), .D(new_n4981_), .Y(new_n5174_));
  NOR4   g04172(.A(new_n5162_), .B(new_n5174_), .C(new_n5156_), .D(new_n5167_), .Y(new_n5175_));
  OAI211 g04173(.A0(new_n5170_), .A1(new_n5167_), .B0(new_n5175_), .B1(new_n5149_), .Y(new_n5176_));
  AOI21  g04174(.A0(new_n5176_), .A1(new_n5173_), .B0(new_n5166_), .Y(new_n5177_));
  NAND2  g04175(.A(new_n5056_), .B(new_n5015_), .Y(new_n5178_));
  NOR3   g04176(.A(new_n5178_), .B(new_n5177_), .C(new_n5159_), .Y(new_n5179_));
  NOR4   g04177(.A(new_n5013_), .B(new_n5010_), .C(new_n5007_), .D(new_n5000_), .Y(new_n5180_));
  NOR4   g04178(.A(new_n5180_), .B(new_n5162_), .C(new_n5174_), .D(new_n5167_), .Y(new_n5181_));
  XOR2   g04179(.A(new_n5157_), .B(new_n5181_), .Y(new_n5182_));
  NAND2  g04180(.A(new_n5182_), .B(new_n5166_), .Y(new_n5183_));
  NAND4  g04181(.A(new_n5123_), .B(new_n5146_), .C(new_n5171_), .D(new_n5133_), .Y(new_n5184_));
  OAI21  g04182(.A0(new_n5170_), .A1(new_n5167_), .B0(new_n5149_), .Y(new_n5185_));
  OAI22  g04183(.A0(new_n5185_), .A1(new_n5184_), .B0(new_n5157_), .B1(new_n5181_), .Y(new_n5186_));
  NAND2  g04184(.A(new_n5186_), .B(new_n5132_), .Y(new_n5187_));
  INV    g04185(.A(new_n5178_), .Y(new_n5188_));
  AOI21  g04186(.A0(new_n5187_), .A1(new_n5183_), .B0(new_n5188_), .Y(new_n5189_));
  NOR2   g04187(.A(new_n5189_), .B(new_n5179_), .Y(new_n5190_));
  NOR2   g04188(.A(new_n5122_), .B(new_n5190_), .Y(new_n5191_));
  NOR2   g04189(.A(new_n5177_), .B(new_n5159_), .Y(new_n5192_));
  NAND3  g04190(.A(new_n5178_), .B(new_n5187_), .C(new_n5183_), .Y(new_n5193_));
  OAI21  g04191(.A0(new_n5192_), .A1(new_n5178_), .B0(new_n5193_), .Y(new_n5194_));
  AOI21  g04192(.A0(new_n5194_), .A1(new_n5122_), .B0(new_n5191_), .Y(new_n5195_));
  NAND2  g04193(.A(new_n5195_), .B(new_n5070_), .Y(new_n5196_));
  NAND2  g04194(.A(new_n5194_), .B(new_n5122_), .Y(new_n5197_));
  OAI21  g04195(.A0(new_n5122_), .A1(new_n5190_), .B0(new_n5197_), .Y(new_n5198_));
  NOR3   g04196(.A(new_n5059_), .B(new_n5068_), .C(new_n4973_), .Y(new_n5199_));
  INV    g04197(.A(new_n5059_), .Y(new_n5200_));
  NOR2   g04198(.A(new_n5069_), .B(new_n5200_), .Y(new_n5201_));
  OAI21  g04199(.A0(new_n5201_), .A1(new_n5199_), .B0(new_n5198_), .Y(new_n5202_));
  NAND2  g04200(.A(new_n5202_), .B(new_n5196_), .Y(new_n5203_));
  INV    g04201(.A(\A[8] ), .Y(new_n5204_));
  NOR2   g04202(.A(new_n5204_), .B(\A[7] ), .Y(new_n5205_));
  INV    g04203(.A(\A[7] ), .Y(new_n5206_));
  OAI21  g04204(.A0(\A[8] ), .A1(new_n5206_), .B0(\A[9] ), .Y(new_n5207_));
  XOR2   g04205(.A(\A[8] ), .B(new_n5206_), .Y(new_n5208_));
  OAI22  g04206(.A0(new_n5208_), .A1(\A[9] ), .B0(new_n5207_), .B1(new_n5205_), .Y(new_n5209_));
  INV    g04207(.A(\A[11] ), .Y(new_n5210_));
  NOR2   g04208(.A(new_n5210_), .B(\A[10] ), .Y(new_n5211_));
  INV    g04209(.A(\A[10] ), .Y(new_n5212_));
  OAI21  g04210(.A0(\A[11] ), .A1(new_n5212_), .B0(\A[12] ), .Y(new_n5213_));
  XOR2   g04211(.A(\A[11] ), .B(new_n5212_), .Y(new_n5214_));
  OAI22  g04212(.A0(new_n5214_), .A1(\A[12] ), .B0(new_n5213_), .B1(new_n5211_), .Y(new_n5215_));
  NAND2  g04213(.A(new_n5215_), .B(new_n5209_), .Y(new_n5216_));
  INV    g04214(.A(\A[12] ), .Y(new_n5217_));
  NAND2  g04215(.A(\A[11] ), .B(\A[10] ), .Y(new_n5218_));
  OAI21  g04216(.A0(new_n5214_), .A1(new_n5217_), .B0(new_n5218_), .Y(new_n5219_));
  XOR2   g04217(.A(\A[8] ), .B(\A[7] ), .Y(new_n5220_));
  NOR2   g04218(.A(new_n5204_), .B(new_n5206_), .Y(new_n5221_));
  AOI21  g04219(.A0(new_n5220_), .A1(\A[9] ), .B0(new_n5221_), .Y(new_n5222_));
  XOR2   g04220(.A(new_n5222_), .B(new_n5219_), .Y(new_n5223_));
  XOR2   g04221(.A(new_n5223_), .B(new_n5216_), .Y(new_n5224_));
  NAND2  g04222(.A(\A[11] ), .B(new_n5212_), .Y(new_n5225_));
  AOI21  g04223(.A0(new_n5210_), .A1(\A[10] ), .B0(new_n5217_), .Y(new_n5226_));
  XOR2   g04224(.A(\A[11] ), .B(\A[10] ), .Y(new_n5227_));
  AOI22  g04225(.A0(new_n5227_), .A1(new_n5217_), .B0(new_n5226_), .B1(new_n5225_), .Y(new_n5228_));
  XOR2   g04226(.A(new_n5228_), .B(new_n5209_), .Y(new_n5229_));
  INV    g04227(.A(\A[9] ), .Y(new_n5230_));
  NAND2  g04228(.A(\A[8] ), .B(new_n5206_), .Y(new_n5231_));
  AOI21  g04229(.A0(new_n5204_), .A1(\A[7] ), .B0(new_n5230_), .Y(new_n5232_));
  AOI22  g04230(.A0(new_n5220_), .A1(new_n5230_), .B0(new_n5232_), .B1(new_n5231_), .Y(new_n5233_));
  NOR2   g04231(.A(new_n5228_), .B(new_n5233_), .Y(new_n5234_));
  NOR2   g04232(.A(new_n5210_), .B(new_n5212_), .Y(new_n5235_));
  AOI21  g04233(.A0(new_n5227_), .A1(\A[12] ), .B0(new_n5235_), .Y(new_n5236_));
  XOR2   g04234(.A(new_n5222_), .B(new_n5236_), .Y(new_n5237_));
  NOR2   g04235(.A(new_n5222_), .B(new_n5236_), .Y(new_n5238_));
  AOI21  g04236(.A0(new_n5237_), .A1(new_n5234_), .B0(new_n5238_), .Y(new_n5239_));
  OAI21  g04237(.A0(new_n5239_), .A1(new_n5229_), .B0(new_n5224_), .Y(new_n5240_));
  XOR2   g04238(.A(new_n5228_), .B(new_n5233_), .Y(new_n5241_));
  NAND2  g04239(.A(\A[17] ), .B(\A[16] ), .Y(new_n5242_));
  XOR2   g04240(.A(\A[17] ), .B(\A[16] ), .Y(new_n5243_));
  NAND2  g04241(.A(new_n5243_), .B(\A[18] ), .Y(new_n5244_));
  NAND2  g04242(.A(new_n5244_), .B(new_n5242_), .Y(new_n5245_));
  NAND2  g04243(.A(\A[14] ), .B(\A[13] ), .Y(new_n5246_));
  XOR2   g04244(.A(\A[14] ), .B(\A[13] ), .Y(new_n5247_));
  NAND2  g04245(.A(new_n5247_), .B(\A[15] ), .Y(new_n5248_));
  NAND2  g04246(.A(new_n5248_), .B(new_n5246_), .Y(new_n5249_));
  INV    g04247(.A(\A[14] ), .Y(new_n5250_));
  NOR2   g04248(.A(new_n5250_), .B(\A[13] ), .Y(new_n5251_));
  INV    g04249(.A(\A[13] ), .Y(new_n5252_));
  OAI21  g04250(.A0(\A[14] ), .A1(new_n5252_), .B0(\A[15] ), .Y(new_n5253_));
  INV    g04251(.A(\A[15] ), .Y(new_n5254_));
  NAND2  g04252(.A(new_n5247_), .B(new_n5254_), .Y(new_n5255_));
  OAI21  g04253(.A0(new_n5253_), .A1(new_n5251_), .B0(new_n5255_), .Y(new_n5256_));
  INV    g04254(.A(\A[17] ), .Y(new_n5257_));
  NOR2   g04255(.A(new_n5257_), .B(\A[16] ), .Y(new_n5258_));
  INV    g04256(.A(\A[16] ), .Y(new_n5259_));
  OAI21  g04257(.A0(\A[17] ), .A1(new_n5259_), .B0(\A[18] ), .Y(new_n5260_));
  INV    g04258(.A(\A[18] ), .Y(new_n5261_));
  NAND2  g04259(.A(new_n5243_), .B(new_n5261_), .Y(new_n5262_));
  OAI21  g04260(.A0(new_n5260_), .A1(new_n5258_), .B0(new_n5262_), .Y(new_n5263_));
  NAND4  g04261(.A(new_n5263_), .B(new_n5256_), .C(new_n5249_), .D(new_n5245_), .Y(new_n5264_));
  NAND2  g04262(.A(\A[8] ), .B(\A[7] ), .Y(new_n5265_));
  OAI21  g04263(.A0(new_n5208_), .A1(new_n5230_), .B0(new_n5265_), .Y(new_n5266_));
  NAND4  g04264(.A(new_n5266_), .B(new_n5219_), .C(new_n5215_), .D(new_n5209_), .Y(new_n5267_));
  NAND2  g04265(.A(\A[14] ), .B(new_n5252_), .Y(new_n5268_));
  AOI21  g04266(.A0(new_n5250_), .A1(\A[13] ), .B0(new_n5254_), .Y(new_n5269_));
  AOI22  g04267(.A0(new_n5269_), .A1(new_n5268_), .B0(new_n5247_), .B1(new_n5254_), .Y(new_n5270_));
  NAND2  g04268(.A(\A[17] ), .B(new_n5259_), .Y(new_n5271_));
  AOI21  g04269(.A0(new_n5257_), .A1(\A[16] ), .B0(new_n5261_), .Y(new_n5272_));
  AOI22  g04270(.A0(new_n5272_), .A1(new_n5271_), .B0(new_n5243_), .B1(new_n5261_), .Y(new_n5273_));
  XOR2   g04271(.A(new_n5273_), .B(new_n5270_), .Y(new_n5274_));
  NAND4  g04272(.A(new_n5274_), .B(new_n5267_), .C(new_n5264_), .D(new_n5241_), .Y(new_n5275_));
  XOR2   g04273(.A(new_n5249_), .B(new_n5245_), .Y(new_n5276_));
  NOR2   g04274(.A(new_n5273_), .B(new_n5270_), .Y(new_n5277_));
  AOI22  g04275(.A0(new_n5248_), .A1(new_n5246_), .B0(new_n5244_), .B1(new_n5242_), .Y(new_n5278_));
  AOI21  g04276(.A0(new_n5277_), .A1(new_n5276_), .B0(new_n5278_), .Y(new_n5279_));
  XOR2   g04277(.A(new_n5277_), .B(new_n5276_), .Y(new_n5280_));
  XOR2   g04278(.A(new_n5273_), .B(new_n5256_), .Y(new_n5281_));
  OAI21  g04279(.A0(new_n5281_), .A1(new_n5279_), .B0(new_n5280_), .Y(new_n5282_));
  XOR2   g04280(.A(new_n5282_), .B(new_n5275_), .Y(new_n5283_));
  NAND2  g04281(.A(new_n5263_), .B(new_n5256_), .Y(new_n5284_));
  XOR2   g04282(.A(new_n5284_), .B(new_n5276_), .Y(new_n5285_));
  NOR2   g04283(.A(new_n5250_), .B(new_n5252_), .Y(new_n5286_));
  AOI221 g04284(.A0(new_n5247_), .A1(\A[15] ), .C0(new_n5286_), .B0(new_n5244_), .B1(new_n5242_), .Y(new_n5287_));
  NOR2   g04285(.A(new_n5257_), .B(new_n5259_), .Y(new_n5288_));
  AOI221 g04286(.A0(new_n5248_), .A1(new_n5246_), .C0(new_n5288_), .B0(new_n5243_), .B1(\A[18] ), .Y(new_n5289_));
  OAI211 g04287(.A0(new_n5289_), .A1(new_n5287_), .B0(new_n5263_), .B1(new_n5256_), .Y(new_n5290_));
  NAND2  g04288(.A(new_n5249_), .B(new_n5245_), .Y(new_n5291_));
  AOI21  g04289(.A0(new_n5291_), .A1(new_n5290_), .B0(new_n5281_), .Y(new_n5292_));
  OAI21  g04290(.A0(new_n5292_), .A1(new_n5285_), .B0(new_n5275_), .Y(new_n5293_));
  NOR2   g04291(.A(new_n5281_), .B(new_n5229_), .Y(new_n5294_));
  OAI211 g04292(.A0(new_n5263_), .A1(new_n5256_), .B0(new_n5249_), .B1(new_n5245_), .Y(new_n5295_));
  NAND4  g04293(.A(new_n5295_), .B(new_n5294_), .C(new_n5267_), .D(new_n5280_), .Y(new_n5296_));
  AOI21  g04294(.A0(new_n5296_), .A1(new_n5293_), .B0(new_n5240_), .Y(new_n5297_));
  AOI21  g04295(.A0(new_n5283_), .A1(new_n5240_), .B0(new_n5297_), .Y(new_n5298_));
  INV    g04296(.A(\A[21] ), .Y(new_n5299_));
  INV    g04297(.A(\A[19] ), .Y(new_n5300_));
  NAND2  g04298(.A(\A[20] ), .B(new_n5300_), .Y(new_n5301_));
  INV    g04299(.A(\A[20] ), .Y(new_n5302_));
  AOI21  g04300(.A0(new_n5302_), .A1(\A[19] ), .B0(new_n5299_), .Y(new_n5303_));
  XOR2   g04301(.A(\A[20] ), .B(\A[19] ), .Y(new_n5304_));
  AOI22  g04302(.A0(new_n5304_), .A1(new_n5299_), .B0(new_n5303_), .B1(new_n5301_), .Y(new_n5305_));
  INV    g04303(.A(\A[24] ), .Y(new_n5306_));
  INV    g04304(.A(\A[22] ), .Y(new_n5307_));
  NAND2  g04305(.A(\A[23] ), .B(new_n5307_), .Y(new_n5308_));
  INV    g04306(.A(\A[23] ), .Y(new_n5309_));
  AOI21  g04307(.A0(new_n5309_), .A1(\A[22] ), .B0(new_n5306_), .Y(new_n5310_));
  XOR2   g04308(.A(\A[23] ), .B(\A[22] ), .Y(new_n5311_));
  AOI22  g04309(.A0(new_n5311_), .A1(new_n5306_), .B0(new_n5310_), .B1(new_n5308_), .Y(new_n5312_));
  NOR2   g04310(.A(new_n5312_), .B(new_n5305_), .Y(new_n5313_));
  XOR2   g04311(.A(\A[23] ), .B(new_n5307_), .Y(new_n5314_));
  NAND2  g04312(.A(\A[23] ), .B(\A[22] ), .Y(new_n5315_));
  OAI21  g04313(.A0(new_n5314_), .A1(new_n5306_), .B0(new_n5315_), .Y(new_n5316_));
  NOR2   g04314(.A(new_n5302_), .B(new_n5300_), .Y(new_n5317_));
  AOI21  g04315(.A0(new_n5304_), .A1(\A[21] ), .B0(new_n5317_), .Y(new_n5318_));
  XOR2   g04316(.A(new_n5318_), .B(new_n5316_), .Y(new_n5319_));
  XOR2   g04317(.A(new_n5319_), .B(new_n5313_), .Y(new_n5320_));
  XOR2   g04318(.A(new_n5312_), .B(new_n5305_), .Y(new_n5321_));
  NOR2   g04319(.A(new_n5302_), .B(\A[19] ), .Y(new_n5322_));
  OAI21  g04320(.A0(\A[20] ), .A1(new_n5300_), .B0(\A[21] ), .Y(new_n5323_));
  XOR2   g04321(.A(\A[20] ), .B(new_n5300_), .Y(new_n5324_));
  OAI22  g04322(.A0(new_n5324_), .A1(\A[21] ), .B0(new_n5323_), .B1(new_n5322_), .Y(new_n5325_));
  NOR2   g04323(.A(new_n5309_), .B(\A[22] ), .Y(new_n5326_));
  OAI21  g04324(.A0(\A[23] ), .A1(new_n5307_), .B0(\A[24] ), .Y(new_n5327_));
  OAI22  g04325(.A0(new_n5314_), .A1(\A[24] ), .B0(new_n5327_), .B1(new_n5326_), .Y(new_n5328_));
  NAND2  g04326(.A(new_n5328_), .B(new_n5325_), .Y(new_n5329_));
  NAND2  g04327(.A(\A[20] ), .B(\A[19] ), .Y(new_n5330_));
  OAI21  g04328(.A0(new_n5324_), .A1(new_n5299_), .B0(new_n5330_), .Y(new_n5331_));
  NAND2  g04329(.A(new_n5331_), .B(new_n5316_), .Y(new_n5332_));
  OAI21  g04330(.A0(new_n5319_), .A1(new_n5329_), .B0(new_n5332_), .Y(new_n5333_));
  AOI21  g04331(.A0(new_n5333_), .A1(new_n5321_), .B0(new_n5320_), .Y(new_n5334_));
  NAND2  g04332(.A(\A[29] ), .B(\A[28] ), .Y(new_n5335_));
  XOR2   g04333(.A(\A[29] ), .B(\A[28] ), .Y(new_n5336_));
  NAND2  g04334(.A(new_n5336_), .B(\A[30] ), .Y(new_n5337_));
  NAND2  g04335(.A(new_n5337_), .B(new_n5335_), .Y(new_n5338_));
  NAND2  g04336(.A(\A[26] ), .B(\A[25] ), .Y(new_n5339_));
  XOR2   g04337(.A(\A[26] ), .B(\A[25] ), .Y(new_n5340_));
  NAND2  g04338(.A(new_n5340_), .B(\A[27] ), .Y(new_n5341_));
  NAND2  g04339(.A(new_n5341_), .B(new_n5339_), .Y(new_n5342_));
  XOR2   g04340(.A(new_n5342_), .B(new_n5338_), .Y(new_n5343_));
  INV    g04341(.A(\A[27] ), .Y(new_n5344_));
  INV    g04342(.A(\A[25] ), .Y(new_n5345_));
  NAND2  g04343(.A(\A[26] ), .B(new_n5345_), .Y(new_n5346_));
  INV    g04344(.A(\A[26] ), .Y(new_n5347_));
  AOI21  g04345(.A0(new_n5347_), .A1(\A[25] ), .B0(new_n5344_), .Y(new_n5348_));
  AOI22  g04346(.A0(new_n5348_), .A1(new_n5346_), .B0(new_n5340_), .B1(new_n5344_), .Y(new_n5349_));
  INV    g04347(.A(\A[30] ), .Y(new_n5350_));
  INV    g04348(.A(\A[28] ), .Y(new_n5351_));
  NAND2  g04349(.A(\A[29] ), .B(new_n5351_), .Y(new_n5352_));
  INV    g04350(.A(\A[29] ), .Y(new_n5353_));
  AOI21  g04351(.A0(new_n5353_), .A1(\A[28] ), .B0(new_n5350_), .Y(new_n5354_));
  AOI22  g04352(.A0(new_n5354_), .A1(new_n5352_), .B0(new_n5336_), .B1(new_n5350_), .Y(new_n5355_));
  NOR2   g04353(.A(new_n5355_), .B(new_n5349_), .Y(new_n5356_));
  AOI22  g04354(.A0(new_n5341_), .A1(new_n5339_), .B0(new_n5337_), .B1(new_n5335_), .Y(new_n5357_));
  AOI21  g04355(.A0(new_n5356_), .A1(new_n5343_), .B0(new_n5357_), .Y(new_n5358_));
  XOR2   g04356(.A(new_n5356_), .B(new_n5343_), .Y(new_n5359_));
  NOR2   g04357(.A(new_n5347_), .B(\A[25] ), .Y(new_n5360_));
  OAI21  g04358(.A0(\A[26] ), .A1(new_n5345_), .B0(\A[27] ), .Y(new_n5361_));
  NAND2  g04359(.A(new_n5340_), .B(new_n5344_), .Y(new_n5362_));
  OAI21  g04360(.A0(new_n5361_), .A1(new_n5360_), .B0(new_n5362_), .Y(new_n5363_));
  XOR2   g04361(.A(new_n5355_), .B(new_n5363_), .Y(new_n5364_));
  NOR2   g04362(.A(new_n5353_), .B(\A[28] ), .Y(new_n5365_));
  OAI21  g04363(.A0(\A[29] ), .A1(new_n5351_), .B0(\A[30] ), .Y(new_n5366_));
  NAND2  g04364(.A(new_n5336_), .B(new_n5350_), .Y(new_n5367_));
  OAI21  g04365(.A0(new_n5366_), .A1(new_n5365_), .B0(new_n5367_), .Y(new_n5368_));
  NAND4  g04366(.A(new_n5368_), .B(new_n5363_), .C(new_n5342_), .D(new_n5338_), .Y(new_n5369_));
  NAND4  g04367(.A(new_n5331_), .B(new_n5316_), .C(new_n5328_), .D(new_n5325_), .Y(new_n5370_));
  XOR2   g04368(.A(new_n5355_), .B(new_n5349_), .Y(new_n5371_));
  NAND4  g04369(.A(new_n5371_), .B(new_n5370_), .C(new_n5369_), .D(new_n5321_), .Y(new_n5372_));
  OAI211 g04370(.A0(new_n5364_), .A1(new_n5358_), .B0(new_n5372_), .B1(new_n5359_), .Y(new_n5373_));
  NOR2   g04371(.A(new_n5347_), .B(new_n5345_), .Y(new_n5374_));
  AOI21  g04372(.A0(new_n5340_), .A1(\A[27] ), .B0(new_n5374_), .Y(new_n5375_));
  XOR2   g04373(.A(new_n5375_), .B(new_n5338_), .Y(new_n5376_));
  XOR2   g04374(.A(new_n5356_), .B(new_n5376_), .Y(new_n5377_));
  XOR2   g04375(.A(new_n5312_), .B(new_n5325_), .Y(new_n5378_));
  NOR2   g04376(.A(new_n5353_), .B(new_n5351_), .Y(new_n5379_));
  AOI21  g04377(.A0(new_n5336_), .A1(\A[30] ), .B0(new_n5379_), .Y(new_n5380_));
  NOR4   g04378(.A(new_n5355_), .B(new_n5349_), .C(new_n5375_), .D(new_n5380_), .Y(new_n5381_));
  NOR2   g04379(.A(new_n5309_), .B(new_n5307_), .Y(new_n5382_));
  AOI21  g04380(.A0(new_n5311_), .A1(\A[24] ), .B0(new_n5382_), .Y(new_n5383_));
  NOR4   g04381(.A(new_n5318_), .B(new_n5383_), .C(new_n5312_), .D(new_n5305_), .Y(new_n5384_));
  NOR4   g04382(.A(new_n5364_), .B(new_n5384_), .C(new_n5381_), .D(new_n5378_), .Y(new_n5385_));
  AOI221 g04383(.A0(new_n5340_), .A1(\A[27] ), .C0(new_n5374_), .B0(new_n5337_), .B1(new_n5335_), .Y(new_n5386_));
  AOI221 g04384(.A0(new_n5341_), .A1(new_n5339_), .C0(new_n5379_), .B0(new_n5336_), .B1(\A[30] ), .Y(new_n5387_));
  OAI211 g04385(.A0(new_n5387_), .A1(new_n5386_), .B0(new_n5368_), .B1(new_n5363_), .Y(new_n5388_));
  NAND2  g04386(.A(new_n5342_), .B(new_n5338_), .Y(new_n5389_));
  AOI21  g04387(.A0(new_n5389_), .A1(new_n5388_), .B0(new_n5364_), .Y(new_n5390_));
  OAI21  g04388(.A0(new_n5390_), .A1(new_n5377_), .B0(new_n5385_), .Y(new_n5391_));
  AOI21  g04389(.A0(new_n5391_), .A1(new_n5373_), .B0(new_n5334_), .Y(new_n5392_));
  XOR2   g04390(.A(new_n5319_), .B(new_n5329_), .Y(new_n5393_));
  XOR2   g04391(.A(new_n5318_), .B(new_n5383_), .Y(new_n5394_));
  NOR2   g04392(.A(new_n5318_), .B(new_n5383_), .Y(new_n5395_));
  AOI21  g04393(.A0(new_n5394_), .A1(new_n5313_), .B0(new_n5395_), .Y(new_n5396_));
  OAI21  g04394(.A0(new_n5396_), .A1(new_n5378_), .B0(new_n5393_), .Y(new_n5397_));
  OAI21  g04395(.A0(new_n5390_), .A1(new_n5377_), .B0(new_n5372_), .Y(new_n5398_));
  NOR2   g04396(.A(new_n5364_), .B(new_n5378_), .Y(new_n5399_));
  OAI211 g04397(.A0(new_n5368_), .A1(new_n5363_), .B0(new_n5342_), .B1(new_n5338_), .Y(new_n5400_));
  NAND4  g04398(.A(new_n5400_), .B(new_n5399_), .C(new_n5370_), .D(new_n5359_), .Y(new_n5401_));
  AOI21  g04399(.A0(new_n5401_), .A1(new_n5398_), .B0(new_n5397_), .Y(new_n5402_));
  NOR2   g04400(.A(new_n5364_), .B(new_n5381_), .Y(new_n5403_));
  XOR2   g04401(.A(new_n5312_), .B(new_n5305_), .Y(new_n5404_));
  XOR2   g04402(.A(new_n5404_), .B(new_n5403_), .Y(new_n5405_));
  NAND2  g04403(.A(new_n5274_), .B(new_n5264_), .Y(new_n5406_));
  XOR2   g04404(.A(new_n5228_), .B(new_n5209_), .Y(new_n5407_));
  XOR2   g04405(.A(new_n5407_), .B(new_n5406_), .Y(new_n5408_));
  NAND2  g04406(.A(new_n5408_), .B(new_n5405_), .Y(new_n5409_));
  NOR3   g04407(.A(new_n5409_), .B(new_n5402_), .C(new_n5392_), .Y(new_n5410_));
  OAI21  g04408(.A0(new_n5364_), .A1(new_n5358_), .B0(new_n5359_), .Y(new_n5411_));
  XOR2   g04409(.A(new_n5411_), .B(new_n5372_), .Y(new_n5412_));
  NAND2  g04410(.A(new_n5412_), .B(new_n5397_), .Y(new_n5413_));
  NAND2  g04411(.A(new_n5401_), .B(new_n5398_), .Y(new_n5414_));
  NAND2  g04412(.A(new_n5414_), .B(new_n5334_), .Y(new_n5415_));
  NAND2  g04413(.A(new_n5371_), .B(new_n5369_), .Y(new_n5416_));
  XOR2   g04414(.A(new_n5404_), .B(new_n5416_), .Y(new_n5417_));
  XOR2   g04415(.A(new_n5228_), .B(new_n5233_), .Y(new_n5418_));
  XOR2   g04416(.A(new_n5418_), .B(new_n5406_), .Y(new_n5419_));
  NOR2   g04417(.A(new_n5419_), .B(new_n5417_), .Y(new_n5420_));
  AOI21  g04418(.A0(new_n5415_), .A1(new_n5413_), .B0(new_n5420_), .Y(new_n5421_));
  OAI21  g04419(.A0(new_n5421_), .A1(new_n5410_), .B0(new_n5298_), .Y(new_n5422_));
  XOR2   g04420(.A(new_n5223_), .B(new_n5234_), .Y(new_n5423_));
  NAND2  g04421(.A(new_n5266_), .B(new_n5219_), .Y(new_n5424_));
  OAI21  g04422(.A0(new_n5223_), .A1(new_n5216_), .B0(new_n5424_), .Y(new_n5425_));
  AOI21  g04423(.A0(new_n5425_), .A1(new_n5241_), .B0(new_n5423_), .Y(new_n5426_));
  NOR2   g04424(.A(new_n5292_), .B(new_n5285_), .Y(new_n5427_));
  XOR2   g04425(.A(new_n5427_), .B(new_n5275_), .Y(new_n5428_));
  NAND2  g04426(.A(new_n5296_), .B(new_n5293_), .Y(new_n5429_));
  NAND2  g04427(.A(new_n5429_), .B(new_n5426_), .Y(new_n5430_));
  OAI21  g04428(.A0(new_n5428_), .A1(new_n5426_), .B0(new_n5430_), .Y(new_n5431_));
  NAND2  g04429(.A(new_n5371_), .B(new_n5321_), .Y(new_n5432_));
  AOI211 g04430(.A0(new_n5355_), .A1(new_n5349_), .B(new_n5375_), .C(new_n5380_), .Y(new_n5433_));
  NOR4   g04431(.A(new_n5433_), .B(new_n5432_), .C(new_n5384_), .D(new_n5377_), .Y(new_n5434_));
  AOI21  g04432(.A0(new_n5411_), .A1(new_n5372_), .B0(new_n5434_), .Y(new_n5435_));
  OAI21  g04433(.A0(new_n5435_), .A1(new_n5397_), .B0(new_n5409_), .Y(new_n5436_));
  OAI21  g04434(.A0(new_n5402_), .A1(new_n5392_), .B0(new_n5420_), .Y(new_n5437_));
  OAI21  g04435(.A0(new_n5436_), .A1(new_n5392_), .B0(new_n5437_), .Y(new_n5438_));
  NAND2  g04436(.A(new_n5438_), .B(new_n5431_), .Y(new_n5439_));
  NAND2  g04437(.A(new_n5419_), .B(new_n5405_), .Y(new_n5440_));
  NAND2  g04438(.A(new_n5408_), .B(new_n5417_), .Y(new_n5441_));
  INV    g04439(.A(\A[993] ), .Y(new_n5442_));
  INV    g04440(.A(\A[992] ), .Y(new_n5443_));
  NAND2  g04441(.A(new_n5443_), .B(\A[991] ), .Y(new_n5444_));
  INV    g04442(.A(\A[991] ), .Y(new_n5445_));
  AOI21  g04443(.A0(\A[992] ), .A1(new_n5445_), .B0(new_n5442_), .Y(new_n5446_));
  XOR2   g04444(.A(\A[992] ), .B(\A[991] ), .Y(new_n5447_));
  AOI22  g04445(.A0(new_n5447_), .A1(new_n5442_), .B0(new_n5446_), .B1(new_n5444_), .Y(new_n5448_));
  INV    g04446(.A(\A[996] ), .Y(new_n5449_));
  INV    g04447(.A(\A[995] ), .Y(new_n5450_));
  NAND2  g04448(.A(new_n5450_), .B(\A[994] ), .Y(new_n5451_));
  INV    g04449(.A(\A[994] ), .Y(new_n5452_));
  AOI21  g04450(.A0(\A[995] ), .A1(new_n5452_), .B0(new_n5449_), .Y(new_n5453_));
  XOR2   g04451(.A(\A[995] ), .B(\A[994] ), .Y(new_n5454_));
  AOI22  g04452(.A0(new_n5454_), .A1(new_n5449_), .B0(new_n5453_), .B1(new_n5451_), .Y(new_n5455_));
  NOR2   g04453(.A(new_n5450_), .B(new_n5452_), .Y(new_n5456_));
  AOI21  g04454(.A0(new_n5454_), .A1(\A[996] ), .B0(new_n5456_), .Y(new_n5457_));
  NOR2   g04455(.A(new_n5443_), .B(new_n5445_), .Y(new_n5458_));
  AOI21  g04456(.A0(new_n5447_), .A1(\A[993] ), .B0(new_n5458_), .Y(new_n5459_));
  XOR2   g04457(.A(new_n5455_), .B(new_n5448_), .Y(new_n5460_));
  INV    g04458(.A(\A[999] ), .Y(new_n5461_));
  INV    g04459(.A(\A[998] ), .Y(new_n5462_));
  NAND2  g04460(.A(new_n5462_), .B(\A[997] ), .Y(new_n5463_));
  INV    g04461(.A(\A[997] ), .Y(new_n5464_));
  AOI21  g04462(.A0(\A[998] ), .A1(new_n5464_), .B0(new_n5461_), .Y(new_n5465_));
  XOR2   g04463(.A(\A[998] ), .B(\A[997] ), .Y(new_n5466_));
  AOI22  g04464(.A0(new_n5466_), .A1(new_n5461_), .B0(new_n5465_), .B1(new_n5463_), .Y(new_n5467_));
  INV    g04465(.A(\A[5] ), .Y(new_n5468_));
  INV    g04466(.A(\A[3] ), .Y(new_n5469_));
  NAND2  g04467(.A(\A[4] ), .B(new_n5469_), .Y(new_n5470_));
  INV    g04468(.A(\A[4] ), .Y(new_n5471_));
  AOI21  g04469(.A0(new_n5471_), .A1(\A[3] ), .B0(new_n5468_), .Y(new_n5472_));
  XOR2   g04470(.A(\A[4] ), .B(\A[3] ), .Y(new_n5473_));
  AOI22  g04471(.A0(new_n5473_), .A1(new_n5468_), .B0(new_n5472_), .B1(new_n5470_), .Y(new_n5474_));
  INV    g04472(.A(\A[6] ), .Y(new_n5475_));
  INV    g04473(.A(\A[0] ), .Y(new_n5476_));
  NOR2   g04474(.A(\A[1] ), .B(new_n5476_), .Y(new_n5477_));
  XOR2   g04475(.A(\A[1] ), .B(new_n5476_), .Y(new_n5478_));
  INV    g04476(.A(\A[1] ), .Y(new_n5479_));
  OAI21  g04477(.A0(new_n5479_), .A1(\A[0] ), .B0(\A[2] ), .Y(new_n5480_));
  OAI22  g04478(.A0(new_n5480_), .A1(new_n5477_), .B0(new_n5478_), .B1(\A[2] ), .Y(new_n5481_));
  INV    g04479(.A(\A[2] ), .Y(new_n5482_));
  NAND2  g04480(.A(new_n5479_), .B(\A[0] ), .Y(new_n5483_));
  XOR2   g04481(.A(\A[1] ), .B(\A[0] ), .Y(new_n5484_));
  AOI21  g04482(.A0(\A[1] ), .A1(new_n5476_), .B0(new_n5482_), .Y(new_n5485_));
  AOI221 g04483(.A0(new_n5485_), .A1(new_n5483_), .C0(new_n5475_), .B0(new_n5484_), .B1(new_n5482_), .Y(new_n5486_));
  AOI211 g04484(.A0(new_n5481_), .A1(new_n5475_), .B(new_n5486_), .C(new_n5474_), .Y(new_n5487_));
  AOI22  g04485(.A0(new_n5485_), .A1(new_n5483_), .B0(new_n5484_), .B1(new_n5482_), .Y(new_n5488_));
  OAI221 g04486(.A0(new_n5480_), .A1(new_n5477_), .C0(\A[6] ), .B0(new_n5478_), .B1(\A[2] ), .Y(new_n5489_));
  OAI21  g04487(.A0(new_n5488_), .A1(\A[6] ), .B0(new_n5489_), .Y(new_n5490_));
  AOI211 g04488(.A0(new_n5490_), .A1(new_n5474_), .B(new_n5467_), .C(new_n5487_), .Y(new_n5491_));
  NOR2   g04489(.A(new_n5471_), .B(\A[3] ), .Y(new_n5492_));
  OAI21  g04490(.A0(\A[4] ), .A1(new_n5469_), .B0(\A[5] ), .Y(new_n5493_));
  XOR2   g04491(.A(\A[4] ), .B(new_n5469_), .Y(new_n5494_));
  OAI22  g04492(.A0(new_n5494_), .A1(\A[5] ), .B0(new_n5493_), .B1(new_n5492_), .Y(new_n5495_));
  OAI211 g04493(.A0(new_n5488_), .A1(\A[6] ), .B0(new_n5489_), .B1(new_n5495_), .Y(new_n5496_));
  AOI21  g04494(.A0(new_n5481_), .A1(new_n5475_), .B0(new_n5486_), .Y(new_n5497_));
  OAI21  g04495(.A0(new_n5497_), .A1(new_n5495_), .B0(new_n5496_), .Y(new_n5498_));
  AOI21  g04496(.A0(new_n5498_), .A1(new_n5467_), .B0(new_n5491_), .Y(new_n5499_));
  XOR2   g04497(.A(new_n5499_), .B(new_n5460_), .Y(new_n5500_));
  AOI21  g04498(.A0(new_n5441_), .A1(new_n5440_), .B0(new_n5500_), .Y(new_n5501_));
  NAND3  g04499(.A(new_n5501_), .B(new_n5439_), .C(new_n5422_), .Y(new_n5502_));
  NAND3  g04500(.A(new_n5420_), .B(new_n5415_), .C(new_n5413_), .Y(new_n5503_));
  OAI21  g04501(.A0(new_n5402_), .A1(new_n5392_), .B0(new_n5409_), .Y(new_n5504_));
  AOI21  g04502(.A0(new_n5504_), .A1(new_n5503_), .B0(new_n5431_), .Y(new_n5505_));
  NAND3  g04503(.A(new_n5409_), .B(new_n5415_), .C(new_n5413_), .Y(new_n5506_));
  AOI21  g04504(.A0(new_n5437_), .A1(new_n5506_), .B0(new_n5298_), .Y(new_n5507_));
  INV    g04505(.A(new_n5501_), .Y(new_n5508_));
  OAI21  g04506(.A0(new_n5507_), .A1(new_n5505_), .B0(new_n5508_), .Y(new_n5509_));
  INV    g04507(.A(new_n5448_), .Y(new_n5510_));
  XOR2   g04508(.A(new_n5455_), .B(new_n5510_), .Y(new_n5511_));
  XOR2   g04509(.A(new_n5459_), .B(new_n5457_), .Y(new_n5512_));
  NOR2   g04510(.A(new_n5455_), .B(new_n5448_), .Y(new_n5513_));
  NOR2   g04511(.A(new_n5459_), .B(new_n5457_), .Y(new_n5514_));
  AOI21  g04512(.A0(new_n5513_), .A1(new_n5512_), .B0(new_n5514_), .Y(new_n5515_));
  XOR2   g04513(.A(new_n5513_), .B(new_n5512_), .Y(new_n5516_));
  OAI21  g04514(.A0(new_n5515_), .A1(new_n5511_), .B0(new_n5516_), .Y(new_n5517_));
  INV    g04515(.A(new_n5515_), .Y(new_n5518_));
  AOI211 g04516(.A0(new_n5516_), .A1(new_n5518_), .B(new_n5499_), .C(new_n5511_), .Y(new_n5519_));
  NOR2   g04517(.A(new_n5462_), .B(new_n5464_), .Y(new_n5520_));
  AOI21  g04518(.A0(new_n5466_), .A1(\A[999] ), .B0(new_n5520_), .Y(new_n5521_));
  NOR2   g04519(.A(new_n5471_), .B(new_n5469_), .Y(new_n5522_));
  AOI21  g04520(.A0(new_n5473_), .A1(\A[5] ), .B0(new_n5522_), .Y(new_n5523_));
  NOR2   g04521(.A(new_n5479_), .B(new_n5476_), .Y(new_n5524_));
  AOI21  g04522(.A0(new_n5484_), .A1(\A[2] ), .B0(new_n5524_), .Y(new_n5525_));
  XOR2   g04523(.A(new_n5525_), .B(new_n5523_), .Y(new_n5526_));
  NOR2   g04524(.A(new_n5488_), .B(new_n5475_), .Y(new_n5527_));
  AOI211 g04525(.A0(new_n5490_), .A1(new_n5495_), .B(new_n5526_), .C(new_n5527_), .Y(new_n5528_));
  NAND2  g04526(.A(new_n5481_), .B(\A[6] ), .Y(new_n5529_));
  OAI21  g04527(.A0(new_n5497_), .A1(new_n5474_), .B0(new_n5529_), .Y(new_n5530_));
  AOI21  g04528(.A0(new_n5530_), .A1(new_n5526_), .B0(new_n5528_), .Y(new_n5531_));
  AOI21  g04529(.A0(new_n5490_), .A1(new_n5474_), .B0(new_n5487_), .Y(new_n5532_));
  NOR2   g04530(.A(new_n5532_), .B(new_n5467_), .Y(new_n5533_));
  NOR2   g04531(.A(new_n5533_), .B(new_n5531_), .Y(new_n5534_));
  NAND2  g04532(.A(\A[4] ), .B(\A[3] ), .Y(new_n5535_));
  OAI21  g04533(.A0(new_n5494_), .A1(new_n5468_), .B0(new_n5535_), .Y(new_n5536_));
  XOR2   g04534(.A(new_n5525_), .B(new_n5536_), .Y(new_n5537_));
  OAI211 g04535(.A0(new_n5497_), .A1(new_n5474_), .B0(new_n5537_), .B1(new_n5529_), .Y(new_n5538_));
  AOI21  g04536(.A0(new_n5490_), .A1(new_n5495_), .B0(new_n5527_), .Y(new_n5539_));
  OAI21  g04537(.A0(new_n5539_), .A1(new_n5537_), .B0(new_n5538_), .Y(new_n5540_));
  INV    g04538(.A(new_n5467_), .Y(new_n5541_));
  NAND2  g04539(.A(new_n5498_), .B(new_n5541_), .Y(new_n5542_));
  XOR2   g04540(.A(new_n5542_), .B(new_n5540_), .Y(new_n5543_));
  OAI21  g04541(.A0(new_n5542_), .A1(new_n5540_), .B0(new_n5521_), .Y(new_n5544_));
  OAI221 g04542(.A0(new_n5544_), .A1(new_n5534_), .C0(new_n5519_), .B0(new_n5543_), .B1(new_n5521_), .Y(new_n5545_));
  INV    g04543(.A(new_n5521_), .Y(new_n5546_));
  NAND2  g04544(.A(new_n5542_), .B(new_n5540_), .Y(new_n5547_));
  XOR2   g04545(.A(new_n5533_), .B(new_n5540_), .Y(new_n5548_));
  AOI21  g04546(.A0(new_n5533_), .A1(new_n5531_), .B0(new_n5546_), .Y(new_n5549_));
  AOI22  g04547(.A0(new_n5549_), .A1(new_n5547_), .B0(new_n5548_), .B1(new_n5546_), .Y(new_n5550_));
  OAI21  g04548(.A0(new_n5550_), .A1(new_n5519_), .B0(new_n5545_), .Y(new_n5551_));
  NAND2  g04549(.A(new_n5551_), .B(new_n5517_), .Y(new_n5552_));
  INV    g04550(.A(new_n5517_), .Y(new_n5553_));
  AOI221 g04551(.A0(new_n5549_), .A1(new_n5547_), .C0(new_n5519_), .B0(new_n5548_), .B1(new_n5546_), .Y(new_n5554_));
  NOR2   g04552(.A(new_n5532_), .B(new_n5541_), .Y(new_n5555_));
  OAI21  g04553(.A0(new_n5555_), .A1(new_n5491_), .B0(new_n5460_), .Y(new_n5556_));
  NOR2   g04554(.A(new_n5550_), .B(new_n5556_), .Y(new_n5557_));
  OAI21  g04555(.A0(new_n5557_), .A1(new_n5554_), .B0(new_n5553_), .Y(new_n5558_));
  NAND2  g04556(.A(new_n5558_), .B(new_n5552_), .Y(new_n5559_));
  AOI21  g04557(.A0(new_n5509_), .A1(new_n5502_), .B0(new_n5559_), .Y(new_n5560_));
  OAI221 g04558(.A0(new_n5544_), .A1(new_n5534_), .C0(new_n5556_), .B0(new_n5543_), .B1(new_n5521_), .Y(new_n5561_));
  OAI22  g04559(.A0(new_n5544_), .A1(new_n5534_), .B0(new_n5543_), .B1(new_n5521_), .Y(new_n5562_));
  NAND2  g04560(.A(new_n5562_), .B(new_n5519_), .Y(new_n5563_));
  AOI21  g04561(.A0(new_n5563_), .A1(new_n5561_), .B0(new_n5517_), .Y(new_n5564_));
  AOI21  g04562(.A0(new_n5551_), .A1(new_n5517_), .B0(new_n5564_), .Y(new_n5565_));
  AOI21  g04563(.A0(new_n5438_), .A1(new_n5431_), .B0(new_n5501_), .Y(new_n5566_));
  NAND2  g04564(.A(new_n5566_), .B(new_n5422_), .Y(new_n5567_));
  OAI21  g04565(.A0(new_n5507_), .A1(new_n5505_), .B0(new_n5501_), .Y(new_n5568_));
  AOI21  g04566(.A0(new_n5568_), .A1(new_n5567_), .B0(new_n5565_), .Y(new_n5569_));
  NOR2   g04567(.A(new_n5569_), .B(new_n5560_), .Y(new_n5570_));
  INV    g04568(.A(\A[45] ), .Y(new_n5571_));
  INV    g04569(.A(\A[43] ), .Y(new_n5572_));
  NAND2  g04570(.A(\A[44] ), .B(new_n5572_), .Y(new_n5573_));
  INV    g04571(.A(\A[44] ), .Y(new_n5574_));
  AOI21  g04572(.A0(new_n5574_), .A1(\A[43] ), .B0(new_n5571_), .Y(new_n5575_));
  XOR2   g04573(.A(\A[44] ), .B(\A[43] ), .Y(new_n5576_));
  AOI22  g04574(.A0(new_n5576_), .A1(new_n5571_), .B0(new_n5575_), .B1(new_n5573_), .Y(new_n5577_));
  INV    g04575(.A(\A[48] ), .Y(new_n5578_));
  INV    g04576(.A(\A[46] ), .Y(new_n5579_));
  NAND2  g04577(.A(\A[47] ), .B(new_n5579_), .Y(new_n5580_));
  INV    g04578(.A(\A[47] ), .Y(new_n5581_));
  AOI21  g04579(.A0(new_n5581_), .A1(\A[46] ), .B0(new_n5578_), .Y(new_n5582_));
  XOR2   g04580(.A(\A[47] ), .B(\A[46] ), .Y(new_n5583_));
  AOI22  g04581(.A0(new_n5583_), .A1(new_n5578_), .B0(new_n5582_), .B1(new_n5580_), .Y(new_n5584_));
  NOR2   g04582(.A(new_n5584_), .B(new_n5577_), .Y(new_n5585_));
  XOR2   g04583(.A(\A[47] ), .B(new_n5579_), .Y(new_n5586_));
  NAND2  g04584(.A(\A[47] ), .B(\A[46] ), .Y(new_n5587_));
  OAI21  g04585(.A0(new_n5586_), .A1(new_n5578_), .B0(new_n5587_), .Y(new_n5588_));
  NOR2   g04586(.A(new_n5574_), .B(new_n5572_), .Y(new_n5589_));
  AOI21  g04587(.A0(new_n5576_), .A1(\A[45] ), .B0(new_n5589_), .Y(new_n5590_));
  XOR2   g04588(.A(new_n5590_), .B(new_n5588_), .Y(new_n5591_));
  XOR2   g04589(.A(new_n5591_), .B(new_n5585_), .Y(new_n5592_));
  XOR2   g04590(.A(new_n5584_), .B(new_n5577_), .Y(new_n5593_));
  NOR2   g04591(.A(new_n5574_), .B(\A[43] ), .Y(new_n5594_));
  OAI21  g04592(.A0(\A[44] ), .A1(new_n5572_), .B0(\A[45] ), .Y(new_n5595_));
  XOR2   g04593(.A(\A[44] ), .B(new_n5572_), .Y(new_n5596_));
  OAI22  g04594(.A0(new_n5596_), .A1(\A[45] ), .B0(new_n5595_), .B1(new_n5594_), .Y(new_n5597_));
  NOR2   g04595(.A(new_n5581_), .B(\A[46] ), .Y(new_n5598_));
  OAI21  g04596(.A0(\A[47] ), .A1(new_n5579_), .B0(\A[48] ), .Y(new_n5599_));
  OAI22  g04597(.A0(new_n5586_), .A1(\A[48] ), .B0(new_n5599_), .B1(new_n5598_), .Y(new_n5600_));
  NAND2  g04598(.A(new_n5600_), .B(new_n5597_), .Y(new_n5601_));
  NAND2  g04599(.A(\A[44] ), .B(\A[43] ), .Y(new_n5602_));
  OAI21  g04600(.A0(new_n5596_), .A1(new_n5571_), .B0(new_n5602_), .Y(new_n5603_));
  NAND2  g04601(.A(new_n5603_), .B(new_n5588_), .Y(new_n5604_));
  OAI21  g04602(.A0(new_n5591_), .A1(new_n5601_), .B0(new_n5604_), .Y(new_n5605_));
  AOI21  g04603(.A0(new_n5605_), .A1(new_n5593_), .B0(new_n5592_), .Y(new_n5606_));
  NAND2  g04604(.A(\A[53] ), .B(\A[52] ), .Y(new_n5607_));
  XOR2   g04605(.A(\A[53] ), .B(\A[52] ), .Y(new_n5608_));
  NAND2  g04606(.A(new_n5608_), .B(\A[54] ), .Y(new_n5609_));
  NAND2  g04607(.A(new_n5609_), .B(new_n5607_), .Y(new_n5610_));
  NAND2  g04608(.A(\A[50] ), .B(\A[49] ), .Y(new_n5611_));
  XOR2   g04609(.A(\A[50] ), .B(\A[49] ), .Y(new_n5612_));
  NAND2  g04610(.A(new_n5612_), .B(\A[51] ), .Y(new_n5613_));
  NAND2  g04611(.A(new_n5613_), .B(new_n5611_), .Y(new_n5614_));
  XOR2   g04612(.A(new_n5614_), .B(new_n5610_), .Y(new_n5615_));
  INV    g04613(.A(\A[51] ), .Y(new_n5616_));
  INV    g04614(.A(\A[49] ), .Y(new_n5617_));
  NAND2  g04615(.A(\A[50] ), .B(new_n5617_), .Y(new_n5618_));
  INV    g04616(.A(\A[50] ), .Y(new_n5619_));
  AOI21  g04617(.A0(new_n5619_), .A1(\A[49] ), .B0(new_n5616_), .Y(new_n5620_));
  AOI22  g04618(.A0(new_n5620_), .A1(new_n5618_), .B0(new_n5612_), .B1(new_n5616_), .Y(new_n5621_));
  INV    g04619(.A(\A[54] ), .Y(new_n5622_));
  INV    g04620(.A(\A[52] ), .Y(new_n5623_));
  NAND2  g04621(.A(\A[53] ), .B(new_n5623_), .Y(new_n5624_));
  INV    g04622(.A(\A[53] ), .Y(new_n5625_));
  AOI21  g04623(.A0(new_n5625_), .A1(\A[52] ), .B0(new_n5622_), .Y(new_n5626_));
  AOI22  g04624(.A0(new_n5626_), .A1(new_n5624_), .B0(new_n5608_), .B1(new_n5622_), .Y(new_n5627_));
  NOR2   g04625(.A(new_n5627_), .B(new_n5621_), .Y(new_n5628_));
  AOI22  g04626(.A0(new_n5613_), .A1(new_n5611_), .B0(new_n5609_), .B1(new_n5607_), .Y(new_n5629_));
  AOI21  g04627(.A0(new_n5628_), .A1(new_n5615_), .B0(new_n5629_), .Y(new_n5630_));
  XOR2   g04628(.A(new_n5628_), .B(new_n5615_), .Y(new_n5631_));
  NOR2   g04629(.A(new_n5619_), .B(\A[49] ), .Y(new_n5632_));
  OAI21  g04630(.A0(\A[50] ), .A1(new_n5617_), .B0(\A[51] ), .Y(new_n5633_));
  NAND2  g04631(.A(new_n5612_), .B(new_n5616_), .Y(new_n5634_));
  OAI21  g04632(.A0(new_n5633_), .A1(new_n5632_), .B0(new_n5634_), .Y(new_n5635_));
  XOR2   g04633(.A(new_n5627_), .B(new_n5635_), .Y(new_n5636_));
  NOR2   g04634(.A(new_n5625_), .B(\A[52] ), .Y(new_n5637_));
  OAI21  g04635(.A0(\A[53] ), .A1(new_n5623_), .B0(\A[54] ), .Y(new_n5638_));
  NAND2  g04636(.A(new_n5608_), .B(new_n5622_), .Y(new_n5639_));
  OAI21  g04637(.A0(new_n5638_), .A1(new_n5637_), .B0(new_n5639_), .Y(new_n5640_));
  NAND4  g04638(.A(new_n5640_), .B(new_n5635_), .C(new_n5614_), .D(new_n5610_), .Y(new_n5641_));
  NAND4  g04639(.A(new_n5603_), .B(new_n5588_), .C(new_n5600_), .D(new_n5597_), .Y(new_n5642_));
  XOR2   g04640(.A(new_n5627_), .B(new_n5621_), .Y(new_n5643_));
  NAND4  g04641(.A(new_n5643_), .B(new_n5642_), .C(new_n5641_), .D(new_n5593_), .Y(new_n5644_));
  OAI211 g04642(.A0(new_n5636_), .A1(new_n5630_), .B0(new_n5644_), .B1(new_n5631_), .Y(new_n5645_));
  NOR2   g04643(.A(new_n5619_), .B(new_n5617_), .Y(new_n5646_));
  AOI21  g04644(.A0(new_n5612_), .A1(\A[51] ), .B0(new_n5646_), .Y(new_n5647_));
  XOR2   g04645(.A(new_n5647_), .B(new_n5610_), .Y(new_n5648_));
  XOR2   g04646(.A(new_n5628_), .B(new_n5648_), .Y(new_n5649_));
  XOR2   g04647(.A(new_n5584_), .B(new_n5597_), .Y(new_n5650_));
  NOR2   g04648(.A(new_n5625_), .B(new_n5623_), .Y(new_n5651_));
  AOI21  g04649(.A0(new_n5608_), .A1(\A[54] ), .B0(new_n5651_), .Y(new_n5652_));
  NOR4   g04650(.A(new_n5627_), .B(new_n5621_), .C(new_n5647_), .D(new_n5652_), .Y(new_n5653_));
  NOR2   g04651(.A(new_n5581_), .B(new_n5579_), .Y(new_n5654_));
  AOI21  g04652(.A0(new_n5583_), .A1(\A[48] ), .B0(new_n5654_), .Y(new_n5655_));
  NOR4   g04653(.A(new_n5590_), .B(new_n5655_), .C(new_n5584_), .D(new_n5577_), .Y(new_n5656_));
  NOR4   g04654(.A(new_n5636_), .B(new_n5656_), .C(new_n5653_), .D(new_n5650_), .Y(new_n5657_));
  AOI221 g04655(.A0(new_n5612_), .A1(\A[51] ), .C0(new_n5646_), .B0(new_n5609_), .B1(new_n5607_), .Y(new_n5658_));
  AOI221 g04656(.A0(new_n5613_), .A1(new_n5611_), .C0(new_n5651_), .B0(new_n5608_), .B1(\A[54] ), .Y(new_n5659_));
  OAI211 g04657(.A0(new_n5659_), .A1(new_n5658_), .B0(new_n5640_), .B1(new_n5635_), .Y(new_n5660_));
  NAND2  g04658(.A(new_n5614_), .B(new_n5610_), .Y(new_n5661_));
  AOI21  g04659(.A0(new_n5661_), .A1(new_n5660_), .B0(new_n5636_), .Y(new_n5662_));
  OAI21  g04660(.A0(new_n5662_), .A1(new_n5649_), .B0(new_n5657_), .Y(new_n5663_));
  AOI21  g04661(.A0(new_n5663_), .A1(new_n5645_), .B0(new_n5606_), .Y(new_n5664_));
  XOR2   g04662(.A(new_n5591_), .B(new_n5601_), .Y(new_n5665_));
  XOR2   g04663(.A(new_n5590_), .B(new_n5655_), .Y(new_n5666_));
  NOR2   g04664(.A(new_n5590_), .B(new_n5655_), .Y(new_n5667_));
  AOI21  g04665(.A0(new_n5666_), .A1(new_n5585_), .B0(new_n5667_), .Y(new_n5668_));
  OAI21  g04666(.A0(new_n5668_), .A1(new_n5650_), .B0(new_n5665_), .Y(new_n5669_));
  OAI21  g04667(.A0(new_n5662_), .A1(new_n5649_), .B0(new_n5644_), .Y(new_n5670_));
  NOR2   g04668(.A(new_n5636_), .B(new_n5650_), .Y(new_n5671_));
  OAI211 g04669(.A0(new_n5640_), .A1(new_n5635_), .B0(new_n5614_), .B1(new_n5610_), .Y(new_n5672_));
  NAND4  g04670(.A(new_n5672_), .B(new_n5671_), .C(new_n5642_), .D(new_n5631_), .Y(new_n5673_));
  AOI21  g04671(.A0(new_n5673_), .A1(new_n5670_), .B0(new_n5669_), .Y(new_n5674_));
  NOR2   g04672(.A(new_n5636_), .B(new_n5653_), .Y(new_n5675_));
  XOR2   g04673(.A(new_n5584_), .B(new_n5577_), .Y(new_n5676_));
  XOR2   g04674(.A(new_n5676_), .B(new_n5675_), .Y(new_n5677_));
  INV    g04675(.A(\A[39] ), .Y(new_n5678_));
  INV    g04676(.A(\A[38] ), .Y(new_n5679_));
  NAND2  g04677(.A(new_n5679_), .B(\A[37] ), .Y(new_n5680_));
  INV    g04678(.A(\A[37] ), .Y(new_n5681_));
  AOI21  g04679(.A0(\A[38] ), .A1(new_n5681_), .B0(new_n5678_), .Y(new_n5682_));
  XOR2   g04680(.A(\A[38] ), .B(\A[37] ), .Y(new_n5683_));
  AOI22  g04681(.A0(new_n5683_), .A1(new_n5678_), .B0(new_n5682_), .B1(new_n5680_), .Y(new_n5684_));
  INV    g04682(.A(\A[42] ), .Y(new_n5685_));
  INV    g04683(.A(\A[41] ), .Y(new_n5686_));
  NAND2  g04684(.A(new_n5686_), .B(\A[40] ), .Y(new_n5687_));
  INV    g04685(.A(\A[40] ), .Y(new_n5688_));
  AOI21  g04686(.A0(\A[41] ), .A1(new_n5688_), .B0(new_n5685_), .Y(new_n5689_));
  XOR2   g04687(.A(\A[41] ), .B(\A[40] ), .Y(new_n5690_));
  AOI22  g04688(.A0(new_n5690_), .A1(new_n5685_), .B0(new_n5689_), .B1(new_n5687_), .Y(new_n5691_));
  NOR2   g04689(.A(new_n5686_), .B(new_n5688_), .Y(new_n5692_));
  AOI21  g04690(.A0(new_n5690_), .A1(\A[42] ), .B0(new_n5692_), .Y(new_n5693_));
  NOR2   g04691(.A(new_n5679_), .B(new_n5681_), .Y(new_n5694_));
  AOI21  g04692(.A0(new_n5683_), .A1(\A[39] ), .B0(new_n5694_), .Y(new_n5695_));
  XOR2   g04693(.A(new_n5691_), .B(new_n5684_), .Y(new_n5696_));
  INV    g04694(.A(\A[33] ), .Y(new_n5697_));
  INV    g04695(.A(\A[32] ), .Y(new_n5698_));
  NAND2  g04696(.A(new_n5698_), .B(\A[31] ), .Y(new_n5699_));
  INV    g04697(.A(\A[31] ), .Y(new_n5700_));
  AOI21  g04698(.A0(\A[32] ), .A1(new_n5700_), .B0(new_n5697_), .Y(new_n5701_));
  XOR2   g04699(.A(\A[32] ), .B(\A[31] ), .Y(new_n5702_));
  AOI22  g04700(.A0(new_n5702_), .A1(new_n5697_), .B0(new_n5701_), .B1(new_n5699_), .Y(new_n5703_));
  INV    g04701(.A(\A[36] ), .Y(new_n5704_));
  INV    g04702(.A(\A[35] ), .Y(new_n5705_));
  NAND2  g04703(.A(new_n5705_), .B(\A[34] ), .Y(new_n5706_));
  INV    g04704(.A(\A[34] ), .Y(new_n5707_));
  AOI21  g04705(.A0(\A[35] ), .A1(new_n5707_), .B0(new_n5704_), .Y(new_n5708_));
  XOR2   g04706(.A(\A[35] ), .B(\A[34] ), .Y(new_n5709_));
  AOI22  g04707(.A0(new_n5709_), .A1(new_n5704_), .B0(new_n5708_), .B1(new_n5706_), .Y(new_n5710_));
  NOR2   g04708(.A(new_n5705_), .B(new_n5707_), .Y(new_n5711_));
  AOI21  g04709(.A0(new_n5709_), .A1(\A[36] ), .B0(new_n5711_), .Y(new_n5712_));
  NOR2   g04710(.A(new_n5698_), .B(new_n5700_), .Y(new_n5713_));
  AOI21  g04711(.A0(new_n5702_), .A1(\A[33] ), .B0(new_n5713_), .Y(new_n5714_));
  XOR2   g04712(.A(new_n5710_), .B(new_n5703_), .Y(new_n5715_));
  XOR2   g04713(.A(new_n5715_), .B(new_n5696_), .Y(new_n5716_));
  NAND2  g04714(.A(new_n5716_), .B(new_n5677_), .Y(new_n5717_));
  NOR3   g04715(.A(new_n5717_), .B(new_n5674_), .C(new_n5664_), .Y(new_n5718_));
  OAI21  g04716(.A0(new_n5636_), .A1(new_n5630_), .B0(new_n5631_), .Y(new_n5719_));
  XOR2   g04717(.A(new_n5719_), .B(new_n5644_), .Y(new_n5720_));
  NAND2  g04718(.A(new_n5720_), .B(new_n5669_), .Y(new_n5721_));
  NAND2  g04719(.A(new_n5673_), .B(new_n5670_), .Y(new_n5722_));
  NAND2  g04720(.A(new_n5722_), .B(new_n5606_), .Y(new_n5723_));
  NAND2  g04721(.A(new_n5643_), .B(new_n5641_), .Y(new_n5724_));
  XOR2   g04722(.A(new_n5676_), .B(new_n5724_), .Y(new_n5725_));
  NOR2   g04723(.A(\A[38] ), .B(new_n5681_), .Y(new_n5726_));
  OAI21  g04724(.A0(new_n5679_), .A1(\A[37] ), .B0(\A[39] ), .Y(new_n5727_));
  NAND2  g04725(.A(new_n5683_), .B(new_n5678_), .Y(new_n5728_));
  OAI21  g04726(.A0(new_n5727_), .A1(new_n5726_), .B0(new_n5728_), .Y(new_n5729_));
  XOR2   g04727(.A(new_n5691_), .B(new_n5729_), .Y(new_n5730_));
  XOR2   g04728(.A(new_n5715_), .B(new_n5730_), .Y(new_n5731_));
  NOR2   g04729(.A(new_n5731_), .B(new_n5725_), .Y(new_n5732_));
  AOI21  g04730(.A0(new_n5723_), .A1(new_n5721_), .B0(new_n5732_), .Y(new_n5733_));
  XOR2   g04731(.A(new_n5710_), .B(new_n5703_), .Y(new_n5734_));
  XOR2   g04732(.A(\A[35] ), .B(new_n5707_), .Y(new_n5735_));
  NAND2  g04733(.A(\A[35] ), .B(\A[34] ), .Y(new_n5736_));
  OAI21  g04734(.A0(new_n5735_), .A1(new_n5704_), .B0(new_n5736_), .Y(new_n5737_));
  XOR2   g04735(.A(new_n5714_), .B(new_n5737_), .Y(new_n5738_));
  NOR2   g04736(.A(\A[32] ), .B(new_n5700_), .Y(new_n5739_));
  OAI21  g04737(.A0(new_n5698_), .A1(\A[31] ), .B0(\A[33] ), .Y(new_n5740_));
  XOR2   g04738(.A(\A[32] ), .B(new_n5700_), .Y(new_n5741_));
  OAI22  g04739(.A0(new_n5741_), .A1(\A[33] ), .B0(new_n5740_), .B1(new_n5739_), .Y(new_n5742_));
  NOR2   g04740(.A(\A[35] ), .B(new_n5707_), .Y(new_n5743_));
  OAI21  g04741(.A0(new_n5705_), .A1(\A[34] ), .B0(\A[36] ), .Y(new_n5744_));
  OAI22  g04742(.A0(new_n5735_), .A1(\A[36] ), .B0(new_n5744_), .B1(new_n5743_), .Y(new_n5745_));
  NAND2  g04743(.A(new_n5745_), .B(new_n5742_), .Y(new_n5746_));
  NAND2  g04744(.A(\A[32] ), .B(\A[31] ), .Y(new_n5747_));
  OAI21  g04745(.A0(new_n5741_), .A1(new_n5697_), .B0(new_n5747_), .Y(new_n5748_));
  NAND2  g04746(.A(new_n5748_), .B(new_n5737_), .Y(new_n5749_));
  OAI21  g04747(.A0(new_n5746_), .A1(new_n5738_), .B0(new_n5749_), .Y(new_n5750_));
  NOR2   g04748(.A(new_n5710_), .B(new_n5703_), .Y(new_n5751_));
  XOR2   g04749(.A(new_n5751_), .B(new_n5738_), .Y(new_n5752_));
  AOI21  g04750(.A0(new_n5750_), .A1(new_n5734_), .B0(new_n5752_), .Y(new_n5753_));
  XOR2   g04751(.A(new_n5691_), .B(new_n5729_), .Y(new_n5754_));
  XOR2   g04752(.A(new_n5695_), .B(new_n5693_), .Y(new_n5755_));
  NOR2   g04753(.A(new_n5691_), .B(new_n5684_), .Y(new_n5756_));
  NAND2  g04754(.A(\A[41] ), .B(\A[40] ), .Y(new_n5757_));
  NAND2  g04755(.A(new_n5690_), .B(\A[42] ), .Y(new_n5758_));
  NAND2  g04756(.A(\A[38] ), .B(\A[37] ), .Y(new_n5759_));
  NAND2  g04757(.A(new_n5683_), .B(\A[39] ), .Y(new_n5760_));
  AOI22  g04758(.A0(new_n5760_), .A1(new_n5759_), .B0(new_n5758_), .B1(new_n5757_), .Y(new_n5761_));
  AOI21  g04759(.A0(new_n5756_), .A1(new_n5755_), .B0(new_n5761_), .Y(new_n5762_));
  XOR2   g04760(.A(new_n5756_), .B(new_n5755_), .Y(new_n5763_));
  XOR2   g04761(.A(new_n5691_), .B(new_n5684_), .Y(new_n5764_));
  NOR2   g04762(.A(\A[41] ), .B(new_n5688_), .Y(new_n5765_));
  OAI21  g04763(.A0(new_n5686_), .A1(\A[40] ), .B0(\A[42] ), .Y(new_n5766_));
  NAND2  g04764(.A(new_n5690_), .B(new_n5685_), .Y(new_n5767_));
  OAI21  g04765(.A0(new_n5766_), .A1(new_n5765_), .B0(new_n5767_), .Y(new_n5768_));
  NAND2  g04766(.A(new_n5758_), .B(new_n5757_), .Y(new_n5769_));
  NAND2  g04767(.A(new_n5760_), .B(new_n5759_), .Y(new_n5770_));
  NAND4  g04768(.A(new_n5770_), .B(new_n5769_), .C(new_n5768_), .D(new_n5729_), .Y(new_n5771_));
  NAND4  g04769(.A(new_n5748_), .B(new_n5737_), .C(new_n5745_), .D(new_n5742_), .Y(new_n5772_));
  NAND4  g04770(.A(new_n5772_), .B(new_n5734_), .C(new_n5771_), .D(new_n5764_), .Y(new_n5773_));
  OAI211 g04771(.A0(new_n5762_), .A1(new_n5754_), .B0(new_n5773_), .B1(new_n5763_), .Y(new_n5774_));
  XOR2   g04772(.A(new_n5695_), .B(new_n5769_), .Y(new_n5775_));
  XOR2   g04773(.A(new_n5756_), .B(new_n5775_), .Y(new_n5776_));
  NOR4   g04774(.A(new_n5695_), .B(new_n5693_), .C(new_n5691_), .D(new_n5684_), .Y(new_n5777_));
  XOR2   g04775(.A(new_n5710_), .B(new_n5742_), .Y(new_n5778_));
  NOR4   g04776(.A(new_n5714_), .B(new_n5712_), .C(new_n5710_), .D(new_n5703_), .Y(new_n5779_));
  NOR4   g04777(.A(new_n5779_), .B(new_n5778_), .C(new_n5777_), .D(new_n5754_), .Y(new_n5780_));
  AOI221 g04778(.A0(new_n5758_), .A1(new_n5757_), .C0(new_n5694_), .B0(new_n5683_), .B1(\A[39] ), .Y(new_n5781_));
  AOI221 g04779(.A0(new_n5760_), .A1(new_n5759_), .C0(new_n5692_), .B0(new_n5690_), .B1(\A[42] ), .Y(new_n5782_));
  OAI211 g04780(.A0(new_n5782_), .A1(new_n5781_), .B0(new_n5768_), .B1(new_n5729_), .Y(new_n5783_));
  NAND2  g04781(.A(new_n5770_), .B(new_n5769_), .Y(new_n5784_));
  AOI21  g04782(.A0(new_n5784_), .A1(new_n5783_), .B0(new_n5754_), .Y(new_n5785_));
  OAI21  g04783(.A0(new_n5785_), .A1(new_n5776_), .B0(new_n5780_), .Y(new_n5786_));
  AOI21  g04784(.A0(new_n5786_), .A1(new_n5774_), .B0(new_n5753_), .Y(new_n5787_));
  NOR2   g04785(.A(new_n5785_), .B(new_n5776_), .Y(new_n5788_));
  NAND4  g04786(.A(new_n5734_), .B(new_n5763_), .C(new_n5762_), .D(new_n5764_), .Y(new_n5789_));
  OAI21  g04787(.A0(new_n5762_), .A1(new_n5754_), .B0(new_n5772_), .Y(new_n5790_));
  OAI22  g04788(.A0(new_n5790_), .A1(new_n5789_), .B0(new_n5788_), .B1(new_n5780_), .Y(new_n5791_));
  AOI21  g04789(.A0(new_n5791_), .A1(new_n5753_), .B0(new_n5787_), .Y(new_n5792_));
  OAI21  g04790(.A0(new_n5733_), .A1(new_n5718_), .B0(new_n5792_), .Y(new_n5793_));
  XOR2   g04791(.A(new_n5788_), .B(new_n5773_), .Y(new_n5794_));
  NAND2  g04792(.A(new_n5791_), .B(new_n5753_), .Y(new_n5795_));
  OAI21  g04793(.A0(new_n5794_), .A1(new_n5753_), .B0(new_n5795_), .Y(new_n5796_));
  NOR3   g04794(.A(new_n5732_), .B(new_n5674_), .C(new_n5664_), .Y(new_n5797_));
  AOI21  g04795(.A0(new_n5723_), .A1(new_n5721_), .B0(new_n5717_), .Y(new_n5798_));
  OAI21  g04796(.A0(new_n5798_), .A1(new_n5797_), .B0(new_n5796_), .Y(new_n5799_));
  NAND2  g04797(.A(new_n5799_), .B(new_n5793_), .Y(new_n5800_));
  INV    g04798(.A(\A[56] ), .Y(new_n5801_));
  NOR2   g04799(.A(new_n5801_), .B(\A[55] ), .Y(new_n5802_));
  INV    g04800(.A(\A[55] ), .Y(new_n5803_));
  OAI21  g04801(.A0(\A[56] ), .A1(new_n5803_), .B0(\A[57] ), .Y(new_n5804_));
  XOR2   g04802(.A(\A[56] ), .B(new_n5803_), .Y(new_n5805_));
  OAI22  g04803(.A0(new_n5805_), .A1(\A[57] ), .B0(new_n5804_), .B1(new_n5802_), .Y(new_n5806_));
  INV    g04804(.A(\A[59] ), .Y(new_n5807_));
  NOR2   g04805(.A(new_n5807_), .B(\A[58] ), .Y(new_n5808_));
  INV    g04806(.A(\A[58] ), .Y(new_n5809_));
  OAI21  g04807(.A0(\A[59] ), .A1(new_n5809_), .B0(\A[60] ), .Y(new_n5810_));
  XOR2   g04808(.A(\A[59] ), .B(new_n5809_), .Y(new_n5811_));
  OAI22  g04809(.A0(new_n5811_), .A1(\A[60] ), .B0(new_n5810_), .B1(new_n5808_), .Y(new_n5812_));
  NAND2  g04810(.A(new_n5812_), .B(new_n5806_), .Y(new_n5813_));
  INV    g04811(.A(\A[60] ), .Y(new_n5814_));
  NAND2  g04812(.A(\A[59] ), .B(\A[58] ), .Y(new_n5815_));
  OAI21  g04813(.A0(new_n5811_), .A1(new_n5814_), .B0(new_n5815_), .Y(new_n5816_));
  XOR2   g04814(.A(\A[56] ), .B(\A[55] ), .Y(new_n5817_));
  NOR2   g04815(.A(new_n5801_), .B(new_n5803_), .Y(new_n5818_));
  AOI21  g04816(.A0(new_n5817_), .A1(\A[57] ), .B0(new_n5818_), .Y(new_n5819_));
  XOR2   g04817(.A(new_n5819_), .B(new_n5816_), .Y(new_n5820_));
  XOR2   g04818(.A(new_n5820_), .B(new_n5813_), .Y(new_n5821_));
  NAND2  g04819(.A(\A[59] ), .B(new_n5809_), .Y(new_n5822_));
  AOI21  g04820(.A0(new_n5807_), .A1(\A[58] ), .B0(new_n5814_), .Y(new_n5823_));
  XOR2   g04821(.A(\A[59] ), .B(\A[58] ), .Y(new_n5824_));
  AOI22  g04822(.A0(new_n5824_), .A1(new_n5814_), .B0(new_n5823_), .B1(new_n5822_), .Y(new_n5825_));
  XOR2   g04823(.A(new_n5825_), .B(new_n5806_), .Y(new_n5826_));
  INV    g04824(.A(\A[57] ), .Y(new_n5827_));
  NAND2  g04825(.A(\A[56] ), .B(new_n5803_), .Y(new_n5828_));
  AOI21  g04826(.A0(new_n5801_), .A1(\A[55] ), .B0(new_n5827_), .Y(new_n5829_));
  AOI22  g04827(.A0(new_n5817_), .A1(new_n5827_), .B0(new_n5829_), .B1(new_n5828_), .Y(new_n5830_));
  NOR2   g04828(.A(new_n5825_), .B(new_n5830_), .Y(new_n5831_));
  NOR2   g04829(.A(new_n5807_), .B(new_n5809_), .Y(new_n5832_));
  AOI21  g04830(.A0(new_n5824_), .A1(\A[60] ), .B0(new_n5832_), .Y(new_n5833_));
  XOR2   g04831(.A(new_n5819_), .B(new_n5833_), .Y(new_n5834_));
  NOR2   g04832(.A(new_n5819_), .B(new_n5833_), .Y(new_n5835_));
  AOI21  g04833(.A0(new_n5834_), .A1(new_n5831_), .B0(new_n5835_), .Y(new_n5836_));
  OAI21  g04834(.A0(new_n5836_), .A1(new_n5826_), .B0(new_n5821_), .Y(new_n5837_));
  XOR2   g04835(.A(new_n5825_), .B(new_n5830_), .Y(new_n5838_));
  NAND2  g04836(.A(\A[65] ), .B(\A[64] ), .Y(new_n5839_));
  XOR2   g04837(.A(\A[65] ), .B(\A[64] ), .Y(new_n5840_));
  NAND2  g04838(.A(new_n5840_), .B(\A[66] ), .Y(new_n5841_));
  NAND2  g04839(.A(new_n5841_), .B(new_n5839_), .Y(new_n5842_));
  NAND2  g04840(.A(\A[62] ), .B(\A[61] ), .Y(new_n5843_));
  XOR2   g04841(.A(\A[62] ), .B(\A[61] ), .Y(new_n5844_));
  NAND2  g04842(.A(new_n5844_), .B(\A[63] ), .Y(new_n5845_));
  NAND2  g04843(.A(new_n5845_), .B(new_n5843_), .Y(new_n5846_));
  INV    g04844(.A(\A[62] ), .Y(new_n5847_));
  NOR2   g04845(.A(new_n5847_), .B(\A[61] ), .Y(new_n5848_));
  INV    g04846(.A(\A[61] ), .Y(new_n5849_));
  OAI21  g04847(.A0(\A[62] ), .A1(new_n5849_), .B0(\A[63] ), .Y(new_n5850_));
  INV    g04848(.A(\A[63] ), .Y(new_n5851_));
  NAND2  g04849(.A(new_n5844_), .B(new_n5851_), .Y(new_n5852_));
  OAI21  g04850(.A0(new_n5850_), .A1(new_n5848_), .B0(new_n5852_), .Y(new_n5853_));
  INV    g04851(.A(\A[65] ), .Y(new_n5854_));
  NOR2   g04852(.A(new_n5854_), .B(\A[64] ), .Y(new_n5855_));
  INV    g04853(.A(\A[64] ), .Y(new_n5856_));
  OAI21  g04854(.A0(\A[65] ), .A1(new_n5856_), .B0(\A[66] ), .Y(new_n5857_));
  INV    g04855(.A(\A[66] ), .Y(new_n5858_));
  NAND2  g04856(.A(new_n5840_), .B(new_n5858_), .Y(new_n5859_));
  OAI21  g04857(.A0(new_n5857_), .A1(new_n5855_), .B0(new_n5859_), .Y(new_n5860_));
  NAND4  g04858(.A(new_n5860_), .B(new_n5853_), .C(new_n5846_), .D(new_n5842_), .Y(new_n5861_));
  NAND2  g04859(.A(\A[56] ), .B(\A[55] ), .Y(new_n5862_));
  OAI21  g04860(.A0(new_n5805_), .A1(new_n5827_), .B0(new_n5862_), .Y(new_n5863_));
  NAND4  g04861(.A(new_n5863_), .B(new_n5816_), .C(new_n5812_), .D(new_n5806_), .Y(new_n5864_));
  NAND2  g04862(.A(\A[62] ), .B(new_n5849_), .Y(new_n5865_));
  AOI21  g04863(.A0(new_n5847_), .A1(\A[61] ), .B0(new_n5851_), .Y(new_n5866_));
  AOI22  g04864(.A0(new_n5866_), .A1(new_n5865_), .B0(new_n5844_), .B1(new_n5851_), .Y(new_n5867_));
  NAND2  g04865(.A(\A[65] ), .B(new_n5856_), .Y(new_n5868_));
  AOI21  g04866(.A0(new_n5854_), .A1(\A[64] ), .B0(new_n5858_), .Y(new_n5869_));
  AOI22  g04867(.A0(new_n5869_), .A1(new_n5868_), .B0(new_n5840_), .B1(new_n5858_), .Y(new_n5870_));
  XOR2   g04868(.A(new_n5870_), .B(new_n5867_), .Y(new_n5871_));
  NAND4  g04869(.A(new_n5871_), .B(new_n5864_), .C(new_n5861_), .D(new_n5838_), .Y(new_n5872_));
  XOR2   g04870(.A(new_n5846_), .B(new_n5842_), .Y(new_n5873_));
  NOR2   g04871(.A(new_n5870_), .B(new_n5867_), .Y(new_n5874_));
  AOI22  g04872(.A0(new_n5845_), .A1(new_n5843_), .B0(new_n5841_), .B1(new_n5839_), .Y(new_n5875_));
  AOI21  g04873(.A0(new_n5874_), .A1(new_n5873_), .B0(new_n5875_), .Y(new_n5876_));
  XOR2   g04874(.A(new_n5874_), .B(new_n5873_), .Y(new_n5877_));
  XOR2   g04875(.A(new_n5870_), .B(new_n5853_), .Y(new_n5878_));
  OAI21  g04876(.A0(new_n5878_), .A1(new_n5876_), .B0(new_n5877_), .Y(new_n5879_));
  XOR2   g04877(.A(new_n5879_), .B(new_n5872_), .Y(new_n5880_));
  NAND2  g04878(.A(new_n5860_), .B(new_n5853_), .Y(new_n5881_));
  XOR2   g04879(.A(new_n5881_), .B(new_n5873_), .Y(new_n5882_));
  NOR2   g04880(.A(new_n5847_), .B(new_n5849_), .Y(new_n5883_));
  AOI221 g04881(.A0(new_n5844_), .A1(\A[63] ), .C0(new_n5883_), .B0(new_n5841_), .B1(new_n5839_), .Y(new_n5884_));
  NOR2   g04882(.A(new_n5854_), .B(new_n5856_), .Y(new_n5885_));
  AOI221 g04883(.A0(new_n5845_), .A1(new_n5843_), .C0(new_n5885_), .B0(new_n5840_), .B1(\A[66] ), .Y(new_n5886_));
  OAI211 g04884(.A0(new_n5886_), .A1(new_n5884_), .B0(new_n5860_), .B1(new_n5853_), .Y(new_n5887_));
  NAND2  g04885(.A(new_n5846_), .B(new_n5842_), .Y(new_n5888_));
  AOI21  g04886(.A0(new_n5888_), .A1(new_n5887_), .B0(new_n5878_), .Y(new_n5889_));
  OAI21  g04887(.A0(new_n5889_), .A1(new_n5882_), .B0(new_n5872_), .Y(new_n5890_));
  NOR2   g04888(.A(new_n5878_), .B(new_n5826_), .Y(new_n5891_));
  OAI211 g04889(.A0(new_n5860_), .A1(new_n5853_), .B0(new_n5846_), .B1(new_n5842_), .Y(new_n5892_));
  NAND4  g04890(.A(new_n5892_), .B(new_n5891_), .C(new_n5864_), .D(new_n5877_), .Y(new_n5893_));
  AOI21  g04891(.A0(new_n5893_), .A1(new_n5890_), .B0(new_n5837_), .Y(new_n5894_));
  AOI21  g04892(.A0(new_n5880_), .A1(new_n5837_), .B0(new_n5894_), .Y(new_n5895_));
  INV    g04893(.A(\A[69] ), .Y(new_n5896_));
  INV    g04894(.A(\A[67] ), .Y(new_n5897_));
  NAND2  g04895(.A(\A[68] ), .B(new_n5897_), .Y(new_n5898_));
  INV    g04896(.A(\A[68] ), .Y(new_n5899_));
  AOI21  g04897(.A0(new_n5899_), .A1(\A[67] ), .B0(new_n5896_), .Y(new_n5900_));
  XOR2   g04898(.A(\A[68] ), .B(\A[67] ), .Y(new_n5901_));
  AOI22  g04899(.A0(new_n5901_), .A1(new_n5896_), .B0(new_n5900_), .B1(new_n5898_), .Y(new_n5902_));
  INV    g04900(.A(\A[72] ), .Y(new_n5903_));
  INV    g04901(.A(\A[70] ), .Y(new_n5904_));
  NAND2  g04902(.A(\A[71] ), .B(new_n5904_), .Y(new_n5905_));
  INV    g04903(.A(\A[71] ), .Y(new_n5906_));
  AOI21  g04904(.A0(new_n5906_), .A1(\A[70] ), .B0(new_n5903_), .Y(new_n5907_));
  XOR2   g04905(.A(\A[71] ), .B(\A[70] ), .Y(new_n5908_));
  AOI22  g04906(.A0(new_n5908_), .A1(new_n5903_), .B0(new_n5907_), .B1(new_n5905_), .Y(new_n5909_));
  NOR2   g04907(.A(new_n5909_), .B(new_n5902_), .Y(new_n5910_));
  XOR2   g04908(.A(\A[71] ), .B(new_n5904_), .Y(new_n5911_));
  NAND2  g04909(.A(\A[71] ), .B(\A[70] ), .Y(new_n5912_));
  OAI21  g04910(.A0(new_n5911_), .A1(new_n5903_), .B0(new_n5912_), .Y(new_n5913_));
  NOR2   g04911(.A(new_n5899_), .B(new_n5897_), .Y(new_n5914_));
  AOI21  g04912(.A0(new_n5901_), .A1(\A[69] ), .B0(new_n5914_), .Y(new_n5915_));
  XOR2   g04913(.A(new_n5915_), .B(new_n5913_), .Y(new_n5916_));
  XOR2   g04914(.A(new_n5916_), .B(new_n5910_), .Y(new_n5917_));
  XOR2   g04915(.A(new_n5909_), .B(new_n5902_), .Y(new_n5918_));
  NOR2   g04916(.A(new_n5899_), .B(\A[67] ), .Y(new_n5919_));
  OAI21  g04917(.A0(\A[68] ), .A1(new_n5897_), .B0(\A[69] ), .Y(new_n5920_));
  XOR2   g04918(.A(\A[68] ), .B(new_n5897_), .Y(new_n5921_));
  OAI22  g04919(.A0(new_n5921_), .A1(\A[69] ), .B0(new_n5920_), .B1(new_n5919_), .Y(new_n5922_));
  NOR2   g04920(.A(new_n5906_), .B(\A[70] ), .Y(new_n5923_));
  OAI21  g04921(.A0(\A[71] ), .A1(new_n5904_), .B0(\A[72] ), .Y(new_n5924_));
  OAI22  g04922(.A0(new_n5911_), .A1(\A[72] ), .B0(new_n5924_), .B1(new_n5923_), .Y(new_n5925_));
  NAND2  g04923(.A(new_n5925_), .B(new_n5922_), .Y(new_n5926_));
  NAND2  g04924(.A(\A[68] ), .B(\A[67] ), .Y(new_n5927_));
  OAI21  g04925(.A0(new_n5921_), .A1(new_n5896_), .B0(new_n5927_), .Y(new_n5928_));
  NAND2  g04926(.A(new_n5928_), .B(new_n5913_), .Y(new_n5929_));
  OAI21  g04927(.A0(new_n5916_), .A1(new_n5926_), .B0(new_n5929_), .Y(new_n5930_));
  AOI21  g04928(.A0(new_n5930_), .A1(new_n5918_), .B0(new_n5917_), .Y(new_n5931_));
  NAND2  g04929(.A(\A[77] ), .B(\A[76] ), .Y(new_n5932_));
  XOR2   g04930(.A(\A[77] ), .B(\A[76] ), .Y(new_n5933_));
  NAND2  g04931(.A(new_n5933_), .B(\A[78] ), .Y(new_n5934_));
  NAND2  g04932(.A(new_n5934_), .B(new_n5932_), .Y(new_n5935_));
  NAND2  g04933(.A(\A[74] ), .B(\A[73] ), .Y(new_n5936_));
  XOR2   g04934(.A(\A[74] ), .B(\A[73] ), .Y(new_n5937_));
  NAND2  g04935(.A(new_n5937_), .B(\A[75] ), .Y(new_n5938_));
  NAND2  g04936(.A(new_n5938_), .B(new_n5936_), .Y(new_n5939_));
  XOR2   g04937(.A(new_n5939_), .B(new_n5935_), .Y(new_n5940_));
  INV    g04938(.A(\A[75] ), .Y(new_n5941_));
  INV    g04939(.A(\A[73] ), .Y(new_n5942_));
  NAND2  g04940(.A(\A[74] ), .B(new_n5942_), .Y(new_n5943_));
  INV    g04941(.A(\A[74] ), .Y(new_n5944_));
  AOI21  g04942(.A0(new_n5944_), .A1(\A[73] ), .B0(new_n5941_), .Y(new_n5945_));
  AOI22  g04943(.A0(new_n5945_), .A1(new_n5943_), .B0(new_n5937_), .B1(new_n5941_), .Y(new_n5946_));
  INV    g04944(.A(\A[78] ), .Y(new_n5947_));
  INV    g04945(.A(\A[76] ), .Y(new_n5948_));
  NAND2  g04946(.A(\A[77] ), .B(new_n5948_), .Y(new_n5949_));
  INV    g04947(.A(\A[77] ), .Y(new_n5950_));
  AOI21  g04948(.A0(new_n5950_), .A1(\A[76] ), .B0(new_n5947_), .Y(new_n5951_));
  AOI22  g04949(.A0(new_n5951_), .A1(new_n5949_), .B0(new_n5933_), .B1(new_n5947_), .Y(new_n5952_));
  NOR2   g04950(.A(new_n5952_), .B(new_n5946_), .Y(new_n5953_));
  AOI22  g04951(.A0(new_n5938_), .A1(new_n5936_), .B0(new_n5934_), .B1(new_n5932_), .Y(new_n5954_));
  AOI21  g04952(.A0(new_n5953_), .A1(new_n5940_), .B0(new_n5954_), .Y(new_n5955_));
  XOR2   g04953(.A(new_n5953_), .B(new_n5940_), .Y(new_n5956_));
  NOR2   g04954(.A(new_n5944_), .B(\A[73] ), .Y(new_n5957_));
  OAI21  g04955(.A0(\A[74] ), .A1(new_n5942_), .B0(\A[75] ), .Y(new_n5958_));
  NAND2  g04956(.A(new_n5937_), .B(new_n5941_), .Y(new_n5959_));
  OAI21  g04957(.A0(new_n5958_), .A1(new_n5957_), .B0(new_n5959_), .Y(new_n5960_));
  XOR2   g04958(.A(new_n5952_), .B(new_n5960_), .Y(new_n5961_));
  NOR2   g04959(.A(new_n5950_), .B(\A[76] ), .Y(new_n5962_));
  OAI21  g04960(.A0(\A[77] ), .A1(new_n5948_), .B0(\A[78] ), .Y(new_n5963_));
  NAND2  g04961(.A(new_n5933_), .B(new_n5947_), .Y(new_n5964_));
  OAI21  g04962(.A0(new_n5963_), .A1(new_n5962_), .B0(new_n5964_), .Y(new_n5965_));
  NAND4  g04963(.A(new_n5965_), .B(new_n5960_), .C(new_n5939_), .D(new_n5935_), .Y(new_n5966_));
  NAND4  g04964(.A(new_n5928_), .B(new_n5913_), .C(new_n5925_), .D(new_n5922_), .Y(new_n5967_));
  XOR2   g04965(.A(new_n5952_), .B(new_n5946_), .Y(new_n5968_));
  NAND4  g04966(.A(new_n5968_), .B(new_n5967_), .C(new_n5966_), .D(new_n5918_), .Y(new_n5969_));
  OAI211 g04967(.A0(new_n5961_), .A1(new_n5955_), .B0(new_n5969_), .B1(new_n5956_), .Y(new_n5970_));
  NOR2   g04968(.A(new_n5944_), .B(new_n5942_), .Y(new_n5971_));
  AOI21  g04969(.A0(new_n5937_), .A1(\A[75] ), .B0(new_n5971_), .Y(new_n5972_));
  XOR2   g04970(.A(new_n5972_), .B(new_n5935_), .Y(new_n5973_));
  XOR2   g04971(.A(new_n5953_), .B(new_n5973_), .Y(new_n5974_));
  XOR2   g04972(.A(new_n5909_), .B(new_n5922_), .Y(new_n5975_));
  NOR2   g04973(.A(new_n5950_), .B(new_n5948_), .Y(new_n5976_));
  AOI21  g04974(.A0(new_n5933_), .A1(\A[78] ), .B0(new_n5976_), .Y(new_n5977_));
  NOR4   g04975(.A(new_n5952_), .B(new_n5946_), .C(new_n5972_), .D(new_n5977_), .Y(new_n5978_));
  NOR2   g04976(.A(new_n5906_), .B(new_n5904_), .Y(new_n5979_));
  AOI21  g04977(.A0(new_n5908_), .A1(\A[72] ), .B0(new_n5979_), .Y(new_n5980_));
  NOR4   g04978(.A(new_n5915_), .B(new_n5980_), .C(new_n5909_), .D(new_n5902_), .Y(new_n5981_));
  NOR4   g04979(.A(new_n5961_), .B(new_n5981_), .C(new_n5978_), .D(new_n5975_), .Y(new_n5982_));
  AOI221 g04980(.A0(new_n5937_), .A1(\A[75] ), .C0(new_n5971_), .B0(new_n5934_), .B1(new_n5932_), .Y(new_n5983_));
  AOI221 g04981(.A0(new_n5938_), .A1(new_n5936_), .C0(new_n5976_), .B0(new_n5933_), .B1(\A[78] ), .Y(new_n5984_));
  OAI211 g04982(.A0(new_n5984_), .A1(new_n5983_), .B0(new_n5965_), .B1(new_n5960_), .Y(new_n5985_));
  NAND2  g04983(.A(new_n5939_), .B(new_n5935_), .Y(new_n5986_));
  AOI21  g04984(.A0(new_n5986_), .A1(new_n5985_), .B0(new_n5961_), .Y(new_n5987_));
  OAI21  g04985(.A0(new_n5987_), .A1(new_n5974_), .B0(new_n5982_), .Y(new_n5988_));
  AOI21  g04986(.A0(new_n5988_), .A1(new_n5970_), .B0(new_n5931_), .Y(new_n5989_));
  XOR2   g04987(.A(new_n5916_), .B(new_n5926_), .Y(new_n5990_));
  XOR2   g04988(.A(new_n5915_), .B(new_n5980_), .Y(new_n5991_));
  NOR2   g04989(.A(new_n5915_), .B(new_n5980_), .Y(new_n5992_));
  AOI21  g04990(.A0(new_n5991_), .A1(new_n5910_), .B0(new_n5992_), .Y(new_n5993_));
  OAI21  g04991(.A0(new_n5993_), .A1(new_n5975_), .B0(new_n5990_), .Y(new_n5994_));
  OAI21  g04992(.A0(new_n5987_), .A1(new_n5974_), .B0(new_n5969_), .Y(new_n5995_));
  NOR2   g04993(.A(new_n5961_), .B(new_n5975_), .Y(new_n5996_));
  OAI211 g04994(.A0(new_n5965_), .A1(new_n5960_), .B0(new_n5939_), .B1(new_n5935_), .Y(new_n5997_));
  NAND4  g04995(.A(new_n5997_), .B(new_n5996_), .C(new_n5967_), .D(new_n5956_), .Y(new_n5998_));
  AOI21  g04996(.A0(new_n5998_), .A1(new_n5995_), .B0(new_n5994_), .Y(new_n5999_));
  NOR2   g04997(.A(new_n5961_), .B(new_n5978_), .Y(new_n6000_));
  XOR2   g04998(.A(new_n5909_), .B(new_n5902_), .Y(new_n6001_));
  XOR2   g04999(.A(new_n6001_), .B(new_n6000_), .Y(new_n6002_));
  NAND2  g05000(.A(new_n5871_), .B(new_n5861_), .Y(new_n6003_));
  XOR2   g05001(.A(new_n5825_), .B(new_n5806_), .Y(new_n6004_));
  XOR2   g05002(.A(new_n6004_), .B(new_n6003_), .Y(new_n6005_));
  NAND2  g05003(.A(new_n6005_), .B(new_n6002_), .Y(new_n6006_));
  NOR3   g05004(.A(new_n6006_), .B(new_n5999_), .C(new_n5989_), .Y(new_n6007_));
  OAI21  g05005(.A0(new_n5961_), .A1(new_n5955_), .B0(new_n5956_), .Y(new_n6008_));
  XOR2   g05006(.A(new_n6008_), .B(new_n5969_), .Y(new_n6009_));
  NAND2  g05007(.A(new_n6009_), .B(new_n5994_), .Y(new_n6010_));
  NAND2  g05008(.A(new_n5998_), .B(new_n5995_), .Y(new_n6011_));
  NAND2  g05009(.A(new_n6011_), .B(new_n5931_), .Y(new_n6012_));
  NAND2  g05010(.A(new_n5968_), .B(new_n5966_), .Y(new_n6013_));
  XOR2   g05011(.A(new_n6001_), .B(new_n6013_), .Y(new_n6014_));
  XOR2   g05012(.A(new_n5825_), .B(new_n5830_), .Y(new_n6015_));
  XOR2   g05013(.A(new_n6015_), .B(new_n6003_), .Y(new_n6016_));
  NOR2   g05014(.A(new_n6016_), .B(new_n6014_), .Y(new_n6017_));
  AOI21  g05015(.A0(new_n6012_), .A1(new_n6010_), .B0(new_n6017_), .Y(new_n6018_));
  OAI21  g05016(.A0(new_n6018_), .A1(new_n6007_), .B0(new_n5895_), .Y(new_n6019_));
  NAND2  g05017(.A(new_n5880_), .B(new_n5837_), .Y(new_n6020_));
  NAND2  g05018(.A(new_n5888_), .B(new_n5887_), .Y(new_n6021_));
  NAND3  g05019(.A(new_n5891_), .B(new_n5864_), .C(new_n5877_), .Y(new_n6022_));
  AOI211 g05020(.A0(new_n5877_), .A1(new_n6021_), .B(new_n6022_), .C(new_n5889_), .Y(new_n6023_));
  AOI21  g05021(.A0(new_n5879_), .A1(new_n5872_), .B0(new_n6023_), .Y(new_n6024_));
  OAI21  g05022(.A0(new_n6024_), .A1(new_n5837_), .B0(new_n6020_), .Y(new_n6025_));
  NAND2  g05023(.A(new_n5968_), .B(new_n5918_), .Y(new_n6026_));
  AOI211 g05024(.A0(new_n5952_), .A1(new_n5946_), .B(new_n5972_), .C(new_n5977_), .Y(new_n6027_));
  NOR4   g05025(.A(new_n6027_), .B(new_n6026_), .C(new_n5981_), .D(new_n5974_), .Y(new_n6028_));
  AOI21  g05026(.A0(new_n6008_), .A1(new_n5969_), .B0(new_n6028_), .Y(new_n6029_));
  OAI21  g05027(.A0(new_n6029_), .A1(new_n5994_), .B0(new_n6006_), .Y(new_n6030_));
  OAI21  g05028(.A0(new_n5999_), .A1(new_n5989_), .B0(new_n6017_), .Y(new_n6031_));
  OAI21  g05029(.A0(new_n6030_), .A1(new_n5989_), .B0(new_n6031_), .Y(new_n6032_));
  NAND2  g05030(.A(new_n6032_), .B(new_n6025_), .Y(new_n6033_));
  XOR2   g05031(.A(new_n6016_), .B(new_n6002_), .Y(new_n6034_));
  XOR2   g05032(.A(new_n5731_), .B(new_n5677_), .Y(new_n6035_));
  NOR2   g05033(.A(new_n6035_), .B(new_n6034_), .Y(new_n6036_));
  NAND3  g05034(.A(new_n6036_), .B(new_n6033_), .C(new_n6019_), .Y(new_n6037_));
  NAND3  g05035(.A(new_n6017_), .B(new_n6012_), .C(new_n6010_), .Y(new_n6038_));
  OAI21  g05036(.A0(new_n5999_), .A1(new_n5989_), .B0(new_n6006_), .Y(new_n6039_));
  AOI21  g05037(.A0(new_n6039_), .A1(new_n6038_), .B0(new_n6025_), .Y(new_n6040_));
  NAND3  g05038(.A(new_n6006_), .B(new_n6012_), .C(new_n6010_), .Y(new_n6041_));
  AOI21  g05039(.A0(new_n6031_), .A1(new_n6041_), .B0(new_n5895_), .Y(new_n6042_));
  INV    g05040(.A(new_n6036_), .Y(new_n6043_));
  OAI21  g05041(.A0(new_n6042_), .A1(new_n6040_), .B0(new_n6043_), .Y(new_n6044_));
  AOI21  g05042(.A0(new_n6044_), .A1(new_n6037_), .B0(new_n5800_), .Y(new_n6045_));
  NAND3  g05043(.A(new_n5732_), .B(new_n5723_), .C(new_n5721_), .Y(new_n6046_));
  OAI21  g05044(.A0(new_n5674_), .A1(new_n5664_), .B0(new_n5717_), .Y(new_n6047_));
  AOI21  g05045(.A0(new_n6047_), .A1(new_n6046_), .B0(new_n5796_), .Y(new_n6048_));
  NAND3  g05046(.A(new_n5717_), .B(new_n5723_), .C(new_n5721_), .Y(new_n6049_));
  OAI21  g05047(.A0(new_n5674_), .A1(new_n5664_), .B0(new_n5732_), .Y(new_n6050_));
  AOI21  g05048(.A0(new_n6050_), .A1(new_n6049_), .B0(new_n5792_), .Y(new_n6051_));
  NOR2   g05049(.A(new_n6051_), .B(new_n6048_), .Y(new_n6052_));
  AOI21  g05050(.A0(new_n6032_), .A1(new_n6025_), .B0(new_n6036_), .Y(new_n6053_));
  NAND2  g05051(.A(new_n6053_), .B(new_n6019_), .Y(new_n6054_));
  OAI21  g05052(.A0(new_n6042_), .A1(new_n6040_), .B0(new_n6036_), .Y(new_n6055_));
  AOI21  g05053(.A0(new_n6055_), .A1(new_n6054_), .B0(new_n6052_), .Y(new_n6056_));
  XOR2   g05054(.A(new_n6035_), .B(new_n6034_), .Y(new_n6057_));
  INV    g05055(.A(new_n6057_), .Y(new_n6058_));
  XOR2   g05056(.A(new_n5419_), .B(new_n5417_), .Y(new_n6059_));
  AOI21  g05057(.A0(new_n5419_), .A1(new_n5405_), .B0(new_n5500_), .Y(new_n6060_));
  AOI22  g05058(.A0(new_n6060_), .A1(new_n5441_), .B0(new_n5500_), .B1(new_n6059_), .Y(new_n6061_));
  NOR2   g05059(.A(new_n6061_), .B(new_n6058_), .Y(new_n6062_));
  INV    g05060(.A(new_n6062_), .Y(new_n6063_));
  NOR3   g05061(.A(new_n6063_), .B(new_n6056_), .C(new_n6045_), .Y(new_n6064_));
  NOR3   g05062(.A(new_n6043_), .B(new_n6042_), .C(new_n6040_), .Y(new_n6065_));
  AOI21  g05063(.A0(new_n6033_), .A1(new_n6019_), .B0(new_n6036_), .Y(new_n6066_));
  OAI21  g05064(.A0(new_n6066_), .A1(new_n6065_), .B0(new_n6052_), .Y(new_n6067_));
  NOR3   g05065(.A(new_n6036_), .B(new_n6042_), .C(new_n6040_), .Y(new_n6068_));
  AOI21  g05066(.A0(new_n6033_), .A1(new_n6019_), .B0(new_n6043_), .Y(new_n6069_));
  OAI21  g05067(.A0(new_n6069_), .A1(new_n6068_), .B0(new_n5800_), .Y(new_n6070_));
  AOI21  g05068(.A0(new_n6070_), .A1(new_n6067_), .B0(new_n6062_), .Y(new_n6071_));
  OAI21  g05069(.A0(new_n6071_), .A1(new_n6064_), .B0(new_n5570_), .Y(new_n6072_));
  NOR3   g05070(.A(new_n5508_), .B(new_n5507_), .C(new_n5505_), .Y(new_n6073_));
  AOI21  g05071(.A0(new_n5439_), .A1(new_n5422_), .B0(new_n5501_), .Y(new_n6074_));
  OAI21  g05072(.A0(new_n6074_), .A1(new_n6073_), .B0(new_n5565_), .Y(new_n6075_));
  NOR3   g05073(.A(new_n5501_), .B(new_n5507_), .C(new_n5505_), .Y(new_n6076_));
  AOI21  g05074(.A0(new_n5439_), .A1(new_n5422_), .B0(new_n5508_), .Y(new_n6077_));
  OAI21  g05075(.A0(new_n6077_), .A1(new_n6076_), .B0(new_n5559_), .Y(new_n6078_));
  NAND2  g05076(.A(new_n6078_), .B(new_n6075_), .Y(new_n6079_));
  NOR3   g05077(.A(new_n6062_), .B(new_n6056_), .C(new_n6045_), .Y(new_n6080_));
  AOI21  g05078(.A0(new_n6070_), .A1(new_n6067_), .B0(new_n6063_), .Y(new_n6081_));
  OAI21  g05079(.A0(new_n6081_), .A1(new_n6080_), .B0(new_n6079_), .Y(new_n6082_));
  XOR2   g05080(.A(new_n6061_), .B(new_n6057_), .Y(new_n6083_));
  INV    g05081(.A(new_n4974_), .Y(new_n6084_));
  XOR2   g05082(.A(new_n5058_), .B(new_n6084_), .Y(new_n6085_));
  NOR2   g05083(.A(new_n6085_), .B(new_n6083_), .Y(new_n6086_));
  NAND3  g05084(.A(new_n6086_), .B(new_n6082_), .C(new_n6072_), .Y(new_n6087_));
  NAND3  g05085(.A(new_n6062_), .B(new_n6070_), .C(new_n6067_), .Y(new_n6088_));
  OAI21  g05086(.A0(new_n6056_), .A1(new_n6045_), .B0(new_n6063_), .Y(new_n6089_));
  AOI21  g05087(.A0(new_n6089_), .A1(new_n6088_), .B0(new_n6079_), .Y(new_n6090_));
  NAND3  g05088(.A(new_n6063_), .B(new_n6070_), .C(new_n6067_), .Y(new_n6091_));
  OAI21  g05089(.A0(new_n6056_), .A1(new_n6045_), .B0(new_n6062_), .Y(new_n6092_));
  AOI21  g05090(.A0(new_n6092_), .A1(new_n6091_), .B0(new_n5570_), .Y(new_n6093_));
  INV    g05091(.A(new_n6086_), .Y(new_n6094_));
  OAI21  g05092(.A0(new_n6093_), .A1(new_n6090_), .B0(new_n6094_), .Y(new_n6095_));
  AOI21  g05093(.A0(new_n6095_), .A1(new_n6087_), .B0(new_n5203_), .Y(new_n6096_));
  NAND2  g05094(.A(new_n4972_), .B(new_n4958_), .Y(new_n6097_));
  NAND2  g05095(.A(new_n6097_), .B(new_n5065_), .Y(new_n6098_));
  NAND3  g05096(.A(new_n5200_), .B(new_n5062_), .C(new_n6098_), .Y(new_n6099_));
  OAI21  g05097(.A0(new_n5068_), .A1(new_n4973_), .B0(new_n5059_), .Y(new_n6100_));
  AOI21  g05098(.A0(new_n6100_), .A1(new_n6099_), .B0(new_n5195_), .Y(new_n6101_));
  AOI21  g05099(.A0(new_n5195_), .A1(new_n5070_), .B0(new_n6101_), .Y(new_n6102_));
  NAND3  g05100(.A(new_n6094_), .B(new_n6082_), .C(new_n6072_), .Y(new_n6103_));
  OAI21  g05101(.A0(new_n6093_), .A1(new_n6090_), .B0(new_n6086_), .Y(new_n6104_));
  AOI21  g05102(.A0(new_n6104_), .A1(new_n6103_), .B0(new_n6102_), .Y(new_n6105_));
  AOI221 g05103(.A0(new_n6060_), .A1(new_n5441_), .C0(new_n6058_), .B0(new_n5500_), .B1(new_n6059_), .Y(new_n6106_));
  NOR2   g05104(.A(new_n6061_), .B(new_n6057_), .Y(new_n6107_));
  OAI21  g05105(.A0(new_n6107_), .A1(new_n6106_), .B0(new_n6085_), .Y(new_n6108_));
  NOR3   g05106(.A(new_n6085_), .B(new_n6107_), .C(new_n6106_), .Y(new_n6109_));
  INV    g05107(.A(new_n6109_), .Y(new_n6110_));
  INV    g05108(.A(\A[939] ), .Y(new_n6111_));
  INV    g05109(.A(\A[938] ), .Y(new_n6112_));
  NAND2  g05110(.A(new_n6112_), .B(\A[937] ), .Y(new_n6113_));
  INV    g05111(.A(\A[937] ), .Y(new_n6114_));
  AOI21  g05112(.A0(\A[938] ), .A1(new_n6114_), .B0(new_n6111_), .Y(new_n6115_));
  XOR2   g05113(.A(\A[938] ), .B(\A[937] ), .Y(new_n6116_));
  AOI22  g05114(.A0(new_n6116_), .A1(new_n6111_), .B0(new_n6115_), .B1(new_n6113_), .Y(new_n6117_));
  INV    g05115(.A(\A[942] ), .Y(new_n6118_));
  INV    g05116(.A(\A[941] ), .Y(new_n6119_));
  NAND2  g05117(.A(new_n6119_), .B(\A[940] ), .Y(new_n6120_));
  INV    g05118(.A(\A[940] ), .Y(new_n6121_));
  AOI21  g05119(.A0(\A[941] ), .A1(new_n6121_), .B0(new_n6118_), .Y(new_n6122_));
  XOR2   g05120(.A(\A[941] ), .B(\A[940] ), .Y(new_n6123_));
  AOI22  g05121(.A0(new_n6123_), .A1(new_n6118_), .B0(new_n6122_), .B1(new_n6120_), .Y(new_n6124_));
  NOR2   g05122(.A(new_n6119_), .B(new_n6121_), .Y(new_n6125_));
  AOI21  g05123(.A0(new_n6123_), .A1(\A[942] ), .B0(new_n6125_), .Y(new_n6126_));
  NOR2   g05124(.A(new_n6112_), .B(new_n6114_), .Y(new_n6127_));
  AOI21  g05125(.A0(new_n6116_), .A1(\A[939] ), .B0(new_n6127_), .Y(new_n6128_));
  XOR2   g05126(.A(new_n6124_), .B(new_n6117_), .Y(new_n6129_));
  INV    g05127(.A(\A[933] ), .Y(new_n6130_));
  INV    g05128(.A(\A[932] ), .Y(new_n6131_));
  NAND2  g05129(.A(new_n6131_), .B(\A[931] ), .Y(new_n6132_));
  INV    g05130(.A(\A[931] ), .Y(new_n6133_));
  AOI21  g05131(.A0(\A[932] ), .A1(new_n6133_), .B0(new_n6130_), .Y(new_n6134_));
  XOR2   g05132(.A(\A[932] ), .B(\A[931] ), .Y(new_n6135_));
  AOI22  g05133(.A0(new_n6135_), .A1(new_n6130_), .B0(new_n6134_), .B1(new_n6132_), .Y(new_n6136_));
  INV    g05134(.A(\A[936] ), .Y(new_n6137_));
  INV    g05135(.A(\A[935] ), .Y(new_n6138_));
  NAND2  g05136(.A(new_n6138_), .B(\A[934] ), .Y(new_n6139_));
  INV    g05137(.A(\A[934] ), .Y(new_n6140_));
  AOI21  g05138(.A0(\A[935] ), .A1(new_n6140_), .B0(new_n6137_), .Y(new_n6141_));
  XOR2   g05139(.A(\A[935] ), .B(\A[934] ), .Y(new_n6142_));
  AOI22  g05140(.A0(new_n6142_), .A1(new_n6137_), .B0(new_n6141_), .B1(new_n6139_), .Y(new_n6143_));
  NAND2  g05141(.A(\A[935] ), .B(\A[934] ), .Y(new_n6144_));
  INV    g05142(.A(new_n6144_), .Y(new_n6145_));
  AOI21  g05143(.A0(new_n6142_), .A1(\A[936] ), .B0(new_n6145_), .Y(new_n6146_));
  NOR2   g05144(.A(new_n6131_), .B(new_n6133_), .Y(new_n6147_));
  AOI21  g05145(.A0(new_n6135_), .A1(\A[933] ), .B0(new_n6147_), .Y(new_n6148_));
  XOR2   g05146(.A(new_n6143_), .B(new_n6136_), .Y(new_n6149_));
  XOR2   g05147(.A(new_n6149_), .B(new_n6129_), .Y(new_n6150_));
  INV    g05148(.A(\A[927] ), .Y(new_n6151_));
  INV    g05149(.A(\A[926] ), .Y(new_n6152_));
  NAND2  g05150(.A(new_n6152_), .B(\A[925] ), .Y(new_n6153_));
  INV    g05151(.A(\A[925] ), .Y(new_n6154_));
  AOI21  g05152(.A0(\A[926] ), .A1(new_n6154_), .B0(new_n6151_), .Y(new_n6155_));
  XOR2   g05153(.A(\A[926] ), .B(\A[925] ), .Y(new_n6156_));
  AOI22  g05154(.A0(new_n6156_), .A1(new_n6151_), .B0(new_n6155_), .B1(new_n6153_), .Y(new_n6157_));
  INV    g05155(.A(\A[930] ), .Y(new_n6158_));
  INV    g05156(.A(\A[929] ), .Y(new_n6159_));
  NAND2  g05157(.A(new_n6159_), .B(\A[928] ), .Y(new_n6160_));
  INV    g05158(.A(\A[928] ), .Y(new_n6161_));
  AOI21  g05159(.A0(\A[929] ), .A1(new_n6161_), .B0(new_n6158_), .Y(new_n6162_));
  XOR2   g05160(.A(\A[929] ), .B(\A[928] ), .Y(new_n6163_));
  AOI22  g05161(.A0(new_n6163_), .A1(new_n6158_), .B0(new_n6162_), .B1(new_n6160_), .Y(new_n6164_));
  NOR2   g05162(.A(new_n6159_), .B(new_n6161_), .Y(new_n6165_));
  AOI21  g05163(.A0(new_n6163_), .A1(\A[930] ), .B0(new_n6165_), .Y(new_n6166_));
  NOR2   g05164(.A(new_n6152_), .B(new_n6154_), .Y(new_n6167_));
  AOI21  g05165(.A0(new_n6156_), .A1(\A[927] ), .B0(new_n6167_), .Y(new_n6168_));
  XOR2   g05166(.A(new_n6164_), .B(new_n6157_), .Y(new_n6169_));
  INV    g05167(.A(\A[921] ), .Y(new_n6170_));
  INV    g05168(.A(\A[920] ), .Y(new_n6171_));
  NAND2  g05169(.A(new_n6171_), .B(\A[919] ), .Y(new_n6172_));
  INV    g05170(.A(\A[919] ), .Y(new_n6173_));
  AOI21  g05171(.A0(\A[920] ), .A1(new_n6173_), .B0(new_n6170_), .Y(new_n6174_));
  XOR2   g05172(.A(\A[920] ), .B(\A[919] ), .Y(new_n6175_));
  AOI22  g05173(.A0(new_n6175_), .A1(new_n6170_), .B0(new_n6174_), .B1(new_n6172_), .Y(new_n6176_));
  INV    g05174(.A(\A[924] ), .Y(new_n6177_));
  INV    g05175(.A(\A[923] ), .Y(new_n6178_));
  NAND2  g05176(.A(new_n6178_), .B(\A[922] ), .Y(new_n6179_));
  INV    g05177(.A(\A[922] ), .Y(new_n6180_));
  AOI21  g05178(.A0(\A[923] ), .A1(new_n6180_), .B0(new_n6177_), .Y(new_n6181_));
  XOR2   g05179(.A(\A[923] ), .B(\A[922] ), .Y(new_n6182_));
  AOI22  g05180(.A0(new_n6182_), .A1(new_n6177_), .B0(new_n6181_), .B1(new_n6179_), .Y(new_n6183_));
  NOR2   g05181(.A(new_n6178_), .B(new_n6180_), .Y(new_n6184_));
  AOI21  g05182(.A0(new_n6182_), .A1(\A[924] ), .B0(new_n6184_), .Y(new_n6185_));
  NOR2   g05183(.A(new_n6171_), .B(new_n6173_), .Y(new_n6186_));
  AOI21  g05184(.A0(new_n6175_), .A1(\A[921] ), .B0(new_n6186_), .Y(new_n6187_));
  XOR2   g05185(.A(new_n6183_), .B(new_n6176_), .Y(new_n6188_));
  XOR2   g05186(.A(new_n6188_), .B(new_n6169_), .Y(new_n6189_));
  INV    g05187(.A(new_n6189_), .Y(new_n6190_));
  XOR2   g05188(.A(new_n6190_), .B(new_n6150_), .Y(new_n6191_));
  INV    g05189(.A(new_n6191_), .Y(new_n6192_));
  INV    g05190(.A(\A[915] ), .Y(new_n6193_));
  INV    g05191(.A(\A[914] ), .Y(new_n6194_));
  NAND2  g05192(.A(new_n6194_), .B(\A[913] ), .Y(new_n6195_));
  INV    g05193(.A(\A[913] ), .Y(new_n6196_));
  AOI21  g05194(.A0(\A[914] ), .A1(new_n6196_), .B0(new_n6193_), .Y(new_n6197_));
  XOR2   g05195(.A(\A[914] ), .B(\A[913] ), .Y(new_n6198_));
  AOI22  g05196(.A0(new_n6198_), .A1(new_n6193_), .B0(new_n6197_), .B1(new_n6195_), .Y(new_n6199_));
  INV    g05197(.A(\A[918] ), .Y(new_n6200_));
  INV    g05198(.A(\A[917] ), .Y(new_n6201_));
  NAND2  g05199(.A(new_n6201_), .B(\A[916] ), .Y(new_n6202_));
  INV    g05200(.A(\A[916] ), .Y(new_n6203_));
  AOI21  g05201(.A0(\A[917] ), .A1(new_n6203_), .B0(new_n6200_), .Y(new_n6204_));
  XOR2   g05202(.A(\A[917] ), .B(\A[916] ), .Y(new_n6205_));
  AOI22  g05203(.A0(new_n6205_), .A1(new_n6200_), .B0(new_n6204_), .B1(new_n6202_), .Y(new_n6206_));
  NOR2   g05204(.A(new_n6201_), .B(new_n6203_), .Y(new_n6207_));
  AOI21  g05205(.A0(new_n6205_), .A1(\A[918] ), .B0(new_n6207_), .Y(new_n6208_));
  NOR2   g05206(.A(new_n6194_), .B(new_n6196_), .Y(new_n6209_));
  AOI21  g05207(.A0(new_n6198_), .A1(\A[915] ), .B0(new_n6209_), .Y(new_n6210_));
  XOR2   g05208(.A(new_n6206_), .B(new_n6199_), .Y(new_n6211_));
  INV    g05209(.A(\A[909] ), .Y(new_n6212_));
  INV    g05210(.A(\A[908] ), .Y(new_n6213_));
  NAND2  g05211(.A(new_n6213_), .B(\A[907] ), .Y(new_n6214_));
  INV    g05212(.A(\A[907] ), .Y(new_n6215_));
  AOI21  g05213(.A0(\A[908] ), .A1(new_n6215_), .B0(new_n6212_), .Y(new_n6216_));
  XOR2   g05214(.A(\A[908] ), .B(\A[907] ), .Y(new_n6217_));
  AOI22  g05215(.A0(new_n6217_), .A1(new_n6212_), .B0(new_n6216_), .B1(new_n6214_), .Y(new_n6218_));
  INV    g05216(.A(\A[912] ), .Y(new_n6219_));
  INV    g05217(.A(\A[911] ), .Y(new_n6220_));
  NAND2  g05218(.A(new_n6220_), .B(\A[910] ), .Y(new_n6221_));
  INV    g05219(.A(\A[910] ), .Y(new_n6222_));
  AOI21  g05220(.A0(\A[911] ), .A1(new_n6222_), .B0(new_n6219_), .Y(new_n6223_));
  XOR2   g05221(.A(\A[911] ), .B(\A[910] ), .Y(new_n6224_));
  AOI22  g05222(.A0(new_n6224_), .A1(new_n6219_), .B0(new_n6223_), .B1(new_n6221_), .Y(new_n6225_));
  NOR2   g05223(.A(new_n6220_), .B(new_n6222_), .Y(new_n6226_));
  AOI21  g05224(.A0(new_n6224_), .A1(\A[912] ), .B0(new_n6226_), .Y(new_n6227_));
  NOR2   g05225(.A(new_n6213_), .B(new_n6215_), .Y(new_n6228_));
  AOI21  g05226(.A0(new_n6217_), .A1(\A[909] ), .B0(new_n6228_), .Y(new_n6229_));
  XOR2   g05227(.A(new_n6225_), .B(new_n6218_), .Y(new_n6230_));
  XOR2   g05228(.A(new_n6230_), .B(new_n6211_), .Y(new_n6231_));
  INV    g05229(.A(\A[903] ), .Y(new_n6232_));
  INV    g05230(.A(\A[902] ), .Y(new_n6233_));
  NAND2  g05231(.A(new_n6233_), .B(\A[901] ), .Y(new_n6234_));
  INV    g05232(.A(\A[901] ), .Y(new_n6235_));
  AOI21  g05233(.A0(\A[902] ), .A1(new_n6235_), .B0(new_n6232_), .Y(new_n6236_));
  XOR2   g05234(.A(\A[902] ), .B(\A[901] ), .Y(new_n6237_));
  AOI22  g05235(.A0(new_n6237_), .A1(new_n6232_), .B0(new_n6236_), .B1(new_n6234_), .Y(new_n6238_));
  INV    g05236(.A(\A[906] ), .Y(new_n6239_));
  INV    g05237(.A(\A[905] ), .Y(new_n6240_));
  NAND2  g05238(.A(new_n6240_), .B(\A[904] ), .Y(new_n6241_));
  INV    g05239(.A(\A[904] ), .Y(new_n6242_));
  AOI21  g05240(.A0(\A[905] ), .A1(new_n6242_), .B0(new_n6239_), .Y(new_n6243_));
  XOR2   g05241(.A(\A[905] ), .B(\A[904] ), .Y(new_n6244_));
  AOI22  g05242(.A0(new_n6244_), .A1(new_n6239_), .B0(new_n6243_), .B1(new_n6241_), .Y(new_n6245_));
  NOR2   g05243(.A(new_n6240_), .B(new_n6242_), .Y(new_n6246_));
  AOI21  g05244(.A0(new_n6244_), .A1(\A[906] ), .B0(new_n6246_), .Y(new_n6247_));
  NOR2   g05245(.A(new_n6233_), .B(new_n6235_), .Y(new_n6248_));
  AOI21  g05246(.A0(new_n6237_), .A1(\A[903] ), .B0(new_n6248_), .Y(new_n6249_));
  XOR2   g05247(.A(new_n6245_), .B(new_n6238_), .Y(new_n6250_));
  INV    g05248(.A(\A[897] ), .Y(new_n6251_));
  INV    g05249(.A(\A[896] ), .Y(new_n6252_));
  NAND2  g05250(.A(new_n6252_), .B(\A[895] ), .Y(new_n6253_));
  INV    g05251(.A(\A[895] ), .Y(new_n6254_));
  AOI21  g05252(.A0(\A[896] ), .A1(new_n6254_), .B0(new_n6251_), .Y(new_n6255_));
  XOR2   g05253(.A(\A[896] ), .B(\A[895] ), .Y(new_n6256_));
  AOI22  g05254(.A0(new_n6256_), .A1(new_n6251_), .B0(new_n6255_), .B1(new_n6253_), .Y(new_n6257_));
  INV    g05255(.A(\A[900] ), .Y(new_n6258_));
  INV    g05256(.A(\A[899] ), .Y(new_n6259_));
  NAND2  g05257(.A(new_n6259_), .B(\A[898] ), .Y(new_n6260_));
  INV    g05258(.A(\A[898] ), .Y(new_n6261_));
  AOI21  g05259(.A0(\A[899] ), .A1(new_n6261_), .B0(new_n6258_), .Y(new_n6262_));
  XOR2   g05260(.A(\A[899] ), .B(\A[898] ), .Y(new_n6263_));
  AOI22  g05261(.A0(new_n6263_), .A1(new_n6258_), .B0(new_n6262_), .B1(new_n6260_), .Y(new_n6264_));
  NOR2   g05262(.A(new_n6259_), .B(new_n6261_), .Y(new_n6265_));
  AOI21  g05263(.A0(new_n6263_), .A1(\A[900] ), .B0(new_n6265_), .Y(new_n6266_));
  NOR2   g05264(.A(new_n6252_), .B(new_n6254_), .Y(new_n6267_));
  AOI21  g05265(.A0(new_n6256_), .A1(\A[897] ), .B0(new_n6267_), .Y(new_n6268_));
  XOR2   g05266(.A(new_n6264_), .B(new_n6257_), .Y(new_n6269_));
  XOR2   g05267(.A(new_n6269_), .B(new_n6250_), .Y(new_n6270_));
  INV    g05268(.A(new_n6270_), .Y(new_n6271_));
  XOR2   g05269(.A(new_n6271_), .B(new_n6231_), .Y(new_n6272_));
  XOR2   g05270(.A(new_n6272_), .B(new_n6192_), .Y(new_n6273_));
  INV    g05271(.A(new_n6273_), .Y(new_n6274_));
  INV    g05272(.A(\A[891] ), .Y(new_n6275_));
  INV    g05273(.A(\A[890] ), .Y(new_n6276_));
  NAND2  g05274(.A(new_n6276_), .B(\A[889] ), .Y(new_n6277_));
  INV    g05275(.A(\A[889] ), .Y(new_n6278_));
  AOI21  g05276(.A0(\A[890] ), .A1(new_n6278_), .B0(new_n6275_), .Y(new_n6279_));
  XOR2   g05277(.A(\A[890] ), .B(\A[889] ), .Y(new_n6280_));
  AOI22  g05278(.A0(new_n6280_), .A1(new_n6275_), .B0(new_n6279_), .B1(new_n6277_), .Y(new_n6281_));
  INV    g05279(.A(\A[894] ), .Y(new_n6282_));
  INV    g05280(.A(\A[893] ), .Y(new_n6283_));
  NAND2  g05281(.A(new_n6283_), .B(\A[892] ), .Y(new_n6284_));
  INV    g05282(.A(\A[892] ), .Y(new_n6285_));
  AOI21  g05283(.A0(\A[893] ), .A1(new_n6285_), .B0(new_n6282_), .Y(new_n6286_));
  XOR2   g05284(.A(\A[893] ), .B(\A[892] ), .Y(new_n6287_));
  AOI22  g05285(.A0(new_n6287_), .A1(new_n6282_), .B0(new_n6286_), .B1(new_n6284_), .Y(new_n6288_));
  NOR2   g05286(.A(new_n6283_), .B(new_n6285_), .Y(new_n6289_));
  AOI21  g05287(.A0(new_n6287_), .A1(\A[894] ), .B0(new_n6289_), .Y(new_n6290_));
  NOR2   g05288(.A(new_n6276_), .B(new_n6278_), .Y(new_n6291_));
  AOI21  g05289(.A0(new_n6280_), .A1(\A[891] ), .B0(new_n6291_), .Y(new_n6292_));
  XOR2   g05290(.A(new_n6288_), .B(new_n6281_), .Y(new_n6293_));
  INV    g05291(.A(\A[885] ), .Y(new_n6294_));
  INV    g05292(.A(\A[884] ), .Y(new_n6295_));
  NAND2  g05293(.A(new_n6295_), .B(\A[883] ), .Y(new_n6296_));
  INV    g05294(.A(\A[883] ), .Y(new_n6297_));
  AOI21  g05295(.A0(\A[884] ), .A1(new_n6297_), .B0(new_n6294_), .Y(new_n6298_));
  XOR2   g05296(.A(\A[884] ), .B(\A[883] ), .Y(new_n6299_));
  AOI22  g05297(.A0(new_n6299_), .A1(new_n6294_), .B0(new_n6298_), .B1(new_n6296_), .Y(new_n6300_));
  INV    g05298(.A(\A[888] ), .Y(new_n6301_));
  INV    g05299(.A(\A[887] ), .Y(new_n6302_));
  NAND2  g05300(.A(new_n6302_), .B(\A[886] ), .Y(new_n6303_));
  INV    g05301(.A(\A[886] ), .Y(new_n6304_));
  AOI21  g05302(.A0(\A[887] ), .A1(new_n6304_), .B0(new_n6301_), .Y(new_n6305_));
  XOR2   g05303(.A(\A[887] ), .B(\A[886] ), .Y(new_n6306_));
  AOI22  g05304(.A0(new_n6306_), .A1(new_n6301_), .B0(new_n6305_), .B1(new_n6303_), .Y(new_n6307_));
  NOR2   g05305(.A(new_n6302_), .B(new_n6304_), .Y(new_n6308_));
  AOI21  g05306(.A0(new_n6306_), .A1(\A[888] ), .B0(new_n6308_), .Y(new_n6309_));
  NOR2   g05307(.A(new_n6295_), .B(new_n6297_), .Y(new_n6310_));
  AOI21  g05308(.A0(new_n6299_), .A1(\A[885] ), .B0(new_n6310_), .Y(new_n6311_));
  XOR2   g05309(.A(new_n6307_), .B(new_n6300_), .Y(new_n6312_));
  XOR2   g05310(.A(new_n6312_), .B(new_n6293_), .Y(new_n6313_));
  INV    g05311(.A(\A[879] ), .Y(new_n6314_));
  INV    g05312(.A(\A[878] ), .Y(new_n6315_));
  NAND2  g05313(.A(new_n6315_), .B(\A[877] ), .Y(new_n6316_));
  INV    g05314(.A(\A[877] ), .Y(new_n6317_));
  AOI21  g05315(.A0(\A[878] ), .A1(new_n6317_), .B0(new_n6314_), .Y(new_n6318_));
  XOR2   g05316(.A(\A[878] ), .B(\A[877] ), .Y(new_n6319_));
  AOI22  g05317(.A0(new_n6319_), .A1(new_n6314_), .B0(new_n6318_), .B1(new_n6316_), .Y(new_n6320_));
  INV    g05318(.A(\A[882] ), .Y(new_n6321_));
  INV    g05319(.A(\A[881] ), .Y(new_n6322_));
  NAND2  g05320(.A(new_n6322_), .B(\A[880] ), .Y(new_n6323_));
  INV    g05321(.A(\A[880] ), .Y(new_n6324_));
  AOI21  g05322(.A0(\A[881] ), .A1(new_n6324_), .B0(new_n6321_), .Y(new_n6325_));
  XOR2   g05323(.A(\A[881] ), .B(\A[880] ), .Y(new_n6326_));
  AOI22  g05324(.A0(new_n6326_), .A1(new_n6321_), .B0(new_n6325_), .B1(new_n6323_), .Y(new_n6327_));
  NOR2   g05325(.A(new_n6322_), .B(new_n6324_), .Y(new_n6328_));
  AOI21  g05326(.A0(new_n6326_), .A1(\A[882] ), .B0(new_n6328_), .Y(new_n6329_));
  NOR2   g05327(.A(new_n6315_), .B(new_n6317_), .Y(new_n6330_));
  AOI21  g05328(.A0(new_n6319_), .A1(\A[879] ), .B0(new_n6330_), .Y(new_n6331_));
  XOR2   g05329(.A(new_n6327_), .B(new_n6320_), .Y(new_n6332_));
  INV    g05330(.A(\A[873] ), .Y(new_n6333_));
  INV    g05331(.A(\A[872] ), .Y(new_n6334_));
  NAND2  g05332(.A(new_n6334_), .B(\A[871] ), .Y(new_n6335_));
  INV    g05333(.A(\A[871] ), .Y(new_n6336_));
  AOI21  g05334(.A0(\A[872] ), .A1(new_n6336_), .B0(new_n6333_), .Y(new_n6337_));
  XOR2   g05335(.A(\A[872] ), .B(\A[871] ), .Y(new_n6338_));
  AOI22  g05336(.A0(new_n6338_), .A1(new_n6333_), .B0(new_n6337_), .B1(new_n6335_), .Y(new_n6339_));
  INV    g05337(.A(\A[876] ), .Y(new_n6340_));
  INV    g05338(.A(\A[875] ), .Y(new_n6341_));
  NAND2  g05339(.A(new_n6341_), .B(\A[874] ), .Y(new_n6342_));
  INV    g05340(.A(\A[874] ), .Y(new_n6343_));
  AOI21  g05341(.A0(\A[875] ), .A1(new_n6343_), .B0(new_n6340_), .Y(new_n6344_));
  XOR2   g05342(.A(\A[875] ), .B(\A[874] ), .Y(new_n6345_));
  AOI22  g05343(.A0(new_n6345_), .A1(new_n6340_), .B0(new_n6344_), .B1(new_n6342_), .Y(new_n6346_));
  NOR2   g05344(.A(new_n6341_), .B(new_n6343_), .Y(new_n6347_));
  AOI21  g05345(.A0(new_n6345_), .A1(\A[876] ), .B0(new_n6347_), .Y(new_n6348_));
  NOR2   g05346(.A(new_n6334_), .B(new_n6336_), .Y(new_n6349_));
  AOI21  g05347(.A0(new_n6338_), .A1(\A[873] ), .B0(new_n6349_), .Y(new_n6350_));
  XOR2   g05348(.A(new_n6346_), .B(new_n6339_), .Y(new_n6351_));
  XOR2   g05349(.A(new_n6351_), .B(new_n6332_), .Y(new_n6352_));
  INV    g05350(.A(new_n6352_), .Y(new_n6353_));
  XOR2   g05351(.A(new_n6353_), .B(new_n6313_), .Y(new_n6354_));
  INV    g05352(.A(new_n6354_), .Y(new_n6355_));
  INV    g05353(.A(\A[867] ), .Y(new_n6356_));
  INV    g05354(.A(\A[866] ), .Y(new_n6357_));
  NAND2  g05355(.A(new_n6357_), .B(\A[865] ), .Y(new_n6358_));
  INV    g05356(.A(\A[865] ), .Y(new_n6359_));
  AOI21  g05357(.A0(\A[866] ), .A1(new_n6359_), .B0(new_n6356_), .Y(new_n6360_));
  XOR2   g05358(.A(\A[866] ), .B(\A[865] ), .Y(new_n6361_));
  AOI22  g05359(.A0(new_n6361_), .A1(new_n6356_), .B0(new_n6360_), .B1(new_n6358_), .Y(new_n6362_));
  INV    g05360(.A(\A[870] ), .Y(new_n6363_));
  INV    g05361(.A(\A[869] ), .Y(new_n6364_));
  NAND2  g05362(.A(new_n6364_), .B(\A[868] ), .Y(new_n6365_));
  INV    g05363(.A(\A[868] ), .Y(new_n6366_));
  AOI21  g05364(.A0(\A[869] ), .A1(new_n6366_), .B0(new_n6363_), .Y(new_n6367_));
  XOR2   g05365(.A(\A[869] ), .B(\A[868] ), .Y(new_n6368_));
  AOI22  g05366(.A0(new_n6368_), .A1(new_n6363_), .B0(new_n6367_), .B1(new_n6365_), .Y(new_n6369_));
  NOR2   g05367(.A(new_n6364_), .B(new_n6366_), .Y(new_n6370_));
  AOI21  g05368(.A0(new_n6368_), .A1(\A[870] ), .B0(new_n6370_), .Y(new_n6371_));
  NOR2   g05369(.A(new_n6357_), .B(new_n6359_), .Y(new_n6372_));
  AOI21  g05370(.A0(new_n6361_), .A1(\A[867] ), .B0(new_n6372_), .Y(new_n6373_));
  XOR2   g05371(.A(new_n6369_), .B(new_n6362_), .Y(new_n6374_));
  INV    g05372(.A(\A[861] ), .Y(new_n6375_));
  INV    g05373(.A(\A[860] ), .Y(new_n6376_));
  NAND2  g05374(.A(new_n6376_), .B(\A[859] ), .Y(new_n6377_));
  INV    g05375(.A(\A[859] ), .Y(new_n6378_));
  AOI21  g05376(.A0(\A[860] ), .A1(new_n6378_), .B0(new_n6375_), .Y(new_n6379_));
  XOR2   g05377(.A(\A[860] ), .B(\A[859] ), .Y(new_n6380_));
  AOI22  g05378(.A0(new_n6380_), .A1(new_n6375_), .B0(new_n6379_), .B1(new_n6377_), .Y(new_n6381_));
  INV    g05379(.A(\A[864] ), .Y(new_n6382_));
  INV    g05380(.A(\A[863] ), .Y(new_n6383_));
  NAND2  g05381(.A(new_n6383_), .B(\A[862] ), .Y(new_n6384_));
  INV    g05382(.A(\A[862] ), .Y(new_n6385_));
  AOI21  g05383(.A0(\A[863] ), .A1(new_n6385_), .B0(new_n6382_), .Y(new_n6386_));
  XOR2   g05384(.A(\A[863] ), .B(\A[862] ), .Y(new_n6387_));
  AOI22  g05385(.A0(new_n6387_), .A1(new_n6382_), .B0(new_n6386_), .B1(new_n6384_), .Y(new_n6388_));
  NOR2   g05386(.A(new_n6383_), .B(new_n6385_), .Y(new_n6389_));
  AOI21  g05387(.A0(new_n6387_), .A1(\A[864] ), .B0(new_n6389_), .Y(new_n6390_));
  NOR2   g05388(.A(new_n6376_), .B(new_n6378_), .Y(new_n6391_));
  AOI21  g05389(.A0(new_n6380_), .A1(\A[861] ), .B0(new_n6391_), .Y(new_n6392_));
  XOR2   g05390(.A(new_n6388_), .B(new_n6381_), .Y(new_n6393_));
  XOR2   g05391(.A(new_n6393_), .B(new_n6374_), .Y(new_n6394_));
  INV    g05392(.A(\A[855] ), .Y(new_n6395_));
  INV    g05393(.A(\A[854] ), .Y(new_n6396_));
  NAND2  g05394(.A(new_n6396_), .B(\A[853] ), .Y(new_n6397_));
  INV    g05395(.A(\A[853] ), .Y(new_n6398_));
  AOI21  g05396(.A0(\A[854] ), .A1(new_n6398_), .B0(new_n6395_), .Y(new_n6399_));
  XOR2   g05397(.A(\A[854] ), .B(\A[853] ), .Y(new_n6400_));
  AOI22  g05398(.A0(new_n6400_), .A1(new_n6395_), .B0(new_n6399_), .B1(new_n6397_), .Y(new_n6401_));
  INV    g05399(.A(\A[858] ), .Y(new_n6402_));
  INV    g05400(.A(\A[857] ), .Y(new_n6403_));
  NAND2  g05401(.A(new_n6403_), .B(\A[856] ), .Y(new_n6404_));
  INV    g05402(.A(\A[856] ), .Y(new_n6405_));
  AOI21  g05403(.A0(\A[857] ), .A1(new_n6405_), .B0(new_n6402_), .Y(new_n6406_));
  XOR2   g05404(.A(\A[857] ), .B(\A[856] ), .Y(new_n6407_));
  AOI22  g05405(.A0(new_n6407_), .A1(new_n6402_), .B0(new_n6406_), .B1(new_n6404_), .Y(new_n6408_));
  NOR2   g05406(.A(new_n6403_), .B(new_n6405_), .Y(new_n6409_));
  AOI21  g05407(.A0(new_n6407_), .A1(\A[858] ), .B0(new_n6409_), .Y(new_n6410_));
  NOR2   g05408(.A(new_n6396_), .B(new_n6398_), .Y(new_n6411_));
  AOI21  g05409(.A0(new_n6400_), .A1(\A[855] ), .B0(new_n6411_), .Y(new_n6412_));
  XOR2   g05410(.A(new_n6408_), .B(new_n6401_), .Y(new_n6413_));
  INV    g05411(.A(\A[849] ), .Y(new_n6414_));
  INV    g05412(.A(\A[848] ), .Y(new_n6415_));
  NAND2  g05413(.A(new_n6415_), .B(\A[847] ), .Y(new_n6416_));
  INV    g05414(.A(\A[847] ), .Y(new_n6417_));
  AOI21  g05415(.A0(\A[848] ), .A1(new_n6417_), .B0(new_n6414_), .Y(new_n6418_));
  XOR2   g05416(.A(\A[848] ), .B(\A[847] ), .Y(new_n6419_));
  AOI22  g05417(.A0(new_n6419_), .A1(new_n6414_), .B0(new_n6418_), .B1(new_n6416_), .Y(new_n6420_));
  INV    g05418(.A(\A[852] ), .Y(new_n6421_));
  INV    g05419(.A(\A[851] ), .Y(new_n6422_));
  NAND2  g05420(.A(new_n6422_), .B(\A[850] ), .Y(new_n6423_));
  INV    g05421(.A(\A[850] ), .Y(new_n6424_));
  AOI21  g05422(.A0(\A[851] ), .A1(new_n6424_), .B0(new_n6421_), .Y(new_n6425_));
  XOR2   g05423(.A(\A[851] ), .B(\A[850] ), .Y(new_n6426_));
  AOI22  g05424(.A0(new_n6426_), .A1(new_n6421_), .B0(new_n6425_), .B1(new_n6423_), .Y(new_n6427_));
  NOR2   g05425(.A(new_n6422_), .B(new_n6424_), .Y(new_n6428_));
  AOI21  g05426(.A0(new_n6426_), .A1(\A[852] ), .B0(new_n6428_), .Y(new_n6429_));
  NOR2   g05427(.A(new_n6415_), .B(new_n6417_), .Y(new_n6430_));
  AOI21  g05428(.A0(new_n6419_), .A1(\A[849] ), .B0(new_n6430_), .Y(new_n6431_));
  XOR2   g05429(.A(new_n6427_), .B(new_n6420_), .Y(new_n6432_));
  XOR2   g05430(.A(new_n6432_), .B(new_n6413_), .Y(new_n6433_));
  INV    g05431(.A(new_n6433_), .Y(new_n6434_));
  XOR2   g05432(.A(new_n6434_), .B(new_n6394_), .Y(new_n6435_));
  XOR2   g05433(.A(new_n6435_), .B(new_n6355_), .Y(new_n6436_));
  XOR2   g05434(.A(new_n6436_), .B(new_n6274_), .Y(new_n6437_));
  AOI21  g05435(.A0(new_n6110_), .A1(new_n6108_), .B0(new_n6437_), .Y(new_n6438_));
  INV    g05436(.A(new_n6438_), .Y(new_n6439_));
  NOR3   g05437(.A(new_n6439_), .B(new_n6105_), .C(new_n6096_), .Y(new_n6440_));
  NOR3   g05438(.A(new_n6094_), .B(new_n6093_), .C(new_n6090_), .Y(new_n6441_));
  AOI21  g05439(.A0(new_n6082_), .A1(new_n6072_), .B0(new_n6086_), .Y(new_n6442_));
  OAI21  g05440(.A0(new_n6442_), .A1(new_n6441_), .B0(new_n6102_), .Y(new_n6443_));
  NOR3   g05441(.A(new_n6086_), .B(new_n6093_), .C(new_n6090_), .Y(new_n6444_));
  AOI21  g05442(.A0(new_n6082_), .A1(new_n6072_), .B0(new_n6094_), .Y(new_n6445_));
  OAI21  g05443(.A0(new_n6445_), .A1(new_n6444_), .B0(new_n5203_), .Y(new_n6446_));
  AOI21  g05444(.A0(new_n6446_), .A1(new_n6443_), .B0(new_n6438_), .Y(new_n6447_));
  NAND2  g05445(.A(new_n6270_), .B(new_n6231_), .Y(new_n6448_));
  XOR2   g05446(.A(new_n6225_), .B(new_n6218_), .Y(new_n6449_));
  XOR2   g05447(.A(\A[911] ), .B(new_n6222_), .Y(new_n6450_));
  NAND2  g05448(.A(\A[911] ), .B(\A[910] ), .Y(new_n6451_));
  OAI21  g05449(.A0(new_n6450_), .A1(new_n6219_), .B0(new_n6451_), .Y(new_n6452_));
  XOR2   g05450(.A(new_n6229_), .B(new_n6452_), .Y(new_n6453_));
  NOR2   g05451(.A(\A[908] ), .B(new_n6215_), .Y(new_n6454_));
  OAI21  g05452(.A0(new_n6213_), .A1(\A[907] ), .B0(\A[909] ), .Y(new_n6455_));
  XOR2   g05453(.A(\A[908] ), .B(new_n6215_), .Y(new_n6456_));
  OAI22  g05454(.A0(new_n6456_), .A1(\A[909] ), .B0(new_n6455_), .B1(new_n6454_), .Y(new_n6457_));
  NOR2   g05455(.A(\A[911] ), .B(new_n6222_), .Y(new_n6458_));
  OAI21  g05456(.A0(new_n6220_), .A1(\A[910] ), .B0(\A[912] ), .Y(new_n6459_));
  OAI22  g05457(.A0(new_n6450_), .A1(\A[912] ), .B0(new_n6459_), .B1(new_n6458_), .Y(new_n6460_));
  NAND2  g05458(.A(new_n6460_), .B(new_n6457_), .Y(new_n6461_));
  NAND2  g05459(.A(\A[908] ), .B(\A[907] ), .Y(new_n6462_));
  OAI21  g05460(.A0(new_n6456_), .A1(new_n6212_), .B0(new_n6462_), .Y(new_n6463_));
  NAND2  g05461(.A(new_n6463_), .B(new_n6452_), .Y(new_n6464_));
  OAI21  g05462(.A0(new_n6461_), .A1(new_n6453_), .B0(new_n6464_), .Y(new_n6465_));
  NOR2   g05463(.A(new_n6225_), .B(new_n6218_), .Y(new_n6466_));
  XOR2   g05464(.A(new_n6466_), .B(new_n6453_), .Y(new_n6467_));
  AOI21  g05465(.A0(new_n6465_), .A1(new_n6449_), .B0(new_n6467_), .Y(new_n6468_));
  XOR2   g05466(.A(new_n6206_), .B(new_n6199_), .Y(new_n6469_));
  NOR2   g05467(.A(\A[914] ), .B(new_n6196_), .Y(new_n6470_));
  OAI21  g05468(.A0(new_n6194_), .A1(\A[913] ), .B0(\A[915] ), .Y(new_n6471_));
  NAND2  g05469(.A(new_n6198_), .B(new_n6193_), .Y(new_n6472_));
  OAI21  g05470(.A0(new_n6471_), .A1(new_n6470_), .B0(new_n6472_), .Y(new_n6473_));
  NOR2   g05471(.A(\A[917] ), .B(new_n6203_), .Y(new_n6474_));
  OAI21  g05472(.A0(new_n6201_), .A1(\A[916] ), .B0(\A[918] ), .Y(new_n6475_));
  NAND2  g05473(.A(new_n6205_), .B(new_n6200_), .Y(new_n6476_));
  OAI21  g05474(.A0(new_n6475_), .A1(new_n6474_), .B0(new_n6476_), .Y(new_n6477_));
  NAND2  g05475(.A(new_n6205_), .B(\A[918] ), .Y(new_n6478_));
  OAI21  g05476(.A0(new_n6201_), .A1(new_n6203_), .B0(new_n6478_), .Y(new_n6479_));
  NAND2  g05477(.A(new_n6198_), .B(\A[915] ), .Y(new_n6480_));
  OAI21  g05478(.A0(new_n6194_), .A1(new_n6196_), .B0(new_n6480_), .Y(new_n6481_));
  NAND4  g05479(.A(new_n6481_), .B(new_n6479_), .C(new_n6477_), .D(new_n6473_), .Y(new_n6482_));
  NAND4  g05480(.A(new_n6463_), .B(new_n6452_), .C(new_n6460_), .D(new_n6457_), .Y(new_n6483_));
  NAND4  g05481(.A(new_n6483_), .B(new_n6449_), .C(new_n6482_), .D(new_n6469_), .Y(new_n6484_));
  XOR2   g05482(.A(new_n6210_), .B(new_n6479_), .Y(new_n6485_));
  NAND2  g05483(.A(new_n6477_), .B(new_n6473_), .Y(new_n6486_));
  NAND2  g05484(.A(new_n6481_), .B(new_n6479_), .Y(new_n6487_));
  OAI21  g05485(.A0(new_n6486_), .A1(new_n6485_), .B0(new_n6487_), .Y(new_n6488_));
  NOR2   g05486(.A(new_n6206_), .B(new_n6199_), .Y(new_n6489_));
  XOR2   g05487(.A(new_n6489_), .B(new_n6485_), .Y(new_n6490_));
  AOI21  g05488(.A0(new_n6488_), .A1(new_n6469_), .B0(new_n6490_), .Y(new_n6491_));
  XOR2   g05489(.A(new_n6491_), .B(new_n6484_), .Y(new_n6492_));
  NOR2   g05490(.A(new_n6492_), .B(new_n6468_), .Y(new_n6493_));
  XOR2   g05491(.A(new_n6206_), .B(new_n6473_), .Y(new_n6494_));
  NOR4   g05492(.A(new_n6210_), .B(new_n6208_), .C(new_n6206_), .D(new_n6199_), .Y(new_n6495_));
  XOR2   g05493(.A(new_n6225_), .B(new_n6457_), .Y(new_n6496_));
  NOR4   g05494(.A(new_n6229_), .B(new_n6227_), .C(new_n6225_), .D(new_n6218_), .Y(new_n6497_));
  NOR4   g05495(.A(new_n6497_), .B(new_n6496_), .C(new_n6495_), .D(new_n6494_), .Y(new_n6498_));
  XOR2   g05496(.A(new_n6210_), .B(new_n6208_), .Y(new_n6499_));
  XOR2   g05497(.A(new_n6489_), .B(new_n6499_), .Y(new_n6500_));
  NAND4  g05498(.A(new_n6449_), .B(new_n6482_), .C(new_n6500_), .D(new_n6469_), .Y(new_n6501_));
  NOR2   g05499(.A(new_n6210_), .B(new_n6208_), .Y(new_n6502_));
  AOI21  g05500(.A0(new_n6489_), .A1(new_n6499_), .B0(new_n6502_), .Y(new_n6503_));
  OAI21  g05501(.A0(new_n6503_), .A1(new_n6494_), .B0(new_n6483_), .Y(new_n6504_));
  OAI22  g05502(.A0(new_n6504_), .A1(new_n6501_), .B0(new_n6491_), .B1(new_n6498_), .Y(new_n6505_));
  AOI211 g05503(.A0(new_n6505_), .A1(new_n6468_), .B(new_n6448_), .C(new_n6493_), .Y(new_n6506_));
  XOR2   g05504(.A(new_n6229_), .B(new_n6227_), .Y(new_n6507_));
  NOR2   g05505(.A(new_n6229_), .B(new_n6227_), .Y(new_n6508_));
  AOI21  g05506(.A0(new_n6466_), .A1(new_n6507_), .B0(new_n6508_), .Y(new_n6509_));
  XOR2   g05507(.A(new_n6466_), .B(new_n6507_), .Y(new_n6510_));
  OAI21  g05508(.A0(new_n6509_), .A1(new_n6496_), .B0(new_n6510_), .Y(new_n6511_));
  XOR2   g05509(.A(new_n6491_), .B(new_n6498_), .Y(new_n6512_));
  NAND2  g05510(.A(new_n6512_), .B(new_n6511_), .Y(new_n6513_));
  NAND2  g05511(.A(new_n6505_), .B(new_n6468_), .Y(new_n6514_));
  NAND2  g05512(.A(new_n6514_), .B(new_n6513_), .Y(new_n6515_));
  AOI21  g05513(.A0(new_n6515_), .A1(new_n6448_), .B0(new_n6506_), .Y(new_n6516_));
  XOR2   g05514(.A(new_n6264_), .B(new_n6257_), .Y(new_n6517_));
  XOR2   g05515(.A(new_n6268_), .B(new_n6266_), .Y(new_n6518_));
  NOR2   g05516(.A(new_n6264_), .B(new_n6257_), .Y(new_n6519_));
  NAND2  g05517(.A(new_n6519_), .B(new_n6518_), .Y(new_n6520_));
  OAI21  g05518(.A0(new_n6268_), .A1(new_n6266_), .B0(new_n6520_), .Y(new_n6521_));
  INV    g05519(.A(new_n6263_), .Y(new_n6522_));
  NAND2  g05520(.A(\A[899] ), .B(\A[898] ), .Y(new_n6523_));
  OAI21  g05521(.A0(new_n6522_), .A1(new_n6258_), .B0(new_n6523_), .Y(new_n6524_));
  XOR2   g05522(.A(new_n6268_), .B(new_n6524_), .Y(new_n6525_));
  XOR2   g05523(.A(new_n6519_), .B(new_n6525_), .Y(new_n6526_));
  AOI21  g05524(.A0(new_n6521_), .A1(new_n6517_), .B0(new_n6526_), .Y(new_n6527_));
  XOR2   g05525(.A(new_n6245_), .B(new_n6238_), .Y(new_n6528_));
  NOR2   g05526(.A(\A[902] ), .B(new_n6235_), .Y(new_n6529_));
  OAI21  g05527(.A0(new_n6233_), .A1(\A[901] ), .B0(\A[903] ), .Y(new_n6530_));
  NAND2  g05528(.A(new_n6237_), .B(new_n6232_), .Y(new_n6531_));
  OAI21  g05529(.A0(new_n6530_), .A1(new_n6529_), .B0(new_n6531_), .Y(new_n6532_));
  NOR2   g05530(.A(\A[905] ), .B(new_n6242_), .Y(new_n6533_));
  OAI21  g05531(.A0(new_n6240_), .A1(\A[904] ), .B0(\A[906] ), .Y(new_n6534_));
  NAND2  g05532(.A(new_n6244_), .B(new_n6239_), .Y(new_n6535_));
  OAI21  g05533(.A0(new_n6534_), .A1(new_n6533_), .B0(new_n6535_), .Y(new_n6536_));
  NAND2  g05534(.A(new_n6244_), .B(\A[906] ), .Y(new_n6537_));
  OAI21  g05535(.A0(new_n6240_), .A1(new_n6242_), .B0(new_n6537_), .Y(new_n6538_));
  NAND2  g05536(.A(new_n6237_), .B(\A[903] ), .Y(new_n6539_));
  OAI21  g05537(.A0(new_n6233_), .A1(new_n6235_), .B0(new_n6539_), .Y(new_n6540_));
  NAND4  g05538(.A(new_n6540_), .B(new_n6538_), .C(new_n6536_), .D(new_n6532_), .Y(new_n6541_));
  INV    g05539(.A(new_n6256_), .Y(new_n6542_));
  NOR2   g05540(.A(new_n6542_), .B(new_n6251_), .Y(new_n6543_));
  OAI211 g05541(.A0(new_n6543_), .A1(new_n6267_), .B0(new_n6519_), .B1(new_n6524_), .Y(new_n6544_));
  NAND4  g05542(.A(new_n6544_), .B(new_n6517_), .C(new_n6541_), .D(new_n6528_), .Y(new_n6545_));
  XOR2   g05543(.A(new_n6249_), .B(new_n6538_), .Y(new_n6546_));
  NAND2  g05544(.A(new_n6536_), .B(new_n6532_), .Y(new_n6547_));
  NAND2  g05545(.A(new_n6540_), .B(new_n6538_), .Y(new_n6548_));
  OAI21  g05546(.A0(new_n6547_), .A1(new_n6546_), .B0(new_n6548_), .Y(new_n6549_));
  NOR2   g05547(.A(new_n6245_), .B(new_n6238_), .Y(new_n6550_));
  XOR2   g05548(.A(new_n6550_), .B(new_n6546_), .Y(new_n6551_));
  AOI21  g05549(.A0(new_n6549_), .A1(new_n6528_), .B0(new_n6551_), .Y(new_n6552_));
  XOR2   g05550(.A(new_n6552_), .B(new_n6545_), .Y(new_n6553_));
  XOR2   g05551(.A(new_n6245_), .B(new_n6532_), .Y(new_n6554_));
  XOR2   g05552(.A(new_n6249_), .B(new_n6247_), .Y(new_n6555_));
  NOR2   g05553(.A(new_n6249_), .B(new_n6247_), .Y(new_n6556_));
  AOI21  g05554(.A0(new_n6550_), .A1(new_n6555_), .B0(new_n6556_), .Y(new_n6557_));
  XOR2   g05555(.A(new_n6550_), .B(new_n6555_), .Y(new_n6558_));
  OAI21  g05556(.A0(new_n6557_), .A1(new_n6554_), .B0(new_n6558_), .Y(new_n6559_));
  NAND2  g05557(.A(new_n6559_), .B(new_n6545_), .Y(new_n6560_));
  NAND2  g05558(.A(new_n6255_), .B(new_n6253_), .Y(new_n6561_));
  OAI21  g05559(.A0(new_n6542_), .A1(\A[897] ), .B0(new_n6561_), .Y(new_n6562_));
  XOR2   g05560(.A(new_n6264_), .B(new_n6562_), .Y(new_n6563_));
  NOR4   g05561(.A(new_n6563_), .B(new_n6551_), .C(new_n6549_), .D(new_n6554_), .Y(new_n6564_));
  OAI211 g05562(.A0(new_n6557_), .A1(new_n6554_), .B0(new_n6564_), .B1(new_n6544_), .Y(new_n6565_));
  NAND2  g05563(.A(new_n6565_), .B(new_n6560_), .Y(new_n6566_));
  NAND2  g05564(.A(new_n6566_), .B(new_n6527_), .Y(new_n6567_));
  OAI21  g05565(.A0(new_n6553_), .A1(new_n6527_), .B0(new_n6567_), .Y(new_n6568_));
  NOR2   g05566(.A(new_n6568_), .B(new_n6516_), .Y(new_n6569_));
  NOR2   g05567(.A(new_n6553_), .B(new_n6527_), .Y(new_n6570_));
  NOR2   g05568(.A(new_n6268_), .B(new_n6266_), .Y(new_n6571_));
  AOI21  g05569(.A0(new_n6519_), .A1(new_n6518_), .B0(new_n6571_), .Y(new_n6572_));
  XOR2   g05570(.A(new_n6519_), .B(new_n6518_), .Y(new_n6573_));
  OAI21  g05571(.A0(new_n6572_), .A1(new_n6563_), .B0(new_n6573_), .Y(new_n6574_));
  AOI21  g05572(.A0(new_n6565_), .A1(new_n6560_), .B0(new_n6574_), .Y(new_n6575_));
  NOR2   g05573(.A(new_n6575_), .B(new_n6570_), .Y(new_n6576_));
  NAND3  g05574(.A(new_n6448_), .B(new_n6514_), .C(new_n6513_), .Y(new_n6577_));
  INV    g05575(.A(new_n6448_), .Y(new_n6578_));
  NAND2  g05576(.A(new_n6515_), .B(new_n6578_), .Y(new_n6579_));
  AOI21  g05577(.A0(new_n6579_), .A1(new_n6577_), .B0(new_n6576_), .Y(new_n6580_));
  NOR2   g05578(.A(new_n6580_), .B(new_n6569_), .Y(new_n6581_));
  XOR2   g05579(.A(new_n6183_), .B(new_n6176_), .Y(new_n6582_));
  XOR2   g05580(.A(new_n6187_), .B(new_n6185_), .Y(new_n6583_));
  NOR2   g05581(.A(new_n6183_), .B(new_n6176_), .Y(new_n6584_));
  NAND2  g05582(.A(new_n6584_), .B(new_n6583_), .Y(new_n6585_));
  OAI21  g05583(.A0(new_n6187_), .A1(new_n6185_), .B0(new_n6585_), .Y(new_n6586_));
  INV    g05584(.A(new_n6182_), .Y(new_n6587_));
  NAND2  g05585(.A(\A[923] ), .B(\A[922] ), .Y(new_n6588_));
  OAI21  g05586(.A0(new_n6587_), .A1(new_n6177_), .B0(new_n6588_), .Y(new_n6589_));
  XOR2   g05587(.A(new_n6187_), .B(new_n6589_), .Y(new_n6590_));
  XOR2   g05588(.A(new_n6584_), .B(new_n6590_), .Y(new_n6591_));
  AOI21  g05589(.A0(new_n6586_), .A1(new_n6582_), .B0(new_n6591_), .Y(new_n6592_));
  XOR2   g05590(.A(new_n6164_), .B(new_n6157_), .Y(new_n6593_));
  NOR2   g05591(.A(\A[926] ), .B(new_n6154_), .Y(new_n6594_));
  OAI21  g05592(.A0(new_n6152_), .A1(\A[925] ), .B0(\A[927] ), .Y(new_n6595_));
  NAND2  g05593(.A(new_n6156_), .B(new_n6151_), .Y(new_n6596_));
  OAI21  g05594(.A0(new_n6595_), .A1(new_n6594_), .B0(new_n6596_), .Y(new_n6597_));
  NOR2   g05595(.A(\A[929] ), .B(new_n6161_), .Y(new_n6598_));
  OAI21  g05596(.A0(new_n6159_), .A1(\A[928] ), .B0(\A[930] ), .Y(new_n6599_));
  NAND2  g05597(.A(new_n6163_), .B(new_n6158_), .Y(new_n6600_));
  OAI21  g05598(.A0(new_n6599_), .A1(new_n6598_), .B0(new_n6600_), .Y(new_n6601_));
  NAND2  g05599(.A(new_n6163_), .B(\A[930] ), .Y(new_n6602_));
  OAI21  g05600(.A0(new_n6159_), .A1(new_n6161_), .B0(new_n6602_), .Y(new_n6603_));
  NAND2  g05601(.A(new_n6156_), .B(\A[927] ), .Y(new_n6604_));
  OAI21  g05602(.A0(new_n6152_), .A1(new_n6154_), .B0(new_n6604_), .Y(new_n6605_));
  NAND4  g05603(.A(new_n6605_), .B(new_n6603_), .C(new_n6601_), .D(new_n6597_), .Y(new_n6606_));
  INV    g05604(.A(new_n6175_), .Y(new_n6607_));
  NOR2   g05605(.A(new_n6607_), .B(new_n6170_), .Y(new_n6608_));
  OAI211 g05606(.A0(new_n6608_), .A1(new_n6186_), .B0(new_n6584_), .B1(new_n6589_), .Y(new_n6609_));
  NAND4  g05607(.A(new_n6609_), .B(new_n6582_), .C(new_n6606_), .D(new_n6593_), .Y(new_n6610_));
  XOR2   g05608(.A(new_n6168_), .B(new_n6603_), .Y(new_n6611_));
  NAND2  g05609(.A(new_n6601_), .B(new_n6597_), .Y(new_n6612_));
  NAND2  g05610(.A(new_n6605_), .B(new_n6603_), .Y(new_n6613_));
  OAI21  g05611(.A0(new_n6612_), .A1(new_n6611_), .B0(new_n6613_), .Y(new_n6614_));
  NOR2   g05612(.A(new_n6164_), .B(new_n6157_), .Y(new_n6615_));
  XOR2   g05613(.A(new_n6615_), .B(new_n6611_), .Y(new_n6616_));
  AOI21  g05614(.A0(new_n6614_), .A1(new_n6593_), .B0(new_n6616_), .Y(new_n6617_));
  XOR2   g05615(.A(new_n6617_), .B(new_n6610_), .Y(new_n6618_));
  XOR2   g05616(.A(new_n6164_), .B(new_n6597_), .Y(new_n6619_));
  XOR2   g05617(.A(new_n6168_), .B(new_n6166_), .Y(new_n6620_));
  NOR2   g05618(.A(new_n6168_), .B(new_n6166_), .Y(new_n6621_));
  AOI21  g05619(.A0(new_n6615_), .A1(new_n6620_), .B0(new_n6621_), .Y(new_n6622_));
  XOR2   g05620(.A(new_n6615_), .B(new_n6620_), .Y(new_n6623_));
  OAI21  g05621(.A0(new_n6622_), .A1(new_n6619_), .B0(new_n6623_), .Y(new_n6624_));
  NAND2  g05622(.A(new_n6624_), .B(new_n6610_), .Y(new_n6625_));
  NAND2  g05623(.A(new_n6174_), .B(new_n6172_), .Y(new_n6626_));
  OAI21  g05624(.A0(new_n6607_), .A1(\A[921] ), .B0(new_n6626_), .Y(new_n6627_));
  XOR2   g05625(.A(new_n6183_), .B(new_n6627_), .Y(new_n6628_));
  NOR4   g05626(.A(new_n6628_), .B(new_n6616_), .C(new_n6614_), .D(new_n6619_), .Y(new_n6629_));
  OAI211 g05627(.A0(new_n6622_), .A1(new_n6619_), .B0(new_n6629_), .B1(new_n6609_), .Y(new_n6630_));
  NAND2  g05628(.A(new_n6630_), .B(new_n6625_), .Y(new_n6631_));
  NAND2  g05629(.A(new_n6631_), .B(new_n6592_), .Y(new_n6632_));
  OAI21  g05630(.A0(new_n6618_), .A1(new_n6592_), .B0(new_n6632_), .Y(new_n6633_));
  NOR2   g05631(.A(\A[932] ), .B(new_n6133_), .Y(new_n6634_));
  OAI21  g05632(.A0(new_n6131_), .A1(\A[931] ), .B0(\A[933] ), .Y(new_n6635_));
  XOR2   g05633(.A(\A[932] ), .B(new_n6133_), .Y(new_n6636_));
  OAI22  g05634(.A0(new_n6636_), .A1(\A[933] ), .B0(new_n6635_), .B1(new_n6634_), .Y(new_n6637_));
  XOR2   g05635(.A(new_n6143_), .B(new_n6637_), .Y(new_n6638_));
  XOR2   g05636(.A(new_n6148_), .B(new_n6146_), .Y(new_n6639_));
  NOR2   g05637(.A(new_n6143_), .B(new_n6136_), .Y(new_n6640_));
  NOR2   g05638(.A(new_n6148_), .B(new_n6146_), .Y(new_n6641_));
  AOI21  g05639(.A0(new_n6640_), .A1(new_n6639_), .B0(new_n6641_), .Y(new_n6642_));
  XOR2   g05640(.A(new_n6640_), .B(new_n6639_), .Y(new_n6643_));
  OAI21  g05641(.A0(new_n6642_), .A1(new_n6638_), .B0(new_n6643_), .Y(new_n6644_));
  NOR2   g05642(.A(\A[938] ), .B(new_n6114_), .Y(new_n6645_));
  OAI21  g05643(.A0(new_n6112_), .A1(\A[937] ), .B0(\A[939] ), .Y(new_n6646_));
  NAND2  g05644(.A(new_n6116_), .B(new_n6111_), .Y(new_n6647_));
  OAI21  g05645(.A0(new_n6646_), .A1(new_n6645_), .B0(new_n6647_), .Y(new_n6648_));
  XOR2   g05646(.A(new_n6124_), .B(new_n6648_), .Y(new_n6649_));
  NOR4   g05647(.A(new_n6128_), .B(new_n6126_), .C(new_n6124_), .D(new_n6117_), .Y(new_n6650_));
  NOR4   g05648(.A(new_n6148_), .B(new_n6146_), .C(new_n6143_), .D(new_n6136_), .Y(new_n6651_));
  NOR4   g05649(.A(new_n6651_), .B(new_n6638_), .C(new_n6650_), .D(new_n6649_), .Y(new_n6652_));
  XOR2   g05650(.A(new_n6124_), .B(new_n6117_), .Y(new_n6653_));
  NAND2  g05651(.A(new_n6123_), .B(\A[942] ), .Y(new_n6654_));
  OAI21  g05652(.A0(new_n6119_), .A1(new_n6121_), .B0(new_n6654_), .Y(new_n6655_));
  XOR2   g05653(.A(new_n6128_), .B(new_n6655_), .Y(new_n6656_));
  NOR2   g05654(.A(\A[941] ), .B(new_n6121_), .Y(new_n6657_));
  OAI21  g05655(.A0(new_n6119_), .A1(\A[940] ), .B0(\A[942] ), .Y(new_n6658_));
  NAND2  g05656(.A(new_n6123_), .B(new_n6118_), .Y(new_n6659_));
  OAI21  g05657(.A0(new_n6658_), .A1(new_n6657_), .B0(new_n6659_), .Y(new_n6660_));
  NAND2  g05658(.A(new_n6660_), .B(new_n6648_), .Y(new_n6661_));
  NAND2  g05659(.A(new_n6116_), .B(\A[939] ), .Y(new_n6662_));
  OAI21  g05660(.A0(new_n6112_), .A1(new_n6114_), .B0(new_n6662_), .Y(new_n6663_));
  NAND2  g05661(.A(new_n6663_), .B(new_n6655_), .Y(new_n6664_));
  OAI21  g05662(.A0(new_n6661_), .A1(new_n6656_), .B0(new_n6664_), .Y(new_n6665_));
  NOR2   g05663(.A(new_n6124_), .B(new_n6117_), .Y(new_n6666_));
  XOR2   g05664(.A(new_n6666_), .B(new_n6656_), .Y(new_n6667_));
  AOI21  g05665(.A0(new_n6665_), .A1(new_n6653_), .B0(new_n6667_), .Y(new_n6668_));
  XOR2   g05666(.A(new_n6668_), .B(new_n6652_), .Y(new_n6669_));
  NAND2  g05667(.A(new_n6669_), .B(new_n6644_), .Y(new_n6670_));
  XOR2   g05668(.A(new_n6143_), .B(new_n6136_), .Y(new_n6671_));
  XOR2   g05669(.A(\A[935] ), .B(new_n6140_), .Y(new_n6672_));
  OAI21  g05670(.A0(new_n6672_), .A1(new_n6137_), .B0(new_n6144_), .Y(new_n6673_));
  XOR2   g05671(.A(new_n6148_), .B(new_n6673_), .Y(new_n6674_));
  NOR2   g05672(.A(\A[935] ), .B(new_n6140_), .Y(new_n6675_));
  OAI21  g05673(.A0(new_n6138_), .A1(\A[934] ), .B0(\A[936] ), .Y(new_n6676_));
  OAI22  g05674(.A0(new_n6672_), .A1(\A[936] ), .B0(new_n6676_), .B1(new_n6675_), .Y(new_n6677_));
  NAND2  g05675(.A(new_n6677_), .B(new_n6637_), .Y(new_n6678_));
  NAND2  g05676(.A(\A[932] ), .B(\A[931] ), .Y(new_n6679_));
  OAI21  g05677(.A0(new_n6636_), .A1(new_n6130_), .B0(new_n6679_), .Y(new_n6680_));
  NAND2  g05678(.A(new_n6680_), .B(new_n6673_), .Y(new_n6681_));
  OAI21  g05679(.A0(new_n6678_), .A1(new_n6674_), .B0(new_n6681_), .Y(new_n6682_));
  XOR2   g05680(.A(new_n6640_), .B(new_n6674_), .Y(new_n6683_));
  AOI21  g05681(.A0(new_n6682_), .A1(new_n6671_), .B0(new_n6683_), .Y(new_n6684_));
  XOR2   g05682(.A(new_n6128_), .B(new_n6126_), .Y(new_n6685_));
  XOR2   g05683(.A(new_n6666_), .B(new_n6685_), .Y(new_n6686_));
  NAND4  g05684(.A(new_n6663_), .B(new_n6655_), .C(new_n6660_), .D(new_n6648_), .Y(new_n6687_));
  NAND4  g05685(.A(new_n6671_), .B(new_n6687_), .C(new_n6686_), .D(new_n6653_), .Y(new_n6688_));
  NOR2   g05686(.A(new_n6128_), .B(new_n6126_), .Y(new_n6689_));
  AOI21  g05687(.A0(new_n6666_), .A1(new_n6685_), .B0(new_n6689_), .Y(new_n6690_));
  NAND4  g05688(.A(new_n6680_), .B(new_n6673_), .C(new_n6677_), .D(new_n6637_), .Y(new_n6691_));
  OAI21  g05689(.A0(new_n6690_), .A1(new_n6649_), .B0(new_n6691_), .Y(new_n6692_));
  OAI22  g05690(.A0(new_n6692_), .A1(new_n6688_), .B0(new_n6668_), .B1(new_n6652_), .Y(new_n6693_));
  NAND2  g05691(.A(new_n6693_), .B(new_n6684_), .Y(new_n6694_));
  NAND2  g05692(.A(new_n6189_), .B(new_n6150_), .Y(new_n6695_));
  INV    g05693(.A(new_n6695_), .Y(new_n6696_));
  NAND3  g05694(.A(new_n6696_), .B(new_n6694_), .C(new_n6670_), .Y(new_n6697_));
  NAND4  g05695(.A(new_n6691_), .B(new_n6671_), .C(new_n6687_), .D(new_n6653_), .Y(new_n6698_));
  XOR2   g05696(.A(new_n6668_), .B(new_n6698_), .Y(new_n6699_));
  NOR2   g05697(.A(new_n6699_), .B(new_n6684_), .Y(new_n6700_));
  NOR2   g05698(.A(new_n6668_), .B(new_n6652_), .Y(new_n6701_));
  NOR2   g05699(.A(new_n6692_), .B(new_n6688_), .Y(new_n6702_));
  NOR2   g05700(.A(new_n6702_), .B(new_n6701_), .Y(new_n6703_));
  NOR2   g05701(.A(new_n6703_), .B(new_n6644_), .Y(new_n6704_));
  OAI21  g05702(.A0(new_n6704_), .A1(new_n6700_), .B0(new_n6695_), .Y(new_n6705_));
  AOI21  g05703(.A0(new_n6705_), .A1(new_n6697_), .B0(new_n6633_), .Y(new_n6706_));
  NOR2   g05704(.A(new_n6618_), .B(new_n6592_), .Y(new_n6707_));
  NOR2   g05705(.A(new_n6187_), .B(new_n6185_), .Y(new_n6708_));
  AOI21  g05706(.A0(new_n6584_), .A1(new_n6583_), .B0(new_n6708_), .Y(new_n6709_));
  XOR2   g05707(.A(new_n6584_), .B(new_n6583_), .Y(new_n6710_));
  OAI21  g05708(.A0(new_n6709_), .A1(new_n6628_), .B0(new_n6710_), .Y(new_n6711_));
  AOI21  g05709(.A0(new_n6630_), .A1(new_n6625_), .B0(new_n6711_), .Y(new_n6712_));
  NOR2   g05710(.A(new_n6712_), .B(new_n6707_), .Y(new_n6713_));
  NAND3  g05711(.A(new_n6695_), .B(new_n6694_), .C(new_n6670_), .Y(new_n6714_));
  OAI21  g05712(.A0(new_n6704_), .A1(new_n6700_), .B0(new_n6696_), .Y(new_n6715_));
  AOI21  g05713(.A0(new_n6715_), .A1(new_n6714_), .B0(new_n6713_), .Y(new_n6716_));
  NOR2   g05714(.A(new_n6272_), .B(new_n6191_), .Y(new_n6717_));
  INV    g05715(.A(new_n6717_), .Y(new_n6718_));
  NOR3   g05716(.A(new_n6718_), .B(new_n6716_), .C(new_n6706_), .Y(new_n6719_));
  AOI21  g05717(.A0(new_n6693_), .A1(new_n6684_), .B0(new_n6700_), .Y(new_n6720_));
  OAI21  g05718(.A0(new_n6720_), .A1(new_n6696_), .B0(new_n6697_), .Y(new_n6721_));
  NAND2  g05719(.A(new_n6721_), .B(new_n6713_), .Y(new_n6722_));
  AOI211 g05720(.A0(new_n6693_), .A1(new_n6684_), .B(new_n6696_), .C(new_n6700_), .Y(new_n6723_));
  AOI21  g05721(.A0(new_n6694_), .A1(new_n6670_), .B0(new_n6695_), .Y(new_n6724_));
  OAI22  g05722(.A0(new_n6724_), .A1(new_n6723_), .B0(new_n6712_), .B1(new_n6707_), .Y(new_n6725_));
  AOI21  g05723(.A0(new_n6725_), .A1(new_n6722_), .B0(new_n6717_), .Y(new_n6726_));
  OAI21  g05724(.A0(new_n6726_), .A1(new_n6719_), .B0(new_n6581_), .Y(new_n6727_));
  AOI211 g05725(.A0(new_n6505_), .A1(new_n6468_), .B(new_n6578_), .C(new_n6493_), .Y(new_n6728_));
  AOI21  g05726(.A0(new_n6514_), .A1(new_n6513_), .B0(new_n6448_), .Y(new_n6729_));
  OAI22  g05727(.A0(new_n6729_), .A1(new_n6728_), .B0(new_n6575_), .B1(new_n6570_), .Y(new_n6730_));
  OAI21  g05728(.A0(new_n6568_), .A1(new_n6516_), .B0(new_n6730_), .Y(new_n6731_));
  NOR3   g05729(.A(new_n6717_), .B(new_n6716_), .C(new_n6706_), .Y(new_n6732_));
  AOI21  g05730(.A0(new_n6725_), .A1(new_n6722_), .B0(new_n6718_), .Y(new_n6733_));
  OAI21  g05731(.A0(new_n6733_), .A1(new_n6732_), .B0(new_n6731_), .Y(new_n6734_));
  NOR2   g05732(.A(new_n6436_), .B(new_n6273_), .Y(new_n6735_));
  NAND3  g05733(.A(new_n6735_), .B(new_n6734_), .C(new_n6727_), .Y(new_n6736_));
  NAND3  g05734(.A(new_n6717_), .B(new_n6725_), .C(new_n6722_), .Y(new_n6737_));
  OAI21  g05735(.A0(new_n6716_), .A1(new_n6706_), .B0(new_n6718_), .Y(new_n6738_));
  AOI21  g05736(.A0(new_n6738_), .A1(new_n6737_), .B0(new_n6731_), .Y(new_n6739_));
  NAND3  g05737(.A(new_n6718_), .B(new_n6725_), .C(new_n6722_), .Y(new_n6740_));
  OAI21  g05738(.A0(new_n6716_), .A1(new_n6706_), .B0(new_n6717_), .Y(new_n6741_));
  AOI21  g05739(.A0(new_n6741_), .A1(new_n6740_), .B0(new_n6581_), .Y(new_n6742_));
  INV    g05740(.A(new_n6735_), .Y(new_n6743_));
  OAI21  g05741(.A0(new_n6742_), .A1(new_n6739_), .B0(new_n6743_), .Y(new_n6744_));
  NAND2  g05742(.A(new_n6744_), .B(new_n6736_), .Y(new_n6745_));
  XOR2   g05743(.A(new_n6346_), .B(new_n6339_), .Y(new_n6746_));
  XOR2   g05744(.A(\A[875] ), .B(new_n6343_), .Y(new_n6747_));
  NAND2  g05745(.A(\A[875] ), .B(\A[874] ), .Y(new_n6748_));
  OAI21  g05746(.A0(new_n6747_), .A1(new_n6340_), .B0(new_n6748_), .Y(new_n6749_));
  XOR2   g05747(.A(new_n6350_), .B(new_n6749_), .Y(new_n6750_));
  NOR2   g05748(.A(\A[872] ), .B(new_n6336_), .Y(new_n6751_));
  OAI21  g05749(.A0(new_n6334_), .A1(\A[871] ), .B0(\A[873] ), .Y(new_n6752_));
  XOR2   g05750(.A(\A[872] ), .B(new_n6336_), .Y(new_n6753_));
  OAI22  g05751(.A0(new_n6753_), .A1(\A[873] ), .B0(new_n6752_), .B1(new_n6751_), .Y(new_n6754_));
  NOR2   g05752(.A(\A[875] ), .B(new_n6343_), .Y(new_n6755_));
  OAI21  g05753(.A0(new_n6341_), .A1(\A[874] ), .B0(\A[876] ), .Y(new_n6756_));
  OAI22  g05754(.A0(new_n6747_), .A1(\A[876] ), .B0(new_n6756_), .B1(new_n6755_), .Y(new_n6757_));
  NAND2  g05755(.A(new_n6757_), .B(new_n6754_), .Y(new_n6758_));
  NAND2  g05756(.A(\A[872] ), .B(\A[871] ), .Y(new_n6759_));
  OAI21  g05757(.A0(new_n6753_), .A1(new_n6333_), .B0(new_n6759_), .Y(new_n6760_));
  NAND2  g05758(.A(new_n6760_), .B(new_n6749_), .Y(new_n6761_));
  OAI21  g05759(.A0(new_n6758_), .A1(new_n6750_), .B0(new_n6761_), .Y(new_n6762_));
  NOR2   g05760(.A(new_n6346_), .B(new_n6339_), .Y(new_n6763_));
  XOR2   g05761(.A(new_n6763_), .B(new_n6750_), .Y(new_n6764_));
  AOI21  g05762(.A0(new_n6762_), .A1(new_n6746_), .B0(new_n6764_), .Y(new_n6765_));
  XOR2   g05763(.A(new_n6327_), .B(new_n6320_), .Y(new_n6766_));
  NOR2   g05764(.A(\A[878] ), .B(new_n6317_), .Y(new_n6767_));
  OAI21  g05765(.A0(new_n6315_), .A1(\A[877] ), .B0(\A[879] ), .Y(new_n6768_));
  NAND2  g05766(.A(new_n6319_), .B(new_n6314_), .Y(new_n6769_));
  OAI21  g05767(.A0(new_n6768_), .A1(new_n6767_), .B0(new_n6769_), .Y(new_n6770_));
  NOR2   g05768(.A(\A[881] ), .B(new_n6324_), .Y(new_n6771_));
  OAI21  g05769(.A0(new_n6322_), .A1(\A[880] ), .B0(\A[882] ), .Y(new_n6772_));
  NAND2  g05770(.A(new_n6326_), .B(new_n6321_), .Y(new_n6773_));
  OAI21  g05771(.A0(new_n6772_), .A1(new_n6771_), .B0(new_n6773_), .Y(new_n6774_));
  NAND2  g05772(.A(new_n6326_), .B(\A[882] ), .Y(new_n6775_));
  OAI21  g05773(.A0(new_n6322_), .A1(new_n6324_), .B0(new_n6775_), .Y(new_n6776_));
  NAND2  g05774(.A(new_n6319_), .B(\A[879] ), .Y(new_n6777_));
  OAI21  g05775(.A0(new_n6315_), .A1(new_n6317_), .B0(new_n6777_), .Y(new_n6778_));
  NAND4  g05776(.A(new_n6778_), .B(new_n6776_), .C(new_n6774_), .D(new_n6770_), .Y(new_n6779_));
  NAND4  g05777(.A(new_n6760_), .B(new_n6749_), .C(new_n6757_), .D(new_n6754_), .Y(new_n6780_));
  NAND4  g05778(.A(new_n6780_), .B(new_n6746_), .C(new_n6779_), .D(new_n6766_), .Y(new_n6781_));
  XOR2   g05779(.A(new_n6331_), .B(new_n6776_), .Y(new_n6782_));
  NAND2  g05780(.A(new_n6774_), .B(new_n6770_), .Y(new_n6783_));
  NAND2  g05781(.A(new_n6778_), .B(new_n6776_), .Y(new_n6784_));
  OAI21  g05782(.A0(new_n6783_), .A1(new_n6782_), .B0(new_n6784_), .Y(new_n6785_));
  NOR2   g05783(.A(new_n6327_), .B(new_n6320_), .Y(new_n6786_));
  XOR2   g05784(.A(new_n6786_), .B(new_n6782_), .Y(new_n6787_));
  AOI21  g05785(.A0(new_n6785_), .A1(new_n6766_), .B0(new_n6787_), .Y(new_n6788_));
  XOR2   g05786(.A(new_n6788_), .B(new_n6781_), .Y(new_n6789_));
  NOR2   g05787(.A(new_n6789_), .B(new_n6765_), .Y(new_n6790_));
  XOR2   g05788(.A(new_n6327_), .B(new_n6770_), .Y(new_n6791_));
  NOR4   g05789(.A(new_n6331_), .B(new_n6329_), .C(new_n6327_), .D(new_n6320_), .Y(new_n6792_));
  XOR2   g05790(.A(new_n6346_), .B(new_n6754_), .Y(new_n6793_));
  NOR4   g05791(.A(new_n6350_), .B(new_n6348_), .C(new_n6346_), .D(new_n6339_), .Y(new_n6794_));
  NOR4   g05792(.A(new_n6794_), .B(new_n6793_), .C(new_n6792_), .D(new_n6791_), .Y(new_n6795_));
  XOR2   g05793(.A(new_n6331_), .B(new_n6329_), .Y(new_n6796_));
  NOR2   g05794(.A(new_n6331_), .B(new_n6329_), .Y(new_n6797_));
  AOI21  g05795(.A0(new_n6786_), .A1(new_n6796_), .B0(new_n6797_), .Y(new_n6798_));
  NOR4   g05796(.A(new_n6793_), .B(new_n6792_), .C(new_n6787_), .D(new_n6791_), .Y(new_n6799_));
  OAI211 g05797(.A0(new_n6798_), .A1(new_n6791_), .B0(new_n6799_), .B1(new_n6780_), .Y(new_n6800_));
  OAI21  g05798(.A0(new_n6788_), .A1(new_n6795_), .B0(new_n6800_), .Y(new_n6801_));
  AOI21  g05799(.A0(new_n6801_), .A1(new_n6765_), .B0(new_n6790_), .Y(new_n6802_));
  NOR2   g05800(.A(\A[884] ), .B(new_n6297_), .Y(new_n6803_));
  OAI21  g05801(.A0(new_n6295_), .A1(\A[883] ), .B0(\A[885] ), .Y(new_n6804_));
  XOR2   g05802(.A(\A[884] ), .B(new_n6297_), .Y(new_n6805_));
  OAI22  g05803(.A0(new_n6805_), .A1(\A[885] ), .B0(new_n6804_), .B1(new_n6803_), .Y(new_n6806_));
  XOR2   g05804(.A(new_n6307_), .B(new_n6806_), .Y(new_n6807_));
  XOR2   g05805(.A(new_n6311_), .B(new_n6309_), .Y(new_n6808_));
  NOR2   g05806(.A(new_n6307_), .B(new_n6300_), .Y(new_n6809_));
  NOR2   g05807(.A(new_n6311_), .B(new_n6309_), .Y(new_n6810_));
  AOI21  g05808(.A0(new_n6809_), .A1(new_n6808_), .B0(new_n6810_), .Y(new_n6811_));
  XOR2   g05809(.A(new_n6809_), .B(new_n6808_), .Y(new_n6812_));
  OAI21  g05810(.A0(new_n6811_), .A1(new_n6807_), .B0(new_n6812_), .Y(new_n6813_));
  NOR2   g05811(.A(\A[890] ), .B(new_n6278_), .Y(new_n6814_));
  OAI21  g05812(.A0(new_n6276_), .A1(\A[889] ), .B0(\A[891] ), .Y(new_n6815_));
  NAND2  g05813(.A(new_n6280_), .B(new_n6275_), .Y(new_n6816_));
  OAI21  g05814(.A0(new_n6815_), .A1(new_n6814_), .B0(new_n6816_), .Y(new_n6817_));
  XOR2   g05815(.A(new_n6288_), .B(new_n6817_), .Y(new_n6818_));
  NOR4   g05816(.A(new_n6292_), .B(new_n6290_), .C(new_n6288_), .D(new_n6281_), .Y(new_n6819_));
  NOR4   g05817(.A(new_n6311_), .B(new_n6309_), .C(new_n6307_), .D(new_n6300_), .Y(new_n6820_));
  NOR4   g05818(.A(new_n6820_), .B(new_n6807_), .C(new_n6819_), .D(new_n6818_), .Y(new_n6821_));
  XOR2   g05819(.A(new_n6288_), .B(new_n6281_), .Y(new_n6822_));
  NAND2  g05820(.A(new_n6287_), .B(\A[894] ), .Y(new_n6823_));
  OAI21  g05821(.A0(new_n6283_), .A1(new_n6285_), .B0(new_n6823_), .Y(new_n6824_));
  XOR2   g05822(.A(new_n6292_), .B(new_n6824_), .Y(new_n6825_));
  NOR2   g05823(.A(\A[893] ), .B(new_n6285_), .Y(new_n6826_));
  OAI21  g05824(.A0(new_n6283_), .A1(\A[892] ), .B0(\A[894] ), .Y(new_n6827_));
  NAND2  g05825(.A(new_n6287_), .B(new_n6282_), .Y(new_n6828_));
  OAI21  g05826(.A0(new_n6827_), .A1(new_n6826_), .B0(new_n6828_), .Y(new_n6829_));
  NAND2  g05827(.A(new_n6829_), .B(new_n6817_), .Y(new_n6830_));
  NAND2  g05828(.A(new_n6280_), .B(\A[891] ), .Y(new_n6831_));
  OAI21  g05829(.A0(new_n6276_), .A1(new_n6278_), .B0(new_n6831_), .Y(new_n6832_));
  NAND2  g05830(.A(new_n6832_), .B(new_n6824_), .Y(new_n6833_));
  OAI21  g05831(.A0(new_n6830_), .A1(new_n6825_), .B0(new_n6833_), .Y(new_n6834_));
  NOR2   g05832(.A(new_n6288_), .B(new_n6281_), .Y(new_n6835_));
  XOR2   g05833(.A(new_n6835_), .B(new_n6825_), .Y(new_n6836_));
  AOI21  g05834(.A0(new_n6834_), .A1(new_n6822_), .B0(new_n6836_), .Y(new_n6837_));
  XOR2   g05835(.A(new_n6837_), .B(new_n6821_), .Y(new_n6838_));
  NAND2  g05836(.A(new_n6838_), .B(new_n6813_), .Y(new_n6839_));
  XOR2   g05837(.A(new_n6307_), .B(new_n6300_), .Y(new_n6840_));
  XOR2   g05838(.A(\A[887] ), .B(new_n6304_), .Y(new_n6841_));
  NAND2  g05839(.A(\A[887] ), .B(\A[886] ), .Y(new_n6842_));
  OAI21  g05840(.A0(new_n6841_), .A1(new_n6301_), .B0(new_n6842_), .Y(new_n6843_));
  XOR2   g05841(.A(new_n6311_), .B(new_n6843_), .Y(new_n6844_));
  NOR2   g05842(.A(\A[887] ), .B(new_n6304_), .Y(new_n6845_));
  OAI21  g05843(.A0(new_n6302_), .A1(\A[886] ), .B0(\A[888] ), .Y(new_n6846_));
  OAI22  g05844(.A0(new_n6841_), .A1(\A[888] ), .B0(new_n6846_), .B1(new_n6845_), .Y(new_n6847_));
  NAND2  g05845(.A(new_n6847_), .B(new_n6806_), .Y(new_n6848_));
  NAND2  g05846(.A(\A[884] ), .B(\A[883] ), .Y(new_n6849_));
  OAI21  g05847(.A0(new_n6805_), .A1(new_n6294_), .B0(new_n6849_), .Y(new_n6850_));
  NAND2  g05848(.A(new_n6850_), .B(new_n6843_), .Y(new_n6851_));
  OAI21  g05849(.A0(new_n6848_), .A1(new_n6844_), .B0(new_n6851_), .Y(new_n6852_));
  XOR2   g05850(.A(new_n6809_), .B(new_n6844_), .Y(new_n6853_));
  AOI21  g05851(.A0(new_n6852_), .A1(new_n6840_), .B0(new_n6853_), .Y(new_n6854_));
  XOR2   g05852(.A(new_n6292_), .B(new_n6290_), .Y(new_n6855_));
  XOR2   g05853(.A(new_n6835_), .B(new_n6855_), .Y(new_n6856_));
  NAND4  g05854(.A(new_n6832_), .B(new_n6824_), .C(new_n6829_), .D(new_n6817_), .Y(new_n6857_));
  NAND4  g05855(.A(new_n6840_), .B(new_n6857_), .C(new_n6856_), .D(new_n6822_), .Y(new_n6858_));
  NOR2   g05856(.A(new_n6292_), .B(new_n6290_), .Y(new_n6859_));
  AOI21  g05857(.A0(new_n6835_), .A1(new_n6855_), .B0(new_n6859_), .Y(new_n6860_));
  NAND4  g05858(.A(new_n6850_), .B(new_n6843_), .C(new_n6847_), .D(new_n6806_), .Y(new_n6861_));
  OAI21  g05859(.A0(new_n6860_), .A1(new_n6818_), .B0(new_n6861_), .Y(new_n6862_));
  OAI22  g05860(.A0(new_n6862_), .A1(new_n6858_), .B0(new_n6837_), .B1(new_n6821_), .Y(new_n6863_));
  NAND2  g05861(.A(new_n6863_), .B(new_n6854_), .Y(new_n6864_));
  NAND2  g05862(.A(new_n6352_), .B(new_n6313_), .Y(new_n6865_));
  INV    g05863(.A(new_n6865_), .Y(new_n6866_));
  NAND3  g05864(.A(new_n6866_), .B(new_n6864_), .C(new_n6839_), .Y(new_n6867_));
  NAND4  g05865(.A(new_n6861_), .B(new_n6840_), .C(new_n6857_), .D(new_n6822_), .Y(new_n6868_));
  XOR2   g05866(.A(new_n6837_), .B(new_n6868_), .Y(new_n6869_));
  NOR2   g05867(.A(new_n6869_), .B(new_n6854_), .Y(new_n6870_));
  OAI21  g05868(.A0(new_n6860_), .A1(new_n6818_), .B0(new_n6856_), .Y(new_n6871_));
  NAND2  g05869(.A(new_n6871_), .B(new_n6868_), .Y(new_n6872_));
  NOR4   g05870(.A(new_n6807_), .B(new_n6819_), .C(new_n6836_), .D(new_n6818_), .Y(new_n6873_));
  OAI211 g05871(.A0(new_n6860_), .A1(new_n6818_), .B0(new_n6873_), .B1(new_n6861_), .Y(new_n6874_));
  AOI21  g05872(.A0(new_n6874_), .A1(new_n6872_), .B0(new_n6813_), .Y(new_n6875_));
  OAI21  g05873(.A0(new_n6875_), .A1(new_n6870_), .B0(new_n6865_), .Y(new_n6876_));
  NAND2  g05874(.A(new_n6876_), .B(new_n6867_), .Y(new_n6877_));
  NAND2  g05875(.A(new_n6877_), .B(new_n6802_), .Y(new_n6878_));
  XOR2   g05876(.A(new_n6786_), .B(new_n6796_), .Y(new_n6879_));
  OAI21  g05877(.A0(new_n6798_), .A1(new_n6791_), .B0(new_n6879_), .Y(new_n6880_));
  NAND2  g05878(.A(new_n6880_), .B(new_n6781_), .Y(new_n6881_));
  AOI221 g05879(.A0(new_n6800_), .A1(new_n6881_), .C0(new_n6764_), .B0(new_n6762_), .B1(new_n6746_), .Y(new_n6882_));
  NOR3   g05880(.A(new_n6866_), .B(new_n6875_), .C(new_n6870_), .Y(new_n6883_));
  AOI21  g05881(.A0(new_n6864_), .A1(new_n6839_), .B0(new_n6865_), .Y(new_n6884_));
  OAI22  g05882(.A0(new_n6884_), .A1(new_n6883_), .B0(new_n6882_), .B1(new_n6790_), .Y(new_n6885_));
  NOR2   g05883(.A(new_n6435_), .B(new_n6354_), .Y(new_n6886_));
  NAND3  g05884(.A(new_n6886_), .B(new_n6885_), .C(new_n6878_), .Y(new_n6887_));
  AOI221 g05885(.A0(new_n6876_), .A1(new_n6867_), .C0(new_n6790_), .B0(new_n6801_), .B1(new_n6765_), .Y(new_n6888_));
  NAND3  g05886(.A(new_n6865_), .B(new_n6864_), .C(new_n6839_), .Y(new_n6889_));
  OAI21  g05887(.A0(new_n6875_), .A1(new_n6870_), .B0(new_n6866_), .Y(new_n6890_));
  AOI21  g05888(.A0(new_n6890_), .A1(new_n6889_), .B0(new_n6802_), .Y(new_n6891_));
  INV    g05889(.A(new_n6886_), .Y(new_n6892_));
  OAI21  g05890(.A0(new_n6891_), .A1(new_n6888_), .B0(new_n6892_), .Y(new_n6893_));
  XOR2   g05891(.A(new_n6388_), .B(new_n6381_), .Y(new_n6894_));
  XOR2   g05892(.A(\A[863] ), .B(new_n6385_), .Y(new_n6895_));
  NAND2  g05893(.A(\A[863] ), .B(\A[862] ), .Y(new_n6896_));
  OAI21  g05894(.A0(new_n6895_), .A1(new_n6382_), .B0(new_n6896_), .Y(new_n6897_));
  XOR2   g05895(.A(new_n6392_), .B(new_n6897_), .Y(new_n6898_));
  NOR2   g05896(.A(\A[860] ), .B(new_n6378_), .Y(new_n6899_));
  OAI21  g05897(.A0(new_n6376_), .A1(\A[859] ), .B0(\A[861] ), .Y(new_n6900_));
  XOR2   g05898(.A(\A[860] ), .B(new_n6378_), .Y(new_n6901_));
  OAI22  g05899(.A0(new_n6901_), .A1(\A[861] ), .B0(new_n6900_), .B1(new_n6899_), .Y(new_n6902_));
  NOR2   g05900(.A(\A[863] ), .B(new_n6385_), .Y(new_n6903_));
  OAI21  g05901(.A0(new_n6383_), .A1(\A[862] ), .B0(\A[864] ), .Y(new_n6904_));
  OAI22  g05902(.A0(new_n6895_), .A1(\A[864] ), .B0(new_n6904_), .B1(new_n6903_), .Y(new_n6905_));
  NAND2  g05903(.A(new_n6905_), .B(new_n6902_), .Y(new_n6906_));
  NAND2  g05904(.A(\A[860] ), .B(\A[859] ), .Y(new_n6907_));
  OAI21  g05905(.A0(new_n6901_), .A1(new_n6375_), .B0(new_n6907_), .Y(new_n6908_));
  NAND2  g05906(.A(new_n6908_), .B(new_n6897_), .Y(new_n6909_));
  OAI21  g05907(.A0(new_n6906_), .A1(new_n6898_), .B0(new_n6909_), .Y(new_n6910_));
  NOR2   g05908(.A(new_n6388_), .B(new_n6381_), .Y(new_n6911_));
  XOR2   g05909(.A(new_n6911_), .B(new_n6898_), .Y(new_n6912_));
  AOI21  g05910(.A0(new_n6910_), .A1(new_n6894_), .B0(new_n6912_), .Y(new_n6913_));
  XOR2   g05911(.A(new_n6369_), .B(new_n6362_), .Y(new_n6914_));
  NOR2   g05912(.A(\A[866] ), .B(new_n6359_), .Y(new_n6915_));
  OAI21  g05913(.A0(new_n6357_), .A1(\A[865] ), .B0(\A[867] ), .Y(new_n6916_));
  NAND2  g05914(.A(new_n6361_), .B(new_n6356_), .Y(new_n6917_));
  OAI21  g05915(.A0(new_n6916_), .A1(new_n6915_), .B0(new_n6917_), .Y(new_n6918_));
  NOR2   g05916(.A(\A[869] ), .B(new_n6366_), .Y(new_n6919_));
  OAI21  g05917(.A0(new_n6364_), .A1(\A[868] ), .B0(\A[870] ), .Y(new_n6920_));
  NAND2  g05918(.A(new_n6368_), .B(new_n6363_), .Y(new_n6921_));
  OAI21  g05919(.A0(new_n6920_), .A1(new_n6919_), .B0(new_n6921_), .Y(new_n6922_));
  NAND2  g05920(.A(new_n6368_), .B(\A[870] ), .Y(new_n6923_));
  OAI21  g05921(.A0(new_n6364_), .A1(new_n6366_), .B0(new_n6923_), .Y(new_n6924_));
  NAND2  g05922(.A(new_n6361_), .B(\A[867] ), .Y(new_n6925_));
  OAI21  g05923(.A0(new_n6357_), .A1(new_n6359_), .B0(new_n6925_), .Y(new_n6926_));
  NAND4  g05924(.A(new_n6926_), .B(new_n6924_), .C(new_n6922_), .D(new_n6918_), .Y(new_n6927_));
  NAND4  g05925(.A(new_n6908_), .B(new_n6897_), .C(new_n6905_), .D(new_n6902_), .Y(new_n6928_));
  NAND4  g05926(.A(new_n6928_), .B(new_n6894_), .C(new_n6927_), .D(new_n6914_), .Y(new_n6929_));
  XOR2   g05927(.A(new_n6373_), .B(new_n6924_), .Y(new_n6930_));
  NAND2  g05928(.A(new_n6922_), .B(new_n6918_), .Y(new_n6931_));
  NAND2  g05929(.A(new_n6926_), .B(new_n6924_), .Y(new_n6932_));
  OAI21  g05930(.A0(new_n6931_), .A1(new_n6930_), .B0(new_n6932_), .Y(new_n6933_));
  NOR2   g05931(.A(new_n6369_), .B(new_n6362_), .Y(new_n6934_));
  XOR2   g05932(.A(new_n6934_), .B(new_n6930_), .Y(new_n6935_));
  AOI21  g05933(.A0(new_n6933_), .A1(new_n6914_), .B0(new_n6935_), .Y(new_n6936_));
  XOR2   g05934(.A(new_n6936_), .B(new_n6929_), .Y(new_n6937_));
  NOR2   g05935(.A(new_n6937_), .B(new_n6913_), .Y(new_n6938_));
  XOR2   g05936(.A(new_n6388_), .B(new_n6902_), .Y(new_n6939_));
  XOR2   g05937(.A(new_n6392_), .B(new_n6390_), .Y(new_n6940_));
  NOR2   g05938(.A(new_n6392_), .B(new_n6390_), .Y(new_n6941_));
  AOI21  g05939(.A0(new_n6911_), .A1(new_n6940_), .B0(new_n6941_), .Y(new_n6942_));
  XOR2   g05940(.A(new_n6911_), .B(new_n6940_), .Y(new_n6943_));
  OAI21  g05941(.A0(new_n6942_), .A1(new_n6939_), .B0(new_n6943_), .Y(new_n6944_));
  XOR2   g05942(.A(new_n6369_), .B(new_n6918_), .Y(new_n6945_));
  XOR2   g05943(.A(new_n6373_), .B(new_n6371_), .Y(new_n6946_));
  NOR2   g05944(.A(new_n6373_), .B(new_n6371_), .Y(new_n6947_));
  AOI21  g05945(.A0(new_n6934_), .A1(new_n6946_), .B0(new_n6947_), .Y(new_n6948_));
  XOR2   g05946(.A(new_n6934_), .B(new_n6946_), .Y(new_n6949_));
  OAI21  g05947(.A0(new_n6948_), .A1(new_n6945_), .B0(new_n6949_), .Y(new_n6950_));
  NAND2  g05948(.A(new_n6950_), .B(new_n6929_), .Y(new_n6951_));
  NOR4   g05949(.A(new_n6373_), .B(new_n6371_), .C(new_n6369_), .D(new_n6362_), .Y(new_n6952_));
  NOR4   g05950(.A(new_n6939_), .B(new_n6952_), .C(new_n6935_), .D(new_n6945_), .Y(new_n6953_));
  OAI211 g05951(.A0(new_n6948_), .A1(new_n6945_), .B0(new_n6953_), .B1(new_n6928_), .Y(new_n6954_));
  AOI21  g05952(.A0(new_n6954_), .A1(new_n6951_), .B0(new_n6944_), .Y(new_n6955_));
  NAND2  g05953(.A(new_n6433_), .B(new_n6394_), .Y(new_n6956_));
  NOR3   g05954(.A(new_n6956_), .B(new_n6955_), .C(new_n6938_), .Y(new_n6957_));
  NOR4   g05955(.A(new_n6392_), .B(new_n6390_), .C(new_n6388_), .D(new_n6381_), .Y(new_n6958_));
  NOR4   g05956(.A(new_n6958_), .B(new_n6939_), .C(new_n6952_), .D(new_n6945_), .Y(new_n6959_));
  XOR2   g05957(.A(new_n6936_), .B(new_n6959_), .Y(new_n6960_));
  NAND2  g05958(.A(new_n6960_), .B(new_n6944_), .Y(new_n6961_));
  NAND4  g05959(.A(new_n6894_), .B(new_n6927_), .C(new_n6949_), .D(new_n6914_), .Y(new_n6962_));
  OAI21  g05960(.A0(new_n6948_), .A1(new_n6945_), .B0(new_n6928_), .Y(new_n6963_));
  OAI22  g05961(.A0(new_n6963_), .A1(new_n6962_), .B0(new_n6936_), .B1(new_n6959_), .Y(new_n6964_));
  NAND2  g05962(.A(new_n6964_), .B(new_n6913_), .Y(new_n6965_));
  INV    g05963(.A(new_n6956_), .Y(new_n6966_));
  AOI21  g05964(.A0(new_n6965_), .A1(new_n6961_), .B0(new_n6966_), .Y(new_n6967_));
  NOR2   g05965(.A(new_n6967_), .B(new_n6957_), .Y(new_n6968_));
  XOR2   g05966(.A(new_n6427_), .B(new_n6420_), .Y(new_n6969_));
  XOR2   g05967(.A(\A[851] ), .B(new_n6424_), .Y(new_n6970_));
  NAND2  g05968(.A(\A[851] ), .B(\A[850] ), .Y(new_n6971_));
  OAI21  g05969(.A0(new_n6970_), .A1(new_n6421_), .B0(new_n6971_), .Y(new_n6972_));
  XOR2   g05970(.A(new_n6431_), .B(new_n6972_), .Y(new_n6973_));
  NOR2   g05971(.A(\A[848] ), .B(new_n6417_), .Y(new_n6974_));
  OAI21  g05972(.A0(new_n6415_), .A1(\A[847] ), .B0(\A[849] ), .Y(new_n6975_));
  XOR2   g05973(.A(\A[848] ), .B(new_n6417_), .Y(new_n6976_));
  OAI22  g05974(.A0(new_n6976_), .A1(\A[849] ), .B0(new_n6975_), .B1(new_n6974_), .Y(new_n6977_));
  NOR2   g05975(.A(\A[851] ), .B(new_n6424_), .Y(new_n6978_));
  OAI21  g05976(.A0(new_n6422_), .A1(\A[850] ), .B0(\A[852] ), .Y(new_n6979_));
  OAI22  g05977(.A0(new_n6970_), .A1(\A[852] ), .B0(new_n6979_), .B1(new_n6978_), .Y(new_n6980_));
  NAND2  g05978(.A(new_n6980_), .B(new_n6977_), .Y(new_n6981_));
  NAND2  g05979(.A(\A[848] ), .B(\A[847] ), .Y(new_n6982_));
  OAI21  g05980(.A0(new_n6976_), .A1(new_n6414_), .B0(new_n6982_), .Y(new_n6983_));
  NAND2  g05981(.A(new_n6983_), .B(new_n6972_), .Y(new_n6984_));
  OAI21  g05982(.A0(new_n6981_), .A1(new_n6973_), .B0(new_n6984_), .Y(new_n6985_));
  NOR2   g05983(.A(new_n6427_), .B(new_n6420_), .Y(new_n6986_));
  XOR2   g05984(.A(new_n6986_), .B(new_n6973_), .Y(new_n6987_));
  AOI21  g05985(.A0(new_n6985_), .A1(new_n6969_), .B0(new_n6987_), .Y(new_n6988_));
  XOR2   g05986(.A(new_n6408_), .B(new_n6401_), .Y(new_n6989_));
  NOR2   g05987(.A(\A[854] ), .B(new_n6398_), .Y(new_n6990_));
  OAI21  g05988(.A0(new_n6396_), .A1(\A[853] ), .B0(\A[855] ), .Y(new_n6991_));
  NAND2  g05989(.A(new_n6400_), .B(new_n6395_), .Y(new_n6992_));
  OAI21  g05990(.A0(new_n6991_), .A1(new_n6990_), .B0(new_n6992_), .Y(new_n6993_));
  NOR2   g05991(.A(\A[857] ), .B(new_n6405_), .Y(new_n6994_));
  OAI21  g05992(.A0(new_n6403_), .A1(\A[856] ), .B0(\A[858] ), .Y(new_n6995_));
  NAND2  g05993(.A(new_n6407_), .B(new_n6402_), .Y(new_n6996_));
  OAI21  g05994(.A0(new_n6995_), .A1(new_n6994_), .B0(new_n6996_), .Y(new_n6997_));
  NAND2  g05995(.A(new_n6407_), .B(\A[858] ), .Y(new_n6998_));
  OAI21  g05996(.A0(new_n6403_), .A1(new_n6405_), .B0(new_n6998_), .Y(new_n6999_));
  NAND2  g05997(.A(new_n6400_), .B(\A[855] ), .Y(new_n7000_));
  OAI21  g05998(.A0(new_n6396_), .A1(new_n6398_), .B0(new_n7000_), .Y(new_n7001_));
  NAND4  g05999(.A(new_n7001_), .B(new_n6999_), .C(new_n6997_), .D(new_n6993_), .Y(new_n7002_));
  NAND4  g06000(.A(new_n6983_), .B(new_n6972_), .C(new_n6980_), .D(new_n6977_), .Y(new_n7003_));
  NAND4  g06001(.A(new_n7003_), .B(new_n6969_), .C(new_n7002_), .D(new_n6989_), .Y(new_n7004_));
  XOR2   g06002(.A(new_n6412_), .B(new_n6999_), .Y(new_n7005_));
  NAND2  g06003(.A(new_n6997_), .B(new_n6993_), .Y(new_n7006_));
  NAND2  g06004(.A(new_n7001_), .B(new_n6999_), .Y(new_n7007_));
  OAI21  g06005(.A0(new_n7006_), .A1(new_n7005_), .B0(new_n7007_), .Y(new_n7008_));
  NOR2   g06006(.A(new_n6408_), .B(new_n6401_), .Y(new_n7009_));
  XOR2   g06007(.A(new_n7009_), .B(new_n7005_), .Y(new_n7010_));
  AOI21  g06008(.A0(new_n7008_), .A1(new_n6989_), .B0(new_n7010_), .Y(new_n7011_));
  XOR2   g06009(.A(new_n7011_), .B(new_n7004_), .Y(new_n7012_));
  XOR2   g06010(.A(new_n6408_), .B(new_n6993_), .Y(new_n7013_));
  NOR4   g06011(.A(new_n6412_), .B(new_n6410_), .C(new_n6408_), .D(new_n6401_), .Y(new_n7014_));
  XOR2   g06012(.A(new_n6427_), .B(new_n6977_), .Y(new_n7015_));
  NOR4   g06013(.A(new_n6431_), .B(new_n6429_), .C(new_n6427_), .D(new_n6420_), .Y(new_n7016_));
  NOR4   g06014(.A(new_n7016_), .B(new_n7015_), .C(new_n7014_), .D(new_n7013_), .Y(new_n7017_));
  XOR2   g06015(.A(new_n6412_), .B(new_n6410_), .Y(new_n7018_));
  NOR2   g06016(.A(new_n6412_), .B(new_n6410_), .Y(new_n7019_));
  AOI21  g06017(.A0(new_n7009_), .A1(new_n7018_), .B0(new_n7019_), .Y(new_n7020_));
  NOR4   g06018(.A(new_n7015_), .B(new_n7014_), .C(new_n7010_), .D(new_n7013_), .Y(new_n7021_));
  OAI211 g06019(.A0(new_n7020_), .A1(new_n7013_), .B0(new_n7021_), .B1(new_n7003_), .Y(new_n7022_));
  OAI21  g06020(.A0(new_n7011_), .A1(new_n7017_), .B0(new_n7022_), .Y(new_n7023_));
  NAND2  g06021(.A(new_n7023_), .B(new_n6988_), .Y(new_n7024_));
  OAI21  g06022(.A0(new_n7012_), .A1(new_n6988_), .B0(new_n7024_), .Y(new_n7025_));
  NOR2   g06023(.A(new_n6955_), .B(new_n6938_), .Y(new_n7026_));
  NAND3  g06024(.A(new_n6956_), .B(new_n6965_), .C(new_n6961_), .Y(new_n7027_));
  OAI21  g06025(.A0(new_n7026_), .A1(new_n6956_), .B0(new_n7027_), .Y(new_n7028_));
  NAND2  g06026(.A(new_n7028_), .B(new_n7025_), .Y(new_n7029_));
  OAI21  g06027(.A0(new_n7025_), .A1(new_n6968_), .B0(new_n7029_), .Y(new_n7030_));
  AOI21  g06028(.A0(new_n6893_), .A1(new_n6887_), .B0(new_n7030_), .Y(new_n7031_));
  NOR2   g06029(.A(new_n7025_), .B(new_n6968_), .Y(new_n7032_));
  AOI21  g06030(.A0(new_n7028_), .A1(new_n7025_), .B0(new_n7032_), .Y(new_n7033_));
  NAND3  g06031(.A(new_n6892_), .B(new_n6885_), .C(new_n6878_), .Y(new_n7034_));
  OAI21  g06032(.A0(new_n6891_), .A1(new_n6888_), .B0(new_n6886_), .Y(new_n7035_));
  AOI21  g06033(.A0(new_n7035_), .A1(new_n7034_), .B0(new_n7033_), .Y(new_n7036_));
  NOR2   g06034(.A(new_n7036_), .B(new_n7031_), .Y(new_n7037_));
  NAND3  g06035(.A(new_n6743_), .B(new_n6734_), .C(new_n6727_), .Y(new_n7038_));
  OAI21  g06036(.A0(new_n6742_), .A1(new_n6739_), .B0(new_n6735_), .Y(new_n7039_));
  AOI21  g06037(.A0(new_n7039_), .A1(new_n7038_), .B0(new_n7037_), .Y(new_n7040_));
  AOI21  g06038(.A0(new_n7037_), .A1(new_n6745_), .B0(new_n7040_), .Y(new_n7041_));
  OAI21  g06039(.A0(new_n6447_), .A1(new_n6440_), .B0(new_n7041_), .Y(new_n7042_));
  NAND2  g06040(.A(new_n7037_), .B(new_n6745_), .Y(new_n7043_));
  NOR3   g06041(.A(new_n6892_), .B(new_n6891_), .C(new_n6888_), .Y(new_n7044_));
  AOI21  g06042(.A0(new_n6885_), .A1(new_n6878_), .B0(new_n6886_), .Y(new_n7045_));
  OAI21  g06043(.A0(new_n7045_), .A1(new_n7044_), .B0(new_n7033_), .Y(new_n7046_));
  NOR3   g06044(.A(new_n6886_), .B(new_n6891_), .C(new_n6888_), .Y(new_n7047_));
  AOI21  g06045(.A0(new_n6885_), .A1(new_n6878_), .B0(new_n6892_), .Y(new_n7048_));
  OAI21  g06046(.A0(new_n7048_), .A1(new_n7047_), .B0(new_n7030_), .Y(new_n7049_));
  NAND2  g06047(.A(new_n7049_), .B(new_n7046_), .Y(new_n7050_));
  NOR3   g06048(.A(new_n6735_), .B(new_n6742_), .C(new_n6739_), .Y(new_n7051_));
  AOI21  g06049(.A0(new_n6734_), .A1(new_n6727_), .B0(new_n6743_), .Y(new_n7052_));
  OAI21  g06050(.A0(new_n7052_), .A1(new_n7051_), .B0(new_n7050_), .Y(new_n7053_));
  NAND2  g06051(.A(new_n7053_), .B(new_n7043_), .Y(new_n7054_));
  NOR3   g06052(.A(new_n6438_), .B(new_n6105_), .C(new_n6096_), .Y(new_n7055_));
  AOI21  g06053(.A0(new_n6446_), .A1(new_n6443_), .B0(new_n6439_), .Y(new_n7056_));
  OAI21  g06054(.A0(new_n7056_), .A1(new_n7055_), .B0(new_n7054_), .Y(new_n7057_));
  NAND2  g06055(.A(new_n7057_), .B(new_n7042_), .Y(new_n7058_));
  INV    g06056(.A(\A[200] ), .Y(new_n7059_));
  NOR2   g06057(.A(new_n7059_), .B(\A[199] ), .Y(new_n7060_));
  INV    g06058(.A(\A[199] ), .Y(new_n7061_));
  OAI21  g06059(.A0(\A[200] ), .A1(new_n7061_), .B0(\A[201] ), .Y(new_n7062_));
  XOR2   g06060(.A(\A[200] ), .B(new_n7061_), .Y(new_n7063_));
  OAI22  g06061(.A0(new_n7063_), .A1(\A[201] ), .B0(new_n7062_), .B1(new_n7060_), .Y(new_n7064_));
  INV    g06062(.A(\A[203] ), .Y(new_n7065_));
  NOR2   g06063(.A(new_n7065_), .B(\A[202] ), .Y(new_n7066_));
  INV    g06064(.A(\A[202] ), .Y(new_n7067_));
  OAI21  g06065(.A0(\A[203] ), .A1(new_n7067_), .B0(\A[204] ), .Y(new_n7068_));
  XOR2   g06066(.A(\A[203] ), .B(new_n7067_), .Y(new_n7069_));
  OAI22  g06067(.A0(new_n7069_), .A1(\A[204] ), .B0(new_n7068_), .B1(new_n7066_), .Y(new_n7070_));
  NAND2  g06068(.A(new_n7070_), .B(new_n7064_), .Y(new_n7071_));
  INV    g06069(.A(\A[204] ), .Y(new_n7072_));
  NAND2  g06070(.A(\A[203] ), .B(\A[202] ), .Y(new_n7073_));
  OAI21  g06071(.A0(new_n7069_), .A1(new_n7072_), .B0(new_n7073_), .Y(new_n7074_));
  XOR2   g06072(.A(\A[200] ), .B(\A[199] ), .Y(new_n7075_));
  NOR2   g06073(.A(new_n7059_), .B(new_n7061_), .Y(new_n7076_));
  AOI21  g06074(.A0(new_n7075_), .A1(\A[201] ), .B0(new_n7076_), .Y(new_n7077_));
  XOR2   g06075(.A(new_n7077_), .B(new_n7074_), .Y(new_n7078_));
  XOR2   g06076(.A(new_n7078_), .B(new_n7071_), .Y(new_n7079_));
  NAND2  g06077(.A(\A[203] ), .B(new_n7067_), .Y(new_n7080_));
  AOI21  g06078(.A0(new_n7065_), .A1(\A[202] ), .B0(new_n7072_), .Y(new_n7081_));
  XOR2   g06079(.A(\A[203] ), .B(\A[202] ), .Y(new_n7082_));
  AOI22  g06080(.A0(new_n7082_), .A1(new_n7072_), .B0(new_n7081_), .B1(new_n7080_), .Y(new_n7083_));
  XOR2   g06081(.A(new_n7083_), .B(new_n7064_), .Y(new_n7084_));
  INV    g06082(.A(\A[201] ), .Y(new_n7085_));
  NAND2  g06083(.A(\A[200] ), .B(new_n7061_), .Y(new_n7086_));
  AOI21  g06084(.A0(new_n7059_), .A1(\A[199] ), .B0(new_n7085_), .Y(new_n7087_));
  AOI22  g06085(.A0(new_n7075_), .A1(new_n7085_), .B0(new_n7087_), .B1(new_n7086_), .Y(new_n7088_));
  NOR2   g06086(.A(new_n7083_), .B(new_n7088_), .Y(new_n7089_));
  NOR2   g06087(.A(new_n7065_), .B(new_n7067_), .Y(new_n7090_));
  AOI21  g06088(.A0(new_n7082_), .A1(\A[204] ), .B0(new_n7090_), .Y(new_n7091_));
  XOR2   g06089(.A(new_n7077_), .B(new_n7091_), .Y(new_n7092_));
  NOR2   g06090(.A(new_n7077_), .B(new_n7091_), .Y(new_n7093_));
  AOI21  g06091(.A0(new_n7092_), .A1(new_n7089_), .B0(new_n7093_), .Y(new_n7094_));
  OAI21  g06092(.A0(new_n7094_), .A1(new_n7084_), .B0(new_n7079_), .Y(new_n7095_));
  XOR2   g06093(.A(new_n7083_), .B(new_n7088_), .Y(new_n7096_));
  NAND2  g06094(.A(\A[209] ), .B(\A[208] ), .Y(new_n7097_));
  XOR2   g06095(.A(\A[209] ), .B(\A[208] ), .Y(new_n7098_));
  NAND2  g06096(.A(new_n7098_), .B(\A[210] ), .Y(new_n7099_));
  NAND2  g06097(.A(new_n7099_), .B(new_n7097_), .Y(new_n7100_));
  NAND2  g06098(.A(\A[206] ), .B(\A[205] ), .Y(new_n7101_));
  XOR2   g06099(.A(\A[206] ), .B(\A[205] ), .Y(new_n7102_));
  NAND2  g06100(.A(new_n7102_), .B(\A[207] ), .Y(new_n7103_));
  NAND2  g06101(.A(new_n7103_), .B(new_n7101_), .Y(new_n7104_));
  INV    g06102(.A(\A[206] ), .Y(new_n7105_));
  NOR2   g06103(.A(new_n7105_), .B(\A[205] ), .Y(new_n7106_));
  INV    g06104(.A(\A[205] ), .Y(new_n7107_));
  OAI21  g06105(.A0(\A[206] ), .A1(new_n7107_), .B0(\A[207] ), .Y(new_n7108_));
  INV    g06106(.A(\A[207] ), .Y(new_n7109_));
  NAND2  g06107(.A(new_n7102_), .B(new_n7109_), .Y(new_n7110_));
  OAI21  g06108(.A0(new_n7108_), .A1(new_n7106_), .B0(new_n7110_), .Y(new_n7111_));
  INV    g06109(.A(\A[209] ), .Y(new_n7112_));
  NOR2   g06110(.A(new_n7112_), .B(\A[208] ), .Y(new_n7113_));
  INV    g06111(.A(\A[208] ), .Y(new_n7114_));
  OAI21  g06112(.A0(\A[209] ), .A1(new_n7114_), .B0(\A[210] ), .Y(new_n7115_));
  INV    g06113(.A(\A[210] ), .Y(new_n7116_));
  NAND2  g06114(.A(new_n7098_), .B(new_n7116_), .Y(new_n7117_));
  OAI21  g06115(.A0(new_n7115_), .A1(new_n7113_), .B0(new_n7117_), .Y(new_n7118_));
  NAND4  g06116(.A(new_n7118_), .B(new_n7111_), .C(new_n7104_), .D(new_n7100_), .Y(new_n7119_));
  NAND2  g06117(.A(\A[200] ), .B(\A[199] ), .Y(new_n7120_));
  OAI21  g06118(.A0(new_n7063_), .A1(new_n7085_), .B0(new_n7120_), .Y(new_n7121_));
  NAND4  g06119(.A(new_n7121_), .B(new_n7074_), .C(new_n7070_), .D(new_n7064_), .Y(new_n7122_));
  NAND2  g06120(.A(\A[206] ), .B(new_n7107_), .Y(new_n7123_));
  AOI21  g06121(.A0(new_n7105_), .A1(\A[205] ), .B0(new_n7109_), .Y(new_n7124_));
  AOI22  g06122(.A0(new_n7124_), .A1(new_n7123_), .B0(new_n7102_), .B1(new_n7109_), .Y(new_n7125_));
  NAND2  g06123(.A(\A[209] ), .B(new_n7114_), .Y(new_n7126_));
  AOI21  g06124(.A0(new_n7112_), .A1(\A[208] ), .B0(new_n7116_), .Y(new_n7127_));
  AOI22  g06125(.A0(new_n7127_), .A1(new_n7126_), .B0(new_n7098_), .B1(new_n7116_), .Y(new_n7128_));
  XOR2   g06126(.A(new_n7128_), .B(new_n7125_), .Y(new_n7129_));
  NAND4  g06127(.A(new_n7129_), .B(new_n7122_), .C(new_n7119_), .D(new_n7096_), .Y(new_n7130_));
  XOR2   g06128(.A(new_n7104_), .B(new_n7100_), .Y(new_n7131_));
  NOR2   g06129(.A(new_n7128_), .B(new_n7125_), .Y(new_n7132_));
  AOI22  g06130(.A0(new_n7103_), .A1(new_n7101_), .B0(new_n7099_), .B1(new_n7097_), .Y(new_n7133_));
  AOI21  g06131(.A0(new_n7132_), .A1(new_n7131_), .B0(new_n7133_), .Y(new_n7134_));
  XOR2   g06132(.A(new_n7132_), .B(new_n7131_), .Y(new_n7135_));
  XOR2   g06133(.A(new_n7128_), .B(new_n7111_), .Y(new_n7136_));
  OAI21  g06134(.A0(new_n7136_), .A1(new_n7134_), .B0(new_n7135_), .Y(new_n7137_));
  XOR2   g06135(.A(new_n7137_), .B(new_n7130_), .Y(new_n7138_));
  NAND2  g06136(.A(new_n7118_), .B(new_n7111_), .Y(new_n7139_));
  XOR2   g06137(.A(new_n7139_), .B(new_n7131_), .Y(new_n7140_));
  NOR2   g06138(.A(new_n7105_), .B(new_n7107_), .Y(new_n7141_));
  AOI221 g06139(.A0(new_n7102_), .A1(\A[207] ), .C0(new_n7141_), .B0(new_n7099_), .B1(new_n7097_), .Y(new_n7142_));
  NOR2   g06140(.A(new_n7112_), .B(new_n7114_), .Y(new_n7143_));
  AOI221 g06141(.A0(new_n7103_), .A1(new_n7101_), .C0(new_n7143_), .B0(new_n7098_), .B1(\A[210] ), .Y(new_n7144_));
  OAI211 g06142(.A0(new_n7144_), .A1(new_n7142_), .B0(new_n7118_), .B1(new_n7111_), .Y(new_n7145_));
  NAND2  g06143(.A(new_n7104_), .B(new_n7100_), .Y(new_n7146_));
  AOI21  g06144(.A0(new_n7146_), .A1(new_n7145_), .B0(new_n7136_), .Y(new_n7147_));
  OAI21  g06145(.A0(new_n7147_), .A1(new_n7140_), .B0(new_n7130_), .Y(new_n7148_));
  NOR2   g06146(.A(new_n7136_), .B(new_n7084_), .Y(new_n7149_));
  OAI211 g06147(.A0(new_n7118_), .A1(new_n7111_), .B0(new_n7104_), .B1(new_n7100_), .Y(new_n7150_));
  NAND4  g06148(.A(new_n7150_), .B(new_n7149_), .C(new_n7122_), .D(new_n7135_), .Y(new_n7151_));
  AOI21  g06149(.A0(new_n7151_), .A1(new_n7148_), .B0(new_n7095_), .Y(new_n7152_));
  AOI21  g06150(.A0(new_n7138_), .A1(new_n7095_), .B0(new_n7152_), .Y(new_n7153_));
  INV    g06151(.A(\A[213] ), .Y(new_n7154_));
  INV    g06152(.A(\A[211] ), .Y(new_n7155_));
  NAND2  g06153(.A(\A[212] ), .B(new_n7155_), .Y(new_n7156_));
  INV    g06154(.A(\A[212] ), .Y(new_n7157_));
  AOI21  g06155(.A0(new_n7157_), .A1(\A[211] ), .B0(new_n7154_), .Y(new_n7158_));
  XOR2   g06156(.A(\A[212] ), .B(\A[211] ), .Y(new_n7159_));
  AOI22  g06157(.A0(new_n7159_), .A1(new_n7154_), .B0(new_n7158_), .B1(new_n7156_), .Y(new_n7160_));
  INV    g06158(.A(\A[216] ), .Y(new_n7161_));
  INV    g06159(.A(\A[214] ), .Y(new_n7162_));
  NAND2  g06160(.A(\A[215] ), .B(new_n7162_), .Y(new_n7163_));
  INV    g06161(.A(\A[215] ), .Y(new_n7164_));
  AOI21  g06162(.A0(new_n7164_), .A1(\A[214] ), .B0(new_n7161_), .Y(new_n7165_));
  XOR2   g06163(.A(\A[215] ), .B(\A[214] ), .Y(new_n7166_));
  AOI22  g06164(.A0(new_n7166_), .A1(new_n7161_), .B0(new_n7165_), .B1(new_n7163_), .Y(new_n7167_));
  NOR2   g06165(.A(new_n7167_), .B(new_n7160_), .Y(new_n7168_));
  XOR2   g06166(.A(\A[215] ), .B(new_n7162_), .Y(new_n7169_));
  NAND2  g06167(.A(\A[215] ), .B(\A[214] ), .Y(new_n7170_));
  OAI21  g06168(.A0(new_n7169_), .A1(new_n7161_), .B0(new_n7170_), .Y(new_n7171_));
  NOR2   g06169(.A(new_n7157_), .B(new_n7155_), .Y(new_n7172_));
  AOI21  g06170(.A0(new_n7159_), .A1(\A[213] ), .B0(new_n7172_), .Y(new_n7173_));
  XOR2   g06171(.A(new_n7173_), .B(new_n7171_), .Y(new_n7174_));
  XOR2   g06172(.A(new_n7174_), .B(new_n7168_), .Y(new_n7175_));
  XOR2   g06173(.A(new_n7167_), .B(new_n7160_), .Y(new_n7176_));
  NOR2   g06174(.A(new_n7157_), .B(\A[211] ), .Y(new_n7177_));
  OAI21  g06175(.A0(\A[212] ), .A1(new_n7155_), .B0(\A[213] ), .Y(new_n7178_));
  XOR2   g06176(.A(\A[212] ), .B(new_n7155_), .Y(new_n7179_));
  OAI22  g06177(.A0(new_n7179_), .A1(\A[213] ), .B0(new_n7178_), .B1(new_n7177_), .Y(new_n7180_));
  NOR2   g06178(.A(new_n7164_), .B(\A[214] ), .Y(new_n7181_));
  OAI21  g06179(.A0(\A[215] ), .A1(new_n7162_), .B0(\A[216] ), .Y(new_n7182_));
  OAI22  g06180(.A0(new_n7169_), .A1(\A[216] ), .B0(new_n7182_), .B1(new_n7181_), .Y(new_n7183_));
  NAND2  g06181(.A(new_n7183_), .B(new_n7180_), .Y(new_n7184_));
  NAND2  g06182(.A(\A[212] ), .B(\A[211] ), .Y(new_n7185_));
  OAI21  g06183(.A0(new_n7179_), .A1(new_n7154_), .B0(new_n7185_), .Y(new_n7186_));
  NAND2  g06184(.A(new_n7186_), .B(new_n7171_), .Y(new_n7187_));
  OAI21  g06185(.A0(new_n7174_), .A1(new_n7184_), .B0(new_n7187_), .Y(new_n7188_));
  AOI21  g06186(.A0(new_n7188_), .A1(new_n7176_), .B0(new_n7175_), .Y(new_n7189_));
  NAND2  g06187(.A(\A[221] ), .B(\A[220] ), .Y(new_n7190_));
  XOR2   g06188(.A(\A[221] ), .B(\A[220] ), .Y(new_n7191_));
  NAND2  g06189(.A(new_n7191_), .B(\A[222] ), .Y(new_n7192_));
  NAND2  g06190(.A(new_n7192_), .B(new_n7190_), .Y(new_n7193_));
  NAND2  g06191(.A(\A[218] ), .B(\A[217] ), .Y(new_n7194_));
  XOR2   g06192(.A(\A[218] ), .B(\A[217] ), .Y(new_n7195_));
  NAND2  g06193(.A(new_n7195_), .B(\A[219] ), .Y(new_n7196_));
  NAND2  g06194(.A(new_n7196_), .B(new_n7194_), .Y(new_n7197_));
  XOR2   g06195(.A(new_n7197_), .B(new_n7193_), .Y(new_n7198_));
  INV    g06196(.A(\A[219] ), .Y(new_n7199_));
  INV    g06197(.A(\A[217] ), .Y(new_n7200_));
  NAND2  g06198(.A(\A[218] ), .B(new_n7200_), .Y(new_n7201_));
  INV    g06199(.A(\A[218] ), .Y(new_n7202_));
  AOI21  g06200(.A0(new_n7202_), .A1(\A[217] ), .B0(new_n7199_), .Y(new_n7203_));
  AOI22  g06201(.A0(new_n7203_), .A1(new_n7201_), .B0(new_n7195_), .B1(new_n7199_), .Y(new_n7204_));
  INV    g06202(.A(\A[222] ), .Y(new_n7205_));
  INV    g06203(.A(\A[220] ), .Y(new_n7206_));
  NAND2  g06204(.A(\A[221] ), .B(new_n7206_), .Y(new_n7207_));
  INV    g06205(.A(\A[221] ), .Y(new_n7208_));
  AOI21  g06206(.A0(new_n7208_), .A1(\A[220] ), .B0(new_n7205_), .Y(new_n7209_));
  AOI22  g06207(.A0(new_n7209_), .A1(new_n7207_), .B0(new_n7191_), .B1(new_n7205_), .Y(new_n7210_));
  NOR2   g06208(.A(new_n7210_), .B(new_n7204_), .Y(new_n7211_));
  AOI22  g06209(.A0(new_n7196_), .A1(new_n7194_), .B0(new_n7192_), .B1(new_n7190_), .Y(new_n7212_));
  AOI21  g06210(.A0(new_n7211_), .A1(new_n7198_), .B0(new_n7212_), .Y(new_n7213_));
  XOR2   g06211(.A(new_n7211_), .B(new_n7198_), .Y(new_n7214_));
  NOR2   g06212(.A(new_n7202_), .B(\A[217] ), .Y(new_n7215_));
  OAI21  g06213(.A0(\A[218] ), .A1(new_n7200_), .B0(\A[219] ), .Y(new_n7216_));
  NAND2  g06214(.A(new_n7195_), .B(new_n7199_), .Y(new_n7217_));
  OAI21  g06215(.A0(new_n7216_), .A1(new_n7215_), .B0(new_n7217_), .Y(new_n7218_));
  XOR2   g06216(.A(new_n7210_), .B(new_n7218_), .Y(new_n7219_));
  NOR2   g06217(.A(new_n7208_), .B(\A[220] ), .Y(new_n7220_));
  OAI21  g06218(.A0(\A[221] ), .A1(new_n7206_), .B0(\A[222] ), .Y(new_n7221_));
  NAND2  g06219(.A(new_n7191_), .B(new_n7205_), .Y(new_n7222_));
  OAI21  g06220(.A0(new_n7221_), .A1(new_n7220_), .B0(new_n7222_), .Y(new_n7223_));
  NAND4  g06221(.A(new_n7223_), .B(new_n7218_), .C(new_n7197_), .D(new_n7193_), .Y(new_n7224_));
  NAND4  g06222(.A(new_n7186_), .B(new_n7171_), .C(new_n7183_), .D(new_n7180_), .Y(new_n7225_));
  XOR2   g06223(.A(new_n7210_), .B(new_n7204_), .Y(new_n7226_));
  NAND4  g06224(.A(new_n7226_), .B(new_n7225_), .C(new_n7224_), .D(new_n7176_), .Y(new_n7227_));
  OAI211 g06225(.A0(new_n7219_), .A1(new_n7213_), .B0(new_n7227_), .B1(new_n7214_), .Y(new_n7228_));
  NOR2   g06226(.A(new_n7202_), .B(new_n7200_), .Y(new_n7229_));
  AOI21  g06227(.A0(new_n7195_), .A1(\A[219] ), .B0(new_n7229_), .Y(new_n7230_));
  XOR2   g06228(.A(new_n7230_), .B(new_n7193_), .Y(new_n7231_));
  XOR2   g06229(.A(new_n7211_), .B(new_n7231_), .Y(new_n7232_));
  XOR2   g06230(.A(new_n7167_), .B(new_n7180_), .Y(new_n7233_));
  NOR2   g06231(.A(new_n7208_), .B(new_n7206_), .Y(new_n7234_));
  AOI21  g06232(.A0(new_n7191_), .A1(\A[222] ), .B0(new_n7234_), .Y(new_n7235_));
  NOR4   g06233(.A(new_n7210_), .B(new_n7204_), .C(new_n7230_), .D(new_n7235_), .Y(new_n7236_));
  NOR2   g06234(.A(new_n7164_), .B(new_n7162_), .Y(new_n7237_));
  AOI21  g06235(.A0(new_n7166_), .A1(\A[216] ), .B0(new_n7237_), .Y(new_n7238_));
  NOR4   g06236(.A(new_n7173_), .B(new_n7238_), .C(new_n7167_), .D(new_n7160_), .Y(new_n7239_));
  NOR4   g06237(.A(new_n7219_), .B(new_n7239_), .C(new_n7236_), .D(new_n7233_), .Y(new_n7240_));
  AOI221 g06238(.A0(new_n7195_), .A1(\A[219] ), .C0(new_n7229_), .B0(new_n7192_), .B1(new_n7190_), .Y(new_n7241_));
  AOI221 g06239(.A0(new_n7196_), .A1(new_n7194_), .C0(new_n7234_), .B0(new_n7191_), .B1(\A[222] ), .Y(new_n7242_));
  OAI211 g06240(.A0(new_n7242_), .A1(new_n7241_), .B0(new_n7223_), .B1(new_n7218_), .Y(new_n7243_));
  NAND2  g06241(.A(new_n7197_), .B(new_n7193_), .Y(new_n7244_));
  AOI21  g06242(.A0(new_n7244_), .A1(new_n7243_), .B0(new_n7219_), .Y(new_n7245_));
  OAI21  g06243(.A0(new_n7245_), .A1(new_n7232_), .B0(new_n7240_), .Y(new_n7246_));
  AOI21  g06244(.A0(new_n7246_), .A1(new_n7228_), .B0(new_n7189_), .Y(new_n7247_));
  XOR2   g06245(.A(new_n7174_), .B(new_n7184_), .Y(new_n7248_));
  XOR2   g06246(.A(new_n7173_), .B(new_n7238_), .Y(new_n7249_));
  NOR2   g06247(.A(new_n7173_), .B(new_n7238_), .Y(new_n7250_));
  AOI21  g06248(.A0(new_n7249_), .A1(new_n7168_), .B0(new_n7250_), .Y(new_n7251_));
  OAI21  g06249(.A0(new_n7251_), .A1(new_n7233_), .B0(new_n7248_), .Y(new_n7252_));
  OAI21  g06250(.A0(new_n7245_), .A1(new_n7232_), .B0(new_n7227_), .Y(new_n7253_));
  NOR2   g06251(.A(new_n7219_), .B(new_n7233_), .Y(new_n7254_));
  OAI211 g06252(.A0(new_n7223_), .A1(new_n7218_), .B0(new_n7197_), .B1(new_n7193_), .Y(new_n7255_));
  NAND4  g06253(.A(new_n7255_), .B(new_n7254_), .C(new_n7225_), .D(new_n7214_), .Y(new_n7256_));
  AOI21  g06254(.A0(new_n7256_), .A1(new_n7253_), .B0(new_n7252_), .Y(new_n7257_));
  NOR2   g06255(.A(new_n7219_), .B(new_n7236_), .Y(new_n7258_));
  XOR2   g06256(.A(new_n7167_), .B(new_n7160_), .Y(new_n7259_));
  XOR2   g06257(.A(new_n7259_), .B(new_n7258_), .Y(new_n7260_));
  NAND2  g06258(.A(new_n7129_), .B(new_n7119_), .Y(new_n7261_));
  XOR2   g06259(.A(new_n7083_), .B(new_n7064_), .Y(new_n7262_));
  XOR2   g06260(.A(new_n7262_), .B(new_n7261_), .Y(new_n7263_));
  NAND2  g06261(.A(new_n7263_), .B(new_n7260_), .Y(new_n7264_));
  NOR3   g06262(.A(new_n7264_), .B(new_n7257_), .C(new_n7247_), .Y(new_n7265_));
  OAI21  g06263(.A0(new_n7219_), .A1(new_n7213_), .B0(new_n7214_), .Y(new_n7266_));
  XOR2   g06264(.A(new_n7266_), .B(new_n7227_), .Y(new_n7267_));
  NAND2  g06265(.A(new_n7267_), .B(new_n7252_), .Y(new_n7268_));
  NAND2  g06266(.A(new_n7256_), .B(new_n7253_), .Y(new_n7269_));
  NAND2  g06267(.A(new_n7269_), .B(new_n7189_), .Y(new_n7270_));
  NAND2  g06268(.A(new_n7226_), .B(new_n7224_), .Y(new_n7271_));
  XOR2   g06269(.A(new_n7259_), .B(new_n7271_), .Y(new_n7272_));
  XOR2   g06270(.A(new_n7083_), .B(new_n7088_), .Y(new_n7273_));
  XOR2   g06271(.A(new_n7273_), .B(new_n7261_), .Y(new_n7274_));
  NOR2   g06272(.A(new_n7274_), .B(new_n7272_), .Y(new_n7275_));
  AOI21  g06273(.A0(new_n7270_), .A1(new_n7268_), .B0(new_n7275_), .Y(new_n7276_));
  OAI21  g06274(.A0(new_n7276_), .A1(new_n7265_), .B0(new_n7153_), .Y(new_n7277_));
  NAND2  g06275(.A(new_n7138_), .B(new_n7095_), .Y(new_n7278_));
  NAND2  g06276(.A(new_n7146_), .B(new_n7145_), .Y(new_n7279_));
  NAND3  g06277(.A(new_n7149_), .B(new_n7122_), .C(new_n7135_), .Y(new_n7280_));
  AOI211 g06278(.A0(new_n7135_), .A1(new_n7279_), .B(new_n7280_), .C(new_n7147_), .Y(new_n7281_));
  AOI21  g06279(.A0(new_n7137_), .A1(new_n7130_), .B0(new_n7281_), .Y(new_n7282_));
  OAI21  g06280(.A0(new_n7282_), .A1(new_n7095_), .B0(new_n7278_), .Y(new_n7283_));
  NAND2  g06281(.A(new_n7226_), .B(new_n7176_), .Y(new_n7284_));
  AOI211 g06282(.A0(new_n7210_), .A1(new_n7204_), .B(new_n7230_), .C(new_n7235_), .Y(new_n7285_));
  NOR4   g06283(.A(new_n7285_), .B(new_n7284_), .C(new_n7239_), .D(new_n7232_), .Y(new_n7286_));
  AOI21  g06284(.A0(new_n7266_), .A1(new_n7227_), .B0(new_n7286_), .Y(new_n7287_));
  OAI21  g06285(.A0(new_n7287_), .A1(new_n7252_), .B0(new_n7264_), .Y(new_n7288_));
  OAI21  g06286(.A0(new_n7257_), .A1(new_n7247_), .B0(new_n7275_), .Y(new_n7289_));
  OAI21  g06287(.A0(new_n7288_), .A1(new_n7247_), .B0(new_n7289_), .Y(new_n7290_));
  NAND2  g06288(.A(new_n7290_), .B(new_n7283_), .Y(new_n7291_));
  XOR2   g06289(.A(new_n7274_), .B(new_n7260_), .Y(new_n7292_));
  INV    g06290(.A(\A[195] ), .Y(new_n7293_));
  INV    g06291(.A(\A[194] ), .Y(new_n7294_));
  NAND2  g06292(.A(new_n7294_), .B(\A[193] ), .Y(new_n7295_));
  INV    g06293(.A(\A[193] ), .Y(new_n7296_));
  AOI21  g06294(.A0(\A[194] ), .A1(new_n7296_), .B0(new_n7293_), .Y(new_n7297_));
  XOR2   g06295(.A(\A[194] ), .B(\A[193] ), .Y(new_n7298_));
  AOI22  g06296(.A0(new_n7298_), .A1(new_n7293_), .B0(new_n7297_), .B1(new_n7295_), .Y(new_n7299_));
  INV    g06297(.A(\A[198] ), .Y(new_n7300_));
  INV    g06298(.A(\A[197] ), .Y(new_n7301_));
  NAND2  g06299(.A(new_n7301_), .B(\A[196] ), .Y(new_n7302_));
  INV    g06300(.A(\A[196] ), .Y(new_n7303_));
  AOI21  g06301(.A0(\A[197] ), .A1(new_n7303_), .B0(new_n7300_), .Y(new_n7304_));
  XOR2   g06302(.A(\A[197] ), .B(\A[196] ), .Y(new_n7305_));
  AOI22  g06303(.A0(new_n7305_), .A1(new_n7300_), .B0(new_n7304_), .B1(new_n7302_), .Y(new_n7306_));
  NOR2   g06304(.A(new_n7301_), .B(new_n7303_), .Y(new_n7307_));
  AOI21  g06305(.A0(new_n7305_), .A1(\A[198] ), .B0(new_n7307_), .Y(new_n7308_));
  NOR2   g06306(.A(new_n7294_), .B(new_n7296_), .Y(new_n7309_));
  AOI21  g06307(.A0(new_n7298_), .A1(\A[195] ), .B0(new_n7309_), .Y(new_n7310_));
  XOR2   g06308(.A(new_n7306_), .B(new_n7299_), .Y(new_n7311_));
  INV    g06309(.A(\A[189] ), .Y(new_n7312_));
  INV    g06310(.A(\A[188] ), .Y(new_n7313_));
  NAND2  g06311(.A(new_n7313_), .B(\A[187] ), .Y(new_n7314_));
  INV    g06312(.A(\A[187] ), .Y(new_n7315_));
  AOI21  g06313(.A0(\A[188] ), .A1(new_n7315_), .B0(new_n7312_), .Y(new_n7316_));
  XOR2   g06314(.A(\A[188] ), .B(\A[187] ), .Y(new_n7317_));
  AOI22  g06315(.A0(new_n7317_), .A1(new_n7312_), .B0(new_n7316_), .B1(new_n7314_), .Y(new_n7318_));
  INV    g06316(.A(\A[192] ), .Y(new_n7319_));
  INV    g06317(.A(\A[191] ), .Y(new_n7320_));
  NAND2  g06318(.A(new_n7320_), .B(\A[190] ), .Y(new_n7321_));
  INV    g06319(.A(\A[190] ), .Y(new_n7322_));
  AOI21  g06320(.A0(\A[191] ), .A1(new_n7322_), .B0(new_n7319_), .Y(new_n7323_));
  XOR2   g06321(.A(\A[191] ), .B(\A[190] ), .Y(new_n7324_));
  AOI22  g06322(.A0(new_n7324_), .A1(new_n7319_), .B0(new_n7323_), .B1(new_n7321_), .Y(new_n7325_));
  NOR2   g06323(.A(new_n7320_), .B(new_n7322_), .Y(new_n7326_));
  AOI21  g06324(.A0(new_n7324_), .A1(\A[192] ), .B0(new_n7326_), .Y(new_n7327_));
  NOR2   g06325(.A(new_n7313_), .B(new_n7315_), .Y(new_n7328_));
  AOI21  g06326(.A0(new_n7317_), .A1(\A[189] ), .B0(new_n7328_), .Y(new_n7329_));
  XOR2   g06327(.A(new_n7325_), .B(new_n7318_), .Y(new_n7330_));
  XOR2   g06328(.A(new_n7330_), .B(new_n7311_), .Y(new_n7331_));
  INV    g06329(.A(\A[181] ), .Y(new_n7332_));
  NOR2   g06330(.A(\A[182] ), .B(new_n7332_), .Y(new_n7333_));
  INV    g06331(.A(\A[182] ), .Y(new_n7334_));
  OAI21  g06332(.A0(new_n7334_), .A1(\A[181] ), .B0(\A[183] ), .Y(new_n7335_));
  INV    g06333(.A(\A[183] ), .Y(new_n7336_));
  XOR2   g06334(.A(\A[182] ), .B(\A[181] ), .Y(new_n7337_));
  NAND2  g06335(.A(new_n7337_), .B(new_n7336_), .Y(new_n7338_));
  OAI21  g06336(.A0(new_n7335_), .A1(new_n7333_), .B0(new_n7338_), .Y(new_n7339_));
  INV    g06337(.A(\A[186] ), .Y(new_n7340_));
  INV    g06338(.A(\A[185] ), .Y(new_n7341_));
  NAND2  g06339(.A(new_n7341_), .B(\A[184] ), .Y(new_n7342_));
  INV    g06340(.A(\A[184] ), .Y(new_n7343_));
  AOI21  g06341(.A0(\A[185] ), .A1(new_n7343_), .B0(new_n7340_), .Y(new_n7344_));
  XOR2   g06342(.A(\A[185] ), .B(\A[184] ), .Y(new_n7345_));
  AOI22  g06343(.A0(new_n7345_), .A1(new_n7340_), .B0(new_n7344_), .B1(new_n7342_), .Y(new_n7346_));
  NOR2   g06344(.A(new_n7341_), .B(new_n7343_), .Y(new_n7347_));
  AOI21  g06345(.A0(new_n7345_), .A1(\A[186] ), .B0(new_n7347_), .Y(new_n7348_));
  NOR2   g06346(.A(new_n7334_), .B(new_n7332_), .Y(new_n7349_));
  AOI21  g06347(.A0(new_n7337_), .A1(\A[183] ), .B0(new_n7349_), .Y(new_n7350_));
  XOR2   g06348(.A(new_n7346_), .B(new_n7339_), .Y(new_n7351_));
  INV    g06349(.A(\A[177] ), .Y(new_n7352_));
  INV    g06350(.A(\A[176] ), .Y(new_n7353_));
  NAND2  g06351(.A(new_n7353_), .B(\A[175] ), .Y(new_n7354_));
  INV    g06352(.A(\A[175] ), .Y(new_n7355_));
  AOI21  g06353(.A0(\A[176] ), .A1(new_n7355_), .B0(new_n7352_), .Y(new_n7356_));
  XOR2   g06354(.A(\A[176] ), .B(\A[175] ), .Y(new_n7357_));
  AOI22  g06355(.A0(new_n7357_), .A1(new_n7352_), .B0(new_n7356_), .B1(new_n7354_), .Y(new_n7358_));
  INV    g06356(.A(\A[180] ), .Y(new_n7359_));
  INV    g06357(.A(\A[179] ), .Y(new_n7360_));
  NAND2  g06358(.A(new_n7360_), .B(\A[178] ), .Y(new_n7361_));
  INV    g06359(.A(\A[178] ), .Y(new_n7362_));
  AOI21  g06360(.A0(\A[179] ), .A1(new_n7362_), .B0(new_n7359_), .Y(new_n7363_));
  XOR2   g06361(.A(\A[179] ), .B(\A[178] ), .Y(new_n7364_));
  AOI22  g06362(.A0(new_n7364_), .A1(new_n7359_), .B0(new_n7363_), .B1(new_n7361_), .Y(new_n7365_));
  NOR2   g06363(.A(new_n7360_), .B(new_n7362_), .Y(new_n7366_));
  AOI21  g06364(.A0(new_n7364_), .A1(\A[180] ), .B0(new_n7366_), .Y(new_n7367_));
  NOR2   g06365(.A(new_n7353_), .B(new_n7355_), .Y(new_n7368_));
  AOI21  g06366(.A0(new_n7357_), .A1(\A[177] ), .B0(new_n7368_), .Y(new_n7369_));
  XOR2   g06367(.A(new_n7365_), .B(new_n7358_), .Y(new_n7370_));
  XOR2   g06368(.A(new_n7370_), .B(new_n7351_), .Y(new_n7371_));
  XOR2   g06369(.A(new_n7371_), .B(new_n7331_), .Y(new_n7372_));
  NOR2   g06370(.A(new_n7372_), .B(new_n7292_), .Y(new_n7373_));
  NAND3  g06371(.A(new_n7373_), .B(new_n7291_), .C(new_n7277_), .Y(new_n7374_));
  NAND3  g06372(.A(new_n7275_), .B(new_n7270_), .C(new_n7268_), .Y(new_n7375_));
  OAI21  g06373(.A0(new_n7257_), .A1(new_n7247_), .B0(new_n7264_), .Y(new_n7376_));
  AOI21  g06374(.A0(new_n7376_), .A1(new_n7375_), .B0(new_n7283_), .Y(new_n7377_));
  NAND3  g06375(.A(new_n7264_), .B(new_n7270_), .C(new_n7268_), .Y(new_n7378_));
  AOI21  g06376(.A0(new_n7289_), .A1(new_n7378_), .B0(new_n7153_), .Y(new_n7379_));
  INV    g06377(.A(new_n7373_), .Y(new_n7380_));
  OAI21  g06378(.A0(new_n7379_), .A1(new_n7377_), .B0(new_n7380_), .Y(new_n7381_));
  XOR2   g06379(.A(new_n7325_), .B(new_n7318_), .Y(new_n7382_));
  XOR2   g06380(.A(\A[191] ), .B(new_n7322_), .Y(new_n7383_));
  NAND2  g06381(.A(\A[191] ), .B(\A[190] ), .Y(new_n7384_));
  OAI21  g06382(.A0(new_n7383_), .A1(new_n7319_), .B0(new_n7384_), .Y(new_n7385_));
  XOR2   g06383(.A(new_n7329_), .B(new_n7385_), .Y(new_n7386_));
  NOR2   g06384(.A(\A[188] ), .B(new_n7315_), .Y(new_n7387_));
  OAI21  g06385(.A0(new_n7313_), .A1(\A[187] ), .B0(\A[189] ), .Y(new_n7388_));
  XOR2   g06386(.A(\A[188] ), .B(new_n7315_), .Y(new_n7389_));
  OAI22  g06387(.A0(new_n7389_), .A1(\A[189] ), .B0(new_n7388_), .B1(new_n7387_), .Y(new_n7390_));
  NOR2   g06388(.A(\A[191] ), .B(new_n7322_), .Y(new_n7391_));
  OAI21  g06389(.A0(new_n7320_), .A1(\A[190] ), .B0(\A[192] ), .Y(new_n7392_));
  OAI22  g06390(.A0(new_n7383_), .A1(\A[192] ), .B0(new_n7392_), .B1(new_n7391_), .Y(new_n7393_));
  NAND2  g06391(.A(new_n7393_), .B(new_n7390_), .Y(new_n7394_));
  NAND2  g06392(.A(\A[188] ), .B(\A[187] ), .Y(new_n7395_));
  OAI21  g06393(.A0(new_n7389_), .A1(new_n7312_), .B0(new_n7395_), .Y(new_n7396_));
  NAND2  g06394(.A(new_n7396_), .B(new_n7385_), .Y(new_n7397_));
  OAI21  g06395(.A0(new_n7394_), .A1(new_n7386_), .B0(new_n7397_), .Y(new_n7398_));
  NOR2   g06396(.A(new_n7325_), .B(new_n7318_), .Y(new_n7399_));
  XOR2   g06397(.A(new_n7399_), .B(new_n7386_), .Y(new_n7400_));
  AOI21  g06398(.A0(new_n7398_), .A1(new_n7382_), .B0(new_n7400_), .Y(new_n7401_));
  NOR2   g06399(.A(\A[194] ), .B(new_n7296_), .Y(new_n7402_));
  OAI21  g06400(.A0(new_n7294_), .A1(\A[193] ), .B0(\A[195] ), .Y(new_n7403_));
  NAND2  g06401(.A(new_n7298_), .B(new_n7293_), .Y(new_n7404_));
  OAI21  g06402(.A0(new_n7403_), .A1(new_n7402_), .B0(new_n7404_), .Y(new_n7405_));
  XOR2   g06403(.A(new_n7306_), .B(new_n7405_), .Y(new_n7406_));
  XOR2   g06404(.A(new_n7310_), .B(new_n7308_), .Y(new_n7407_));
  NOR2   g06405(.A(new_n7306_), .B(new_n7299_), .Y(new_n7408_));
  NAND2  g06406(.A(\A[197] ), .B(\A[196] ), .Y(new_n7409_));
  NAND2  g06407(.A(new_n7305_), .B(\A[198] ), .Y(new_n7410_));
  NAND2  g06408(.A(\A[194] ), .B(\A[193] ), .Y(new_n7411_));
  NAND2  g06409(.A(new_n7298_), .B(\A[195] ), .Y(new_n7412_));
  AOI22  g06410(.A0(new_n7412_), .A1(new_n7411_), .B0(new_n7410_), .B1(new_n7409_), .Y(new_n7413_));
  AOI21  g06411(.A0(new_n7408_), .A1(new_n7407_), .B0(new_n7413_), .Y(new_n7414_));
  XOR2   g06412(.A(new_n7408_), .B(new_n7407_), .Y(new_n7415_));
  XOR2   g06413(.A(new_n7306_), .B(new_n7299_), .Y(new_n7416_));
  NOR2   g06414(.A(\A[197] ), .B(new_n7303_), .Y(new_n7417_));
  OAI21  g06415(.A0(new_n7301_), .A1(\A[196] ), .B0(\A[198] ), .Y(new_n7418_));
  NAND2  g06416(.A(new_n7305_), .B(new_n7300_), .Y(new_n7419_));
  OAI21  g06417(.A0(new_n7418_), .A1(new_n7417_), .B0(new_n7419_), .Y(new_n7420_));
  NAND2  g06418(.A(new_n7410_), .B(new_n7409_), .Y(new_n7421_));
  NAND2  g06419(.A(new_n7412_), .B(new_n7411_), .Y(new_n7422_));
  NAND4  g06420(.A(new_n7422_), .B(new_n7421_), .C(new_n7420_), .D(new_n7405_), .Y(new_n7423_));
  NAND4  g06421(.A(new_n7396_), .B(new_n7385_), .C(new_n7393_), .D(new_n7390_), .Y(new_n7424_));
  NAND4  g06422(.A(new_n7424_), .B(new_n7382_), .C(new_n7423_), .D(new_n7416_), .Y(new_n7425_));
  OAI211 g06423(.A0(new_n7414_), .A1(new_n7406_), .B0(new_n7425_), .B1(new_n7415_), .Y(new_n7426_));
  XOR2   g06424(.A(new_n7310_), .B(new_n7421_), .Y(new_n7427_));
  XOR2   g06425(.A(new_n7408_), .B(new_n7427_), .Y(new_n7428_));
  NOR4   g06426(.A(new_n7310_), .B(new_n7308_), .C(new_n7306_), .D(new_n7299_), .Y(new_n7429_));
  XOR2   g06427(.A(new_n7325_), .B(new_n7390_), .Y(new_n7430_));
  NOR4   g06428(.A(new_n7329_), .B(new_n7327_), .C(new_n7325_), .D(new_n7318_), .Y(new_n7431_));
  NOR4   g06429(.A(new_n7431_), .B(new_n7430_), .C(new_n7429_), .D(new_n7406_), .Y(new_n7432_));
  AOI221 g06430(.A0(new_n7410_), .A1(new_n7409_), .C0(new_n7309_), .B0(new_n7298_), .B1(\A[195] ), .Y(new_n7433_));
  AOI221 g06431(.A0(new_n7412_), .A1(new_n7411_), .C0(new_n7307_), .B0(new_n7305_), .B1(\A[198] ), .Y(new_n7434_));
  OAI211 g06432(.A0(new_n7434_), .A1(new_n7433_), .B0(new_n7420_), .B1(new_n7405_), .Y(new_n7435_));
  NAND2  g06433(.A(new_n7422_), .B(new_n7421_), .Y(new_n7436_));
  AOI21  g06434(.A0(new_n7436_), .A1(new_n7435_), .B0(new_n7406_), .Y(new_n7437_));
  OAI21  g06435(.A0(new_n7437_), .A1(new_n7428_), .B0(new_n7432_), .Y(new_n7438_));
  AOI21  g06436(.A0(new_n7438_), .A1(new_n7426_), .B0(new_n7401_), .Y(new_n7439_));
  OAI21  g06437(.A0(new_n7437_), .A1(new_n7428_), .B0(new_n7425_), .Y(new_n7440_));
  NAND4  g06438(.A(new_n7382_), .B(new_n7415_), .C(new_n7414_), .D(new_n7416_), .Y(new_n7441_));
  OAI21  g06439(.A0(new_n7414_), .A1(new_n7406_), .B0(new_n7424_), .Y(new_n7442_));
  OAI21  g06440(.A0(new_n7442_), .A1(new_n7441_), .B0(new_n7440_), .Y(new_n7443_));
  NAND2  g06441(.A(new_n7334_), .B(\A[181] ), .Y(new_n7444_));
  AOI21  g06442(.A0(\A[182] ), .A1(new_n7332_), .B0(new_n7336_), .Y(new_n7445_));
  AOI22  g06443(.A0(new_n7337_), .A1(new_n7336_), .B0(new_n7445_), .B1(new_n7444_), .Y(new_n7446_));
  XOR2   g06444(.A(new_n7346_), .B(new_n7446_), .Y(new_n7447_));
  XOR2   g06445(.A(new_n7370_), .B(new_n7447_), .Y(new_n7448_));
  NAND2  g06446(.A(new_n7448_), .B(new_n7331_), .Y(new_n7449_));
  AOI211 g06447(.A0(new_n7443_), .A1(new_n7401_), .B(new_n7449_), .C(new_n7439_), .Y(new_n7450_));
  XOR2   g06448(.A(new_n7306_), .B(new_n7405_), .Y(new_n7451_));
  XOR2   g06449(.A(new_n7330_), .B(new_n7451_), .Y(new_n7452_));
  NOR2   g06450(.A(new_n7371_), .B(new_n7452_), .Y(new_n7453_));
  AOI21  g06451(.A0(new_n7443_), .A1(new_n7401_), .B0(new_n7439_), .Y(new_n7454_));
  NOR2   g06452(.A(new_n7454_), .B(new_n7453_), .Y(new_n7455_));
  XOR2   g06453(.A(new_n7365_), .B(new_n7358_), .Y(new_n7456_));
  XOR2   g06454(.A(\A[179] ), .B(new_n7362_), .Y(new_n7457_));
  NAND2  g06455(.A(\A[179] ), .B(\A[178] ), .Y(new_n7458_));
  OAI21  g06456(.A0(new_n7457_), .A1(new_n7359_), .B0(new_n7458_), .Y(new_n7459_));
  XOR2   g06457(.A(new_n7369_), .B(new_n7459_), .Y(new_n7460_));
  NOR2   g06458(.A(\A[176] ), .B(new_n7355_), .Y(new_n7461_));
  OAI21  g06459(.A0(new_n7353_), .A1(\A[175] ), .B0(\A[177] ), .Y(new_n7462_));
  XOR2   g06460(.A(\A[176] ), .B(new_n7355_), .Y(new_n7463_));
  OAI22  g06461(.A0(new_n7463_), .A1(\A[177] ), .B0(new_n7462_), .B1(new_n7461_), .Y(new_n7464_));
  NOR2   g06462(.A(\A[179] ), .B(new_n7362_), .Y(new_n7465_));
  OAI21  g06463(.A0(new_n7360_), .A1(\A[178] ), .B0(\A[180] ), .Y(new_n7466_));
  OAI22  g06464(.A0(new_n7457_), .A1(\A[180] ), .B0(new_n7466_), .B1(new_n7465_), .Y(new_n7467_));
  NAND2  g06465(.A(new_n7467_), .B(new_n7464_), .Y(new_n7468_));
  NAND2  g06466(.A(\A[176] ), .B(\A[175] ), .Y(new_n7469_));
  OAI21  g06467(.A0(new_n7463_), .A1(new_n7352_), .B0(new_n7469_), .Y(new_n7470_));
  NAND2  g06468(.A(new_n7470_), .B(new_n7459_), .Y(new_n7471_));
  OAI21  g06469(.A0(new_n7468_), .A1(new_n7460_), .B0(new_n7471_), .Y(new_n7472_));
  NOR2   g06470(.A(new_n7365_), .B(new_n7358_), .Y(new_n7473_));
  XOR2   g06471(.A(new_n7473_), .B(new_n7460_), .Y(new_n7474_));
  AOI21  g06472(.A0(new_n7472_), .A1(new_n7456_), .B0(new_n7474_), .Y(new_n7475_));
  XOR2   g06473(.A(new_n7346_), .B(new_n7339_), .Y(new_n7476_));
  XOR2   g06474(.A(new_n7350_), .B(new_n7348_), .Y(new_n7477_));
  NOR2   g06475(.A(new_n7346_), .B(new_n7446_), .Y(new_n7478_));
  NAND2  g06476(.A(\A[185] ), .B(\A[184] ), .Y(new_n7479_));
  NAND2  g06477(.A(new_n7345_), .B(\A[186] ), .Y(new_n7480_));
  NAND2  g06478(.A(\A[182] ), .B(\A[181] ), .Y(new_n7481_));
  NAND2  g06479(.A(new_n7337_), .B(\A[183] ), .Y(new_n7482_));
  AOI22  g06480(.A0(new_n7482_), .A1(new_n7481_), .B0(new_n7480_), .B1(new_n7479_), .Y(new_n7483_));
  AOI21  g06481(.A0(new_n7478_), .A1(new_n7477_), .B0(new_n7483_), .Y(new_n7484_));
  XOR2   g06482(.A(new_n7478_), .B(new_n7477_), .Y(new_n7485_));
  XOR2   g06483(.A(new_n7346_), .B(new_n7446_), .Y(new_n7486_));
  NOR2   g06484(.A(\A[185] ), .B(new_n7343_), .Y(new_n7487_));
  OAI21  g06485(.A0(new_n7341_), .A1(\A[184] ), .B0(\A[186] ), .Y(new_n7488_));
  NAND2  g06486(.A(new_n7345_), .B(new_n7340_), .Y(new_n7489_));
  OAI21  g06487(.A0(new_n7488_), .A1(new_n7487_), .B0(new_n7489_), .Y(new_n7490_));
  NAND2  g06488(.A(new_n7480_), .B(new_n7479_), .Y(new_n7491_));
  NAND2  g06489(.A(new_n7482_), .B(new_n7481_), .Y(new_n7492_));
  NAND4  g06490(.A(new_n7492_), .B(new_n7491_), .C(new_n7490_), .D(new_n7339_), .Y(new_n7493_));
  NAND4  g06491(.A(new_n7470_), .B(new_n7459_), .C(new_n7467_), .D(new_n7464_), .Y(new_n7494_));
  NAND4  g06492(.A(new_n7494_), .B(new_n7456_), .C(new_n7493_), .D(new_n7486_), .Y(new_n7495_));
  OAI211 g06493(.A0(new_n7484_), .A1(new_n7476_), .B0(new_n7495_), .B1(new_n7485_), .Y(new_n7496_));
  XOR2   g06494(.A(new_n7350_), .B(new_n7491_), .Y(new_n7497_));
  XOR2   g06495(.A(new_n7478_), .B(new_n7497_), .Y(new_n7498_));
  NOR4   g06496(.A(new_n7350_), .B(new_n7348_), .C(new_n7346_), .D(new_n7446_), .Y(new_n7499_));
  XOR2   g06497(.A(new_n7365_), .B(new_n7464_), .Y(new_n7500_));
  NOR4   g06498(.A(new_n7369_), .B(new_n7367_), .C(new_n7365_), .D(new_n7358_), .Y(new_n7501_));
  NOR4   g06499(.A(new_n7501_), .B(new_n7500_), .C(new_n7499_), .D(new_n7476_), .Y(new_n7502_));
  AOI221 g06500(.A0(new_n7480_), .A1(new_n7479_), .C0(new_n7349_), .B0(new_n7337_), .B1(\A[183] ), .Y(new_n7503_));
  AOI221 g06501(.A0(new_n7482_), .A1(new_n7481_), .C0(new_n7347_), .B0(new_n7345_), .B1(\A[186] ), .Y(new_n7504_));
  OAI211 g06502(.A0(new_n7504_), .A1(new_n7503_), .B0(new_n7490_), .B1(new_n7339_), .Y(new_n7505_));
  NAND2  g06503(.A(new_n7492_), .B(new_n7491_), .Y(new_n7506_));
  AOI21  g06504(.A0(new_n7506_), .A1(new_n7505_), .B0(new_n7476_), .Y(new_n7507_));
  OAI21  g06505(.A0(new_n7507_), .A1(new_n7498_), .B0(new_n7502_), .Y(new_n7508_));
  AOI21  g06506(.A0(new_n7508_), .A1(new_n7496_), .B0(new_n7475_), .Y(new_n7509_));
  NOR2   g06507(.A(new_n7507_), .B(new_n7498_), .Y(new_n7510_));
  NAND4  g06508(.A(new_n7456_), .B(new_n7485_), .C(new_n7484_), .D(new_n7486_), .Y(new_n7511_));
  OAI21  g06509(.A0(new_n7484_), .A1(new_n7476_), .B0(new_n7494_), .Y(new_n7512_));
  OAI22  g06510(.A0(new_n7512_), .A1(new_n7511_), .B0(new_n7510_), .B1(new_n7502_), .Y(new_n7513_));
  AOI21  g06511(.A0(new_n7513_), .A1(new_n7475_), .B0(new_n7509_), .Y(new_n7514_));
  OAI21  g06512(.A0(new_n7455_), .A1(new_n7450_), .B0(new_n7514_), .Y(new_n7515_));
  XOR2   g06513(.A(new_n7510_), .B(new_n7495_), .Y(new_n7516_));
  NAND2  g06514(.A(new_n7513_), .B(new_n7475_), .Y(new_n7517_));
  OAI21  g06515(.A0(new_n7516_), .A1(new_n7475_), .B0(new_n7517_), .Y(new_n7518_));
  AOI211 g06516(.A0(new_n7443_), .A1(new_n7401_), .B(new_n7453_), .C(new_n7439_), .Y(new_n7519_));
  NOR2   g06517(.A(new_n7454_), .B(new_n7449_), .Y(new_n7520_));
  OAI21  g06518(.A0(new_n7520_), .A1(new_n7519_), .B0(new_n7518_), .Y(new_n7521_));
  NAND2  g06519(.A(new_n7521_), .B(new_n7515_), .Y(new_n7522_));
  AOI21  g06520(.A0(new_n7381_), .A1(new_n7374_), .B0(new_n7522_), .Y(new_n7523_));
  XOR2   g06521(.A(new_n7329_), .B(new_n7327_), .Y(new_n7524_));
  NOR2   g06522(.A(new_n7329_), .B(new_n7327_), .Y(new_n7525_));
  AOI21  g06523(.A0(new_n7399_), .A1(new_n7524_), .B0(new_n7525_), .Y(new_n7526_));
  XOR2   g06524(.A(new_n7399_), .B(new_n7524_), .Y(new_n7527_));
  OAI21  g06525(.A0(new_n7526_), .A1(new_n7430_), .B0(new_n7527_), .Y(new_n7528_));
  OAI21  g06526(.A0(new_n7414_), .A1(new_n7406_), .B0(new_n7415_), .Y(new_n7529_));
  XOR2   g06527(.A(new_n7529_), .B(new_n7425_), .Y(new_n7530_));
  NAND2  g06528(.A(new_n7530_), .B(new_n7528_), .Y(new_n7531_));
  NAND2  g06529(.A(new_n7443_), .B(new_n7401_), .Y(new_n7532_));
  NAND3  g06530(.A(new_n7453_), .B(new_n7532_), .C(new_n7531_), .Y(new_n7533_));
  NAND2  g06531(.A(new_n7436_), .B(new_n7435_), .Y(new_n7534_));
  NOR4   g06532(.A(new_n7430_), .B(new_n7428_), .C(new_n7534_), .D(new_n7406_), .Y(new_n7535_));
  OAI211 g06533(.A0(new_n7414_), .A1(new_n7406_), .B0(new_n7535_), .B1(new_n7424_), .Y(new_n7536_));
  AOI21  g06534(.A0(new_n7536_), .A1(new_n7440_), .B0(new_n7528_), .Y(new_n7537_));
  OAI21  g06535(.A0(new_n7537_), .A1(new_n7439_), .B0(new_n7449_), .Y(new_n7538_));
  AOI21  g06536(.A0(new_n7538_), .A1(new_n7533_), .B0(new_n7518_), .Y(new_n7539_));
  NAND3  g06537(.A(new_n7449_), .B(new_n7532_), .C(new_n7531_), .Y(new_n7540_));
  OAI21  g06538(.A0(new_n7454_), .A1(new_n7449_), .B0(new_n7540_), .Y(new_n7541_));
  AOI21  g06539(.A0(new_n7541_), .A1(new_n7518_), .B0(new_n7539_), .Y(new_n7542_));
  AOI21  g06540(.A0(new_n7290_), .A1(new_n7283_), .B0(new_n7373_), .Y(new_n7543_));
  NAND2  g06541(.A(new_n7543_), .B(new_n7277_), .Y(new_n7544_));
  OAI21  g06542(.A0(new_n7379_), .A1(new_n7377_), .B0(new_n7373_), .Y(new_n7545_));
  AOI21  g06543(.A0(new_n7545_), .A1(new_n7544_), .B0(new_n7542_), .Y(new_n7546_));
  NOR2   g06544(.A(new_n7546_), .B(new_n7523_), .Y(new_n7547_));
  INV    g06545(.A(\A[237] ), .Y(new_n7548_));
  INV    g06546(.A(\A[235] ), .Y(new_n7549_));
  NAND2  g06547(.A(\A[236] ), .B(new_n7549_), .Y(new_n7550_));
  INV    g06548(.A(\A[236] ), .Y(new_n7551_));
  AOI21  g06549(.A0(new_n7551_), .A1(\A[235] ), .B0(new_n7548_), .Y(new_n7552_));
  XOR2   g06550(.A(\A[236] ), .B(\A[235] ), .Y(new_n7553_));
  AOI22  g06551(.A0(new_n7553_), .A1(new_n7548_), .B0(new_n7552_), .B1(new_n7550_), .Y(new_n7554_));
  INV    g06552(.A(\A[240] ), .Y(new_n7555_));
  INV    g06553(.A(\A[238] ), .Y(new_n7556_));
  NAND2  g06554(.A(\A[239] ), .B(new_n7556_), .Y(new_n7557_));
  INV    g06555(.A(\A[239] ), .Y(new_n7558_));
  AOI21  g06556(.A0(new_n7558_), .A1(\A[238] ), .B0(new_n7555_), .Y(new_n7559_));
  XOR2   g06557(.A(\A[239] ), .B(\A[238] ), .Y(new_n7560_));
  AOI22  g06558(.A0(new_n7560_), .A1(new_n7555_), .B0(new_n7559_), .B1(new_n7557_), .Y(new_n7561_));
  NOR2   g06559(.A(new_n7561_), .B(new_n7554_), .Y(new_n7562_));
  XOR2   g06560(.A(\A[239] ), .B(new_n7556_), .Y(new_n7563_));
  NAND2  g06561(.A(\A[239] ), .B(\A[238] ), .Y(new_n7564_));
  OAI21  g06562(.A0(new_n7563_), .A1(new_n7555_), .B0(new_n7564_), .Y(new_n7565_));
  NOR2   g06563(.A(new_n7551_), .B(new_n7549_), .Y(new_n7566_));
  AOI21  g06564(.A0(new_n7553_), .A1(\A[237] ), .B0(new_n7566_), .Y(new_n7567_));
  XOR2   g06565(.A(new_n7567_), .B(new_n7565_), .Y(new_n7568_));
  XOR2   g06566(.A(new_n7568_), .B(new_n7562_), .Y(new_n7569_));
  XOR2   g06567(.A(new_n7561_), .B(new_n7554_), .Y(new_n7570_));
  NOR2   g06568(.A(new_n7551_), .B(\A[235] ), .Y(new_n7571_));
  OAI21  g06569(.A0(\A[236] ), .A1(new_n7549_), .B0(\A[237] ), .Y(new_n7572_));
  XOR2   g06570(.A(\A[236] ), .B(new_n7549_), .Y(new_n7573_));
  OAI22  g06571(.A0(new_n7573_), .A1(\A[237] ), .B0(new_n7572_), .B1(new_n7571_), .Y(new_n7574_));
  NOR2   g06572(.A(new_n7558_), .B(\A[238] ), .Y(new_n7575_));
  OAI21  g06573(.A0(\A[239] ), .A1(new_n7556_), .B0(\A[240] ), .Y(new_n7576_));
  OAI22  g06574(.A0(new_n7563_), .A1(\A[240] ), .B0(new_n7576_), .B1(new_n7575_), .Y(new_n7577_));
  NAND2  g06575(.A(new_n7577_), .B(new_n7574_), .Y(new_n7578_));
  NAND2  g06576(.A(\A[236] ), .B(\A[235] ), .Y(new_n7579_));
  OAI21  g06577(.A0(new_n7573_), .A1(new_n7548_), .B0(new_n7579_), .Y(new_n7580_));
  NAND2  g06578(.A(new_n7580_), .B(new_n7565_), .Y(new_n7581_));
  OAI21  g06579(.A0(new_n7568_), .A1(new_n7578_), .B0(new_n7581_), .Y(new_n7582_));
  AOI21  g06580(.A0(new_n7582_), .A1(new_n7570_), .B0(new_n7569_), .Y(new_n7583_));
  NAND2  g06581(.A(\A[245] ), .B(\A[244] ), .Y(new_n7584_));
  XOR2   g06582(.A(\A[245] ), .B(\A[244] ), .Y(new_n7585_));
  NAND2  g06583(.A(new_n7585_), .B(\A[246] ), .Y(new_n7586_));
  NAND2  g06584(.A(new_n7586_), .B(new_n7584_), .Y(new_n7587_));
  NAND2  g06585(.A(\A[242] ), .B(\A[241] ), .Y(new_n7588_));
  XOR2   g06586(.A(\A[242] ), .B(\A[241] ), .Y(new_n7589_));
  NAND2  g06587(.A(new_n7589_), .B(\A[243] ), .Y(new_n7590_));
  NAND2  g06588(.A(new_n7590_), .B(new_n7588_), .Y(new_n7591_));
  XOR2   g06589(.A(new_n7591_), .B(new_n7587_), .Y(new_n7592_));
  INV    g06590(.A(\A[243] ), .Y(new_n7593_));
  INV    g06591(.A(\A[241] ), .Y(new_n7594_));
  NAND2  g06592(.A(\A[242] ), .B(new_n7594_), .Y(new_n7595_));
  INV    g06593(.A(\A[242] ), .Y(new_n7596_));
  AOI21  g06594(.A0(new_n7596_), .A1(\A[241] ), .B0(new_n7593_), .Y(new_n7597_));
  AOI22  g06595(.A0(new_n7597_), .A1(new_n7595_), .B0(new_n7589_), .B1(new_n7593_), .Y(new_n7598_));
  INV    g06596(.A(\A[246] ), .Y(new_n7599_));
  INV    g06597(.A(\A[244] ), .Y(new_n7600_));
  NAND2  g06598(.A(\A[245] ), .B(new_n7600_), .Y(new_n7601_));
  INV    g06599(.A(\A[245] ), .Y(new_n7602_));
  AOI21  g06600(.A0(new_n7602_), .A1(\A[244] ), .B0(new_n7599_), .Y(new_n7603_));
  AOI22  g06601(.A0(new_n7603_), .A1(new_n7601_), .B0(new_n7585_), .B1(new_n7599_), .Y(new_n7604_));
  NOR2   g06602(.A(new_n7604_), .B(new_n7598_), .Y(new_n7605_));
  AOI22  g06603(.A0(new_n7590_), .A1(new_n7588_), .B0(new_n7586_), .B1(new_n7584_), .Y(new_n7606_));
  AOI21  g06604(.A0(new_n7605_), .A1(new_n7592_), .B0(new_n7606_), .Y(new_n7607_));
  XOR2   g06605(.A(new_n7605_), .B(new_n7592_), .Y(new_n7608_));
  NOR2   g06606(.A(new_n7596_), .B(\A[241] ), .Y(new_n7609_));
  OAI21  g06607(.A0(\A[242] ), .A1(new_n7594_), .B0(\A[243] ), .Y(new_n7610_));
  NAND2  g06608(.A(new_n7589_), .B(new_n7593_), .Y(new_n7611_));
  OAI21  g06609(.A0(new_n7610_), .A1(new_n7609_), .B0(new_n7611_), .Y(new_n7612_));
  XOR2   g06610(.A(new_n7604_), .B(new_n7612_), .Y(new_n7613_));
  NOR2   g06611(.A(new_n7602_), .B(\A[244] ), .Y(new_n7614_));
  OAI21  g06612(.A0(\A[245] ), .A1(new_n7600_), .B0(\A[246] ), .Y(new_n7615_));
  NAND2  g06613(.A(new_n7585_), .B(new_n7599_), .Y(new_n7616_));
  OAI21  g06614(.A0(new_n7615_), .A1(new_n7614_), .B0(new_n7616_), .Y(new_n7617_));
  NAND4  g06615(.A(new_n7617_), .B(new_n7612_), .C(new_n7591_), .D(new_n7587_), .Y(new_n7618_));
  NAND4  g06616(.A(new_n7580_), .B(new_n7565_), .C(new_n7577_), .D(new_n7574_), .Y(new_n7619_));
  XOR2   g06617(.A(new_n7604_), .B(new_n7598_), .Y(new_n7620_));
  NAND4  g06618(.A(new_n7620_), .B(new_n7619_), .C(new_n7618_), .D(new_n7570_), .Y(new_n7621_));
  OAI211 g06619(.A0(new_n7613_), .A1(new_n7607_), .B0(new_n7621_), .B1(new_n7608_), .Y(new_n7622_));
  NOR2   g06620(.A(new_n7596_), .B(new_n7594_), .Y(new_n7623_));
  AOI21  g06621(.A0(new_n7589_), .A1(\A[243] ), .B0(new_n7623_), .Y(new_n7624_));
  XOR2   g06622(.A(new_n7624_), .B(new_n7587_), .Y(new_n7625_));
  XOR2   g06623(.A(new_n7605_), .B(new_n7625_), .Y(new_n7626_));
  XOR2   g06624(.A(new_n7561_), .B(new_n7574_), .Y(new_n7627_));
  NOR2   g06625(.A(new_n7602_), .B(new_n7600_), .Y(new_n7628_));
  AOI21  g06626(.A0(new_n7585_), .A1(\A[246] ), .B0(new_n7628_), .Y(new_n7629_));
  NOR4   g06627(.A(new_n7604_), .B(new_n7598_), .C(new_n7624_), .D(new_n7629_), .Y(new_n7630_));
  NOR2   g06628(.A(new_n7558_), .B(new_n7556_), .Y(new_n7631_));
  AOI21  g06629(.A0(new_n7560_), .A1(\A[240] ), .B0(new_n7631_), .Y(new_n7632_));
  NOR4   g06630(.A(new_n7567_), .B(new_n7632_), .C(new_n7561_), .D(new_n7554_), .Y(new_n7633_));
  NOR4   g06631(.A(new_n7613_), .B(new_n7633_), .C(new_n7630_), .D(new_n7627_), .Y(new_n7634_));
  AOI221 g06632(.A0(new_n7589_), .A1(\A[243] ), .C0(new_n7623_), .B0(new_n7586_), .B1(new_n7584_), .Y(new_n7635_));
  AOI221 g06633(.A0(new_n7590_), .A1(new_n7588_), .C0(new_n7628_), .B0(new_n7585_), .B1(\A[246] ), .Y(new_n7636_));
  OAI211 g06634(.A0(new_n7636_), .A1(new_n7635_), .B0(new_n7617_), .B1(new_n7612_), .Y(new_n7637_));
  NAND2  g06635(.A(new_n7591_), .B(new_n7587_), .Y(new_n7638_));
  AOI21  g06636(.A0(new_n7638_), .A1(new_n7637_), .B0(new_n7613_), .Y(new_n7639_));
  OAI21  g06637(.A0(new_n7639_), .A1(new_n7626_), .B0(new_n7634_), .Y(new_n7640_));
  AOI21  g06638(.A0(new_n7640_), .A1(new_n7622_), .B0(new_n7583_), .Y(new_n7641_));
  XOR2   g06639(.A(new_n7568_), .B(new_n7578_), .Y(new_n7642_));
  XOR2   g06640(.A(new_n7567_), .B(new_n7632_), .Y(new_n7643_));
  NOR2   g06641(.A(new_n7567_), .B(new_n7632_), .Y(new_n7644_));
  AOI21  g06642(.A0(new_n7643_), .A1(new_n7562_), .B0(new_n7644_), .Y(new_n7645_));
  OAI21  g06643(.A0(new_n7645_), .A1(new_n7627_), .B0(new_n7642_), .Y(new_n7646_));
  OAI21  g06644(.A0(new_n7639_), .A1(new_n7626_), .B0(new_n7621_), .Y(new_n7647_));
  NOR2   g06645(.A(new_n7613_), .B(new_n7627_), .Y(new_n7648_));
  OAI211 g06646(.A0(new_n7617_), .A1(new_n7612_), .B0(new_n7591_), .B1(new_n7587_), .Y(new_n7649_));
  NAND4  g06647(.A(new_n7649_), .B(new_n7648_), .C(new_n7619_), .D(new_n7608_), .Y(new_n7650_));
  AOI21  g06648(.A0(new_n7650_), .A1(new_n7647_), .B0(new_n7646_), .Y(new_n7651_));
  NOR2   g06649(.A(new_n7613_), .B(new_n7630_), .Y(new_n7652_));
  XOR2   g06650(.A(new_n7561_), .B(new_n7554_), .Y(new_n7653_));
  XOR2   g06651(.A(new_n7653_), .B(new_n7652_), .Y(new_n7654_));
  INV    g06652(.A(\A[231] ), .Y(new_n7655_));
  INV    g06653(.A(\A[230] ), .Y(new_n7656_));
  NAND2  g06654(.A(new_n7656_), .B(\A[229] ), .Y(new_n7657_));
  INV    g06655(.A(\A[229] ), .Y(new_n7658_));
  AOI21  g06656(.A0(\A[230] ), .A1(new_n7658_), .B0(new_n7655_), .Y(new_n7659_));
  XOR2   g06657(.A(\A[230] ), .B(\A[229] ), .Y(new_n7660_));
  AOI22  g06658(.A0(new_n7660_), .A1(new_n7655_), .B0(new_n7659_), .B1(new_n7657_), .Y(new_n7661_));
  INV    g06659(.A(\A[234] ), .Y(new_n7662_));
  INV    g06660(.A(\A[233] ), .Y(new_n7663_));
  NAND2  g06661(.A(new_n7663_), .B(\A[232] ), .Y(new_n7664_));
  INV    g06662(.A(\A[232] ), .Y(new_n7665_));
  AOI21  g06663(.A0(\A[233] ), .A1(new_n7665_), .B0(new_n7662_), .Y(new_n7666_));
  XOR2   g06664(.A(\A[233] ), .B(\A[232] ), .Y(new_n7667_));
  AOI22  g06665(.A0(new_n7667_), .A1(new_n7662_), .B0(new_n7666_), .B1(new_n7664_), .Y(new_n7668_));
  NOR2   g06666(.A(new_n7663_), .B(new_n7665_), .Y(new_n7669_));
  AOI21  g06667(.A0(new_n7667_), .A1(\A[234] ), .B0(new_n7669_), .Y(new_n7670_));
  NOR2   g06668(.A(new_n7656_), .B(new_n7658_), .Y(new_n7671_));
  AOI21  g06669(.A0(new_n7660_), .A1(\A[231] ), .B0(new_n7671_), .Y(new_n7672_));
  XOR2   g06670(.A(new_n7668_), .B(new_n7661_), .Y(new_n7673_));
  INV    g06671(.A(\A[225] ), .Y(new_n7674_));
  INV    g06672(.A(\A[224] ), .Y(new_n7675_));
  NAND2  g06673(.A(new_n7675_), .B(\A[223] ), .Y(new_n7676_));
  INV    g06674(.A(\A[223] ), .Y(new_n7677_));
  AOI21  g06675(.A0(\A[224] ), .A1(new_n7677_), .B0(new_n7674_), .Y(new_n7678_));
  XOR2   g06676(.A(\A[224] ), .B(\A[223] ), .Y(new_n7679_));
  AOI22  g06677(.A0(new_n7679_), .A1(new_n7674_), .B0(new_n7678_), .B1(new_n7676_), .Y(new_n7680_));
  INV    g06678(.A(\A[228] ), .Y(new_n7681_));
  INV    g06679(.A(\A[227] ), .Y(new_n7682_));
  NAND2  g06680(.A(new_n7682_), .B(\A[226] ), .Y(new_n7683_));
  INV    g06681(.A(\A[226] ), .Y(new_n7684_));
  AOI21  g06682(.A0(\A[227] ), .A1(new_n7684_), .B0(new_n7681_), .Y(new_n7685_));
  XOR2   g06683(.A(\A[227] ), .B(\A[226] ), .Y(new_n7686_));
  AOI22  g06684(.A0(new_n7686_), .A1(new_n7681_), .B0(new_n7685_), .B1(new_n7683_), .Y(new_n7687_));
  NOR2   g06685(.A(new_n7682_), .B(new_n7684_), .Y(new_n7688_));
  AOI21  g06686(.A0(new_n7686_), .A1(\A[228] ), .B0(new_n7688_), .Y(new_n7689_));
  NOR2   g06687(.A(new_n7675_), .B(new_n7677_), .Y(new_n7690_));
  AOI21  g06688(.A0(new_n7679_), .A1(\A[225] ), .B0(new_n7690_), .Y(new_n7691_));
  XOR2   g06689(.A(new_n7687_), .B(new_n7680_), .Y(new_n7692_));
  XOR2   g06690(.A(new_n7692_), .B(new_n7673_), .Y(new_n7693_));
  NAND2  g06691(.A(new_n7693_), .B(new_n7654_), .Y(new_n7694_));
  NOR3   g06692(.A(new_n7694_), .B(new_n7651_), .C(new_n7641_), .Y(new_n7695_));
  OAI21  g06693(.A0(new_n7613_), .A1(new_n7607_), .B0(new_n7608_), .Y(new_n7696_));
  XOR2   g06694(.A(new_n7696_), .B(new_n7621_), .Y(new_n7697_));
  NAND2  g06695(.A(new_n7697_), .B(new_n7646_), .Y(new_n7698_));
  NAND2  g06696(.A(new_n7650_), .B(new_n7647_), .Y(new_n7699_));
  NAND2  g06697(.A(new_n7699_), .B(new_n7583_), .Y(new_n7700_));
  NAND2  g06698(.A(new_n7620_), .B(new_n7618_), .Y(new_n7701_));
  XOR2   g06699(.A(new_n7653_), .B(new_n7701_), .Y(new_n7702_));
  NOR2   g06700(.A(\A[230] ), .B(new_n7658_), .Y(new_n7703_));
  OAI21  g06701(.A0(new_n7656_), .A1(\A[229] ), .B0(\A[231] ), .Y(new_n7704_));
  NAND2  g06702(.A(new_n7660_), .B(new_n7655_), .Y(new_n7705_));
  OAI21  g06703(.A0(new_n7704_), .A1(new_n7703_), .B0(new_n7705_), .Y(new_n7706_));
  XOR2   g06704(.A(new_n7668_), .B(new_n7706_), .Y(new_n7707_));
  XOR2   g06705(.A(new_n7692_), .B(new_n7707_), .Y(new_n7708_));
  NOR2   g06706(.A(new_n7708_), .B(new_n7702_), .Y(new_n7709_));
  AOI21  g06707(.A0(new_n7700_), .A1(new_n7698_), .B0(new_n7709_), .Y(new_n7710_));
  XOR2   g06708(.A(new_n7687_), .B(new_n7680_), .Y(new_n7711_));
  XOR2   g06709(.A(\A[227] ), .B(new_n7684_), .Y(new_n7712_));
  NAND2  g06710(.A(\A[227] ), .B(\A[226] ), .Y(new_n7713_));
  OAI21  g06711(.A0(new_n7712_), .A1(new_n7681_), .B0(new_n7713_), .Y(new_n7714_));
  XOR2   g06712(.A(new_n7691_), .B(new_n7714_), .Y(new_n7715_));
  NOR2   g06713(.A(\A[224] ), .B(new_n7677_), .Y(new_n7716_));
  OAI21  g06714(.A0(new_n7675_), .A1(\A[223] ), .B0(\A[225] ), .Y(new_n7717_));
  XOR2   g06715(.A(\A[224] ), .B(new_n7677_), .Y(new_n7718_));
  OAI22  g06716(.A0(new_n7718_), .A1(\A[225] ), .B0(new_n7717_), .B1(new_n7716_), .Y(new_n7719_));
  NOR2   g06717(.A(\A[227] ), .B(new_n7684_), .Y(new_n7720_));
  OAI21  g06718(.A0(new_n7682_), .A1(\A[226] ), .B0(\A[228] ), .Y(new_n7721_));
  OAI22  g06719(.A0(new_n7712_), .A1(\A[228] ), .B0(new_n7721_), .B1(new_n7720_), .Y(new_n7722_));
  NAND2  g06720(.A(new_n7722_), .B(new_n7719_), .Y(new_n7723_));
  NAND2  g06721(.A(\A[224] ), .B(\A[223] ), .Y(new_n7724_));
  OAI21  g06722(.A0(new_n7718_), .A1(new_n7674_), .B0(new_n7724_), .Y(new_n7725_));
  NAND2  g06723(.A(new_n7725_), .B(new_n7714_), .Y(new_n7726_));
  OAI21  g06724(.A0(new_n7723_), .A1(new_n7715_), .B0(new_n7726_), .Y(new_n7727_));
  NOR2   g06725(.A(new_n7687_), .B(new_n7680_), .Y(new_n7728_));
  XOR2   g06726(.A(new_n7728_), .B(new_n7715_), .Y(new_n7729_));
  AOI21  g06727(.A0(new_n7727_), .A1(new_n7711_), .B0(new_n7729_), .Y(new_n7730_));
  XOR2   g06728(.A(new_n7668_), .B(new_n7706_), .Y(new_n7731_));
  XOR2   g06729(.A(new_n7672_), .B(new_n7670_), .Y(new_n7732_));
  NOR2   g06730(.A(new_n7668_), .B(new_n7661_), .Y(new_n7733_));
  NAND2  g06731(.A(\A[233] ), .B(\A[232] ), .Y(new_n7734_));
  NAND2  g06732(.A(new_n7667_), .B(\A[234] ), .Y(new_n7735_));
  NAND2  g06733(.A(\A[230] ), .B(\A[229] ), .Y(new_n7736_));
  NAND2  g06734(.A(new_n7660_), .B(\A[231] ), .Y(new_n7737_));
  AOI22  g06735(.A0(new_n7737_), .A1(new_n7736_), .B0(new_n7735_), .B1(new_n7734_), .Y(new_n7738_));
  AOI21  g06736(.A0(new_n7733_), .A1(new_n7732_), .B0(new_n7738_), .Y(new_n7739_));
  XOR2   g06737(.A(new_n7733_), .B(new_n7732_), .Y(new_n7740_));
  XOR2   g06738(.A(new_n7668_), .B(new_n7661_), .Y(new_n7741_));
  NOR2   g06739(.A(\A[233] ), .B(new_n7665_), .Y(new_n7742_));
  OAI21  g06740(.A0(new_n7663_), .A1(\A[232] ), .B0(\A[234] ), .Y(new_n7743_));
  NAND2  g06741(.A(new_n7667_), .B(new_n7662_), .Y(new_n7744_));
  OAI21  g06742(.A0(new_n7743_), .A1(new_n7742_), .B0(new_n7744_), .Y(new_n7745_));
  NAND2  g06743(.A(new_n7735_), .B(new_n7734_), .Y(new_n7746_));
  NAND2  g06744(.A(new_n7737_), .B(new_n7736_), .Y(new_n7747_));
  NAND4  g06745(.A(new_n7747_), .B(new_n7746_), .C(new_n7745_), .D(new_n7706_), .Y(new_n7748_));
  NAND4  g06746(.A(new_n7725_), .B(new_n7714_), .C(new_n7722_), .D(new_n7719_), .Y(new_n7749_));
  NAND4  g06747(.A(new_n7749_), .B(new_n7711_), .C(new_n7748_), .D(new_n7741_), .Y(new_n7750_));
  OAI211 g06748(.A0(new_n7739_), .A1(new_n7731_), .B0(new_n7750_), .B1(new_n7740_), .Y(new_n7751_));
  XOR2   g06749(.A(new_n7672_), .B(new_n7746_), .Y(new_n7752_));
  XOR2   g06750(.A(new_n7733_), .B(new_n7752_), .Y(new_n7753_));
  NOR4   g06751(.A(new_n7672_), .B(new_n7670_), .C(new_n7668_), .D(new_n7661_), .Y(new_n7754_));
  XOR2   g06752(.A(new_n7687_), .B(new_n7719_), .Y(new_n7755_));
  NOR3   g06753(.A(new_n7755_), .B(new_n7754_), .C(new_n7731_), .Y(new_n7756_));
  AOI221 g06754(.A0(new_n7735_), .A1(new_n7734_), .C0(new_n7671_), .B0(new_n7660_), .B1(\A[231] ), .Y(new_n7757_));
  AOI221 g06755(.A0(new_n7737_), .A1(new_n7736_), .C0(new_n7669_), .B0(new_n7667_), .B1(\A[234] ), .Y(new_n7758_));
  OAI211 g06756(.A0(new_n7758_), .A1(new_n7757_), .B0(new_n7745_), .B1(new_n7706_), .Y(new_n7759_));
  NAND2  g06757(.A(new_n7747_), .B(new_n7746_), .Y(new_n7760_));
  AOI21  g06758(.A0(new_n7760_), .A1(new_n7759_), .B0(new_n7731_), .Y(new_n7761_));
  OAI211 g06759(.A0(new_n7761_), .A1(new_n7753_), .B0(new_n7756_), .B1(new_n7749_), .Y(new_n7762_));
  AOI21  g06760(.A0(new_n7762_), .A1(new_n7751_), .B0(new_n7730_), .Y(new_n7763_));
  OAI21  g06761(.A0(new_n7761_), .A1(new_n7753_), .B0(new_n7750_), .Y(new_n7764_));
  NAND4  g06762(.A(new_n7711_), .B(new_n7740_), .C(new_n7739_), .D(new_n7741_), .Y(new_n7765_));
  OAI21  g06763(.A0(new_n7739_), .A1(new_n7731_), .B0(new_n7749_), .Y(new_n7766_));
  OAI21  g06764(.A0(new_n7766_), .A1(new_n7765_), .B0(new_n7764_), .Y(new_n7767_));
  AOI21  g06765(.A0(new_n7767_), .A1(new_n7730_), .B0(new_n7763_), .Y(new_n7768_));
  OAI21  g06766(.A0(new_n7710_), .A1(new_n7695_), .B0(new_n7768_), .Y(new_n7769_));
  XOR2   g06767(.A(new_n7691_), .B(new_n7689_), .Y(new_n7770_));
  NOR2   g06768(.A(new_n7691_), .B(new_n7689_), .Y(new_n7771_));
  AOI21  g06769(.A0(new_n7728_), .A1(new_n7770_), .B0(new_n7771_), .Y(new_n7772_));
  XOR2   g06770(.A(new_n7728_), .B(new_n7770_), .Y(new_n7773_));
  OAI21  g06771(.A0(new_n7772_), .A1(new_n7755_), .B0(new_n7773_), .Y(new_n7774_));
  OAI21  g06772(.A0(new_n7739_), .A1(new_n7731_), .B0(new_n7740_), .Y(new_n7775_));
  XOR2   g06773(.A(new_n7775_), .B(new_n7750_), .Y(new_n7776_));
  NAND2  g06774(.A(new_n7776_), .B(new_n7774_), .Y(new_n7777_));
  NAND2  g06775(.A(new_n7767_), .B(new_n7730_), .Y(new_n7778_));
  NAND2  g06776(.A(new_n7778_), .B(new_n7777_), .Y(new_n7779_));
  NAND2  g06777(.A(new_n7620_), .B(new_n7570_), .Y(new_n7780_));
  AOI211 g06778(.A0(new_n7604_), .A1(new_n7598_), .B(new_n7624_), .C(new_n7629_), .Y(new_n7781_));
  NOR4   g06779(.A(new_n7781_), .B(new_n7780_), .C(new_n7633_), .D(new_n7626_), .Y(new_n7782_));
  AOI21  g06780(.A0(new_n7696_), .A1(new_n7621_), .B0(new_n7782_), .Y(new_n7783_));
  OAI21  g06781(.A0(new_n7783_), .A1(new_n7646_), .B0(new_n7694_), .Y(new_n7784_));
  OAI21  g06782(.A0(new_n7651_), .A1(new_n7641_), .B0(new_n7709_), .Y(new_n7785_));
  OAI21  g06783(.A0(new_n7784_), .A1(new_n7641_), .B0(new_n7785_), .Y(new_n7786_));
  NAND2  g06784(.A(new_n7786_), .B(new_n7779_), .Y(new_n7787_));
  NAND2  g06785(.A(new_n7787_), .B(new_n7769_), .Y(new_n7788_));
  INV    g06786(.A(\A[248] ), .Y(new_n7789_));
  NOR2   g06787(.A(new_n7789_), .B(\A[247] ), .Y(new_n7790_));
  INV    g06788(.A(\A[247] ), .Y(new_n7791_));
  OAI21  g06789(.A0(\A[248] ), .A1(new_n7791_), .B0(\A[249] ), .Y(new_n7792_));
  XOR2   g06790(.A(\A[248] ), .B(new_n7791_), .Y(new_n7793_));
  OAI22  g06791(.A0(new_n7793_), .A1(\A[249] ), .B0(new_n7792_), .B1(new_n7790_), .Y(new_n7794_));
  INV    g06792(.A(\A[251] ), .Y(new_n7795_));
  NOR2   g06793(.A(new_n7795_), .B(\A[250] ), .Y(new_n7796_));
  INV    g06794(.A(\A[250] ), .Y(new_n7797_));
  OAI21  g06795(.A0(\A[251] ), .A1(new_n7797_), .B0(\A[252] ), .Y(new_n7798_));
  XOR2   g06796(.A(\A[251] ), .B(new_n7797_), .Y(new_n7799_));
  OAI22  g06797(.A0(new_n7799_), .A1(\A[252] ), .B0(new_n7798_), .B1(new_n7796_), .Y(new_n7800_));
  NAND2  g06798(.A(new_n7800_), .B(new_n7794_), .Y(new_n7801_));
  INV    g06799(.A(\A[252] ), .Y(new_n7802_));
  NAND2  g06800(.A(\A[251] ), .B(\A[250] ), .Y(new_n7803_));
  OAI21  g06801(.A0(new_n7799_), .A1(new_n7802_), .B0(new_n7803_), .Y(new_n7804_));
  XOR2   g06802(.A(\A[248] ), .B(\A[247] ), .Y(new_n7805_));
  NOR2   g06803(.A(new_n7789_), .B(new_n7791_), .Y(new_n7806_));
  AOI21  g06804(.A0(new_n7805_), .A1(\A[249] ), .B0(new_n7806_), .Y(new_n7807_));
  XOR2   g06805(.A(new_n7807_), .B(new_n7804_), .Y(new_n7808_));
  XOR2   g06806(.A(new_n7808_), .B(new_n7801_), .Y(new_n7809_));
  NAND2  g06807(.A(\A[251] ), .B(new_n7797_), .Y(new_n7810_));
  AOI21  g06808(.A0(new_n7795_), .A1(\A[250] ), .B0(new_n7802_), .Y(new_n7811_));
  XOR2   g06809(.A(\A[251] ), .B(\A[250] ), .Y(new_n7812_));
  AOI22  g06810(.A0(new_n7812_), .A1(new_n7802_), .B0(new_n7811_), .B1(new_n7810_), .Y(new_n7813_));
  XOR2   g06811(.A(new_n7813_), .B(new_n7794_), .Y(new_n7814_));
  INV    g06812(.A(\A[249] ), .Y(new_n7815_));
  NAND2  g06813(.A(\A[248] ), .B(new_n7791_), .Y(new_n7816_));
  AOI21  g06814(.A0(new_n7789_), .A1(\A[247] ), .B0(new_n7815_), .Y(new_n7817_));
  AOI22  g06815(.A0(new_n7805_), .A1(new_n7815_), .B0(new_n7817_), .B1(new_n7816_), .Y(new_n7818_));
  NOR2   g06816(.A(new_n7813_), .B(new_n7818_), .Y(new_n7819_));
  NOR2   g06817(.A(new_n7795_), .B(new_n7797_), .Y(new_n7820_));
  AOI21  g06818(.A0(new_n7812_), .A1(\A[252] ), .B0(new_n7820_), .Y(new_n7821_));
  XOR2   g06819(.A(new_n7807_), .B(new_n7821_), .Y(new_n7822_));
  NOR2   g06820(.A(new_n7807_), .B(new_n7821_), .Y(new_n7823_));
  AOI21  g06821(.A0(new_n7822_), .A1(new_n7819_), .B0(new_n7823_), .Y(new_n7824_));
  OAI21  g06822(.A0(new_n7824_), .A1(new_n7814_), .B0(new_n7809_), .Y(new_n7825_));
  XOR2   g06823(.A(new_n7813_), .B(new_n7818_), .Y(new_n7826_));
  NAND2  g06824(.A(\A[257] ), .B(\A[256] ), .Y(new_n7827_));
  XOR2   g06825(.A(\A[257] ), .B(\A[256] ), .Y(new_n7828_));
  NAND2  g06826(.A(new_n7828_), .B(\A[258] ), .Y(new_n7829_));
  NAND2  g06827(.A(new_n7829_), .B(new_n7827_), .Y(new_n7830_));
  NAND2  g06828(.A(\A[254] ), .B(\A[253] ), .Y(new_n7831_));
  XOR2   g06829(.A(\A[254] ), .B(\A[253] ), .Y(new_n7832_));
  NAND2  g06830(.A(new_n7832_), .B(\A[255] ), .Y(new_n7833_));
  NAND2  g06831(.A(new_n7833_), .B(new_n7831_), .Y(new_n7834_));
  INV    g06832(.A(\A[254] ), .Y(new_n7835_));
  NOR2   g06833(.A(new_n7835_), .B(\A[253] ), .Y(new_n7836_));
  INV    g06834(.A(\A[253] ), .Y(new_n7837_));
  OAI21  g06835(.A0(\A[254] ), .A1(new_n7837_), .B0(\A[255] ), .Y(new_n7838_));
  INV    g06836(.A(\A[255] ), .Y(new_n7839_));
  NAND2  g06837(.A(new_n7832_), .B(new_n7839_), .Y(new_n7840_));
  OAI21  g06838(.A0(new_n7838_), .A1(new_n7836_), .B0(new_n7840_), .Y(new_n7841_));
  INV    g06839(.A(\A[257] ), .Y(new_n7842_));
  NOR2   g06840(.A(new_n7842_), .B(\A[256] ), .Y(new_n7843_));
  INV    g06841(.A(\A[256] ), .Y(new_n7844_));
  OAI21  g06842(.A0(\A[257] ), .A1(new_n7844_), .B0(\A[258] ), .Y(new_n7845_));
  INV    g06843(.A(\A[258] ), .Y(new_n7846_));
  NAND2  g06844(.A(new_n7828_), .B(new_n7846_), .Y(new_n7847_));
  OAI21  g06845(.A0(new_n7845_), .A1(new_n7843_), .B0(new_n7847_), .Y(new_n7848_));
  NAND4  g06846(.A(new_n7848_), .B(new_n7841_), .C(new_n7834_), .D(new_n7830_), .Y(new_n7849_));
  NAND2  g06847(.A(\A[248] ), .B(\A[247] ), .Y(new_n7850_));
  OAI21  g06848(.A0(new_n7793_), .A1(new_n7815_), .B0(new_n7850_), .Y(new_n7851_));
  NAND4  g06849(.A(new_n7851_), .B(new_n7804_), .C(new_n7800_), .D(new_n7794_), .Y(new_n7852_));
  NAND2  g06850(.A(\A[254] ), .B(new_n7837_), .Y(new_n7853_));
  AOI21  g06851(.A0(new_n7835_), .A1(\A[253] ), .B0(new_n7839_), .Y(new_n7854_));
  AOI22  g06852(.A0(new_n7854_), .A1(new_n7853_), .B0(new_n7832_), .B1(new_n7839_), .Y(new_n7855_));
  NAND2  g06853(.A(\A[257] ), .B(new_n7844_), .Y(new_n7856_));
  AOI21  g06854(.A0(new_n7842_), .A1(\A[256] ), .B0(new_n7846_), .Y(new_n7857_));
  AOI22  g06855(.A0(new_n7857_), .A1(new_n7856_), .B0(new_n7828_), .B1(new_n7846_), .Y(new_n7858_));
  XOR2   g06856(.A(new_n7858_), .B(new_n7855_), .Y(new_n7859_));
  NAND4  g06857(.A(new_n7859_), .B(new_n7852_), .C(new_n7849_), .D(new_n7826_), .Y(new_n7860_));
  XOR2   g06858(.A(new_n7834_), .B(new_n7830_), .Y(new_n7861_));
  NOR2   g06859(.A(new_n7858_), .B(new_n7855_), .Y(new_n7862_));
  AOI22  g06860(.A0(new_n7833_), .A1(new_n7831_), .B0(new_n7829_), .B1(new_n7827_), .Y(new_n7863_));
  AOI21  g06861(.A0(new_n7862_), .A1(new_n7861_), .B0(new_n7863_), .Y(new_n7864_));
  XOR2   g06862(.A(new_n7862_), .B(new_n7861_), .Y(new_n7865_));
  XOR2   g06863(.A(new_n7858_), .B(new_n7841_), .Y(new_n7866_));
  OAI21  g06864(.A0(new_n7866_), .A1(new_n7864_), .B0(new_n7865_), .Y(new_n7867_));
  XOR2   g06865(.A(new_n7867_), .B(new_n7860_), .Y(new_n7868_));
  NAND2  g06866(.A(new_n7848_), .B(new_n7841_), .Y(new_n7869_));
  XOR2   g06867(.A(new_n7869_), .B(new_n7861_), .Y(new_n7870_));
  NOR2   g06868(.A(new_n7835_), .B(new_n7837_), .Y(new_n7871_));
  AOI221 g06869(.A0(new_n7832_), .A1(\A[255] ), .C0(new_n7871_), .B0(new_n7829_), .B1(new_n7827_), .Y(new_n7872_));
  NOR2   g06870(.A(new_n7842_), .B(new_n7844_), .Y(new_n7873_));
  AOI221 g06871(.A0(new_n7833_), .A1(new_n7831_), .C0(new_n7873_), .B0(new_n7828_), .B1(\A[258] ), .Y(new_n7874_));
  OAI211 g06872(.A0(new_n7874_), .A1(new_n7872_), .B0(new_n7848_), .B1(new_n7841_), .Y(new_n7875_));
  NAND2  g06873(.A(new_n7834_), .B(new_n7830_), .Y(new_n7876_));
  AOI21  g06874(.A0(new_n7876_), .A1(new_n7875_), .B0(new_n7866_), .Y(new_n7877_));
  OAI21  g06875(.A0(new_n7877_), .A1(new_n7870_), .B0(new_n7860_), .Y(new_n7878_));
  NOR2   g06876(.A(new_n7866_), .B(new_n7814_), .Y(new_n7879_));
  OAI211 g06877(.A0(new_n7848_), .A1(new_n7841_), .B0(new_n7834_), .B1(new_n7830_), .Y(new_n7880_));
  NAND4  g06878(.A(new_n7880_), .B(new_n7879_), .C(new_n7852_), .D(new_n7865_), .Y(new_n7881_));
  AOI21  g06879(.A0(new_n7881_), .A1(new_n7878_), .B0(new_n7825_), .Y(new_n7882_));
  AOI21  g06880(.A0(new_n7868_), .A1(new_n7825_), .B0(new_n7882_), .Y(new_n7883_));
  INV    g06881(.A(\A[261] ), .Y(new_n7884_));
  INV    g06882(.A(\A[259] ), .Y(new_n7885_));
  NAND2  g06883(.A(\A[260] ), .B(new_n7885_), .Y(new_n7886_));
  INV    g06884(.A(\A[260] ), .Y(new_n7887_));
  AOI21  g06885(.A0(new_n7887_), .A1(\A[259] ), .B0(new_n7884_), .Y(new_n7888_));
  XOR2   g06886(.A(\A[260] ), .B(\A[259] ), .Y(new_n7889_));
  AOI22  g06887(.A0(new_n7889_), .A1(new_n7884_), .B0(new_n7888_), .B1(new_n7886_), .Y(new_n7890_));
  INV    g06888(.A(\A[264] ), .Y(new_n7891_));
  INV    g06889(.A(\A[262] ), .Y(new_n7892_));
  NAND2  g06890(.A(\A[263] ), .B(new_n7892_), .Y(new_n7893_));
  INV    g06891(.A(\A[263] ), .Y(new_n7894_));
  AOI21  g06892(.A0(new_n7894_), .A1(\A[262] ), .B0(new_n7891_), .Y(new_n7895_));
  XOR2   g06893(.A(\A[263] ), .B(\A[262] ), .Y(new_n7896_));
  AOI22  g06894(.A0(new_n7896_), .A1(new_n7891_), .B0(new_n7895_), .B1(new_n7893_), .Y(new_n7897_));
  NOR2   g06895(.A(new_n7897_), .B(new_n7890_), .Y(new_n7898_));
  XOR2   g06896(.A(\A[263] ), .B(new_n7892_), .Y(new_n7899_));
  NAND2  g06897(.A(\A[263] ), .B(\A[262] ), .Y(new_n7900_));
  OAI21  g06898(.A0(new_n7899_), .A1(new_n7891_), .B0(new_n7900_), .Y(new_n7901_));
  NOR2   g06899(.A(new_n7887_), .B(new_n7885_), .Y(new_n7902_));
  AOI21  g06900(.A0(new_n7889_), .A1(\A[261] ), .B0(new_n7902_), .Y(new_n7903_));
  XOR2   g06901(.A(new_n7903_), .B(new_n7901_), .Y(new_n7904_));
  XOR2   g06902(.A(new_n7904_), .B(new_n7898_), .Y(new_n7905_));
  XOR2   g06903(.A(new_n7897_), .B(new_n7890_), .Y(new_n7906_));
  NOR2   g06904(.A(new_n7887_), .B(\A[259] ), .Y(new_n7907_));
  OAI21  g06905(.A0(\A[260] ), .A1(new_n7885_), .B0(\A[261] ), .Y(new_n7908_));
  XOR2   g06906(.A(\A[260] ), .B(new_n7885_), .Y(new_n7909_));
  OAI22  g06907(.A0(new_n7909_), .A1(\A[261] ), .B0(new_n7908_), .B1(new_n7907_), .Y(new_n7910_));
  NOR2   g06908(.A(new_n7894_), .B(\A[262] ), .Y(new_n7911_));
  OAI21  g06909(.A0(\A[263] ), .A1(new_n7892_), .B0(\A[264] ), .Y(new_n7912_));
  OAI22  g06910(.A0(new_n7899_), .A1(\A[264] ), .B0(new_n7912_), .B1(new_n7911_), .Y(new_n7913_));
  NAND2  g06911(.A(new_n7913_), .B(new_n7910_), .Y(new_n7914_));
  NAND2  g06912(.A(\A[260] ), .B(\A[259] ), .Y(new_n7915_));
  OAI21  g06913(.A0(new_n7909_), .A1(new_n7884_), .B0(new_n7915_), .Y(new_n7916_));
  NAND2  g06914(.A(new_n7916_), .B(new_n7901_), .Y(new_n7917_));
  OAI21  g06915(.A0(new_n7904_), .A1(new_n7914_), .B0(new_n7917_), .Y(new_n7918_));
  AOI21  g06916(.A0(new_n7918_), .A1(new_n7906_), .B0(new_n7905_), .Y(new_n7919_));
  NAND2  g06917(.A(\A[269] ), .B(\A[268] ), .Y(new_n7920_));
  XOR2   g06918(.A(\A[269] ), .B(\A[268] ), .Y(new_n7921_));
  NAND2  g06919(.A(new_n7921_), .B(\A[270] ), .Y(new_n7922_));
  NAND2  g06920(.A(new_n7922_), .B(new_n7920_), .Y(new_n7923_));
  NAND2  g06921(.A(\A[266] ), .B(\A[265] ), .Y(new_n7924_));
  XOR2   g06922(.A(\A[266] ), .B(\A[265] ), .Y(new_n7925_));
  NAND2  g06923(.A(new_n7925_), .B(\A[267] ), .Y(new_n7926_));
  NAND2  g06924(.A(new_n7926_), .B(new_n7924_), .Y(new_n7927_));
  XOR2   g06925(.A(new_n7927_), .B(new_n7923_), .Y(new_n7928_));
  INV    g06926(.A(\A[267] ), .Y(new_n7929_));
  INV    g06927(.A(\A[265] ), .Y(new_n7930_));
  NAND2  g06928(.A(\A[266] ), .B(new_n7930_), .Y(new_n7931_));
  INV    g06929(.A(\A[266] ), .Y(new_n7932_));
  AOI21  g06930(.A0(new_n7932_), .A1(\A[265] ), .B0(new_n7929_), .Y(new_n7933_));
  AOI22  g06931(.A0(new_n7933_), .A1(new_n7931_), .B0(new_n7925_), .B1(new_n7929_), .Y(new_n7934_));
  INV    g06932(.A(\A[270] ), .Y(new_n7935_));
  INV    g06933(.A(\A[268] ), .Y(new_n7936_));
  NAND2  g06934(.A(\A[269] ), .B(new_n7936_), .Y(new_n7937_));
  INV    g06935(.A(\A[269] ), .Y(new_n7938_));
  AOI21  g06936(.A0(new_n7938_), .A1(\A[268] ), .B0(new_n7935_), .Y(new_n7939_));
  AOI22  g06937(.A0(new_n7939_), .A1(new_n7937_), .B0(new_n7921_), .B1(new_n7935_), .Y(new_n7940_));
  NOR2   g06938(.A(new_n7940_), .B(new_n7934_), .Y(new_n7941_));
  AOI22  g06939(.A0(new_n7926_), .A1(new_n7924_), .B0(new_n7922_), .B1(new_n7920_), .Y(new_n7942_));
  AOI21  g06940(.A0(new_n7941_), .A1(new_n7928_), .B0(new_n7942_), .Y(new_n7943_));
  XOR2   g06941(.A(new_n7941_), .B(new_n7928_), .Y(new_n7944_));
  NOR2   g06942(.A(new_n7932_), .B(\A[265] ), .Y(new_n7945_));
  OAI21  g06943(.A0(\A[266] ), .A1(new_n7930_), .B0(\A[267] ), .Y(new_n7946_));
  NAND2  g06944(.A(new_n7925_), .B(new_n7929_), .Y(new_n7947_));
  OAI21  g06945(.A0(new_n7946_), .A1(new_n7945_), .B0(new_n7947_), .Y(new_n7948_));
  XOR2   g06946(.A(new_n7940_), .B(new_n7948_), .Y(new_n7949_));
  NOR2   g06947(.A(new_n7938_), .B(\A[268] ), .Y(new_n7950_));
  OAI21  g06948(.A0(\A[269] ), .A1(new_n7936_), .B0(\A[270] ), .Y(new_n7951_));
  NAND2  g06949(.A(new_n7921_), .B(new_n7935_), .Y(new_n7952_));
  OAI21  g06950(.A0(new_n7951_), .A1(new_n7950_), .B0(new_n7952_), .Y(new_n7953_));
  NAND4  g06951(.A(new_n7953_), .B(new_n7948_), .C(new_n7927_), .D(new_n7923_), .Y(new_n7954_));
  NAND4  g06952(.A(new_n7916_), .B(new_n7901_), .C(new_n7913_), .D(new_n7910_), .Y(new_n7955_));
  XOR2   g06953(.A(new_n7940_), .B(new_n7934_), .Y(new_n7956_));
  NAND4  g06954(.A(new_n7956_), .B(new_n7955_), .C(new_n7954_), .D(new_n7906_), .Y(new_n7957_));
  OAI211 g06955(.A0(new_n7949_), .A1(new_n7943_), .B0(new_n7957_), .B1(new_n7944_), .Y(new_n7958_));
  NOR2   g06956(.A(new_n7932_), .B(new_n7930_), .Y(new_n7959_));
  AOI21  g06957(.A0(new_n7925_), .A1(\A[267] ), .B0(new_n7959_), .Y(new_n7960_));
  XOR2   g06958(.A(new_n7960_), .B(new_n7923_), .Y(new_n7961_));
  XOR2   g06959(.A(new_n7941_), .B(new_n7961_), .Y(new_n7962_));
  XOR2   g06960(.A(new_n7897_), .B(new_n7910_), .Y(new_n7963_));
  NOR2   g06961(.A(new_n7938_), .B(new_n7936_), .Y(new_n7964_));
  AOI21  g06962(.A0(new_n7921_), .A1(\A[270] ), .B0(new_n7964_), .Y(new_n7965_));
  NOR4   g06963(.A(new_n7940_), .B(new_n7934_), .C(new_n7960_), .D(new_n7965_), .Y(new_n7966_));
  NOR2   g06964(.A(new_n7894_), .B(new_n7892_), .Y(new_n7967_));
  AOI21  g06965(.A0(new_n7896_), .A1(\A[264] ), .B0(new_n7967_), .Y(new_n7968_));
  NOR4   g06966(.A(new_n7903_), .B(new_n7968_), .C(new_n7897_), .D(new_n7890_), .Y(new_n7969_));
  NOR4   g06967(.A(new_n7949_), .B(new_n7969_), .C(new_n7966_), .D(new_n7963_), .Y(new_n7970_));
  AOI221 g06968(.A0(new_n7925_), .A1(\A[267] ), .C0(new_n7959_), .B0(new_n7922_), .B1(new_n7920_), .Y(new_n7971_));
  AOI221 g06969(.A0(new_n7926_), .A1(new_n7924_), .C0(new_n7964_), .B0(new_n7921_), .B1(\A[270] ), .Y(new_n7972_));
  OAI211 g06970(.A0(new_n7972_), .A1(new_n7971_), .B0(new_n7953_), .B1(new_n7948_), .Y(new_n7973_));
  NAND2  g06971(.A(new_n7927_), .B(new_n7923_), .Y(new_n7974_));
  AOI21  g06972(.A0(new_n7974_), .A1(new_n7973_), .B0(new_n7949_), .Y(new_n7975_));
  OAI21  g06973(.A0(new_n7975_), .A1(new_n7962_), .B0(new_n7970_), .Y(new_n7976_));
  AOI21  g06974(.A0(new_n7976_), .A1(new_n7958_), .B0(new_n7919_), .Y(new_n7977_));
  XOR2   g06975(.A(new_n7904_), .B(new_n7914_), .Y(new_n7978_));
  XOR2   g06976(.A(new_n7903_), .B(new_n7968_), .Y(new_n7979_));
  NOR2   g06977(.A(new_n7903_), .B(new_n7968_), .Y(new_n7980_));
  AOI21  g06978(.A0(new_n7979_), .A1(new_n7898_), .B0(new_n7980_), .Y(new_n7981_));
  OAI21  g06979(.A0(new_n7981_), .A1(new_n7963_), .B0(new_n7978_), .Y(new_n7982_));
  OAI21  g06980(.A0(new_n7975_), .A1(new_n7962_), .B0(new_n7957_), .Y(new_n7983_));
  NOR2   g06981(.A(new_n7949_), .B(new_n7963_), .Y(new_n7984_));
  OAI211 g06982(.A0(new_n7953_), .A1(new_n7948_), .B0(new_n7927_), .B1(new_n7923_), .Y(new_n7985_));
  NAND4  g06983(.A(new_n7985_), .B(new_n7984_), .C(new_n7955_), .D(new_n7944_), .Y(new_n7986_));
  AOI21  g06984(.A0(new_n7986_), .A1(new_n7983_), .B0(new_n7982_), .Y(new_n7987_));
  NOR2   g06985(.A(new_n7949_), .B(new_n7966_), .Y(new_n7988_));
  XOR2   g06986(.A(new_n7897_), .B(new_n7890_), .Y(new_n7989_));
  XOR2   g06987(.A(new_n7989_), .B(new_n7988_), .Y(new_n7990_));
  NAND2  g06988(.A(new_n7859_), .B(new_n7849_), .Y(new_n7991_));
  XOR2   g06989(.A(new_n7813_), .B(new_n7794_), .Y(new_n7992_));
  XOR2   g06990(.A(new_n7992_), .B(new_n7991_), .Y(new_n7993_));
  NAND2  g06991(.A(new_n7993_), .B(new_n7990_), .Y(new_n7994_));
  NOR3   g06992(.A(new_n7994_), .B(new_n7987_), .C(new_n7977_), .Y(new_n7995_));
  OAI21  g06993(.A0(new_n7949_), .A1(new_n7943_), .B0(new_n7944_), .Y(new_n7996_));
  XOR2   g06994(.A(new_n7996_), .B(new_n7957_), .Y(new_n7997_));
  NAND2  g06995(.A(new_n7997_), .B(new_n7982_), .Y(new_n7998_));
  NAND2  g06996(.A(new_n7986_), .B(new_n7983_), .Y(new_n7999_));
  NAND2  g06997(.A(new_n7999_), .B(new_n7919_), .Y(new_n8000_));
  NAND2  g06998(.A(new_n7956_), .B(new_n7954_), .Y(new_n8001_));
  XOR2   g06999(.A(new_n7989_), .B(new_n8001_), .Y(new_n8002_));
  XOR2   g07000(.A(new_n7813_), .B(new_n7818_), .Y(new_n8003_));
  XOR2   g07001(.A(new_n8003_), .B(new_n7991_), .Y(new_n8004_));
  NOR2   g07002(.A(new_n8004_), .B(new_n8002_), .Y(new_n8005_));
  AOI21  g07003(.A0(new_n8000_), .A1(new_n7998_), .B0(new_n8005_), .Y(new_n8006_));
  OAI21  g07004(.A0(new_n8006_), .A1(new_n7995_), .B0(new_n7883_), .Y(new_n8007_));
  XOR2   g07005(.A(new_n7808_), .B(new_n7819_), .Y(new_n8008_));
  NAND2  g07006(.A(new_n7851_), .B(new_n7804_), .Y(new_n8009_));
  OAI21  g07007(.A0(new_n7808_), .A1(new_n7801_), .B0(new_n8009_), .Y(new_n8010_));
  AOI21  g07008(.A0(new_n8010_), .A1(new_n7826_), .B0(new_n8008_), .Y(new_n8011_));
  NOR2   g07009(.A(new_n7877_), .B(new_n7870_), .Y(new_n8012_));
  XOR2   g07010(.A(new_n8012_), .B(new_n7860_), .Y(new_n8013_));
  NAND2  g07011(.A(new_n7881_), .B(new_n7878_), .Y(new_n8014_));
  NAND2  g07012(.A(new_n8014_), .B(new_n8011_), .Y(new_n8015_));
  OAI21  g07013(.A0(new_n8013_), .A1(new_n8011_), .B0(new_n8015_), .Y(new_n8016_));
  NAND2  g07014(.A(new_n7956_), .B(new_n7906_), .Y(new_n8017_));
  AOI211 g07015(.A0(new_n7940_), .A1(new_n7934_), .B(new_n7960_), .C(new_n7965_), .Y(new_n8018_));
  NOR4   g07016(.A(new_n8018_), .B(new_n8017_), .C(new_n7969_), .D(new_n7962_), .Y(new_n8019_));
  AOI21  g07017(.A0(new_n7996_), .A1(new_n7957_), .B0(new_n8019_), .Y(new_n8020_));
  OAI21  g07018(.A0(new_n8020_), .A1(new_n7982_), .B0(new_n7994_), .Y(new_n8021_));
  OAI21  g07019(.A0(new_n7987_), .A1(new_n7977_), .B0(new_n8005_), .Y(new_n8022_));
  OAI21  g07020(.A0(new_n8021_), .A1(new_n7977_), .B0(new_n8022_), .Y(new_n8023_));
  NAND2  g07021(.A(new_n8023_), .B(new_n8016_), .Y(new_n8024_));
  XOR2   g07022(.A(new_n8004_), .B(new_n7990_), .Y(new_n8025_));
  XOR2   g07023(.A(new_n7708_), .B(new_n7654_), .Y(new_n8026_));
  NOR2   g07024(.A(new_n8026_), .B(new_n8025_), .Y(new_n8027_));
  NAND3  g07025(.A(new_n8027_), .B(new_n8024_), .C(new_n8007_), .Y(new_n8028_));
  NAND3  g07026(.A(new_n8005_), .B(new_n8000_), .C(new_n7998_), .Y(new_n8029_));
  OAI21  g07027(.A0(new_n7987_), .A1(new_n7977_), .B0(new_n7994_), .Y(new_n8030_));
  AOI21  g07028(.A0(new_n8030_), .A1(new_n8029_), .B0(new_n8016_), .Y(new_n8031_));
  NAND3  g07029(.A(new_n7994_), .B(new_n8000_), .C(new_n7998_), .Y(new_n8032_));
  AOI21  g07030(.A0(new_n8022_), .A1(new_n8032_), .B0(new_n7883_), .Y(new_n8033_));
  INV    g07031(.A(new_n8027_), .Y(new_n8034_));
  OAI21  g07032(.A0(new_n8033_), .A1(new_n8031_), .B0(new_n8034_), .Y(new_n8035_));
  AOI21  g07033(.A0(new_n8035_), .A1(new_n8028_), .B0(new_n7788_), .Y(new_n8036_));
  NAND3  g07034(.A(new_n7709_), .B(new_n7700_), .C(new_n7698_), .Y(new_n8037_));
  OAI21  g07035(.A0(new_n7651_), .A1(new_n7641_), .B0(new_n7694_), .Y(new_n8038_));
  AOI21  g07036(.A0(new_n8038_), .A1(new_n8037_), .B0(new_n7779_), .Y(new_n8039_));
  AOI21  g07037(.A0(new_n7786_), .A1(new_n7779_), .B0(new_n8039_), .Y(new_n8040_));
  AOI21  g07038(.A0(new_n8023_), .A1(new_n8016_), .B0(new_n8027_), .Y(new_n8041_));
  NAND2  g07039(.A(new_n8041_), .B(new_n8007_), .Y(new_n8042_));
  OAI21  g07040(.A0(new_n8033_), .A1(new_n8031_), .B0(new_n8027_), .Y(new_n8043_));
  AOI21  g07041(.A0(new_n8043_), .A1(new_n8042_), .B0(new_n8040_), .Y(new_n8044_));
  XOR2   g07042(.A(new_n8026_), .B(new_n8025_), .Y(new_n8045_));
  INV    g07043(.A(new_n8045_), .Y(new_n8046_));
  XOR2   g07044(.A(new_n7372_), .B(new_n7292_), .Y(new_n8047_));
  INV    g07045(.A(new_n8047_), .Y(new_n8048_));
  NOR2   g07046(.A(new_n8048_), .B(new_n8046_), .Y(new_n8049_));
  INV    g07047(.A(new_n8049_), .Y(new_n8050_));
  NOR3   g07048(.A(new_n8050_), .B(new_n8044_), .C(new_n8036_), .Y(new_n8051_));
  NOR3   g07049(.A(new_n8034_), .B(new_n8033_), .C(new_n8031_), .Y(new_n8052_));
  AOI21  g07050(.A0(new_n8024_), .A1(new_n8007_), .B0(new_n8027_), .Y(new_n8053_));
  OAI21  g07051(.A0(new_n8053_), .A1(new_n8052_), .B0(new_n8040_), .Y(new_n8054_));
  NOR3   g07052(.A(new_n8027_), .B(new_n8033_), .C(new_n8031_), .Y(new_n8055_));
  AOI21  g07053(.A0(new_n8024_), .A1(new_n8007_), .B0(new_n8034_), .Y(new_n8056_));
  OAI21  g07054(.A0(new_n8056_), .A1(new_n8055_), .B0(new_n7788_), .Y(new_n8057_));
  AOI21  g07055(.A0(new_n8057_), .A1(new_n8054_), .B0(new_n8049_), .Y(new_n8058_));
  OAI21  g07056(.A0(new_n8058_), .A1(new_n8051_), .B0(new_n7547_), .Y(new_n8059_));
  NOR3   g07057(.A(new_n7380_), .B(new_n7379_), .C(new_n7377_), .Y(new_n8060_));
  AOI21  g07058(.A0(new_n7291_), .A1(new_n7277_), .B0(new_n7373_), .Y(new_n8061_));
  OAI21  g07059(.A0(new_n8061_), .A1(new_n8060_), .B0(new_n7542_), .Y(new_n8062_));
  NOR3   g07060(.A(new_n7373_), .B(new_n7379_), .C(new_n7377_), .Y(new_n8063_));
  AOI21  g07061(.A0(new_n7291_), .A1(new_n7277_), .B0(new_n7380_), .Y(new_n8064_));
  OAI21  g07062(.A0(new_n8064_), .A1(new_n8063_), .B0(new_n7522_), .Y(new_n8065_));
  NAND2  g07063(.A(new_n8065_), .B(new_n8062_), .Y(new_n8066_));
  NOR3   g07064(.A(new_n8049_), .B(new_n8044_), .C(new_n8036_), .Y(new_n8067_));
  AOI21  g07065(.A0(new_n8057_), .A1(new_n8054_), .B0(new_n8050_), .Y(new_n8068_));
  OAI21  g07066(.A0(new_n8068_), .A1(new_n8067_), .B0(new_n8066_), .Y(new_n8069_));
  XOR2   g07067(.A(new_n8048_), .B(new_n8045_), .Y(new_n8070_));
  INV    g07068(.A(\A[171] ), .Y(new_n8071_));
  INV    g07069(.A(\A[170] ), .Y(new_n8072_));
  NAND2  g07070(.A(new_n8072_), .B(\A[169] ), .Y(new_n8073_));
  INV    g07071(.A(\A[169] ), .Y(new_n8074_));
  AOI21  g07072(.A0(\A[170] ), .A1(new_n8074_), .B0(new_n8071_), .Y(new_n8075_));
  XOR2   g07073(.A(\A[170] ), .B(\A[169] ), .Y(new_n8076_));
  AOI22  g07074(.A0(new_n8076_), .A1(new_n8071_), .B0(new_n8075_), .B1(new_n8073_), .Y(new_n8077_));
  INV    g07075(.A(\A[174] ), .Y(new_n8078_));
  INV    g07076(.A(\A[173] ), .Y(new_n8079_));
  NAND2  g07077(.A(new_n8079_), .B(\A[172] ), .Y(new_n8080_));
  INV    g07078(.A(\A[172] ), .Y(new_n8081_));
  AOI21  g07079(.A0(\A[173] ), .A1(new_n8081_), .B0(new_n8078_), .Y(new_n8082_));
  XOR2   g07080(.A(\A[173] ), .B(\A[172] ), .Y(new_n8083_));
  AOI22  g07081(.A0(new_n8083_), .A1(new_n8078_), .B0(new_n8082_), .B1(new_n8080_), .Y(new_n8084_));
  NOR2   g07082(.A(new_n8079_), .B(new_n8081_), .Y(new_n8085_));
  AOI21  g07083(.A0(new_n8083_), .A1(\A[174] ), .B0(new_n8085_), .Y(new_n8086_));
  NOR2   g07084(.A(new_n8072_), .B(new_n8074_), .Y(new_n8087_));
  AOI21  g07085(.A0(new_n8076_), .A1(\A[171] ), .B0(new_n8087_), .Y(new_n8088_));
  XOR2   g07086(.A(new_n8084_), .B(new_n8077_), .Y(new_n8089_));
  INV    g07087(.A(\A[165] ), .Y(new_n8090_));
  INV    g07088(.A(\A[164] ), .Y(new_n8091_));
  NAND2  g07089(.A(new_n8091_), .B(\A[163] ), .Y(new_n8092_));
  INV    g07090(.A(\A[163] ), .Y(new_n8093_));
  AOI21  g07091(.A0(\A[164] ), .A1(new_n8093_), .B0(new_n8090_), .Y(new_n8094_));
  XOR2   g07092(.A(\A[164] ), .B(\A[163] ), .Y(new_n8095_));
  AOI22  g07093(.A0(new_n8095_), .A1(new_n8090_), .B0(new_n8094_), .B1(new_n8092_), .Y(new_n8096_));
  INV    g07094(.A(\A[168] ), .Y(new_n8097_));
  INV    g07095(.A(\A[167] ), .Y(new_n8098_));
  NAND2  g07096(.A(new_n8098_), .B(\A[166] ), .Y(new_n8099_));
  INV    g07097(.A(\A[166] ), .Y(new_n8100_));
  AOI21  g07098(.A0(\A[167] ), .A1(new_n8100_), .B0(new_n8097_), .Y(new_n8101_));
  XOR2   g07099(.A(\A[167] ), .B(\A[166] ), .Y(new_n8102_));
  AOI22  g07100(.A0(new_n8102_), .A1(new_n8097_), .B0(new_n8101_), .B1(new_n8099_), .Y(new_n8103_));
  NOR2   g07101(.A(new_n8098_), .B(new_n8100_), .Y(new_n8104_));
  AOI21  g07102(.A0(new_n8102_), .A1(\A[168] ), .B0(new_n8104_), .Y(new_n8105_));
  NOR2   g07103(.A(new_n8091_), .B(new_n8093_), .Y(new_n8106_));
  AOI21  g07104(.A0(new_n8095_), .A1(\A[165] ), .B0(new_n8106_), .Y(new_n8107_));
  XOR2   g07105(.A(new_n8103_), .B(new_n8096_), .Y(new_n8108_));
  XOR2   g07106(.A(new_n8108_), .B(new_n8089_), .Y(new_n8109_));
  INV    g07107(.A(\A[157] ), .Y(new_n8110_));
  NOR2   g07108(.A(\A[158] ), .B(new_n8110_), .Y(new_n8111_));
  INV    g07109(.A(\A[158] ), .Y(new_n8112_));
  OAI21  g07110(.A0(new_n8112_), .A1(\A[157] ), .B0(\A[159] ), .Y(new_n8113_));
  INV    g07111(.A(\A[159] ), .Y(new_n8114_));
  XOR2   g07112(.A(\A[158] ), .B(\A[157] ), .Y(new_n8115_));
  NAND2  g07113(.A(new_n8115_), .B(new_n8114_), .Y(new_n8116_));
  OAI21  g07114(.A0(new_n8113_), .A1(new_n8111_), .B0(new_n8116_), .Y(new_n8117_));
  INV    g07115(.A(\A[162] ), .Y(new_n8118_));
  INV    g07116(.A(\A[161] ), .Y(new_n8119_));
  NAND2  g07117(.A(new_n8119_), .B(\A[160] ), .Y(new_n8120_));
  INV    g07118(.A(\A[160] ), .Y(new_n8121_));
  AOI21  g07119(.A0(\A[161] ), .A1(new_n8121_), .B0(new_n8118_), .Y(new_n8122_));
  XOR2   g07120(.A(\A[161] ), .B(\A[160] ), .Y(new_n8123_));
  AOI22  g07121(.A0(new_n8123_), .A1(new_n8118_), .B0(new_n8122_), .B1(new_n8120_), .Y(new_n8124_));
  NOR2   g07122(.A(new_n8119_), .B(new_n8121_), .Y(new_n8125_));
  AOI21  g07123(.A0(new_n8123_), .A1(\A[162] ), .B0(new_n8125_), .Y(new_n8126_));
  NOR2   g07124(.A(new_n8112_), .B(new_n8110_), .Y(new_n8127_));
  AOI21  g07125(.A0(new_n8115_), .A1(\A[159] ), .B0(new_n8127_), .Y(new_n8128_));
  XOR2   g07126(.A(new_n8124_), .B(new_n8117_), .Y(new_n8129_));
  INV    g07127(.A(\A[153] ), .Y(new_n8130_));
  INV    g07128(.A(\A[152] ), .Y(new_n8131_));
  NAND2  g07129(.A(new_n8131_), .B(\A[151] ), .Y(new_n8132_));
  INV    g07130(.A(\A[151] ), .Y(new_n8133_));
  AOI21  g07131(.A0(\A[152] ), .A1(new_n8133_), .B0(new_n8130_), .Y(new_n8134_));
  XOR2   g07132(.A(\A[152] ), .B(\A[151] ), .Y(new_n8135_));
  AOI22  g07133(.A0(new_n8135_), .A1(new_n8130_), .B0(new_n8134_), .B1(new_n8132_), .Y(new_n8136_));
  INV    g07134(.A(\A[156] ), .Y(new_n8137_));
  INV    g07135(.A(\A[155] ), .Y(new_n8138_));
  NAND2  g07136(.A(new_n8138_), .B(\A[154] ), .Y(new_n8139_));
  INV    g07137(.A(\A[154] ), .Y(new_n8140_));
  AOI21  g07138(.A0(\A[155] ), .A1(new_n8140_), .B0(new_n8137_), .Y(new_n8141_));
  XOR2   g07139(.A(\A[155] ), .B(\A[154] ), .Y(new_n8142_));
  AOI22  g07140(.A0(new_n8142_), .A1(new_n8137_), .B0(new_n8141_), .B1(new_n8139_), .Y(new_n8143_));
  NOR2   g07141(.A(new_n8138_), .B(new_n8140_), .Y(new_n8144_));
  AOI21  g07142(.A0(new_n8142_), .A1(\A[156] ), .B0(new_n8144_), .Y(new_n8145_));
  NOR2   g07143(.A(new_n8131_), .B(new_n8133_), .Y(new_n8146_));
  AOI21  g07144(.A0(new_n8135_), .A1(\A[153] ), .B0(new_n8146_), .Y(new_n8147_));
  XOR2   g07145(.A(new_n8143_), .B(new_n8136_), .Y(new_n8148_));
  XOR2   g07146(.A(new_n8148_), .B(new_n8129_), .Y(new_n8149_));
  XOR2   g07147(.A(new_n8149_), .B(new_n8109_), .Y(new_n8150_));
  INV    g07148(.A(new_n8150_), .Y(new_n8151_));
  INV    g07149(.A(\A[147] ), .Y(new_n8152_));
  INV    g07150(.A(\A[146] ), .Y(new_n8153_));
  NAND2  g07151(.A(new_n8153_), .B(\A[145] ), .Y(new_n8154_));
  INV    g07152(.A(\A[145] ), .Y(new_n8155_));
  AOI21  g07153(.A0(\A[146] ), .A1(new_n8155_), .B0(new_n8152_), .Y(new_n8156_));
  XOR2   g07154(.A(\A[146] ), .B(\A[145] ), .Y(new_n8157_));
  AOI22  g07155(.A0(new_n8157_), .A1(new_n8152_), .B0(new_n8156_), .B1(new_n8154_), .Y(new_n8158_));
  INV    g07156(.A(\A[150] ), .Y(new_n8159_));
  INV    g07157(.A(\A[149] ), .Y(new_n8160_));
  NAND2  g07158(.A(new_n8160_), .B(\A[148] ), .Y(new_n8161_));
  INV    g07159(.A(\A[148] ), .Y(new_n8162_));
  AOI21  g07160(.A0(\A[149] ), .A1(new_n8162_), .B0(new_n8159_), .Y(new_n8163_));
  XOR2   g07161(.A(\A[149] ), .B(\A[148] ), .Y(new_n8164_));
  AOI22  g07162(.A0(new_n8164_), .A1(new_n8159_), .B0(new_n8163_), .B1(new_n8161_), .Y(new_n8165_));
  NOR2   g07163(.A(new_n8160_), .B(new_n8162_), .Y(new_n8166_));
  AOI21  g07164(.A0(new_n8164_), .A1(\A[150] ), .B0(new_n8166_), .Y(new_n8167_));
  NOR2   g07165(.A(new_n8153_), .B(new_n8155_), .Y(new_n8168_));
  AOI21  g07166(.A0(new_n8157_), .A1(\A[147] ), .B0(new_n8168_), .Y(new_n8169_));
  XOR2   g07167(.A(new_n8165_), .B(new_n8158_), .Y(new_n8170_));
  INV    g07168(.A(\A[141] ), .Y(new_n8171_));
  INV    g07169(.A(\A[140] ), .Y(new_n8172_));
  NAND2  g07170(.A(new_n8172_), .B(\A[139] ), .Y(new_n8173_));
  INV    g07171(.A(\A[139] ), .Y(new_n8174_));
  AOI21  g07172(.A0(\A[140] ), .A1(new_n8174_), .B0(new_n8171_), .Y(new_n8175_));
  XOR2   g07173(.A(\A[140] ), .B(\A[139] ), .Y(new_n8176_));
  AOI22  g07174(.A0(new_n8176_), .A1(new_n8171_), .B0(new_n8175_), .B1(new_n8173_), .Y(new_n8177_));
  INV    g07175(.A(\A[144] ), .Y(new_n8178_));
  INV    g07176(.A(\A[143] ), .Y(new_n8179_));
  NAND2  g07177(.A(new_n8179_), .B(\A[142] ), .Y(new_n8180_));
  INV    g07178(.A(\A[142] ), .Y(new_n8181_));
  AOI21  g07179(.A0(\A[143] ), .A1(new_n8181_), .B0(new_n8178_), .Y(new_n8182_));
  XOR2   g07180(.A(\A[143] ), .B(\A[142] ), .Y(new_n8183_));
  AOI22  g07181(.A0(new_n8183_), .A1(new_n8178_), .B0(new_n8182_), .B1(new_n8180_), .Y(new_n8184_));
  NOR2   g07182(.A(new_n8179_), .B(new_n8181_), .Y(new_n8185_));
  AOI21  g07183(.A0(new_n8183_), .A1(\A[144] ), .B0(new_n8185_), .Y(new_n8186_));
  NOR2   g07184(.A(new_n8172_), .B(new_n8174_), .Y(new_n8187_));
  AOI21  g07185(.A0(new_n8176_), .A1(\A[141] ), .B0(new_n8187_), .Y(new_n8188_));
  XOR2   g07186(.A(new_n8184_), .B(new_n8177_), .Y(new_n8189_));
  XOR2   g07187(.A(new_n8189_), .B(new_n8170_), .Y(new_n8190_));
  INV    g07188(.A(\A[133] ), .Y(new_n8191_));
  NOR2   g07189(.A(\A[134] ), .B(new_n8191_), .Y(new_n8192_));
  INV    g07190(.A(\A[134] ), .Y(new_n8193_));
  OAI21  g07191(.A0(new_n8193_), .A1(\A[133] ), .B0(\A[135] ), .Y(new_n8194_));
  INV    g07192(.A(\A[135] ), .Y(new_n8195_));
  XOR2   g07193(.A(\A[134] ), .B(\A[133] ), .Y(new_n8196_));
  NAND2  g07194(.A(new_n8196_), .B(new_n8195_), .Y(new_n8197_));
  OAI21  g07195(.A0(new_n8194_), .A1(new_n8192_), .B0(new_n8197_), .Y(new_n8198_));
  INV    g07196(.A(\A[138] ), .Y(new_n8199_));
  INV    g07197(.A(\A[137] ), .Y(new_n8200_));
  NAND2  g07198(.A(new_n8200_), .B(\A[136] ), .Y(new_n8201_));
  INV    g07199(.A(\A[136] ), .Y(new_n8202_));
  AOI21  g07200(.A0(\A[137] ), .A1(new_n8202_), .B0(new_n8199_), .Y(new_n8203_));
  XOR2   g07201(.A(\A[137] ), .B(\A[136] ), .Y(new_n8204_));
  AOI22  g07202(.A0(new_n8204_), .A1(new_n8199_), .B0(new_n8203_), .B1(new_n8201_), .Y(new_n8205_));
  NOR2   g07203(.A(new_n8200_), .B(new_n8202_), .Y(new_n8206_));
  AOI21  g07204(.A0(new_n8204_), .A1(\A[138] ), .B0(new_n8206_), .Y(new_n8207_));
  NOR2   g07205(.A(new_n8193_), .B(new_n8191_), .Y(new_n8208_));
  AOI21  g07206(.A0(new_n8196_), .A1(\A[135] ), .B0(new_n8208_), .Y(new_n8209_));
  XOR2   g07207(.A(new_n8205_), .B(new_n8198_), .Y(new_n8210_));
  INV    g07208(.A(\A[129] ), .Y(new_n8211_));
  INV    g07209(.A(\A[128] ), .Y(new_n8212_));
  NAND2  g07210(.A(new_n8212_), .B(\A[127] ), .Y(new_n8213_));
  INV    g07211(.A(\A[127] ), .Y(new_n8214_));
  AOI21  g07212(.A0(\A[128] ), .A1(new_n8214_), .B0(new_n8211_), .Y(new_n8215_));
  XOR2   g07213(.A(\A[128] ), .B(\A[127] ), .Y(new_n8216_));
  AOI22  g07214(.A0(new_n8216_), .A1(new_n8211_), .B0(new_n8215_), .B1(new_n8213_), .Y(new_n8217_));
  INV    g07215(.A(\A[132] ), .Y(new_n8218_));
  INV    g07216(.A(\A[131] ), .Y(new_n8219_));
  NAND2  g07217(.A(new_n8219_), .B(\A[130] ), .Y(new_n8220_));
  INV    g07218(.A(\A[130] ), .Y(new_n8221_));
  AOI21  g07219(.A0(\A[131] ), .A1(new_n8221_), .B0(new_n8218_), .Y(new_n8222_));
  XOR2   g07220(.A(\A[131] ), .B(\A[130] ), .Y(new_n8223_));
  AOI22  g07221(.A0(new_n8223_), .A1(new_n8218_), .B0(new_n8222_), .B1(new_n8220_), .Y(new_n8224_));
  NOR2   g07222(.A(new_n8219_), .B(new_n8221_), .Y(new_n8225_));
  AOI21  g07223(.A0(new_n8223_), .A1(\A[132] ), .B0(new_n8225_), .Y(new_n8226_));
  NOR2   g07224(.A(new_n8212_), .B(new_n8214_), .Y(new_n8227_));
  AOI21  g07225(.A0(new_n8216_), .A1(\A[129] ), .B0(new_n8227_), .Y(new_n8228_));
  XOR2   g07226(.A(new_n8224_), .B(new_n8217_), .Y(new_n8229_));
  XOR2   g07227(.A(new_n8229_), .B(new_n8210_), .Y(new_n8230_));
  XOR2   g07228(.A(new_n8230_), .B(new_n8190_), .Y(new_n8231_));
  XOR2   g07229(.A(new_n8231_), .B(new_n8151_), .Y(new_n8232_));
  INV    g07230(.A(new_n8232_), .Y(new_n8233_));
  INV    g07231(.A(\A[123] ), .Y(new_n8234_));
  INV    g07232(.A(\A[122] ), .Y(new_n8235_));
  NAND2  g07233(.A(new_n8235_), .B(\A[121] ), .Y(new_n8236_));
  INV    g07234(.A(\A[121] ), .Y(new_n8237_));
  AOI21  g07235(.A0(\A[122] ), .A1(new_n8237_), .B0(new_n8234_), .Y(new_n8238_));
  XOR2   g07236(.A(\A[122] ), .B(\A[121] ), .Y(new_n8239_));
  AOI22  g07237(.A0(new_n8239_), .A1(new_n8234_), .B0(new_n8238_), .B1(new_n8236_), .Y(new_n8240_));
  INV    g07238(.A(\A[126] ), .Y(new_n8241_));
  INV    g07239(.A(\A[125] ), .Y(new_n8242_));
  NAND2  g07240(.A(new_n8242_), .B(\A[124] ), .Y(new_n8243_));
  INV    g07241(.A(\A[124] ), .Y(new_n8244_));
  AOI21  g07242(.A0(\A[125] ), .A1(new_n8244_), .B0(new_n8241_), .Y(new_n8245_));
  XOR2   g07243(.A(\A[125] ), .B(\A[124] ), .Y(new_n8246_));
  AOI22  g07244(.A0(new_n8246_), .A1(new_n8241_), .B0(new_n8245_), .B1(new_n8243_), .Y(new_n8247_));
  NOR2   g07245(.A(new_n8242_), .B(new_n8244_), .Y(new_n8248_));
  AOI21  g07246(.A0(new_n8246_), .A1(\A[126] ), .B0(new_n8248_), .Y(new_n8249_));
  NOR2   g07247(.A(new_n8235_), .B(new_n8237_), .Y(new_n8250_));
  AOI21  g07248(.A0(new_n8239_), .A1(\A[123] ), .B0(new_n8250_), .Y(new_n8251_));
  XOR2   g07249(.A(new_n8247_), .B(new_n8240_), .Y(new_n8252_));
  INV    g07250(.A(\A[117] ), .Y(new_n8253_));
  INV    g07251(.A(\A[116] ), .Y(new_n8254_));
  NAND2  g07252(.A(new_n8254_), .B(\A[115] ), .Y(new_n8255_));
  INV    g07253(.A(\A[115] ), .Y(new_n8256_));
  AOI21  g07254(.A0(\A[116] ), .A1(new_n8256_), .B0(new_n8253_), .Y(new_n8257_));
  XOR2   g07255(.A(\A[116] ), .B(\A[115] ), .Y(new_n8258_));
  AOI22  g07256(.A0(new_n8258_), .A1(new_n8253_), .B0(new_n8257_), .B1(new_n8255_), .Y(new_n8259_));
  INV    g07257(.A(\A[120] ), .Y(new_n8260_));
  INV    g07258(.A(\A[119] ), .Y(new_n8261_));
  NAND2  g07259(.A(new_n8261_), .B(\A[118] ), .Y(new_n8262_));
  INV    g07260(.A(\A[118] ), .Y(new_n8263_));
  AOI21  g07261(.A0(\A[119] ), .A1(new_n8263_), .B0(new_n8260_), .Y(new_n8264_));
  XOR2   g07262(.A(\A[119] ), .B(\A[118] ), .Y(new_n8265_));
  AOI22  g07263(.A0(new_n8265_), .A1(new_n8260_), .B0(new_n8264_), .B1(new_n8262_), .Y(new_n8266_));
  NOR2   g07264(.A(new_n8261_), .B(new_n8263_), .Y(new_n8267_));
  AOI21  g07265(.A0(new_n8265_), .A1(\A[120] ), .B0(new_n8267_), .Y(new_n8268_));
  NOR2   g07266(.A(new_n8254_), .B(new_n8256_), .Y(new_n8269_));
  AOI21  g07267(.A0(new_n8258_), .A1(\A[117] ), .B0(new_n8269_), .Y(new_n8270_));
  XOR2   g07268(.A(new_n8266_), .B(new_n8259_), .Y(new_n8271_));
  XOR2   g07269(.A(new_n8271_), .B(new_n8252_), .Y(new_n8272_));
  INV    g07270(.A(\A[109] ), .Y(new_n8273_));
  NOR2   g07271(.A(\A[110] ), .B(new_n8273_), .Y(new_n8274_));
  INV    g07272(.A(\A[110] ), .Y(new_n8275_));
  OAI21  g07273(.A0(new_n8275_), .A1(\A[109] ), .B0(\A[111] ), .Y(new_n8276_));
  INV    g07274(.A(\A[111] ), .Y(new_n8277_));
  XOR2   g07275(.A(\A[110] ), .B(\A[109] ), .Y(new_n8278_));
  NAND2  g07276(.A(new_n8278_), .B(new_n8277_), .Y(new_n8279_));
  OAI21  g07277(.A0(new_n8276_), .A1(new_n8274_), .B0(new_n8279_), .Y(new_n8280_));
  INV    g07278(.A(\A[114] ), .Y(new_n8281_));
  INV    g07279(.A(\A[113] ), .Y(new_n8282_));
  NAND2  g07280(.A(new_n8282_), .B(\A[112] ), .Y(new_n8283_));
  INV    g07281(.A(\A[112] ), .Y(new_n8284_));
  AOI21  g07282(.A0(\A[113] ), .A1(new_n8284_), .B0(new_n8281_), .Y(new_n8285_));
  XOR2   g07283(.A(\A[113] ), .B(\A[112] ), .Y(new_n8286_));
  AOI22  g07284(.A0(new_n8286_), .A1(new_n8281_), .B0(new_n8285_), .B1(new_n8283_), .Y(new_n8287_));
  NOR2   g07285(.A(new_n8282_), .B(new_n8284_), .Y(new_n8288_));
  AOI21  g07286(.A0(new_n8286_), .A1(\A[114] ), .B0(new_n8288_), .Y(new_n8289_));
  NOR2   g07287(.A(new_n8275_), .B(new_n8273_), .Y(new_n8290_));
  AOI21  g07288(.A0(new_n8278_), .A1(\A[111] ), .B0(new_n8290_), .Y(new_n8291_));
  XOR2   g07289(.A(new_n8287_), .B(new_n8280_), .Y(new_n8292_));
  INV    g07290(.A(\A[105] ), .Y(new_n8293_));
  INV    g07291(.A(\A[104] ), .Y(new_n8294_));
  NAND2  g07292(.A(new_n8294_), .B(\A[103] ), .Y(new_n8295_));
  INV    g07293(.A(\A[103] ), .Y(new_n8296_));
  AOI21  g07294(.A0(\A[104] ), .A1(new_n8296_), .B0(new_n8293_), .Y(new_n8297_));
  XOR2   g07295(.A(\A[104] ), .B(\A[103] ), .Y(new_n8298_));
  AOI22  g07296(.A0(new_n8298_), .A1(new_n8293_), .B0(new_n8297_), .B1(new_n8295_), .Y(new_n8299_));
  INV    g07297(.A(\A[108] ), .Y(new_n8300_));
  INV    g07298(.A(\A[107] ), .Y(new_n8301_));
  NAND2  g07299(.A(new_n8301_), .B(\A[106] ), .Y(new_n8302_));
  INV    g07300(.A(\A[106] ), .Y(new_n8303_));
  AOI21  g07301(.A0(\A[107] ), .A1(new_n8303_), .B0(new_n8300_), .Y(new_n8304_));
  XOR2   g07302(.A(\A[107] ), .B(\A[106] ), .Y(new_n8305_));
  AOI22  g07303(.A0(new_n8305_), .A1(new_n8300_), .B0(new_n8304_), .B1(new_n8302_), .Y(new_n8306_));
  NOR2   g07304(.A(new_n8301_), .B(new_n8303_), .Y(new_n8307_));
  AOI21  g07305(.A0(new_n8305_), .A1(\A[108] ), .B0(new_n8307_), .Y(new_n8308_));
  NOR2   g07306(.A(new_n8294_), .B(new_n8296_), .Y(new_n8309_));
  AOI21  g07307(.A0(new_n8298_), .A1(\A[105] ), .B0(new_n8309_), .Y(new_n8310_));
  XOR2   g07308(.A(new_n8306_), .B(new_n8299_), .Y(new_n8311_));
  XOR2   g07309(.A(new_n8311_), .B(new_n8292_), .Y(new_n8312_));
  XOR2   g07310(.A(new_n8312_), .B(new_n8272_), .Y(new_n8313_));
  INV    g07311(.A(new_n8313_), .Y(new_n8314_));
  INV    g07312(.A(\A[99] ), .Y(new_n8315_));
  INV    g07313(.A(\A[98] ), .Y(new_n8316_));
  NAND2  g07314(.A(new_n8316_), .B(\A[97] ), .Y(new_n8317_));
  INV    g07315(.A(\A[97] ), .Y(new_n8318_));
  AOI21  g07316(.A0(\A[98] ), .A1(new_n8318_), .B0(new_n8315_), .Y(new_n8319_));
  XOR2   g07317(.A(\A[98] ), .B(\A[97] ), .Y(new_n8320_));
  AOI22  g07318(.A0(new_n8320_), .A1(new_n8315_), .B0(new_n8319_), .B1(new_n8317_), .Y(new_n8321_));
  INV    g07319(.A(\A[102] ), .Y(new_n8322_));
  INV    g07320(.A(\A[101] ), .Y(new_n8323_));
  NAND2  g07321(.A(new_n8323_), .B(\A[100] ), .Y(new_n8324_));
  INV    g07322(.A(\A[100] ), .Y(new_n8325_));
  AOI21  g07323(.A0(\A[101] ), .A1(new_n8325_), .B0(new_n8322_), .Y(new_n8326_));
  XOR2   g07324(.A(\A[101] ), .B(\A[100] ), .Y(new_n8327_));
  AOI22  g07325(.A0(new_n8327_), .A1(new_n8322_), .B0(new_n8326_), .B1(new_n8324_), .Y(new_n8328_));
  NOR2   g07326(.A(new_n8323_), .B(new_n8325_), .Y(new_n8329_));
  AOI21  g07327(.A0(new_n8327_), .A1(\A[102] ), .B0(new_n8329_), .Y(new_n8330_));
  NOR2   g07328(.A(new_n8316_), .B(new_n8318_), .Y(new_n8331_));
  AOI21  g07329(.A0(new_n8320_), .A1(\A[99] ), .B0(new_n8331_), .Y(new_n8332_));
  XOR2   g07330(.A(new_n8328_), .B(new_n8321_), .Y(new_n8333_));
  INV    g07331(.A(\A[93] ), .Y(new_n8334_));
  INV    g07332(.A(\A[92] ), .Y(new_n8335_));
  NAND2  g07333(.A(new_n8335_), .B(\A[91] ), .Y(new_n8336_));
  INV    g07334(.A(\A[91] ), .Y(new_n8337_));
  AOI21  g07335(.A0(\A[92] ), .A1(new_n8337_), .B0(new_n8334_), .Y(new_n8338_));
  XOR2   g07336(.A(\A[92] ), .B(\A[91] ), .Y(new_n8339_));
  AOI22  g07337(.A0(new_n8339_), .A1(new_n8334_), .B0(new_n8338_), .B1(new_n8336_), .Y(new_n8340_));
  INV    g07338(.A(\A[96] ), .Y(new_n8341_));
  INV    g07339(.A(\A[95] ), .Y(new_n8342_));
  NAND2  g07340(.A(new_n8342_), .B(\A[94] ), .Y(new_n8343_));
  INV    g07341(.A(\A[94] ), .Y(new_n8344_));
  AOI21  g07342(.A0(\A[95] ), .A1(new_n8344_), .B0(new_n8341_), .Y(new_n8345_));
  XOR2   g07343(.A(\A[95] ), .B(\A[94] ), .Y(new_n8346_));
  AOI22  g07344(.A0(new_n8346_), .A1(new_n8341_), .B0(new_n8345_), .B1(new_n8343_), .Y(new_n8347_));
  NOR2   g07345(.A(new_n8342_), .B(new_n8344_), .Y(new_n8348_));
  AOI21  g07346(.A0(new_n8346_), .A1(\A[96] ), .B0(new_n8348_), .Y(new_n8349_));
  NOR2   g07347(.A(new_n8335_), .B(new_n8337_), .Y(new_n8350_));
  AOI21  g07348(.A0(new_n8339_), .A1(\A[93] ), .B0(new_n8350_), .Y(new_n8351_));
  XOR2   g07349(.A(new_n8347_), .B(new_n8340_), .Y(new_n8352_));
  XOR2   g07350(.A(new_n8352_), .B(new_n8333_), .Y(new_n8353_));
  INV    g07351(.A(\A[85] ), .Y(new_n8354_));
  NOR2   g07352(.A(\A[86] ), .B(new_n8354_), .Y(new_n8355_));
  INV    g07353(.A(\A[86] ), .Y(new_n8356_));
  OAI21  g07354(.A0(new_n8356_), .A1(\A[85] ), .B0(\A[87] ), .Y(new_n8357_));
  INV    g07355(.A(\A[87] ), .Y(new_n8358_));
  XOR2   g07356(.A(\A[86] ), .B(\A[85] ), .Y(new_n8359_));
  NAND2  g07357(.A(new_n8359_), .B(new_n8358_), .Y(new_n8360_));
  OAI21  g07358(.A0(new_n8357_), .A1(new_n8355_), .B0(new_n8360_), .Y(new_n8361_));
  INV    g07359(.A(\A[90] ), .Y(new_n8362_));
  INV    g07360(.A(\A[89] ), .Y(new_n8363_));
  NAND2  g07361(.A(new_n8363_), .B(\A[88] ), .Y(new_n8364_));
  INV    g07362(.A(\A[88] ), .Y(new_n8365_));
  AOI21  g07363(.A0(\A[89] ), .A1(new_n8365_), .B0(new_n8362_), .Y(new_n8366_));
  XOR2   g07364(.A(\A[89] ), .B(\A[88] ), .Y(new_n8367_));
  AOI22  g07365(.A0(new_n8367_), .A1(new_n8362_), .B0(new_n8366_), .B1(new_n8364_), .Y(new_n8368_));
  NOR2   g07366(.A(new_n8363_), .B(new_n8365_), .Y(new_n8369_));
  AOI21  g07367(.A0(new_n8367_), .A1(\A[90] ), .B0(new_n8369_), .Y(new_n8370_));
  NOR2   g07368(.A(new_n8356_), .B(new_n8354_), .Y(new_n8371_));
  AOI21  g07369(.A0(new_n8359_), .A1(\A[87] ), .B0(new_n8371_), .Y(new_n8372_));
  XOR2   g07370(.A(new_n8368_), .B(new_n8361_), .Y(new_n8373_));
  INV    g07371(.A(\A[81] ), .Y(new_n8374_));
  INV    g07372(.A(\A[80] ), .Y(new_n8375_));
  NAND2  g07373(.A(new_n8375_), .B(\A[79] ), .Y(new_n8376_));
  INV    g07374(.A(\A[79] ), .Y(new_n8377_));
  AOI21  g07375(.A0(\A[80] ), .A1(new_n8377_), .B0(new_n8374_), .Y(new_n8378_));
  XOR2   g07376(.A(\A[80] ), .B(\A[79] ), .Y(new_n8379_));
  AOI22  g07377(.A0(new_n8379_), .A1(new_n8374_), .B0(new_n8378_), .B1(new_n8376_), .Y(new_n8380_));
  INV    g07378(.A(\A[84] ), .Y(new_n8381_));
  INV    g07379(.A(\A[83] ), .Y(new_n8382_));
  NAND2  g07380(.A(new_n8382_), .B(\A[82] ), .Y(new_n8383_));
  INV    g07381(.A(\A[82] ), .Y(new_n8384_));
  AOI21  g07382(.A0(\A[83] ), .A1(new_n8384_), .B0(new_n8381_), .Y(new_n8385_));
  XOR2   g07383(.A(\A[83] ), .B(\A[82] ), .Y(new_n8386_));
  AOI22  g07384(.A0(new_n8386_), .A1(new_n8381_), .B0(new_n8385_), .B1(new_n8383_), .Y(new_n8387_));
  NOR2   g07385(.A(new_n8382_), .B(new_n8384_), .Y(new_n8388_));
  AOI21  g07386(.A0(new_n8386_), .A1(\A[84] ), .B0(new_n8388_), .Y(new_n8389_));
  NOR2   g07387(.A(new_n8375_), .B(new_n8377_), .Y(new_n8390_));
  AOI21  g07388(.A0(new_n8379_), .A1(\A[81] ), .B0(new_n8390_), .Y(new_n8391_));
  XOR2   g07389(.A(new_n8387_), .B(new_n8380_), .Y(new_n8392_));
  XOR2   g07390(.A(new_n8392_), .B(new_n8373_), .Y(new_n8393_));
  XOR2   g07391(.A(new_n8393_), .B(new_n8353_), .Y(new_n8394_));
  XOR2   g07392(.A(new_n8394_), .B(new_n8314_), .Y(new_n8395_));
  XOR2   g07393(.A(new_n8395_), .B(new_n8233_), .Y(new_n8396_));
  NOR2   g07394(.A(new_n8396_), .B(new_n8070_), .Y(new_n8397_));
  NAND3  g07395(.A(new_n8397_), .B(new_n8069_), .C(new_n8059_), .Y(new_n8398_));
  NAND3  g07396(.A(new_n8049_), .B(new_n8057_), .C(new_n8054_), .Y(new_n8399_));
  OAI21  g07397(.A0(new_n8044_), .A1(new_n8036_), .B0(new_n8050_), .Y(new_n8400_));
  AOI21  g07398(.A0(new_n8400_), .A1(new_n8399_), .B0(new_n8066_), .Y(new_n8401_));
  NAND3  g07399(.A(new_n8050_), .B(new_n8057_), .C(new_n8054_), .Y(new_n8402_));
  OAI21  g07400(.A0(new_n8044_), .A1(new_n8036_), .B0(new_n8049_), .Y(new_n8403_));
  AOI21  g07401(.A0(new_n8403_), .A1(new_n8402_), .B0(new_n7547_), .Y(new_n8404_));
  INV    g07402(.A(new_n8397_), .Y(new_n8405_));
  OAI21  g07403(.A0(new_n8404_), .A1(new_n8401_), .B0(new_n8405_), .Y(new_n8406_));
  XOR2   g07404(.A(new_n8184_), .B(new_n8177_), .Y(new_n8407_));
  XOR2   g07405(.A(\A[143] ), .B(new_n8181_), .Y(new_n8408_));
  NAND2  g07406(.A(\A[143] ), .B(\A[142] ), .Y(new_n8409_));
  OAI21  g07407(.A0(new_n8408_), .A1(new_n8178_), .B0(new_n8409_), .Y(new_n8410_));
  XOR2   g07408(.A(new_n8188_), .B(new_n8410_), .Y(new_n8411_));
  NOR2   g07409(.A(\A[140] ), .B(new_n8174_), .Y(new_n8412_));
  OAI21  g07410(.A0(new_n8172_), .A1(\A[139] ), .B0(\A[141] ), .Y(new_n8413_));
  XOR2   g07411(.A(\A[140] ), .B(new_n8174_), .Y(new_n8414_));
  OAI22  g07412(.A0(new_n8414_), .A1(\A[141] ), .B0(new_n8413_), .B1(new_n8412_), .Y(new_n8415_));
  NOR2   g07413(.A(\A[143] ), .B(new_n8181_), .Y(new_n8416_));
  OAI21  g07414(.A0(new_n8179_), .A1(\A[142] ), .B0(\A[144] ), .Y(new_n8417_));
  OAI22  g07415(.A0(new_n8408_), .A1(\A[144] ), .B0(new_n8417_), .B1(new_n8416_), .Y(new_n8418_));
  NAND2  g07416(.A(new_n8418_), .B(new_n8415_), .Y(new_n8419_));
  NAND2  g07417(.A(\A[140] ), .B(\A[139] ), .Y(new_n8420_));
  OAI21  g07418(.A0(new_n8414_), .A1(new_n8171_), .B0(new_n8420_), .Y(new_n8421_));
  NAND2  g07419(.A(new_n8421_), .B(new_n8410_), .Y(new_n8422_));
  OAI21  g07420(.A0(new_n8419_), .A1(new_n8411_), .B0(new_n8422_), .Y(new_n8423_));
  NOR2   g07421(.A(new_n8184_), .B(new_n8177_), .Y(new_n8424_));
  XOR2   g07422(.A(new_n8424_), .B(new_n8411_), .Y(new_n8425_));
  AOI21  g07423(.A0(new_n8423_), .A1(new_n8407_), .B0(new_n8425_), .Y(new_n8426_));
  NOR2   g07424(.A(\A[146] ), .B(new_n8155_), .Y(new_n8427_));
  OAI21  g07425(.A0(new_n8153_), .A1(\A[145] ), .B0(\A[147] ), .Y(new_n8428_));
  NAND2  g07426(.A(new_n8157_), .B(new_n8152_), .Y(new_n8429_));
  OAI21  g07427(.A0(new_n8428_), .A1(new_n8427_), .B0(new_n8429_), .Y(new_n8430_));
  XOR2   g07428(.A(new_n8165_), .B(new_n8430_), .Y(new_n8431_));
  XOR2   g07429(.A(new_n8169_), .B(new_n8167_), .Y(new_n8432_));
  NOR2   g07430(.A(new_n8165_), .B(new_n8158_), .Y(new_n8433_));
  NAND2  g07431(.A(\A[149] ), .B(\A[148] ), .Y(new_n8434_));
  NAND2  g07432(.A(new_n8164_), .B(\A[150] ), .Y(new_n8435_));
  NAND2  g07433(.A(\A[146] ), .B(\A[145] ), .Y(new_n8436_));
  NAND2  g07434(.A(new_n8157_), .B(\A[147] ), .Y(new_n8437_));
  AOI22  g07435(.A0(new_n8437_), .A1(new_n8436_), .B0(new_n8435_), .B1(new_n8434_), .Y(new_n8438_));
  AOI21  g07436(.A0(new_n8433_), .A1(new_n8432_), .B0(new_n8438_), .Y(new_n8439_));
  XOR2   g07437(.A(new_n8433_), .B(new_n8432_), .Y(new_n8440_));
  XOR2   g07438(.A(new_n8165_), .B(new_n8158_), .Y(new_n8441_));
  NOR2   g07439(.A(\A[149] ), .B(new_n8162_), .Y(new_n8442_));
  OAI21  g07440(.A0(new_n8160_), .A1(\A[148] ), .B0(\A[150] ), .Y(new_n8443_));
  NAND2  g07441(.A(new_n8164_), .B(new_n8159_), .Y(new_n8444_));
  OAI21  g07442(.A0(new_n8443_), .A1(new_n8442_), .B0(new_n8444_), .Y(new_n8445_));
  NAND2  g07443(.A(new_n8435_), .B(new_n8434_), .Y(new_n8446_));
  NAND2  g07444(.A(new_n8437_), .B(new_n8436_), .Y(new_n8447_));
  NAND4  g07445(.A(new_n8447_), .B(new_n8446_), .C(new_n8445_), .D(new_n8430_), .Y(new_n8448_));
  NAND4  g07446(.A(new_n8421_), .B(new_n8410_), .C(new_n8418_), .D(new_n8415_), .Y(new_n8449_));
  NAND4  g07447(.A(new_n8449_), .B(new_n8407_), .C(new_n8448_), .D(new_n8441_), .Y(new_n8450_));
  OAI211 g07448(.A0(new_n8439_), .A1(new_n8431_), .B0(new_n8450_), .B1(new_n8440_), .Y(new_n8451_));
  XOR2   g07449(.A(new_n8169_), .B(new_n8446_), .Y(new_n8452_));
  XOR2   g07450(.A(new_n8433_), .B(new_n8452_), .Y(new_n8453_));
  NOR4   g07451(.A(new_n8169_), .B(new_n8167_), .C(new_n8165_), .D(new_n8158_), .Y(new_n8454_));
  XOR2   g07452(.A(new_n8184_), .B(new_n8415_), .Y(new_n8455_));
  NOR4   g07453(.A(new_n8188_), .B(new_n8186_), .C(new_n8184_), .D(new_n8177_), .Y(new_n8456_));
  NOR4   g07454(.A(new_n8456_), .B(new_n8455_), .C(new_n8454_), .D(new_n8431_), .Y(new_n8457_));
  AOI221 g07455(.A0(new_n8435_), .A1(new_n8434_), .C0(new_n8168_), .B0(new_n8157_), .B1(\A[147] ), .Y(new_n8458_));
  AOI221 g07456(.A0(new_n8437_), .A1(new_n8436_), .C0(new_n8166_), .B0(new_n8164_), .B1(\A[150] ), .Y(new_n8459_));
  OAI211 g07457(.A0(new_n8459_), .A1(new_n8458_), .B0(new_n8445_), .B1(new_n8430_), .Y(new_n8460_));
  NAND2  g07458(.A(new_n8447_), .B(new_n8446_), .Y(new_n8461_));
  AOI21  g07459(.A0(new_n8461_), .A1(new_n8460_), .B0(new_n8431_), .Y(new_n8462_));
  OAI21  g07460(.A0(new_n8462_), .A1(new_n8453_), .B0(new_n8457_), .Y(new_n8463_));
  AOI21  g07461(.A0(new_n8463_), .A1(new_n8451_), .B0(new_n8426_), .Y(new_n8464_));
  OAI21  g07462(.A0(new_n8462_), .A1(new_n8453_), .B0(new_n8450_), .Y(new_n8465_));
  NAND4  g07463(.A(new_n8407_), .B(new_n8440_), .C(new_n8439_), .D(new_n8441_), .Y(new_n8466_));
  OAI21  g07464(.A0(new_n8439_), .A1(new_n8431_), .B0(new_n8449_), .Y(new_n8467_));
  OAI21  g07465(.A0(new_n8467_), .A1(new_n8466_), .B0(new_n8465_), .Y(new_n8468_));
  NAND2  g07466(.A(new_n8193_), .B(\A[133] ), .Y(new_n8469_));
  AOI21  g07467(.A0(\A[134] ), .A1(new_n8191_), .B0(new_n8195_), .Y(new_n8470_));
  AOI22  g07468(.A0(new_n8196_), .A1(new_n8195_), .B0(new_n8470_), .B1(new_n8469_), .Y(new_n8471_));
  XOR2   g07469(.A(new_n8205_), .B(new_n8471_), .Y(new_n8472_));
  XOR2   g07470(.A(new_n8229_), .B(new_n8472_), .Y(new_n8473_));
  NAND2  g07471(.A(new_n8473_), .B(new_n8190_), .Y(new_n8474_));
  AOI211 g07472(.A0(new_n8468_), .A1(new_n8426_), .B(new_n8474_), .C(new_n8464_), .Y(new_n8475_));
  XOR2   g07473(.A(new_n8165_), .B(new_n8430_), .Y(new_n8476_));
  XOR2   g07474(.A(new_n8189_), .B(new_n8476_), .Y(new_n8477_));
  NOR2   g07475(.A(new_n8230_), .B(new_n8477_), .Y(new_n8478_));
  AOI21  g07476(.A0(new_n8468_), .A1(new_n8426_), .B0(new_n8464_), .Y(new_n8479_));
  NOR2   g07477(.A(new_n8479_), .B(new_n8478_), .Y(new_n8480_));
  XOR2   g07478(.A(new_n8224_), .B(new_n8217_), .Y(new_n8481_));
  XOR2   g07479(.A(\A[131] ), .B(new_n8221_), .Y(new_n8482_));
  NAND2  g07480(.A(\A[131] ), .B(\A[130] ), .Y(new_n8483_));
  OAI21  g07481(.A0(new_n8482_), .A1(new_n8218_), .B0(new_n8483_), .Y(new_n8484_));
  XOR2   g07482(.A(new_n8228_), .B(new_n8484_), .Y(new_n8485_));
  NOR2   g07483(.A(\A[128] ), .B(new_n8214_), .Y(new_n8486_));
  OAI21  g07484(.A0(new_n8212_), .A1(\A[127] ), .B0(\A[129] ), .Y(new_n8487_));
  XOR2   g07485(.A(\A[128] ), .B(new_n8214_), .Y(new_n8488_));
  OAI22  g07486(.A0(new_n8488_), .A1(\A[129] ), .B0(new_n8487_), .B1(new_n8486_), .Y(new_n8489_));
  NOR2   g07487(.A(\A[131] ), .B(new_n8221_), .Y(new_n8490_));
  OAI21  g07488(.A0(new_n8219_), .A1(\A[130] ), .B0(\A[132] ), .Y(new_n8491_));
  OAI22  g07489(.A0(new_n8482_), .A1(\A[132] ), .B0(new_n8491_), .B1(new_n8490_), .Y(new_n8492_));
  NAND2  g07490(.A(new_n8492_), .B(new_n8489_), .Y(new_n8493_));
  NAND2  g07491(.A(\A[128] ), .B(\A[127] ), .Y(new_n8494_));
  OAI21  g07492(.A0(new_n8488_), .A1(new_n8211_), .B0(new_n8494_), .Y(new_n8495_));
  NAND2  g07493(.A(new_n8495_), .B(new_n8484_), .Y(new_n8496_));
  OAI21  g07494(.A0(new_n8493_), .A1(new_n8485_), .B0(new_n8496_), .Y(new_n8497_));
  NOR2   g07495(.A(new_n8224_), .B(new_n8217_), .Y(new_n8498_));
  XOR2   g07496(.A(new_n8498_), .B(new_n8485_), .Y(new_n8499_));
  AOI21  g07497(.A0(new_n8497_), .A1(new_n8481_), .B0(new_n8499_), .Y(new_n8500_));
  XOR2   g07498(.A(new_n8205_), .B(new_n8198_), .Y(new_n8501_));
  XOR2   g07499(.A(new_n8209_), .B(new_n8207_), .Y(new_n8502_));
  NOR2   g07500(.A(new_n8205_), .B(new_n8471_), .Y(new_n8503_));
  NAND2  g07501(.A(\A[137] ), .B(\A[136] ), .Y(new_n8504_));
  NAND2  g07502(.A(new_n8204_), .B(\A[138] ), .Y(new_n8505_));
  NAND2  g07503(.A(\A[134] ), .B(\A[133] ), .Y(new_n8506_));
  NAND2  g07504(.A(new_n8196_), .B(\A[135] ), .Y(new_n8507_));
  AOI22  g07505(.A0(new_n8507_), .A1(new_n8506_), .B0(new_n8505_), .B1(new_n8504_), .Y(new_n8508_));
  AOI21  g07506(.A0(new_n8503_), .A1(new_n8502_), .B0(new_n8508_), .Y(new_n8509_));
  XOR2   g07507(.A(new_n8503_), .B(new_n8502_), .Y(new_n8510_));
  XOR2   g07508(.A(new_n8205_), .B(new_n8471_), .Y(new_n8511_));
  NOR2   g07509(.A(\A[137] ), .B(new_n8202_), .Y(new_n8512_));
  OAI21  g07510(.A0(new_n8200_), .A1(\A[136] ), .B0(\A[138] ), .Y(new_n8513_));
  NAND2  g07511(.A(new_n8204_), .B(new_n8199_), .Y(new_n8514_));
  OAI21  g07512(.A0(new_n8513_), .A1(new_n8512_), .B0(new_n8514_), .Y(new_n8515_));
  NAND2  g07513(.A(new_n8505_), .B(new_n8504_), .Y(new_n8516_));
  NAND2  g07514(.A(new_n8507_), .B(new_n8506_), .Y(new_n8517_));
  NAND4  g07515(.A(new_n8517_), .B(new_n8516_), .C(new_n8515_), .D(new_n8198_), .Y(new_n8518_));
  NAND4  g07516(.A(new_n8495_), .B(new_n8484_), .C(new_n8492_), .D(new_n8489_), .Y(new_n8519_));
  NAND4  g07517(.A(new_n8519_), .B(new_n8481_), .C(new_n8518_), .D(new_n8511_), .Y(new_n8520_));
  OAI211 g07518(.A0(new_n8509_), .A1(new_n8501_), .B0(new_n8520_), .B1(new_n8510_), .Y(new_n8521_));
  XOR2   g07519(.A(new_n8209_), .B(new_n8516_), .Y(new_n8522_));
  XOR2   g07520(.A(new_n8503_), .B(new_n8522_), .Y(new_n8523_));
  NOR4   g07521(.A(new_n8209_), .B(new_n8207_), .C(new_n8205_), .D(new_n8471_), .Y(new_n8524_));
  XOR2   g07522(.A(new_n8224_), .B(new_n8489_), .Y(new_n8525_));
  NOR3   g07523(.A(new_n8525_), .B(new_n8524_), .C(new_n8501_), .Y(new_n8526_));
  AOI221 g07524(.A0(new_n8505_), .A1(new_n8504_), .C0(new_n8208_), .B0(new_n8196_), .B1(\A[135] ), .Y(new_n8527_));
  AOI221 g07525(.A0(new_n8507_), .A1(new_n8506_), .C0(new_n8206_), .B0(new_n8204_), .B1(\A[138] ), .Y(new_n8528_));
  OAI211 g07526(.A0(new_n8528_), .A1(new_n8527_), .B0(new_n8515_), .B1(new_n8198_), .Y(new_n8529_));
  NAND2  g07527(.A(new_n8517_), .B(new_n8516_), .Y(new_n8530_));
  AOI21  g07528(.A0(new_n8530_), .A1(new_n8529_), .B0(new_n8501_), .Y(new_n8531_));
  OAI211 g07529(.A0(new_n8531_), .A1(new_n8523_), .B0(new_n8526_), .B1(new_n8519_), .Y(new_n8532_));
  AOI21  g07530(.A0(new_n8532_), .A1(new_n8521_), .B0(new_n8500_), .Y(new_n8533_));
  OAI21  g07531(.A0(new_n8531_), .A1(new_n8523_), .B0(new_n8520_), .Y(new_n8534_));
  NAND4  g07532(.A(new_n8481_), .B(new_n8510_), .C(new_n8509_), .D(new_n8511_), .Y(new_n8535_));
  OAI21  g07533(.A0(new_n8509_), .A1(new_n8501_), .B0(new_n8519_), .Y(new_n8536_));
  OAI21  g07534(.A0(new_n8536_), .A1(new_n8535_), .B0(new_n8534_), .Y(new_n8537_));
  AOI21  g07535(.A0(new_n8537_), .A1(new_n8500_), .B0(new_n8533_), .Y(new_n8538_));
  OAI21  g07536(.A0(new_n8480_), .A1(new_n8475_), .B0(new_n8538_), .Y(new_n8539_));
  XOR2   g07537(.A(new_n8228_), .B(new_n8226_), .Y(new_n8540_));
  NOR2   g07538(.A(new_n8228_), .B(new_n8226_), .Y(new_n8541_));
  AOI21  g07539(.A0(new_n8498_), .A1(new_n8540_), .B0(new_n8541_), .Y(new_n8542_));
  XOR2   g07540(.A(new_n8498_), .B(new_n8540_), .Y(new_n8543_));
  OAI21  g07541(.A0(new_n8542_), .A1(new_n8525_), .B0(new_n8543_), .Y(new_n8544_));
  OAI21  g07542(.A0(new_n8509_), .A1(new_n8501_), .B0(new_n8510_), .Y(new_n8545_));
  XOR2   g07543(.A(new_n8545_), .B(new_n8520_), .Y(new_n8546_));
  NAND2  g07544(.A(new_n8546_), .B(new_n8544_), .Y(new_n8547_));
  NAND2  g07545(.A(new_n8537_), .B(new_n8500_), .Y(new_n8548_));
  NAND2  g07546(.A(new_n8548_), .B(new_n8547_), .Y(new_n8549_));
  XOR2   g07547(.A(new_n8188_), .B(new_n8186_), .Y(new_n8550_));
  NOR2   g07548(.A(new_n8188_), .B(new_n8186_), .Y(new_n8551_));
  AOI21  g07549(.A0(new_n8424_), .A1(new_n8550_), .B0(new_n8551_), .Y(new_n8552_));
  XOR2   g07550(.A(new_n8424_), .B(new_n8550_), .Y(new_n8553_));
  OAI21  g07551(.A0(new_n8552_), .A1(new_n8455_), .B0(new_n8553_), .Y(new_n8554_));
  OAI21  g07552(.A0(new_n8439_), .A1(new_n8431_), .B0(new_n8440_), .Y(new_n8555_));
  NAND2  g07553(.A(new_n8461_), .B(new_n8460_), .Y(new_n8556_));
  NOR4   g07554(.A(new_n8455_), .B(new_n8453_), .C(new_n8556_), .D(new_n8431_), .Y(new_n8557_));
  NOR2   g07555(.A(new_n8462_), .B(new_n8456_), .Y(new_n8558_));
  AOI22  g07556(.A0(new_n8558_), .A1(new_n8557_), .B0(new_n8555_), .B1(new_n8450_), .Y(new_n8559_));
  OAI21  g07557(.A0(new_n8559_), .A1(new_n8554_), .B0(new_n8474_), .Y(new_n8560_));
  OAI22  g07558(.A0(new_n8560_), .A1(new_n8464_), .B0(new_n8479_), .B1(new_n8474_), .Y(new_n8561_));
  NAND2  g07559(.A(new_n8561_), .B(new_n8549_), .Y(new_n8562_));
  NAND2  g07560(.A(new_n8562_), .B(new_n8539_), .Y(new_n8563_));
  XOR2   g07561(.A(new_n8143_), .B(new_n8136_), .Y(new_n8564_));
  XOR2   g07562(.A(\A[155] ), .B(new_n8140_), .Y(new_n8565_));
  NAND2  g07563(.A(\A[155] ), .B(\A[154] ), .Y(new_n8566_));
  OAI21  g07564(.A0(new_n8565_), .A1(new_n8137_), .B0(new_n8566_), .Y(new_n8567_));
  XOR2   g07565(.A(new_n8147_), .B(new_n8567_), .Y(new_n8568_));
  NOR2   g07566(.A(\A[152] ), .B(new_n8133_), .Y(new_n8569_));
  OAI21  g07567(.A0(new_n8131_), .A1(\A[151] ), .B0(\A[153] ), .Y(new_n8570_));
  XOR2   g07568(.A(\A[152] ), .B(new_n8133_), .Y(new_n8571_));
  OAI22  g07569(.A0(new_n8571_), .A1(\A[153] ), .B0(new_n8570_), .B1(new_n8569_), .Y(new_n8572_));
  NOR2   g07570(.A(\A[155] ), .B(new_n8140_), .Y(new_n8573_));
  OAI21  g07571(.A0(new_n8138_), .A1(\A[154] ), .B0(\A[156] ), .Y(new_n8574_));
  OAI22  g07572(.A0(new_n8565_), .A1(\A[156] ), .B0(new_n8574_), .B1(new_n8573_), .Y(new_n8575_));
  NAND2  g07573(.A(new_n8575_), .B(new_n8572_), .Y(new_n8576_));
  NAND2  g07574(.A(\A[152] ), .B(\A[151] ), .Y(new_n8577_));
  OAI21  g07575(.A0(new_n8571_), .A1(new_n8130_), .B0(new_n8577_), .Y(new_n8578_));
  NAND2  g07576(.A(new_n8578_), .B(new_n8567_), .Y(new_n8579_));
  OAI21  g07577(.A0(new_n8576_), .A1(new_n8568_), .B0(new_n8579_), .Y(new_n8580_));
  NOR2   g07578(.A(new_n8143_), .B(new_n8136_), .Y(new_n8581_));
  XOR2   g07579(.A(new_n8581_), .B(new_n8568_), .Y(new_n8582_));
  AOI21  g07580(.A0(new_n8580_), .A1(new_n8564_), .B0(new_n8582_), .Y(new_n8583_));
  XOR2   g07581(.A(new_n8124_), .B(new_n8117_), .Y(new_n8584_));
  XOR2   g07582(.A(new_n8128_), .B(new_n8126_), .Y(new_n8585_));
  NAND2  g07583(.A(new_n8112_), .B(\A[157] ), .Y(new_n8586_));
  AOI21  g07584(.A0(\A[158] ), .A1(new_n8110_), .B0(new_n8114_), .Y(new_n8587_));
  AOI22  g07585(.A0(new_n8115_), .A1(new_n8114_), .B0(new_n8587_), .B1(new_n8586_), .Y(new_n8588_));
  NOR2   g07586(.A(new_n8124_), .B(new_n8588_), .Y(new_n8589_));
  NAND2  g07587(.A(\A[161] ), .B(\A[160] ), .Y(new_n8590_));
  NAND2  g07588(.A(new_n8123_), .B(\A[162] ), .Y(new_n8591_));
  NAND2  g07589(.A(\A[158] ), .B(\A[157] ), .Y(new_n8592_));
  NAND2  g07590(.A(new_n8115_), .B(\A[159] ), .Y(new_n8593_));
  AOI22  g07591(.A0(new_n8593_), .A1(new_n8592_), .B0(new_n8591_), .B1(new_n8590_), .Y(new_n8594_));
  AOI21  g07592(.A0(new_n8589_), .A1(new_n8585_), .B0(new_n8594_), .Y(new_n8595_));
  XOR2   g07593(.A(new_n8589_), .B(new_n8585_), .Y(new_n8596_));
  XOR2   g07594(.A(new_n8124_), .B(new_n8588_), .Y(new_n8597_));
  NOR2   g07595(.A(\A[161] ), .B(new_n8121_), .Y(new_n8598_));
  OAI21  g07596(.A0(new_n8119_), .A1(\A[160] ), .B0(\A[162] ), .Y(new_n8599_));
  NAND2  g07597(.A(new_n8123_), .B(new_n8118_), .Y(new_n8600_));
  OAI21  g07598(.A0(new_n8599_), .A1(new_n8598_), .B0(new_n8600_), .Y(new_n8601_));
  NAND2  g07599(.A(new_n8591_), .B(new_n8590_), .Y(new_n8602_));
  NAND2  g07600(.A(new_n8593_), .B(new_n8592_), .Y(new_n8603_));
  NAND4  g07601(.A(new_n8603_), .B(new_n8602_), .C(new_n8601_), .D(new_n8117_), .Y(new_n8604_));
  NAND4  g07602(.A(new_n8578_), .B(new_n8567_), .C(new_n8575_), .D(new_n8572_), .Y(new_n8605_));
  NAND4  g07603(.A(new_n8605_), .B(new_n8564_), .C(new_n8604_), .D(new_n8597_), .Y(new_n8606_));
  OAI211 g07604(.A0(new_n8595_), .A1(new_n8584_), .B0(new_n8606_), .B1(new_n8596_), .Y(new_n8607_));
  XOR2   g07605(.A(new_n8128_), .B(new_n8602_), .Y(new_n8608_));
  XOR2   g07606(.A(new_n8589_), .B(new_n8608_), .Y(new_n8609_));
  NOR4   g07607(.A(new_n8128_), .B(new_n8126_), .C(new_n8124_), .D(new_n8588_), .Y(new_n8610_));
  XOR2   g07608(.A(new_n8143_), .B(new_n8572_), .Y(new_n8611_));
  NOR3   g07609(.A(new_n8611_), .B(new_n8610_), .C(new_n8584_), .Y(new_n8612_));
  AOI221 g07610(.A0(new_n8591_), .A1(new_n8590_), .C0(new_n8127_), .B0(new_n8115_), .B1(\A[159] ), .Y(new_n8613_));
  AOI221 g07611(.A0(new_n8593_), .A1(new_n8592_), .C0(new_n8125_), .B0(new_n8123_), .B1(\A[162] ), .Y(new_n8614_));
  OAI211 g07612(.A0(new_n8614_), .A1(new_n8613_), .B0(new_n8601_), .B1(new_n8117_), .Y(new_n8615_));
  NAND2  g07613(.A(new_n8603_), .B(new_n8602_), .Y(new_n8616_));
  AOI21  g07614(.A0(new_n8616_), .A1(new_n8615_), .B0(new_n8584_), .Y(new_n8617_));
  OAI211 g07615(.A0(new_n8617_), .A1(new_n8609_), .B0(new_n8612_), .B1(new_n8605_), .Y(new_n8618_));
  AOI21  g07616(.A0(new_n8618_), .A1(new_n8607_), .B0(new_n8583_), .Y(new_n8619_));
  OAI21  g07617(.A0(new_n8617_), .A1(new_n8609_), .B0(new_n8606_), .Y(new_n8620_));
  NAND4  g07618(.A(new_n8564_), .B(new_n8596_), .C(new_n8595_), .D(new_n8597_), .Y(new_n8621_));
  OAI21  g07619(.A0(new_n8595_), .A1(new_n8584_), .B0(new_n8605_), .Y(new_n8622_));
  OAI21  g07620(.A0(new_n8622_), .A1(new_n8621_), .B0(new_n8620_), .Y(new_n8623_));
  AOI21  g07621(.A0(new_n8623_), .A1(new_n8583_), .B0(new_n8619_), .Y(new_n8624_));
  XOR2   g07622(.A(new_n8103_), .B(new_n8096_), .Y(new_n8625_));
  XOR2   g07623(.A(\A[167] ), .B(new_n8100_), .Y(new_n8626_));
  NAND2  g07624(.A(\A[167] ), .B(\A[166] ), .Y(new_n8627_));
  OAI21  g07625(.A0(new_n8626_), .A1(new_n8097_), .B0(new_n8627_), .Y(new_n8628_));
  XOR2   g07626(.A(new_n8107_), .B(new_n8628_), .Y(new_n8629_));
  NOR2   g07627(.A(\A[164] ), .B(new_n8093_), .Y(new_n8630_));
  OAI21  g07628(.A0(new_n8091_), .A1(\A[163] ), .B0(\A[165] ), .Y(new_n8631_));
  XOR2   g07629(.A(\A[164] ), .B(new_n8093_), .Y(new_n8632_));
  OAI22  g07630(.A0(new_n8632_), .A1(\A[165] ), .B0(new_n8631_), .B1(new_n8630_), .Y(new_n8633_));
  NOR2   g07631(.A(\A[167] ), .B(new_n8100_), .Y(new_n8634_));
  OAI21  g07632(.A0(new_n8098_), .A1(\A[166] ), .B0(\A[168] ), .Y(new_n8635_));
  OAI22  g07633(.A0(new_n8626_), .A1(\A[168] ), .B0(new_n8635_), .B1(new_n8634_), .Y(new_n8636_));
  NAND2  g07634(.A(new_n8636_), .B(new_n8633_), .Y(new_n8637_));
  NAND2  g07635(.A(\A[164] ), .B(\A[163] ), .Y(new_n8638_));
  OAI21  g07636(.A0(new_n8632_), .A1(new_n8090_), .B0(new_n8638_), .Y(new_n8639_));
  NAND2  g07637(.A(new_n8639_), .B(new_n8628_), .Y(new_n8640_));
  OAI21  g07638(.A0(new_n8637_), .A1(new_n8629_), .B0(new_n8640_), .Y(new_n8641_));
  NOR2   g07639(.A(new_n8103_), .B(new_n8096_), .Y(new_n8642_));
  XOR2   g07640(.A(new_n8642_), .B(new_n8629_), .Y(new_n8643_));
  AOI21  g07641(.A0(new_n8641_), .A1(new_n8625_), .B0(new_n8643_), .Y(new_n8644_));
  NOR2   g07642(.A(\A[170] ), .B(new_n8074_), .Y(new_n8645_));
  OAI21  g07643(.A0(new_n8072_), .A1(\A[169] ), .B0(\A[171] ), .Y(new_n8646_));
  NAND2  g07644(.A(new_n8076_), .B(new_n8071_), .Y(new_n8647_));
  OAI21  g07645(.A0(new_n8646_), .A1(new_n8645_), .B0(new_n8647_), .Y(new_n8648_));
  XOR2   g07646(.A(new_n8084_), .B(new_n8648_), .Y(new_n8649_));
  XOR2   g07647(.A(new_n8088_), .B(new_n8086_), .Y(new_n8650_));
  NOR2   g07648(.A(new_n8084_), .B(new_n8077_), .Y(new_n8651_));
  NAND2  g07649(.A(\A[173] ), .B(\A[172] ), .Y(new_n8652_));
  NAND2  g07650(.A(new_n8083_), .B(\A[174] ), .Y(new_n8653_));
  NAND2  g07651(.A(\A[170] ), .B(\A[169] ), .Y(new_n8654_));
  NAND2  g07652(.A(new_n8076_), .B(\A[171] ), .Y(new_n8655_));
  AOI22  g07653(.A0(new_n8655_), .A1(new_n8654_), .B0(new_n8653_), .B1(new_n8652_), .Y(new_n8656_));
  AOI21  g07654(.A0(new_n8651_), .A1(new_n8650_), .B0(new_n8656_), .Y(new_n8657_));
  XOR2   g07655(.A(new_n8651_), .B(new_n8650_), .Y(new_n8658_));
  XOR2   g07656(.A(new_n8084_), .B(new_n8077_), .Y(new_n8659_));
  NOR2   g07657(.A(\A[173] ), .B(new_n8081_), .Y(new_n8660_));
  OAI21  g07658(.A0(new_n8079_), .A1(\A[172] ), .B0(\A[174] ), .Y(new_n8661_));
  NAND2  g07659(.A(new_n8083_), .B(new_n8078_), .Y(new_n8662_));
  OAI21  g07660(.A0(new_n8661_), .A1(new_n8660_), .B0(new_n8662_), .Y(new_n8663_));
  NAND2  g07661(.A(new_n8653_), .B(new_n8652_), .Y(new_n8664_));
  NAND2  g07662(.A(new_n8655_), .B(new_n8654_), .Y(new_n8665_));
  NAND4  g07663(.A(new_n8665_), .B(new_n8664_), .C(new_n8663_), .D(new_n8648_), .Y(new_n8666_));
  NAND4  g07664(.A(new_n8639_), .B(new_n8628_), .C(new_n8636_), .D(new_n8633_), .Y(new_n8667_));
  NAND4  g07665(.A(new_n8667_), .B(new_n8625_), .C(new_n8666_), .D(new_n8659_), .Y(new_n8668_));
  OAI211 g07666(.A0(new_n8657_), .A1(new_n8649_), .B0(new_n8668_), .B1(new_n8658_), .Y(new_n8669_));
  XOR2   g07667(.A(new_n8088_), .B(new_n8664_), .Y(new_n8670_));
  XOR2   g07668(.A(new_n8651_), .B(new_n8670_), .Y(new_n8671_));
  NOR4   g07669(.A(new_n8088_), .B(new_n8086_), .C(new_n8084_), .D(new_n8077_), .Y(new_n8672_));
  XOR2   g07670(.A(new_n8103_), .B(new_n8633_), .Y(new_n8673_));
  NOR4   g07671(.A(new_n8107_), .B(new_n8105_), .C(new_n8103_), .D(new_n8096_), .Y(new_n8674_));
  NOR4   g07672(.A(new_n8674_), .B(new_n8673_), .C(new_n8672_), .D(new_n8649_), .Y(new_n8675_));
  AOI221 g07673(.A0(new_n8653_), .A1(new_n8652_), .C0(new_n8087_), .B0(new_n8076_), .B1(\A[171] ), .Y(new_n8676_));
  AOI221 g07674(.A0(new_n8655_), .A1(new_n8654_), .C0(new_n8085_), .B0(new_n8083_), .B1(\A[174] ), .Y(new_n8677_));
  OAI211 g07675(.A0(new_n8677_), .A1(new_n8676_), .B0(new_n8663_), .B1(new_n8648_), .Y(new_n8678_));
  NAND2  g07676(.A(new_n8665_), .B(new_n8664_), .Y(new_n8679_));
  AOI21  g07677(.A0(new_n8679_), .A1(new_n8678_), .B0(new_n8649_), .Y(new_n8680_));
  OAI21  g07678(.A0(new_n8680_), .A1(new_n8671_), .B0(new_n8675_), .Y(new_n8681_));
  AOI21  g07679(.A0(new_n8681_), .A1(new_n8669_), .B0(new_n8644_), .Y(new_n8682_));
  OAI21  g07680(.A0(new_n8680_), .A1(new_n8671_), .B0(new_n8668_), .Y(new_n8683_));
  NAND4  g07681(.A(new_n8625_), .B(new_n8658_), .C(new_n8657_), .D(new_n8659_), .Y(new_n8684_));
  OAI21  g07682(.A0(new_n8657_), .A1(new_n8649_), .B0(new_n8667_), .Y(new_n8685_));
  OAI21  g07683(.A0(new_n8685_), .A1(new_n8684_), .B0(new_n8683_), .Y(new_n8686_));
  XOR2   g07684(.A(new_n8124_), .B(new_n8588_), .Y(new_n8687_));
  XOR2   g07685(.A(new_n8148_), .B(new_n8687_), .Y(new_n8688_));
  NAND2  g07686(.A(new_n8688_), .B(new_n8109_), .Y(new_n8689_));
  AOI211 g07687(.A0(new_n8686_), .A1(new_n8644_), .B(new_n8689_), .C(new_n8682_), .Y(new_n8690_));
  XOR2   g07688(.A(new_n8084_), .B(new_n8648_), .Y(new_n8691_));
  XOR2   g07689(.A(new_n8108_), .B(new_n8691_), .Y(new_n8692_));
  NOR2   g07690(.A(new_n8149_), .B(new_n8692_), .Y(new_n8693_));
  AOI21  g07691(.A0(new_n8686_), .A1(new_n8644_), .B0(new_n8682_), .Y(new_n8694_));
  NOR2   g07692(.A(new_n8694_), .B(new_n8693_), .Y(new_n8695_));
  OAI21  g07693(.A0(new_n8695_), .A1(new_n8690_), .B0(new_n8624_), .Y(new_n8696_));
  XOR2   g07694(.A(new_n8147_), .B(new_n8145_), .Y(new_n8697_));
  NOR2   g07695(.A(new_n8147_), .B(new_n8145_), .Y(new_n8698_));
  AOI21  g07696(.A0(new_n8581_), .A1(new_n8697_), .B0(new_n8698_), .Y(new_n8699_));
  XOR2   g07697(.A(new_n8581_), .B(new_n8697_), .Y(new_n8700_));
  OAI21  g07698(.A0(new_n8699_), .A1(new_n8611_), .B0(new_n8700_), .Y(new_n8701_));
  OAI21  g07699(.A0(new_n8595_), .A1(new_n8584_), .B0(new_n8596_), .Y(new_n8702_));
  XOR2   g07700(.A(new_n8702_), .B(new_n8606_), .Y(new_n8703_));
  NAND2  g07701(.A(new_n8703_), .B(new_n8701_), .Y(new_n8704_));
  NAND2  g07702(.A(new_n8623_), .B(new_n8583_), .Y(new_n8705_));
  NAND2  g07703(.A(new_n8705_), .B(new_n8704_), .Y(new_n8706_));
  XOR2   g07704(.A(new_n8107_), .B(new_n8105_), .Y(new_n8707_));
  NOR2   g07705(.A(new_n8107_), .B(new_n8105_), .Y(new_n8708_));
  AOI21  g07706(.A0(new_n8642_), .A1(new_n8707_), .B0(new_n8708_), .Y(new_n8709_));
  XOR2   g07707(.A(new_n8642_), .B(new_n8707_), .Y(new_n8710_));
  OAI21  g07708(.A0(new_n8709_), .A1(new_n8673_), .B0(new_n8710_), .Y(new_n8711_));
  OAI21  g07709(.A0(new_n8657_), .A1(new_n8649_), .B0(new_n8658_), .Y(new_n8712_));
  NAND2  g07710(.A(new_n8679_), .B(new_n8678_), .Y(new_n8713_));
  NOR4   g07711(.A(new_n8673_), .B(new_n8671_), .C(new_n8713_), .D(new_n8649_), .Y(new_n8714_));
  NOR2   g07712(.A(new_n8680_), .B(new_n8674_), .Y(new_n8715_));
  AOI22  g07713(.A0(new_n8715_), .A1(new_n8714_), .B0(new_n8712_), .B1(new_n8668_), .Y(new_n8716_));
  OAI21  g07714(.A0(new_n8716_), .A1(new_n8711_), .B0(new_n8689_), .Y(new_n8717_));
  OAI22  g07715(.A0(new_n8717_), .A1(new_n8682_), .B0(new_n8694_), .B1(new_n8689_), .Y(new_n8718_));
  NAND2  g07716(.A(new_n8718_), .B(new_n8706_), .Y(new_n8719_));
  NOR2   g07717(.A(new_n8231_), .B(new_n8150_), .Y(new_n8720_));
  NAND3  g07718(.A(new_n8720_), .B(new_n8719_), .C(new_n8696_), .Y(new_n8721_));
  XOR2   g07719(.A(new_n8712_), .B(new_n8668_), .Y(new_n8722_));
  NAND2  g07720(.A(new_n8722_), .B(new_n8711_), .Y(new_n8723_));
  NAND2  g07721(.A(new_n8686_), .B(new_n8644_), .Y(new_n8724_));
  NAND3  g07722(.A(new_n8693_), .B(new_n8724_), .C(new_n8723_), .Y(new_n8725_));
  NOR2   g07723(.A(new_n8716_), .B(new_n8711_), .Y(new_n8726_));
  OAI21  g07724(.A0(new_n8726_), .A1(new_n8682_), .B0(new_n8689_), .Y(new_n8727_));
  AOI21  g07725(.A0(new_n8727_), .A1(new_n8725_), .B0(new_n8706_), .Y(new_n8728_));
  NAND3  g07726(.A(new_n8689_), .B(new_n8724_), .C(new_n8723_), .Y(new_n8729_));
  OAI21  g07727(.A0(new_n8726_), .A1(new_n8682_), .B0(new_n8693_), .Y(new_n8730_));
  AOI21  g07728(.A0(new_n8730_), .A1(new_n8729_), .B0(new_n8624_), .Y(new_n8731_));
  INV    g07729(.A(new_n8720_), .Y(new_n8732_));
  OAI21  g07730(.A0(new_n8731_), .A1(new_n8728_), .B0(new_n8732_), .Y(new_n8733_));
  AOI21  g07731(.A0(new_n8733_), .A1(new_n8721_), .B0(new_n8563_), .Y(new_n8734_));
  XOR2   g07732(.A(new_n8555_), .B(new_n8457_), .Y(new_n8735_));
  AOI21  g07733(.A0(new_n8468_), .A1(new_n8426_), .B0(new_n8474_), .Y(new_n8736_));
  OAI21  g07734(.A0(new_n8735_), .A1(new_n8426_), .B0(new_n8736_), .Y(new_n8737_));
  NOR2   g07735(.A(new_n8559_), .B(new_n8554_), .Y(new_n8738_));
  OAI21  g07736(.A0(new_n8738_), .A1(new_n8464_), .B0(new_n8474_), .Y(new_n8739_));
  AOI21  g07737(.A0(new_n8739_), .A1(new_n8737_), .B0(new_n8549_), .Y(new_n8740_));
  AOI21  g07738(.A0(new_n8561_), .A1(new_n8549_), .B0(new_n8740_), .Y(new_n8741_));
  AOI21  g07739(.A0(new_n8718_), .A1(new_n8706_), .B0(new_n8720_), .Y(new_n8742_));
  NAND2  g07740(.A(new_n8742_), .B(new_n8696_), .Y(new_n8743_));
  OAI21  g07741(.A0(new_n8731_), .A1(new_n8728_), .B0(new_n8720_), .Y(new_n8744_));
  AOI21  g07742(.A0(new_n8744_), .A1(new_n8743_), .B0(new_n8741_), .Y(new_n8745_));
  NOR2   g07743(.A(new_n8395_), .B(new_n8232_), .Y(new_n8746_));
  INV    g07744(.A(new_n8746_), .Y(new_n8747_));
  NOR3   g07745(.A(new_n8747_), .B(new_n8745_), .C(new_n8734_), .Y(new_n8748_));
  NOR3   g07746(.A(new_n8732_), .B(new_n8731_), .C(new_n8728_), .Y(new_n8749_));
  AOI21  g07747(.A0(new_n8719_), .A1(new_n8696_), .B0(new_n8720_), .Y(new_n8750_));
  OAI21  g07748(.A0(new_n8750_), .A1(new_n8749_), .B0(new_n8741_), .Y(new_n8751_));
  NOR3   g07749(.A(new_n8720_), .B(new_n8731_), .C(new_n8728_), .Y(new_n8752_));
  AOI21  g07750(.A0(new_n8719_), .A1(new_n8696_), .B0(new_n8732_), .Y(new_n8753_));
  OAI21  g07751(.A0(new_n8753_), .A1(new_n8752_), .B0(new_n8563_), .Y(new_n8754_));
  AOI21  g07752(.A0(new_n8754_), .A1(new_n8751_), .B0(new_n8746_), .Y(new_n8755_));
  XOR2   g07753(.A(new_n8306_), .B(new_n8299_), .Y(new_n8756_));
  XOR2   g07754(.A(\A[107] ), .B(new_n8303_), .Y(new_n8757_));
  NAND2  g07755(.A(\A[107] ), .B(\A[106] ), .Y(new_n8758_));
  OAI21  g07756(.A0(new_n8757_), .A1(new_n8300_), .B0(new_n8758_), .Y(new_n8759_));
  XOR2   g07757(.A(new_n8310_), .B(new_n8759_), .Y(new_n8760_));
  NOR2   g07758(.A(\A[104] ), .B(new_n8296_), .Y(new_n8761_));
  OAI21  g07759(.A0(new_n8294_), .A1(\A[103] ), .B0(\A[105] ), .Y(new_n8762_));
  XOR2   g07760(.A(\A[104] ), .B(new_n8296_), .Y(new_n8763_));
  OAI22  g07761(.A0(new_n8763_), .A1(\A[105] ), .B0(new_n8762_), .B1(new_n8761_), .Y(new_n8764_));
  NOR2   g07762(.A(\A[107] ), .B(new_n8303_), .Y(new_n8765_));
  OAI21  g07763(.A0(new_n8301_), .A1(\A[106] ), .B0(\A[108] ), .Y(new_n8766_));
  OAI22  g07764(.A0(new_n8757_), .A1(\A[108] ), .B0(new_n8766_), .B1(new_n8765_), .Y(new_n8767_));
  NAND2  g07765(.A(new_n8767_), .B(new_n8764_), .Y(new_n8768_));
  NAND2  g07766(.A(\A[104] ), .B(\A[103] ), .Y(new_n8769_));
  OAI21  g07767(.A0(new_n8763_), .A1(new_n8293_), .B0(new_n8769_), .Y(new_n8770_));
  NAND2  g07768(.A(new_n8770_), .B(new_n8759_), .Y(new_n8771_));
  OAI21  g07769(.A0(new_n8768_), .A1(new_n8760_), .B0(new_n8771_), .Y(new_n8772_));
  NOR2   g07770(.A(new_n8306_), .B(new_n8299_), .Y(new_n8773_));
  XOR2   g07771(.A(new_n8773_), .B(new_n8760_), .Y(new_n8774_));
  AOI21  g07772(.A0(new_n8772_), .A1(new_n8756_), .B0(new_n8774_), .Y(new_n8775_));
  XOR2   g07773(.A(new_n8287_), .B(new_n8280_), .Y(new_n8776_));
  XOR2   g07774(.A(new_n8291_), .B(new_n8289_), .Y(new_n8777_));
  NAND2  g07775(.A(new_n8275_), .B(\A[109] ), .Y(new_n8778_));
  AOI21  g07776(.A0(\A[110] ), .A1(new_n8273_), .B0(new_n8277_), .Y(new_n8779_));
  AOI22  g07777(.A0(new_n8278_), .A1(new_n8277_), .B0(new_n8779_), .B1(new_n8778_), .Y(new_n8780_));
  NOR2   g07778(.A(new_n8287_), .B(new_n8780_), .Y(new_n8781_));
  NAND2  g07779(.A(\A[113] ), .B(\A[112] ), .Y(new_n8782_));
  NAND2  g07780(.A(new_n8286_), .B(\A[114] ), .Y(new_n8783_));
  NAND2  g07781(.A(\A[110] ), .B(\A[109] ), .Y(new_n8784_));
  NAND2  g07782(.A(new_n8278_), .B(\A[111] ), .Y(new_n8785_));
  AOI22  g07783(.A0(new_n8785_), .A1(new_n8784_), .B0(new_n8783_), .B1(new_n8782_), .Y(new_n8786_));
  AOI21  g07784(.A0(new_n8781_), .A1(new_n8777_), .B0(new_n8786_), .Y(new_n8787_));
  XOR2   g07785(.A(new_n8781_), .B(new_n8777_), .Y(new_n8788_));
  XOR2   g07786(.A(new_n8287_), .B(new_n8780_), .Y(new_n8789_));
  NOR2   g07787(.A(\A[113] ), .B(new_n8284_), .Y(new_n8790_));
  OAI21  g07788(.A0(new_n8282_), .A1(\A[112] ), .B0(\A[114] ), .Y(new_n8791_));
  NAND2  g07789(.A(new_n8286_), .B(new_n8281_), .Y(new_n8792_));
  OAI21  g07790(.A0(new_n8791_), .A1(new_n8790_), .B0(new_n8792_), .Y(new_n8793_));
  NAND2  g07791(.A(new_n8783_), .B(new_n8782_), .Y(new_n8794_));
  NAND2  g07792(.A(new_n8785_), .B(new_n8784_), .Y(new_n8795_));
  NAND4  g07793(.A(new_n8795_), .B(new_n8794_), .C(new_n8793_), .D(new_n8280_), .Y(new_n8796_));
  NAND4  g07794(.A(new_n8770_), .B(new_n8759_), .C(new_n8767_), .D(new_n8764_), .Y(new_n8797_));
  NAND4  g07795(.A(new_n8797_), .B(new_n8756_), .C(new_n8796_), .D(new_n8789_), .Y(new_n8798_));
  OAI211 g07796(.A0(new_n8787_), .A1(new_n8776_), .B0(new_n8798_), .B1(new_n8788_), .Y(new_n8799_));
  XOR2   g07797(.A(new_n8291_), .B(new_n8794_), .Y(new_n8800_));
  XOR2   g07798(.A(new_n8781_), .B(new_n8800_), .Y(new_n8801_));
  NOR4   g07799(.A(new_n8291_), .B(new_n8289_), .C(new_n8287_), .D(new_n8780_), .Y(new_n8802_));
  XOR2   g07800(.A(new_n8306_), .B(new_n8764_), .Y(new_n8803_));
  NOR4   g07801(.A(new_n8310_), .B(new_n8308_), .C(new_n8306_), .D(new_n8299_), .Y(new_n8804_));
  NOR4   g07802(.A(new_n8804_), .B(new_n8803_), .C(new_n8802_), .D(new_n8776_), .Y(new_n8805_));
  AOI221 g07803(.A0(new_n8783_), .A1(new_n8782_), .C0(new_n8290_), .B0(new_n8278_), .B1(\A[111] ), .Y(new_n8806_));
  AOI221 g07804(.A0(new_n8785_), .A1(new_n8784_), .C0(new_n8288_), .B0(new_n8286_), .B1(\A[114] ), .Y(new_n8807_));
  OAI211 g07805(.A0(new_n8807_), .A1(new_n8806_), .B0(new_n8793_), .B1(new_n8280_), .Y(new_n8808_));
  NAND2  g07806(.A(new_n8795_), .B(new_n8794_), .Y(new_n8809_));
  AOI21  g07807(.A0(new_n8809_), .A1(new_n8808_), .B0(new_n8776_), .Y(new_n8810_));
  OAI21  g07808(.A0(new_n8810_), .A1(new_n8801_), .B0(new_n8805_), .Y(new_n8811_));
  AOI21  g07809(.A0(new_n8811_), .A1(new_n8799_), .B0(new_n8775_), .Y(new_n8812_));
  NOR2   g07810(.A(new_n8810_), .B(new_n8801_), .Y(new_n8813_));
  NAND4  g07811(.A(new_n8756_), .B(new_n8788_), .C(new_n8787_), .D(new_n8789_), .Y(new_n8814_));
  OAI21  g07812(.A0(new_n8787_), .A1(new_n8776_), .B0(new_n8797_), .Y(new_n8815_));
  OAI22  g07813(.A0(new_n8815_), .A1(new_n8814_), .B0(new_n8813_), .B1(new_n8805_), .Y(new_n8816_));
  AOI21  g07814(.A0(new_n8816_), .A1(new_n8775_), .B0(new_n8812_), .Y(new_n8817_));
  XOR2   g07815(.A(new_n8266_), .B(new_n8259_), .Y(new_n8818_));
  XOR2   g07816(.A(\A[119] ), .B(new_n8263_), .Y(new_n8819_));
  NAND2  g07817(.A(\A[119] ), .B(\A[118] ), .Y(new_n8820_));
  OAI21  g07818(.A0(new_n8819_), .A1(new_n8260_), .B0(new_n8820_), .Y(new_n8821_));
  XOR2   g07819(.A(new_n8270_), .B(new_n8821_), .Y(new_n8822_));
  NOR2   g07820(.A(\A[116] ), .B(new_n8256_), .Y(new_n8823_));
  OAI21  g07821(.A0(new_n8254_), .A1(\A[115] ), .B0(\A[117] ), .Y(new_n8824_));
  XOR2   g07822(.A(\A[116] ), .B(new_n8256_), .Y(new_n8825_));
  OAI22  g07823(.A0(new_n8825_), .A1(\A[117] ), .B0(new_n8824_), .B1(new_n8823_), .Y(new_n8826_));
  NOR2   g07824(.A(\A[119] ), .B(new_n8263_), .Y(new_n8827_));
  OAI21  g07825(.A0(new_n8261_), .A1(\A[118] ), .B0(\A[120] ), .Y(new_n8828_));
  OAI22  g07826(.A0(new_n8819_), .A1(\A[120] ), .B0(new_n8828_), .B1(new_n8827_), .Y(new_n8829_));
  NAND2  g07827(.A(new_n8829_), .B(new_n8826_), .Y(new_n8830_));
  NAND2  g07828(.A(\A[116] ), .B(\A[115] ), .Y(new_n8831_));
  OAI21  g07829(.A0(new_n8825_), .A1(new_n8253_), .B0(new_n8831_), .Y(new_n8832_));
  NAND2  g07830(.A(new_n8832_), .B(new_n8821_), .Y(new_n8833_));
  OAI21  g07831(.A0(new_n8830_), .A1(new_n8822_), .B0(new_n8833_), .Y(new_n8834_));
  NOR2   g07832(.A(new_n8266_), .B(new_n8259_), .Y(new_n8835_));
  XOR2   g07833(.A(new_n8835_), .B(new_n8822_), .Y(new_n8836_));
  AOI21  g07834(.A0(new_n8834_), .A1(new_n8818_), .B0(new_n8836_), .Y(new_n8837_));
  NOR2   g07835(.A(\A[122] ), .B(new_n8237_), .Y(new_n8838_));
  OAI21  g07836(.A0(new_n8235_), .A1(\A[121] ), .B0(\A[123] ), .Y(new_n8839_));
  NAND2  g07837(.A(new_n8239_), .B(new_n8234_), .Y(new_n8840_));
  OAI21  g07838(.A0(new_n8839_), .A1(new_n8838_), .B0(new_n8840_), .Y(new_n8841_));
  XOR2   g07839(.A(new_n8247_), .B(new_n8841_), .Y(new_n8842_));
  XOR2   g07840(.A(new_n8251_), .B(new_n8249_), .Y(new_n8843_));
  NOR2   g07841(.A(new_n8247_), .B(new_n8240_), .Y(new_n8844_));
  NAND2  g07842(.A(\A[125] ), .B(\A[124] ), .Y(new_n8845_));
  NAND2  g07843(.A(new_n8246_), .B(\A[126] ), .Y(new_n8846_));
  NAND2  g07844(.A(\A[122] ), .B(\A[121] ), .Y(new_n8847_));
  NAND2  g07845(.A(new_n8239_), .B(\A[123] ), .Y(new_n8848_));
  AOI22  g07846(.A0(new_n8848_), .A1(new_n8847_), .B0(new_n8846_), .B1(new_n8845_), .Y(new_n8849_));
  AOI21  g07847(.A0(new_n8844_), .A1(new_n8843_), .B0(new_n8849_), .Y(new_n8850_));
  XOR2   g07848(.A(new_n8844_), .B(new_n8843_), .Y(new_n8851_));
  XOR2   g07849(.A(new_n8247_), .B(new_n8240_), .Y(new_n8852_));
  NOR2   g07850(.A(\A[125] ), .B(new_n8244_), .Y(new_n8853_));
  OAI21  g07851(.A0(new_n8242_), .A1(\A[124] ), .B0(\A[126] ), .Y(new_n8854_));
  NAND2  g07852(.A(new_n8246_), .B(new_n8241_), .Y(new_n8855_));
  OAI21  g07853(.A0(new_n8854_), .A1(new_n8853_), .B0(new_n8855_), .Y(new_n8856_));
  NAND2  g07854(.A(new_n8846_), .B(new_n8845_), .Y(new_n8857_));
  NAND2  g07855(.A(new_n8848_), .B(new_n8847_), .Y(new_n8858_));
  NAND4  g07856(.A(new_n8858_), .B(new_n8857_), .C(new_n8856_), .D(new_n8841_), .Y(new_n8859_));
  NAND4  g07857(.A(new_n8832_), .B(new_n8821_), .C(new_n8829_), .D(new_n8826_), .Y(new_n8860_));
  NAND4  g07858(.A(new_n8860_), .B(new_n8818_), .C(new_n8859_), .D(new_n8852_), .Y(new_n8861_));
  OAI211 g07859(.A0(new_n8850_), .A1(new_n8842_), .B0(new_n8861_), .B1(new_n8851_), .Y(new_n8862_));
  XOR2   g07860(.A(new_n8251_), .B(new_n8857_), .Y(new_n8863_));
  XOR2   g07861(.A(new_n8844_), .B(new_n8863_), .Y(new_n8864_));
  NOR4   g07862(.A(new_n8251_), .B(new_n8249_), .C(new_n8247_), .D(new_n8240_), .Y(new_n8865_));
  XOR2   g07863(.A(new_n8266_), .B(new_n8826_), .Y(new_n8866_));
  NOR4   g07864(.A(new_n8270_), .B(new_n8268_), .C(new_n8266_), .D(new_n8259_), .Y(new_n8867_));
  NOR4   g07865(.A(new_n8867_), .B(new_n8866_), .C(new_n8865_), .D(new_n8842_), .Y(new_n8868_));
  AOI221 g07866(.A0(new_n8846_), .A1(new_n8845_), .C0(new_n8250_), .B0(new_n8239_), .B1(\A[123] ), .Y(new_n8869_));
  AOI221 g07867(.A0(new_n8848_), .A1(new_n8847_), .C0(new_n8248_), .B0(new_n8246_), .B1(\A[126] ), .Y(new_n8870_));
  OAI211 g07868(.A0(new_n8870_), .A1(new_n8869_), .B0(new_n8856_), .B1(new_n8841_), .Y(new_n8871_));
  NAND2  g07869(.A(new_n8858_), .B(new_n8857_), .Y(new_n8872_));
  AOI21  g07870(.A0(new_n8872_), .A1(new_n8871_), .B0(new_n8842_), .Y(new_n8873_));
  OAI21  g07871(.A0(new_n8873_), .A1(new_n8864_), .B0(new_n8868_), .Y(new_n8874_));
  AOI21  g07872(.A0(new_n8874_), .A1(new_n8862_), .B0(new_n8837_), .Y(new_n8875_));
  OAI21  g07873(.A0(new_n8873_), .A1(new_n8864_), .B0(new_n8861_), .Y(new_n8876_));
  NAND4  g07874(.A(new_n8818_), .B(new_n8851_), .C(new_n8850_), .D(new_n8852_), .Y(new_n8877_));
  OAI21  g07875(.A0(new_n8850_), .A1(new_n8842_), .B0(new_n8860_), .Y(new_n8878_));
  OAI21  g07876(.A0(new_n8878_), .A1(new_n8877_), .B0(new_n8876_), .Y(new_n8879_));
  XOR2   g07877(.A(new_n8287_), .B(new_n8780_), .Y(new_n8880_));
  XOR2   g07878(.A(new_n8311_), .B(new_n8880_), .Y(new_n8881_));
  NAND2  g07879(.A(new_n8881_), .B(new_n8272_), .Y(new_n8882_));
  AOI211 g07880(.A0(new_n8879_), .A1(new_n8837_), .B(new_n8882_), .C(new_n8875_), .Y(new_n8883_));
  XOR2   g07881(.A(new_n8247_), .B(new_n8841_), .Y(new_n8884_));
  XOR2   g07882(.A(new_n8271_), .B(new_n8884_), .Y(new_n8885_));
  NOR2   g07883(.A(new_n8312_), .B(new_n8885_), .Y(new_n8886_));
  AOI21  g07884(.A0(new_n8879_), .A1(new_n8837_), .B0(new_n8875_), .Y(new_n8887_));
  NOR2   g07885(.A(new_n8887_), .B(new_n8886_), .Y(new_n8888_));
  OAI21  g07886(.A0(new_n8888_), .A1(new_n8883_), .B0(new_n8817_), .Y(new_n8889_));
  XOR2   g07887(.A(new_n8813_), .B(new_n8798_), .Y(new_n8890_));
  NAND2  g07888(.A(new_n8816_), .B(new_n8775_), .Y(new_n8891_));
  OAI21  g07889(.A0(new_n8890_), .A1(new_n8775_), .B0(new_n8891_), .Y(new_n8892_));
  XOR2   g07890(.A(new_n8270_), .B(new_n8268_), .Y(new_n8893_));
  NOR2   g07891(.A(new_n8270_), .B(new_n8268_), .Y(new_n8894_));
  AOI21  g07892(.A0(new_n8835_), .A1(new_n8893_), .B0(new_n8894_), .Y(new_n8895_));
  XOR2   g07893(.A(new_n8835_), .B(new_n8893_), .Y(new_n8896_));
  OAI21  g07894(.A0(new_n8895_), .A1(new_n8866_), .B0(new_n8896_), .Y(new_n8897_));
  OAI21  g07895(.A0(new_n8850_), .A1(new_n8842_), .B0(new_n8851_), .Y(new_n8898_));
  NAND2  g07896(.A(new_n8872_), .B(new_n8871_), .Y(new_n8899_));
  NOR4   g07897(.A(new_n8866_), .B(new_n8864_), .C(new_n8899_), .D(new_n8842_), .Y(new_n8900_));
  NOR2   g07898(.A(new_n8873_), .B(new_n8867_), .Y(new_n8901_));
  AOI22  g07899(.A0(new_n8901_), .A1(new_n8900_), .B0(new_n8898_), .B1(new_n8861_), .Y(new_n8902_));
  OAI21  g07900(.A0(new_n8902_), .A1(new_n8897_), .B0(new_n8882_), .Y(new_n8903_));
  OAI22  g07901(.A0(new_n8903_), .A1(new_n8875_), .B0(new_n8887_), .B1(new_n8882_), .Y(new_n8904_));
  NAND2  g07902(.A(new_n8904_), .B(new_n8892_), .Y(new_n8905_));
  NOR2   g07903(.A(new_n8394_), .B(new_n8313_), .Y(new_n8906_));
  NAND3  g07904(.A(new_n8906_), .B(new_n8905_), .C(new_n8889_), .Y(new_n8907_));
  XOR2   g07905(.A(new_n8898_), .B(new_n8861_), .Y(new_n8908_));
  NAND2  g07906(.A(new_n8908_), .B(new_n8897_), .Y(new_n8909_));
  NAND2  g07907(.A(new_n8879_), .B(new_n8837_), .Y(new_n8910_));
  NAND3  g07908(.A(new_n8886_), .B(new_n8910_), .C(new_n8909_), .Y(new_n8911_));
  NOR2   g07909(.A(new_n8902_), .B(new_n8897_), .Y(new_n8912_));
  OAI21  g07910(.A0(new_n8912_), .A1(new_n8875_), .B0(new_n8882_), .Y(new_n8913_));
  AOI21  g07911(.A0(new_n8913_), .A1(new_n8911_), .B0(new_n8892_), .Y(new_n8914_));
  NAND3  g07912(.A(new_n8882_), .B(new_n8910_), .C(new_n8909_), .Y(new_n8915_));
  OAI21  g07913(.A0(new_n8912_), .A1(new_n8875_), .B0(new_n8886_), .Y(new_n8916_));
  AOI21  g07914(.A0(new_n8916_), .A1(new_n8915_), .B0(new_n8817_), .Y(new_n8917_));
  INV    g07915(.A(new_n8906_), .Y(new_n8918_));
  OAI21  g07916(.A0(new_n8917_), .A1(new_n8914_), .B0(new_n8918_), .Y(new_n8919_));
  XOR2   g07917(.A(new_n8347_), .B(new_n8340_), .Y(new_n8920_));
  XOR2   g07918(.A(\A[95] ), .B(new_n8344_), .Y(new_n8921_));
  NAND2  g07919(.A(\A[95] ), .B(\A[94] ), .Y(new_n8922_));
  OAI21  g07920(.A0(new_n8921_), .A1(new_n8341_), .B0(new_n8922_), .Y(new_n8923_));
  XOR2   g07921(.A(new_n8351_), .B(new_n8923_), .Y(new_n8924_));
  NOR2   g07922(.A(\A[92] ), .B(new_n8337_), .Y(new_n8925_));
  OAI21  g07923(.A0(new_n8335_), .A1(\A[91] ), .B0(\A[93] ), .Y(new_n8926_));
  XOR2   g07924(.A(\A[92] ), .B(new_n8337_), .Y(new_n8927_));
  OAI22  g07925(.A0(new_n8927_), .A1(\A[93] ), .B0(new_n8926_), .B1(new_n8925_), .Y(new_n8928_));
  NOR2   g07926(.A(\A[95] ), .B(new_n8344_), .Y(new_n8929_));
  OAI21  g07927(.A0(new_n8342_), .A1(\A[94] ), .B0(\A[96] ), .Y(new_n8930_));
  OAI22  g07928(.A0(new_n8921_), .A1(\A[96] ), .B0(new_n8930_), .B1(new_n8929_), .Y(new_n8931_));
  NAND2  g07929(.A(new_n8931_), .B(new_n8928_), .Y(new_n8932_));
  NAND2  g07930(.A(\A[92] ), .B(\A[91] ), .Y(new_n8933_));
  OAI21  g07931(.A0(new_n8927_), .A1(new_n8334_), .B0(new_n8933_), .Y(new_n8934_));
  NAND2  g07932(.A(new_n8934_), .B(new_n8923_), .Y(new_n8935_));
  OAI21  g07933(.A0(new_n8932_), .A1(new_n8924_), .B0(new_n8935_), .Y(new_n8936_));
  NOR2   g07934(.A(new_n8347_), .B(new_n8340_), .Y(new_n8937_));
  XOR2   g07935(.A(new_n8937_), .B(new_n8924_), .Y(new_n8938_));
  AOI21  g07936(.A0(new_n8936_), .A1(new_n8920_), .B0(new_n8938_), .Y(new_n8939_));
  NOR2   g07937(.A(\A[98] ), .B(new_n8318_), .Y(new_n8940_));
  OAI21  g07938(.A0(new_n8316_), .A1(\A[97] ), .B0(\A[99] ), .Y(new_n8941_));
  NAND2  g07939(.A(new_n8320_), .B(new_n8315_), .Y(new_n8942_));
  OAI21  g07940(.A0(new_n8941_), .A1(new_n8940_), .B0(new_n8942_), .Y(new_n8943_));
  XOR2   g07941(.A(new_n8328_), .B(new_n8943_), .Y(new_n8944_));
  XOR2   g07942(.A(new_n8332_), .B(new_n8330_), .Y(new_n8945_));
  NOR2   g07943(.A(new_n8328_), .B(new_n8321_), .Y(new_n8946_));
  NAND2  g07944(.A(\A[101] ), .B(\A[100] ), .Y(new_n8947_));
  NAND2  g07945(.A(new_n8327_), .B(\A[102] ), .Y(new_n8948_));
  NAND2  g07946(.A(\A[98] ), .B(\A[97] ), .Y(new_n8949_));
  NAND2  g07947(.A(new_n8320_), .B(\A[99] ), .Y(new_n8950_));
  AOI22  g07948(.A0(new_n8950_), .A1(new_n8949_), .B0(new_n8948_), .B1(new_n8947_), .Y(new_n8951_));
  AOI21  g07949(.A0(new_n8946_), .A1(new_n8945_), .B0(new_n8951_), .Y(new_n8952_));
  XOR2   g07950(.A(new_n8946_), .B(new_n8945_), .Y(new_n8953_));
  XOR2   g07951(.A(new_n8328_), .B(new_n8321_), .Y(new_n8954_));
  NOR2   g07952(.A(\A[101] ), .B(new_n8325_), .Y(new_n8955_));
  OAI21  g07953(.A0(new_n8323_), .A1(\A[100] ), .B0(\A[102] ), .Y(new_n8956_));
  NAND2  g07954(.A(new_n8327_), .B(new_n8322_), .Y(new_n8957_));
  OAI21  g07955(.A0(new_n8956_), .A1(new_n8955_), .B0(new_n8957_), .Y(new_n8958_));
  NAND2  g07956(.A(new_n8948_), .B(new_n8947_), .Y(new_n8959_));
  NAND2  g07957(.A(new_n8950_), .B(new_n8949_), .Y(new_n8960_));
  NAND4  g07958(.A(new_n8960_), .B(new_n8959_), .C(new_n8958_), .D(new_n8943_), .Y(new_n8961_));
  NAND4  g07959(.A(new_n8934_), .B(new_n8923_), .C(new_n8931_), .D(new_n8928_), .Y(new_n8962_));
  NAND4  g07960(.A(new_n8962_), .B(new_n8920_), .C(new_n8961_), .D(new_n8954_), .Y(new_n8963_));
  OAI211 g07961(.A0(new_n8952_), .A1(new_n8944_), .B0(new_n8963_), .B1(new_n8953_), .Y(new_n8964_));
  XOR2   g07962(.A(new_n8332_), .B(new_n8959_), .Y(new_n8965_));
  XOR2   g07963(.A(new_n8946_), .B(new_n8965_), .Y(new_n8966_));
  NOR4   g07964(.A(new_n8332_), .B(new_n8330_), .C(new_n8328_), .D(new_n8321_), .Y(new_n8967_));
  XOR2   g07965(.A(new_n8347_), .B(new_n8928_), .Y(new_n8968_));
  NOR4   g07966(.A(new_n8351_), .B(new_n8349_), .C(new_n8347_), .D(new_n8340_), .Y(new_n8969_));
  NOR4   g07967(.A(new_n8969_), .B(new_n8968_), .C(new_n8967_), .D(new_n8944_), .Y(new_n8970_));
  AOI221 g07968(.A0(new_n8948_), .A1(new_n8947_), .C0(new_n8331_), .B0(new_n8320_), .B1(\A[99] ), .Y(new_n8971_));
  AOI221 g07969(.A0(new_n8950_), .A1(new_n8949_), .C0(new_n8329_), .B0(new_n8327_), .B1(\A[102] ), .Y(new_n8972_));
  OAI211 g07970(.A0(new_n8972_), .A1(new_n8971_), .B0(new_n8958_), .B1(new_n8943_), .Y(new_n8973_));
  NAND2  g07971(.A(new_n8960_), .B(new_n8959_), .Y(new_n8974_));
  AOI21  g07972(.A0(new_n8974_), .A1(new_n8973_), .B0(new_n8944_), .Y(new_n8975_));
  OAI21  g07973(.A0(new_n8975_), .A1(new_n8966_), .B0(new_n8970_), .Y(new_n8976_));
  AOI21  g07974(.A0(new_n8976_), .A1(new_n8964_), .B0(new_n8939_), .Y(new_n8977_));
  OAI21  g07975(.A0(new_n8975_), .A1(new_n8966_), .B0(new_n8963_), .Y(new_n8978_));
  NAND4  g07976(.A(new_n8920_), .B(new_n8953_), .C(new_n8952_), .D(new_n8954_), .Y(new_n8979_));
  OAI21  g07977(.A0(new_n8952_), .A1(new_n8944_), .B0(new_n8962_), .Y(new_n8980_));
  OAI21  g07978(.A0(new_n8980_), .A1(new_n8979_), .B0(new_n8978_), .Y(new_n8981_));
  NAND2  g07979(.A(new_n8356_), .B(\A[85] ), .Y(new_n8982_));
  AOI21  g07980(.A0(\A[86] ), .A1(new_n8354_), .B0(new_n8358_), .Y(new_n8983_));
  AOI22  g07981(.A0(new_n8359_), .A1(new_n8358_), .B0(new_n8983_), .B1(new_n8982_), .Y(new_n8984_));
  XOR2   g07982(.A(new_n8368_), .B(new_n8984_), .Y(new_n8985_));
  XOR2   g07983(.A(new_n8392_), .B(new_n8985_), .Y(new_n8986_));
  NAND2  g07984(.A(new_n8986_), .B(new_n8353_), .Y(new_n8987_));
  AOI211 g07985(.A0(new_n8981_), .A1(new_n8939_), .B(new_n8987_), .C(new_n8977_), .Y(new_n8988_));
  XOR2   g07986(.A(new_n8328_), .B(new_n8943_), .Y(new_n8989_));
  XOR2   g07987(.A(new_n8352_), .B(new_n8989_), .Y(new_n8990_));
  NOR2   g07988(.A(new_n8393_), .B(new_n8990_), .Y(new_n8991_));
  AOI21  g07989(.A0(new_n8981_), .A1(new_n8939_), .B0(new_n8977_), .Y(new_n8992_));
  NOR2   g07990(.A(new_n8992_), .B(new_n8991_), .Y(new_n8993_));
  XOR2   g07991(.A(new_n8387_), .B(new_n8380_), .Y(new_n8994_));
  XOR2   g07992(.A(\A[83] ), .B(new_n8384_), .Y(new_n8995_));
  NAND2  g07993(.A(\A[83] ), .B(\A[82] ), .Y(new_n8996_));
  OAI21  g07994(.A0(new_n8995_), .A1(new_n8381_), .B0(new_n8996_), .Y(new_n8997_));
  XOR2   g07995(.A(new_n8391_), .B(new_n8997_), .Y(new_n8998_));
  NOR2   g07996(.A(\A[80] ), .B(new_n8377_), .Y(new_n8999_));
  OAI21  g07997(.A0(new_n8375_), .A1(\A[79] ), .B0(\A[81] ), .Y(new_n9000_));
  XOR2   g07998(.A(\A[80] ), .B(new_n8377_), .Y(new_n9001_));
  OAI22  g07999(.A0(new_n9001_), .A1(\A[81] ), .B0(new_n9000_), .B1(new_n8999_), .Y(new_n9002_));
  NOR2   g08000(.A(\A[83] ), .B(new_n8384_), .Y(new_n9003_));
  OAI21  g08001(.A0(new_n8382_), .A1(\A[82] ), .B0(\A[84] ), .Y(new_n9004_));
  OAI22  g08002(.A0(new_n8995_), .A1(\A[84] ), .B0(new_n9004_), .B1(new_n9003_), .Y(new_n9005_));
  NAND2  g08003(.A(new_n9005_), .B(new_n9002_), .Y(new_n9006_));
  NAND2  g08004(.A(\A[80] ), .B(\A[79] ), .Y(new_n9007_));
  OAI21  g08005(.A0(new_n9001_), .A1(new_n8374_), .B0(new_n9007_), .Y(new_n9008_));
  NAND2  g08006(.A(new_n9008_), .B(new_n8997_), .Y(new_n9009_));
  OAI21  g08007(.A0(new_n9006_), .A1(new_n8998_), .B0(new_n9009_), .Y(new_n9010_));
  NOR2   g08008(.A(new_n8387_), .B(new_n8380_), .Y(new_n9011_));
  XOR2   g08009(.A(new_n9011_), .B(new_n8998_), .Y(new_n9012_));
  AOI21  g08010(.A0(new_n9010_), .A1(new_n8994_), .B0(new_n9012_), .Y(new_n9013_));
  XOR2   g08011(.A(new_n8368_), .B(new_n8361_), .Y(new_n9014_));
  XOR2   g08012(.A(new_n8372_), .B(new_n8370_), .Y(new_n9015_));
  NOR2   g08013(.A(new_n8368_), .B(new_n8984_), .Y(new_n9016_));
  NAND2  g08014(.A(\A[89] ), .B(\A[88] ), .Y(new_n9017_));
  NAND2  g08015(.A(new_n8367_), .B(\A[90] ), .Y(new_n9018_));
  NAND2  g08016(.A(\A[86] ), .B(\A[85] ), .Y(new_n9019_));
  NAND2  g08017(.A(new_n8359_), .B(\A[87] ), .Y(new_n9020_));
  AOI22  g08018(.A0(new_n9020_), .A1(new_n9019_), .B0(new_n9018_), .B1(new_n9017_), .Y(new_n9021_));
  AOI21  g08019(.A0(new_n9016_), .A1(new_n9015_), .B0(new_n9021_), .Y(new_n9022_));
  XOR2   g08020(.A(new_n9016_), .B(new_n9015_), .Y(new_n9023_));
  XOR2   g08021(.A(new_n8368_), .B(new_n8984_), .Y(new_n9024_));
  NOR2   g08022(.A(\A[89] ), .B(new_n8365_), .Y(new_n9025_));
  OAI21  g08023(.A0(new_n8363_), .A1(\A[88] ), .B0(\A[90] ), .Y(new_n9026_));
  NAND2  g08024(.A(new_n8367_), .B(new_n8362_), .Y(new_n9027_));
  OAI21  g08025(.A0(new_n9026_), .A1(new_n9025_), .B0(new_n9027_), .Y(new_n9028_));
  NAND2  g08026(.A(new_n9018_), .B(new_n9017_), .Y(new_n9029_));
  NAND2  g08027(.A(new_n9020_), .B(new_n9019_), .Y(new_n9030_));
  NAND4  g08028(.A(new_n9030_), .B(new_n9029_), .C(new_n9028_), .D(new_n8361_), .Y(new_n9031_));
  NAND4  g08029(.A(new_n9008_), .B(new_n8997_), .C(new_n9005_), .D(new_n9002_), .Y(new_n9032_));
  NAND4  g08030(.A(new_n9032_), .B(new_n8994_), .C(new_n9031_), .D(new_n9024_), .Y(new_n9033_));
  OAI211 g08031(.A0(new_n9022_), .A1(new_n9014_), .B0(new_n9033_), .B1(new_n9023_), .Y(new_n9034_));
  XOR2   g08032(.A(new_n8372_), .B(new_n9029_), .Y(new_n9035_));
  XOR2   g08033(.A(new_n9016_), .B(new_n9035_), .Y(new_n9036_));
  NOR4   g08034(.A(new_n8372_), .B(new_n8370_), .C(new_n8368_), .D(new_n8984_), .Y(new_n9037_));
  XOR2   g08035(.A(new_n8387_), .B(new_n9002_), .Y(new_n9038_));
  NOR4   g08036(.A(new_n8391_), .B(new_n8389_), .C(new_n8387_), .D(new_n8380_), .Y(new_n9039_));
  NOR4   g08037(.A(new_n9039_), .B(new_n9038_), .C(new_n9037_), .D(new_n9014_), .Y(new_n9040_));
  AOI221 g08038(.A0(new_n9018_), .A1(new_n9017_), .C0(new_n8371_), .B0(new_n8359_), .B1(\A[87] ), .Y(new_n9041_));
  AOI221 g08039(.A0(new_n9020_), .A1(new_n9019_), .C0(new_n8369_), .B0(new_n8367_), .B1(\A[90] ), .Y(new_n9042_));
  OAI211 g08040(.A0(new_n9042_), .A1(new_n9041_), .B0(new_n9028_), .B1(new_n8361_), .Y(new_n9043_));
  NAND2  g08041(.A(new_n9030_), .B(new_n9029_), .Y(new_n9044_));
  AOI21  g08042(.A0(new_n9044_), .A1(new_n9043_), .B0(new_n9014_), .Y(new_n9045_));
  OAI21  g08043(.A0(new_n9045_), .A1(new_n9036_), .B0(new_n9040_), .Y(new_n9046_));
  AOI21  g08044(.A0(new_n9046_), .A1(new_n9034_), .B0(new_n9013_), .Y(new_n9047_));
  NOR2   g08045(.A(new_n9045_), .B(new_n9036_), .Y(new_n9048_));
  NAND4  g08046(.A(new_n8994_), .B(new_n9023_), .C(new_n9022_), .D(new_n9024_), .Y(new_n9049_));
  OAI21  g08047(.A0(new_n9022_), .A1(new_n9014_), .B0(new_n9032_), .Y(new_n9050_));
  OAI22  g08048(.A0(new_n9050_), .A1(new_n9049_), .B0(new_n9048_), .B1(new_n9040_), .Y(new_n9051_));
  AOI21  g08049(.A0(new_n9051_), .A1(new_n9013_), .B0(new_n9047_), .Y(new_n9052_));
  OAI21  g08050(.A0(new_n8993_), .A1(new_n8988_), .B0(new_n9052_), .Y(new_n9053_));
  XOR2   g08051(.A(new_n9048_), .B(new_n9033_), .Y(new_n9054_));
  NAND2  g08052(.A(new_n9051_), .B(new_n9013_), .Y(new_n9055_));
  OAI21  g08053(.A0(new_n9054_), .A1(new_n9013_), .B0(new_n9055_), .Y(new_n9056_));
  AOI211 g08054(.A0(new_n8981_), .A1(new_n8939_), .B(new_n8991_), .C(new_n8977_), .Y(new_n9057_));
  NOR2   g08055(.A(new_n8992_), .B(new_n8987_), .Y(new_n9058_));
  OAI21  g08056(.A0(new_n9058_), .A1(new_n9057_), .B0(new_n9056_), .Y(new_n9059_));
  NAND2  g08057(.A(new_n9059_), .B(new_n9053_), .Y(new_n9060_));
  AOI21  g08058(.A0(new_n8919_), .A1(new_n8907_), .B0(new_n9060_), .Y(new_n9061_));
  XOR2   g08059(.A(new_n8351_), .B(new_n8349_), .Y(new_n9062_));
  NOR2   g08060(.A(new_n8351_), .B(new_n8349_), .Y(new_n9063_));
  AOI21  g08061(.A0(new_n8937_), .A1(new_n9062_), .B0(new_n9063_), .Y(new_n9064_));
  XOR2   g08062(.A(new_n8937_), .B(new_n9062_), .Y(new_n9065_));
  OAI21  g08063(.A0(new_n9064_), .A1(new_n8968_), .B0(new_n9065_), .Y(new_n9066_));
  OAI21  g08064(.A0(new_n8952_), .A1(new_n8944_), .B0(new_n8953_), .Y(new_n9067_));
  XOR2   g08065(.A(new_n9067_), .B(new_n8963_), .Y(new_n9068_));
  NAND2  g08066(.A(new_n9068_), .B(new_n9066_), .Y(new_n9069_));
  NAND2  g08067(.A(new_n8981_), .B(new_n8939_), .Y(new_n9070_));
  NAND3  g08068(.A(new_n8991_), .B(new_n9070_), .C(new_n9069_), .Y(new_n9071_));
  NAND2  g08069(.A(new_n8974_), .B(new_n8973_), .Y(new_n9072_));
  NOR4   g08070(.A(new_n8968_), .B(new_n8966_), .C(new_n9072_), .D(new_n8944_), .Y(new_n9073_));
  OAI211 g08071(.A0(new_n8952_), .A1(new_n8944_), .B0(new_n9073_), .B1(new_n8962_), .Y(new_n9074_));
  AOI21  g08072(.A0(new_n9074_), .A1(new_n8978_), .B0(new_n9066_), .Y(new_n9075_));
  OAI21  g08073(.A0(new_n9075_), .A1(new_n8977_), .B0(new_n8987_), .Y(new_n9076_));
  AOI21  g08074(.A0(new_n9076_), .A1(new_n9071_), .B0(new_n9056_), .Y(new_n9077_));
  NAND3  g08075(.A(new_n8987_), .B(new_n9070_), .C(new_n9069_), .Y(new_n9078_));
  OAI21  g08076(.A0(new_n8992_), .A1(new_n8987_), .B0(new_n9078_), .Y(new_n9079_));
  AOI21  g08077(.A0(new_n9079_), .A1(new_n9056_), .B0(new_n9077_), .Y(new_n9080_));
  AOI21  g08078(.A0(new_n8904_), .A1(new_n8892_), .B0(new_n8906_), .Y(new_n9081_));
  NAND2  g08079(.A(new_n9081_), .B(new_n8889_), .Y(new_n9082_));
  OAI21  g08080(.A0(new_n8917_), .A1(new_n8914_), .B0(new_n8906_), .Y(new_n9083_));
  AOI21  g08081(.A0(new_n9083_), .A1(new_n9082_), .B0(new_n9080_), .Y(new_n9084_));
  NOR2   g08082(.A(new_n9084_), .B(new_n9061_), .Y(new_n9085_));
  OAI21  g08083(.A0(new_n8755_), .A1(new_n8748_), .B0(new_n9085_), .Y(new_n9086_));
  NOR3   g08084(.A(new_n8918_), .B(new_n8917_), .C(new_n8914_), .Y(new_n9087_));
  AOI21  g08085(.A0(new_n8905_), .A1(new_n8889_), .B0(new_n8906_), .Y(new_n9088_));
  OAI21  g08086(.A0(new_n9088_), .A1(new_n9087_), .B0(new_n9080_), .Y(new_n9089_));
  NOR3   g08087(.A(new_n8906_), .B(new_n8917_), .C(new_n8914_), .Y(new_n9090_));
  AOI21  g08088(.A0(new_n8905_), .A1(new_n8889_), .B0(new_n8918_), .Y(new_n9091_));
  OAI21  g08089(.A0(new_n9091_), .A1(new_n9090_), .B0(new_n9060_), .Y(new_n9092_));
  NAND2  g08090(.A(new_n9092_), .B(new_n9089_), .Y(new_n9093_));
  NOR3   g08091(.A(new_n8746_), .B(new_n8745_), .C(new_n8734_), .Y(new_n9094_));
  AOI21  g08092(.A0(new_n8754_), .A1(new_n8751_), .B0(new_n8747_), .Y(new_n9095_));
  OAI21  g08093(.A0(new_n9095_), .A1(new_n9094_), .B0(new_n9093_), .Y(new_n9096_));
  NAND2  g08094(.A(new_n9096_), .B(new_n9086_), .Y(new_n9097_));
  AOI21  g08095(.A0(new_n8406_), .A1(new_n8398_), .B0(new_n9097_), .Y(new_n9098_));
  NAND3  g08096(.A(new_n8746_), .B(new_n8754_), .C(new_n8751_), .Y(new_n9099_));
  OAI21  g08097(.A0(new_n8745_), .A1(new_n8734_), .B0(new_n8747_), .Y(new_n9100_));
  AOI21  g08098(.A0(new_n9100_), .A1(new_n9099_), .B0(new_n9093_), .Y(new_n9101_));
  NAND3  g08099(.A(new_n8747_), .B(new_n8754_), .C(new_n8751_), .Y(new_n9102_));
  OAI21  g08100(.A0(new_n8745_), .A1(new_n8734_), .B0(new_n8746_), .Y(new_n9103_));
  AOI21  g08101(.A0(new_n9103_), .A1(new_n9102_), .B0(new_n9085_), .Y(new_n9104_));
  NOR2   g08102(.A(new_n9104_), .B(new_n9101_), .Y(new_n9105_));
  NAND3  g08103(.A(new_n8405_), .B(new_n8069_), .C(new_n8059_), .Y(new_n9106_));
  OAI21  g08104(.A0(new_n8404_), .A1(new_n8401_), .B0(new_n8397_), .Y(new_n9107_));
  AOI21  g08105(.A0(new_n9107_), .A1(new_n9106_), .B0(new_n9105_), .Y(new_n9108_));
  NOR2   g08106(.A(new_n9108_), .B(new_n9098_), .Y(new_n9109_));
  INV    g08107(.A(\A[333] ), .Y(new_n9110_));
  INV    g08108(.A(\A[331] ), .Y(new_n9111_));
  NAND2  g08109(.A(\A[332] ), .B(new_n9111_), .Y(new_n9112_));
  INV    g08110(.A(\A[332] ), .Y(new_n9113_));
  AOI21  g08111(.A0(new_n9113_), .A1(\A[331] ), .B0(new_n9110_), .Y(new_n9114_));
  XOR2   g08112(.A(\A[332] ), .B(\A[331] ), .Y(new_n9115_));
  AOI22  g08113(.A0(new_n9115_), .A1(new_n9110_), .B0(new_n9114_), .B1(new_n9112_), .Y(new_n9116_));
  INV    g08114(.A(\A[336] ), .Y(new_n9117_));
  INV    g08115(.A(\A[334] ), .Y(new_n9118_));
  NAND2  g08116(.A(\A[335] ), .B(new_n9118_), .Y(new_n9119_));
  INV    g08117(.A(\A[335] ), .Y(new_n9120_));
  AOI21  g08118(.A0(new_n9120_), .A1(\A[334] ), .B0(new_n9117_), .Y(new_n9121_));
  XOR2   g08119(.A(\A[335] ), .B(\A[334] ), .Y(new_n9122_));
  AOI22  g08120(.A0(new_n9122_), .A1(new_n9117_), .B0(new_n9121_), .B1(new_n9119_), .Y(new_n9123_));
  NOR2   g08121(.A(new_n9123_), .B(new_n9116_), .Y(new_n9124_));
  XOR2   g08122(.A(\A[335] ), .B(new_n9118_), .Y(new_n9125_));
  NAND2  g08123(.A(\A[335] ), .B(\A[334] ), .Y(new_n9126_));
  OAI21  g08124(.A0(new_n9125_), .A1(new_n9117_), .B0(new_n9126_), .Y(new_n9127_));
  NOR2   g08125(.A(new_n9113_), .B(new_n9111_), .Y(new_n9128_));
  AOI21  g08126(.A0(new_n9115_), .A1(\A[333] ), .B0(new_n9128_), .Y(new_n9129_));
  XOR2   g08127(.A(new_n9129_), .B(new_n9127_), .Y(new_n9130_));
  XOR2   g08128(.A(new_n9130_), .B(new_n9124_), .Y(new_n9131_));
  XOR2   g08129(.A(new_n9123_), .B(new_n9116_), .Y(new_n9132_));
  NOR2   g08130(.A(new_n9113_), .B(\A[331] ), .Y(new_n9133_));
  OAI21  g08131(.A0(\A[332] ), .A1(new_n9111_), .B0(\A[333] ), .Y(new_n9134_));
  XOR2   g08132(.A(\A[332] ), .B(new_n9111_), .Y(new_n9135_));
  OAI22  g08133(.A0(new_n9135_), .A1(\A[333] ), .B0(new_n9134_), .B1(new_n9133_), .Y(new_n9136_));
  NOR2   g08134(.A(new_n9120_), .B(\A[334] ), .Y(new_n9137_));
  OAI21  g08135(.A0(\A[335] ), .A1(new_n9118_), .B0(\A[336] ), .Y(new_n9138_));
  OAI22  g08136(.A0(new_n9125_), .A1(\A[336] ), .B0(new_n9138_), .B1(new_n9137_), .Y(new_n9139_));
  NAND2  g08137(.A(new_n9139_), .B(new_n9136_), .Y(new_n9140_));
  NAND2  g08138(.A(\A[332] ), .B(\A[331] ), .Y(new_n9141_));
  OAI21  g08139(.A0(new_n9135_), .A1(new_n9110_), .B0(new_n9141_), .Y(new_n9142_));
  NAND2  g08140(.A(new_n9142_), .B(new_n9127_), .Y(new_n9143_));
  OAI21  g08141(.A0(new_n9130_), .A1(new_n9140_), .B0(new_n9143_), .Y(new_n9144_));
  AOI21  g08142(.A0(new_n9144_), .A1(new_n9132_), .B0(new_n9131_), .Y(new_n9145_));
  NAND2  g08143(.A(\A[341] ), .B(\A[340] ), .Y(new_n9146_));
  XOR2   g08144(.A(\A[341] ), .B(\A[340] ), .Y(new_n9147_));
  NAND2  g08145(.A(new_n9147_), .B(\A[342] ), .Y(new_n9148_));
  NAND2  g08146(.A(new_n9148_), .B(new_n9146_), .Y(new_n9149_));
  NAND2  g08147(.A(\A[338] ), .B(\A[337] ), .Y(new_n9150_));
  XOR2   g08148(.A(\A[338] ), .B(\A[337] ), .Y(new_n9151_));
  NAND2  g08149(.A(new_n9151_), .B(\A[339] ), .Y(new_n9152_));
  NAND2  g08150(.A(new_n9152_), .B(new_n9150_), .Y(new_n9153_));
  XOR2   g08151(.A(new_n9153_), .B(new_n9149_), .Y(new_n9154_));
  INV    g08152(.A(\A[339] ), .Y(new_n9155_));
  INV    g08153(.A(\A[337] ), .Y(new_n9156_));
  NAND2  g08154(.A(\A[338] ), .B(new_n9156_), .Y(new_n9157_));
  INV    g08155(.A(\A[338] ), .Y(new_n9158_));
  AOI21  g08156(.A0(new_n9158_), .A1(\A[337] ), .B0(new_n9155_), .Y(new_n9159_));
  AOI22  g08157(.A0(new_n9159_), .A1(new_n9157_), .B0(new_n9151_), .B1(new_n9155_), .Y(new_n9160_));
  INV    g08158(.A(\A[342] ), .Y(new_n9161_));
  INV    g08159(.A(\A[340] ), .Y(new_n9162_));
  NAND2  g08160(.A(\A[341] ), .B(new_n9162_), .Y(new_n9163_));
  INV    g08161(.A(\A[341] ), .Y(new_n9164_));
  AOI21  g08162(.A0(new_n9164_), .A1(\A[340] ), .B0(new_n9161_), .Y(new_n9165_));
  AOI22  g08163(.A0(new_n9165_), .A1(new_n9163_), .B0(new_n9147_), .B1(new_n9161_), .Y(new_n9166_));
  NOR2   g08164(.A(new_n9166_), .B(new_n9160_), .Y(new_n9167_));
  AOI22  g08165(.A0(new_n9152_), .A1(new_n9150_), .B0(new_n9148_), .B1(new_n9146_), .Y(new_n9168_));
  AOI21  g08166(.A0(new_n9167_), .A1(new_n9154_), .B0(new_n9168_), .Y(new_n9169_));
  XOR2   g08167(.A(new_n9167_), .B(new_n9154_), .Y(new_n9170_));
  NOR2   g08168(.A(new_n9158_), .B(\A[337] ), .Y(new_n9171_));
  OAI21  g08169(.A0(\A[338] ), .A1(new_n9156_), .B0(\A[339] ), .Y(new_n9172_));
  NAND2  g08170(.A(new_n9151_), .B(new_n9155_), .Y(new_n9173_));
  OAI21  g08171(.A0(new_n9172_), .A1(new_n9171_), .B0(new_n9173_), .Y(new_n9174_));
  XOR2   g08172(.A(new_n9166_), .B(new_n9174_), .Y(new_n9175_));
  NOR2   g08173(.A(new_n9164_), .B(\A[340] ), .Y(new_n9176_));
  OAI21  g08174(.A0(\A[341] ), .A1(new_n9162_), .B0(\A[342] ), .Y(new_n9177_));
  NAND2  g08175(.A(new_n9147_), .B(new_n9161_), .Y(new_n9178_));
  OAI21  g08176(.A0(new_n9177_), .A1(new_n9176_), .B0(new_n9178_), .Y(new_n9179_));
  NAND4  g08177(.A(new_n9179_), .B(new_n9174_), .C(new_n9153_), .D(new_n9149_), .Y(new_n9180_));
  NAND4  g08178(.A(new_n9142_), .B(new_n9127_), .C(new_n9139_), .D(new_n9136_), .Y(new_n9181_));
  XOR2   g08179(.A(new_n9166_), .B(new_n9160_), .Y(new_n9182_));
  NAND4  g08180(.A(new_n9182_), .B(new_n9181_), .C(new_n9180_), .D(new_n9132_), .Y(new_n9183_));
  OAI211 g08181(.A0(new_n9175_), .A1(new_n9169_), .B0(new_n9183_), .B1(new_n9170_), .Y(new_n9184_));
  NOR2   g08182(.A(new_n9158_), .B(new_n9156_), .Y(new_n9185_));
  AOI21  g08183(.A0(new_n9151_), .A1(\A[339] ), .B0(new_n9185_), .Y(new_n9186_));
  XOR2   g08184(.A(new_n9186_), .B(new_n9149_), .Y(new_n9187_));
  XOR2   g08185(.A(new_n9167_), .B(new_n9187_), .Y(new_n9188_));
  XOR2   g08186(.A(new_n9123_), .B(new_n9136_), .Y(new_n9189_));
  NOR2   g08187(.A(new_n9164_), .B(new_n9162_), .Y(new_n9190_));
  AOI21  g08188(.A0(new_n9147_), .A1(\A[342] ), .B0(new_n9190_), .Y(new_n9191_));
  NOR4   g08189(.A(new_n9166_), .B(new_n9160_), .C(new_n9186_), .D(new_n9191_), .Y(new_n9192_));
  NOR2   g08190(.A(new_n9120_), .B(new_n9118_), .Y(new_n9193_));
  AOI21  g08191(.A0(new_n9122_), .A1(\A[336] ), .B0(new_n9193_), .Y(new_n9194_));
  NOR4   g08192(.A(new_n9129_), .B(new_n9194_), .C(new_n9123_), .D(new_n9116_), .Y(new_n9195_));
  NOR4   g08193(.A(new_n9175_), .B(new_n9195_), .C(new_n9192_), .D(new_n9189_), .Y(new_n9196_));
  AOI221 g08194(.A0(new_n9151_), .A1(\A[339] ), .C0(new_n9185_), .B0(new_n9148_), .B1(new_n9146_), .Y(new_n9197_));
  AOI221 g08195(.A0(new_n9152_), .A1(new_n9150_), .C0(new_n9190_), .B0(new_n9147_), .B1(\A[342] ), .Y(new_n9198_));
  OAI211 g08196(.A0(new_n9198_), .A1(new_n9197_), .B0(new_n9179_), .B1(new_n9174_), .Y(new_n9199_));
  NAND2  g08197(.A(new_n9153_), .B(new_n9149_), .Y(new_n9200_));
  AOI21  g08198(.A0(new_n9200_), .A1(new_n9199_), .B0(new_n9175_), .Y(new_n9201_));
  OAI21  g08199(.A0(new_n9201_), .A1(new_n9188_), .B0(new_n9196_), .Y(new_n9202_));
  AOI21  g08200(.A0(new_n9202_), .A1(new_n9184_), .B0(new_n9145_), .Y(new_n9203_));
  XOR2   g08201(.A(new_n9130_), .B(new_n9140_), .Y(new_n9204_));
  XOR2   g08202(.A(new_n9129_), .B(new_n9194_), .Y(new_n9205_));
  NOR2   g08203(.A(new_n9129_), .B(new_n9194_), .Y(new_n9206_));
  AOI21  g08204(.A0(new_n9205_), .A1(new_n9124_), .B0(new_n9206_), .Y(new_n9207_));
  OAI21  g08205(.A0(new_n9207_), .A1(new_n9189_), .B0(new_n9204_), .Y(new_n9208_));
  OAI21  g08206(.A0(new_n9201_), .A1(new_n9188_), .B0(new_n9183_), .Y(new_n9209_));
  NOR2   g08207(.A(new_n9175_), .B(new_n9189_), .Y(new_n9210_));
  OAI211 g08208(.A0(new_n9179_), .A1(new_n9174_), .B0(new_n9153_), .B1(new_n9149_), .Y(new_n9211_));
  NAND4  g08209(.A(new_n9211_), .B(new_n9210_), .C(new_n9181_), .D(new_n9170_), .Y(new_n9212_));
  AOI21  g08210(.A0(new_n9212_), .A1(new_n9209_), .B0(new_n9208_), .Y(new_n9213_));
  NOR2   g08211(.A(new_n9175_), .B(new_n9192_), .Y(new_n9214_));
  XOR2   g08212(.A(new_n9123_), .B(new_n9116_), .Y(new_n9215_));
  XOR2   g08213(.A(new_n9215_), .B(new_n9214_), .Y(new_n9216_));
  INV    g08214(.A(\A[327] ), .Y(new_n9217_));
  INV    g08215(.A(\A[326] ), .Y(new_n9218_));
  NAND2  g08216(.A(new_n9218_), .B(\A[325] ), .Y(new_n9219_));
  INV    g08217(.A(\A[325] ), .Y(new_n9220_));
  AOI21  g08218(.A0(\A[326] ), .A1(new_n9220_), .B0(new_n9217_), .Y(new_n9221_));
  XOR2   g08219(.A(\A[326] ), .B(\A[325] ), .Y(new_n9222_));
  AOI22  g08220(.A0(new_n9222_), .A1(new_n9217_), .B0(new_n9221_), .B1(new_n9219_), .Y(new_n9223_));
  INV    g08221(.A(\A[330] ), .Y(new_n9224_));
  INV    g08222(.A(\A[329] ), .Y(new_n9225_));
  NAND2  g08223(.A(new_n9225_), .B(\A[328] ), .Y(new_n9226_));
  INV    g08224(.A(\A[328] ), .Y(new_n9227_));
  AOI21  g08225(.A0(\A[329] ), .A1(new_n9227_), .B0(new_n9224_), .Y(new_n9228_));
  XOR2   g08226(.A(\A[329] ), .B(\A[328] ), .Y(new_n9229_));
  AOI22  g08227(.A0(new_n9229_), .A1(new_n9224_), .B0(new_n9228_), .B1(new_n9226_), .Y(new_n9230_));
  NOR2   g08228(.A(new_n9225_), .B(new_n9227_), .Y(new_n9231_));
  AOI21  g08229(.A0(new_n9229_), .A1(\A[330] ), .B0(new_n9231_), .Y(new_n9232_));
  NOR2   g08230(.A(new_n9218_), .B(new_n9220_), .Y(new_n9233_));
  AOI21  g08231(.A0(new_n9222_), .A1(\A[327] ), .B0(new_n9233_), .Y(new_n9234_));
  XOR2   g08232(.A(new_n9230_), .B(new_n9223_), .Y(new_n9235_));
  INV    g08233(.A(\A[321] ), .Y(new_n9236_));
  INV    g08234(.A(\A[320] ), .Y(new_n9237_));
  NAND2  g08235(.A(new_n9237_), .B(\A[319] ), .Y(new_n9238_));
  INV    g08236(.A(\A[319] ), .Y(new_n9239_));
  AOI21  g08237(.A0(\A[320] ), .A1(new_n9239_), .B0(new_n9236_), .Y(new_n9240_));
  XOR2   g08238(.A(\A[320] ), .B(\A[319] ), .Y(new_n9241_));
  AOI22  g08239(.A0(new_n9241_), .A1(new_n9236_), .B0(new_n9240_), .B1(new_n9238_), .Y(new_n9242_));
  INV    g08240(.A(\A[324] ), .Y(new_n9243_));
  INV    g08241(.A(\A[323] ), .Y(new_n9244_));
  NAND2  g08242(.A(new_n9244_), .B(\A[322] ), .Y(new_n9245_));
  INV    g08243(.A(\A[322] ), .Y(new_n9246_));
  AOI21  g08244(.A0(\A[323] ), .A1(new_n9246_), .B0(new_n9243_), .Y(new_n9247_));
  XOR2   g08245(.A(\A[323] ), .B(\A[322] ), .Y(new_n9248_));
  AOI22  g08246(.A0(new_n9248_), .A1(new_n9243_), .B0(new_n9247_), .B1(new_n9245_), .Y(new_n9249_));
  NOR2   g08247(.A(new_n9244_), .B(new_n9246_), .Y(new_n9250_));
  AOI21  g08248(.A0(new_n9248_), .A1(\A[324] ), .B0(new_n9250_), .Y(new_n9251_));
  NOR2   g08249(.A(new_n9237_), .B(new_n9239_), .Y(new_n9252_));
  AOI21  g08250(.A0(new_n9241_), .A1(\A[321] ), .B0(new_n9252_), .Y(new_n9253_));
  XOR2   g08251(.A(new_n9249_), .B(new_n9242_), .Y(new_n9254_));
  XOR2   g08252(.A(new_n9254_), .B(new_n9235_), .Y(new_n9255_));
  NAND2  g08253(.A(new_n9255_), .B(new_n9216_), .Y(new_n9256_));
  NOR3   g08254(.A(new_n9256_), .B(new_n9213_), .C(new_n9203_), .Y(new_n9257_));
  OAI21  g08255(.A0(new_n9175_), .A1(new_n9169_), .B0(new_n9170_), .Y(new_n9258_));
  XOR2   g08256(.A(new_n9258_), .B(new_n9183_), .Y(new_n9259_));
  NAND2  g08257(.A(new_n9259_), .B(new_n9208_), .Y(new_n9260_));
  NAND2  g08258(.A(new_n9212_), .B(new_n9209_), .Y(new_n9261_));
  NAND2  g08259(.A(new_n9261_), .B(new_n9145_), .Y(new_n9262_));
  NAND2  g08260(.A(new_n9182_), .B(new_n9180_), .Y(new_n9263_));
  XOR2   g08261(.A(new_n9215_), .B(new_n9263_), .Y(new_n9264_));
  NOR2   g08262(.A(\A[326] ), .B(new_n9220_), .Y(new_n9265_));
  OAI21  g08263(.A0(new_n9218_), .A1(\A[325] ), .B0(\A[327] ), .Y(new_n9266_));
  NAND2  g08264(.A(new_n9222_), .B(new_n9217_), .Y(new_n9267_));
  OAI21  g08265(.A0(new_n9266_), .A1(new_n9265_), .B0(new_n9267_), .Y(new_n9268_));
  XOR2   g08266(.A(new_n9230_), .B(new_n9268_), .Y(new_n9269_));
  XOR2   g08267(.A(new_n9254_), .B(new_n9269_), .Y(new_n9270_));
  NOR2   g08268(.A(new_n9270_), .B(new_n9264_), .Y(new_n9271_));
  AOI21  g08269(.A0(new_n9262_), .A1(new_n9260_), .B0(new_n9271_), .Y(new_n9272_));
  XOR2   g08270(.A(new_n9249_), .B(new_n9242_), .Y(new_n9273_));
  XOR2   g08271(.A(\A[323] ), .B(new_n9246_), .Y(new_n9274_));
  NAND2  g08272(.A(\A[323] ), .B(\A[322] ), .Y(new_n9275_));
  OAI21  g08273(.A0(new_n9274_), .A1(new_n9243_), .B0(new_n9275_), .Y(new_n9276_));
  XOR2   g08274(.A(new_n9253_), .B(new_n9276_), .Y(new_n9277_));
  NOR2   g08275(.A(\A[320] ), .B(new_n9239_), .Y(new_n9278_));
  OAI21  g08276(.A0(new_n9237_), .A1(\A[319] ), .B0(\A[321] ), .Y(new_n9279_));
  XOR2   g08277(.A(\A[320] ), .B(new_n9239_), .Y(new_n9280_));
  OAI22  g08278(.A0(new_n9280_), .A1(\A[321] ), .B0(new_n9279_), .B1(new_n9278_), .Y(new_n9281_));
  NOR2   g08279(.A(\A[323] ), .B(new_n9246_), .Y(new_n9282_));
  OAI21  g08280(.A0(new_n9244_), .A1(\A[322] ), .B0(\A[324] ), .Y(new_n9283_));
  OAI22  g08281(.A0(new_n9274_), .A1(\A[324] ), .B0(new_n9283_), .B1(new_n9282_), .Y(new_n9284_));
  NAND2  g08282(.A(new_n9284_), .B(new_n9281_), .Y(new_n9285_));
  NAND2  g08283(.A(\A[320] ), .B(\A[319] ), .Y(new_n9286_));
  OAI21  g08284(.A0(new_n9280_), .A1(new_n9236_), .B0(new_n9286_), .Y(new_n9287_));
  NAND2  g08285(.A(new_n9287_), .B(new_n9276_), .Y(new_n9288_));
  OAI21  g08286(.A0(new_n9285_), .A1(new_n9277_), .B0(new_n9288_), .Y(new_n9289_));
  NOR2   g08287(.A(new_n9249_), .B(new_n9242_), .Y(new_n9290_));
  XOR2   g08288(.A(new_n9290_), .B(new_n9277_), .Y(new_n9291_));
  AOI21  g08289(.A0(new_n9289_), .A1(new_n9273_), .B0(new_n9291_), .Y(new_n9292_));
  XOR2   g08290(.A(new_n9230_), .B(new_n9268_), .Y(new_n9293_));
  XOR2   g08291(.A(new_n9234_), .B(new_n9232_), .Y(new_n9294_));
  NOR2   g08292(.A(new_n9230_), .B(new_n9223_), .Y(new_n9295_));
  NAND2  g08293(.A(\A[329] ), .B(\A[328] ), .Y(new_n9296_));
  NAND2  g08294(.A(new_n9229_), .B(\A[330] ), .Y(new_n9297_));
  NAND2  g08295(.A(\A[326] ), .B(\A[325] ), .Y(new_n9298_));
  NAND2  g08296(.A(new_n9222_), .B(\A[327] ), .Y(new_n9299_));
  AOI22  g08297(.A0(new_n9299_), .A1(new_n9298_), .B0(new_n9297_), .B1(new_n9296_), .Y(new_n9300_));
  AOI21  g08298(.A0(new_n9295_), .A1(new_n9294_), .B0(new_n9300_), .Y(new_n9301_));
  XOR2   g08299(.A(new_n9295_), .B(new_n9294_), .Y(new_n9302_));
  XOR2   g08300(.A(new_n9230_), .B(new_n9223_), .Y(new_n9303_));
  NOR2   g08301(.A(\A[329] ), .B(new_n9227_), .Y(new_n9304_));
  OAI21  g08302(.A0(new_n9225_), .A1(\A[328] ), .B0(\A[330] ), .Y(new_n9305_));
  NAND2  g08303(.A(new_n9229_), .B(new_n9224_), .Y(new_n9306_));
  OAI21  g08304(.A0(new_n9305_), .A1(new_n9304_), .B0(new_n9306_), .Y(new_n9307_));
  NAND2  g08305(.A(new_n9297_), .B(new_n9296_), .Y(new_n9308_));
  NAND2  g08306(.A(new_n9299_), .B(new_n9298_), .Y(new_n9309_));
  NAND4  g08307(.A(new_n9309_), .B(new_n9308_), .C(new_n9307_), .D(new_n9268_), .Y(new_n9310_));
  NAND4  g08308(.A(new_n9287_), .B(new_n9276_), .C(new_n9284_), .D(new_n9281_), .Y(new_n9311_));
  NAND4  g08309(.A(new_n9311_), .B(new_n9273_), .C(new_n9310_), .D(new_n9303_), .Y(new_n9312_));
  OAI211 g08310(.A0(new_n9301_), .A1(new_n9293_), .B0(new_n9312_), .B1(new_n9302_), .Y(new_n9313_));
  XOR2   g08311(.A(new_n9234_), .B(new_n9308_), .Y(new_n9314_));
  XOR2   g08312(.A(new_n9295_), .B(new_n9314_), .Y(new_n9315_));
  NOR4   g08313(.A(new_n9234_), .B(new_n9232_), .C(new_n9230_), .D(new_n9223_), .Y(new_n9316_));
  XOR2   g08314(.A(new_n9249_), .B(new_n9281_), .Y(new_n9317_));
  NOR3   g08315(.A(new_n9317_), .B(new_n9316_), .C(new_n9293_), .Y(new_n9318_));
  AOI221 g08316(.A0(new_n9297_), .A1(new_n9296_), .C0(new_n9233_), .B0(new_n9222_), .B1(\A[327] ), .Y(new_n9319_));
  AOI221 g08317(.A0(new_n9299_), .A1(new_n9298_), .C0(new_n9231_), .B0(new_n9229_), .B1(\A[330] ), .Y(new_n9320_));
  OAI211 g08318(.A0(new_n9320_), .A1(new_n9319_), .B0(new_n9307_), .B1(new_n9268_), .Y(new_n9321_));
  NAND2  g08319(.A(new_n9309_), .B(new_n9308_), .Y(new_n9322_));
  AOI21  g08320(.A0(new_n9322_), .A1(new_n9321_), .B0(new_n9293_), .Y(new_n9323_));
  OAI211 g08321(.A0(new_n9323_), .A1(new_n9315_), .B0(new_n9318_), .B1(new_n9311_), .Y(new_n9324_));
  AOI21  g08322(.A0(new_n9324_), .A1(new_n9313_), .B0(new_n9292_), .Y(new_n9325_));
  OAI21  g08323(.A0(new_n9323_), .A1(new_n9315_), .B0(new_n9312_), .Y(new_n9326_));
  NAND4  g08324(.A(new_n9273_), .B(new_n9302_), .C(new_n9301_), .D(new_n9303_), .Y(new_n9327_));
  OAI21  g08325(.A0(new_n9301_), .A1(new_n9293_), .B0(new_n9311_), .Y(new_n9328_));
  OAI21  g08326(.A0(new_n9328_), .A1(new_n9327_), .B0(new_n9326_), .Y(new_n9329_));
  AOI21  g08327(.A0(new_n9329_), .A1(new_n9292_), .B0(new_n9325_), .Y(new_n9330_));
  OAI21  g08328(.A0(new_n9272_), .A1(new_n9257_), .B0(new_n9330_), .Y(new_n9331_));
  XOR2   g08329(.A(new_n9253_), .B(new_n9251_), .Y(new_n9332_));
  NOR2   g08330(.A(new_n9253_), .B(new_n9251_), .Y(new_n9333_));
  AOI21  g08331(.A0(new_n9290_), .A1(new_n9332_), .B0(new_n9333_), .Y(new_n9334_));
  XOR2   g08332(.A(new_n9290_), .B(new_n9332_), .Y(new_n9335_));
  OAI21  g08333(.A0(new_n9334_), .A1(new_n9317_), .B0(new_n9335_), .Y(new_n9336_));
  OAI21  g08334(.A0(new_n9301_), .A1(new_n9293_), .B0(new_n9302_), .Y(new_n9337_));
  XOR2   g08335(.A(new_n9337_), .B(new_n9312_), .Y(new_n9338_));
  NAND2  g08336(.A(new_n9338_), .B(new_n9336_), .Y(new_n9339_));
  NAND2  g08337(.A(new_n9329_), .B(new_n9292_), .Y(new_n9340_));
  NAND2  g08338(.A(new_n9340_), .B(new_n9339_), .Y(new_n9341_));
  NAND2  g08339(.A(new_n9182_), .B(new_n9132_), .Y(new_n9342_));
  AOI211 g08340(.A0(new_n9166_), .A1(new_n9160_), .B(new_n9186_), .C(new_n9191_), .Y(new_n9343_));
  NOR4   g08341(.A(new_n9343_), .B(new_n9342_), .C(new_n9195_), .D(new_n9188_), .Y(new_n9344_));
  AOI21  g08342(.A0(new_n9258_), .A1(new_n9183_), .B0(new_n9344_), .Y(new_n9345_));
  OAI21  g08343(.A0(new_n9345_), .A1(new_n9208_), .B0(new_n9256_), .Y(new_n9346_));
  OAI21  g08344(.A0(new_n9213_), .A1(new_n9203_), .B0(new_n9271_), .Y(new_n9347_));
  OAI21  g08345(.A0(new_n9346_), .A1(new_n9203_), .B0(new_n9347_), .Y(new_n9348_));
  NAND2  g08346(.A(new_n9348_), .B(new_n9341_), .Y(new_n9349_));
  NAND2  g08347(.A(new_n9349_), .B(new_n9331_), .Y(new_n9350_));
  INV    g08348(.A(\A[344] ), .Y(new_n9351_));
  NOR2   g08349(.A(new_n9351_), .B(\A[343] ), .Y(new_n9352_));
  INV    g08350(.A(\A[343] ), .Y(new_n9353_));
  OAI21  g08351(.A0(\A[344] ), .A1(new_n9353_), .B0(\A[345] ), .Y(new_n9354_));
  XOR2   g08352(.A(\A[344] ), .B(new_n9353_), .Y(new_n9355_));
  OAI22  g08353(.A0(new_n9355_), .A1(\A[345] ), .B0(new_n9354_), .B1(new_n9352_), .Y(new_n9356_));
  INV    g08354(.A(\A[347] ), .Y(new_n9357_));
  NOR2   g08355(.A(new_n9357_), .B(\A[346] ), .Y(new_n9358_));
  INV    g08356(.A(\A[346] ), .Y(new_n9359_));
  OAI21  g08357(.A0(\A[347] ), .A1(new_n9359_), .B0(\A[348] ), .Y(new_n9360_));
  XOR2   g08358(.A(\A[347] ), .B(new_n9359_), .Y(new_n9361_));
  OAI22  g08359(.A0(new_n9361_), .A1(\A[348] ), .B0(new_n9360_), .B1(new_n9358_), .Y(new_n9362_));
  NAND2  g08360(.A(new_n9362_), .B(new_n9356_), .Y(new_n9363_));
  INV    g08361(.A(\A[348] ), .Y(new_n9364_));
  NAND2  g08362(.A(\A[347] ), .B(\A[346] ), .Y(new_n9365_));
  OAI21  g08363(.A0(new_n9361_), .A1(new_n9364_), .B0(new_n9365_), .Y(new_n9366_));
  XOR2   g08364(.A(\A[344] ), .B(\A[343] ), .Y(new_n9367_));
  NOR2   g08365(.A(new_n9351_), .B(new_n9353_), .Y(new_n9368_));
  AOI21  g08366(.A0(new_n9367_), .A1(\A[345] ), .B0(new_n9368_), .Y(new_n9369_));
  XOR2   g08367(.A(new_n9369_), .B(new_n9366_), .Y(new_n9370_));
  XOR2   g08368(.A(new_n9370_), .B(new_n9363_), .Y(new_n9371_));
  NAND2  g08369(.A(\A[347] ), .B(new_n9359_), .Y(new_n9372_));
  AOI21  g08370(.A0(new_n9357_), .A1(\A[346] ), .B0(new_n9364_), .Y(new_n9373_));
  XOR2   g08371(.A(\A[347] ), .B(\A[346] ), .Y(new_n9374_));
  AOI22  g08372(.A0(new_n9374_), .A1(new_n9364_), .B0(new_n9373_), .B1(new_n9372_), .Y(new_n9375_));
  XOR2   g08373(.A(new_n9375_), .B(new_n9356_), .Y(new_n9376_));
  INV    g08374(.A(\A[345] ), .Y(new_n9377_));
  NAND2  g08375(.A(\A[344] ), .B(new_n9353_), .Y(new_n9378_));
  AOI21  g08376(.A0(new_n9351_), .A1(\A[343] ), .B0(new_n9377_), .Y(new_n9379_));
  AOI22  g08377(.A0(new_n9367_), .A1(new_n9377_), .B0(new_n9379_), .B1(new_n9378_), .Y(new_n9380_));
  NOR2   g08378(.A(new_n9375_), .B(new_n9380_), .Y(new_n9381_));
  NOR2   g08379(.A(new_n9357_), .B(new_n9359_), .Y(new_n9382_));
  AOI21  g08380(.A0(new_n9374_), .A1(\A[348] ), .B0(new_n9382_), .Y(new_n9383_));
  XOR2   g08381(.A(new_n9369_), .B(new_n9383_), .Y(new_n9384_));
  NOR2   g08382(.A(new_n9369_), .B(new_n9383_), .Y(new_n9385_));
  AOI21  g08383(.A0(new_n9384_), .A1(new_n9381_), .B0(new_n9385_), .Y(new_n9386_));
  OAI21  g08384(.A0(new_n9386_), .A1(new_n9376_), .B0(new_n9371_), .Y(new_n9387_));
  XOR2   g08385(.A(new_n9375_), .B(new_n9380_), .Y(new_n9388_));
  NAND2  g08386(.A(\A[353] ), .B(\A[352] ), .Y(new_n9389_));
  XOR2   g08387(.A(\A[353] ), .B(\A[352] ), .Y(new_n9390_));
  NAND2  g08388(.A(new_n9390_), .B(\A[354] ), .Y(new_n9391_));
  NAND2  g08389(.A(new_n9391_), .B(new_n9389_), .Y(new_n9392_));
  NAND2  g08390(.A(\A[350] ), .B(\A[349] ), .Y(new_n9393_));
  XOR2   g08391(.A(\A[350] ), .B(\A[349] ), .Y(new_n9394_));
  NAND2  g08392(.A(new_n9394_), .B(\A[351] ), .Y(new_n9395_));
  NAND2  g08393(.A(new_n9395_), .B(new_n9393_), .Y(new_n9396_));
  INV    g08394(.A(\A[350] ), .Y(new_n9397_));
  NOR2   g08395(.A(new_n9397_), .B(\A[349] ), .Y(new_n9398_));
  INV    g08396(.A(\A[349] ), .Y(new_n9399_));
  OAI21  g08397(.A0(\A[350] ), .A1(new_n9399_), .B0(\A[351] ), .Y(new_n9400_));
  INV    g08398(.A(\A[351] ), .Y(new_n9401_));
  NAND2  g08399(.A(new_n9394_), .B(new_n9401_), .Y(new_n9402_));
  OAI21  g08400(.A0(new_n9400_), .A1(new_n9398_), .B0(new_n9402_), .Y(new_n9403_));
  INV    g08401(.A(\A[353] ), .Y(new_n9404_));
  NOR2   g08402(.A(new_n9404_), .B(\A[352] ), .Y(new_n9405_));
  INV    g08403(.A(\A[352] ), .Y(new_n9406_));
  OAI21  g08404(.A0(\A[353] ), .A1(new_n9406_), .B0(\A[354] ), .Y(new_n9407_));
  INV    g08405(.A(\A[354] ), .Y(new_n9408_));
  NAND2  g08406(.A(new_n9390_), .B(new_n9408_), .Y(new_n9409_));
  OAI21  g08407(.A0(new_n9407_), .A1(new_n9405_), .B0(new_n9409_), .Y(new_n9410_));
  NAND4  g08408(.A(new_n9410_), .B(new_n9403_), .C(new_n9396_), .D(new_n9392_), .Y(new_n9411_));
  NAND2  g08409(.A(\A[344] ), .B(\A[343] ), .Y(new_n9412_));
  OAI21  g08410(.A0(new_n9355_), .A1(new_n9377_), .B0(new_n9412_), .Y(new_n9413_));
  NAND4  g08411(.A(new_n9413_), .B(new_n9366_), .C(new_n9362_), .D(new_n9356_), .Y(new_n9414_));
  NAND2  g08412(.A(\A[350] ), .B(new_n9399_), .Y(new_n9415_));
  AOI21  g08413(.A0(new_n9397_), .A1(\A[349] ), .B0(new_n9401_), .Y(new_n9416_));
  AOI22  g08414(.A0(new_n9416_), .A1(new_n9415_), .B0(new_n9394_), .B1(new_n9401_), .Y(new_n9417_));
  NAND2  g08415(.A(\A[353] ), .B(new_n9406_), .Y(new_n9418_));
  AOI21  g08416(.A0(new_n9404_), .A1(\A[352] ), .B0(new_n9408_), .Y(new_n9419_));
  AOI22  g08417(.A0(new_n9419_), .A1(new_n9418_), .B0(new_n9390_), .B1(new_n9408_), .Y(new_n9420_));
  XOR2   g08418(.A(new_n9420_), .B(new_n9417_), .Y(new_n9421_));
  NAND4  g08419(.A(new_n9421_), .B(new_n9414_), .C(new_n9411_), .D(new_n9388_), .Y(new_n9422_));
  XOR2   g08420(.A(new_n9396_), .B(new_n9392_), .Y(new_n9423_));
  NOR2   g08421(.A(new_n9420_), .B(new_n9417_), .Y(new_n9424_));
  AOI22  g08422(.A0(new_n9395_), .A1(new_n9393_), .B0(new_n9391_), .B1(new_n9389_), .Y(new_n9425_));
  AOI21  g08423(.A0(new_n9424_), .A1(new_n9423_), .B0(new_n9425_), .Y(new_n9426_));
  XOR2   g08424(.A(new_n9424_), .B(new_n9423_), .Y(new_n9427_));
  XOR2   g08425(.A(new_n9420_), .B(new_n9403_), .Y(new_n9428_));
  OAI21  g08426(.A0(new_n9428_), .A1(new_n9426_), .B0(new_n9427_), .Y(new_n9429_));
  XOR2   g08427(.A(new_n9429_), .B(new_n9422_), .Y(new_n9430_));
  NAND2  g08428(.A(new_n9410_), .B(new_n9403_), .Y(new_n9431_));
  XOR2   g08429(.A(new_n9431_), .B(new_n9423_), .Y(new_n9432_));
  NOR2   g08430(.A(new_n9397_), .B(new_n9399_), .Y(new_n9433_));
  AOI221 g08431(.A0(new_n9394_), .A1(\A[351] ), .C0(new_n9433_), .B0(new_n9391_), .B1(new_n9389_), .Y(new_n9434_));
  NOR2   g08432(.A(new_n9404_), .B(new_n9406_), .Y(new_n9435_));
  AOI221 g08433(.A0(new_n9395_), .A1(new_n9393_), .C0(new_n9435_), .B0(new_n9390_), .B1(\A[354] ), .Y(new_n9436_));
  OAI211 g08434(.A0(new_n9436_), .A1(new_n9434_), .B0(new_n9410_), .B1(new_n9403_), .Y(new_n9437_));
  NAND2  g08435(.A(new_n9396_), .B(new_n9392_), .Y(new_n9438_));
  AOI21  g08436(.A0(new_n9438_), .A1(new_n9437_), .B0(new_n9428_), .Y(new_n9439_));
  OAI21  g08437(.A0(new_n9439_), .A1(new_n9432_), .B0(new_n9422_), .Y(new_n9440_));
  NOR2   g08438(.A(new_n9428_), .B(new_n9376_), .Y(new_n9441_));
  OAI211 g08439(.A0(new_n9410_), .A1(new_n9403_), .B0(new_n9396_), .B1(new_n9392_), .Y(new_n9442_));
  NAND4  g08440(.A(new_n9442_), .B(new_n9441_), .C(new_n9414_), .D(new_n9427_), .Y(new_n9443_));
  AOI21  g08441(.A0(new_n9443_), .A1(new_n9440_), .B0(new_n9387_), .Y(new_n9444_));
  AOI21  g08442(.A0(new_n9430_), .A1(new_n9387_), .B0(new_n9444_), .Y(new_n9445_));
  INV    g08443(.A(\A[357] ), .Y(new_n9446_));
  INV    g08444(.A(\A[355] ), .Y(new_n9447_));
  NAND2  g08445(.A(\A[356] ), .B(new_n9447_), .Y(new_n9448_));
  INV    g08446(.A(\A[356] ), .Y(new_n9449_));
  AOI21  g08447(.A0(new_n9449_), .A1(\A[355] ), .B0(new_n9446_), .Y(new_n9450_));
  XOR2   g08448(.A(\A[356] ), .B(\A[355] ), .Y(new_n9451_));
  AOI22  g08449(.A0(new_n9451_), .A1(new_n9446_), .B0(new_n9450_), .B1(new_n9448_), .Y(new_n9452_));
  INV    g08450(.A(\A[360] ), .Y(new_n9453_));
  INV    g08451(.A(\A[358] ), .Y(new_n9454_));
  NAND2  g08452(.A(\A[359] ), .B(new_n9454_), .Y(new_n9455_));
  INV    g08453(.A(\A[359] ), .Y(new_n9456_));
  AOI21  g08454(.A0(new_n9456_), .A1(\A[358] ), .B0(new_n9453_), .Y(new_n9457_));
  XOR2   g08455(.A(\A[359] ), .B(\A[358] ), .Y(new_n9458_));
  AOI22  g08456(.A0(new_n9458_), .A1(new_n9453_), .B0(new_n9457_), .B1(new_n9455_), .Y(new_n9459_));
  NOR2   g08457(.A(new_n9459_), .B(new_n9452_), .Y(new_n9460_));
  XOR2   g08458(.A(\A[359] ), .B(new_n9454_), .Y(new_n9461_));
  NAND2  g08459(.A(\A[359] ), .B(\A[358] ), .Y(new_n9462_));
  OAI21  g08460(.A0(new_n9461_), .A1(new_n9453_), .B0(new_n9462_), .Y(new_n9463_));
  NOR2   g08461(.A(new_n9449_), .B(new_n9447_), .Y(new_n9464_));
  AOI21  g08462(.A0(new_n9451_), .A1(\A[357] ), .B0(new_n9464_), .Y(new_n9465_));
  XOR2   g08463(.A(new_n9465_), .B(new_n9463_), .Y(new_n9466_));
  XOR2   g08464(.A(new_n9466_), .B(new_n9460_), .Y(new_n9467_));
  XOR2   g08465(.A(new_n9459_), .B(new_n9452_), .Y(new_n9468_));
  NOR2   g08466(.A(new_n9449_), .B(\A[355] ), .Y(new_n9469_));
  OAI21  g08467(.A0(\A[356] ), .A1(new_n9447_), .B0(\A[357] ), .Y(new_n9470_));
  XOR2   g08468(.A(\A[356] ), .B(new_n9447_), .Y(new_n9471_));
  OAI22  g08469(.A0(new_n9471_), .A1(\A[357] ), .B0(new_n9470_), .B1(new_n9469_), .Y(new_n9472_));
  NOR2   g08470(.A(new_n9456_), .B(\A[358] ), .Y(new_n9473_));
  OAI21  g08471(.A0(\A[359] ), .A1(new_n9454_), .B0(\A[360] ), .Y(new_n9474_));
  OAI22  g08472(.A0(new_n9461_), .A1(\A[360] ), .B0(new_n9474_), .B1(new_n9473_), .Y(new_n9475_));
  NAND2  g08473(.A(new_n9475_), .B(new_n9472_), .Y(new_n9476_));
  NAND2  g08474(.A(\A[356] ), .B(\A[355] ), .Y(new_n9477_));
  OAI21  g08475(.A0(new_n9471_), .A1(new_n9446_), .B0(new_n9477_), .Y(new_n9478_));
  NAND2  g08476(.A(new_n9478_), .B(new_n9463_), .Y(new_n9479_));
  OAI21  g08477(.A0(new_n9466_), .A1(new_n9476_), .B0(new_n9479_), .Y(new_n9480_));
  AOI21  g08478(.A0(new_n9480_), .A1(new_n9468_), .B0(new_n9467_), .Y(new_n9481_));
  NAND2  g08479(.A(\A[365] ), .B(\A[364] ), .Y(new_n9482_));
  XOR2   g08480(.A(\A[365] ), .B(\A[364] ), .Y(new_n9483_));
  NAND2  g08481(.A(new_n9483_), .B(\A[366] ), .Y(new_n9484_));
  NAND2  g08482(.A(new_n9484_), .B(new_n9482_), .Y(new_n9485_));
  NAND2  g08483(.A(\A[362] ), .B(\A[361] ), .Y(new_n9486_));
  XOR2   g08484(.A(\A[362] ), .B(\A[361] ), .Y(new_n9487_));
  NAND2  g08485(.A(new_n9487_), .B(\A[363] ), .Y(new_n9488_));
  NAND2  g08486(.A(new_n9488_), .B(new_n9486_), .Y(new_n9489_));
  XOR2   g08487(.A(new_n9489_), .B(new_n9485_), .Y(new_n9490_));
  INV    g08488(.A(\A[363] ), .Y(new_n9491_));
  INV    g08489(.A(\A[361] ), .Y(new_n9492_));
  NAND2  g08490(.A(\A[362] ), .B(new_n9492_), .Y(new_n9493_));
  INV    g08491(.A(\A[362] ), .Y(new_n9494_));
  AOI21  g08492(.A0(new_n9494_), .A1(\A[361] ), .B0(new_n9491_), .Y(new_n9495_));
  AOI22  g08493(.A0(new_n9495_), .A1(new_n9493_), .B0(new_n9487_), .B1(new_n9491_), .Y(new_n9496_));
  INV    g08494(.A(\A[366] ), .Y(new_n9497_));
  INV    g08495(.A(\A[364] ), .Y(new_n9498_));
  NAND2  g08496(.A(\A[365] ), .B(new_n9498_), .Y(new_n9499_));
  INV    g08497(.A(\A[365] ), .Y(new_n9500_));
  AOI21  g08498(.A0(new_n9500_), .A1(\A[364] ), .B0(new_n9497_), .Y(new_n9501_));
  AOI22  g08499(.A0(new_n9501_), .A1(new_n9499_), .B0(new_n9483_), .B1(new_n9497_), .Y(new_n9502_));
  NOR2   g08500(.A(new_n9502_), .B(new_n9496_), .Y(new_n9503_));
  AOI22  g08501(.A0(new_n9488_), .A1(new_n9486_), .B0(new_n9484_), .B1(new_n9482_), .Y(new_n9504_));
  AOI21  g08502(.A0(new_n9503_), .A1(new_n9490_), .B0(new_n9504_), .Y(new_n9505_));
  XOR2   g08503(.A(new_n9503_), .B(new_n9490_), .Y(new_n9506_));
  NOR2   g08504(.A(new_n9494_), .B(\A[361] ), .Y(new_n9507_));
  OAI21  g08505(.A0(\A[362] ), .A1(new_n9492_), .B0(\A[363] ), .Y(new_n9508_));
  NAND2  g08506(.A(new_n9487_), .B(new_n9491_), .Y(new_n9509_));
  OAI21  g08507(.A0(new_n9508_), .A1(new_n9507_), .B0(new_n9509_), .Y(new_n9510_));
  XOR2   g08508(.A(new_n9502_), .B(new_n9510_), .Y(new_n9511_));
  NOR2   g08509(.A(new_n9500_), .B(\A[364] ), .Y(new_n9512_));
  OAI21  g08510(.A0(\A[365] ), .A1(new_n9498_), .B0(\A[366] ), .Y(new_n9513_));
  NAND2  g08511(.A(new_n9483_), .B(new_n9497_), .Y(new_n9514_));
  OAI21  g08512(.A0(new_n9513_), .A1(new_n9512_), .B0(new_n9514_), .Y(new_n9515_));
  NAND4  g08513(.A(new_n9515_), .B(new_n9510_), .C(new_n9489_), .D(new_n9485_), .Y(new_n9516_));
  NAND4  g08514(.A(new_n9478_), .B(new_n9463_), .C(new_n9475_), .D(new_n9472_), .Y(new_n9517_));
  XOR2   g08515(.A(new_n9502_), .B(new_n9496_), .Y(new_n9518_));
  NAND4  g08516(.A(new_n9518_), .B(new_n9517_), .C(new_n9516_), .D(new_n9468_), .Y(new_n9519_));
  OAI211 g08517(.A0(new_n9511_), .A1(new_n9505_), .B0(new_n9519_), .B1(new_n9506_), .Y(new_n9520_));
  NOR2   g08518(.A(new_n9494_), .B(new_n9492_), .Y(new_n9521_));
  AOI21  g08519(.A0(new_n9487_), .A1(\A[363] ), .B0(new_n9521_), .Y(new_n9522_));
  XOR2   g08520(.A(new_n9522_), .B(new_n9485_), .Y(new_n9523_));
  XOR2   g08521(.A(new_n9503_), .B(new_n9523_), .Y(new_n9524_));
  XOR2   g08522(.A(new_n9459_), .B(new_n9472_), .Y(new_n9525_));
  NOR2   g08523(.A(new_n9500_), .B(new_n9498_), .Y(new_n9526_));
  AOI21  g08524(.A0(new_n9483_), .A1(\A[366] ), .B0(new_n9526_), .Y(new_n9527_));
  NOR4   g08525(.A(new_n9502_), .B(new_n9496_), .C(new_n9522_), .D(new_n9527_), .Y(new_n9528_));
  NOR2   g08526(.A(new_n9456_), .B(new_n9454_), .Y(new_n9529_));
  AOI21  g08527(.A0(new_n9458_), .A1(\A[360] ), .B0(new_n9529_), .Y(new_n9530_));
  NOR4   g08528(.A(new_n9465_), .B(new_n9530_), .C(new_n9459_), .D(new_n9452_), .Y(new_n9531_));
  NOR4   g08529(.A(new_n9511_), .B(new_n9531_), .C(new_n9528_), .D(new_n9525_), .Y(new_n9532_));
  AOI221 g08530(.A0(new_n9487_), .A1(\A[363] ), .C0(new_n9521_), .B0(new_n9484_), .B1(new_n9482_), .Y(new_n9533_));
  AOI221 g08531(.A0(new_n9488_), .A1(new_n9486_), .C0(new_n9526_), .B0(new_n9483_), .B1(\A[366] ), .Y(new_n9534_));
  OAI211 g08532(.A0(new_n9534_), .A1(new_n9533_), .B0(new_n9515_), .B1(new_n9510_), .Y(new_n9535_));
  NAND2  g08533(.A(new_n9489_), .B(new_n9485_), .Y(new_n9536_));
  AOI21  g08534(.A0(new_n9536_), .A1(new_n9535_), .B0(new_n9511_), .Y(new_n9537_));
  OAI21  g08535(.A0(new_n9537_), .A1(new_n9524_), .B0(new_n9532_), .Y(new_n9538_));
  AOI21  g08536(.A0(new_n9538_), .A1(new_n9520_), .B0(new_n9481_), .Y(new_n9539_));
  XOR2   g08537(.A(new_n9466_), .B(new_n9476_), .Y(new_n9540_));
  XOR2   g08538(.A(new_n9465_), .B(new_n9530_), .Y(new_n9541_));
  NOR2   g08539(.A(new_n9465_), .B(new_n9530_), .Y(new_n9542_));
  AOI21  g08540(.A0(new_n9541_), .A1(new_n9460_), .B0(new_n9542_), .Y(new_n9543_));
  OAI21  g08541(.A0(new_n9543_), .A1(new_n9525_), .B0(new_n9540_), .Y(new_n9544_));
  OAI21  g08542(.A0(new_n9537_), .A1(new_n9524_), .B0(new_n9519_), .Y(new_n9545_));
  NOR2   g08543(.A(new_n9511_), .B(new_n9525_), .Y(new_n9546_));
  OAI211 g08544(.A0(new_n9515_), .A1(new_n9510_), .B0(new_n9489_), .B1(new_n9485_), .Y(new_n9547_));
  NAND4  g08545(.A(new_n9547_), .B(new_n9546_), .C(new_n9517_), .D(new_n9506_), .Y(new_n9548_));
  AOI21  g08546(.A0(new_n9548_), .A1(new_n9545_), .B0(new_n9544_), .Y(new_n9549_));
  NOR2   g08547(.A(new_n9511_), .B(new_n9528_), .Y(new_n9550_));
  XOR2   g08548(.A(new_n9459_), .B(new_n9452_), .Y(new_n9551_));
  XOR2   g08549(.A(new_n9551_), .B(new_n9550_), .Y(new_n9552_));
  NAND2  g08550(.A(new_n9421_), .B(new_n9411_), .Y(new_n9553_));
  XOR2   g08551(.A(new_n9375_), .B(new_n9356_), .Y(new_n9554_));
  XOR2   g08552(.A(new_n9554_), .B(new_n9553_), .Y(new_n9555_));
  NAND2  g08553(.A(new_n9555_), .B(new_n9552_), .Y(new_n9556_));
  NOR3   g08554(.A(new_n9556_), .B(new_n9549_), .C(new_n9539_), .Y(new_n9557_));
  OAI21  g08555(.A0(new_n9511_), .A1(new_n9505_), .B0(new_n9506_), .Y(new_n9558_));
  XOR2   g08556(.A(new_n9558_), .B(new_n9519_), .Y(new_n9559_));
  NAND2  g08557(.A(new_n9559_), .B(new_n9544_), .Y(new_n9560_));
  NAND2  g08558(.A(new_n9548_), .B(new_n9545_), .Y(new_n9561_));
  NAND2  g08559(.A(new_n9561_), .B(new_n9481_), .Y(new_n9562_));
  NAND2  g08560(.A(new_n9518_), .B(new_n9516_), .Y(new_n9563_));
  XOR2   g08561(.A(new_n9551_), .B(new_n9563_), .Y(new_n9564_));
  XOR2   g08562(.A(new_n9375_), .B(new_n9380_), .Y(new_n9565_));
  XOR2   g08563(.A(new_n9565_), .B(new_n9553_), .Y(new_n9566_));
  NOR2   g08564(.A(new_n9566_), .B(new_n9564_), .Y(new_n9567_));
  AOI21  g08565(.A0(new_n9562_), .A1(new_n9560_), .B0(new_n9567_), .Y(new_n9568_));
  OAI21  g08566(.A0(new_n9568_), .A1(new_n9557_), .B0(new_n9445_), .Y(new_n9569_));
  XOR2   g08567(.A(new_n9370_), .B(new_n9381_), .Y(new_n9570_));
  NAND2  g08568(.A(new_n9413_), .B(new_n9366_), .Y(new_n9571_));
  OAI21  g08569(.A0(new_n9370_), .A1(new_n9363_), .B0(new_n9571_), .Y(new_n9572_));
  AOI21  g08570(.A0(new_n9572_), .A1(new_n9388_), .B0(new_n9570_), .Y(new_n9573_));
  NOR2   g08571(.A(new_n9439_), .B(new_n9432_), .Y(new_n9574_));
  XOR2   g08572(.A(new_n9574_), .B(new_n9422_), .Y(new_n9575_));
  NAND2  g08573(.A(new_n9443_), .B(new_n9440_), .Y(new_n9576_));
  NAND2  g08574(.A(new_n9576_), .B(new_n9573_), .Y(new_n9577_));
  OAI21  g08575(.A0(new_n9575_), .A1(new_n9573_), .B0(new_n9577_), .Y(new_n9578_));
  NAND2  g08576(.A(new_n9518_), .B(new_n9468_), .Y(new_n9579_));
  AOI211 g08577(.A0(new_n9502_), .A1(new_n9496_), .B(new_n9522_), .C(new_n9527_), .Y(new_n9580_));
  NOR4   g08578(.A(new_n9580_), .B(new_n9579_), .C(new_n9531_), .D(new_n9524_), .Y(new_n9581_));
  AOI21  g08579(.A0(new_n9558_), .A1(new_n9519_), .B0(new_n9581_), .Y(new_n9582_));
  OAI21  g08580(.A0(new_n9582_), .A1(new_n9544_), .B0(new_n9556_), .Y(new_n9583_));
  OAI21  g08581(.A0(new_n9549_), .A1(new_n9539_), .B0(new_n9567_), .Y(new_n9584_));
  OAI21  g08582(.A0(new_n9583_), .A1(new_n9539_), .B0(new_n9584_), .Y(new_n9585_));
  NAND2  g08583(.A(new_n9585_), .B(new_n9578_), .Y(new_n9586_));
  XOR2   g08584(.A(new_n9566_), .B(new_n9552_), .Y(new_n9587_));
  XOR2   g08585(.A(new_n9270_), .B(new_n9216_), .Y(new_n9588_));
  NOR2   g08586(.A(new_n9588_), .B(new_n9587_), .Y(new_n9589_));
  NAND3  g08587(.A(new_n9589_), .B(new_n9586_), .C(new_n9569_), .Y(new_n9590_));
  NAND3  g08588(.A(new_n9567_), .B(new_n9562_), .C(new_n9560_), .Y(new_n9591_));
  OAI21  g08589(.A0(new_n9549_), .A1(new_n9539_), .B0(new_n9556_), .Y(new_n9592_));
  AOI21  g08590(.A0(new_n9592_), .A1(new_n9591_), .B0(new_n9578_), .Y(new_n9593_));
  NAND3  g08591(.A(new_n9556_), .B(new_n9562_), .C(new_n9560_), .Y(new_n9594_));
  AOI21  g08592(.A0(new_n9584_), .A1(new_n9594_), .B0(new_n9445_), .Y(new_n9595_));
  INV    g08593(.A(new_n9589_), .Y(new_n9596_));
  OAI21  g08594(.A0(new_n9595_), .A1(new_n9593_), .B0(new_n9596_), .Y(new_n9597_));
  AOI21  g08595(.A0(new_n9597_), .A1(new_n9590_), .B0(new_n9350_), .Y(new_n9598_));
  NAND3  g08596(.A(new_n9271_), .B(new_n9262_), .C(new_n9260_), .Y(new_n9599_));
  OAI21  g08597(.A0(new_n9213_), .A1(new_n9203_), .B0(new_n9256_), .Y(new_n9600_));
  AOI21  g08598(.A0(new_n9600_), .A1(new_n9599_), .B0(new_n9341_), .Y(new_n9601_));
  AOI21  g08599(.A0(new_n9348_), .A1(new_n9341_), .B0(new_n9601_), .Y(new_n9602_));
  AOI21  g08600(.A0(new_n9585_), .A1(new_n9578_), .B0(new_n9589_), .Y(new_n9603_));
  NAND2  g08601(.A(new_n9603_), .B(new_n9569_), .Y(new_n9604_));
  OAI21  g08602(.A0(new_n9595_), .A1(new_n9593_), .B0(new_n9589_), .Y(new_n9605_));
  AOI21  g08603(.A0(new_n9605_), .A1(new_n9604_), .B0(new_n9602_), .Y(new_n9606_));
  XOR2   g08604(.A(new_n9588_), .B(new_n9587_), .Y(new_n9607_));
  INV    g08605(.A(new_n9607_), .Y(new_n9608_));
  INV    g08606(.A(\A[315] ), .Y(new_n9609_));
  INV    g08607(.A(\A[314] ), .Y(new_n9610_));
  NAND2  g08608(.A(new_n9610_), .B(\A[313] ), .Y(new_n9611_));
  INV    g08609(.A(\A[313] ), .Y(new_n9612_));
  AOI21  g08610(.A0(\A[314] ), .A1(new_n9612_), .B0(new_n9609_), .Y(new_n9613_));
  XOR2   g08611(.A(\A[314] ), .B(\A[313] ), .Y(new_n9614_));
  AOI22  g08612(.A0(new_n9614_), .A1(new_n9609_), .B0(new_n9613_), .B1(new_n9611_), .Y(new_n9615_));
  INV    g08613(.A(\A[318] ), .Y(new_n9616_));
  INV    g08614(.A(\A[317] ), .Y(new_n9617_));
  NAND2  g08615(.A(new_n9617_), .B(\A[316] ), .Y(new_n9618_));
  INV    g08616(.A(\A[316] ), .Y(new_n9619_));
  AOI21  g08617(.A0(\A[317] ), .A1(new_n9619_), .B0(new_n9616_), .Y(new_n9620_));
  XOR2   g08618(.A(\A[317] ), .B(\A[316] ), .Y(new_n9621_));
  AOI22  g08619(.A0(new_n9621_), .A1(new_n9616_), .B0(new_n9620_), .B1(new_n9618_), .Y(new_n9622_));
  NOR2   g08620(.A(new_n9617_), .B(new_n9619_), .Y(new_n9623_));
  AOI21  g08621(.A0(new_n9621_), .A1(\A[318] ), .B0(new_n9623_), .Y(new_n9624_));
  NOR2   g08622(.A(new_n9610_), .B(new_n9612_), .Y(new_n9625_));
  AOI21  g08623(.A0(new_n9614_), .A1(\A[315] ), .B0(new_n9625_), .Y(new_n9626_));
  XOR2   g08624(.A(new_n9622_), .B(new_n9615_), .Y(new_n9627_));
  INV    g08625(.A(\A[309] ), .Y(new_n9628_));
  INV    g08626(.A(\A[308] ), .Y(new_n9629_));
  NAND2  g08627(.A(new_n9629_), .B(\A[307] ), .Y(new_n9630_));
  INV    g08628(.A(\A[307] ), .Y(new_n9631_));
  AOI21  g08629(.A0(\A[308] ), .A1(new_n9631_), .B0(new_n9628_), .Y(new_n9632_));
  XOR2   g08630(.A(\A[308] ), .B(\A[307] ), .Y(new_n9633_));
  AOI22  g08631(.A0(new_n9633_), .A1(new_n9628_), .B0(new_n9632_), .B1(new_n9630_), .Y(new_n9634_));
  INV    g08632(.A(\A[312] ), .Y(new_n9635_));
  INV    g08633(.A(\A[311] ), .Y(new_n9636_));
  NAND2  g08634(.A(new_n9636_), .B(\A[310] ), .Y(new_n9637_));
  INV    g08635(.A(\A[310] ), .Y(new_n9638_));
  AOI21  g08636(.A0(\A[311] ), .A1(new_n9638_), .B0(new_n9635_), .Y(new_n9639_));
  XOR2   g08637(.A(\A[311] ), .B(\A[310] ), .Y(new_n9640_));
  AOI22  g08638(.A0(new_n9640_), .A1(new_n9635_), .B0(new_n9639_), .B1(new_n9637_), .Y(new_n9641_));
  NOR2   g08639(.A(new_n9636_), .B(new_n9638_), .Y(new_n9642_));
  AOI21  g08640(.A0(new_n9640_), .A1(\A[312] ), .B0(new_n9642_), .Y(new_n9643_));
  NOR2   g08641(.A(new_n9629_), .B(new_n9631_), .Y(new_n9644_));
  AOI21  g08642(.A0(new_n9633_), .A1(\A[309] ), .B0(new_n9644_), .Y(new_n9645_));
  XOR2   g08643(.A(new_n9641_), .B(new_n9634_), .Y(new_n9646_));
  XOR2   g08644(.A(new_n9646_), .B(new_n9627_), .Y(new_n9647_));
  INV    g08645(.A(\A[301] ), .Y(new_n9648_));
  NOR2   g08646(.A(\A[302] ), .B(new_n9648_), .Y(new_n9649_));
  INV    g08647(.A(\A[302] ), .Y(new_n9650_));
  OAI21  g08648(.A0(new_n9650_), .A1(\A[301] ), .B0(\A[303] ), .Y(new_n9651_));
  INV    g08649(.A(\A[303] ), .Y(new_n9652_));
  XOR2   g08650(.A(\A[302] ), .B(\A[301] ), .Y(new_n9653_));
  NAND2  g08651(.A(new_n9653_), .B(new_n9652_), .Y(new_n9654_));
  OAI21  g08652(.A0(new_n9651_), .A1(new_n9649_), .B0(new_n9654_), .Y(new_n9655_));
  INV    g08653(.A(\A[306] ), .Y(new_n9656_));
  INV    g08654(.A(\A[305] ), .Y(new_n9657_));
  NAND2  g08655(.A(new_n9657_), .B(\A[304] ), .Y(new_n9658_));
  INV    g08656(.A(\A[304] ), .Y(new_n9659_));
  AOI21  g08657(.A0(\A[305] ), .A1(new_n9659_), .B0(new_n9656_), .Y(new_n9660_));
  XOR2   g08658(.A(\A[305] ), .B(\A[304] ), .Y(new_n9661_));
  AOI22  g08659(.A0(new_n9661_), .A1(new_n9656_), .B0(new_n9660_), .B1(new_n9658_), .Y(new_n9662_));
  NOR2   g08660(.A(new_n9657_), .B(new_n9659_), .Y(new_n9663_));
  AOI21  g08661(.A0(new_n9661_), .A1(\A[306] ), .B0(new_n9663_), .Y(new_n9664_));
  NOR2   g08662(.A(new_n9650_), .B(new_n9648_), .Y(new_n9665_));
  AOI21  g08663(.A0(new_n9653_), .A1(\A[303] ), .B0(new_n9665_), .Y(new_n9666_));
  XOR2   g08664(.A(new_n9662_), .B(new_n9655_), .Y(new_n9667_));
  INV    g08665(.A(\A[297] ), .Y(new_n9668_));
  INV    g08666(.A(\A[296] ), .Y(new_n9669_));
  NAND2  g08667(.A(new_n9669_), .B(\A[295] ), .Y(new_n9670_));
  INV    g08668(.A(\A[295] ), .Y(new_n9671_));
  AOI21  g08669(.A0(\A[296] ), .A1(new_n9671_), .B0(new_n9668_), .Y(new_n9672_));
  XOR2   g08670(.A(\A[296] ), .B(\A[295] ), .Y(new_n9673_));
  AOI22  g08671(.A0(new_n9673_), .A1(new_n9668_), .B0(new_n9672_), .B1(new_n9670_), .Y(new_n9674_));
  INV    g08672(.A(\A[300] ), .Y(new_n9675_));
  INV    g08673(.A(\A[299] ), .Y(new_n9676_));
  NAND2  g08674(.A(new_n9676_), .B(\A[298] ), .Y(new_n9677_));
  INV    g08675(.A(\A[298] ), .Y(new_n9678_));
  AOI21  g08676(.A0(\A[299] ), .A1(new_n9678_), .B0(new_n9675_), .Y(new_n9679_));
  XOR2   g08677(.A(\A[299] ), .B(\A[298] ), .Y(new_n9680_));
  AOI22  g08678(.A0(new_n9680_), .A1(new_n9675_), .B0(new_n9679_), .B1(new_n9677_), .Y(new_n9681_));
  NOR2   g08679(.A(new_n9676_), .B(new_n9678_), .Y(new_n9682_));
  AOI21  g08680(.A0(new_n9680_), .A1(\A[300] ), .B0(new_n9682_), .Y(new_n9683_));
  NOR2   g08681(.A(new_n9669_), .B(new_n9671_), .Y(new_n9684_));
  AOI21  g08682(.A0(new_n9673_), .A1(\A[297] ), .B0(new_n9684_), .Y(new_n9685_));
  XOR2   g08683(.A(new_n9681_), .B(new_n9674_), .Y(new_n9686_));
  XOR2   g08684(.A(new_n9686_), .B(new_n9667_), .Y(new_n9687_));
  XOR2   g08685(.A(new_n9687_), .B(new_n9647_), .Y(new_n9688_));
  INV    g08686(.A(new_n9688_), .Y(new_n9689_));
  INV    g08687(.A(\A[291] ), .Y(new_n9690_));
  INV    g08688(.A(\A[290] ), .Y(new_n9691_));
  NAND2  g08689(.A(new_n9691_), .B(\A[289] ), .Y(new_n9692_));
  INV    g08690(.A(\A[289] ), .Y(new_n9693_));
  AOI21  g08691(.A0(\A[290] ), .A1(new_n9693_), .B0(new_n9690_), .Y(new_n9694_));
  XOR2   g08692(.A(\A[290] ), .B(\A[289] ), .Y(new_n9695_));
  AOI22  g08693(.A0(new_n9695_), .A1(new_n9690_), .B0(new_n9694_), .B1(new_n9692_), .Y(new_n9696_));
  INV    g08694(.A(\A[294] ), .Y(new_n9697_));
  INV    g08695(.A(\A[293] ), .Y(new_n9698_));
  NAND2  g08696(.A(new_n9698_), .B(\A[292] ), .Y(new_n9699_));
  INV    g08697(.A(\A[292] ), .Y(new_n9700_));
  AOI21  g08698(.A0(\A[293] ), .A1(new_n9700_), .B0(new_n9697_), .Y(new_n9701_));
  XOR2   g08699(.A(\A[293] ), .B(\A[292] ), .Y(new_n9702_));
  AOI22  g08700(.A0(new_n9702_), .A1(new_n9697_), .B0(new_n9701_), .B1(new_n9699_), .Y(new_n9703_));
  NOR2   g08701(.A(new_n9698_), .B(new_n9700_), .Y(new_n9704_));
  AOI21  g08702(.A0(new_n9702_), .A1(\A[294] ), .B0(new_n9704_), .Y(new_n9705_));
  NOR2   g08703(.A(new_n9691_), .B(new_n9693_), .Y(new_n9706_));
  AOI21  g08704(.A0(new_n9695_), .A1(\A[291] ), .B0(new_n9706_), .Y(new_n9707_));
  XOR2   g08705(.A(new_n9703_), .B(new_n9696_), .Y(new_n9708_));
  INV    g08706(.A(\A[285] ), .Y(new_n9709_));
  INV    g08707(.A(\A[284] ), .Y(new_n9710_));
  NAND2  g08708(.A(new_n9710_), .B(\A[283] ), .Y(new_n9711_));
  INV    g08709(.A(\A[283] ), .Y(new_n9712_));
  AOI21  g08710(.A0(\A[284] ), .A1(new_n9712_), .B0(new_n9709_), .Y(new_n9713_));
  XOR2   g08711(.A(\A[284] ), .B(\A[283] ), .Y(new_n9714_));
  AOI22  g08712(.A0(new_n9714_), .A1(new_n9709_), .B0(new_n9713_), .B1(new_n9711_), .Y(new_n9715_));
  INV    g08713(.A(\A[288] ), .Y(new_n9716_));
  INV    g08714(.A(\A[287] ), .Y(new_n9717_));
  NAND2  g08715(.A(new_n9717_), .B(\A[286] ), .Y(new_n9718_));
  INV    g08716(.A(\A[286] ), .Y(new_n9719_));
  AOI21  g08717(.A0(\A[287] ), .A1(new_n9719_), .B0(new_n9716_), .Y(new_n9720_));
  XOR2   g08718(.A(\A[287] ), .B(\A[286] ), .Y(new_n9721_));
  AOI22  g08719(.A0(new_n9721_), .A1(new_n9716_), .B0(new_n9720_), .B1(new_n9718_), .Y(new_n9722_));
  NOR2   g08720(.A(new_n9717_), .B(new_n9719_), .Y(new_n9723_));
  AOI21  g08721(.A0(new_n9721_), .A1(\A[288] ), .B0(new_n9723_), .Y(new_n9724_));
  NOR2   g08722(.A(new_n9710_), .B(new_n9712_), .Y(new_n9725_));
  AOI21  g08723(.A0(new_n9714_), .A1(\A[285] ), .B0(new_n9725_), .Y(new_n9726_));
  XOR2   g08724(.A(new_n9722_), .B(new_n9715_), .Y(new_n9727_));
  XOR2   g08725(.A(new_n9727_), .B(new_n9708_), .Y(new_n9728_));
  INV    g08726(.A(\A[277] ), .Y(new_n9729_));
  NOR2   g08727(.A(\A[278] ), .B(new_n9729_), .Y(new_n9730_));
  INV    g08728(.A(\A[278] ), .Y(new_n9731_));
  OAI21  g08729(.A0(new_n9731_), .A1(\A[277] ), .B0(\A[279] ), .Y(new_n9732_));
  INV    g08730(.A(\A[279] ), .Y(new_n9733_));
  XOR2   g08731(.A(\A[278] ), .B(\A[277] ), .Y(new_n9734_));
  NAND2  g08732(.A(new_n9734_), .B(new_n9733_), .Y(new_n9735_));
  OAI21  g08733(.A0(new_n9732_), .A1(new_n9730_), .B0(new_n9735_), .Y(new_n9736_));
  INV    g08734(.A(\A[282] ), .Y(new_n9737_));
  INV    g08735(.A(\A[281] ), .Y(new_n9738_));
  NAND2  g08736(.A(new_n9738_), .B(\A[280] ), .Y(new_n9739_));
  INV    g08737(.A(\A[280] ), .Y(new_n9740_));
  AOI21  g08738(.A0(\A[281] ), .A1(new_n9740_), .B0(new_n9737_), .Y(new_n9741_));
  XOR2   g08739(.A(\A[281] ), .B(\A[280] ), .Y(new_n9742_));
  AOI22  g08740(.A0(new_n9742_), .A1(new_n9737_), .B0(new_n9741_), .B1(new_n9739_), .Y(new_n9743_));
  NOR2   g08741(.A(new_n9738_), .B(new_n9740_), .Y(new_n9744_));
  AOI21  g08742(.A0(new_n9742_), .A1(\A[282] ), .B0(new_n9744_), .Y(new_n9745_));
  NOR2   g08743(.A(new_n9731_), .B(new_n9729_), .Y(new_n9746_));
  AOI21  g08744(.A0(new_n9734_), .A1(\A[279] ), .B0(new_n9746_), .Y(new_n9747_));
  XOR2   g08745(.A(new_n9743_), .B(new_n9736_), .Y(new_n9748_));
  INV    g08746(.A(\A[273] ), .Y(new_n9749_));
  INV    g08747(.A(\A[272] ), .Y(new_n9750_));
  NAND2  g08748(.A(new_n9750_), .B(\A[271] ), .Y(new_n9751_));
  INV    g08749(.A(\A[271] ), .Y(new_n9752_));
  AOI21  g08750(.A0(\A[272] ), .A1(new_n9752_), .B0(new_n9749_), .Y(new_n9753_));
  XOR2   g08751(.A(\A[272] ), .B(\A[271] ), .Y(new_n9754_));
  AOI22  g08752(.A0(new_n9754_), .A1(new_n9749_), .B0(new_n9753_), .B1(new_n9751_), .Y(new_n9755_));
  INV    g08753(.A(\A[276] ), .Y(new_n9756_));
  INV    g08754(.A(\A[275] ), .Y(new_n9757_));
  NAND2  g08755(.A(new_n9757_), .B(\A[274] ), .Y(new_n9758_));
  INV    g08756(.A(\A[274] ), .Y(new_n9759_));
  AOI21  g08757(.A0(\A[275] ), .A1(new_n9759_), .B0(new_n9756_), .Y(new_n9760_));
  XOR2   g08758(.A(\A[275] ), .B(\A[274] ), .Y(new_n9761_));
  AOI22  g08759(.A0(new_n9761_), .A1(new_n9756_), .B0(new_n9760_), .B1(new_n9758_), .Y(new_n9762_));
  NOR2   g08760(.A(new_n9757_), .B(new_n9759_), .Y(new_n9763_));
  AOI21  g08761(.A0(new_n9761_), .A1(\A[276] ), .B0(new_n9763_), .Y(new_n9764_));
  NOR2   g08762(.A(new_n9750_), .B(new_n9752_), .Y(new_n9765_));
  AOI21  g08763(.A0(new_n9754_), .A1(\A[273] ), .B0(new_n9765_), .Y(new_n9766_));
  XOR2   g08764(.A(new_n9762_), .B(new_n9755_), .Y(new_n9767_));
  XOR2   g08765(.A(new_n9767_), .B(new_n9748_), .Y(new_n9768_));
  XOR2   g08766(.A(new_n9768_), .B(new_n9728_), .Y(new_n9769_));
  XOR2   g08767(.A(new_n9769_), .B(new_n9689_), .Y(new_n9770_));
  NOR2   g08768(.A(new_n9770_), .B(new_n9608_), .Y(new_n9771_));
  INV    g08769(.A(new_n9771_), .Y(new_n9772_));
  NOR3   g08770(.A(new_n9772_), .B(new_n9606_), .C(new_n9598_), .Y(new_n9773_));
  NOR3   g08771(.A(new_n9596_), .B(new_n9595_), .C(new_n9593_), .Y(new_n9774_));
  AOI21  g08772(.A0(new_n9586_), .A1(new_n9569_), .B0(new_n9589_), .Y(new_n9775_));
  OAI21  g08773(.A0(new_n9775_), .A1(new_n9774_), .B0(new_n9602_), .Y(new_n9776_));
  NOR3   g08774(.A(new_n9589_), .B(new_n9595_), .C(new_n9593_), .Y(new_n9777_));
  AOI21  g08775(.A0(new_n9586_), .A1(new_n9569_), .B0(new_n9596_), .Y(new_n9778_));
  OAI21  g08776(.A0(new_n9778_), .A1(new_n9777_), .B0(new_n9350_), .Y(new_n9779_));
  AOI21  g08777(.A0(new_n9779_), .A1(new_n9776_), .B0(new_n9771_), .Y(new_n9780_));
  XOR2   g08778(.A(new_n9681_), .B(new_n9674_), .Y(new_n9781_));
  XOR2   g08779(.A(\A[299] ), .B(new_n9678_), .Y(new_n9782_));
  NAND2  g08780(.A(\A[299] ), .B(\A[298] ), .Y(new_n9783_));
  OAI21  g08781(.A0(new_n9782_), .A1(new_n9675_), .B0(new_n9783_), .Y(new_n9784_));
  XOR2   g08782(.A(new_n9685_), .B(new_n9784_), .Y(new_n9785_));
  NOR2   g08783(.A(\A[296] ), .B(new_n9671_), .Y(new_n9786_));
  OAI21  g08784(.A0(new_n9669_), .A1(\A[295] ), .B0(\A[297] ), .Y(new_n9787_));
  XOR2   g08785(.A(\A[296] ), .B(new_n9671_), .Y(new_n9788_));
  OAI22  g08786(.A0(new_n9788_), .A1(\A[297] ), .B0(new_n9787_), .B1(new_n9786_), .Y(new_n9789_));
  NOR2   g08787(.A(\A[299] ), .B(new_n9678_), .Y(new_n9790_));
  OAI21  g08788(.A0(new_n9676_), .A1(\A[298] ), .B0(\A[300] ), .Y(new_n9791_));
  OAI22  g08789(.A0(new_n9782_), .A1(\A[300] ), .B0(new_n9791_), .B1(new_n9790_), .Y(new_n9792_));
  NAND2  g08790(.A(new_n9792_), .B(new_n9789_), .Y(new_n9793_));
  NAND2  g08791(.A(\A[296] ), .B(\A[295] ), .Y(new_n9794_));
  OAI21  g08792(.A0(new_n9788_), .A1(new_n9668_), .B0(new_n9794_), .Y(new_n9795_));
  NAND2  g08793(.A(new_n9795_), .B(new_n9784_), .Y(new_n9796_));
  OAI21  g08794(.A0(new_n9793_), .A1(new_n9785_), .B0(new_n9796_), .Y(new_n9797_));
  NOR2   g08795(.A(new_n9681_), .B(new_n9674_), .Y(new_n9798_));
  XOR2   g08796(.A(new_n9798_), .B(new_n9785_), .Y(new_n9799_));
  AOI21  g08797(.A0(new_n9797_), .A1(new_n9781_), .B0(new_n9799_), .Y(new_n9800_));
  XOR2   g08798(.A(new_n9662_), .B(new_n9655_), .Y(new_n9801_));
  XOR2   g08799(.A(new_n9666_), .B(new_n9664_), .Y(new_n9802_));
  NAND2  g08800(.A(new_n9650_), .B(\A[301] ), .Y(new_n9803_));
  AOI21  g08801(.A0(\A[302] ), .A1(new_n9648_), .B0(new_n9652_), .Y(new_n9804_));
  AOI22  g08802(.A0(new_n9653_), .A1(new_n9652_), .B0(new_n9804_), .B1(new_n9803_), .Y(new_n9805_));
  NOR2   g08803(.A(new_n9662_), .B(new_n9805_), .Y(new_n9806_));
  NAND2  g08804(.A(\A[305] ), .B(\A[304] ), .Y(new_n9807_));
  NAND2  g08805(.A(new_n9661_), .B(\A[306] ), .Y(new_n9808_));
  NAND2  g08806(.A(\A[302] ), .B(\A[301] ), .Y(new_n9809_));
  NAND2  g08807(.A(new_n9653_), .B(\A[303] ), .Y(new_n9810_));
  AOI22  g08808(.A0(new_n9810_), .A1(new_n9809_), .B0(new_n9808_), .B1(new_n9807_), .Y(new_n9811_));
  AOI21  g08809(.A0(new_n9806_), .A1(new_n9802_), .B0(new_n9811_), .Y(new_n9812_));
  XOR2   g08810(.A(new_n9806_), .B(new_n9802_), .Y(new_n9813_));
  XOR2   g08811(.A(new_n9662_), .B(new_n9805_), .Y(new_n9814_));
  NOR2   g08812(.A(\A[305] ), .B(new_n9659_), .Y(new_n9815_));
  OAI21  g08813(.A0(new_n9657_), .A1(\A[304] ), .B0(\A[306] ), .Y(new_n9816_));
  NAND2  g08814(.A(new_n9661_), .B(new_n9656_), .Y(new_n9817_));
  OAI21  g08815(.A0(new_n9816_), .A1(new_n9815_), .B0(new_n9817_), .Y(new_n9818_));
  NAND2  g08816(.A(new_n9808_), .B(new_n9807_), .Y(new_n9819_));
  NAND2  g08817(.A(new_n9810_), .B(new_n9809_), .Y(new_n9820_));
  NAND4  g08818(.A(new_n9820_), .B(new_n9819_), .C(new_n9818_), .D(new_n9655_), .Y(new_n9821_));
  NAND4  g08819(.A(new_n9795_), .B(new_n9784_), .C(new_n9792_), .D(new_n9789_), .Y(new_n9822_));
  NAND4  g08820(.A(new_n9822_), .B(new_n9781_), .C(new_n9821_), .D(new_n9814_), .Y(new_n9823_));
  OAI211 g08821(.A0(new_n9812_), .A1(new_n9801_), .B0(new_n9823_), .B1(new_n9813_), .Y(new_n9824_));
  XOR2   g08822(.A(new_n9666_), .B(new_n9819_), .Y(new_n9825_));
  XOR2   g08823(.A(new_n9806_), .B(new_n9825_), .Y(new_n9826_));
  NOR4   g08824(.A(new_n9666_), .B(new_n9664_), .C(new_n9662_), .D(new_n9805_), .Y(new_n9827_));
  XOR2   g08825(.A(new_n9681_), .B(new_n9789_), .Y(new_n9828_));
  NOR4   g08826(.A(new_n9685_), .B(new_n9683_), .C(new_n9681_), .D(new_n9674_), .Y(new_n9829_));
  NOR4   g08827(.A(new_n9829_), .B(new_n9828_), .C(new_n9827_), .D(new_n9801_), .Y(new_n9830_));
  AOI221 g08828(.A0(new_n9808_), .A1(new_n9807_), .C0(new_n9665_), .B0(new_n9653_), .B1(\A[303] ), .Y(new_n9831_));
  AOI221 g08829(.A0(new_n9810_), .A1(new_n9809_), .C0(new_n9663_), .B0(new_n9661_), .B1(\A[306] ), .Y(new_n9832_));
  OAI211 g08830(.A0(new_n9832_), .A1(new_n9831_), .B0(new_n9818_), .B1(new_n9655_), .Y(new_n9833_));
  NAND2  g08831(.A(new_n9820_), .B(new_n9819_), .Y(new_n9834_));
  AOI21  g08832(.A0(new_n9834_), .A1(new_n9833_), .B0(new_n9801_), .Y(new_n9835_));
  OAI21  g08833(.A0(new_n9835_), .A1(new_n9826_), .B0(new_n9830_), .Y(new_n9836_));
  AOI21  g08834(.A0(new_n9836_), .A1(new_n9824_), .B0(new_n9800_), .Y(new_n9837_));
  NOR2   g08835(.A(new_n9835_), .B(new_n9826_), .Y(new_n9838_));
  NAND4  g08836(.A(new_n9781_), .B(new_n9813_), .C(new_n9812_), .D(new_n9814_), .Y(new_n9839_));
  OAI21  g08837(.A0(new_n9812_), .A1(new_n9801_), .B0(new_n9822_), .Y(new_n9840_));
  OAI22  g08838(.A0(new_n9840_), .A1(new_n9839_), .B0(new_n9838_), .B1(new_n9830_), .Y(new_n9841_));
  AOI21  g08839(.A0(new_n9841_), .A1(new_n9800_), .B0(new_n9837_), .Y(new_n9842_));
  XOR2   g08840(.A(new_n9641_), .B(new_n9634_), .Y(new_n9843_));
  XOR2   g08841(.A(\A[311] ), .B(new_n9638_), .Y(new_n9844_));
  NAND2  g08842(.A(\A[311] ), .B(\A[310] ), .Y(new_n9845_));
  OAI21  g08843(.A0(new_n9844_), .A1(new_n9635_), .B0(new_n9845_), .Y(new_n9846_));
  XOR2   g08844(.A(new_n9645_), .B(new_n9846_), .Y(new_n9847_));
  NOR2   g08845(.A(\A[308] ), .B(new_n9631_), .Y(new_n9848_));
  OAI21  g08846(.A0(new_n9629_), .A1(\A[307] ), .B0(\A[309] ), .Y(new_n9849_));
  XOR2   g08847(.A(\A[308] ), .B(new_n9631_), .Y(new_n9850_));
  OAI22  g08848(.A0(new_n9850_), .A1(\A[309] ), .B0(new_n9849_), .B1(new_n9848_), .Y(new_n9851_));
  NOR2   g08849(.A(\A[311] ), .B(new_n9638_), .Y(new_n9852_));
  OAI21  g08850(.A0(new_n9636_), .A1(\A[310] ), .B0(\A[312] ), .Y(new_n9853_));
  OAI22  g08851(.A0(new_n9844_), .A1(\A[312] ), .B0(new_n9853_), .B1(new_n9852_), .Y(new_n9854_));
  NAND2  g08852(.A(new_n9854_), .B(new_n9851_), .Y(new_n9855_));
  NAND2  g08853(.A(\A[308] ), .B(\A[307] ), .Y(new_n9856_));
  OAI21  g08854(.A0(new_n9850_), .A1(new_n9628_), .B0(new_n9856_), .Y(new_n9857_));
  NAND2  g08855(.A(new_n9857_), .B(new_n9846_), .Y(new_n9858_));
  OAI21  g08856(.A0(new_n9855_), .A1(new_n9847_), .B0(new_n9858_), .Y(new_n9859_));
  NOR2   g08857(.A(new_n9641_), .B(new_n9634_), .Y(new_n9860_));
  XOR2   g08858(.A(new_n9860_), .B(new_n9847_), .Y(new_n9861_));
  AOI21  g08859(.A0(new_n9859_), .A1(new_n9843_), .B0(new_n9861_), .Y(new_n9862_));
  NOR2   g08860(.A(\A[314] ), .B(new_n9612_), .Y(new_n9863_));
  OAI21  g08861(.A0(new_n9610_), .A1(\A[313] ), .B0(\A[315] ), .Y(new_n9864_));
  NAND2  g08862(.A(new_n9614_), .B(new_n9609_), .Y(new_n9865_));
  OAI21  g08863(.A0(new_n9864_), .A1(new_n9863_), .B0(new_n9865_), .Y(new_n9866_));
  XOR2   g08864(.A(new_n9622_), .B(new_n9866_), .Y(new_n9867_));
  XOR2   g08865(.A(new_n9626_), .B(new_n9624_), .Y(new_n9868_));
  NOR2   g08866(.A(new_n9622_), .B(new_n9615_), .Y(new_n9869_));
  NAND2  g08867(.A(\A[317] ), .B(\A[316] ), .Y(new_n9870_));
  NAND2  g08868(.A(new_n9621_), .B(\A[318] ), .Y(new_n9871_));
  NAND2  g08869(.A(\A[314] ), .B(\A[313] ), .Y(new_n9872_));
  NAND2  g08870(.A(new_n9614_), .B(\A[315] ), .Y(new_n9873_));
  AOI22  g08871(.A0(new_n9873_), .A1(new_n9872_), .B0(new_n9871_), .B1(new_n9870_), .Y(new_n9874_));
  AOI21  g08872(.A0(new_n9869_), .A1(new_n9868_), .B0(new_n9874_), .Y(new_n9875_));
  XOR2   g08873(.A(new_n9869_), .B(new_n9868_), .Y(new_n9876_));
  XOR2   g08874(.A(new_n9622_), .B(new_n9615_), .Y(new_n9877_));
  NOR2   g08875(.A(\A[317] ), .B(new_n9619_), .Y(new_n9878_));
  OAI21  g08876(.A0(new_n9617_), .A1(\A[316] ), .B0(\A[318] ), .Y(new_n9879_));
  NAND2  g08877(.A(new_n9621_), .B(new_n9616_), .Y(new_n9880_));
  OAI21  g08878(.A0(new_n9879_), .A1(new_n9878_), .B0(new_n9880_), .Y(new_n9881_));
  NAND2  g08879(.A(new_n9871_), .B(new_n9870_), .Y(new_n9882_));
  NAND2  g08880(.A(new_n9873_), .B(new_n9872_), .Y(new_n9883_));
  NAND4  g08881(.A(new_n9883_), .B(new_n9882_), .C(new_n9881_), .D(new_n9866_), .Y(new_n9884_));
  NAND4  g08882(.A(new_n9857_), .B(new_n9846_), .C(new_n9854_), .D(new_n9851_), .Y(new_n9885_));
  NAND4  g08883(.A(new_n9885_), .B(new_n9843_), .C(new_n9884_), .D(new_n9877_), .Y(new_n9886_));
  OAI211 g08884(.A0(new_n9875_), .A1(new_n9867_), .B0(new_n9886_), .B1(new_n9876_), .Y(new_n9887_));
  XOR2   g08885(.A(new_n9626_), .B(new_n9882_), .Y(new_n9888_));
  XOR2   g08886(.A(new_n9869_), .B(new_n9888_), .Y(new_n9889_));
  NOR4   g08887(.A(new_n9626_), .B(new_n9624_), .C(new_n9622_), .D(new_n9615_), .Y(new_n9890_));
  XOR2   g08888(.A(new_n9641_), .B(new_n9851_), .Y(new_n9891_));
  NOR4   g08889(.A(new_n9645_), .B(new_n9643_), .C(new_n9641_), .D(new_n9634_), .Y(new_n9892_));
  NOR4   g08890(.A(new_n9892_), .B(new_n9891_), .C(new_n9890_), .D(new_n9867_), .Y(new_n9893_));
  AOI221 g08891(.A0(new_n9871_), .A1(new_n9870_), .C0(new_n9625_), .B0(new_n9614_), .B1(\A[315] ), .Y(new_n9894_));
  AOI221 g08892(.A0(new_n9873_), .A1(new_n9872_), .C0(new_n9623_), .B0(new_n9621_), .B1(\A[318] ), .Y(new_n9895_));
  OAI211 g08893(.A0(new_n9895_), .A1(new_n9894_), .B0(new_n9881_), .B1(new_n9866_), .Y(new_n9896_));
  NAND2  g08894(.A(new_n9883_), .B(new_n9882_), .Y(new_n9897_));
  AOI21  g08895(.A0(new_n9897_), .A1(new_n9896_), .B0(new_n9867_), .Y(new_n9898_));
  OAI21  g08896(.A0(new_n9898_), .A1(new_n9889_), .B0(new_n9893_), .Y(new_n9899_));
  AOI21  g08897(.A0(new_n9899_), .A1(new_n9887_), .B0(new_n9862_), .Y(new_n9900_));
  OAI21  g08898(.A0(new_n9898_), .A1(new_n9889_), .B0(new_n9886_), .Y(new_n9901_));
  NAND4  g08899(.A(new_n9843_), .B(new_n9876_), .C(new_n9875_), .D(new_n9877_), .Y(new_n9902_));
  OAI21  g08900(.A0(new_n9875_), .A1(new_n9867_), .B0(new_n9885_), .Y(new_n9903_));
  OAI21  g08901(.A0(new_n9903_), .A1(new_n9902_), .B0(new_n9901_), .Y(new_n9904_));
  XOR2   g08902(.A(new_n9662_), .B(new_n9805_), .Y(new_n9905_));
  XOR2   g08903(.A(new_n9686_), .B(new_n9905_), .Y(new_n9906_));
  NAND2  g08904(.A(new_n9906_), .B(new_n9647_), .Y(new_n9907_));
  AOI211 g08905(.A0(new_n9904_), .A1(new_n9862_), .B(new_n9907_), .C(new_n9900_), .Y(new_n9908_));
  XOR2   g08906(.A(new_n9622_), .B(new_n9866_), .Y(new_n9909_));
  XOR2   g08907(.A(new_n9646_), .B(new_n9909_), .Y(new_n9910_));
  NOR2   g08908(.A(new_n9687_), .B(new_n9910_), .Y(new_n9911_));
  AOI21  g08909(.A0(new_n9904_), .A1(new_n9862_), .B0(new_n9900_), .Y(new_n9912_));
  NOR2   g08910(.A(new_n9912_), .B(new_n9911_), .Y(new_n9913_));
  OAI21  g08911(.A0(new_n9913_), .A1(new_n9908_), .B0(new_n9842_), .Y(new_n9914_));
  XOR2   g08912(.A(new_n9838_), .B(new_n9823_), .Y(new_n9915_));
  NAND2  g08913(.A(new_n9841_), .B(new_n9800_), .Y(new_n9916_));
  OAI21  g08914(.A0(new_n9915_), .A1(new_n9800_), .B0(new_n9916_), .Y(new_n9917_));
  XOR2   g08915(.A(new_n9645_), .B(new_n9643_), .Y(new_n9918_));
  NOR2   g08916(.A(new_n9645_), .B(new_n9643_), .Y(new_n9919_));
  AOI21  g08917(.A0(new_n9860_), .A1(new_n9918_), .B0(new_n9919_), .Y(new_n9920_));
  XOR2   g08918(.A(new_n9860_), .B(new_n9918_), .Y(new_n9921_));
  OAI21  g08919(.A0(new_n9920_), .A1(new_n9891_), .B0(new_n9921_), .Y(new_n9922_));
  OAI21  g08920(.A0(new_n9875_), .A1(new_n9867_), .B0(new_n9876_), .Y(new_n9923_));
  NAND2  g08921(.A(new_n9897_), .B(new_n9896_), .Y(new_n9924_));
  NOR4   g08922(.A(new_n9891_), .B(new_n9889_), .C(new_n9924_), .D(new_n9867_), .Y(new_n9925_));
  NOR2   g08923(.A(new_n9898_), .B(new_n9892_), .Y(new_n9926_));
  AOI22  g08924(.A0(new_n9926_), .A1(new_n9925_), .B0(new_n9923_), .B1(new_n9886_), .Y(new_n9927_));
  OAI21  g08925(.A0(new_n9927_), .A1(new_n9922_), .B0(new_n9907_), .Y(new_n9928_));
  OAI22  g08926(.A0(new_n9928_), .A1(new_n9900_), .B0(new_n9912_), .B1(new_n9907_), .Y(new_n9929_));
  NAND2  g08927(.A(new_n9929_), .B(new_n9917_), .Y(new_n9930_));
  NOR2   g08928(.A(new_n9769_), .B(new_n9688_), .Y(new_n9931_));
  NAND3  g08929(.A(new_n9931_), .B(new_n9930_), .C(new_n9914_), .Y(new_n9932_));
  XOR2   g08930(.A(new_n9923_), .B(new_n9886_), .Y(new_n9933_));
  NAND2  g08931(.A(new_n9933_), .B(new_n9922_), .Y(new_n9934_));
  NAND2  g08932(.A(new_n9904_), .B(new_n9862_), .Y(new_n9935_));
  NAND3  g08933(.A(new_n9911_), .B(new_n9935_), .C(new_n9934_), .Y(new_n9936_));
  NOR2   g08934(.A(new_n9927_), .B(new_n9922_), .Y(new_n9937_));
  OAI21  g08935(.A0(new_n9937_), .A1(new_n9900_), .B0(new_n9907_), .Y(new_n9938_));
  AOI21  g08936(.A0(new_n9938_), .A1(new_n9936_), .B0(new_n9917_), .Y(new_n9939_));
  NAND3  g08937(.A(new_n9907_), .B(new_n9935_), .C(new_n9934_), .Y(new_n9940_));
  OAI21  g08938(.A0(new_n9937_), .A1(new_n9900_), .B0(new_n9911_), .Y(new_n9941_));
  AOI21  g08939(.A0(new_n9941_), .A1(new_n9940_), .B0(new_n9842_), .Y(new_n9942_));
  INV    g08940(.A(new_n9931_), .Y(new_n9943_));
  OAI21  g08941(.A0(new_n9942_), .A1(new_n9939_), .B0(new_n9943_), .Y(new_n9944_));
  XOR2   g08942(.A(new_n9722_), .B(new_n9715_), .Y(new_n9945_));
  XOR2   g08943(.A(\A[287] ), .B(new_n9719_), .Y(new_n9946_));
  NAND2  g08944(.A(\A[287] ), .B(\A[286] ), .Y(new_n9947_));
  OAI21  g08945(.A0(new_n9946_), .A1(new_n9716_), .B0(new_n9947_), .Y(new_n9948_));
  XOR2   g08946(.A(new_n9726_), .B(new_n9948_), .Y(new_n9949_));
  NOR2   g08947(.A(\A[284] ), .B(new_n9712_), .Y(new_n9950_));
  OAI21  g08948(.A0(new_n9710_), .A1(\A[283] ), .B0(\A[285] ), .Y(new_n9951_));
  XOR2   g08949(.A(\A[284] ), .B(new_n9712_), .Y(new_n9952_));
  OAI22  g08950(.A0(new_n9952_), .A1(\A[285] ), .B0(new_n9951_), .B1(new_n9950_), .Y(new_n9953_));
  NOR2   g08951(.A(\A[287] ), .B(new_n9719_), .Y(new_n9954_));
  OAI21  g08952(.A0(new_n9717_), .A1(\A[286] ), .B0(\A[288] ), .Y(new_n9955_));
  OAI22  g08953(.A0(new_n9946_), .A1(\A[288] ), .B0(new_n9955_), .B1(new_n9954_), .Y(new_n9956_));
  NAND2  g08954(.A(new_n9956_), .B(new_n9953_), .Y(new_n9957_));
  NAND2  g08955(.A(\A[284] ), .B(\A[283] ), .Y(new_n9958_));
  OAI21  g08956(.A0(new_n9952_), .A1(new_n9709_), .B0(new_n9958_), .Y(new_n9959_));
  NAND2  g08957(.A(new_n9959_), .B(new_n9948_), .Y(new_n9960_));
  OAI21  g08958(.A0(new_n9957_), .A1(new_n9949_), .B0(new_n9960_), .Y(new_n9961_));
  NOR2   g08959(.A(new_n9722_), .B(new_n9715_), .Y(new_n9962_));
  XOR2   g08960(.A(new_n9962_), .B(new_n9949_), .Y(new_n9963_));
  AOI21  g08961(.A0(new_n9961_), .A1(new_n9945_), .B0(new_n9963_), .Y(new_n9964_));
  NOR2   g08962(.A(\A[290] ), .B(new_n9693_), .Y(new_n9965_));
  OAI21  g08963(.A0(new_n9691_), .A1(\A[289] ), .B0(\A[291] ), .Y(new_n9966_));
  NAND2  g08964(.A(new_n9695_), .B(new_n9690_), .Y(new_n9967_));
  OAI21  g08965(.A0(new_n9966_), .A1(new_n9965_), .B0(new_n9967_), .Y(new_n9968_));
  XOR2   g08966(.A(new_n9703_), .B(new_n9968_), .Y(new_n9969_));
  XOR2   g08967(.A(new_n9707_), .B(new_n9705_), .Y(new_n9970_));
  NOR2   g08968(.A(new_n9703_), .B(new_n9696_), .Y(new_n9971_));
  NAND2  g08969(.A(\A[293] ), .B(\A[292] ), .Y(new_n9972_));
  NAND2  g08970(.A(new_n9702_), .B(\A[294] ), .Y(new_n9973_));
  NAND2  g08971(.A(\A[290] ), .B(\A[289] ), .Y(new_n9974_));
  NAND2  g08972(.A(new_n9695_), .B(\A[291] ), .Y(new_n9975_));
  AOI22  g08973(.A0(new_n9975_), .A1(new_n9974_), .B0(new_n9973_), .B1(new_n9972_), .Y(new_n9976_));
  AOI21  g08974(.A0(new_n9971_), .A1(new_n9970_), .B0(new_n9976_), .Y(new_n9977_));
  XOR2   g08975(.A(new_n9971_), .B(new_n9970_), .Y(new_n9978_));
  XOR2   g08976(.A(new_n9703_), .B(new_n9696_), .Y(new_n9979_));
  NOR2   g08977(.A(\A[293] ), .B(new_n9700_), .Y(new_n9980_));
  OAI21  g08978(.A0(new_n9698_), .A1(\A[292] ), .B0(\A[294] ), .Y(new_n9981_));
  NAND2  g08979(.A(new_n9702_), .B(new_n9697_), .Y(new_n9982_));
  OAI21  g08980(.A0(new_n9981_), .A1(new_n9980_), .B0(new_n9982_), .Y(new_n9983_));
  NAND2  g08981(.A(new_n9973_), .B(new_n9972_), .Y(new_n9984_));
  NAND2  g08982(.A(new_n9975_), .B(new_n9974_), .Y(new_n9985_));
  NAND4  g08983(.A(new_n9985_), .B(new_n9984_), .C(new_n9983_), .D(new_n9968_), .Y(new_n9986_));
  NAND4  g08984(.A(new_n9959_), .B(new_n9948_), .C(new_n9956_), .D(new_n9953_), .Y(new_n9987_));
  NAND4  g08985(.A(new_n9987_), .B(new_n9945_), .C(new_n9986_), .D(new_n9979_), .Y(new_n9988_));
  OAI211 g08986(.A0(new_n9977_), .A1(new_n9969_), .B0(new_n9988_), .B1(new_n9978_), .Y(new_n9989_));
  XOR2   g08987(.A(new_n9707_), .B(new_n9984_), .Y(new_n9990_));
  XOR2   g08988(.A(new_n9971_), .B(new_n9990_), .Y(new_n9991_));
  NOR4   g08989(.A(new_n9707_), .B(new_n9705_), .C(new_n9703_), .D(new_n9696_), .Y(new_n9992_));
  XOR2   g08990(.A(new_n9722_), .B(new_n9953_), .Y(new_n9993_));
  NOR4   g08991(.A(new_n9726_), .B(new_n9724_), .C(new_n9722_), .D(new_n9715_), .Y(new_n9994_));
  NOR4   g08992(.A(new_n9994_), .B(new_n9993_), .C(new_n9992_), .D(new_n9969_), .Y(new_n9995_));
  AOI221 g08993(.A0(new_n9973_), .A1(new_n9972_), .C0(new_n9706_), .B0(new_n9695_), .B1(\A[291] ), .Y(new_n9996_));
  AOI221 g08994(.A0(new_n9975_), .A1(new_n9974_), .C0(new_n9704_), .B0(new_n9702_), .B1(\A[294] ), .Y(new_n9997_));
  OAI211 g08995(.A0(new_n9997_), .A1(new_n9996_), .B0(new_n9983_), .B1(new_n9968_), .Y(new_n9998_));
  NAND2  g08996(.A(new_n9985_), .B(new_n9984_), .Y(new_n9999_));
  AOI21  g08997(.A0(new_n9999_), .A1(new_n9998_), .B0(new_n9969_), .Y(new_n10000_));
  OAI21  g08998(.A0(new_n10000_), .A1(new_n9991_), .B0(new_n9995_), .Y(new_n10001_));
  AOI21  g08999(.A0(new_n10001_), .A1(new_n9989_), .B0(new_n9964_), .Y(new_n10002_));
  OAI21  g09000(.A0(new_n10000_), .A1(new_n9991_), .B0(new_n9988_), .Y(new_n10003_));
  NAND4  g09001(.A(new_n9945_), .B(new_n9978_), .C(new_n9977_), .D(new_n9979_), .Y(new_n10004_));
  OAI21  g09002(.A0(new_n9977_), .A1(new_n9969_), .B0(new_n9987_), .Y(new_n10005_));
  OAI21  g09003(.A0(new_n10005_), .A1(new_n10004_), .B0(new_n10003_), .Y(new_n10006_));
  NAND2  g09004(.A(new_n9731_), .B(\A[277] ), .Y(new_n10007_));
  AOI21  g09005(.A0(\A[278] ), .A1(new_n9729_), .B0(new_n9733_), .Y(new_n10008_));
  AOI22  g09006(.A0(new_n9734_), .A1(new_n9733_), .B0(new_n10008_), .B1(new_n10007_), .Y(new_n10009_));
  XOR2   g09007(.A(new_n9743_), .B(new_n10009_), .Y(new_n10010_));
  XOR2   g09008(.A(new_n9767_), .B(new_n10010_), .Y(new_n10011_));
  NAND2  g09009(.A(new_n10011_), .B(new_n9728_), .Y(new_n10012_));
  AOI211 g09010(.A0(new_n10006_), .A1(new_n9964_), .B(new_n10012_), .C(new_n10002_), .Y(new_n10013_));
  XOR2   g09011(.A(new_n9703_), .B(new_n9968_), .Y(new_n10014_));
  XOR2   g09012(.A(new_n9727_), .B(new_n10014_), .Y(new_n10015_));
  NOR2   g09013(.A(new_n9768_), .B(new_n10015_), .Y(new_n10016_));
  AOI21  g09014(.A0(new_n10006_), .A1(new_n9964_), .B0(new_n10002_), .Y(new_n10017_));
  NOR2   g09015(.A(new_n10017_), .B(new_n10016_), .Y(new_n10018_));
  XOR2   g09016(.A(new_n9762_), .B(new_n9755_), .Y(new_n10019_));
  XOR2   g09017(.A(\A[275] ), .B(new_n9759_), .Y(new_n10020_));
  NAND2  g09018(.A(\A[275] ), .B(\A[274] ), .Y(new_n10021_));
  OAI21  g09019(.A0(new_n10020_), .A1(new_n9756_), .B0(new_n10021_), .Y(new_n10022_));
  XOR2   g09020(.A(new_n9766_), .B(new_n10022_), .Y(new_n10023_));
  NOR2   g09021(.A(\A[272] ), .B(new_n9752_), .Y(new_n10024_));
  OAI21  g09022(.A0(new_n9750_), .A1(\A[271] ), .B0(\A[273] ), .Y(new_n10025_));
  XOR2   g09023(.A(\A[272] ), .B(new_n9752_), .Y(new_n10026_));
  OAI22  g09024(.A0(new_n10026_), .A1(\A[273] ), .B0(new_n10025_), .B1(new_n10024_), .Y(new_n10027_));
  NOR2   g09025(.A(\A[275] ), .B(new_n9759_), .Y(new_n10028_));
  OAI21  g09026(.A0(new_n9757_), .A1(\A[274] ), .B0(\A[276] ), .Y(new_n10029_));
  OAI22  g09027(.A0(new_n10020_), .A1(\A[276] ), .B0(new_n10029_), .B1(new_n10028_), .Y(new_n10030_));
  NAND2  g09028(.A(new_n10030_), .B(new_n10027_), .Y(new_n10031_));
  NAND2  g09029(.A(\A[272] ), .B(\A[271] ), .Y(new_n10032_));
  OAI21  g09030(.A0(new_n10026_), .A1(new_n9749_), .B0(new_n10032_), .Y(new_n10033_));
  NAND2  g09031(.A(new_n10033_), .B(new_n10022_), .Y(new_n10034_));
  OAI21  g09032(.A0(new_n10031_), .A1(new_n10023_), .B0(new_n10034_), .Y(new_n10035_));
  NOR2   g09033(.A(new_n9762_), .B(new_n9755_), .Y(new_n10036_));
  XOR2   g09034(.A(new_n10036_), .B(new_n10023_), .Y(new_n10037_));
  AOI21  g09035(.A0(new_n10035_), .A1(new_n10019_), .B0(new_n10037_), .Y(new_n10038_));
  XOR2   g09036(.A(new_n9743_), .B(new_n9736_), .Y(new_n10039_));
  XOR2   g09037(.A(new_n9747_), .B(new_n9745_), .Y(new_n10040_));
  NOR2   g09038(.A(new_n9743_), .B(new_n10009_), .Y(new_n10041_));
  NAND2  g09039(.A(\A[281] ), .B(\A[280] ), .Y(new_n10042_));
  NAND2  g09040(.A(new_n9742_), .B(\A[282] ), .Y(new_n10043_));
  NAND2  g09041(.A(\A[278] ), .B(\A[277] ), .Y(new_n10044_));
  NAND2  g09042(.A(new_n9734_), .B(\A[279] ), .Y(new_n10045_));
  AOI22  g09043(.A0(new_n10045_), .A1(new_n10044_), .B0(new_n10043_), .B1(new_n10042_), .Y(new_n10046_));
  AOI21  g09044(.A0(new_n10041_), .A1(new_n10040_), .B0(new_n10046_), .Y(new_n10047_));
  XOR2   g09045(.A(new_n10041_), .B(new_n10040_), .Y(new_n10048_));
  XOR2   g09046(.A(new_n9743_), .B(new_n10009_), .Y(new_n10049_));
  NOR2   g09047(.A(\A[281] ), .B(new_n9740_), .Y(new_n10050_));
  OAI21  g09048(.A0(new_n9738_), .A1(\A[280] ), .B0(\A[282] ), .Y(new_n10051_));
  NAND2  g09049(.A(new_n9742_), .B(new_n9737_), .Y(new_n10052_));
  OAI21  g09050(.A0(new_n10051_), .A1(new_n10050_), .B0(new_n10052_), .Y(new_n10053_));
  NAND2  g09051(.A(new_n10043_), .B(new_n10042_), .Y(new_n10054_));
  NAND2  g09052(.A(new_n10045_), .B(new_n10044_), .Y(new_n10055_));
  NAND4  g09053(.A(new_n10055_), .B(new_n10054_), .C(new_n10053_), .D(new_n9736_), .Y(new_n10056_));
  NAND4  g09054(.A(new_n10033_), .B(new_n10022_), .C(new_n10030_), .D(new_n10027_), .Y(new_n10057_));
  NAND4  g09055(.A(new_n10057_), .B(new_n10019_), .C(new_n10056_), .D(new_n10049_), .Y(new_n10058_));
  OAI211 g09056(.A0(new_n10047_), .A1(new_n10039_), .B0(new_n10058_), .B1(new_n10048_), .Y(new_n10059_));
  XOR2   g09057(.A(new_n9747_), .B(new_n10054_), .Y(new_n10060_));
  XOR2   g09058(.A(new_n10041_), .B(new_n10060_), .Y(new_n10061_));
  NOR4   g09059(.A(new_n9747_), .B(new_n9745_), .C(new_n9743_), .D(new_n10009_), .Y(new_n10062_));
  XOR2   g09060(.A(new_n9762_), .B(new_n10027_), .Y(new_n10063_));
  NOR4   g09061(.A(new_n9766_), .B(new_n9764_), .C(new_n9762_), .D(new_n9755_), .Y(new_n10064_));
  NOR4   g09062(.A(new_n10064_), .B(new_n10063_), .C(new_n10062_), .D(new_n10039_), .Y(new_n10065_));
  AOI221 g09063(.A0(new_n10043_), .A1(new_n10042_), .C0(new_n9746_), .B0(new_n9734_), .B1(\A[279] ), .Y(new_n10066_));
  AOI221 g09064(.A0(new_n10045_), .A1(new_n10044_), .C0(new_n9744_), .B0(new_n9742_), .B1(\A[282] ), .Y(new_n10067_));
  OAI211 g09065(.A0(new_n10067_), .A1(new_n10066_), .B0(new_n10053_), .B1(new_n9736_), .Y(new_n10068_));
  NAND2  g09066(.A(new_n10055_), .B(new_n10054_), .Y(new_n10069_));
  AOI21  g09067(.A0(new_n10069_), .A1(new_n10068_), .B0(new_n10039_), .Y(new_n10070_));
  OAI21  g09068(.A0(new_n10070_), .A1(new_n10061_), .B0(new_n10065_), .Y(new_n10071_));
  AOI21  g09069(.A0(new_n10071_), .A1(new_n10059_), .B0(new_n10038_), .Y(new_n10072_));
  NOR2   g09070(.A(new_n10070_), .B(new_n10061_), .Y(new_n10073_));
  NAND4  g09071(.A(new_n10019_), .B(new_n10048_), .C(new_n10047_), .D(new_n10049_), .Y(new_n10074_));
  OAI21  g09072(.A0(new_n10047_), .A1(new_n10039_), .B0(new_n10057_), .Y(new_n10075_));
  OAI22  g09073(.A0(new_n10075_), .A1(new_n10074_), .B0(new_n10073_), .B1(new_n10065_), .Y(new_n10076_));
  AOI21  g09074(.A0(new_n10076_), .A1(new_n10038_), .B0(new_n10072_), .Y(new_n10077_));
  OAI21  g09075(.A0(new_n10018_), .A1(new_n10013_), .B0(new_n10077_), .Y(new_n10078_));
  XOR2   g09076(.A(new_n10073_), .B(new_n10058_), .Y(new_n10079_));
  NAND2  g09077(.A(new_n10076_), .B(new_n10038_), .Y(new_n10080_));
  OAI21  g09078(.A0(new_n10079_), .A1(new_n10038_), .B0(new_n10080_), .Y(new_n10081_));
  AOI211 g09079(.A0(new_n10006_), .A1(new_n9964_), .B(new_n10016_), .C(new_n10002_), .Y(new_n10082_));
  NOR2   g09080(.A(new_n10017_), .B(new_n10012_), .Y(new_n10083_));
  OAI21  g09081(.A0(new_n10083_), .A1(new_n10082_), .B0(new_n10081_), .Y(new_n10084_));
  NAND2  g09082(.A(new_n10084_), .B(new_n10078_), .Y(new_n10085_));
  AOI21  g09083(.A0(new_n9944_), .A1(new_n9932_), .B0(new_n10085_), .Y(new_n10086_));
  XOR2   g09084(.A(new_n9726_), .B(new_n9724_), .Y(new_n10087_));
  NOR2   g09085(.A(new_n9726_), .B(new_n9724_), .Y(new_n10088_));
  AOI21  g09086(.A0(new_n9962_), .A1(new_n10087_), .B0(new_n10088_), .Y(new_n10089_));
  XOR2   g09087(.A(new_n9962_), .B(new_n10087_), .Y(new_n10090_));
  OAI21  g09088(.A0(new_n10089_), .A1(new_n9993_), .B0(new_n10090_), .Y(new_n10091_));
  OAI21  g09089(.A0(new_n9977_), .A1(new_n9969_), .B0(new_n9978_), .Y(new_n10092_));
  XOR2   g09090(.A(new_n10092_), .B(new_n9988_), .Y(new_n10093_));
  NAND2  g09091(.A(new_n10093_), .B(new_n10091_), .Y(new_n10094_));
  NAND2  g09092(.A(new_n10006_), .B(new_n9964_), .Y(new_n10095_));
  NAND3  g09093(.A(new_n10016_), .B(new_n10095_), .C(new_n10094_), .Y(new_n10096_));
  NAND2  g09094(.A(new_n9999_), .B(new_n9998_), .Y(new_n10097_));
  NOR4   g09095(.A(new_n9993_), .B(new_n9991_), .C(new_n10097_), .D(new_n9969_), .Y(new_n10098_));
  OAI211 g09096(.A0(new_n9977_), .A1(new_n9969_), .B0(new_n10098_), .B1(new_n9987_), .Y(new_n10099_));
  AOI21  g09097(.A0(new_n10099_), .A1(new_n10003_), .B0(new_n10091_), .Y(new_n10100_));
  OAI21  g09098(.A0(new_n10100_), .A1(new_n10002_), .B0(new_n10012_), .Y(new_n10101_));
  AOI21  g09099(.A0(new_n10101_), .A1(new_n10096_), .B0(new_n10081_), .Y(new_n10102_));
  NAND3  g09100(.A(new_n10012_), .B(new_n10095_), .C(new_n10094_), .Y(new_n10103_));
  OAI21  g09101(.A0(new_n10017_), .A1(new_n10012_), .B0(new_n10103_), .Y(new_n10104_));
  AOI21  g09102(.A0(new_n10104_), .A1(new_n10081_), .B0(new_n10102_), .Y(new_n10105_));
  AOI21  g09103(.A0(new_n9929_), .A1(new_n9917_), .B0(new_n9931_), .Y(new_n10106_));
  NAND2  g09104(.A(new_n10106_), .B(new_n9914_), .Y(new_n10107_));
  OAI21  g09105(.A0(new_n9942_), .A1(new_n9939_), .B0(new_n9931_), .Y(new_n10108_));
  AOI21  g09106(.A0(new_n10108_), .A1(new_n10107_), .B0(new_n10105_), .Y(new_n10109_));
  NOR2   g09107(.A(new_n10109_), .B(new_n10086_), .Y(new_n10110_));
  OAI21  g09108(.A0(new_n9780_), .A1(new_n9773_), .B0(new_n10110_), .Y(new_n10111_));
  NOR3   g09109(.A(new_n9943_), .B(new_n9942_), .C(new_n9939_), .Y(new_n10112_));
  AOI21  g09110(.A0(new_n9930_), .A1(new_n9914_), .B0(new_n9931_), .Y(new_n10113_));
  OAI21  g09111(.A0(new_n10113_), .A1(new_n10112_), .B0(new_n10105_), .Y(new_n10114_));
  NOR3   g09112(.A(new_n9931_), .B(new_n9942_), .C(new_n9939_), .Y(new_n10115_));
  AOI21  g09113(.A0(new_n9930_), .A1(new_n9914_), .B0(new_n9943_), .Y(new_n10116_));
  OAI21  g09114(.A0(new_n10116_), .A1(new_n10115_), .B0(new_n10085_), .Y(new_n10117_));
  NAND2  g09115(.A(new_n10117_), .B(new_n10114_), .Y(new_n10118_));
  NOR3   g09116(.A(new_n9771_), .B(new_n9606_), .C(new_n9598_), .Y(new_n10119_));
  AOI21  g09117(.A0(new_n9779_), .A1(new_n9776_), .B0(new_n9772_), .Y(new_n10120_));
  OAI21  g09118(.A0(new_n10120_), .A1(new_n10119_), .B0(new_n10118_), .Y(new_n10121_));
  NAND2  g09119(.A(new_n10121_), .B(new_n10111_), .Y(new_n10122_));
  INV    g09120(.A(\A[392] ), .Y(new_n10123_));
  NOR2   g09121(.A(new_n10123_), .B(\A[391] ), .Y(new_n10124_));
  INV    g09122(.A(\A[391] ), .Y(new_n10125_));
  OAI21  g09123(.A0(\A[392] ), .A1(new_n10125_), .B0(\A[393] ), .Y(new_n10126_));
  XOR2   g09124(.A(\A[392] ), .B(new_n10125_), .Y(new_n10127_));
  OAI22  g09125(.A0(new_n10127_), .A1(\A[393] ), .B0(new_n10126_), .B1(new_n10124_), .Y(new_n10128_));
  INV    g09126(.A(\A[395] ), .Y(new_n10129_));
  NOR2   g09127(.A(new_n10129_), .B(\A[394] ), .Y(new_n10130_));
  INV    g09128(.A(\A[394] ), .Y(new_n10131_));
  OAI21  g09129(.A0(\A[395] ), .A1(new_n10131_), .B0(\A[396] ), .Y(new_n10132_));
  XOR2   g09130(.A(\A[395] ), .B(new_n10131_), .Y(new_n10133_));
  OAI22  g09131(.A0(new_n10133_), .A1(\A[396] ), .B0(new_n10132_), .B1(new_n10130_), .Y(new_n10134_));
  NAND2  g09132(.A(new_n10134_), .B(new_n10128_), .Y(new_n10135_));
  INV    g09133(.A(\A[396] ), .Y(new_n10136_));
  NAND2  g09134(.A(\A[395] ), .B(\A[394] ), .Y(new_n10137_));
  OAI21  g09135(.A0(new_n10133_), .A1(new_n10136_), .B0(new_n10137_), .Y(new_n10138_));
  XOR2   g09136(.A(\A[392] ), .B(\A[391] ), .Y(new_n10139_));
  NOR2   g09137(.A(new_n10123_), .B(new_n10125_), .Y(new_n10140_));
  AOI21  g09138(.A0(new_n10139_), .A1(\A[393] ), .B0(new_n10140_), .Y(new_n10141_));
  XOR2   g09139(.A(new_n10141_), .B(new_n10138_), .Y(new_n10142_));
  XOR2   g09140(.A(new_n10142_), .B(new_n10135_), .Y(new_n10143_));
  NAND2  g09141(.A(\A[395] ), .B(new_n10131_), .Y(new_n10144_));
  AOI21  g09142(.A0(new_n10129_), .A1(\A[394] ), .B0(new_n10136_), .Y(new_n10145_));
  XOR2   g09143(.A(\A[395] ), .B(\A[394] ), .Y(new_n10146_));
  AOI22  g09144(.A0(new_n10146_), .A1(new_n10136_), .B0(new_n10145_), .B1(new_n10144_), .Y(new_n10147_));
  XOR2   g09145(.A(new_n10147_), .B(new_n10128_), .Y(new_n10148_));
  INV    g09146(.A(\A[393] ), .Y(new_n10149_));
  NAND2  g09147(.A(\A[392] ), .B(new_n10125_), .Y(new_n10150_));
  AOI21  g09148(.A0(new_n10123_), .A1(\A[391] ), .B0(new_n10149_), .Y(new_n10151_));
  AOI22  g09149(.A0(new_n10139_), .A1(new_n10149_), .B0(new_n10151_), .B1(new_n10150_), .Y(new_n10152_));
  NOR2   g09150(.A(new_n10147_), .B(new_n10152_), .Y(new_n10153_));
  NOR2   g09151(.A(new_n10129_), .B(new_n10131_), .Y(new_n10154_));
  AOI21  g09152(.A0(new_n10146_), .A1(\A[396] ), .B0(new_n10154_), .Y(new_n10155_));
  XOR2   g09153(.A(new_n10141_), .B(new_n10155_), .Y(new_n10156_));
  NOR2   g09154(.A(new_n10141_), .B(new_n10155_), .Y(new_n10157_));
  AOI21  g09155(.A0(new_n10156_), .A1(new_n10153_), .B0(new_n10157_), .Y(new_n10158_));
  OAI21  g09156(.A0(new_n10158_), .A1(new_n10148_), .B0(new_n10143_), .Y(new_n10159_));
  XOR2   g09157(.A(new_n10147_), .B(new_n10152_), .Y(new_n10160_));
  NAND2  g09158(.A(\A[401] ), .B(\A[400] ), .Y(new_n10161_));
  XOR2   g09159(.A(\A[401] ), .B(\A[400] ), .Y(new_n10162_));
  NAND2  g09160(.A(new_n10162_), .B(\A[402] ), .Y(new_n10163_));
  NAND2  g09161(.A(new_n10163_), .B(new_n10161_), .Y(new_n10164_));
  NAND2  g09162(.A(\A[398] ), .B(\A[397] ), .Y(new_n10165_));
  XOR2   g09163(.A(\A[398] ), .B(\A[397] ), .Y(new_n10166_));
  NAND2  g09164(.A(new_n10166_), .B(\A[399] ), .Y(new_n10167_));
  NAND2  g09165(.A(new_n10167_), .B(new_n10165_), .Y(new_n10168_));
  INV    g09166(.A(\A[398] ), .Y(new_n10169_));
  NOR2   g09167(.A(new_n10169_), .B(\A[397] ), .Y(new_n10170_));
  INV    g09168(.A(\A[397] ), .Y(new_n10171_));
  OAI21  g09169(.A0(\A[398] ), .A1(new_n10171_), .B0(\A[399] ), .Y(new_n10172_));
  INV    g09170(.A(\A[399] ), .Y(new_n10173_));
  NAND2  g09171(.A(new_n10166_), .B(new_n10173_), .Y(new_n10174_));
  OAI21  g09172(.A0(new_n10172_), .A1(new_n10170_), .B0(new_n10174_), .Y(new_n10175_));
  INV    g09173(.A(\A[401] ), .Y(new_n10176_));
  NOR2   g09174(.A(new_n10176_), .B(\A[400] ), .Y(new_n10177_));
  INV    g09175(.A(\A[400] ), .Y(new_n10178_));
  OAI21  g09176(.A0(\A[401] ), .A1(new_n10178_), .B0(\A[402] ), .Y(new_n10179_));
  INV    g09177(.A(\A[402] ), .Y(new_n10180_));
  NAND2  g09178(.A(new_n10162_), .B(new_n10180_), .Y(new_n10181_));
  OAI21  g09179(.A0(new_n10179_), .A1(new_n10177_), .B0(new_n10181_), .Y(new_n10182_));
  NAND4  g09180(.A(new_n10182_), .B(new_n10175_), .C(new_n10168_), .D(new_n10164_), .Y(new_n10183_));
  NAND2  g09181(.A(\A[392] ), .B(\A[391] ), .Y(new_n10184_));
  OAI21  g09182(.A0(new_n10127_), .A1(new_n10149_), .B0(new_n10184_), .Y(new_n10185_));
  NAND4  g09183(.A(new_n10185_), .B(new_n10138_), .C(new_n10134_), .D(new_n10128_), .Y(new_n10186_));
  NAND2  g09184(.A(\A[398] ), .B(new_n10171_), .Y(new_n10187_));
  AOI21  g09185(.A0(new_n10169_), .A1(\A[397] ), .B0(new_n10173_), .Y(new_n10188_));
  AOI22  g09186(.A0(new_n10188_), .A1(new_n10187_), .B0(new_n10166_), .B1(new_n10173_), .Y(new_n10189_));
  NAND2  g09187(.A(\A[401] ), .B(new_n10178_), .Y(new_n10190_));
  AOI21  g09188(.A0(new_n10176_), .A1(\A[400] ), .B0(new_n10180_), .Y(new_n10191_));
  AOI22  g09189(.A0(new_n10191_), .A1(new_n10190_), .B0(new_n10162_), .B1(new_n10180_), .Y(new_n10192_));
  XOR2   g09190(.A(new_n10192_), .B(new_n10189_), .Y(new_n10193_));
  NAND4  g09191(.A(new_n10193_), .B(new_n10186_), .C(new_n10183_), .D(new_n10160_), .Y(new_n10194_));
  XOR2   g09192(.A(new_n10168_), .B(new_n10164_), .Y(new_n10195_));
  NOR2   g09193(.A(new_n10192_), .B(new_n10189_), .Y(new_n10196_));
  AOI22  g09194(.A0(new_n10167_), .A1(new_n10165_), .B0(new_n10163_), .B1(new_n10161_), .Y(new_n10197_));
  AOI21  g09195(.A0(new_n10196_), .A1(new_n10195_), .B0(new_n10197_), .Y(new_n10198_));
  XOR2   g09196(.A(new_n10196_), .B(new_n10195_), .Y(new_n10199_));
  XOR2   g09197(.A(new_n10192_), .B(new_n10175_), .Y(new_n10200_));
  OAI21  g09198(.A0(new_n10200_), .A1(new_n10198_), .B0(new_n10199_), .Y(new_n10201_));
  XOR2   g09199(.A(new_n10201_), .B(new_n10194_), .Y(new_n10202_));
  NAND2  g09200(.A(new_n10182_), .B(new_n10175_), .Y(new_n10203_));
  XOR2   g09201(.A(new_n10203_), .B(new_n10195_), .Y(new_n10204_));
  NOR2   g09202(.A(new_n10169_), .B(new_n10171_), .Y(new_n10205_));
  AOI221 g09203(.A0(new_n10166_), .A1(\A[399] ), .C0(new_n10205_), .B0(new_n10163_), .B1(new_n10161_), .Y(new_n10206_));
  NOR2   g09204(.A(new_n10176_), .B(new_n10178_), .Y(new_n10207_));
  AOI221 g09205(.A0(new_n10167_), .A1(new_n10165_), .C0(new_n10207_), .B0(new_n10162_), .B1(\A[402] ), .Y(new_n10208_));
  OAI211 g09206(.A0(new_n10208_), .A1(new_n10206_), .B0(new_n10182_), .B1(new_n10175_), .Y(new_n10209_));
  NAND2  g09207(.A(new_n10168_), .B(new_n10164_), .Y(new_n10210_));
  AOI21  g09208(.A0(new_n10210_), .A1(new_n10209_), .B0(new_n10200_), .Y(new_n10211_));
  OAI21  g09209(.A0(new_n10211_), .A1(new_n10204_), .B0(new_n10194_), .Y(new_n10212_));
  NOR2   g09210(.A(new_n10200_), .B(new_n10148_), .Y(new_n10213_));
  OAI211 g09211(.A0(new_n10182_), .A1(new_n10175_), .B0(new_n10168_), .B1(new_n10164_), .Y(new_n10214_));
  NAND4  g09212(.A(new_n10214_), .B(new_n10213_), .C(new_n10186_), .D(new_n10199_), .Y(new_n10215_));
  AOI21  g09213(.A0(new_n10215_), .A1(new_n10212_), .B0(new_n10159_), .Y(new_n10216_));
  AOI21  g09214(.A0(new_n10202_), .A1(new_n10159_), .B0(new_n10216_), .Y(new_n10217_));
  INV    g09215(.A(\A[405] ), .Y(new_n10218_));
  INV    g09216(.A(\A[403] ), .Y(new_n10219_));
  NAND2  g09217(.A(\A[404] ), .B(new_n10219_), .Y(new_n10220_));
  INV    g09218(.A(\A[404] ), .Y(new_n10221_));
  AOI21  g09219(.A0(new_n10221_), .A1(\A[403] ), .B0(new_n10218_), .Y(new_n10222_));
  XOR2   g09220(.A(\A[404] ), .B(\A[403] ), .Y(new_n10223_));
  AOI22  g09221(.A0(new_n10223_), .A1(new_n10218_), .B0(new_n10222_), .B1(new_n10220_), .Y(new_n10224_));
  INV    g09222(.A(\A[408] ), .Y(new_n10225_));
  INV    g09223(.A(\A[406] ), .Y(new_n10226_));
  NAND2  g09224(.A(\A[407] ), .B(new_n10226_), .Y(new_n10227_));
  INV    g09225(.A(\A[407] ), .Y(new_n10228_));
  AOI21  g09226(.A0(new_n10228_), .A1(\A[406] ), .B0(new_n10225_), .Y(new_n10229_));
  XOR2   g09227(.A(\A[407] ), .B(\A[406] ), .Y(new_n10230_));
  AOI22  g09228(.A0(new_n10230_), .A1(new_n10225_), .B0(new_n10229_), .B1(new_n10227_), .Y(new_n10231_));
  NOR2   g09229(.A(new_n10231_), .B(new_n10224_), .Y(new_n10232_));
  XOR2   g09230(.A(\A[407] ), .B(new_n10226_), .Y(new_n10233_));
  NAND2  g09231(.A(\A[407] ), .B(\A[406] ), .Y(new_n10234_));
  OAI21  g09232(.A0(new_n10233_), .A1(new_n10225_), .B0(new_n10234_), .Y(new_n10235_));
  NOR2   g09233(.A(new_n10221_), .B(new_n10219_), .Y(new_n10236_));
  AOI21  g09234(.A0(new_n10223_), .A1(\A[405] ), .B0(new_n10236_), .Y(new_n10237_));
  XOR2   g09235(.A(new_n10237_), .B(new_n10235_), .Y(new_n10238_));
  XOR2   g09236(.A(new_n10238_), .B(new_n10232_), .Y(new_n10239_));
  XOR2   g09237(.A(new_n10231_), .B(new_n10224_), .Y(new_n10240_));
  NOR2   g09238(.A(new_n10221_), .B(\A[403] ), .Y(new_n10241_));
  OAI21  g09239(.A0(\A[404] ), .A1(new_n10219_), .B0(\A[405] ), .Y(new_n10242_));
  XOR2   g09240(.A(\A[404] ), .B(new_n10219_), .Y(new_n10243_));
  OAI22  g09241(.A0(new_n10243_), .A1(\A[405] ), .B0(new_n10242_), .B1(new_n10241_), .Y(new_n10244_));
  NOR2   g09242(.A(new_n10228_), .B(\A[406] ), .Y(new_n10245_));
  OAI21  g09243(.A0(\A[407] ), .A1(new_n10226_), .B0(\A[408] ), .Y(new_n10246_));
  OAI22  g09244(.A0(new_n10233_), .A1(\A[408] ), .B0(new_n10246_), .B1(new_n10245_), .Y(new_n10247_));
  NAND2  g09245(.A(new_n10247_), .B(new_n10244_), .Y(new_n10248_));
  NAND2  g09246(.A(\A[404] ), .B(\A[403] ), .Y(new_n10249_));
  OAI21  g09247(.A0(new_n10243_), .A1(new_n10218_), .B0(new_n10249_), .Y(new_n10250_));
  NAND2  g09248(.A(new_n10250_), .B(new_n10235_), .Y(new_n10251_));
  OAI21  g09249(.A0(new_n10238_), .A1(new_n10248_), .B0(new_n10251_), .Y(new_n10252_));
  AOI21  g09250(.A0(new_n10252_), .A1(new_n10240_), .B0(new_n10239_), .Y(new_n10253_));
  NAND2  g09251(.A(\A[413] ), .B(\A[412] ), .Y(new_n10254_));
  XOR2   g09252(.A(\A[413] ), .B(\A[412] ), .Y(new_n10255_));
  NAND2  g09253(.A(new_n10255_), .B(\A[414] ), .Y(new_n10256_));
  NAND2  g09254(.A(new_n10256_), .B(new_n10254_), .Y(new_n10257_));
  NAND2  g09255(.A(\A[410] ), .B(\A[409] ), .Y(new_n10258_));
  XOR2   g09256(.A(\A[410] ), .B(\A[409] ), .Y(new_n10259_));
  NAND2  g09257(.A(new_n10259_), .B(\A[411] ), .Y(new_n10260_));
  NAND2  g09258(.A(new_n10260_), .B(new_n10258_), .Y(new_n10261_));
  XOR2   g09259(.A(new_n10261_), .B(new_n10257_), .Y(new_n10262_));
  INV    g09260(.A(\A[411] ), .Y(new_n10263_));
  INV    g09261(.A(\A[409] ), .Y(new_n10264_));
  NAND2  g09262(.A(\A[410] ), .B(new_n10264_), .Y(new_n10265_));
  INV    g09263(.A(\A[410] ), .Y(new_n10266_));
  AOI21  g09264(.A0(new_n10266_), .A1(\A[409] ), .B0(new_n10263_), .Y(new_n10267_));
  AOI22  g09265(.A0(new_n10267_), .A1(new_n10265_), .B0(new_n10259_), .B1(new_n10263_), .Y(new_n10268_));
  INV    g09266(.A(\A[414] ), .Y(new_n10269_));
  INV    g09267(.A(\A[412] ), .Y(new_n10270_));
  NAND2  g09268(.A(\A[413] ), .B(new_n10270_), .Y(new_n10271_));
  INV    g09269(.A(\A[413] ), .Y(new_n10272_));
  AOI21  g09270(.A0(new_n10272_), .A1(\A[412] ), .B0(new_n10269_), .Y(new_n10273_));
  AOI22  g09271(.A0(new_n10273_), .A1(new_n10271_), .B0(new_n10255_), .B1(new_n10269_), .Y(new_n10274_));
  NOR2   g09272(.A(new_n10274_), .B(new_n10268_), .Y(new_n10275_));
  AOI22  g09273(.A0(new_n10260_), .A1(new_n10258_), .B0(new_n10256_), .B1(new_n10254_), .Y(new_n10276_));
  AOI21  g09274(.A0(new_n10275_), .A1(new_n10262_), .B0(new_n10276_), .Y(new_n10277_));
  XOR2   g09275(.A(new_n10275_), .B(new_n10262_), .Y(new_n10278_));
  NOR2   g09276(.A(new_n10266_), .B(\A[409] ), .Y(new_n10279_));
  OAI21  g09277(.A0(\A[410] ), .A1(new_n10264_), .B0(\A[411] ), .Y(new_n10280_));
  NAND2  g09278(.A(new_n10259_), .B(new_n10263_), .Y(new_n10281_));
  OAI21  g09279(.A0(new_n10280_), .A1(new_n10279_), .B0(new_n10281_), .Y(new_n10282_));
  XOR2   g09280(.A(new_n10274_), .B(new_n10282_), .Y(new_n10283_));
  NOR2   g09281(.A(new_n10272_), .B(\A[412] ), .Y(new_n10284_));
  OAI21  g09282(.A0(\A[413] ), .A1(new_n10270_), .B0(\A[414] ), .Y(new_n10285_));
  NAND2  g09283(.A(new_n10255_), .B(new_n10269_), .Y(new_n10286_));
  OAI21  g09284(.A0(new_n10285_), .A1(new_n10284_), .B0(new_n10286_), .Y(new_n10287_));
  NAND4  g09285(.A(new_n10287_), .B(new_n10282_), .C(new_n10261_), .D(new_n10257_), .Y(new_n10288_));
  NAND4  g09286(.A(new_n10250_), .B(new_n10235_), .C(new_n10247_), .D(new_n10244_), .Y(new_n10289_));
  XOR2   g09287(.A(new_n10274_), .B(new_n10268_), .Y(new_n10290_));
  NAND4  g09288(.A(new_n10290_), .B(new_n10289_), .C(new_n10288_), .D(new_n10240_), .Y(new_n10291_));
  OAI211 g09289(.A0(new_n10283_), .A1(new_n10277_), .B0(new_n10291_), .B1(new_n10278_), .Y(new_n10292_));
  NOR2   g09290(.A(new_n10266_), .B(new_n10264_), .Y(new_n10293_));
  AOI21  g09291(.A0(new_n10259_), .A1(\A[411] ), .B0(new_n10293_), .Y(new_n10294_));
  XOR2   g09292(.A(new_n10294_), .B(new_n10257_), .Y(new_n10295_));
  XOR2   g09293(.A(new_n10275_), .B(new_n10295_), .Y(new_n10296_));
  XOR2   g09294(.A(new_n10231_), .B(new_n10244_), .Y(new_n10297_));
  NOR2   g09295(.A(new_n10272_), .B(new_n10270_), .Y(new_n10298_));
  AOI21  g09296(.A0(new_n10255_), .A1(\A[414] ), .B0(new_n10298_), .Y(new_n10299_));
  NOR4   g09297(.A(new_n10274_), .B(new_n10268_), .C(new_n10294_), .D(new_n10299_), .Y(new_n10300_));
  NOR2   g09298(.A(new_n10228_), .B(new_n10226_), .Y(new_n10301_));
  AOI21  g09299(.A0(new_n10230_), .A1(\A[408] ), .B0(new_n10301_), .Y(new_n10302_));
  NOR4   g09300(.A(new_n10237_), .B(new_n10302_), .C(new_n10231_), .D(new_n10224_), .Y(new_n10303_));
  NOR4   g09301(.A(new_n10283_), .B(new_n10303_), .C(new_n10300_), .D(new_n10297_), .Y(new_n10304_));
  AOI221 g09302(.A0(new_n10259_), .A1(\A[411] ), .C0(new_n10293_), .B0(new_n10256_), .B1(new_n10254_), .Y(new_n10305_));
  AOI221 g09303(.A0(new_n10260_), .A1(new_n10258_), .C0(new_n10298_), .B0(new_n10255_), .B1(\A[414] ), .Y(new_n10306_));
  OAI211 g09304(.A0(new_n10306_), .A1(new_n10305_), .B0(new_n10287_), .B1(new_n10282_), .Y(new_n10307_));
  NAND2  g09305(.A(new_n10261_), .B(new_n10257_), .Y(new_n10308_));
  AOI21  g09306(.A0(new_n10308_), .A1(new_n10307_), .B0(new_n10283_), .Y(new_n10309_));
  OAI21  g09307(.A0(new_n10309_), .A1(new_n10296_), .B0(new_n10304_), .Y(new_n10310_));
  AOI21  g09308(.A0(new_n10310_), .A1(new_n10292_), .B0(new_n10253_), .Y(new_n10311_));
  XOR2   g09309(.A(new_n10238_), .B(new_n10248_), .Y(new_n10312_));
  XOR2   g09310(.A(new_n10237_), .B(new_n10302_), .Y(new_n10313_));
  NOR2   g09311(.A(new_n10237_), .B(new_n10302_), .Y(new_n10314_));
  AOI21  g09312(.A0(new_n10313_), .A1(new_n10232_), .B0(new_n10314_), .Y(new_n10315_));
  OAI21  g09313(.A0(new_n10315_), .A1(new_n10297_), .B0(new_n10312_), .Y(new_n10316_));
  OAI21  g09314(.A0(new_n10309_), .A1(new_n10296_), .B0(new_n10291_), .Y(new_n10317_));
  NOR2   g09315(.A(new_n10283_), .B(new_n10297_), .Y(new_n10318_));
  OAI211 g09316(.A0(new_n10287_), .A1(new_n10282_), .B0(new_n10261_), .B1(new_n10257_), .Y(new_n10319_));
  NAND4  g09317(.A(new_n10319_), .B(new_n10318_), .C(new_n10289_), .D(new_n10278_), .Y(new_n10320_));
  AOI21  g09318(.A0(new_n10320_), .A1(new_n10317_), .B0(new_n10316_), .Y(new_n10321_));
  NOR2   g09319(.A(new_n10283_), .B(new_n10300_), .Y(new_n10322_));
  XOR2   g09320(.A(new_n10231_), .B(new_n10224_), .Y(new_n10323_));
  XOR2   g09321(.A(new_n10323_), .B(new_n10322_), .Y(new_n10324_));
  NAND2  g09322(.A(new_n10193_), .B(new_n10183_), .Y(new_n10325_));
  XOR2   g09323(.A(new_n10147_), .B(new_n10128_), .Y(new_n10326_));
  XOR2   g09324(.A(new_n10326_), .B(new_n10325_), .Y(new_n10327_));
  NAND2  g09325(.A(new_n10327_), .B(new_n10324_), .Y(new_n10328_));
  NOR3   g09326(.A(new_n10328_), .B(new_n10321_), .C(new_n10311_), .Y(new_n10329_));
  OAI21  g09327(.A0(new_n10283_), .A1(new_n10277_), .B0(new_n10278_), .Y(new_n10330_));
  XOR2   g09328(.A(new_n10330_), .B(new_n10291_), .Y(new_n10331_));
  NAND2  g09329(.A(new_n10331_), .B(new_n10316_), .Y(new_n10332_));
  NAND2  g09330(.A(new_n10320_), .B(new_n10317_), .Y(new_n10333_));
  NAND2  g09331(.A(new_n10333_), .B(new_n10253_), .Y(new_n10334_));
  NAND2  g09332(.A(new_n10290_), .B(new_n10288_), .Y(new_n10335_));
  XOR2   g09333(.A(new_n10323_), .B(new_n10335_), .Y(new_n10336_));
  XOR2   g09334(.A(new_n10147_), .B(new_n10152_), .Y(new_n10337_));
  XOR2   g09335(.A(new_n10337_), .B(new_n10325_), .Y(new_n10338_));
  NOR2   g09336(.A(new_n10338_), .B(new_n10336_), .Y(new_n10339_));
  AOI21  g09337(.A0(new_n10334_), .A1(new_n10332_), .B0(new_n10339_), .Y(new_n10340_));
  OAI21  g09338(.A0(new_n10340_), .A1(new_n10329_), .B0(new_n10217_), .Y(new_n10341_));
  NAND2  g09339(.A(new_n10202_), .B(new_n10159_), .Y(new_n10342_));
  NAND2  g09340(.A(new_n10210_), .B(new_n10209_), .Y(new_n10343_));
  NAND3  g09341(.A(new_n10213_), .B(new_n10186_), .C(new_n10199_), .Y(new_n10344_));
  AOI211 g09342(.A0(new_n10199_), .A1(new_n10343_), .B(new_n10344_), .C(new_n10211_), .Y(new_n10345_));
  AOI21  g09343(.A0(new_n10201_), .A1(new_n10194_), .B0(new_n10345_), .Y(new_n10346_));
  OAI21  g09344(.A0(new_n10346_), .A1(new_n10159_), .B0(new_n10342_), .Y(new_n10347_));
  NAND2  g09345(.A(new_n10290_), .B(new_n10240_), .Y(new_n10348_));
  AOI211 g09346(.A0(new_n10274_), .A1(new_n10268_), .B(new_n10294_), .C(new_n10299_), .Y(new_n10349_));
  NOR4   g09347(.A(new_n10349_), .B(new_n10348_), .C(new_n10303_), .D(new_n10296_), .Y(new_n10350_));
  AOI21  g09348(.A0(new_n10330_), .A1(new_n10291_), .B0(new_n10350_), .Y(new_n10351_));
  OAI21  g09349(.A0(new_n10351_), .A1(new_n10316_), .B0(new_n10328_), .Y(new_n10352_));
  OAI21  g09350(.A0(new_n10321_), .A1(new_n10311_), .B0(new_n10339_), .Y(new_n10353_));
  OAI21  g09351(.A0(new_n10352_), .A1(new_n10311_), .B0(new_n10353_), .Y(new_n10354_));
  NAND2  g09352(.A(new_n10354_), .B(new_n10347_), .Y(new_n10355_));
  XOR2   g09353(.A(new_n10338_), .B(new_n10324_), .Y(new_n10356_));
  INV    g09354(.A(\A[387] ), .Y(new_n10357_));
  INV    g09355(.A(\A[386] ), .Y(new_n10358_));
  NAND2  g09356(.A(new_n10358_), .B(\A[385] ), .Y(new_n10359_));
  INV    g09357(.A(\A[385] ), .Y(new_n10360_));
  AOI21  g09358(.A0(\A[386] ), .A1(new_n10360_), .B0(new_n10357_), .Y(new_n10361_));
  XOR2   g09359(.A(\A[386] ), .B(\A[385] ), .Y(new_n10362_));
  AOI22  g09360(.A0(new_n10362_), .A1(new_n10357_), .B0(new_n10361_), .B1(new_n10359_), .Y(new_n10363_));
  INV    g09361(.A(\A[390] ), .Y(new_n10364_));
  INV    g09362(.A(\A[389] ), .Y(new_n10365_));
  NAND2  g09363(.A(new_n10365_), .B(\A[388] ), .Y(new_n10366_));
  INV    g09364(.A(\A[388] ), .Y(new_n10367_));
  AOI21  g09365(.A0(\A[389] ), .A1(new_n10367_), .B0(new_n10364_), .Y(new_n10368_));
  XOR2   g09366(.A(\A[389] ), .B(\A[388] ), .Y(new_n10369_));
  AOI22  g09367(.A0(new_n10369_), .A1(new_n10364_), .B0(new_n10368_), .B1(new_n10366_), .Y(new_n10370_));
  NOR2   g09368(.A(new_n10365_), .B(new_n10367_), .Y(new_n10371_));
  AOI21  g09369(.A0(new_n10369_), .A1(\A[390] ), .B0(new_n10371_), .Y(new_n10372_));
  NOR2   g09370(.A(new_n10358_), .B(new_n10360_), .Y(new_n10373_));
  AOI21  g09371(.A0(new_n10362_), .A1(\A[387] ), .B0(new_n10373_), .Y(new_n10374_));
  XOR2   g09372(.A(new_n10370_), .B(new_n10363_), .Y(new_n10375_));
  INV    g09373(.A(\A[381] ), .Y(new_n10376_));
  INV    g09374(.A(\A[380] ), .Y(new_n10377_));
  NAND2  g09375(.A(new_n10377_), .B(\A[379] ), .Y(new_n10378_));
  INV    g09376(.A(\A[379] ), .Y(new_n10379_));
  AOI21  g09377(.A0(\A[380] ), .A1(new_n10379_), .B0(new_n10376_), .Y(new_n10380_));
  XOR2   g09378(.A(\A[380] ), .B(\A[379] ), .Y(new_n10381_));
  AOI22  g09379(.A0(new_n10381_), .A1(new_n10376_), .B0(new_n10380_), .B1(new_n10378_), .Y(new_n10382_));
  INV    g09380(.A(\A[384] ), .Y(new_n10383_));
  INV    g09381(.A(\A[383] ), .Y(new_n10384_));
  NAND2  g09382(.A(new_n10384_), .B(\A[382] ), .Y(new_n10385_));
  INV    g09383(.A(\A[382] ), .Y(new_n10386_));
  AOI21  g09384(.A0(\A[383] ), .A1(new_n10386_), .B0(new_n10383_), .Y(new_n10387_));
  XOR2   g09385(.A(\A[383] ), .B(\A[382] ), .Y(new_n10388_));
  AOI22  g09386(.A0(new_n10388_), .A1(new_n10383_), .B0(new_n10387_), .B1(new_n10385_), .Y(new_n10389_));
  NOR2   g09387(.A(new_n10384_), .B(new_n10386_), .Y(new_n10390_));
  AOI21  g09388(.A0(new_n10388_), .A1(\A[384] ), .B0(new_n10390_), .Y(new_n10391_));
  NOR2   g09389(.A(new_n10377_), .B(new_n10379_), .Y(new_n10392_));
  AOI21  g09390(.A0(new_n10381_), .A1(\A[381] ), .B0(new_n10392_), .Y(new_n10393_));
  XOR2   g09391(.A(new_n10389_), .B(new_n10382_), .Y(new_n10394_));
  XOR2   g09392(.A(new_n10394_), .B(new_n10375_), .Y(new_n10395_));
  INV    g09393(.A(\A[373] ), .Y(new_n10396_));
  NOR2   g09394(.A(\A[374] ), .B(new_n10396_), .Y(new_n10397_));
  INV    g09395(.A(\A[374] ), .Y(new_n10398_));
  OAI21  g09396(.A0(new_n10398_), .A1(\A[373] ), .B0(\A[375] ), .Y(new_n10399_));
  INV    g09397(.A(\A[375] ), .Y(new_n10400_));
  XOR2   g09398(.A(\A[374] ), .B(\A[373] ), .Y(new_n10401_));
  NAND2  g09399(.A(new_n10401_), .B(new_n10400_), .Y(new_n10402_));
  OAI21  g09400(.A0(new_n10399_), .A1(new_n10397_), .B0(new_n10402_), .Y(new_n10403_));
  INV    g09401(.A(\A[378] ), .Y(new_n10404_));
  INV    g09402(.A(\A[377] ), .Y(new_n10405_));
  NAND2  g09403(.A(new_n10405_), .B(\A[376] ), .Y(new_n10406_));
  INV    g09404(.A(\A[376] ), .Y(new_n10407_));
  AOI21  g09405(.A0(\A[377] ), .A1(new_n10407_), .B0(new_n10404_), .Y(new_n10408_));
  XOR2   g09406(.A(\A[377] ), .B(\A[376] ), .Y(new_n10409_));
  AOI22  g09407(.A0(new_n10409_), .A1(new_n10404_), .B0(new_n10408_), .B1(new_n10406_), .Y(new_n10410_));
  NOR2   g09408(.A(new_n10405_), .B(new_n10407_), .Y(new_n10411_));
  AOI21  g09409(.A0(new_n10409_), .A1(\A[378] ), .B0(new_n10411_), .Y(new_n10412_));
  NOR2   g09410(.A(new_n10398_), .B(new_n10396_), .Y(new_n10413_));
  AOI21  g09411(.A0(new_n10401_), .A1(\A[375] ), .B0(new_n10413_), .Y(new_n10414_));
  XOR2   g09412(.A(new_n10410_), .B(new_n10403_), .Y(new_n10415_));
  INV    g09413(.A(\A[369] ), .Y(new_n10416_));
  INV    g09414(.A(\A[368] ), .Y(new_n10417_));
  NAND2  g09415(.A(new_n10417_), .B(\A[367] ), .Y(new_n10418_));
  INV    g09416(.A(\A[367] ), .Y(new_n10419_));
  AOI21  g09417(.A0(\A[368] ), .A1(new_n10419_), .B0(new_n10416_), .Y(new_n10420_));
  XOR2   g09418(.A(\A[368] ), .B(\A[367] ), .Y(new_n10421_));
  AOI22  g09419(.A0(new_n10421_), .A1(new_n10416_), .B0(new_n10420_), .B1(new_n10418_), .Y(new_n10422_));
  INV    g09420(.A(\A[372] ), .Y(new_n10423_));
  INV    g09421(.A(\A[371] ), .Y(new_n10424_));
  NAND2  g09422(.A(new_n10424_), .B(\A[370] ), .Y(new_n10425_));
  INV    g09423(.A(\A[370] ), .Y(new_n10426_));
  AOI21  g09424(.A0(\A[371] ), .A1(new_n10426_), .B0(new_n10423_), .Y(new_n10427_));
  XOR2   g09425(.A(\A[371] ), .B(\A[370] ), .Y(new_n10428_));
  AOI22  g09426(.A0(new_n10428_), .A1(new_n10423_), .B0(new_n10427_), .B1(new_n10425_), .Y(new_n10429_));
  NOR2   g09427(.A(new_n10424_), .B(new_n10426_), .Y(new_n10430_));
  AOI21  g09428(.A0(new_n10428_), .A1(\A[372] ), .B0(new_n10430_), .Y(new_n10431_));
  NOR2   g09429(.A(new_n10417_), .B(new_n10419_), .Y(new_n10432_));
  AOI21  g09430(.A0(new_n10421_), .A1(\A[369] ), .B0(new_n10432_), .Y(new_n10433_));
  XOR2   g09431(.A(new_n10429_), .B(new_n10422_), .Y(new_n10434_));
  XOR2   g09432(.A(new_n10434_), .B(new_n10415_), .Y(new_n10435_));
  XOR2   g09433(.A(new_n10435_), .B(new_n10395_), .Y(new_n10436_));
  NOR2   g09434(.A(new_n10436_), .B(new_n10356_), .Y(new_n10437_));
  NAND3  g09435(.A(new_n10437_), .B(new_n10355_), .C(new_n10341_), .Y(new_n10438_));
  NAND3  g09436(.A(new_n10339_), .B(new_n10334_), .C(new_n10332_), .Y(new_n10439_));
  OAI21  g09437(.A0(new_n10321_), .A1(new_n10311_), .B0(new_n10328_), .Y(new_n10440_));
  AOI21  g09438(.A0(new_n10440_), .A1(new_n10439_), .B0(new_n10347_), .Y(new_n10441_));
  NAND3  g09439(.A(new_n10328_), .B(new_n10334_), .C(new_n10332_), .Y(new_n10442_));
  AOI21  g09440(.A0(new_n10353_), .A1(new_n10442_), .B0(new_n10217_), .Y(new_n10443_));
  INV    g09441(.A(new_n10437_), .Y(new_n10444_));
  OAI21  g09442(.A0(new_n10443_), .A1(new_n10441_), .B0(new_n10444_), .Y(new_n10445_));
  XOR2   g09443(.A(new_n10389_), .B(new_n10382_), .Y(new_n10446_));
  XOR2   g09444(.A(\A[383] ), .B(new_n10386_), .Y(new_n10447_));
  NAND2  g09445(.A(\A[383] ), .B(\A[382] ), .Y(new_n10448_));
  OAI21  g09446(.A0(new_n10447_), .A1(new_n10383_), .B0(new_n10448_), .Y(new_n10449_));
  XOR2   g09447(.A(new_n10393_), .B(new_n10449_), .Y(new_n10450_));
  NOR2   g09448(.A(\A[380] ), .B(new_n10379_), .Y(new_n10451_));
  OAI21  g09449(.A0(new_n10377_), .A1(\A[379] ), .B0(\A[381] ), .Y(new_n10452_));
  XOR2   g09450(.A(\A[380] ), .B(new_n10379_), .Y(new_n10453_));
  OAI22  g09451(.A0(new_n10453_), .A1(\A[381] ), .B0(new_n10452_), .B1(new_n10451_), .Y(new_n10454_));
  NOR2   g09452(.A(\A[383] ), .B(new_n10386_), .Y(new_n10455_));
  OAI21  g09453(.A0(new_n10384_), .A1(\A[382] ), .B0(\A[384] ), .Y(new_n10456_));
  OAI22  g09454(.A0(new_n10447_), .A1(\A[384] ), .B0(new_n10456_), .B1(new_n10455_), .Y(new_n10457_));
  NAND2  g09455(.A(new_n10457_), .B(new_n10454_), .Y(new_n10458_));
  NAND2  g09456(.A(\A[380] ), .B(\A[379] ), .Y(new_n10459_));
  OAI21  g09457(.A0(new_n10453_), .A1(new_n10376_), .B0(new_n10459_), .Y(new_n10460_));
  NAND2  g09458(.A(new_n10460_), .B(new_n10449_), .Y(new_n10461_));
  OAI21  g09459(.A0(new_n10458_), .A1(new_n10450_), .B0(new_n10461_), .Y(new_n10462_));
  NOR2   g09460(.A(new_n10389_), .B(new_n10382_), .Y(new_n10463_));
  XOR2   g09461(.A(new_n10463_), .B(new_n10450_), .Y(new_n10464_));
  AOI21  g09462(.A0(new_n10462_), .A1(new_n10446_), .B0(new_n10464_), .Y(new_n10465_));
  NOR2   g09463(.A(\A[386] ), .B(new_n10360_), .Y(new_n10466_));
  OAI21  g09464(.A0(new_n10358_), .A1(\A[385] ), .B0(\A[387] ), .Y(new_n10467_));
  NAND2  g09465(.A(new_n10362_), .B(new_n10357_), .Y(new_n10468_));
  OAI21  g09466(.A0(new_n10467_), .A1(new_n10466_), .B0(new_n10468_), .Y(new_n10469_));
  XOR2   g09467(.A(new_n10370_), .B(new_n10469_), .Y(new_n10470_));
  XOR2   g09468(.A(new_n10374_), .B(new_n10372_), .Y(new_n10471_));
  NOR2   g09469(.A(new_n10370_), .B(new_n10363_), .Y(new_n10472_));
  NAND2  g09470(.A(\A[389] ), .B(\A[388] ), .Y(new_n10473_));
  NAND2  g09471(.A(new_n10369_), .B(\A[390] ), .Y(new_n10474_));
  NAND2  g09472(.A(\A[386] ), .B(\A[385] ), .Y(new_n10475_));
  NAND2  g09473(.A(new_n10362_), .B(\A[387] ), .Y(new_n10476_));
  AOI22  g09474(.A0(new_n10476_), .A1(new_n10475_), .B0(new_n10474_), .B1(new_n10473_), .Y(new_n10477_));
  AOI21  g09475(.A0(new_n10472_), .A1(new_n10471_), .B0(new_n10477_), .Y(new_n10478_));
  XOR2   g09476(.A(new_n10472_), .B(new_n10471_), .Y(new_n10479_));
  XOR2   g09477(.A(new_n10370_), .B(new_n10363_), .Y(new_n10480_));
  NOR2   g09478(.A(\A[389] ), .B(new_n10367_), .Y(new_n10481_));
  OAI21  g09479(.A0(new_n10365_), .A1(\A[388] ), .B0(\A[390] ), .Y(new_n10482_));
  NAND2  g09480(.A(new_n10369_), .B(new_n10364_), .Y(new_n10483_));
  OAI21  g09481(.A0(new_n10482_), .A1(new_n10481_), .B0(new_n10483_), .Y(new_n10484_));
  NAND2  g09482(.A(new_n10474_), .B(new_n10473_), .Y(new_n10485_));
  NAND2  g09483(.A(new_n10476_), .B(new_n10475_), .Y(new_n10486_));
  NAND4  g09484(.A(new_n10486_), .B(new_n10485_), .C(new_n10484_), .D(new_n10469_), .Y(new_n10487_));
  NAND4  g09485(.A(new_n10460_), .B(new_n10449_), .C(new_n10457_), .D(new_n10454_), .Y(new_n10488_));
  NAND4  g09486(.A(new_n10488_), .B(new_n10446_), .C(new_n10487_), .D(new_n10480_), .Y(new_n10489_));
  OAI211 g09487(.A0(new_n10478_), .A1(new_n10470_), .B0(new_n10489_), .B1(new_n10479_), .Y(new_n10490_));
  XOR2   g09488(.A(new_n10374_), .B(new_n10485_), .Y(new_n10491_));
  XOR2   g09489(.A(new_n10472_), .B(new_n10491_), .Y(new_n10492_));
  NOR4   g09490(.A(new_n10374_), .B(new_n10372_), .C(new_n10370_), .D(new_n10363_), .Y(new_n10493_));
  XOR2   g09491(.A(new_n10389_), .B(new_n10454_), .Y(new_n10494_));
  NOR4   g09492(.A(new_n10393_), .B(new_n10391_), .C(new_n10389_), .D(new_n10382_), .Y(new_n10495_));
  NOR4   g09493(.A(new_n10495_), .B(new_n10494_), .C(new_n10493_), .D(new_n10470_), .Y(new_n10496_));
  AOI221 g09494(.A0(new_n10474_), .A1(new_n10473_), .C0(new_n10373_), .B0(new_n10362_), .B1(\A[387] ), .Y(new_n10497_));
  AOI221 g09495(.A0(new_n10476_), .A1(new_n10475_), .C0(new_n10371_), .B0(new_n10369_), .B1(\A[390] ), .Y(new_n10498_));
  OAI211 g09496(.A0(new_n10498_), .A1(new_n10497_), .B0(new_n10484_), .B1(new_n10469_), .Y(new_n10499_));
  NAND2  g09497(.A(new_n10486_), .B(new_n10485_), .Y(new_n10500_));
  AOI21  g09498(.A0(new_n10500_), .A1(new_n10499_), .B0(new_n10470_), .Y(new_n10501_));
  OAI21  g09499(.A0(new_n10501_), .A1(new_n10492_), .B0(new_n10496_), .Y(new_n10502_));
  AOI21  g09500(.A0(new_n10502_), .A1(new_n10490_), .B0(new_n10465_), .Y(new_n10503_));
  OAI21  g09501(.A0(new_n10501_), .A1(new_n10492_), .B0(new_n10489_), .Y(new_n10504_));
  NAND4  g09502(.A(new_n10446_), .B(new_n10479_), .C(new_n10478_), .D(new_n10480_), .Y(new_n10505_));
  OAI21  g09503(.A0(new_n10478_), .A1(new_n10470_), .B0(new_n10488_), .Y(new_n10506_));
  OAI21  g09504(.A0(new_n10506_), .A1(new_n10505_), .B0(new_n10504_), .Y(new_n10507_));
  NAND2  g09505(.A(new_n10398_), .B(\A[373] ), .Y(new_n10508_));
  AOI21  g09506(.A0(\A[374] ), .A1(new_n10396_), .B0(new_n10400_), .Y(new_n10509_));
  AOI22  g09507(.A0(new_n10401_), .A1(new_n10400_), .B0(new_n10509_), .B1(new_n10508_), .Y(new_n10510_));
  XOR2   g09508(.A(new_n10410_), .B(new_n10510_), .Y(new_n10511_));
  XOR2   g09509(.A(new_n10434_), .B(new_n10511_), .Y(new_n10512_));
  NAND2  g09510(.A(new_n10512_), .B(new_n10395_), .Y(new_n10513_));
  AOI211 g09511(.A0(new_n10507_), .A1(new_n10465_), .B(new_n10513_), .C(new_n10503_), .Y(new_n10514_));
  XOR2   g09512(.A(new_n10370_), .B(new_n10469_), .Y(new_n10515_));
  XOR2   g09513(.A(new_n10394_), .B(new_n10515_), .Y(new_n10516_));
  NOR2   g09514(.A(new_n10435_), .B(new_n10516_), .Y(new_n10517_));
  AOI21  g09515(.A0(new_n10507_), .A1(new_n10465_), .B0(new_n10503_), .Y(new_n10518_));
  NOR2   g09516(.A(new_n10518_), .B(new_n10517_), .Y(new_n10519_));
  XOR2   g09517(.A(new_n10429_), .B(new_n10422_), .Y(new_n10520_));
  XOR2   g09518(.A(\A[371] ), .B(new_n10426_), .Y(new_n10521_));
  NAND2  g09519(.A(\A[371] ), .B(\A[370] ), .Y(new_n10522_));
  OAI21  g09520(.A0(new_n10521_), .A1(new_n10423_), .B0(new_n10522_), .Y(new_n10523_));
  XOR2   g09521(.A(new_n10433_), .B(new_n10523_), .Y(new_n10524_));
  NOR2   g09522(.A(\A[368] ), .B(new_n10419_), .Y(new_n10525_));
  OAI21  g09523(.A0(new_n10417_), .A1(\A[367] ), .B0(\A[369] ), .Y(new_n10526_));
  XOR2   g09524(.A(\A[368] ), .B(new_n10419_), .Y(new_n10527_));
  OAI22  g09525(.A0(new_n10527_), .A1(\A[369] ), .B0(new_n10526_), .B1(new_n10525_), .Y(new_n10528_));
  NOR2   g09526(.A(\A[371] ), .B(new_n10426_), .Y(new_n10529_));
  OAI21  g09527(.A0(new_n10424_), .A1(\A[370] ), .B0(\A[372] ), .Y(new_n10530_));
  OAI22  g09528(.A0(new_n10521_), .A1(\A[372] ), .B0(new_n10530_), .B1(new_n10529_), .Y(new_n10531_));
  NAND2  g09529(.A(new_n10531_), .B(new_n10528_), .Y(new_n10532_));
  NAND2  g09530(.A(\A[368] ), .B(\A[367] ), .Y(new_n10533_));
  OAI21  g09531(.A0(new_n10527_), .A1(new_n10416_), .B0(new_n10533_), .Y(new_n10534_));
  NAND2  g09532(.A(new_n10534_), .B(new_n10523_), .Y(new_n10535_));
  OAI21  g09533(.A0(new_n10532_), .A1(new_n10524_), .B0(new_n10535_), .Y(new_n10536_));
  NOR2   g09534(.A(new_n10429_), .B(new_n10422_), .Y(new_n10537_));
  XOR2   g09535(.A(new_n10537_), .B(new_n10524_), .Y(new_n10538_));
  AOI21  g09536(.A0(new_n10536_), .A1(new_n10520_), .B0(new_n10538_), .Y(new_n10539_));
  XOR2   g09537(.A(new_n10410_), .B(new_n10403_), .Y(new_n10540_));
  XOR2   g09538(.A(new_n10414_), .B(new_n10412_), .Y(new_n10541_));
  NOR2   g09539(.A(new_n10410_), .B(new_n10510_), .Y(new_n10542_));
  NAND2  g09540(.A(\A[377] ), .B(\A[376] ), .Y(new_n10543_));
  NAND2  g09541(.A(new_n10409_), .B(\A[378] ), .Y(new_n10544_));
  NAND2  g09542(.A(\A[374] ), .B(\A[373] ), .Y(new_n10545_));
  NAND2  g09543(.A(new_n10401_), .B(\A[375] ), .Y(new_n10546_));
  AOI22  g09544(.A0(new_n10546_), .A1(new_n10545_), .B0(new_n10544_), .B1(new_n10543_), .Y(new_n10547_));
  AOI21  g09545(.A0(new_n10542_), .A1(new_n10541_), .B0(new_n10547_), .Y(new_n10548_));
  XOR2   g09546(.A(new_n10542_), .B(new_n10541_), .Y(new_n10549_));
  XOR2   g09547(.A(new_n10410_), .B(new_n10510_), .Y(new_n10550_));
  NOR2   g09548(.A(\A[377] ), .B(new_n10407_), .Y(new_n10551_));
  OAI21  g09549(.A0(new_n10405_), .A1(\A[376] ), .B0(\A[378] ), .Y(new_n10552_));
  NAND2  g09550(.A(new_n10409_), .B(new_n10404_), .Y(new_n10553_));
  OAI21  g09551(.A0(new_n10552_), .A1(new_n10551_), .B0(new_n10553_), .Y(new_n10554_));
  NAND2  g09552(.A(new_n10544_), .B(new_n10543_), .Y(new_n10555_));
  NAND2  g09553(.A(new_n10546_), .B(new_n10545_), .Y(new_n10556_));
  NAND4  g09554(.A(new_n10556_), .B(new_n10555_), .C(new_n10554_), .D(new_n10403_), .Y(new_n10557_));
  NAND4  g09555(.A(new_n10534_), .B(new_n10523_), .C(new_n10531_), .D(new_n10528_), .Y(new_n10558_));
  NAND4  g09556(.A(new_n10558_), .B(new_n10520_), .C(new_n10557_), .D(new_n10550_), .Y(new_n10559_));
  OAI211 g09557(.A0(new_n10548_), .A1(new_n10540_), .B0(new_n10559_), .B1(new_n10549_), .Y(new_n10560_));
  XOR2   g09558(.A(new_n10414_), .B(new_n10555_), .Y(new_n10561_));
  XOR2   g09559(.A(new_n10542_), .B(new_n10561_), .Y(new_n10562_));
  NOR4   g09560(.A(new_n10414_), .B(new_n10412_), .C(new_n10410_), .D(new_n10510_), .Y(new_n10563_));
  XOR2   g09561(.A(new_n10429_), .B(new_n10528_), .Y(new_n10564_));
  NOR4   g09562(.A(new_n10433_), .B(new_n10431_), .C(new_n10429_), .D(new_n10422_), .Y(new_n10565_));
  NOR4   g09563(.A(new_n10565_), .B(new_n10564_), .C(new_n10563_), .D(new_n10540_), .Y(new_n10566_));
  AOI221 g09564(.A0(new_n10544_), .A1(new_n10543_), .C0(new_n10413_), .B0(new_n10401_), .B1(\A[375] ), .Y(new_n10567_));
  AOI221 g09565(.A0(new_n10546_), .A1(new_n10545_), .C0(new_n10411_), .B0(new_n10409_), .B1(\A[378] ), .Y(new_n10568_));
  OAI211 g09566(.A0(new_n10568_), .A1(new_n10567_), .B0(new_n10554_), .B1(new_n10403_), .Y(new_n10569_));
  NAND2  g09567(.A(new_n10556_), .B(new_n10555_), .Y(new_n10570_));
  AOI21  g09568(.A0(new_n10570_), .A1(new_n10569_), .B0(new_n10540_), .Y(new_n10571_));
  OAI21  g09569(.A0(new_n10571_), .A1(new_n10562_), .B0(new_n10566_), .Y(new_n10572_));
  AOI21  g09570(.A0(new_n10572_), .A1(new_n10560_), .B0(new_n10539_), .Y(new_n10573_));
  NOR2   g09571(.A(new_n10571_), .B(new_n10562_), .Y(new_n10574_));
  NAND4  g09572(.A(new_n10520_), .B(new_n10549_), .C(new_n10548_), .D(new_n10550_), .Y(new_n10575_));
  OAI21  g09573(.A0(new_n10548_), .A1(new_n10540_), .B0(new_n10558_), .Y(new_n10576_));
  OAI22  g09574(.A0(new_n10576_), .A1(new_n10575_), .B0(new_n10574_), .B1(new_n10566_), .Y(new_n10577_));
  AOI21  g09575(.A0(new_n10577_), .A1(new_n10539_), .B0(new_n10573_), .Y(new_n10578_));
  OAI21  g09576(.A0(new_n10519_), .A1(new_n10514_), .B0(new_n10578_), .Y(new_n10579_));
  XOR2   g09577(.A(new_n10574_), .B(new_n10559_), .Y(new_n10580_));
  NAND2  g09578(.A(new_n10577_), .B(new_n10539_), .Y(new_n10581_));
  OAI21  g09579(.A0(new_n10580_), .A1(new_n10539_), .B0(new_n10581_), .Y(new_n10582_));
  AOI211 g09580(.A0(new_n10507_), .A1(new_n10465_), .B(new_n10517_), .C(new_n10503_), .Y(new_n10583_));
  NOR2   g09581(.A(new_n10518_), .B(new_n10513_), .Y(new_n10584_));
  OAI21  g09582(.A0(new_n10584_), .A1(new_n10583_), .B0(new_n10582_), .Y(new_n10585_));
  NAND2  g09583(.A(new_n10585_), .B(new_n10579_), .Y(new_n10586_));
  AOI21  g09584(.A0(new_n10445_), .A1(new_n10438_), .B0(new_n10586_), .Y(new_n10587_));
  XOR2   g09585(.A(new_n10393_), .B(new_n10391_), .Y(new_n10588_));
  NOR2   g09586(.A(new_n10393_), .B(new_n10391_), .Y(new_n10589_));
  AOI21  g09587(.A0(new_n10463_), .A1(new_n10588_), .B0(new_n10589_), .Y(new_n10590_));
  XOR2   g09588(.A(new_n10463_), .B(new_n10588_), .Y(new_n10591_));
  OAI21  g09589(.A0(new_n10590_), .A1(new_n10494_), .B0(new_n10591_), .Y(new_n10592_));
  OAI21  g09590(.A0(new_n10478_), .A1(new_n10470_), .B0(new_n10479_), .Y(new_n10593_));
  XOR2   g09591(.A(new_n10593_), .B(new_n10489_), .Y(new_n10594_));
  NAND2  g09592(.A(new_n10594_), .B(new_n10592_), .Y(new_n10595_));
  NAND2  g09593(.A(new_n10507_), .B(new_n10465_), .Y(new_n10596_));
  NAND3  g09594(.A(new_n10517_), .B(new_n10596_), .C(new_n10595_), .Y(new_n10597_));
  NAND2  g09595(.A(new_n10500_), .B(new_n10499_), .Y(new_n10598_));
  NOR4   g09596(.A(new_n10494_), .B(new_n10492_), .C(new_n10598_), .D(new_n10470_), .Y(new_n10599_));
  OAI211 g09597(.A0(new_n10478_), .A1(new_n10470_), .B0(new_n10599_), .B1(new_n10488_), .Y(new_n10600_));
  AOI21  g09598(.A0(new_n10600_), .A1(new_n10504_), .B0(new_n10592_), .Y(new_n10601_));
  OAI21  g09599(.A0(new_n10601_), .A1(new_n10503_), .B0(new_n10513_), .Y(new_n10602_));
  AOI21  g09600(.A0(new_n10602_), .A1(new_n10597_), .B0(new_n10582_), .Y(new_n10603_));
  NAND3  g09601(.A(new_n10513_), .B(new_n10596_), .C(new_n10595_), .Y(new_n10604_));
  OAI21  g09602(.A0(new_n10518_), .A1(new_n10513_), .B0(new_n10604_), .Y(new_n10605_));
  AOI21  g09603(.A0(new_n10605_), .A1(new_n10582_), .B0(new_n10603_), .Y(new_n10606_));
  AOI21  g09604(.A0(new_n10354_), .A1(new_n10347_), .B0(new_n10437_), .Y(new_n10607_));
  NAND2  g09605(.A(new_n10607_), .B(new_n10341_), .Y(new_n10608_));
  OAI21  g09606(.A0(new_n10443_), .A1(new_n10441_), .B0(new_n10437_), .Y(new_n10609_));
  AOI21  g09607(.A0(new_n10609_), .A1(new_n10608_), .B0(new_n10606_), .Y(new_n10610_));
  NOR2   g09608(.A(new_n10610_), .B(new_n10587_), .Y(new_n10611_));
  INV    g09609(.A(\A[429] ), .Y(new_n10612_));
  INV    g09610(.A(\A[427] ), .Y(new_n10613_));
  NAND2  g09611(.A(\A[428] ), .B(new_n10613_), .Y(new_n10614_));
  INV    g09612(.A(\A[428] ), .Y(new_n10615_));
  AOI21  g09613(.A0(new_n10615_), .A1(\A[427] ), .B0(new_n10612_), .Y(new_n10616_));
  XOR2   g09614(.A(\A[428] ), .B(\A[427] ), .Y(new_n10617_));
  AOI22  g09615(.A0(new_n10617_), .A1(new_n10612_), .B0(new_n10616_), .B1(new_n10614_), .Y(new_n10618_));
  INV    g09616(.A(\A[432] ), .Y(new_n10619_));
  INV    g09617(.A(\A[430] ), .Y(new_n10620_));
  NAND2  g09618(.A(\A[431] ), .B(new_n10620_), .Y(new_n10621_));
  INV    g09619(.A(\A[431] ), .Y(new_n10622_));
  AOI21  g09620(.A0(new_n10622_), .A1(\A[430] ), .B0(new_n10619_), .Y(new_n10623_));
  XOR2   g09621(.A(\A[431] ), .B(\A[430] ), .Y(new_n10624_));
  AOI22  g09622(.A0(new_n10624_), .A1(new_n10619_), .B0(new_n10623_), .B1(new_n10621_), .Y(new_n10625_));
  NOR2   g09623(.A(new_n10625_), .B(new_n10618_), .Y(new_n10626_));
  XOR2   g09624(.A(\A[431] ), .B(new_n10620_), .Y(new_n10627_));
  NAND2  g09625(.A(\A[431] ), .B(\A[430] ), .Y(new_n10628_));
  OAI21  g09626(.A0(new_n10627_), .A1(new_n10619_), .B0(new_n10628_), .Y(new_n10629_));
  NOR2   g09627(.A(new_n10615_), .B(new_n10613_), .Y(new_n10630_));
  AOI21  g09628(.A0(new_n10617_), .A1(\A[429] ), .B0(new_n10630_), .Y(new_n10631_));
  XOR2   g09629(.A(new_n10631_), .B(new_n10629_), .Y(new_n10632_));
  XOR2   g09630(.A(new_n10632_), .B(new_n10626_), .Y(new_n10633_));
  XOR2   g09631(.A(new_n10625_), .B(new_n10618_), .Y(new_n10634_));
  NOR2   g09632(.A(new_n10615_), .B(\A[427] ), .Y(new_n10635_));
  OAI21  g09633(.A0(\A[428] ), .A1(new_n10613_), .B0(\A[429] ), .Y(new_n10636_));
  XOR2   g09634(.A(\A[428] ), .B(new_n10613_), .Y(new_n10637_));
  OAI22  g09635(.A0(new_n10637_), .A1(\A[429] ), .B0(new_n10636_), .B1(new_n10635_), .Y(new_n10638_));
  NOR2   g09636(.A(new_n10622_), .B(\A[430] ), .Y(new_n10639_));
  OAI21  g09637(.A0(\A[431] ), .A1(new_n10620_), .B0(\A[432] ), .Y(new_n10640_));
  OAI22  g09638(.A0(new_n10627_), .A1(\A[432] ), .B0(new_n10640_), .B1(new_n10639_), .Y(new_n10641_));
  NAND2  g09639(.A(new_n10641_), .B(new_n10638_), .Y(new_n10642_));
  NAND2  g09640(.A(\A[428] ), .B(\A[427] ), .Y(new_n10643_));
  OAI21  g09641(.A0(new_n10637_), .A1(new_n10612_), .B0(new_n10643_), .Y(new_n10644_));
  NAND2  g09642(.A(new_n10644_), .B(new_n10629_), .Y(new_n10645_));
  OAI21  g09643(.A0(new_n10632_), .A1(new_n10642_), .B0(new_n10645_), .Y(new_n10646_));
  AOI21  g09644(.A0(new_n10646_), .A1(new_n10634_), .B0(new_n10633_), .Y(new_n10647_));
  NAND2  g09645(.A(\A[437] ), .B(\A[436] ), .Y(new_n10648_));
  XOR2   g09646(.A(\A[437] ), .B(\A[436] ), .Y(new_n10649_));
  NAND2  g09647(.A(new_n10649_), .B(\A[438] ), .Y(new_n10650_));
  NAND2  g09648(.A(new_n10650_), .B(new_n10648_), .Y(new_n10651_));
  NAND2  g09649(.A(\A[434] ), .B(\A[433] ), .Y(new_n10652_));
  XOR2   g09650(.A(\A[434] ), .B(\A[433] ), .Y(new_n10653_));
  NAND2  g09651(.A(new_n10653_), .B(\A[435] ), .Y(new_n10654_));
  NAND2  g09652(.A(new_n10654_), .B(new_n10652_), .Y(new_n10655_));
  XOR2   g09653(.A(new_n10655_), .B(new_n10651_), .Y(new_n10656_));
  INV    g09654(.A(\A[435] ), .Y(new_n10657_));
  INV    g09655(.A(\A[433] ), .Y(new_n10658_));
  NAND2  g09656(.A(\A[434] ), .B(new_n10658_), .Y(new_n10659_));
  INV    g09657(.A(\A[434] ), .Y(new_n10660_));
  AOI21  g09658(.A0(new_n10660_), .A1(\A[433] ), .B0(new_n10657_), .Y(new_n10661_));
  AOI22  g09659(.A0(new_n10661_), .A1(new_n10659_), .B0(new_n10653_), .B1(new_n10657_), .Y(new_n10662_));
  INV    g09660(.A(\A[438] ), .Y(new_n10663_));
  INV    g09661(.A(\A[436] ), .Y(new_n10664_));
  NAND2  g09662(.A(\A[437] ), .B(new_n10664_), .Y(new_n10665_));
  INV    g09663(.A(\A[437] ), .Y(new_n10666_));
  AOI21  g09664(.A0(new_n10666_), .A1(\A[436] ), .B0(new_n10663_), .Y(new_n10667_));
  AOI22  g09665(.A0(new_n10667_), .A1(new_n10665_), .B0(new_n10649_), .B1(new_n10663_), .Y(new_n10668_));
  NOR2   g09666(.A(new_n10668_), .B(new_n10662_), .Y(new_n10669_));
  AOI22  g09667(.A0(new_n10654_), .A1(new_n10652_), .B0(new_n10650_), .B1(new_n10648_), .Y(new_n10670_));
  AOI21  g09668(.A0(new_n10669_), .A1(new_n10656_), .B0(new_n10670_), .Y(new_n10671_));
  XOR2   g09669(.A(new_n10669_), .B(new_n10656_), .Y(new_n10672_));
  NOR2   g09670(.A(new_n10660_), .B(\A[433] ), .Y(new_n10673_));
  OAI21  g09671(.A0(\A[434] ), .A1(new_n10658_), .B0(\A[435] ), .Y(new_n10674_));
  NAND2  g09672(.A(new_n10653_), .B(new_n10657_), .Y(new_n10675_));
  OAI21  g09673(.A0(new_n10674_), .A1(new_n10673_), .B0(new_n10675_), .Y(new_n10676_));
  XOR2   g09674(.A(new_n10668_), .B(new_n10676_), .Y(new_n10677_));
  NOR2   g09675(.A(new_n10666_), .B(\A[436] ), .Y(new_n10678_));
  OAI21  g09676(.A0(\A[437] ), .A1(new_n10664_), .B0(\A[438] ), .Y(new_n10679_));
  NAND2  g09677(.A(new_n10649_), .B(new_n10663_), .Y(new_n10680_));
  OAI21  g09678(.A0(new_n10679_), .A1(new_n10678_), .B0(new_n10680_), .Y(new_n10681_));
  NAND4  g09679(.A(new_n10681_), .B(new_n10676_), .C(new_n10655_), .D(new_n10651_), .Y(new_n10682_));
  NAND4  g09680(.A(new_n10644_), .B(new_n10629_), .C(new_n10641_), .D(new_n10638_), .Y(new_n10683_));
  XOR2   g09681(.A(new_n10668_), .B(new_n10662_), .Y(new_n10684_));
  NAND4  g09682(.A(new_n10684_), .B(new_n10683_), .C(new_n10682_), .D(new_n10634_), .Y(new_n10685_));
  OAI211 g09683(.A0(new_n10677_), .A1(new_n10671_), .B0(new_n10685_), .B1(new_n10672_), .Y(new_n10686_));
  NOR2   g09684(.A(new_n10660_), .B(new_n10658_), .Y(new_n10687_));
  AOI21  g09685(.A0(new_n10653_), .A1(\A[435] ), .B0(new_n10687_), .Y(new_n10688_));
  XOR2   g09686(.A(new_n10688_), .B(new_n10651_), .Y(new_n10689_));
  XOR2   g09687(.A(new_n10669_), .B(new_n10689_), .Y(new_n10690_));
  XOR2   g09688(.A(new_n10625_), .B(new_n10638_), .Y(new_n10691_));
  NOR2   g09689(.A(new_n10666_), .B(new_n10664_), .Y(new_n10692_));
  AOI21  g09690(.A0(new_n10649_), .A1(\A[438] ), .B0(new_n10692_), .Y(new_n10693_));
  NOR4   g09691(.A(new_n10668_), .B(new_n10662_), .C(new_n10688_), .D(new_n10693_), .Y(new_n10694_));
  NOR2   g09692(.A(new_n10622_), .B(new_n10620_), .Y(new_n10695_));
  AOI21  g09693(.A0(new_n10624_), .A1(\A[432] ), .B0(new_n10695_), .Y(new_n10696_));
  NOR4   g09694(.A(new_n10631_), .B(new_n10696_), .C(new_n10625_), .D(new_n10618_), .Y(new_n10697_));
  NOR4   g09695(.A(new_n10677_), .B(new_n10697_), .C(new_n10694_), .D(new_n10691_), .Y(new_n10698_));
  AOI221 g09696(.A0(new_n10653_), .A1(\A[435] ), .C0(new_n10687_), .B0(new_n10650_), .B1(new_n10648_), .Y(new_n10699_));
  AOI221 g09697(.A0(new_n10654_), .A1(new_n10652_), .C0(new_n10692_), .B0(new_n10649_), .B1(\A[438] ), .Y(new_n10700_));
  OAI211 g09698(.A0(new_n10700_), .A1(new_n10699_), .B0(new_n10681_), .B1(new_n10676_), .Y(new_n10701_));
  NAND2  g09699(.A(new_n10655_), .B(new_n10651_), .Y(new_n10702_));
  AOI21  g09700(.A0(new_n10702_), .A1(new_n10701_), .B0(new_n10677_), .Y(new_n10703_));
  OAI21  g09701(.A0(new_n10703_), .A1(new_n10690_), .B0(new_n10698_), .Y(new_n10704_));
  AOI21  g09702(.A0(new_n10704_), .A1(new_n10686_), .B0(new_n10647_), .Y(new_n10705_));
  XOR2   g09703(.A(new_n10632_), .B(new_n10642_), .Y(new_n10706_));
  XOR2   g09704(.A(new_n10631_), .B(new_n10696_), .Y(new_n10707_));
  NOR2   g09705(.A(new_n10631_), .B(new_n10696_), .Y(new_n10708_));
  AOI21  g09706(.A0(new_n10707_), .A1(new_n10626_), .B0(new_n10708_), .Y(new_n10709_));
  OAI21  g09707(.A0(new_n10709_), .A1(new_n10691_), .B0(new_n10706_), .Y(new_n10710_));
  OAI21  g09708(.A0(new_n10703_), .A1(new_n10690_), .B0(new_n10685_), .Y(new_n10711_));
  NOR2   g09709(.A(new_n10677_), .B(new_n10691_), .Y(new_n10712_));
  OAI211 g09710(.A0(new_n10681_), .A1(new_n10676_), .B0(new_n10655_), .B1(new_n10651_), .Y(new_n10713_));
  NAND4  g09711(.A(new_n10713_), .B(new_n10712_), .C(new_n10683_), .D(new_n10672_), .Y(new_n10714_));
  AOI21  g09712(.A0(new_n10714_), .A1(new_n10711_), .B0(new_n10710_), .Y(new_n10715_));
  NOR2   g09713(.A(new_n10677_), .B(new_n10694_), .Y(new_n10716_));
  XOR2   g09714(.A(new_n10625_), .B(new_n10618_), .Y(new_n10717_));
  XOR2   g09715(.A(new_n10717_), .B(new_n10716_), .Y(new_n10718_));
  INV    g09716(.A(\A[423] ), .Y(new_n10719_));
  INV    g09717(.A(\A[422] ), .Y(new_n10720_));
  NAND2  g09718(.A(new_n10720_), .B(\A[421] ), .Y(new_n10721_));
  INV    g09719(.A(\A[421] ), .Y(new_n10722_));
  AOI21  g09720(.A0(\A[422] ), .A1(new_n10722_), .B0(new_n10719_), .Y(new_n10723_));
  XOR2   g09721(.A(\A[422] ), .B(\A[421] ), .Y(new_n10724_));
  AOI22  g09722(.A0(new_n10724_), .A1(new_n10719_), .B0(new_n10723_), .B1(new_n10721_), .Y(new_n10725_));
  INV    g09723(.A(\A[426] ), .Y(new_n10726_));
  INV    g09724(.A(\A[425] ), .Y(new_n10727_));
  NAND2  g09725(.A(new_n10727_), .B(\A[424] ), .Y(new_n10728_));
  INV    g09726(.A(\A[424] ), .Y(new_n10729_));
  AOI21  g09727(.A0(\A[425] ), .A1(new_n10729_), .B0(new_n10726_), .Y(new_n10730_));
  XOR2   g09728(.A(\A[425] ), .B(\A[424] ), .Y(new_n10731_));
  AOI22  g09729(.A0(new_n10731_), .A1(new_n10726_), .B0(new_n10730_), .B1(new_n10728_), .Y(new_n10732_));
  NOR2   g09730(.A(new_n10727_), .B(new_n10729_), .Y(new_n10733_));
  AOI21  g09731(.A0(new_n10731_), .A1(\A[426] ), .B0(new_n10733_), .Y(new_n10734_));
  NOR2   g09732(.A(new_n10720_), .B(new_n10722_), .Y(new_n10735_));
  AOI21  g09733(.A0(new_n10724_), .A1(\A[423] ), .B0(new_n10735_), .Y(new_n10736_));
  XOR2   g09734(.A(new_n10732_), .B(new_n10725_), .Y(new_n10737_));
  INV    g09735(.A(\A[417] ), .Y(new_n10738_));
  INV    g09736(.A(\A[416] ), .Y(new_n10739_));
  NAND2  g09737(.A(new_n10739_), .B(\A[415] ), .Y(new_n10740_));
  INV    g09738(.A(\A[415] ), .Y(new_n10741_));
  AOI21  g09739(.A0(\A[416] ), .A1(new_n10741_), .B0(new_n10738_), .Y(new_n10742_));
  XOR2   g09740(.A(\A[416] ), .B(\A[415] ), .Y(new_n10743_));
  AOI22  g09741(.A0(new_n10743_), .A1(new_n10738_), .B0(new_n10742_), .B1(new_n10740_), .Y(new_n10744_));
  INV    g09742(.A(\A[420] ), .Y(new_n10745_));
  INV    g09743(.A(\A[419] ), .Y(new_n10746_));
  NAND2  g09744(.A(new_n10746_), .B(\A[418] ), .Y(new_n10747_));
  INV    g09745(.A(\A[418] ), .Y(new_n10748_));
  AOI21  g09746(.A0(\A[419] ), .A1(new_n10748_), .B0(new_n10745_), .Y(new_n10749_));
  XOR2   g09747(.A(\A[419] ), .B(\A[418] ), .Y(new_n10750_));
  AOI22  g09748(.A0(new_n10750_), .A1(new_n10745_), .B0(new_n10749_), .B1(new_n10747_), .Y(new_n10751_));
  NOR2   g09749(.A(new_n10746_), .B(new_n10748_), .Y(new_n10752_));
  AOI21  g09750(.A0(new_n10750_), .A1(\A[420] ), .B0(new_n10752_), .Y(new_n10753_));
  NOR2   g09751(.A(new_n10739_), .B(new_n10741_), .Y(new_n10754_));
  AOI21  g09752(.A0(new_n10743_), .A1(\A[417] ), .B0(new_n10754_), .Y(new_n10755_));
  XOR2   g09753(.A(new_n10751_), .B(new_n10744_), .Y(new_n10756_));
  XOR2   g09754(.A(new_n10756_), .B(new_n10737_), .Y(new_n10757_));
  NAND2  g09755(.A(new_n10757_), .B(new_n10718_), .Y(new_n10758_));
  NOR3   g09756(.A(new_n10758_), .B(new_n10715_), .C(new_n10705_), .Y(new_n10759_));
  OAI21  g09757(.A0(new_n10677_), .A1(new_n10671_), .B0(new_n10672_), .Y(new_n10760_));
  XOR2   g09758(.A(new_n10760_), .B(new_n10685_), .Y(new_n10761_));
  NAND2  g09759(.A(new_n10761_), .B(new_n10710_), .Y(new_n10762_));
  NAND2  g09760(.A(new_n10714_), .B(new_n10711_), .Y(new_n10763_));
  NAND2  g09761(.A(new_n10763_), .B(new_n10647_), .Y(new_n10764_));
  NAND2  g09762(.A(new_n10684_), .B(new_n10682_), .Y(new_n10765_));
  XOR2   g09763(.A(new_n10717_), .B(new_n10765_), .Y(new_n10766_));
  NOR2   g09764(.A(\A[422] ), .B(new_n10722_), .Y(new_n10767_));
  OAI21  g09765(.A0(new_n10720_), .A1(\A[421] ), .B0(\A[423] ), .Y(new_n10768_));
  NAND2  g09766(.A(new_n10724_), .B(new_n10719_), .Y(new_n10769_));
  OAI21  g09767(.A0(new_n10768_), .A1(new_n10767_), .B0(new_n10769_), .Y(new_n10770_));
  XOR2   g09768(.A(new_n10732_), .B(new_n10770_), .Y(new_n10771_));
  XOR2   g09769(.A(new_n10756_), .B(new_n10771_), .Y(new_n10772_));
  NOR2   g09770(.A(new_n10772_), .B(new_n10766_), .Y(new_n10773_));
  AOI21  g09771(.A0(new_n10764_), .A1(new_n10762_), .B0(new_n10773_), .Y(new_n10774_));
  XOR2   g09772(.A(new_n10751_), .B(new_n10744_), .Y(new_n10775_));
  XOR2   g09773(.A(\A[419] ), .B(new_n10748_), .Y(new_n10776_));
  NAND2  g09774(.A(\A[419] ), .B(\A[418] ), .Y(new_n10777_));
  OAI21  g09775(.A0(new_n10776_), .A1(new_n10745_), .B0(new_n10777_), .Y(new_n10778_));
  XOR2   g09776(.A(new_n10755_), .B(new_n10778_), .Y(new_n10779_));
  NOR2   g09777(.A(\A[416] ), .B(new_n10741_), .Y(new_n10780_));
  OAI21  g09778(.A0(new_n10739_), .A1(\A[415] ), .B0(\A[417] ), .Y(new_n10781_));
  XOR2   g09779(.A(\A[416] ), .B(new_n10741_), .Y(new_n10782_));
  OAI22  g09780(.A0(new_n10782_), .A1(\A[417] ), .B0(new_n10781_), .B1(new_n10780_), .Y(new_n10783_));
  NOR2   g09781(.A(\A[419] ), .B(new_n10748_), .Y(new_n10784_));
  OAI21  g09782(.A0(new_n10746_), .A1(\A[418] ), .B0(\A[420] ), .Y(new_n10785_));
  OAI22  g09783(.A0(new_n10776_), .A1(\A[420] ), .B0(new_n10785_), .B1(new_n10784_), .Y(new_n10786_));
  NAND2  g09784(.A(new_n10786_), .B(new_n10783_), .Y(new_n10787_));
  NAND2  g09785(.A(\A[416] ), .B(\A[415] ), .Y(new_n10788_));
  OAI21  g09786(.A0(new_n10782_), .A1(new_n10738_), .B0(new_n10788_), .Y(new_n10789_));
  NAND2  g09787(.A(new_n10789_), .B(new_n10778_), .Y(new_n10790_));
  OAI21  g09788(.A0(new_n10787_), .A1(new_n10779_), .B0(new_n10790_), .Y(new_n10791_));
  NOR2   g09789(.A(new_n10751_), .B(new_n10744_), .Y(new_n10792_));
  XOR2   g09790(.A(new_n10792_), .B(new_n10779_), .Y(new_n10793_));
  AOI21  g09791(.A0(new_n10791_), .A1(new_n10775_), .B0(new_n10793_), .Y(new_n10794_));
  XOR2   g09792(.A(new_n10732_), .B(new_n10770_), .Y(new_n10795_));
  XOR2   g09793(.A(new_n10736_), .B(new_n10734_), .Y(new_n10796_));
  NOR2   g09794(.A(new_n10732_), .B(new_n10725_), .Y(new_n10797_));
  NAND2  g09795(.A(\A[425] ), .B(\A[424] ), .Y(new_n10798_));
  NAND2  g09796(.A(new_n10731_), .B(\A[426] ), .Y(new_n10799_));
  NAND2  g09797(.A(\A[422] ), .B(\A[421] ), .Y(new_n10800_));
  NAND2  g09798(.A(new_n10724_), .B(\A[423] ), .Y(new_n10801_));
  AOI22  g09799(.A0(new_n10801_), .A1(new_n10800_), .B0(new_n10799_), .B1(new_n10798_), .Y(new_n10802_));
  AOI21  g09800(.A0(new_n10797_), .A1(new_n10796_), .B0(new_n10802_), .Y(new_n10803_));
  XOR2   g09801(.A(new_n10797_), .B(new_n10796_), .Y(new_n10804_));
  XOR2   g09802(.A(new_n10732_), .B(new_n10725_), .Y(new_n10805_));
  NOR2   g09803(.A(\A[425] ), .B(new_n10729_), .Y(new_n10806_));
  OAI21  g09804(.A0(new_n10727_), .A1(\A[424] ), .B0(\A[426] ), .Y(new_n10807_));
  NAND2  g09805(.A(new_n10731_), .B(new_n10726_), .Y(new_n10808_));
  OAI21  g09806(.A0(new_n10807_), .A1(new_n10806_), .B0(new_n10808_), .Y(new_n10809_));
  NAND2  g09807(.A(new_n10799_), .B(new_n10798_), .Y(new_n10810_));
  NAND2  g09808(.A(new_n10801_), .B(new_n10800_), .Y(new_n10811_));
  NAND4  g09809(.A(new_n10811_), .B(new_n10810_), .C(new_n10809_), .D(new_n10770_), .Y(new_n10812_));
  NAND4  g09810(.A(new_n10789_), .B(new_n10778_), .C(new_n10786_), .D(new_n10783_), .Y(new_n10813_));
  NAND4  g09811(.A(new_n10813_), .B(new_n10775_), .C(new_n10812_), .D(new_n10805_), .Y(new_n10814_));
  OAI211 g09812(.A0(new_n10803_), .A1(new_n10795_), .B0(new_n10814_), .B1(new_n10804_), .Y(new_n10815_));
  XOR2   g09813(.A(new_n10736_), .B(new_n10810_), .Y(new_n10816_));
  XOR2   g09814(.A(new_n10797_), .B(new_n10816_), .Y(new_n10817_));
  NOR4   g09815(.A(new_n10736_), .B(new_n10734_), .C(new_n10732_), .D(new_n10725_), .Y(new_n10818_));
  XOR2   g09816(.A(new_n10751_), .B(new_n10783_), .Y(new_n10819_));
  NOR3   g09817(.A(new_n10819_), .B(new_n10818_), .C(new_n10795_), .Y(new_n10820_));
  AOI221 g09818(.A0(new_n10799_), .A1(new_n10798_), .C0(new_n10735_), .B0(new_n10724_), .B1(\A[423] ), .Y(new_n10821_));
  AOI221 g09819(.A0(new_n10801_), .A1(new_n10800_), .C0(new_n10733_), .B0(new_n10731_), .B1(\A[426] ), .Y(new_n10822_));
  OAI211 g09820(.A0(new_n10822_), .A1(new_n10821_), .B0(new_n10809_), .B1(new_n10770_), .Y(new_n10823_));
  NAND2  g09821(.A(new_n10811_), .B(new_n10810_), .Y(new_n10824_));
  AOI21  g09822(.A0(new_n10824_), .A1(new_n10823_), .B0(new_n10795_), .Y(new_n10825_));
  OAI211 g09823(.A0(new_n10825_), .A1(new_n10817_), .B0(new_n10820_), .B1(new_n10813_), .Y(new_n10826_));
  AOI21  g09824(.A0(new_n10826_), .A1(new_n10815_), .B0(new_n10794_), .Y(new_n10827_));
  OAI21  g09825(.A0(new_n10825_), .A1(new_n10817_), .B0(new_n10814_), .Y(new_n10828_));
  NAND4  g09826(.A(new_n10775_), .B(new_n10804_), .C(new_n10803_), .D(new_n10805_), .Y(new_n10829_));
  OAI21  g09827(.A0(new_n10803_), .A1(new_n10795_), .B0(new_n10813_), .Y(new_n10830_));
  OAI21  g09828(.A0(new_n10830_), .A1(new_n10829_), .B0(new_n10828_), .Y(new_n10831_));
  AOI21  g09829(.A0(new_n10831_), .A1(new_n10794_), .B0(new_n10827_), .Y(new_n10832_));
  OAI21  g09830(.A0(new_n10774_), .A1(new_n10759_), .B0(new_n10832_), .Y(new_n10833_));
  XOR2   g09831(.A(new_n10755_), .B(new_n10753_), .Y(new_n10834_));
  NOR2   g09832(.A(new_n10755_), .B(new_n10753_), .Y(new_n10835_));
  AOI21  g09833(.A0(new_n10792_), .A1(new_n10834_), .B0(new_n10835_), .Y(new_n10836_));
  XOR2   g09834(.A(new_n10792_), .B(new_n10834_), .Y(new_n10837_));
  OAI21  g09835(.A0(new_n10836_), .A1(new_n10819_), .B0(new_n10837_), .Y(new_n10838_));
  OAI21  g09836(.A0(new_n10803_), .A1(new_n10795_), .B0(new_n10804_), .Y(new_n10839_));
  XOR2   g09837(.A(new_n10839_), .B(new_n10814_), .Y(new_n10840_));
  NAND2  g09838(.A(new_n10840_), .B(new_n10838_), .Y(new_n10841_));
  NAND2  g09839(.A(new_n10831_), .B(new_n10794_), .Y(new_n10842_));
  NAND2  g09840(.A(new_n10842_), .B(new_n10841_), .Y(new_n10843_));
  NAND2  g09841(.A(new_n10684_), .B(new_n10634_), .Y(new_n10844_));
  AOI211 g09842(.A0(new_n10668_), .A1(new_n10662_), .B(new_n10688_), .C(new_n10693_), .Y(new_n10845_));
  NOR4   g09843(.A(new_n10845_), .B(new_n10844_), .C(new_n10697_), .D(new_n10690_), .Y(new_n10846_));
  AOI21  g09844(.A0(new_n10760_), .A1(new_n10685_), .B0(new_n10846_), .Y(new_n10847_));
  OAI21  g09845(.A0(new_n10847_), .A1(new_n10710_), .B0(new_n10758_), .Y(new_n10848_));
  OAI21  g09846(.A0(new_n10715_), .A1(new_n10705_), .B0(new_n10773_), .Y(new_n10849_));
  OAI21  g09847(.A0(new_n10848_), .A1(new_n10705_), .B0(new_n10849_), .Y(new_n10850_));
  NAND2  g09848(.A(new_n10850_), .B(new_n10843_), .Y(new_n10851_));
  NAND2  g09849(.A(new_n10851_), .B(new_n10833_), .Y(new_n10852_));
  INV    g09850(.A(\A[440] ), .Y(new_n10853_));
  NOR2   g09851(.A(new_n10853_), .B(\A[439] ), .Y(new_n10854_));
  INV    g09852(.A(\A[439] ), .Y(new_n10855_));
  OAI21  g09853(.A0(\A[440] ), .A1(new_n10855_), .B0(\A[441] ), .Y(new_n10856_));
  XOR2   g09854(.A(\A[440] ), .B(new_n10855_), .Y(new_n10857_));
  OAI22  g09855(.A0(new_n10857_), .A1(\A[441] ), .B0(new_n10856_), .B1(new_n10854_), .Y(new_n10858_));
  INV    g09856(.A(\A[443] ), .Y(new_n10859_));
  NOR2   g09857(.A(new_n10859_), .B(\A[442] ), .Y(new_n10860_));
  INV    g09858(.A(\A[442] ), .Y(new_n10861_));
  OAI21  g09859(.A0(\A[443] ), .A1(new_n10861_), .B0(\A[444] ), .Y(new_n10862_));
  XOR2   g09860(.A(\A[443] ), .B(new_n10861_), .Y(new_n10863_));
  OAI22  g09861(.A0(new_n10863_), .A1(\A[444] ), .B0(new_n10862_), .B1(new_n10860_), .Y(new_n10864_));
  NAND2  g09862(.A(new_n10864_), .B(new_n10858_), .Y(new_n10865_));
  INV    g09863(.A(\A[444] ), .Y(new_n10866_));
  NAND2  g09864(.A(\A[443] ), .B(\A[442] ), .Y(new_n10867_));
  OAI21  g09865(.A0(new_n10863_), .A1(new_n10866_), .B0(new_n10867_), .Y(new_n10868_));
  XOR2   g09866(.A(\A[440] ), .B(\A[439] ), .Y(new_n10869_));
  NOR2   g09867(.A(new_n10853_), .B(new_n10855_), .Y(new_n10870_));
  AOI21  g09868(.A0(new_n10869_), .A1(\A[441] ), .B0(new_n10870_), .Y(new_n10871_));
  XOR2   g09869(.A(new_n10871_), .B(new_n10868_), .Y(new_n10872_));
  XOR2   g09870(.A(new_n10872_), .B(new_n10865_), .Y(new_n10873_));
  NAND2  g09871(.A(\A[443] ), .B(new_n10861_), .Y(new_n10874_));
  AOI21  g09872(.A0(new_n10859_), .A1(\A[442] ), .B0(new_n10866_), .Y(new_n10875_));
  XOR2   g09873(.A(\A[443] ), .B(\A[442] ), .Y(new_n10876_));
  AOI22  g09874(.A0(new_n10876_), .A1(new_n10866_), .B0(new_n10875_), .B1(new_n10874_), .Y(new_n10877_));
  XOR2   g09875(.A(new_n10877_), .B(new_n10858_), .Y(new_n10878_));
  INV    g09876(.A(\A[441] ), .Y(new_n10879_));
  NAND2  g09877(.A(\A[440] ), .B(new_n10855_), .Y(new_n10880_));
  AOI21  g09878(.A0(new_n10853_), .A1(\A[439] ), .B0(new_n10879_), .Y(new_n10881_));
  AOI22  g09879(.A0(new_n10869_), .A1(new_n10879_), .B0(new_n10881_), .B1(new_n10880_), .Y(new_n10882_));
  NOR2   g09880(.A(new_n10877_), .B(new_n10882_), .Y(new_n10883_));
  NOR2   g09881(.A(new_n10859_), .B(new_n10861_), .Y(new_n10884_));
  AOI21  g09882(.A0(new_n10876_), .A1(\A[444] ), .B0(new_n10884_), .Y(new_n10885_));
  XOR2   g09883(.A(new_n10871_), .B(new_n10885_), .Y(new_n10886_));
  NOR2   g09884(.A(new_n10871_), .B(new_n10885_), .Y(new_n10887_));
  AOI21  g09885(.A0(new_n10886_), .A1(new_n10883_), .B0(new_n10887_), .Y(new_n10888_));
  OAI21  g09886(.A0(new_n10888_), .A1(new_n10878_), .B0(new_n10873_), .Y(new_n10889_));
  XOR2   g09887(.A(new_n10877_), .B(new_n10882_), .Y(new_n10890_));
  NAND2  g09888(.A(\A[449] ), .B(\A[448] ), .Y(new_n10891_));
  XOR2   g09889(.A(\A[449] ), .B(\A[448] ), .Y(new_n10892_));
  NAND2  g09890(.A(new_n10892_), .B(\A[450] ), .Y(new_n10893_));
  NAND2  g09891(.A(new_n10893_), .B(new_n10891_), .Y(new_n10894_));
  NAND2  g09892(.A(\A[446] ), .B(\A[445] ), .Y(new_n10895_));
  XOR2   g09893(.A(\A[446] ), .B(\A[445] ), .Y(new_n10896_));
  NAND2  g09894(.A(new_n10896_), .B(\A[447] ), .Y(new_n10897_));
  NAND2  g09895(.A(new_n10897_), .B(new_n10895_), .Y(new_n10898_));
  INV    g09896(.A(\A[446] ), .Y(new_n10899_));
  NOR2   g09897(.A(new_n10899_), .B(\A[445] ), .Y(new_n10900_));
  INV    g09898(.A(\A[445] ), .Y(new_n10901_));
  OAI21  g09899(.A0(\A[446] ), .A1(new_n10901_), .B0(\A[447] ), .Y(new_n10902_));
  INV    g09900(.A(\A[447] ), .Y(new_n10903_));
  NAND2  g09901(.A(new_n10896_), .B(new_n10903_), .Y(new_n10904_));
  OAI21  g09902(.A0(new_n10902_), .A1(new_n10900_), .B0(new_n10904_), .Y(new_n10905_));
  INV    g09903(.A(\A[449] ), .Y(new_n10906_));
  NOR2   g09904(.A(new_n10906_), .B(\A[448] ), .Y(new_n10907_));
  INV    g09905(.A(\A[448] ), .Y(new_n10908_));
  OAI21  g09906(.A0(\A[449] ), .A1(new_n10908_), .B0(\A[450] ), .Y(new_n10909_));
  INV    g09907(.A(\A[450] ), .Y(new_n10910_));
  NAND2  g09908(.A(new_n10892_), .B(new_n10910_), .Y(new_n10911_));
  OAI21  g09909(.A0(new_n10909_), .A1(new_n10907_), .B0(new_n10911_), .Y(new_n10912_));
  NAND4  g09910(.A(new_n10912_), .B(new_n10905_), .C(new_n10898_), .D(new_n10894_), .Y(new_n10913_));
  NAND2  g09911(.A(\A[440] ), .B(\A[439] ), .Y(new_n10914_));
  OAI21  g09912(.A0(new_n10857_), .A1(new_n10879_), .B0(new_n10914_), .Y(new_n10915_));
  NAND4  g09913(.A(new_n10915_), .B(new_n10868_), .C(new_n10864_), .D(new_n10858_), .Y(new_n10916_));
  NAND2  g09914(.A(\A[446] ), .B(new_n10901_), .Y(new_n10917_));
  AOI21  g09915(.A0(new_n10899_), .A1(\A[445] ), .B0(new_n10903_), .Y(new_n10918_));
  AOI22  g09916(.A0(new_n10918_), .A1(new_n10917_), .B0(new_n10896_), .B1(new_n10903_), .Y(new_n10919_));
  NAND2  g09917(.A(\A[449] ), .B(new_n10908_), .Y(new_n10920_));
  AOI21  g09918(.A0(new_n10906_), .A1(\A[448] ), .B0(new_n10910_), .Y(new_n10921_));
  AOI22  g09919(.A0(new_n10921_), .A1(new_n10920_), .B0(new_n10892_), .B1(new_n10910_), .Y(new_n10922_));
  XOR2   g09920(.A(new_n10922_), .B(new_n10919_), .Y(new_n10923_));
  NAND4  g09921(.A(new_n10923_), .B(new_n10916_), .C(new_n10913_), .D(new_n10890_), .Y(new_n10924_));
  XOR2   g09922(.A(new_n10898_), .B(new_n10894_), .Y(new_n10925_));
  NOR2   g09923(.A(new_n10922_), .B(new_n10919_), .Y(new_n10926_));
  AOI22  g09924(.A0(new_n10897_), .A1(new_n10895_), .B0(new_n10893_), .B1(new_n10891_), .Y(new_n10927_));
  AOI21  g09925(.A0(new_n10926_), .A1(new_n10925_), .B0(new_n10927_), .Y(new_n10928_));
  XOR2   g09926(.A(new_n10926_), .B(new_n10925_), .Y(new_n10929_));
  XOR2   g09927(.A(new_n10922_), .B(new_n10905_), .Y(new_n10930_));
  OAI21  g09928(.A0(new_n10930_), .A1(new_n10928_), .B0(new_n10929_), .Y(new_n10931_));
  XOR2   g09929(.A(new_n10931_), .B(new_n10924_), .Y(new_n10932_));
  NAND2  g09930(.A(new_n10912_), .B(new_n10905_), .Y(new_n10933_));
  XOR2   g09931(.A(new_n10933_), .B(new_n10925_), .Y(new_n10934_));
  NOR2   g09932(.A(new_n10899_), .B(new_n10901_), .Y(new_n10935_));
  AOI221 g09933(.A0(new_n10896_), .A1(\A[447] ), .C0(new_n10935_), .B0(new_n10893_), .B1(new_n10891_), .Y(new_n10936_));
  NOR2   g09934(.A(new_n10906_), .B(new_n10908_), .Y(new_n10937_));
  AOI221 g09935(.A0(new_n10897_), .A1(new_n10895_), .C0(new_n10937_), .B0(new_n10892_), .B1(\A[450] ), .Y(new_n10938_));
  OAI211 g09936(.A0(new_n10938_), .A1(new_n10936_), .B0(new_n10912_), .B1(new_n10905_), .Y(new_n10939_));
  NAND2  g09937(.A(new_n10898_), .B(new_n10894_), .Y(new_n10940_));
  AOI21  g09938(.A0(new_n10940_), .A1(new_n10939_), .B0(new_n10930_), .Y(new_n10941_));
  OAI21  g09939(.A0(new_n10941_), .A1(new_n10934_), .B0(new_n10924_), .Y(new_n10942_));
  NOR2   g09940(.A(new_n10930_), .B(new_n10878_), .Y(new_n10943_));
  OAI211 g09941(.A0(new_n10912_), .A1(new_n10905_), .B0(new_n10898_), .B1(new_n10894_), .Y(new_n10944_));
  NAND4  g09942(.A(new_n10944_), .B(new_n10943_), .C(new_n10916_), .D(new_n10929_), .Y(new_n10945_));
  AOI21  g09943(.A0(new_n10945_), .A1(new_n10942_), .B0(new_n10889_), .Y(new_n10946_));
  AOI21  g09944(.A0(new_n10932_), .A1(new_n10889_), .B0(new_n10946_), .Y(new_n10947_));
  INV    g09945(.A(\A[453] ), .Y(new_n10948_));
  INV    g09946(.A(\A[451] ), .Y(new_n10949_));
  NAND2  g09947(.A(\A[452] ), .B(new_n10949_), .Y(new_n10950_));
  INV    g09948(.A(\A[452] ), .Y(new_n10951_));
  AOI21  g09949(.A0(new_n10951_), .A1(\A[451] ), .B0(new_n10948_), .Y(new_n10952_));
  XOR2   g09950(.A(\A[452] ), .B(\A[451] ), .Y(new_n10953_));
  AOI22  g09951(.A0(new_n10953_), .A1(new_n10948_), .B0(new_n10952_), .B1(new_n10950_), .Y(new_n10954_));
  INV    g09952(.A(\A[456] ), .Y(new_n10955_));
  INV    g09953(.A(\A[454] ), .Y(new_n10956_));
  NAND2  g09954(.A(\A[455] ), .B(new_n10956_), .Y(new_n10957_));
  INV    g09955(.A(\A[455] ), .Y(new_n10958_));
  AOI21  g09956(.A0(new_n10958_), .A1(\A[454] ), .B0(new_n10955_), .Y(new_n10959_));
  XOR2   g09957(.A(\A[455] ), .B(\A[454] ), .Y(new_n10960_));
  AOI22  g09958(.A0(new_n10960_), .A1(new_n10955_), .B0(new_n10959_), .B1(new_n10957_), .Y(new_n10961_));
  NOR2   g09959(.A(new_n10961_), .B(new_n10954_), .Y(new_n10962_));
  XOR2   g09960(.A(\A[455] ), .B(new_n10956_), .Y(new_n10963_));
  NAND2  g09961(.A(\A[455] ), .B(\A[454] ), .Y(new_n10964_));
  OAI21  g09962(.A0(new_n10963_), .A1(new_n10955_), .B0(new_n10964_), .Y(new_n10965_));
  NOR2   g09963(.A(new_n10951_), .B(new_n10949_), .Y(new_n10966_));
  AOI21  g09964(.A0(new_n10953_), .A1(\A[453] ), .B0(new_n10966_), .Y(new_n10967_));
  XOR2   g09965(.A(new_n10967_), .B(new_n10965_), .Y(new_n10968_));
  XOR2   g09966(.A(new_n10968_), .B(new_n10962_), .Y(new_n10969_));
  XOR2   g09967(.A(new_n10961_), .B(new_n10954_), .Y(new_n10970_));
  NOR2   g09968(.A(new_n10951_), .B(\A[451] ), .Y(new_n10971_));
  OAI21  g09969(.A0(\A[452] ), .A1(new_n10949_), .B0(\A[453] ), .Y(new_n10972_));
  XOR2   g09970(.A(\A[452] ), .B(new_n10949_), .Y(new_n10973_));
  OAI22  g09971(.A0(new_n10973_), .A1(\A[453] ), .B0(new_n10972_), .B1(new_n10971_), .Y(new_n10974_));
  NOR2   g09972(.A(new_n10958_), .B(\A[454] ), .Y(new_n10975_));
  OAI21  g09973(.A0(\A[455] ), .A1(new_n10956_), .B0(\A[456] ), .Y(new_n10976_));
  OAI22  g09974(.A0(new_n10963_), .A1(\A[456] ), .B0(new_n10976_), .B1(new_n10975_), .Y(new_n10977_));
  NAND2  g09975(.A(new_n10977_), .B(new_n10974_), .Y(new_n10978_));
  NAND2  g09976(.A(\A[452] ), .B(\A[451] ), .Y(new_n10979_));
  OAI21  g09977(.A0(new_n10973_), .A1(new_n10948_), .B0(new_n10979_), .Y(new_n10980_));
  NAND2  g09978(.A(new_n10980_), .B(new_n10965_), .Y(new_n10981_));
  OAI21  g09979(.A0(new_n10968_), .A1(new_n10978_), .B0(new_n10981_), .Y(new_n10982_));
  AOI21  g09980(.A0(new_n10982_), .A1(new_n10970_), .B0(new_n10969_), .Y(new_n10983_));
  NAND2  g09981(.A(\A[461] ), .B(\A[460] ), .Y(new_n10984_));
  XOR2   g09982(.A(\A[461] ), .B(\A[460] ), .Y(new_n10985_));
  NAND2  g09983(.A(new_n10985_), .B(\A[462] ), .Y(new_n10986_));
  NAND2  g09984(.A(new_n10986_), .B(new_n10984_), .Y(new_n10987_));
  NAND2  g09985(.A(\A[458] ), .B(\A[457] ), .Y(new_n10988_));
  XOR2   g09986(.A(\A[458] ), .B(\A[457] ), .Y(new_n10989_));
  NAND2  g09987(.A(new_n10989_), .B(\A[459] ), .Y(new_n10990_));
  NAND2  g09988(.A(new_n10990_), .B(new_n10988_), .Y(new_n10991_));
  XOR2   g09989(.A(new_n10991_), .B(new_n10987_), .Y(new_n10992_));
  INV    g09990(.A(\A[459] ), .Y(new_n10993_));
  INV    g09991(.A(\A[457] ), .Y(new_n10994_));
  NAND2  g09992(.A(\A[458] ), .B(new_n10994_), .Y(new_n10995_));
  INV    g09993(.A(\A[458] ), .Y(new_n10996_));
  AOI21  g09994(.A0(new_n10996_), .A1(\A[457] ), .B0(new_n10993_), .Y(new_n10997_));
  AOI22  g09995(.A0(new_n10997_), .A1(new_n10995_), .B0(new_n10989_), .B1(new_n10993_), .Y(new_n10998_));
  INV    g09996(.A(\A[462] ), .Y(new_n10999_));
  INV    g09997(.A(\A[460] ), .Y(new_n11000_));
  NAND2  g09998(.A(\A[461] ), .B(new_n11000_), .Y(new_n11001_));
  INV    g09999(.A(\A[461] ), .Y(new_n11002_));
  AOI21  g10000(.A0(new_n11002_), .A1(\A[460] ), .B0(new_n10999_), .Y(new_n11003_));
  AOI22  g10001(.A0(new_n11003_), .A1(new_n11001_), .B0(new_n10985_), .B1(new_n10999_), .Y(new_n11004_));
  NOR2   g10002(.A(new_n11004_), .B(new_n10998_), .Y(new_n11005_));
  AOI22  g10003(.A0(new_n10990_), .A1(new_n10988_), .B0(new_n10986_), .B1(new_n10984_), .Y(new_n11006_));
  AOI21  g10004(.A0(new_n11005_), .A1(new_n10992_), .B0(new_n11006_), .Y(new_n11007_));
  XOR2   g10005(.A(new_n11005_), .B(new_n10992_), .Y(new_n11008_));
  NOR2   g10006(.A(new_n10996_), .B(\A[457] ), .Y(new_n11009_));
  OAI21  g10007(.A0(\A[458] ), .A1(new_n10994_), .B0(\A[459] ), .Y(new_n11010_));
  NAND2  g10008(.A(new_n10989_), .B(new_n10993_), .Y(new_n11011_));
  OAI21  g10009(.A0(new_n11010_), .A1(new_n11009_), .B0(new_n11011_), .Y(new_n11012_));
  XOR2   g10010(.A(new_n11004_), .B(new_n11012_), .Y(new_n11013_));
  NOR2   g10011(.A(new_n11002_), .B(\A[460] ), .Y(new_n11014_));
  OAI21  g10012(.A0(\A[461] ), .A1(new_n11000_), .B0(\A[462] ), .Y(new_n11015_));
  NAND2  g10013(.A(new_n10985_), .B(new_n10999_), .Y(new_n11016_));
  OAI21  g10014(.A0(new_n11015_), .A1(new_n11014_), .B0(new_n11016_), .Y(new_n11017_));
  NAND4  g10015(.A(new_n11017_), .B(new_n11012_), .C(new_n10991_), .D(new_n10987_), .Y(new_n11018_));
  NAND4  g10016(.A(new_n10980_), .B(new_n10965_), .C(new_n10977_), .D(new_n10974_), .Y(new_n11019_));
  XOR2   g10017(.A(new_n11004_), .B(new_n10998_), .Y(new_n11020_));
  NAND4  g10018(.A(new_n11020_), .B(new_n11019_), .C(new_n11018_), .D(new_n10970_), .Y(new_n11021_));
  OAI211 g10019(.A0(new_n11013_), .A1(new_n11007_), .B0(new_n11021_), .B1(new_n11008_), .Y(new_n11022_));
  NOR2   g10020(.A(new_n10996_), .B(new_n10994_), .Y(new_n11023_));
  AOI21  g10021(.A0(new_n10989_), .A1(\A[459] ), .B0(new_n11023_), .Y(new_n11024_));
  XOR2   g10022(.A(new_n11024_), .B(new_n10987_), .Y(new_n11025_));
  XOR2   g10023(.A(new_n11005_), .B(new_n11025_), .Y(new_n11026_));
  XOR2   g10024(.A(new_n10961_), .B(new_n10974_), .Y(new_n11027_));
  NOR2   g10025(.A(new_n11002_), .B(new_n11000_), .Y(new_n11028_));
  AOI21  g10026(.A0(new_n10985_), .A1(\A[462] ), .B0(new_n11028_), .Y(new_n11029_));
  NOR4   g10027(.A(new_n11004_), .B(new_n10998_), .C(new_n11024_), .D(new_n11029_), .Y(new_n11030_));
  NOR2   g10028(.A(new_n10958_), .B(new_n10956_), .Y(new_n11031_));
  AOI21  g10029(.A0(new_n10960_), .A1(\A[456] ), .B0(new_n11031_), .Y(new_n11032_));
  NOR4   g10030(.A(new_n10967_), .B(new_n11032_), .C(new_n10961_), .D(new_n10954_), .Y(new_n11033_));
  NOR4   g10031(.A(new_n11013_), .B(new_n11033_), .C(new_n11030_), .D(new_n11027_), .Y(new_n11034_));
  AOI221 g10032(.A0(new_n10989_), .A1(\A[459] ), .C0(new_n11023_), .B0(new_n10986_), .B1(new_n10984_), .Y(new_n11035_));
  AOI221 g10033(.A0(new_n10990_), .A1(new_n10988_), .C0(new_n11028_), .B0(new_n10985_), .B1(\A[462] ), .Y(new_n11036_));
  OAI211 g10034(.A0(new_n11036_), .A1(new_n11035_), .B0(new_n11017_), .B1(new_n11012_), .Y(new_n11037_));
  NAND2  g10035(.A(new_n10991_), .B(new_n10987_), .Y(new_n11038_));
  AOI21  g10036(.A0(new_n11038_), .A1(new_n11037_), .B0(new_n11013_), .Y(new_n11039_));
  OAI21  g10037(.A0(new_n11039_), .A1(new_n11026_), .B0(new_n11034_), .Y(new_n11040_));
  AOI21  g10038(.A0(new_n11040_), .A1(new_n11022_), .B0(new_n10983_), .Y(new_n11041_));
  XOR2   g10039(.A(new_n10968_), .B(new_n10978_), .Y(new_n11042_));
  XOR2   g10040(.A(new_n10967_), .B(new_n11032_), .Y(new_n11043_));
  NOR2   g10041(.A(new_n10967_), .B(new_n11032_), .Y(new_n11044_));
  AOI21  g10042(.A0(new_n11043_), .A1(new_n10962_), .B0(new_n11044_), .Y(new_n11045_));
  OAI21  g10043(.A0(new_n11045_), .A1(new_n11027_), .B0(new_n11042_), .Y(new_n11046_));
  OAI21  g10044(.A0(new_n11039_), .A1(new_n11026_), .B0(new_n11021_), .Y(new_n11047_));
  NOR2   g10045(.A(new_n11013_), .B(new_n11027_), .Y(new_n11048_));
  OAI211 g10046(.A0(new_n11017_), .A1(new_n11012_), .B0(new_n10991_), .B1(new_n10987_), .Y(new_n11049_));
  NAND4  g10047(.A(new_n11049_), .B(new_n11048_), .C(new_n11019_), .D(new_n11008_), .Y(new_n11050_));
  AOI21  g10048(.A0(new_n11050_), .A1(new_n11047_), .B0(new_n11046_), .Y(new_n11051_));
  NOR2   g10049(.A(new_n11013_), .B(new_n11030_), .Y(new_n11052_));
  XOR2   g10050(.A(new_n10961_), .B(new_n10954_), .Y(new_n11053_));
  XOR2   g10051(.A(new_n11053_), .B(new_n11052_), .Y(new_n11054_));
  NAND2  g10052(.A(new_n10923_), .B(new_n10913_), .Y(new_n11055_));
  XOR2   g10053(.A(new_n10877_), .B(new_n10858_), .Y(new_n11056_));
  XOR2   g10054(.A(new_n11056_), .B(new_n11055_), .Y(new_n11057_));
  NAND2  g10055(.A(new_n11057_), .B(new_n11054_), .Y(new_n11058_));
  NOR3   g10056(.A(new_n11058_), .B(new_n11051_), .C(new_n11041_), .Y(new_n11059_));
  OAI21  g10057(.A0(new_n11013_), .A1(new_n11007_), .B0(new_n11008_), .Y(new_n11060_));
  XOR2   g10058(.A(new_n11060_), .B(new_n11021_), .Y(new_n11061_));
  NAND2  g10059(.A(new_n11061_), .B(new_n11046_), .Y(new_n11062_));
  NAND2  g10060(.A(new_n11050_), .B(new_n11047_), .Y(new_n11063_));
  NAND2  g10061(.A(new_n11063_), .B(new_n10983_), .Y(new_n11064_));
  NAND2  g10062(.A(new_n11020_), .B(new_n11018_), .Y(new_n11065_));
  XOR2   g10063(.A(new_n11053_), .B(new_n11065_), .Y(new_n11066_));
  XOR2   g10064(.A(new_n10877_), .B(new_n10882_), .Y(new_n11067_));
  XOR2   g10065(.A(new_n11067_), .B(new_n11055_), .Y(new_n11068_));
  NOR2   g10066(.A(new_n11068_), .B(new_n11066_), .Y(new_n11069_));
  AOI21  g10067(.A0(new_n11064_), .A1(new_n11062_), .B0(new_n11069_), .Y(new_n11070_));
  OAI21  g10068(.A0(new_n11070_), .A1(new_n11059_), .B0(new_n10947_), .Y(new_n11071_));
  XOR2   g10069(.A(new_n10872_), .B(new_n10883_), .Y(new_n11072_));
  NAND2  g10070(.A(new_n10915_), .B(new_n10868_), .Y(new_n11073_));
  OAI21  g10071(.A0(new_n10872_), .A1(new_n10865_), .B0(new_n11073_), .Y(new_n11074_));
  AOI21  g10072(.A0(new_n11074_), .A1(new_n10890_), .B0(new_n11072_), .Y(new_n11075_));
  NOR2   g10073(.A(new_n10941_), .B(new_n10934_), .Y(new_n11076_));
  XOR2   g10074(.A(new_n11076_), .B(new_n10924_), .Y(new_n11077_));
  NAND2  g10075(.A(new_n10945_), .B(new_n10942_), .Y(new_n11078_));
  NAND2  g10076(.A(new_n11078_), .B(new_n11075_), .Y(new_n11079_));
  OAI21  g10077(.A0(new_n11077_), .A1(new_n11075_), .B0(new_n11079_), .Y(new_n11080_));
  NAND2  g10078(.A(new_n11020_), .B(new_n10970_), .Y(new_n11081_));
  AOI211 g10079(.A0(new_n11004_), .A1(new_n10998_), .B(new_n11024_), .C(new_n11029_), .Y(new_n11082_));
  NOR4   g10080(.A(new_n11082_), .B(new_n11081_), .C(new_n11033_), .D(new_n11026_), .Y(new_n11083_));
  AOI21  g10081(.A0(new_n11060_), .A1(new_n11021_), .B0(new_n11083_), .Y(new_n11084_));
  OAI21  g10082(.A0(new_n11084_), .A1(new_n11046_), .B0(new_n11058_), .Y(new_n11085_));
  OAI21  g10083(.A0(new_n11051_), .A1(new_n11041_), .B0(new_n11069_), .Y(new_n11086_));
  OAI21  g10084(.A0(new_n11085_), .A1(new_n11041_), .B0(new_n11086_), .Y(new_n11087_));
  NAND2  g10085(.A(new_n11087_), .B(new_n11080_), .Y(new_n11088_));
  XOR2   g10086(.A(new_n11068_), .B(new_n11054_), .Y(new_n11089_));
  XOR2   g10087(.A(new_n10772_), .B(new_n10718_), .Y(new_n11090_));
  NOR2   g10088(.A(new_n11090_), .B(new_n11089_), .Y(new_n11091_));
  NAND3  g10089(.A(new_n11091_), .B(new_n11088_), .C(new_n11071_), .Y(new_n11092_));
  NAND3  g10090(.A(new_n11069_), .B(new_n11064_), .C(new_n11062_), .Y(new_n11093_));
  OAI21  g10091(.A0(new_n11051_), .A1(new_n11041_), .B0(new_n11058_), .Y(new_n11094_));
  AOI21  g10092(.A0(new_n11094_), .A1(new_n11093_), .B0(new_n11080_), .Y(new_n11095_));
  NAND3  g10093(.A(new_n11058_), .B(new_n11064_), .C(new_n11062_), .Y(new_n11096_));
  AOI21  g10094(.A0(new_n11086_), .A1(new_n11096_), .B0(new_n10947_), .Y(new_n11097_));
  INV    g10095(.A(new_n11091_), .Y(new_n11098_));
  OAI21  g10096(.A0(new_n11097_), .A1(new_n11095_), .B0(new_n11098_), .Y(new_n11099_));
  AOI21  g10097(.A0(new_n11099_), .A1(new_n11092_), .B0(new_n10852_), .Y(new_n11100_));
  NAND3  g10098(.A(new_n10773_), .B(new_n10764_), .C(new_n10762_), .Y(new_n11101_));
  OAI21  g10099(.A0(new_n10715_), .A1(new_n10705_), .B0(new_n10758_), .Y(new_n11102_));
  AOI21  g10100(.A0(new_n11102_), .A1(new_n11101_), .B0(new_n10843_), .Y(new_n11103_));
  AOI21  g10101(.A0(new_n10850_), .A1(new_n10843_), .B0(new_n11103_), .Y(new_n11104_));
  AOI21  g10102(.A0(new_n11087_), .A1(new_n11080_), .B0(new_n11091_), .Y(new_n11105_));
  NAND2  g10103(.A(new_n11105_), .B(new_n11071_), .Y(new_n11106_));
  OAI21  g10104(.A0(new_n11097_), .A1(new_n11095_), .B0(new_n11091_), .Y(new_n11107_));
  AOI21  g10105(.A0(new_n11107_), .A1(new_n11106_), .B0(new_n11104_), .Y(new_n11108_));
  XOR2   g10106(.A(new_n11090_), .B(new_n11089_), .Y(new_n11109_));
  INV    g10107(.A(new_n11109_), .Y(new_n11110_));
  XOR2   g10108(.A(new_n10436_), .B(new_n10356_), .Y(new_n11111_));
  INV    g10109(.A(new_n11111_), .Y(new_n11112_));
  NOR2   g10110(.A(new_n11112_), .B(new_n11110_), .Y(new_n11113_));
  INV    g10111(.A(new_n11113_), .Y(new_n11114_));
  NOR3   g10112(.A(new_n11114_), .B(new_n11108_), .C(new_n11100_), .Y(new_n11115_));
  NOR3   g10113(.A(new_n11098_), .B(new_n11097_), .C(new_n11095_), .Y(new_n11116_));
  AOI21  g10114(.A0(new_n11088_), .A1(new_n11071_), .B0(new_n11091_), .Y(new_n11117_));
  OAI21  g10115(.A0(new_n11117_), .A1(new_n11116_), .B0(new_n11104_), .Y(new_n11118_));
  NOR3   g10116(.A(new_n11091_), .B(new_n11097_), .C(new_n11095_), .Y(new_n11119_));
  AOI21  g10117(.A0(new_n11088_), .A1(new_n11071_), .B0(new_n11098_), .Y(new_n11120_));
  OAI21  g10118(.A0(new_n11120_), .A1(new_n11119_), .B0(new_n10852_), .Y(new_n11121_));
  AOI21  g10119(.A0(new_n11121_), .A1(new_n11118_), .B0(new_n11113_), .Y(new_n11122_));
  OAI21  g10120(.A0(new_n11122_), .A1(new_n11115_), .B0(new_n10611_), .Y(new_n11123_));
  NOR3   g10121(.A(new_n10444_), .B(new_n10443_), .C(new_n10441_), .Y(new_n11124_));
  AOI21  g10122(.A0(new_n10355_), .A1(new_n10341_), .B0(new_n10437_), .Y(new_n11125_));
  OAI21  g10123(.A0(new_n11125_), .A1(new_n11124_), .B0(new_n10606_), .Y(new_n11126_));
  NOR3   g10124(.A(new_n10437_), .B(new_n10443_), .C(new_n10441_), .Y(new_n11127_));
  AOI21  g10125(.A0(new_n10355_), .A1(new_n10341_), .B0(new_n10444_), .Y(new_n11128_));
  OAI21  g10126(.A0(new_n11128_), .A1(new_n11127_), .B0(new_n10586_), .Y(new_n11129_));
  NAND2  g10127(.A(new_n11129_), .B(new_n11126_), .Y(new_n11130_));
  NOR3   g10128(.A(new_n11113_), .B(new_n11108_), .C(new_n11100_), .Y(new_n11131_));
  AOI21  g10129(.A0(new_n11121_), .A1(new_n11118_), .B0(new_n11114_), .Y(new_n11132_));
  OAI21  g10130(.A0(new_n11132_), .A1(new_n11131_), .B0(new_n11130_), .Y(new_n11133_));
  XOR2   g10131(.A(new_n11112_), .B(new_n11109_), .Y(new_n11134_));
  XOR2   g10132(.A(new_n9770_), .B(new_n9607_), .Y(new_n11135_));
  NOR2   g10133(.A(new_n11135_), .B(new_n11134_), .Y(new_n11136_));
  NAND3  g10134(.A(new_n11136_), .B(new_n11133_), .C(new_n11123_), .Y(new_n11137_));
  NAND3  g10135(.A(new_n11113_), .B(new_n11121_), .C(new_n11118_), .Y(new_n11138_));
  OAI21  g10136(.A0(new_n11108_), .A1(new_n11100_), .B0(new_n11114_), .Y(new_n11139_));
  AOI21  g10137(.A0(new_n11139_), .A1(new_n11138_), .B0(new_n11130_), .Y(new_n11140_));
  NAND3  g10138(.A(new_n11114_), .B(new_n11121_), .C(new_n11118_), .Y(new_n11141_));
  OAI21  g10139(.A0(new_n11108_), .A1(new_n11100_), .B0(new_n11113_), .Y(new_n11142_));
  AOI21  g10140(.A0(new_n11142_), .A1(new_n11141_), .B0(new_n10611_), .Y(new_n11143_));
  INV    g10141(.A(new_n11136_), .Y(new_n11144_));
  OAI21  g10142(.A0(new_n11143_), .A1(new_n11140_), .B0(new_n11144_), .Y(new_n11145_));
  AOI21  g10143(.A0(new_n11145_), .A1(new_n11137_), .B0(new_n10122_), .Y(new_n11146_));
  NAND3  g10144(.A(new_n9771_), .B(new_n9779_), .C(new_n9776_), .Y(new_n11147_));
  OAI21  g10145(.A0(new_n9606_), .A1(new_n9598_), .B0(new_n9772_), .Y(new_n11148_));
  AOI21  g10146(.A0(new_n11148_), .A1(new_n11147_), .B0(new_n10118_), .Y(new_n11149_));
  NAND3  g10147(.A(new_n9772_), .B(new_n9779_), .C(new_n9776_), .Y(new_n11150_));
  OAI21  g10148(.A0(new_n9606_), .A1(new_n9598_), .B0(new_n9771_), .Y(new_n11151_));
  AOI21  g10149(.A0(new_n11151_), .A1(new_n11150_), .B0(new_n10110_), .Y(new_n11152_));
  NOR2   g10150(.A(new_n11152_), .B(new_n11149_), .Y(new_n11153_));
  NAND3  g10151(.A(new_n11144_), .B(new_n11133_), .C(new_n11123_), .Y(new_n11154_));
  OAI21  g10152(.A0(new_n11143_), .A1(new_n11140_), .B0(new_n11136_), .Y(new_n11155_));
  AOI21  g10153(.A0(new_n11155_), .A1(new_n11154_), .B0(new_n11153_), .Y(new_n11156_));
  INV    g10154(.A(new_n11135_), .Y(new_n11157_));
  XOR2   g10155(.A(new_n11157_), .B(new_n11134_), .Y(new_n11158_));
  INV    g10156(.A(new_n8070_), .Y(new_n11159_));
  XOR2   g10157(.A(new_n8396_), .B(new_n11159_), .Y(new_n11160_));
  NOR2   g10158(.A(new_n11160_), .B(new_n11158_), .Y(new_n11161_));
  INV    g10159(.A(new_n11161_), .Y(new_n11162_));
  NOR3   g10160(.A(new_n11162_), .B(new_n11156_), .C(new_n11146_), .Y(new_n11163_));
  NOR3   g10161(.A(new_n11144_), .B(new_n11143_), .C(new_n11140_), .Y(new_n11164_));
  AOI21  g10162(.A0(new_n11133_), .A1(new_n11123_), .B0(new_n11136_), .Y(new_n11165_));
  OAI21  g10163(.A0(new_n11165_), .A1(new_n11164_), .B0(new_n11153_), .Y(new_n11166_));
  NOR3   g10164(.A(new_n11136_), .B(new_n11143_), .C(new_n11140_), .Y(new_n11167_));
  AOI21  g10165(.A0(new_n11133_), .A1(new_n11123_), .B0(new_n11144_), .Y(new_n11168_));
  OAI21  g10166(.A0(new_n11168_), .A1(new_n11167_), .B0(new_n10122_), .Y(new_n11169_));
  AOI21  g10167(.A0(new_n11169_), .A1(new_n11166_), .B0(new_n11161_), .Y(new_n11170_));
  OAI21  g10168(.A0(new_n11170_), .A1(new_n11163_), .B0(new_n9109_), .Y(new_n11171_));
  NOR3   g10169(.A(new_n8405_), .B(new_n8404_), .C(new_n8401_), .Y(new_n11172_));
  AOI21  g10170(.A0(new_n8069_), .A1(new_n8059_), .B0(new_n8397_), .Y(new_n11173_));
  OAI21  g10171(.A0(new_n11173_), .A1(new_n11172_), .B0(new_n9105_), .Y(new_n11174_));
  NOR3   g10172(.A(new_n8397_), .B(new_n8404_), .C(new_n8401_), .Y(new_n11175_));
  AOI21  g10173(.A0(new_n8069_), .A1(new_n8059_), .B0(new_n8405_), .Y(new_n11176_));
  OAI21  g10174(.A0(new_n11176_), .A1(new_n11175_), .B0(new_n9097_), .Y(new_n11177_));
  NAND2  g10175(.A(new_n11177_), .B(new_n11174_), .Y(new_n11178_));
  NOR3   g10176(.A(new_n11161_), .B(new_n11156_), .C(new_n11146_), .Y(new_n11179_));
  AOI21  g10177(.A0(new_n11169_), .A1(new_n11166_), .B0(new_n11162_), .Y(new_n11180_));
  OAI21  g10178(.A0(new_n11180_), .A1(new_n11179_), .B0(new_n11178_), .Y(new_n11181_));
  XOR2   g10179(.A(new_n11160_), .B(new_n11158_), .Y(new_n11182_));
  INV    g10180(.A(new_n11182_), .Y(new_n11183_));
  INV    g10181(.A(new_n6437_), .Y(new_n11184_));
  AOI21  g10182(.A0(new_n6110_), .A1(new_n6108_), .B0(new_n11184_), .Y(new_n11185_));
  INV    g10183(.A(new_n11185_), .Y(new_n11186_));
  NAND3  g10184(.A(new_n11184_), .B(new_n6110_), .C(new_n6108_), .Y(new_n11187_));
  AOI21  g10185(.A0(new_n11187_), .A1(new_n11186_), .B0(new_n11183_), .Y(new_n11188_));
  NAND3  g10186(.A(new_n11188_), .B(new_n11181_), .C(new_n11171_), .Y(new_n11189_));
  NAND3  g10187(.A(new_n11161_), .B(new_n11169_), .C(new_n11166_), .Y(new_n11190_));
  OAI21  g10188(.A0(new_n11156_), .A1(new_n11146_), .B0(new_n11162_), .Y(new_n11191_));
  AOI21  g10189(.A0(new_n11191_), .A1(new_n11190_), .B0(new_n11178_), .Y(new_n11192_));
  NAND3  g10190(.A(new_n11162_), .B(new_n11169_), .C(new_n11166_), .Y(new_n11193_));
  OAI21  g10191(.A0(new_n11156_), .A1(new_n11146_), .B0(new_n11161_), .Y(new_n11194_));
  AOI21  g10192(.A0(new_n11194_), .A1(new_n11193_), .B0(new_n9109_), .Y(new_n11195_));
  INV    g10193(.A(new_n11188_), .Y(new_n11196_));
  OAI21  g10194(.A0(new_n11195_), .A1(new_n11192_), .B0(new_n11196_), .Y(new_n11197_));
  AOI21  g10195(.A0(new_n11197_), .A1(new_n11189_), .B0(new_n7058_), .Y(new_n11198_));
  NAND3  g10196(.A(new_n6438_), .B(new_n6446_), .C(new_n6443_), .Y(new_n11199_));
  OAI21  g10197(.A0(new_n6105_), .A1(new_n6096_), .B0(new_n6439_), .Y(new_n11200_));
  AOI21  g10198(.A0(new_n11200_), .A1(new_n11199_), .B0(new_n7054_), .Y(new_n11201_));
  NAND3  g10199(.A(new_n6439_), .B(new_n6446_), .C(new_n6443_), .Y(new_n11202_));
  OAI21  g10200(.A0(new_n6105_), .A1(new_n6096_), .B0(new_n6438_), .Y(new_n11203_));
  AOI21  g10201(.A0(new_n11203_), .A1(new_n11202_), .B0(new_n7041_), .Y(new_n11204_));
  NOR2   g10202(.A(new_n11204_), .B(new_n11201_), .Y(new_n11205_));
  NAND3  g10203(.A(new_n11196_), .B(new_n11181_), .C(new_n11171_), .Y(new_n11206_));
  OAI21  g10204(.A0(new_n11195_), .A1(new_n11192_), .B0(new_n11188_), .Y(new_n11207_));
  AOI21  g10205(.A0(new_n11207_), .A1(new_n11206_), .B0(new_n11205_), .Y(new_n11208_));
  XOR2   g10206(.A(new_n3545_), .B(new_n3544_), .Y(new_n11209_));
  INV    g10207(.A(new_n11187_), .Y(new_n11210_));
  NOR3   g10208(.A(new_n11210_), .B(new_n11185_), .C(new_n11183_), .Y(new_n11211_));
  AOI21  g10209(.A0(new_n11187_), .A1(new_n11186_), .B0(new_n11182_), .Y(new_n11212_));
  NOR2   g10210(.A(new_n11212_), .B(new_n11211_), .Y(new_n11213_));
  NOR2   g10211(.A(new_n11213_), .B(new_n11209_), .Y(new_n11214_));
  NOR3   g10212(.A(new_n11214_), .B(new_n11208_), .C(new_n11198_), .Y(new_n11215_));
  OAI21  g10213(.A0(new_n11208_), .A1(new_n11198_), .B0(new_n11214_), .Y(new_n11216_));
  OAI21  g10214(.A0(new_n11215_), .A1(new_n4771_), .B0(new_n11216_), .Y(new_n11217_));
  NOR3   g10215(.A(new_n11188_), .B(new_n11195_), .C(new_n11192_), .Y(new_n11218_));
  OAI21  g10216(.A0(new_n11218_), .A1(new_n11205_), .B0(new_n11207_), .Y(new_n11219_));
  OAI21  g10217(.A0(new_n7055_), .A1(new_n7041_), .B0(new_n11203_), .Y(new_n11220_));
  AOI21  g10218(.A0(new_n6103_), .A1(new_n5203_), .B0(new_n6445_), .Y(new_n11221_));
  OAI21  g10219(.A0(new_n6080_), .A1(new_n5570_), .B0(new_n6092_), .Y(new_n11222_));
  AOI22  g10220(.A0(new_n5566_), .A1(new_n5422_), .B0(new_n5558_), .B1(new_n5552_), .Y(new_n11223_));
  NOR2   g10221(.A(new_n11223_), .B(new_n6077_), .Y(new_n11224_));
  NAND2  g10222(.A(new_n5561_), .B(new_n5553_), .Y(new_n11225_));
  NOR2   g10223(.A(new_n5542_), .B(new_n5540_), .Y(new_n11226_));
  AOI21  g10224(.A0(new_n5542_), .A1(new_n5540_), .B0(new_n5521_), .Y(new_n11227_));
  NOR2   g10225(.A(new_n5525_), .B(new_n5523_), .Y(new_n11228_));
  AOI21  g10226(.A0(new_n5530_), .A1(new_n5526_), .B0(new_n11228_), .Y(new_n11229_));
  OAI21  g10227(.A0(new_n11227_), .A1(new_n11226_), .B0(new_n11229_), .Y(new_n11230_));
  NAND2  g10228(.A(new_n5533_), .B(new_n5531_), .Y(new_n11231_));
  OAI21  g10229(.A0(new_n5533_), .A1(new_n5531_), .B0(new_n5546_), .Y(new_n11232_));
  INV    g10230(.A(new_n11228_), .Y(new_n11233_));
  OAI21  g10231(.A0(new_n5539_), .A1(new_n5537_), .B0(new_n11233_), .Y(new_n11234_));
  NAND3  g10232(.A(new_n11234_), .B(new_n11232_), .C(new_n11231_), .Y(new_n11235_));
  INV    g10233(.A(new_n5511_), .Y(new_n11236_));
  AOI21  g10234(.A0(new_n5516_), .A1(new_n11236_), .B0(new_n5515_), .Y(new_n11237_));
  NAND3  g10235(.A(new_n11237_), .B(new_n11235_), .C(new_n11230_), .Y(new_n11238_));
  AOI21  g10236(.A0(new_n11232_), .A1(new_n11231_), .B0(new_n11234_), .Y(new_n11239_));
  NOR3   g10237(.A(new_n11229_), .B(new_n11227_), .C(new_n11226_), .Y(new_n11240_));
  INV    g10238(.A(new_n5516_), .Y(new_n11241_));
  OAI21  g10239(.A0(new_n11241_), .A1(new_n5511_), .B0(new_n5518_), .Y(new_n11242_));
  OAI21  g10240(.A0(new_n11240_), .A1(new_n11239_), .B0(new_n11242_), .Y(new_n11243_));
  AOI22  g10241(.A0(new_n11243_), .A1(new_n11238_), .B0(new_n11225_), .B1(new_n5563_), .Y(new_n11244_));
  NOR2   g10242(.A(new_n5554_), .B(new_n5517_), .Y(new_n11245_));
  NOR3   g10243(.A(new_n11242_), .B(new_n11240_), .C(new_n11239_), .Y(new_n11246_));
  AOI21  g10244(.A0(new_n11235_), .A1(new_n11230_), .B0(new_n11237_), .Y(new_n11247_));
  NOR4   g10245(.A(new_n11247_), .B(new_n11246_), .C(new_n11245_), .D(new_n5557_), .Y(new_n11248_));
  NOR2   g10246(.A(new_n11248_), .B(new_n11244_), .Y(new_n11249_));
  AOI21  g10247(.A0(new_n5415_), .A1(new_n5413_), .B0(new_n5409_), .Y(new_n11250_));
  AOI21  g10248(.A0(new_n5506_), .A1(new_n5431_), .B0(new_n11250_), .Y(new_n11251_));
  NAND2  g10249(.A(new_n5291_), .B(new_n5290_), .Y(new_n11252_));
  NAND3  g10250(.A(new_n5294_), .B(new_n5267_), .C(new_n5280_), .Y(new_n11253_));
  AOI211 g10251(.A0(new_n5280_), .A1(new_n11252_), .B(new_n11253_), .C(new_n5292_), .Y(new_n11254_));
  AOI21  g10252(.A0(new_n5282_), .A1(new_n5275_), .B0(new_n5240_), .Y(new_n11255_));
  AOI21  g10253(.A0(new_n5274_), .A1(new_n5280_), .B0(new_n5279_), .Y(new_n11256_));
  OAI21  g10254(.A0(new_n5229_), .A1(new_n5423_), .B0(new_n5425_), .Y(new_n11257_));
  NOR2   g10255(.A(new_n11257_), .B(new_n11256_), .Y(new_n11258_));
  OAI21  g10256(.A0(new_n5281_), .A1(new_n5285_), .B0(new_n11252_), .Y(new_n11259_));
  AOI21  g10257(.A0(new_n5241_), .A1(new_n5224_), .B0(new_n5239_), .Y(new_n11260_));
  NOR2   g10258(.A(new_n11260_), .B(new_n11259_), .Y(new_n11261_));
  OAI22  g10259(.A0(new_n11261_), .A1(new_n11258_), .B0(new_n11255_), .B1(new_n11254_), .Y(new_n11262_));
  NAND2  g10260(.A(new_n5293_), .B(new_n5426_), .Y(new_n11263_));
  NAND2  g10261(.A(new_n11260_), .B(new_n11259_), .Y(new_n11264_));
  NAND2  g10262(.A(new_n11257_), .B(new_n11256_), .Y(new_n11265_));
  NAND4  g10263(.A(new_n11265_), .B(new_n11264_), .C(new_n11263_), .D(new_n5296_), .Y(new_n11266_));
  NAND2  g10264(.A(new_n11266_), .B(new_n11262_), .Y(new_n11267_));
  AOI21  g10265(.A0(new_n5411_), .A1(new_n5372_), .B0(new_n5397_), .Y(new_n11268_));
  AOI21  g10266(.A0(new_n5371_), .A1(new_n5359_), .B0(new_n5358_), .Y(new_n11269_));
  OAI21  g10267(.A0(new_n5378_), .A1(new_n5320_), .B0(new_n5333_), .Y(new_n11270_));
  NOR2   g10268(.A(new_n11270_), .B(new_n11269_), .Y(new_n11271_));
  NAND2  g10269(.A(new_n5389_), .B(new_n5388_), .Y(new_n11272_));
  OAI21  g10270(.A0(new_n5364_), .A1(new_n5377_), .B0(new_n11272_), .Y(new_n11273_));
  AOI21  g10271(.A0(new_n5321_), .A1(new_n5393_), .B0(new_n5396_), .Y(new_n11274_));
  NOR2   g10272(.A(new_n11274_), .B(new_n11273_), .Y(new_n11275_));
  OAI22  g10273(.A0(new_n11275_), .A1(new_n11271_), .B0(new_n11268_), .B1(new_n5434_), .Y(new_n11276_));
  NAND2  g10274(.A(new_n5398_), .B(new_n5334_), .Y(new_n11277_));
  NAND2  g10275(.A(new_n11274_), .B(new_n11273_), .Y(new_n11278_));
  NAND2  g10276(.A(new_n11270_), .B(new_n11269_), .Y(new_n11279_));
  NAND4  g10277(.A(new_n11279_), .B(new_n11278_), .C(new_n11277_), .D(new_n5401_), .Y(new_n11280_));
  NAND2  g10278(.A(new_n11280_), .B(new_n11276_), .Y(new_n11281_));
  XOR2   g10279(.A(new_n11281_), .B(new_n11267_), .Y(new_n11282_));
  XOR2   g10280(.A(new_n11282_), .B(new_n11251_), .Y(new_n11283_));
  XOR2   g10281(.A(new_n11283_), .B(new_n11249_), .Y(new_n11284_));
  XOR2   g10282(.A(new_n11284_), .B(new_n11224_), .Y(new_n11285_));
  AOI22  g10283(.A0(new_n6053_), .A1(new_n6019_), .B0(new_n5799_), .B1(new_n5793_), .Y(new_n11286_));
  NOR2   g10284(.A(new_n11286_), .B(new_n6069_), .Y(new_n11287_));
  OAI21  g10285(.A0(new_n5797_), .A1(new_n5792_), .B0(new_n6050_), .Y(new_n11288_));
  NOR2   g10286(.A(new_n5790_), .B(new_n5789_), .Y(new_n11289_));
  OAI21  g10287(.A0(new_n5762_), .A1(new_n5754_), .B0(new_n5763_), .Y(new_n11290_));
  AOI221 g10288(.A0(new_n11290_), .A1(new_n5773_), .C0(new_n5752_), .B0(new_n5750_), .B1(new_n5734_), .Y(new_n11291_));
  AOI21  g10289(.A0(new_n5763_), .A1(new_n5764_), .B0(new_n5762_), .Y(new_n11292_));
  OAI21  g10290(.A0(new_n5752_), .A1(new_n5778_), .B0(new_n5750_), .Y(new_n11293_));
  NOR2   g10291(.A(new_n11293_), .B(new_n11292_), .Y(new_n11294_));
  NAND2  g10292(.A(new_n5784_), .B(new_n5783_), .Y(new_n11295_));
  OAI21  g10293(.A0(new_n5776_), .A1(new_n5754_), .B0(new_n11295_), .Y(new_n11296_));
  XOR2   g10294(.A(new_n5714_), .B(new_n5712_), .Y(new_n11297_));
  NAND2  g10295(.A(new_n5751_), .B(new_n11297_), .Y(new_n11298_));
  XOR2   g10296(.A(new_n5751_), .B(new_n11297_), .Y(new_n11299_));
  AOI22  g10297(.A0(new_n11299_), .A1(new_n5734_), .B0(new_n5749_), .B1(new_n11298_), .Y(new_n11300_));
  NOR2   g10298(.A(new_n11300_), .B(new_n11296_), .Y(new_n11301_));
  OAI22  g10299(.A0(new_n11301_), .A1(new_n11294_), .B0(new_n11291_), .B1(new_n11289_), .Y(new_n11302_));
  NOR4   g10300(.A(new_n5778_), .B(new_n5776_), .C(new_n11295_), .D(new_n5754_), .Y(new_n11303_));
  OAI211 g10301(.A0(new_n5762_), .A1(new_n5754_), .B0(new_n11303_), .B1(new_n5772_), .Y(new_n11304_));
  OAI21  g10302(.A0(new_n5788_), .A1(new_n5780_), .B0(new_n5753_), .Y(new_n11305_));
  NAND2  g10303(.A(new_n11300_), .B(new_n11296_), .Y(new_n11306_));
  NAND2  g10304(.A(new_n11293_), .B(new_n11292_), .Y(new_n11307_));
  NAND4  g10305(.A(new_n11307_), .B(new_n11306_), .C(new_n11305_), .D(new_n11304_), .Y(new_n11308_));
  NAND2  g10306(.A(new_n11308_), .B(new_n11302_), .Y(new_n11309_));
  NAND2  g10307(.A(new_n5670_), .B(new_n5606_), .Y(new_n11310_));
  NAND2  g10308(.A(new_n5661_), .B(new_n5660_), .Y(new_n11311_));
  OAI21  g10309(.A0(new_n5636_), .A1(new_n5649_), .B0(new_n11311_), .Y(new_n11312_));
  AOI21  g10310(.A0(new_n5593_), .A1(new_n5665_), .B0(new_n5668_), .Y(new_n11313_));
  NAND2  g10311(.A(new_n11313_), .B(new_n11312_), .Y(new_n11314_));
  AOI21  g10312(.A0(new_n5643_), .A1(new_n5631_), .B0(new_n5630_), .Y(new_n11315_));
  OAI21  g10313(.A0(new_n5650_), .A1(new_n5592_), .B0(new_n5605_), .Y(new_n11316_));
  NAND2  g10314(.A(new_n11316_), .B(new_n11315_), .Y(new_n11317_));
  AOI22  g10315(.A0(new_n11317_), .A1(new_n11314_), .B0(new_n11310_), .B1(new_n5673_), .Y(new_n11318_));
  NAND3  g10316(.A(new_n5671_), .B(new_n5642_), .C(new_n5631_), .Y(new_n11319_));
  NOR3   g10317(.A(new_n11319_), .B(new_n5662_), .C(new_n5653_), .Y(new_n11320_));
  AOI21  g10318(.A0(new_n5719_), .A1(new_n5644_), .B0(new_n5669_), .Y(new_n11321_));
  NOR2   g10319(.A(new_n11316_), .B(new_n11315_), .Y(new_n11322_));
  NOR2   g10320(.A(new_n11313_), .B(new_n11312_), .Y(new_n11323_));
  NOR4   g10321(.A(new_n11323_), .B(new_n11322_), .C(new_n11321_), .D(new_n11320_), .Y(new_n11324_));
  NOR2   g10322(.A(new_n11324_), .B(new_n11318_), .Y(new_n11325_));
  XOR2   g10323(.A(new_n11325_), .B(new_n11309_), .Y(new_n11326_));
  XOR2   g10324(.A(new_n11326_), .B(new_n11288_), .Y(new_n11327_));
  NOR3   g10325(.A(new_n6017_), .B(new_n5999_), .C(new_n5989_), .Y(new_n11328_));
  OAI21  g10326(.A0(new_n11328_), .A1(new_n5895_), .B0(new_n6031_), .Y(new_n11329_));
  AOI21  g10327(.A0(new_n5879_), .A1(new_n5872_), .B0(new_n5837_), .Y(new_n11330_));
  AOI21  g10328(.A0(new_n5871_), .A1(new_n5877_), .B0(new_n5876_), .Y(new_n11331_));
  XOR2   g10329(.A(new_n5820_), .B(new_n5831_), .Y(new_n11332_));
  NOR2   g10330(.A(new_n5820_), .B(new_n5813_), .Y(new_n11333_));
  OAI22  g10331(.A0(new_n5835_), .A1(new_n11333_), .B0(new_n5826_), .B1(new_n11332_), .Y(new_n11334_));
  NOR2   g10332(.A(new_n11334_), .B(new_n11331_), .Y(new_n11335_));
  OAI21  g10333(.A0(new_n5878_), .A1(new_n5882_), .B0(new_n6021_), .Y(new_n11336_));
  AOI21  g10334(.A0(new_n5838_), .A1(new_n5821_), .B0(new_n5836_), .Y(new_n11337_));
  NOR2   g10335(.A(new_n11337_), .B(new_n11336_), .Y(new_n11338_));
  OAI22  g10336(.A0(new_n11338_), .A1(new_n11335_), .B0(new_n11330_), .B1(new_n6023_), .Y(new_n11339_));
  OAI211 g10337(.A0(new_n5836_), .A1(new_n5826_), .B0(new_n5890_), .B1(new_n5821_), .Y(new_n11340_));
  NAND2  g10338(.A(new_n11337_), .B(new_n11336_), .Y(new_n11341_));
  NAND2  g10339(.A(new_n11334_), .B(new_n11331_), .Y(new_n11342_));
  NAND4  g10340(.A(new_n11342_), .B(new_n11341_), .C(new_n11340_), .D(new_n5893_), .Y(new_n11343_));
  NAND2  g10341(.A(new_n11343_), .B(new_n11339_), .Y(new_n11344_));
  AOI21  g10342(.A0(new_n6008_), .A1(new_n5969_), .B0(new_n5994_), .Y(new_n11345_));
  AOI21  g10343(.A0(new_n5968_), .A1(new_n5956_), .B0(new_n5955_), .Y(new_n11346_));
  OAI21  g10344(.A0(new_n5975_), .A1(new_n5917_), .B0(new_n5930_), .Y(new_n11347_));
  NOR2   g10345(.A(new_n11347_), .B(new_n11346_), .Y(new_n11348_));
  NAND2  g10346(.A(new_n5986_), .B(new_n5985_), .Y(new_n11349_));
  OAI21  g10347(.A0(new_n5961_), .A1(new_n5974_), .B0(new_n11349_), .Y(new_n11350_));
  AOI21  g10348(.A0(new_n5918_), .A1(new_n5990_), .B0(new_n5993_), .Y(new_n11351_));
  NOR2   g10349(.A(new_n11351_), .B(new_n11350_), .Y(new_n11352_));
  OAI22  g10350(.A0(new_n11352_), .A1(new_n11348_), .B0(new_n11345_), .B1(new_n6028_), .Y(new_n11353_));
  NAND2  g10351(.A(new_n5995_), .B(new_n5931_), .Y(new_n11354_));
  NAND2  g10352(.A(new_n11351_), .B(new_n11350_), .Y(new_n11355_));
  NAND2  g10353(.A(new_n11347_), .B(new_n11346_), .Y(new_n11356_));
  NAND4  g10354(.A(new_n11356_), .B(new_n11355_), .C(new_n11354_), .D(new_n5998_), .Y(new_n11357_));
  NAND2  g10355(.A(new_n11357_), .B(new_n11353_), .Y(new_n11358_));
  XOR2   g10356(.A(new_n11358_), .B(new_n11344_), .Y(new_n11359_));
  XOR2   g10357(.A(new_n11359_), .B(new_n11329_), .Y(new_n11360_));
  XOR2   g10358(.A(new_n11360_), .B(new_n11327_), .Y(new_n11361_));
  XOR2   g10359(.A(new_n11361_), .B(new_n11287_), .Y(new_n11362_));
  XOR2   g10360(.A(new_n11362_), .B(new_n11285_), .Y(new_n11363_));
  NAND2  g10361(.A(new_n11363_), .B(new_n11222_), .Y(new_n11364_));
  OAI21  g10362(.A0(new_n5199_), .A1(new_n5195_), .B0(new_n6100_), .Y(new_n11365_));
  NOR2   g10363(.A(new_n5107_), .B(new_n5083_), .Y(new_n11366_));
  AOI21  g10364(.A0(new_n5120_), .A1(new_n5083_), .B0(new_n11366_), .Y(new_n11367_));
  NOR3   g10365(.A(new_n5188_), .B(new_n5177_), .C(new_n5159_), .Y(new_n11368_));
  OAI22  g10366(.A0(new_n11368_), .A1(new_n11367_), .B0(new_n5192_), .B1(new_n5178_), .Y(new_n11369_));
  XOR2   g10367(.A(new_n5104_), .B(new_n5115_), .Y(new_n11370_));
  NAND4  g10368(.A(new_n5071_), .B(new_n5097_), .C(new_n11370_), .D(new_n5084_), .Y(new_n11371_));
  AOI211 g10369(.A0(new_n5103_), .A1(new_n5084_), .B(new_n11371_), .C(new_n5113_), .Y(new_n11372_));
  OAI21  g10370(.A0(new_n5117_), .A1(new_n5108_), .B0(new_n11370_), .Y(new_n11373_));
  AOI221 g10371(.A0(new_n11373_), .A1(new_n5099_), .C0(new_n5082_), .B0(new_n5080_), .B1(new_n5071_), .Y(new_n11374_));
  XOR2   g10372(.A(new_n5073_), .B(new_n5072_), .Y(new_n11375_));
  AOI21  g10373(.A0(new_n11370_), .A1(new_n5084_), .B0(new_n5117_), .Y(new_n11376_));
  AOI221 g10374(.A0(new_n11375_), .A1(new_n5071_), .C0(new_n11376_), .B0(new_n5079_), .B1(new_n5074_), .Y(new_n11377_));
  OAI21  g10375(.A0(new_n5105_), .A1(new_n5108_), .B0(new_n5103_), .Y(new_n11378_));
  AOI22  g10376(.A0(new_n11375_), .A1(new_n5071_), .B0(new_n5079_), .B1(new_n5074_), .Y(new_n11379_));
  NOR2   g10377(.A(new_n11379_), .B(new_n11378_), .Y(new_n11380_));
  OAI22  g10378(.A0(new_n11380_), .A1(new_n11377_), .B0(new_n11374_), .B1(new_n11372_), .Y(new_n11381_));
  OAI21  g10379(.A0(new_n5106_), .A1(new_n5114_), .B0(new_n5083_), .Y(new_n11382_));
  NAND2  g10380(.A(new_n11379_), .B(new_n11378_), .Y(new_n11383_));
  OAI21  g10381(.A0(new_n5082_), .A1(new_n5112_), .B0(new_n5080_), .Y(new_n11384_));
  NAND2  g10382(.A(new_n11384_), .B(new_n11376_), .Y(new_n11385_));
  NAND4  g10383(.A(new_n11385_), .B(new_n11383_), .C(new_n11382_), .D(new_n5119_), .Y(new_n11386_));
  NAND2  g10384(.A(new_n11386_), .B(new_n11381_), .Y(new_n11387_));
  OAI221 g10385(.A0(new_n5157_), .A1(new_n5181_), .C0(new_n5165_), .B0(new_n5164_), .B1(new_n5162_), .Y(new_n11388_));
  OAI21  g10386(.A0(new_n5156_), .A1(new_n5167_), .B0(new_n5154_), .Y(new_n11389_));
  AOI21  g10387(.A0(new_n5165_), .A1(new_n5123_), .B0(new_n5164_), .Y(new_n11390_));
  NAND2  g10388(.A(new_n11390_), .B(new_n11389_), .Y(new_n11391_));
  AOI21  g10389(.A0(new_n5171_), .A1(new_n5133_), .B0(new_n5170_), .Y(new_n11392_));
  OAI21  g10390(.A0(new_n5131_), .A1(new_n5162_), .B0(new_n5127_), .Y(new_n11393_));
  NAND2  g10391(.A(new_n11393_), .B(new_n11392_), .Y(new_n11394_));
  AOI22  g10392(.A0(new_n11394_), .A1(new_n11391_), .B0(new_n11388_), .B1(new_n5176_), .Y(new_n11395_));
  NOR2   g10393(.A(new_n5185_), .B(new_n5184_), .Y(new_n11396_));
  AOI21  g10394(.A0(new_n5172_), .A1(new_n5150_), .B0(new_n5166_), .Y(new_n11397_));
  AOI211 g10395(.A0(new_n5165_), .A1(new_n5123_), .B(new_n11392_), .C(new_n5164_), .Y(new_n11398_));
  NOR2   g10396(.A(new_n11390_), .B(new_n11389_), .Y(new_n11399_));
  NOR4   g10397(.A(new_n11399_), .B(new_n11398_), .C(new_n11397_), .D(new_n11396_), .Y(new_n11400_));
  NOR2   g10398(.A(new_n11400_), .B(new_n11395_), .Y(new_n11401_));
  XOR2   g10399(.A(new_n11401_), .B(new_n11387_), .Y(new_n11402_));
  XOR2   g10400(.A(new_n11402_), .B(new_n11369_), .Y(new_n11403_));
  AOI21  g10401(.A0(new_n5066_), .A1(new_n4858_), .B0(new_n5061_), .Y(new_n11404_));
  AOI21  g10402(.A0(new_n4854_), .A1(new_n4850_), .B0(new_n4799_), .Y(new_n11405_));
  OAI21  g10403(.A0(new_n4853_), .A1(new_n4841_), .B0(new_n4826_), .Y(new_n11406_));
  XOR2   g10404(.A(new_n4790_), .B(new_n4847_), .Y(new_n11407_));
  XOR2   g10405(.A(new_n11407_), .B(new_n4786_), .Y(new_n11408_));
  NOR3   g10406(.A(new_n11407_), .B(new_n4785_), .C(new_n4778_), .Y(new_n11409_));
  OAI22  g10407(.A0(new_n4797_), .A1(new_n11409_), .B0(new_n4796_), .B1(new_n11408_), .Y(new_n11410_));
  XOR2   g10408(.A(new_n11410_), .B(new_n11406_), .Y(new_n11411_));
  OAI21  g10409(.A0(new_n11405_), .A1(new_n4856_), .B0(new_n11411_), .Y(new_n11412_));
  OAI221 g10410(.A0(new_n4842_), .A1(new_n4840_), .C0(new_n4792_), .B0(new_n4798_), .B1(new_n4796_), .Y(new_n11413_));
  AOI21  g10411(.A0(new_n4837_), .A1(new_n4792_), .B0(new_n4798_), .Y(new_n11414_));
  AOI21  g10412(.A0(new_n11414_), .A1(new_n11406_), .B0(new_n4856_), .Y(new_n11415_));
  OAI211 g10413(.A0(new_n11414_), .A1(new_n11406_), .B0(new_n11415_), .B1(new_n11413_), .Y(new_n11416_));
  NAND2  g10414(.A(new_n11416_), .B(new_n11412_), .Y(new_n11417_));
  NAND3  g10415(.A(new_n4945_), .B(new_n4944_), .C(new_n4942_), .Y(new_n11418_));
  AOI211 g10416(.A0(new_n4928_), .A1(new_n4925_), .B(new_n11418_), .C(new_n4906_), .Y(new_n11419_));
  AOI21  g10417(.A0(new_n4964_), .A1(new_n4959_), .B0(new_n4887_), .Y(new_n11420_));
  AOI21  g10418(.A0(new_n4928_), .A1(new_n4942_), .B0(new_n4963_), .Y(new_n11421_));
  AOI211 g10419(.A0(new_n4937_), .A1(new_n4879_), .B(new_n11421_), .C(new_n4886_), .Y(new_n11422_));
  OAI21  g10420(.A0(new_n4912_), .A1(new_n4927_), .B0(new_n4925_), .Y(new_n11423_));
  AOI21  g10421(.A0(new_n4937_), .A1(new_n4879_), .B0(new_n4886_), .Y(new_n11424_));
  NOR2   g10422(.A(new_n11424_), .B(new_n11423_), .Y(new_n11425_));
  OAI22  g10423(.A0(new_n11425_), .A1(new_n11422_), .B0(new_n11420_), .B1(new_n11419_), .Y(new_n11426_));
  OAI221 g10424(.A0(new_n4929_), .A1(new_n4913_), .C0(new_n4879_), .B0(new_n4886_), .B1(new_n4884_), .Y(new_n11427_));
  NAND2  g10425(.A(new_n11424_), .B(new_n11423_), .Y(new_n11428_));
  OAI21  g10426(.A0(new_n4884_), .A1(new_n4936_), .B0(new_n4939_), .Y(new_n11429_));
  NAND2  g10427(.A(new_n11429_), .B(new_n11421_), .Y(new_n11430_));
  NAND4  g10428(.A(new_n11430_), .B(new_n11428_), .C(new_n11427_), .D(new_n4947_), .Y(new_n11431_));
  NAND2  g10429(.A(new_n11431_), .B(new_n11426_), .Y(new_n11432_));
  XOR2   g10430(.A(new_n11432_), .B(new_n11417_), .Y(new_n11433_));
  XOR2   g10431(.A(new_n11433_), .B(new_n11404_), .Y(new_n11434_));
  XOR2   g10432(.A(new_n11434_), .B(new_n11403_), .Y(new_n11435_));
  XOR2   g10433(.A(new_n11435_), .B(new_n11365_), .Y(new_n11436_));
  AOI21  g10434(.A0(new_n6091_), .A1(new_n6079_), .B0(new_n6081_), .Y(new_n11437_));
  OAI21  g10435(.A0(new_n6068_), .A1(new_n6052_), .B0(new_n6055_), .Y(new_n11438_));
  XOR2   g10436(.A(new_n11361_), .B(new_n11438_), .Y(new_n11439_));
  XOR2   g10437(.A(new_n11439_), .B(new_n11285_), .Y(new_n11440_));
  AOI21  g10438(.A0(new_n11440_), .A1(new_n11437_), .B0(new_n11436_), .Y(new_n11441_));
  XOR2   g10439(.A(new_n11440_), .B(new_n11222_), .Y(new_n11442_));
  AOI22  g10440(.A0(new_n11442_), .A1(new_n11436_), .B0(new_n11441_), .B1(new_n11364_), .Y(new_n11443_));
  NOR2   g10441(.A(new_n11443_), .B(new_n11221_), .Y(new_n11444_));
  AOI21  g10442(.A0(new_n7038_), .A1(new_n7050_), .B0(new_n7052_), .Y(new_n11445_));
  OAI21  g10443(.A0(new_n7047_), .A1(new_n7033_), .B0(new_n7035_), .Y(new_n11446_));
  NOR2   g10444(.A(new_n7012_), .B(new_n6988_), .Y(new_n11447_));
  AOI21  g10445(.A0(new_n7023_), .A1(new_n6988_), .B0(new_n11447_), .Y(new_n11448_));
  NOR3   g10446(.A(new_n6966_), .B(new_n6955_), .C(new_n6938_), .Y(new_n11449_));
  OAI22  g10447(.A0(new_n11449_), .A1(new_n11448_), .B0(new_n7026_), .B1(new_n6956_), .Y(new_n11450_));
  XOR2   g10448(.A(new_n7009_), .B(new_n7018_), .Y(new_n11451_));
  NAND4  g10449(.A(new_n6969_), .B(new_n7002_), .C(new_n11451_), .D(new_n6989_), .Y(new_n11452_));
  AOI211 g10450(.A0(new_n7008_), .A1(new_n6989_), .B(new_n11452_), .C(new_n7016_), .Y(new_n11453_));
  OAI21  g10451(.A0(new_n7020_), .A1(new_n7013_), .B0(new_n11451_), .Y(new_n11454_));
  AOI221 g10452(.A0(new_n11454_), .A1(new_n7004_), .C0(new_n6987_), .B0(new_n6985_), .B1(new_n6969_), .Y(new_n11455_));
  AOI21  g10453(.A0(new_n11451_), .A1(new_n6989_), .B0(new_n7020_), .Y(new_n11456_));
  OAI21  g10454(.A0(new_n6987_), .A1(new_n7015_), .B0(new_n6985_), .Y(new_n11457_));
  NOR2   g10455(.A(new_n11457_), .B(new_n11456_), .Y(new_n11458_));
  OAI21  g10456(.A0(new_n7010_), .A1(new_n7013_), .B0(new_n7008_), .Y(new_n11459_));
  XOR2   g10457(.A(new_n6431_), .B(new_n6429_), .Y(new_n11460_));
  NAND2  g10458(.A(new_n6986_), .B(new_n11460_), .Y(new_n11461_));
  XOR2   g10459(.A(new_n6986_), .B(new_n11460_), .Y(new_n11462_));
  AOI22  g10460(.A0(new_n11462_), .A1(new_n6969_), .B0(new_n6984_), .B1(new_n11461_), .Y(new_n11463_));
  NOR2   g10461(.A(new_n11463_), .B(new_n11459_), .Y(new_n11464_));
  OAI22  g10462(.A0(new_n11464_), .A1(new_n11458_), .B0(new_n11455_), .B1(new_n11453_), .Y(new_n11465_));
  OAI21  g10463(.A0(new_n7011_), .A1(new_n7017_), .B0(new_n6988_), .Y(new_n11466_));
  NAND2  g10464(.A(new_n11463_), .B(new_n11459_), .Y(new_n11467_));
  NAND2  g10465(.A(new_n11457_), .B(new_n11456_), .Y(new_n11468_));
  NAND4  g10466(.A(new_n11468_), .B(new_n11467_), .C(new_n11466_), .D(new_n7022_), .Y(new_n11469_));
  NAND2  g10467(.A(new_n11469_), .B(new_n11465_), .Y(new_n11470_));
  OAI21  g10468(.A0(new_n6936_), .A1(new_n6959_), .B0(new_n6913_), .Y(new_n11471_));
  OAI21  g10469(.A0(new_n6935_), .A1(new_n6945_), .B0(new_n6933_), .Y(new_n11472_));
  AOI21  g10470(.A0(new_n6943_), .A1(new_n6894_), .B0(new_n6942_), .Y(new_n11473_));
  NAND2  g10471(.A(new_n11473_), .B(new_n11472_), .Y(new_n11474_));
  AOI21  g10472(.A0(new_n6949_), .A1(new_n6914_), .B0(new_n6948_), .Y(new_n11475_));
  OAI21  g10473(.A0(new_n6912_), .A1(new_n6939_), .B0(new_n6910_), .Y(new_n11476_));
  NAND2  g10474(.A(new_n11476_), .B(new_n11475_), .Y(new_n11477_));
  AOI22  g10475(.A0(new_n11477_), .A1(new_n11474_), .B0(new_n11471_), .B1(new_n6954_), .Y(new_n11478_));
  NOR2   g10476(.A(new_n6963_), .B(new_n6962_), .Y(new_n11479_));
  AOI21  g10477(.A0(new_n6950_), .A1(new_n6929_), .B0(new_n6944_), .Y(new_n11480_));
  NOR2   g10478(.A(new_n11476_), .B(new_n11475_), .Y(new_n11481_));
  NOR2   g10479(.A(new_n11473_), .B(new_n11472_), .Y(new_n11482_));
  NOR4   g10480(.A(new_n11482_), .B(new_n11481_), .C(new_n11480_), .D(new_n11479_), .Y(new_n11483_));
  NOR2   g10481(.A(new_n11483_), .B(new_n11478_), .Y(new_n11484_));
  XOR2   g10482(.A(new_n11484_), .B(new_n11470_), .Y(new_n11485_));
  XOR2   g10483(.A(new_n11485_), .B(new_n11450_), .Y(new_n11486_));
  OAI21  g10484(.A0(new_n6883_), .A1(new_n6802_), .B0(new_n6890_), .Y(new_n11487_));
  NAND4  g10485(.A(new_n6746_), .B(new_n6779_), .C(new_n6879_), .D(new_n6766_), .Y(new_n11488_));
  AOI211 g10486(.A0(new_n6785_), .A1(new_n6766_), .B(new_n11488_), .C(new_n6794_), .Y(new_n11489_));
  AOI221 g10487(.A0(new_n6880_), .A1(new_n6781_), .C0(new_n6764_), .B0(new_n6762_), .B1(new_n6746_), .Y(new_n11490_));
  AOI21  g10488(.A0(new_n6879_), .A1(new_n6766_), .B0(new_n6798_), .Y(new_n11491_));
  OAI21  g10489(.A0(new_n6764_), .A1(new_n6793_), .B0(new_n6762_), .Y(new_n11492_));
  NOR2   g10490(.A(new_n11492_), .B(new_n11491_), .Y(new_n11493_));
  OAI21  g10491(.A0(new_n6787_), .A1(new_n6791_), .B0(new_n6785_), .Y(new_n11494_));
  XOR2   g10492(.A(new_n6350_), .B(new_n6348_), .Y(new_n11495_));
  NAND2  g10493(.A(new_n6763_), .B(new_n11495_), .Y(new_n11496_));
  XOR2   g10494(.A(new_n6763_), .B(new_n11495_), .Y(new_n11497_));
  AOI22  g10495(.A0(new_n11497_), .A1(new_n6746_), .B0(new_n6761_), .B1(new_n11496_), .Y(new_n11498_));
  NOR2   g10496(.A(new_n11498_), .B(new_n11494_), .Y(new_n11499_));
  OAI22  g10497(.A0(new_n11499_), .A1(new_n11493_), .B0(new_n11490_), .B1(new_n11489_), .Y(new_n11500_));
  OAI21  g10498(.A0(new_n6788_), .A1(new_n6795_), .B0(new_n6765_), .Y(new_n11501_));
  NAND2  g10499(.A(new_n11498_), .B(new_n11494_), .Y(new_n11502_));
  NAND2  g10500(.A(new_n11492_), .B(new_n11491_), .Y(new_n11503_));
  NAND4  g10501(.A(new_n11503_), .B(new_n11502_), .C(new_n11501_), .D(new_n6800_), .Y(new_n11504_));
  NAND2  g10502(.A(new_n11504_), .B(new_n11500_), .Y(new_n11505_));
  OAI21  g10503(.A0(new_n6837_), .A1(new_n6821_), .B0(new_n6854_), .Y(new_n11506_));
  OAI21  g10504(.A0(new_n6836_), .A1(new_n6818_), .B0(new_n6834_), .Y(new_n11507_));
  AOI21  g10505(.A0(new_n6812_), .A1(new_n6840_), .B0(new_n6811_), .Y(new_n11508_));
  NAND2  g10506(.A(new_n11508_), .B(new_n11507_), .Y(new_n11509_));
  AOI21  g10507(.A0(new_n6856_), .A1(new_n6822_), .B0(new_n6860_), .Y(new_n11510_));
  OAI21  g10508(.A0(new_n6853_), .A1(new_n6807_), .B0(new_n6852_), .Y(new_n11511_));
  NAND2  g10509(.A(new_n11511_), .B(new_n11510_), .Y(new_n11512_));
  AOI22  g10510(.A0(new_n11512_), .A1(new_n11509_), .B0(new_n11506_), .B1(new_n6874_), .Y(new_n11513_));
  NOR2   g10511(.A(new_n6862_), .B(new_n6858_), .Y(new_n11514_));
  AOI21  g10512(.A0(new_n6871_), .A1(new_n6868_), .B0(new_n6813_), .Y(new_n11515_));
  NOR2   g10513(.A(new_n11511_), .B(new_n11510_), .Y(new_n11516_));
  NOR2   g10514(.A(new_n11508_), .B(new_n11507_), .Y(new_n11517_));
  NOR4   g10515(.A(new_n11517_), .B(new_n11516_), .C(new_n11515_), .D(new_n11514_), .Y(new_n11518_));
  NOR2   g10516(.A(new_n11518_), .B(new_n11513_), .Y(new_n11519_));
  XOR2   g10517(.A(new_n11519_), .B(new_n11505_), .Y(new_n11520_));
  XOR2   g10518(.A(new_n11520_), .B(new_n11487_), .Y(new_n11521_));
  XOR2   g10519(.A(new_n11521_), .B(new_n11486_), .Y(new_n11522_));
  XOR2   g10520(.A(new_n11522_), .B(new_n11446_), .Y(new_n11523_));
  OAI21  g10521(.A0(new_n6732_), .A1(new_n6581_), .B0(new_n6741_), .Y(new_n11524_));
  AOI21  g10522(.A0(new_n6505_), .A1(new_n6468_), .B0(new_n6493_), .Y(new_n11525_));
  OAI22  g10523(.A0(new_n6728_), .A1(new_n6576_), .B0(new_n11525_), .B1(new_n6448_), .Y(new_n11526_));
  NAND4  g10524(.A(new_n6517_), .B(new_n6541_), .C(new_n6558_), .D(new_n6528_), .Y(new_n11527_));
  AOI221 g10525(.A0(new_n6573_), .A1(new_n6521_), .C0(new_n11527_), .B0(new_n6549_), .B1(new_n6528_), .Y(new_n11528_));
  AOI21  g10526(.A0(new_n6559_), .A1(new_n6545_), .B0(new_n6574_), .Y(new_n11529_));
  AOI21  g10527(.A0(new_n6558_), .A1(new_n6528_), .B0(new_n6557_), .Y(new_n11530_));
  AOI211 g10528(.A0(new_n6573_), .A1(new_n6517_), .B(new_n11530_), .C(new_n6572_), .Y(new_n11531_));
  OAI21  g10529(.A0(new_n6551_), .A1(new_n6554_), .B0(new_n6549_), .Y(new_n11532_));
  AOI21  g10530(.A0(new_n6573_), .A1(new_n6517_), .B0(new_n6572_), .Y(new_n11533_));
  NOR2   g10531(.A(new_n11533_), .B(new_n11532_), .Y(new_n11534_));
  OAI22  g10532(.A0(new_n11534_), .A1(new_n11531_), .B0(new_n11529_), .B1(new_n11528_), .Y(new_n11535_));
  NAND2  g10533(.A(new_n6560_), .B(new_n6527_), .Y(new_n11536_));
  NAND2  g10534(.A(new_n11533_), .B(new_n11532_), .Y(new_n11537_));
  OAI21  g10535(.A0(new_n6526_), .A1(new_n6563_), .B0(new_n6521_), .Y(new_n11538_));
  NAND2  g10536(.A(new_n11538_), .B(new_n11530_), .Y(new_n11539_));
  NAND4  g10537(.A(new_n11539_), .B(new_n11537_), .C(new_n11536_), .D(new_n6565_), .Y(new_n11540_));
  NAND2  g10538(.A(new_n11540_), .B(new_n11535_), .Y(new_n11541_));
  NOR4   g10539(.A(new_n6496_), .B(new_n6495_), .C(new_n6490_), .D(new_n6494_), .Y(new_n11542_));
  OAI211 g10540(.A0(new_n6503_), .A1(new_n6494_), .B0(new_n11542_), .B1(new_n6483_), .Y(new_n11543_));
  OAI21  g10541(.A0(new_n6491_), .A1(new_n6498_), .B0(new_n6468_), .Y(new_n11544_));
  OAI21  g10542(.A0(new_n6490_), .A1(new_n6494_), .B0(new_n6488_), .Y(new_n11545_));
  AOI21  g10543(.A0(new_n6510_), .A1(new_n6449_), .B0(new_n6509_), .Y(new_n11546_));
  NAND2  g10544(.A(new_n11546_), .B(new_n11545_), .Y(new_n11547_));
  AOI21  g10545(.A0(new_n6500_), .A1(new_n6469_), .B0(new_n6503_), .Y(new_n11548_));
  OAI21  g10546(.A0(new_n6467_), .A1(new_n6496_), .B0(new_n6465_), .Y(new_n11549_));
  NAND2  g10547(.A(new_n11549_), .B(new_n11548_), .Y(new_n11550_));
  AOI22  g10548(.A0(new_n11550_), .A1(new_n11547_), .B0(new_n11544_), .B1(new_n11543_), .Y(new_n11551_));
  NOR2   g10549(.A(new_n6504_), .B(new_n6501_), .Y(new_n11552_));
  OAI21  g10550(.A0(new_n6503_), .A1(new_n6494_), .B0(new_n6500_), .Y(new_n11553_));
  AOI21  g10551(.A0(new_n11553_), .A1(new_n6484_), .B0(new_n6511_), .Y(new_n11554_));
  NOR2   g10552(.A(new_n11549_), .B(new_n11548_), .Y(new_n11555_));
  NOR2   g10553(.A(new_n11546_), .B(new_n11545_), .Y(new_n11556_));
  NOR4   g10554(.A(new_n11556_), .B(new_n11555_), .C(new_n11554_), .D(new_n11552_), .Y(new_n11557_));
  NOR2   g10555(.A(new_n11557_), .B(new_n11551_), .Y(new_n11558_));
  XOR2   g10556(.A(new_n11558_), .B(new_n11541_), .Y(new_n11559_));
  XOR2   g10557(.A(new_n11559_), .B(new_n11526_), .Y(new_n11560_));
  OAI22  g10558(.A0(new_n6723_), .A1(new_n6713_), .B0(new_n6720_), .B1(new_n6695_), .Y(new_n11561_));
  NAND4  g10559(.A(new_n6582_), .B(new_n6606_), .C(new_n6623_), .D(new_n6593_), .Y(new_n11562_));
  AOI221 g10560(.A0(new_n6710_), .A1(new_n6586_), .C0(new_n11562_), .B0(new_n6614_), .B1(new_n6593_), .Y(new_n11563_));
  AOI21  g10561(.A0(new_n6624_), .A1(new_n6610_), .B0(new_n6711_), .Y(new_n11564_));
  AOI21  g10562(.A0(new_n6623_), .A1(new_n6593_), .B0(new_n6622_), .Y(new_n11565_));
  AOI211 g10563(.A0(new_n6710_), .A1(new_n6582_), .B(new_n11565_), .C(new_n6709_), .Y(new_n11566_));
  OAI21  g10564(.A0(new_n6616_), .A1(new_n6619_), .B0(new_n6614_), .Y(new_n11567_));
  AOI21  g10565(.A0(new_n6710_), .A1(new_n6582_), .B0(new_n6709_), .Y(new_n11568_));
  NOR2   g10566(.A(new_n11568_), .B(new_n11567_), .Y(new_n11569_));
  OAI22  g10567(.A0(new_n11569_), .A1(new_n11566_), .B0(new_n11564_), .B1(new_n11563_), .Y(new_n11570_));
  NAND2  g10568(.A(new_n6625_), .B(new_n6592_), .Y(new_n11571_));
  NAND2  g10569(.A(new_n11568_), .B(new_n11567_), .Y(new_n11572_));
  OAI21  g10570(.A0(new_n6591_), .A1(new_n6628_), .B0(new_n6586_), .Y(new_n11573_));
  NAND2  g10571(.A(new_n11573_), .B(new_n11565_), .Y(new_n11574_));
  NAND4  g10572(.A(new_n11574_), .B(new_n11572_), .C(new_n11571_), .D(new_n6630_), .Y(new_n11575_));
  NAND2  g10573(.A(new_n11575_), .B(new_n11570_), .Y(new_n11576_));
  NOR4   g10574(.A(new_n6638_), .B(new_n6650_), .C(new_n6667_), .D(new_n6649_), .Y(new_n11577_));
  OAI211 g10575(.A0(new_n6690_), .A1(new_n6649_), .B0(new_n11577_), .B1(new_n6691_), .Y(new_n11578_));
  OAI21  g10576(.A0(new_n6668_), .A1(new_n6652_), .B0(new_n6684_), .Y(new_n11579_));
  OAI21  g10577(.A0(new_n6667_), .A1(new_n6649_), .B0(new_n6665_), .Y(new_n11580_));
  AOI21  g10578(.A0(new_n6643_), .A1(new_n6671_), .B0(new_n6642_), .Y(new_n11581_));
  NAND2  g10579(.A(new_n11581_), .B(new_n11580_), .Y(new_n11582_));
  AOI21  g10580(.A0(new_n6686_), .A1(new_n6653_), .B0(new_n6690_), .Y(new_n11583_));
  OAI21  g10581(.A0(new_n6683_), .A1(new_n6638_), .B0(new_n6682_), .Y(new_n11584_));
  NAND2  g10582(.A(new_n11584_), .B(new_n11583_), .Y(new_n11585_));
  AOI22  g10583(.A0(new_n11585_), .A1(new_n11582_), .B0(new_n11579_), .B1(new_n11578_), .Y(new_n11586_));
  NOR2   g10584(.A(new_n6701_), .B(new_n6644_), .Y(new_n11587_));
  NOR2   g10585(.A(new_n11584_), .B(new_n11583_), .Y(new_n11588_));
  NOR2   g10586(.A(new_n11581_), .B(new_n11580_), .Y(new_n11589_));
  NOR4   g10587(.A(new_n11589_), .B(new_n11588_), .C(new_n11587_), .D(new_n6702_), .Y(new_n11590_));
  NOR2   g10588(.A(new_n11590_), .B(new_n11586_), .Y(new_n11591_));
  XOR2   g10589(.A(new_n11591_), .B(new_n11576_), .Y(new_n11592_));
  XOR2   g10590(.A(new_n11592_), .B(new_n11561_), .Y(new_n11593_));
  XOR2   g10591(.A(new_n11593_), .B(new_n11560_), .Y(new_n11594_));
  XOR2   g10592(.A(new_n11594_), .B(new_n11524_), .Y(new_n11595_));
  XOR2   g10593(.A(new_n11595_), .B(new_n11523_), .Y(new_n11596_));
  XOR2   g10594(.A(new_n11596_), .B(new_n11445_), .Y(new_n11597_));
  OAI21  g10595(.A0(new_n6444_), .A1(new_n6102_), .B0(new_n6104_), .Y(new_n11598_));
  NOR2   g10596(.A(new_n11440_), .B(new_n11437_), .Y(new_n11599_));
  AOI21  g10597(.A0(new_n6099_), .A1(new_n5198_), .B0(new_n5201_), .Y(new_n11600_));
  XOR2   g10598(.A(new_n11435_), .B(new_n11600_), .Y(new_n11601_));
  OAI21  g10599(.A0(new_n11363_), .A1(new_n11222_), .B0(new_n11601_), .Y(new_n11602_));
  XOR2   g10600(.A(new_n11363_), .B(new_n11222_), .Y(new_n11603_));
  OAI22  g10601(.A0(new_n11603_), .A1(new_n11601_), .B0(new_n11602_), .B1(new_n11599_), .Y(new_n11604_));
  OAI21  g10602(.A0(new_n11604_), .A1(new_n11598_), .B0(new_n11597_), .Y(new_n11605_));
  XOR2   g10603(.A(new_n11604_), .B(new_n11598_), .Y(new_n11606_));
  OAI22  g10604(.A0(new_n11606_), .A1(new_n11597_), .B0(new_n11605_), .B1(new_n11444_), .Y(new_n11607_));
  XOR2   g10605(.A(new_n11607_), .B(new_n11220_), .Y(new_n11608_));
  OAI21  g10606(.A0(new_n11179_), .A1(new_n9109_), .B0(new_n11194_), .Y(new_n11609_));
  AOI21  g10607(.A0(new_n9106_), .A1(new_n9097_), .B0(new_n11176_), .Y(new_n11610_));
  OAI21  g10608(.A0(new_n9094_), .A1(new_n9085_), .B0(new_n9103_), .Y(new_n11611_));
  OAI21  g10609(.A0(new_n9090_), .A1(new_n9080_), .B0(new_n9083_), .Y(new_n11612_));
  OAI22  g10610(.A0(new_n9057_), .A1(new_n9052_), .B0(new_n8992_), .B1(new_n8987_), .Y(new_n11613_));
  NOR2   g10611(.A(new_n9050_), .B(new_n9049_), .Y(new_n11614_));
  OAI21  g10612(.A0(new_n9022_), .A1(new_n9014_), .B0(new_n9023_), .Y(new_n11615_));
  AOI221 g10613(.A0(new_n11615_), .A1(new_n9033_), .C0(new_n9012_), .B0(new_n9010_), .B1(new_n8994_), .Y(new_n11616_));
  AOI21  g10614(.A0(new_n9023_), .A1(new_n9024_), .B0(new_n9022_), .Y(new_n11617_));
  OAI21  g10615(.A0(new_n9012_), .A1(new_n9038_), .B0(new_n9010_), .Y(new_n11618_));
  NOR2   g10616(.A(new_n11618_), .B(new_n11617_), .Y(new_n11619_));
  NAND2  g10617(.A(new_n9044_), .B(new_n9043_), .Y(new_n11620_));
  OAI21  g10618(.A0(new_n9036_), .A1(new_n9014_), .B0(new_n11620_), .Y(new_n11621_));
  XOR2   g10619(.A(new_n8391_), .B(new_n8389_), .Y(new_n11622_));
  NAND2  g10620(.A(new_n9011_), .B(new_n11622_), .Y(new_n11623_));
  XOR2   g10621(.A(new_n9011_), .B(new_n11622_), .Y(new_n11624_));
  AOI22  g10622(.A0(new_n11624_), .A1(new_n8994_), .B0(new_n9009_), .B1(new_n11623_), .Y(new_n11625_));
  NOR2   g10623(.A(new_n11625_), .B(new_n11621_), .Y(new_n11626_));
  OAI22  g10624(.A0(new_n11626_), .A1(new_n11619_), .B0(new_n11616_), .B1(new_n11614_), .Y(new_n11627_));
  NOR4   g10625(.A(new_n9038_), .B(new_n9036_), .C(new_n11620_), .D(new_n9014_), .Y(new_n11628_));
  OAI211 g10626(.A0(new_n9022_), .A1(new_n9014_), .B0(new_n11628_), .B1(new_n9032_), .Y(new_n11629_));
  OAI21  g10627(.A0(new_n9048_), .A1(new_n9040_), .B0(new_n9013_), .Y(new_n11630_));
  NAND2  g10628(.A(new_n11625_), .B(new_n11621_), .Y(new_n11631_));
  NAND2  g10629(.A(new_n11618_), .B(new_n11617_), .Y(new_n11632_));
  NAND4  g10630(.A(new_n11632_), .B(new_n11631_), .C(new_n11630_), .D(new_n11629_), .Y(new_n11633_));
  NAND2  g10631(.A(new_n11633_), .B(new_n11627_), .Y(new_n11634_));
  NAND2  g10632(.A(new_n8978_), .B(new_n8939_), .Y(new_n11635_));
  OAI21  g10633(.A0(new_n8966_), .A1(new_n8944_), .B0(new_n9072_), .Y(new_n11636_));
  AOI21  g10634(.A0(new_n9065_), .A1(new_n8920_), .B0(new_n9064_), .Y(new_n11637_));
  NAND2  g10635(.A(new_n11637_), .B(new_n11636_), .Y(new_n11638_));
  AOI21  g10636(.A0(new_n8953_), .A1(new_n8954_), .B0(new_n8952_), .Y(new_n11639_));
  OAI21  g10637(.A0(new_n8938_), .A1(new_n8968_), .B0(new_n8936_), .Y(new_n11640_));
  NAND2  g10638(.A(new_n11640_), .B(new_n11639_), .Y(new_n11641_));
  AOI22  g10639(.A0(new_n11641_), .A1(new_n11638_), .B0(new_n11635_), .B1(new_n9074_), .Y(new_n11642_));
  NOR2   g10640(.A(new_n8980_), .B(new_n8979_), .Y(new_n11643_));
  AOI21  g10641(.A0(new_n9067_), .A1(new_n8963_), .B0(new_n9066_), .Y(new_n11644_));
  NOR2   g10642(.A(new_n11640_), .B(new_n11639_), .Y(new_n11645_));
  NOR2   g10643(.A(new_n11637_), .B(new_n11636_), .Y(new_n11646_));
  NOR4   g10644(.A(new_n11646_), .B(new_n11645_), .C(new_n11644_), .D(new_n11643_), .Y(new_n11647_));
  NOR2   g10645(.A(new_n11647_), .B(new_n11642_), .Y(new_n11648_));
  XOR2   g10646(.A(new_n11648_), .B(new_n11634_), .Y(new_n11649_));
  XOR2   g10647(.A(new_n11649_), .B(new_n11613_), .Y(new_n11650_));
  AOI211 g10648(.A0(new_n8879_), .A1(new_n8837_), .B(new_n8886_), .C(new_n8875_), .Y(new_n11651_));
  OAI22  g10649(.A0(new_n11651_), .A1(new_n8817_), .B0(new_n8887_), .B1(new_n8882_), .Y(new_n11652_));
  NOR2   g10650(.A(new_n8815_), .B(new_n8814_), .Y(new_n11653_));
  OAI21  g10651(.A0(new_n8787_), .A1(new_n8776_), .B0(new_n8788_), .Y(new_n11654_));
  AOI221 g10652(.A0(new_n11654_), .A1(new_n8798_), .C0(new_n8774_), .B0(new_n8772_), .B1(new_n8756_), .Y(new_n11655_));
  AOI21  g10653(.A0(new_n8788_), .A1(new_n8789_), .B0(new_n8787_), .Y(new_n11656_));
  OAI21  g10654(.A0(new_n8774_), .A1(new_n8803_), .B0(new_n8772_), .Y(new_n11657_));
  NOR2   g10655(.A(new_n11657_), .B(new_n11656_), .Y(new_n11658_));
  NAND2  g10656(.A(new_n8809_), .B(new_n8808_), .Y(new_n11659_));
  OAI21  g10657(.A0(new_n8801_), .A1(new_n8776_), .B0(new_n11659_), .Y(new_n11660_));
  XOR2   g10658(.A(new_n8310_), .B(new_n8308_), .Y(new_n11661_));
  NAND2  g10659(.A(new_n8773_), .B(new_n11661_), .Y(new_n11662_));
  XOR2   g10660(.A(new_n8773_), .B(new_n11661_), .Y(new_n11663_));
  AOI22  g10661(.A0(new_n11663_), .A1(new_n8756_), .B0(new_n8771_), .B1(new_n11662_), .Y(new_n11664_));
  NOR2   g10662(.A(new_n11664_), .B(new_n11660_), .Y(new_n11665_));
  OAI22  g10663(.A0(new_n11665_), .A1(new_n11658_), .B0(new_n11655_), .B1(new_n11653_), .Y(new_n11666_));
  NOR4   g10664(.A(new_n8803_), .B(new_n8801_), .C(new_n11659_), .D(new_n8776_), .Y(new_n11667_));
  OAI211 g10665(.A0(new_n8787_), .A1(new_n8776_), .B0(new_n11667_), .B1(new_n8797_), .Y(new_n11668_));
  OAI21  g10666(.A0(new_n8813_), .A1(new_n8805_), .B0(new_n8775_), .Y(new_n11669_));
  NAND2  g10667(.A(new_n11664_), .B(new_n11660_), .Y(new_n11670_));
  NAND2  g10668(.A(new_n11657_), .B(new_n11656_), .Y(new_n11671_));
  NAND4  g10669(.A(new_n11671_), .B(new_n11670_), .C(new_n11669_), .D(new_n11668_), .Y(new_n11672_));
  NAND2  g10670(.A(new_n11672_), .B(new_n11666_), .Y(new_n11673_));
  AOI22  g10671(.A0(new_n8901_), .A1(new_n8900_), .B0(new_n8876_), .B1(new_n8837_), .Y(new_n11674_));
  OAI21  g10672(.A0(new_n8864_), .A1(new_n8842_), .B0(new_n8899_), .Y(new_n11675_));
  AOI21  g10673(.A0(new_n8896_), .A1(new_n8818_), .B0(new_n8895_), .Y(new_n11676_));
  NAND2  g10674(.A(new_n11676_), .B(new_n11675_), .Y(new_n11677_));
  AOI21  g10675(.A0(new_n8851_), .A1(new_n8852_), .B0(new_n8850_), .Y(new_n11678_));
  OAI21  g10676(.A0(new_n8836_), .A1(new_n8866_), .B0(new_n8834_), .Y(new_n11679_));
  NAND2  g10677(.A(new_n11679_), .B(new_n11678_), .Y(new_n11680_));
  AOI21  g10678(.A0(new_n11680_), .A1(new_n11677_), .B0(new_n11674_), .Y(new_n11681_));
  NOR2   g10679(.A(new_n8878_), .B(new_n8877_), .Y(new_n11682_));
  AOI21  g10680(.A0(new_n8898_), .A1(new_n8861_), .B0(new_n8897_), .Y(new_n11683_));
  NOR2   g10681(.A(new_n11679_), .B(new_n11678_), .Y(new_n11684_));
  NOR2   g10682(.A(new_n11676_), .B(new_n11675_), .Y(new_n11685_));
  NOR4   g10683(.A(new_n11685_), .B(new_n11684_), .C(new_n11683_), .D(new_n11682_), .Y(new_n11686_));
  NOR2   g10684(.A(new_n11686_), .B(new_n11681_), .Y(new_n11687_));
  XOR2   g10685(.A(new_n11687_), .B(new_n11673_), .Y(new_n11688_));
  XOR2   g10686(.A(new_n11688_), .B(new_n11652_), .Y(new_n11689_));
  XOR2   g10687(.A(new_n11689_), .B(new_n11650_), .Y(new_n11690_));
  XOR2   g10688(.A(new_n11690_), .B(new_n11612_), .Y(new_n11691_));
  OAI21  g10689(.A0(new_n8752_), .A1(new_n8741_), .B0(new_n8744_), .Y(new_n11692_));
  AOI211 g10690(.A0(new_n8468_), .A1(new_n8426_), .B(new_n8478_), .C(new_n8464_), .Y(new_n11693_));
  OAI22  g10691(.A0(new_n11693_), .A1(new_n8538_), .B0(new_n8479_), .B1(new_n8474_), .Y(new_n11694_));
  NOR2   g10692(.A(new_n8536_), .B(new_n8535_), .Y(new_n11695_));
  AOI21  g10693(.A0(new_n8545_), .A1(new_n8520_), .B0(new_n8544_), .Y(new_n11696_));
  AOI21  g10694(.A0(new_n8510_), .A1(new_n8511_), .B0(new_n8509_), .Y(new_n11697_));
  OAI21  g10695(.A0(new_n8499_), .A1(new_n8525_), .B0(new_n8497_), .Y(new_n11698_));
  NOR2   g10696(.A(new_n11698_), .B(new_n11697_), .Y(new_n11699_));
  NAND2  g10697(.A(new_n8530_), .B(new_n8529_), .Y(new_n11700_));
  OAI21  g10698(.A0(new_n8523_), .A1(new_n8501_), .B0(new_n11700_), .Y(new_n11701_));
  AOI21  g10699(.A0(new_n8543_), .A1(new_n8481_), .B0(new_n8542_), .Y(new_n11702_));
  NOR2   g10700(.A(new_n11702_), .B(new_n11701_), .Y(new_n11703_));
  OAI22  g10701(.A0(new_n11703_), .A1(new_n11699_), .B0(new_n11696_), .B1(new_n11695_), .Y(new_n11704_));
  NOR4   g10702(.A(new_n8525_), .B(new_n8523_), .C(new_n11700_), .D(new_n8501_), .Y(new_n11705_));
  OAI211 g10703(.A0(new_n8509_), .A1(new_n8501_), .B0(new_n11705_), .B1(new_n8519_), .Y(new_n11706_));
  NAND2  g10704(.A(new_n8534_), .B(new_n8500_), .Y(new_n11707_));
  NAND2  g10705(.A(new_n11702_), .B(new_n11701_), .Y(new_n11708_));
  NAND2  g10706(.A(new_n11698_), .B(new_n11697_), .Y(new_n11709_));
  NAND4  g10707(.A(new_n11709_), .B(new_n11708_), .C(new_n11707_), .D(new_n11706_), .Y(new_n11710_));
  NAND2  g10708(.A(new_n11710_), .B(new_n11704_), .Y(new_n11711_));
  AOI22  g10709(.A0(new_n8558_), .A1(new_n8557_), .B0(new_n8465_), .B1(new_n8426_), .Y(new_n11712_));
  OAI21  g10710(.A0(new_n8453_), .A1(new_n8431_), .B0(new_n8556_), .Y(new_n11713_));
  AOI21  g10711(.A0(new_n8553_), .A1(new_n8407_), .B0(new_n8552_), .Y(new_n11714_));
  NAND2  g10712(.A(new_n11714_), .B(new_n11713_), .Y(new_n11715_));
  AOI21  g10713(.A0(new_n8440_), .A1(new_n8441_), .B0(new_n8439_), .Y(new_n11716_));
  OAI21  g10714(.A0(new_n8425_), .A1(new_n8455_), .B0(new_n8423_), .Y(new_n11717_));
  NAND2  g10715(.A(new_n11717_), .B(new_n11716_), .Y(new_n11718_));
  AOI21  g10716(.A0(new_n11718_), .A1(new_n11715_), .B0(new_n11712_), .Y(new_n11719_));
  NOR2   g10717(.A(new_n8467_), .B(new_n8466_), .Y(new_n11720_));
  AOI21  g10718(.A0(new_n8555_), .A1(new_n8450_), .B0(new_n8554_), .Y(new_n11721_));
  NOR2   g10719(.A(new_n11717_), .B(new_n11716_), .Y(new_n11722_));
  NOR2   g10720(.A(new_n11714_), .B(new_n11713_), .Y(new_n11723_));
  NOR4   g10721(.A(new_n11723_), .B(new_n11722_), .C(new_n11721_), .D(new_n11720_), .Y(new_n11724_));
  NOR2   g10722(.A(new_n11724_), .B(new_n11719_), .Y(new_n11725_));
  XOR2   g10723(.A(new_n11725_), .B(new_n11711_), .Y(new_n11726_));
  XOR2   g10724(.A(new_n11726_), .B(new_n11694_), .Y(new_n11727_));
  AOI211 g10725(.A0(new_n8686_), .A1(new_n8644_), .B(new_n8693_), .C(new_n8682_), .Y(new_n11728_));
  OAI22  g10726(.A0(new_n11728_), .A1(new_n8624_), .B0(new_n8694_), .B1(new_n8689_), .Y(new_n11729_));
  NOR2   g10727(.A(new_n8622_), .B(new_n8621_), .Y(new_n11730_));
  AOI21  g10728(.A0(new_n8702_), .A1(new_n8606_), .B0(new_n8701_), .Y(new_n11731_));
  AOI21  g10729(.A0(new_n8596_), .A1(new_n8597_), .B0(new_n8595_), .Y(new_n11732_));
  OAI21  g10730(.A0(new_n8582_), .A1(new_n8611_), .B0(new_n8580_), .Y(new_n11733_));
  NOR2   g10731(.A(new_n11733_), .B(new_n11732_), .Y(new_n11734_));
  NAND2  g10732(.A(new_n8616_), .B(new_n8615_), .Y(new_n11735_));
  OAI21  g10733(.A0(new_n8609_), .A1(new_n8584_), .B0(new_n11735_), .Y(new_n11736_));
  AOI21  g10734(.A0(new_n8700_), .A1(new_n8564_), .B0(new_n8699_), .Y(new_n11737_));
  NOR2   g10735(.A(new_n11737_), .B(new_n11736_), .Y(new_n11738_));
  OAI22  g10736(.A0(new_n11738_), .A1(new_n11734_), .B0(new_n11731_), .B1(new_n11730_), .Y(new_n11739_));
  NOR4   g10737(.A(new_n8611_), .B(new_n8609_), .C(new_n11735_), .D(new_n8584_), .Y(new_n11740_));
  OAI211 g10738(.A0(new_n8595_), .A1(new_n8584_), .B0(new_n11740_), .B1(new_n8605_), .Y(new_n11741_));
  NAND2  g10739(.A(new_n8620_), .B(new_n8583_), .Y(new_n11742_));
  NAND2  g10740(.A(new_n11737_), .B(new_n11736_), .Y(new_n11743_));
  NAND2  g10741(.A(new_n11733_), .B(new_n11732_), .Y(new_n11744_));
  NAND4  g10742(.A(new_n11744_), .B(new_n11743_), .C(new_n11742_), .D(new_n11741_), .Y(new_n11745_));
  NAND2  g10743(.A(new_n11745_), .B(new_n11739_), .Y(new_n11746_));
  AOI22  g10744(.A0(new_n8715_), .A1(new_n8714_), .B0(new_n8683_), .B1(new_n8644_), .Y(new_n11747_));
  OAI21  g10745(.A0(new_n8671_), .A1(new_n8649_), .B0(new_n8713_), .Y(new_n11748_));
  AOI21  g10746(.A0(new_n8710_), .A1(new_n8625_), .B0(new_n8709_), .Y(new_n11749_));
  NAND2  g10747(.A(new_n11749_), .B(new_n11748_), .Y(new_n11750_));
  AOI21  g10748(.A0(new_n8658_), .A1(new_n8659_), .B0(new_n8657_), .Y(new_n11751_));
  OAI21  g10749(.A0(new_n8643_), .A1(new_n8673_), .B0(new_n8641_), .Y(new_n11752_));
  NAND2  g10750(.A(new_n11752_), .B(new_n11751_), .Y(new_n11753_));
  AOI21  g10751(.A0(new_n11753_), .A1(new_n11750_), .B0(new_n11747_), .Y(new_n11754_));
  NOR2   g10752(.A(new_n8685_), .B(new_n8684_), .Y(new_n11755_));
  AOI21  g10753(.A0(new_n8712_), .A1(new_n8668_), .B0(new_n8711_), .Y(new_n11756_));
  NOR2   g10754(.A(new_n11752_), .B(new_n11751_), .Y(new_n11757_));
  NOR2   g10755(.A(new_n11749_), .B(new_n11748_), .Y(new_n11758_));
  NOR4   g10756(.A(new_n11758_), .B(new_n11757_), .C(new_n11756_), .D(new_n11755_), .Y(new_n11759_));
  NOR2   g10757(.A(new_n11759_), .B(new_n11754_), .Y(new_n11760_));
  XOR2   g10758(.A(new_n11760_), .B(new_n11746_), .Y(new_n11761_));
  XOR2   g10759(.A(new_n11761_), .B(new_n11729_), .Y(new_n11762_));
  XOR2   g10760(.A(new_n11762_), .B(new_n11727_), .Y(new_n11763_));
  XOR2   g10761(.A(new_n11763_), .B(new_n11692_), .Y(new_n11764_));
  XOR2   g10762(.A(new_n11764_), .B(new_n11691_), .Y(new_n11765_));
  XOR2   g10763(.A(new_n11765_), .B(new_n11611_), .Y(new_n11766_));
  OAI21  g10764(.A0(new_n8067_), .A1(new_n7547_), .B0(new_n8403_), .Y(new_n11767_));
  OAI21  g10765(.A0(new_n8063_), .A1(new_n7542_), .B0(new_n7545_), .Y(new_n11768_));
  OAI22  g10766(.A0(new_n7519_), .A1(new_n7514_), .B0(new_n7454_), .B1(new_n7449_), .Y(new_n11769_));
  NOR2   g10767(.A(new_n7512_), .B(new_n7511_), .Y(new_n11770_));
  OAI21  g10768(.A0(new_n7484_), .A1(new_n7476_), .B0(new_n7485_), .Y(new_n11771_));
  AOI221 g10769(.A0(new_n11771_), .A1(new_n7495_), .C0(new_n7474_), .B0(new_n7472_), .B1(new_n7456_), .Y(new_n11772_));
  AOI21  g10770(.A0(new_n7485_), .A1(new_n7486_), .B0(new_n7484_), .Y(new_n11773_));
  OAI21  g10771(.A0(new_n7474_), .A1(new_n7500_), .B0(new_n7472_), .Y(new_n11774_));
  NOR2   g10772(.A(new_n11774_), .B(new_n11773_), .Y(new_n11775_));
  NAND2  g10773(.A(new_n7506_), .B(new_n7505_), .Y(new_n11776_));
  OAI21  g10774(.A0(new_n7498_), .A1(new_n7476_), .B0(new_n11776_), .Y(new_n11777_));
  XOR2   g10775(.A(new_n7369_), .B(new_n7367_), .Y(new_n11778_));
  NAND2  g10776(.A(new_n7473_), .B(new_n11778_), .Y(new_n11779_));
  XOR2   g10777(.A(new_n7473_), .B(new_n11778_), .Y(new_n11780_));
  AOI22  g10778(.A0(new_n11780_), .A1(new_n7456_), .B0(new_n7471_), .B1(new_n11779_), .Y(new_n11781_));
  NOR2   g10779(.A(new_n11781_), .B(new_n11777_), .Y(new_n11782_));
  OAI22  g10780(.A0(new_n11782_), .A1(new_n11775_), .B0(new_n11772_), .B1(new_n11770_), .Y(new_n11783_));
  NOR4   g10781(.A(new_n7500_), .B(new_n7498_), .C(new_n11776_), .D(new_n7476_), .Y(new_n11784_));
  OAI211 g10782(.A0(new_n7484_), .A1(new_n7476_), .B0(new_n11784_), .B1(new_n7494_), .Y(new_n11785_));
  OAI21  g10783(.A0(new_n7510_), .A1(new_n7502_), .B0(new_n7475_), .Y(new_n11786_));
  NAND2  g10784(.A(new_n11781_), .B(new_n11777_), .Y(new_n11787_));
  NAND2  g10785(.A(new_n11774_), .B(new_n11773_), .Y(new_n11788_));
  NAND4  g10786(.A(new_n11788_), .B(new_n11787_), .C(new_n11786_), .D(new_n11785_), .Y(new_n11789_));
  NAND2  g10787(.A(new_n11789_), .B(new_n11783_), .Y(new_n11790_));
  NAND2  g10788(.A(new_n7440_), .B(new_n7401_), .Y(new_n11791_));
  OAI21  g10789(.A0(new_n7428_), .A1(new_n7406_), .B0(new_n7534_), .Y(new_n11792_));
  AOI21  g10790(.A0(new_n7527_), .A1(new_n7382_), .B0(new_n7526_), .Y(new_n11793_));
  NAND2  g10791(.A(new_n11793_), .B(new_n11792_), .Y(new_n11794_));
  AOI21  g10792(.A0(new_n7415_), .A1(new_n7416_), .B0(new_n7414_), .Y(new_n11795_));
  OAI21  g10793(.A0(new_n7400_), .A1(new_n7430_), .B0(new_n7398_), .Y(new_n11796_));
  NAND2  g10794(.A(new_n11796_), .B(new_n11795_), .Y(new_n11797_));
  AOI22  g10795(.A0(new_n11797_), .A1(new_n11794_), .B0(new_n11791_), .B1(new_n7536_), .Y(new_n11798_));
  NOR2   g10796(.A(new_n7442_), .B(new_n7441_), .Y(new_n11799_));
  AOI21  g10797(.A0(new_n7529_), .A1(new_n7425_), .B0(new_n7528_), .Y(new_n11800_));
  NOR2   g10798(.A(new_n11796_), .B(new_n11795_), .Y(new_n11801_));
  NOR2   g10799(.A(new_n11793_), .B(new_n11792_), .Y(new_n11802_));
  NOR4   g10800(.A(new_n11802_), .B(new_n11801_), .C(new_n11800_), .D(new_n11799_), .Y(new_n11803_));
  NOR2   g10801(.A(new_n11803_), .B(new_n11798_), .Y(new_n11804_));
  XOR2   g10802(.A(new_n11804_), .B(new_n11790_), .Y(new_n11805_));
  XOR2   g10803(.A(new_n11805_), .B(new_n11769_), .Y(new_n11806_));
  NOR3   g10804(.A(new_n7275_), .B(new_n7257_), .C(new_n7247_), .Y(new_n11807_));
  OAI21  g10805(.A0(new_n11807_), .A1(new_n7153_), .B0(new_n7289_), .Y(new_n11808_));
  AOI21  g10806(.A0(new_n7137_), .A1(new_n7130_), .B0(new_n7095_), .Y(new_n11809_));
  AOI21  g10807(.A0(new_n7129_), .A1(new_n7135_), .B0(new_n7134_), .Y(new_n11810_));
  XOR2   g10808(.A(new_n7078_), .B(new_n7089_), .Y(new_n11811_));
  NOR2   g10809(.A(new_n7078_), .B(new_n7071_), .Y(new_n11812_));
  OAI22  g10810(.A0(new_n7093_), .A1(new_n11812_), .B0(new_n7084_), .B1(new_n11811_), .Y(new_n11813_));
  NOR2   g10811(.A(new_n11813_), .B(new_n11810_), .Y(new_n11814_));
  OAI21  g10812(.A0(new_n7136_), .A1(new_n7140_), .B0(new_n7279_), .Y(new_n11815_));
  AOI21  g10813(.A0(new_n7096_), .A1(new_n7079_), .B0(new_n7094_), .Y(new_n11816_));
  NOR2   g10814(.A(new_n11816_), .B(new_n11815_), .Y(new_n11817_));
  OAI22  g10815(.A0(new_n11817_), .A1(new_n11814_), .B0(new_n11809_), .B1(new_n7281_), .Y(new_n11818_));
  OAI211 g10816(.A0(new_n7094_), .A1(new_n7084_), .B0(new_n7148_), .B1(new_n7079_), .Y(new_n11819_));
  NAND2  g10817(.A(new_n11816_), .B(new_n11815_), .Y(new_n11820_));
  NAND2  g10818(.A(new_n11813_), .B(new_n11810_), .Y(new_n11821_));
  NAND4  g10819(.A(new_n11821_), .B(new_n11820_), .C(new_n11819_), .D(new_n7151_), .Y(new_n11822_));
  NAND2  g10820(.A(new_n11822_), .B(new_n11818_), .Y(new_n11823_));
  AOI21  g10821(.A0(new_n7253_), .A1(new_n7189_), .B0(new_n7286_), .Y(new_n11824_));
  NAND2  g10822(.A(new_n7244_), .B(new_n7243_), .Y(new_n11825_));
  OAI21  g10823(.A0(new_n7219_), .A1(new_n7232_), .B0(new_n11825_), .Y(new_n11826_));
  AOI21  g10824(.A0(new_n7176_), .A1(new_n7248_), .B0(new_n7251_), .Y(new_n11827_));
  NAND2  g10825(.A(new_n11827_), .B(new_n11826_), .Y(new_n11828_));
  AOI21  g10826(.A0(new_n7226_), .A1(new_n7214_), .B0(new_n7213_), .Y(new_n11829_));
  OAI21  g10827(.A0(new_n7233_), .A1(new_n7175_), .B0(new_n7188_), .Y(new_n11830_));
  NAND2  g10828(.A(new_n11830_), .B(new_n11829_), .Y(new_n11831_));
  AOI21  g10829(.A0(new_n11831_), .A1(new_n11828_), .B0(new_n11824_), .Y(new_n11832_));
  AOI21  g10830(.A0(new_n7266_), .A1(new_n7227_), .B0(new_n7252_), .Y(new_n11833_));
  NOR2   g10831(.A(new_n11830_), .B(new_n11829_), .Y(new_n11834_));
  NOR2   g10832(.A(new_n11827_), .B(new_n11826_), .Y(new_n11835_));
  NOR4   g10833(.A(new_n11835_), .B(new_n11834_), .C(new_n11833_), .D(new_n7286_), .Y(new_n11836_));
  NOR2   g10834(.A(new_n11836_), .B(new_n11832_), .Y(new_n11837_));
  XOR2   g10835(.A(new_n11837_), .B(new_n11823_), .Y(new_n11838_));
  XOR2   g10836(.A(new_n11838_), .B(new_n11808_), .Y(new_n11839_));
  XOR2   g10837(.A(new_n11839_), .B(new_n11806_), .Y(new_n11840_));
  XOR2   g10838(.A(new_n11840_), .B(new_n11768_), .Y(new_n11841_));
  AOI22  g10839(.A0(new_n8041_), .A1(new_n8007_), .B0(new_n7787_), .B1(new_n7769_), .Y(new_n11842_));
  NOR2   g10840(.A(new_n11842_), .B(new_n8056_), .Y(new_n11843_));
  NOR3   g10841(.A(new_n7709_), .B(new_n7651_), .C(new_n7641_), .Y(new_n11844_));
  OAI21  g10842(.A0(new_n11844_), .A1(new_n7768_), .B0(new_n7785_), .Y(new_n11845_));
  NOR2   g10843(.A(new_n7766_), .B(new_n7765_), .Y(new_n11846_));
  AOI21  g10844(.A0(new_n7775_), .A1(new_n7750_), .B0(new_n7774_), .Y(new_n11847_));
  AOI21  g10845(.A0(new_n7740_), .A1(new_n7741_), .B0(new_n7739_), .Y(new_n11848_));
  OAI21  g10846(.A0(new_n7729_), .A1(new_n7755_), .B0(new_n7727_), .Y(new_n11849_));
  NOR2   g10847(.A(new_n11849_), .B(new_n11848_), .Y(new_n11850_));
  NAND2  g10848(.A(new_n7760_), .B(new_n7759_), .Y(new_n11851_));
  OAI21  g10849(.A0(new_n7753_), .A1(new_n7731_), .B0(new_n11851_), .Y(new_n11852_));
  AOI21  g10850(.A0(new_n7773_), .A1(new_n7711_), .B0(new_n7772_), .Y(new_n11853_));
  NOR2   g10851(.A(new_n11853_), .B(new_n11852_), .Y(new_n11854_));
  OAI22  g10852(.A0(new_n11854_), .A1(new_n11850_), .B0(new_n11847_), .B1(new_n11846_), .Y(new_n11855_));
  NOR4   g10853(.A(new_n7755_), .B(new_n7753_), .C(new_n11851_), .D(new_n7731_), .Y(new_n11856_));
  OAI211 g10854(.A0(new_n7739_), .A1(new_n7731_), .B0(new_n11856_), .B1(new_n7749_), .Y(new_n11857_));
  NAND2  g10855(.A(new_n7764_), .B(new_n7730_), .Y(new_n11858_));
  NAND2  g10856(.A(new_n11853_), .B(new_n11852_), .Y(new_n11859_));
  NAND2  g10857(.A(new_n11849_), .B(new_n11848_), .Y(new_n11860_));
  NAND4  g10858(.A(new_n11860_), .B(new_n11859_), .C(new_n11858_), .D(new_n11857_), .Y(new_n11861_));
  NAND2  g10859(.A(new_n11861_), .B(new_n11855_), .Y(new_n11862_));
  AOI21  g10860(.A0(new_n7647_), .A1(new_n7583_), .B0(new_n7782_), .Y(new_n11863_));
  NAND2  g10861(.A(new_n7638_), .B(new_n7637_), .Y(new_n11864_));
  OAI21  g10862(.A0(new_n7613_), .A1(new_n7626_), .B0(new_n11864_), .Y(new_n11865_));
  AOI21  g10863(.A0(new_n7570_), .A1(new_n7642_), .B0(new_n7645_), .Y(new_n11866_));
  NAND2  g10864(.A(new_n11866_), .B(new_n11865_), .Y(new_n11867_));
  AOI21  g10865(.A0(new_n7620_), .A1(new_n7608_), .B0(new_n7607_), .Y(new_n11868_));
  OAI21  g10866(.A0(new_n7627_), .A1(new_n7569_), .B0(new_n7582_), .Y(new_n11869_));
  NAND2  g10867(.A(new_n11869_), .B(new_n11868_), .Y(new_n11870_));
  AOI21  g10868(.A0(new_n11870_), .A1(new_n11867_), .B0(new_n11863_), .Y(new_n11871_));
  AOI21  g10869(.A0(new_n7696_), .A1(new_n7621_), .B0(new_n7646_), .Y(new_n11872_));
  NOR2   g10870(.A(new_n11869_), .B(new_n11868_), .Y(new_n11873_));
  NOR2   g10871(.A(new_n11866_), .B(new_n11865_), .Y(new_n11874_));
  NOR4   g10872(.A(new_n11874_), .B(new_n11873_), .C(new_n11872_), .D(new_n7782_), .Y(new_n11875_));
  NOR2   g10873(.A(new_n11875_), .B(new_n11871_), .Y(new_n11876_));
  XOR2   g10874(.A(new_n11876_), .B(new_n11862_), .Y(new_n11877_));
  XOR2   g10875(.A(new_n11877_), .B(new_n11845_), .Y(new_n11878_));
  NOR3   g10876(.A(new_n8005_), .B(new_n7987_), .C(new_n7977_), .Y(new_n11879_));
  OAI21  g10877(.A0(new_n11879_), .A1(new_n7883_), .B0(new_n8022_), .Y(new_n11880_));
  NAND2  g10878(.A(new_n7876_), .B(new_n7875_), .Y(new_n11881_));
  NAND3  g10879(.A(new_n7879_), .B(new_n7852_), .C(new_n7865_), .Y(new_n11882_));
  AOI211 g10880(.A0(new_n7865_), .A1(new_n11881_), .B(new_n11882_), .C(new_n7877_), .Y(new_n11883_));
  AOI21  g10881(.A0(new_n7867_), .A1(new_n7860_), .B0(new_n7825_), .Y(new_n11884_));
  AOI21  g10882(.A0(new_n7859_), .A1(new_n7865_), .B0(new_n7864_), .Y(new_n11885_));
  OAI21  g10883(.A0(new_n7814_), .A1(new_n8008_), .B0(new_n8010_), .Y(new_n11886_));
  NOR2   g10884(.A(new_n11886_), .B(new_n11885_), .Y(new_n11887_));
  OAI21  g10885(.A0(new_n7866_), .A1(new_n7870_), .B0(new_n11881_), .Y(new_n11888_));
  AOI21  g10886(.A0(new_n7826_), .A1(new_n7809_), .B0(new_n7824_), .Y(new_n11889_));
  NOR2   g10887(.A(new_n11889_), .B(new_n11888_), .Y(new_n11890_));
  OAI22  g10888(.A0(new_n11890_), .A1(new_n11887_), .B0(new_n11884_), .B1(new_n11883_), .Y(new_n11891_));
  NAND2  g10889(.A(new_n7878_), .B(new_n8011_), .Y(new_n11892_));
  NAND2  g10890(.A(new_n11889_), .B(new_n11888_), .Y(new_n11893_));
  NAND2  g10891(.A(new_n11886_), .B(new_n11885_), .Y(new_n11894_));
  NAND4  g10892(.A(new_n11894_), .B(new_n11893_), .C(new_n11892_), .D(new_n7881_), .Y(new_n11895_));
  NAND2  g10893(.A(new_n11895_), .B(new_n11891_), .Y(new_n11896_));
  AOI21  g10894(.A0(new_n7996_), .A1(new_n7957_), .B0(new_n7982_), .Y(new_n11897_));
  AOI21  g10895(.A0(new_n7956_), .A1(new_n7944_), .B0(new_n7943_), .Y(new_n11898_));
  OAI21  g10896(.A0(new_n7963_), .A1(new_n7905_), .B0(new_n7918_), .Y(new_n11899_));
  NOR2   g10897(.A(new_n11899_), .B(new_n11898_), .Y(new_n11900_));
  NAND2  g10898(.A(new_n7974_), .B(new_n7973_), .Y(new_n11901_));
  OAI21  g10899(.A0(new_n7949_), .A1(new_n7962_), .B0(new_n11901_), .Y(new_n11902_));
  AOI21  g10900(.A0(new_n7906_), .A1(new_n7978_), .B0(new_n7981_), .Y(new_n11903_));
  NOR2   g10901(.A(new_n11903_), .B(new_n11902_), .Y(new_n11904_));
  OAI22  g10902(.A0(new_n11904_), .A1(new_n11900_), .B0(new_n11897_), .B1(new_n8019_), .Y(new_n11905_));
  NAND2  g10903(.A(new_n7983_), .B(new_n7919_), .Y(new_n11906_));
  NAND2  g10904(.A(new_n11903_), .B(new_n11902_), .Y(new_n11907_));
  NAND2  g10905(.A(new_n11899_), .B(new_n11898_), .Y(new_n11908_));
  NAND4  g10906(.A(new_n11908_), .B(new_n11907_), .C(new_n11906_), .D(new_n7986_), .Y(new_n11909_));
  NAND2  g10907(.A(new_n11909_), .B(new_n11905_), .Y(new_n11910_));
  XOR2   g10908(.A(new_n11910_), .B(new_n11896_), .Y(new_n11911_));
  XOR2   g10909(.A(new_n11911_), .B(new_n11880_), .Y(new_n11912_));
  XOR2   g10910(.A(new_n11912_), .B(new_n11878_), .Y(new_n11913_));
  XOR2   g10911(.A(new_n11913_), .B(new_n11843_), .Y(new_n11914_));
  XOR2   g10912(.A(new_n11914_), .B(new_n11841_), .Y(new_n11915_));
  XOR2   g10913(.A(new_n11915_), .B(new_n11767_), .Y(new_n11916_));
  XOR2   g10914(.A(new_n11916_), .B(new_n11766_), .Y(new_n11917_));
  XOR2   g10915(.A(new_n11917_), .B(new_n11610_), .Y(new_n11918_));
  OAI21  g10916(.A0(new_n11167_), .A1(new_n11153_), .B0(new_n11155_), .Y(new_n11919_));
  OAI21  g10917(.A0(new_n10119_), .A1(new_n10110_), .B0(new_n11151_), .Y(new_n11920_));
  OAI21  g10918(.A0(new_n10115_), .A1(new_n10105_), .B0(new_n10108_), .Y(new_n11921_));
  OAI22  g10919(.A0(new_n10082_), .A1(new_n10077_), .B0(new_n10017_), .B1(new_n10012_), .Y(new_n11922_));
  NOR2   g10920(.A(new_n10075_), .B(new_n10074_), .Y(new_n11923_));
  OAI21  g10921(.A0(new_n10047_), .A1(new_n10039_), .B0(new_n10048_), .Y(new_n11924_));
  AOI221 g10922(.A0(new_n11924_), .A1(new_n10058_), .C0(new_n10037_), .B0(new_n10035_), .B1(new_n10019_), .Y(new_n11925_));
  AOI21  g10923(.A0(new_n10048_), .A1(new_n10049_), .B0(new_n10047_), .Y(new_n11926_));
  OAI21  g10924(.A0(new_n10037_), .A1(new_n10063_), .B0(new_n10035_), .Y(new_n11927_));
  NOR2   g10925(.A(new_n11927_), .B(new_n11926_), .Y(new_n11928_));
  NAND2  g10926(.A(new_n10069_), .B(new_n10068_), .Y(new_n11929_));
  OAI21  g10927(.A0(new_n10061_), .A1(new_n10039_), .B0(new_n11929_), .Y(new_n11930_));
  XOR2   g10928(.A(new_n9766_), .B(new_n9764_), .Y(new_n11931_));
  NAND2  g10929(.A(new_n10036_), .B(new_n11931_), .Y(new_n11932_));
  XOR2   g10930(.A(new_n10036_), .B(new_n11931_), .Y(new_n11933_));
  AOI22  g10931(.A0(new_n11933_), .A1(new_n10019_), .B0(new_n10034_), .B1(new_n11932_), .Y(new_n11934_));
  NOR2   g10932(.A(new_n11934_), .B(new_n11930_), .Y(new_n11935_));
  OAI22  g10933(.A0(new_n11935_), .A1(new_n11928_), .B0(new_n11925_), .B1(new_n11923_), .Y(new_n11936_));
  NOR4   g10934(.A(new_n10063_), .B(new_n10061_), .C(new_n11929_), .D(new_n10039_), .Y(new_n11937_));
  OAI211 g10935(.A0(new_n10047_), .A1(new_n10039_), .B0(new_n11937_), .B1(new_n10057_), .Y(new_n11938_));
  OAI21  g10936(.A0(new_n10073_), .A1(new_n10065_), .B0(new_n10038_), .Y(new_n11939_));
  NAND2  g10937(.A(new_n11934_), .B(new_n11930_), .Y(new_n11940_));
  NAND2  g10938(.A(new_n11927_), .B(new_n11926_), .Y(new_n11941_));
  NAND4  g10939(.A(new_n11941_), .B(new_n11940_), .C(new_n11939_), .D(new_n11938_), .Y(new_n11942_));
  NAND2  g10940(.A(new_n11942_), .B(new_n11936_), .Y(new_n11943_));
  NAND2  g10941(.A(new_n10003_), .B(new_n9964_), .Y(new_n11944_));
  OAI21  g10942(.A0(new_n9991_), .A1(new_n9969_), .B0(new_n10097_), .Y(new_n11945_));
  AOI21  g10943(.A0(new_n10090_), .A1(new_n9945_), .B0(new_n10089_), .Y(new_n11946_));
  NAND2  g10944(.A(new_n11946_), .B(new_n11945_), .Y(new_n11947_));
  AOI21  g10945(.A0(new_n9978_), .A1(new_n9979_), .B0(new_n9977_), .Y(new_n11948_));
  OAI21  g10946(.A0(new_n9963_), .A1(new_n9993_), .B0(new_n9961_), .Y(new_n11949_));
  NAND2  g10947(.A(new_n11949_), .B(new_n11948_), .Y(new_n11950_));
  AOI22  g10948(.A0(new_n11950_), .A1(new_n11947_), .B0(new_n11944_), .B1(new_n10099_), .Y(new_n11951_));
  NOR2   g10949(.A(new_n10005_), .B(new_n10004_), .Y(new_n11952_));
  AOI21  g10950(.A0(new_n10092_), .A1(new_n9988_), .B0(new_n10091_), .Y(new_n11953_));
  NOR2   g10951(.A(new_n11949_), .B(new_n11948_), .Y(new_n11954_));
  NOR2   g10952(.A(new_n11946_), .B(new_n11945_), .Y(new_n11955_));
  NOR4   g10953(.A(new_n11955_), .B(new_n11954_), .C(new_n11953_), .D(new_n11952_), .Y(new_n11956_));
  NOR2   g10954(.A(new_n11956_), .B(new_n11951_), .Y(new_n11957_));
  XOR2   g10955(.A(new_n11957_), .B(new_n11943_), .Y(new_n11958_));
  XOR2   g10956(.A(new_n11958_), .B(new_n11922_), .Y(new_n11959_));
  AOI211 g10957(.A0(new_n9904_), .A1(new_n9862_), .B(new_n9911_), .C(new_n9900_), .Y(new_n11960_));
  OAI22  g10958(.A0(new_n11960_), .A1(new_n9842_), .B0(new_n9912_), .B1(new_n9907_), .Y(new_n11961_));
  NOR2   g10959(.A(new_n9840_), .B(new_n9839_), .Y(new_n11962_));
  OAI21  g10960(.A0(new_n9812_), .A1(new_n9801_), .B0(new_n9813_), .Y(new_n11963_));
  AOI221 g10961(.A0(new_n11963_), .A1(new_n9823_), .C0(new_n9799_), .B0(new_n9797_), .B1(new_n9781_), .Y(new_n11964_));
  AOI21  g10962(.A0(new_n9813_), .A1(new_n9814_), .B0(new_n9812_), .Y(new_n11965_));
  OAI21  g10963(.A0(new_n9799_), .A1(new_n9828_), .B0(new_n9797_), .Y(new_n11966_));
  NOR2   g10964(.A(new_n11966_), .B(new_n11965_), .Y(new_n11967_));
  NAND2  g10965(.A(new_n9834_), .B(new_n9833_), .Y(new_n11968_));
  OAI21  g10966(.A0(new_n9826_), .A1(new_n9801_), .B0(new_n11968_), .Y(new_n11969_));
  XOR2   g10967(.A(new_n9685_), .B(new_n9683_), .Y(new_n11970_));
  NAND2  g10968(.A(new_n9798_), .B(new_n11970_), .Y(new_n11971_));
  XOR2   g10969(.A(new_n9798_), .B(new_n11970_), .Y(new_n11972_));
  AOI22  g10970(.A0(new_n11972_), .A1(new_n9781_), .B0(new_n9796_), .B1(new_n11971_), .Y(new_n11973_));
  NOR2   g10971(.A(new_n11973_), .B(new_n11969_), .Y(new_n11974_));
  OAI22  g10972(.A0(new_n11974_), .A1(new_n11967_), .B0(new_n11964_), .B1(new_n11962_), .Y(new_n11975_));
  NOR4   g10973(.A(new_n9828_), .B(new_n9826_), .C(new_n11968_), .D(new_n9801_), .Y(new_n11976_));
  OAI211 g10974(.A0(new_n9812_), .A1(new_n9801_), .B0(new_n11976_), .B1(new_n9822_), .Y(new_n11977_));
  OAI21  g10975(.A0(new_n9838_), .A1(new_n9830_), .B0(new_n9800_), .Y(new_n11978_));
  NAND2  g10976(.A(new_n11973_), .B(new_n11969_), .Y(new_n11979_));
  NAND2  g10977(.A(new_n11966_), .B(new_n11965_), .Y(new_n11980_));
  NAND4  g10978(.A(new_n11980_), .B(new_n11979_), .C(new_n11978_), .D(new_n11977_), .Y(new_n11981_));
  NAND2  g10979(.A(new_n11981_), .B(new_n11975_), .Y(new_n11982_));
  AOI22  g10980(.A0(new_n9926_), .A1(new_n9925_), .B0(new_n9901_), .B1(new_n9862_), .Y(new_n11983_));
  OAI21  g10981(.A0(new_n9889_), .A1(new_n9867_), .B0(new_n9924_), .Y(new_n11984_));
  AOI21  g10982(.A0(new_n9921_), .A1(new_n9843_), .B0(new_n9920_), .Y(new_n11985_));
  NAND2  g10983(.A(new_n11985_), .B(new_n11984_), .Y(new_n11986_));
  AOI21  g10984(.A0(new_n9876_), .A1(new_n9877_), .B0(new_n9875_), .Y(new_n11987_));
  OAI21  g10985(.A0(new_n9861_), .A1(new_n9891_), .B0(new_n9859_), .Y(new_n11988_));
  NAND2  g10986(.A(new_n11988_), .B(new_n11987_), .Y(new_n11989_));
  AOI21  g10987(.A0(new_n11989_), .A1(new_n11986_), .B0(new_n11983_), .Y(new_n11990_));
  NOR2   g10988(.A(new_n9903_), .B(new_n9902_), .Y(new_n11991_));
  AOI21  g10989(.A0(new_n9923_), .A1(new_n9886_), .B0(new_n9922_), .Y(new_n11992_));
  NOR2   g10990(.A(new_n11988_), .B(new_n11987_), .Y(new_n11993_));
  NOR2   g10991(.A(new_n11985_), .B(new_n11984_), .Y(new_n11994_));
  NOR4   g10992(.A(new_n11994_), .B(new_n11993_), .C(new_n11992_), .D(new_n11991_), .Y(new_n11995_));
  NOR2   g10993(.A(new_n11995_), .B(new_n11990_), .Y(new_n11996_));
  XOR2   g10994(.A(new_n11996_), .B(new_n11982_), .Y(new_n11997_));
  XOR2   g10995(.A(new_n11997_), .B(new_n11961_), .Y(new_n11998_));
  XOR2   g10996(.A(new_n11998_), .B(new_n11959_), .Y(new_n11999_));
  XOR2   g10997(.A(new_n11999_), .B(new_n11921_), .Y(new_n12000_));
  AOI22  g10998(.A0(new_n9603_), .A1(new_n9569_), .B0(new_n9349_), .B1(new_n9331_), .Y(new_n12001_));
  NOR2   g10999(.A(new_n12001_), .B(new_n9778_), .Y(new_n12002_));
  NOR3   g11000(.A(new_n9271_), .B(new_n9213_), .C(new_n9203_), .Y(new_n12003_));
  OAI21  g11001(.A0(new_n12003_), .A1(new_n9330_), .B0(new_n9347_), .Y(new_n12004_));
  NOR2   g11002(.A(new_n9328_), .B(new_n9327_), .Y(new_n12005_));
  AOI21  g11003(.A0(new_n9337_), .A1(new_n9312_), .B0(new_n9336_), .Y(new_n12006_));
  AOI21  g11004(.A0(new_n9302_), .A1(new_n9303_), .B0(new_n9301_), .Y(new_n12007_));
  OAI21  g11005(.A0(new_n9291_), .A1(new_n9317_), .B0(new_n9289_), .Y(new_n12008_));
  NOR2   g11006(.A(new_n12008_), .B(new_n12007_), .Y(new_n12009_));
  NAND2  g11007(.A(new_n9322_), .B(new_n9321_), .Y(new_n12010_));
  OAI21  g11008(.A0(new_n9315_), .A1(new_n9293_), .B0(new_n12010_), .Y(new_n12011_));
  AOI21  g11009(.A0(new_n9335_), .A1(new_n9273_), .B0(new_n9334_), .Y(new_n12012_));
  NOR2   g11010(.A(new_n12012_), .B(new_n12011_), .Y(new_n12013_));
  OAI22  g11011(.A0(new_n12013_), .A1(new_n12009_), .B0(new_n12006_), .B1(new_n12005_), .Y(new_n12014_));
  NOR4   g11012(.A(new_n9317_), .B(new_n9315_), .C(new_n12010_), .D(new_n9293_), .Y(new_n12015_));
  OAI211 g11013(.A0(new_n9301_), .A1(new_n9293_), .B0(new_n12015_), .B1(new_n9311_), .Y(new_n12016_));
  NAND2  g11014(.A(new_n9326_), .B(new_n9292_), .Y(new_n12017_));
  NAND2  g11015(.A(new_n12012_), .B(new_n12011_), .Y(new_n12018_));
  NAND2  g11016(.A(new_n12008_), .B(new_n12007_), .Y(new_n12019_));
  NAND4  g11017(.A(new_n12019_), .B(new_n12018_), .C(new_n12017_), .D(new_n12016_), .Y(new_n12020_));
  NAND2  g11018(.A(new_n12020_), .B(new_n12014_), .Y(new_n12021_));
  AOI21  g11019(.A0(new_n9209_), .A1(new_n9145_), .B0(new_n9344_), .Y(new_n12022_));
  NAND2  g11020(.A(new_n9200_), .B(new_n9199_), .Y(new_n12023_));
  OAI21  g11021(.A0(new_n9175_), .A1(new_n9188_), .B0(new_n12023_), .Y(new_n12024_));
  AOI21  g11022(.A0(new_n9132_), .A1(new_n9204_), .B0(new_n9207_), .Y(new_n12025_));
  NAND2  g11023(.A(new_n12025_), .B(new_n12024_), .Y(new_n12026_));
  AOI21  g11024(.A0(new_n9182_), .A1(new_n9170_), .B0(new_n9169_), .Y(new_n12027_));
  OAI21  g11025(.A0(new_n9189_), .A1(new_n9131_), .B0(new_n9144_), .Y(new_n12028_));
  NAND2  g11026(.A(new_n12028_), .B(new_n12027_), .Y(new_n12029_));
  AOI21  g11027(.A0(new_n12029_), .A1(new_n12026_), .B0(new_n12022_), .Y(new_n12030_));
  AOI21  g11028(.A0(new_n9258_), .A1(new_n9183_), .B0(new_n9208_), .Y(new_n12031_));
  NOR2   g11029(.A(new_n12028_), .B(new_n12027_), .Y(new_n12032_));
  NOR2   g11030(.A(new_n12025_), .B(new_n12024_), .Y(new_n12033_));
  NOR4   g11031(.A(new_n12033_), .B(new_n12032_), .C(new_n12031_), .D(new_n9344_), .Y(new_n12034_));
  NOR2   g11032(.A(new_n12034_), .B(new_n12030_), .Y(new_n12035_));
  XOR2   g11033(.A(new_n12035_), .B(new_n12021_), .Y(new_n12036_));
  XOR2   g11034(.A(new_n12036_), .B(new_n12004_), .Y(new_n12037_));
  NOR3   g11035(.A(new_n9567_), .B(new_n9549_), .C(new_n9539_), .Y(new_n12038_));
  OAI21  g11036(.A0(new_n12038_), .A1(new_n9445_), .B0(new_n9584_), .Y(new_n12039_));
  NAND2  g11037(.A(new_n9438_), .B(new_n9437_), .Y(new_n12040_));
  NAND3  g11038(.A(new_n9441_), .B(new_n9414_), .C(new_n9427_), .Y(new_n12041_));
  AOI211 g11039(.A0(new_n9427_), .A1(new_n12040_), .B(new_n12041_), .C(new_n9439_), .Y(new_n12042_));
  AOI21  g11040(.A0(new_n9429_), .A1(new_n9422_), .B0(new_n9387_), .Y(new_n12043_));
  AOI21  g11041(.A0(new_n9421_), .A1(new_n9427_), .B0(new_n9426_), .Y(new_n12044_));
  OAI21  g11042(.A0(new_n9376_), .A1(new_n9570_), .B0(new_n9572_), .Y(new_n12045_));
  NOR2   g11043(.A(new_n12045_), .B(new_n12044_), .Y(new_n12046_));
  OAI21  g11044(.A0(new_n9428_), .A1(new_n9432_), .B0(new_n12040_), .Y(new_n12047_));
  AOI21  g11045(.A0(new_n9388_), .A1(new_n9371_), .B0(new_n9386_), .Y(new_n12048_));
  NOR2   g11046(.A(new_n12048_), .B(new_n12047_), .Y(new_n12049_));
  OAI22  g11047(.A0(new_n12049_), .A1(new_n12046_), .B0(new_n12043_), .B1(new_n12042_), .Y(new_n12050_));
  NAND2  g11048(.A(new_n9440_), .B(new_n9573_), .Y(new_n12051_));
  NAND2  g11049(.A(new_n12048_), .B(new_n12047_), .Y(new_n12052_));
  NAND2  g11050(.A(new_n12045_), .B(new_n12044_), .Y(new_n12053_));
  NAND4  g11051(.A(new_n12053_), .B(new_n12052_), .C(new_n12051_), .D(new_n9443_), .Y(new_n12054_));
  NAND2  g11052(.A(new_n12054_), .B(new_n12050_), .Y(new_n12055_));
  AOI21  g11053(.A0(new_n9558_), .A1(new_n9519_), .B0(new_n9544_), .Y(new_n12056_));
  AOI21  g11054(.A0(new_n9518_), .A1(new_n9506_), .B0(new_n9505_), .Y(new_n12057_));
  OAI21  g11055(.A0(new_n9525_), .A1(new_n9467_), .B0(new_n9480_), .Y(new_n12058_));
  NOR2   g11056(.A(new_n12058_), .B(new_n12057_), .Y(new_n12059_));
  NAND2  g11057(.A(new_n9536_), .B(new_n9535_), .Y(new_n12060_));
  OAI21  g11058(.A0(new_n9511_), .A1(new_n9524_), .B0(new_n12060_), .Y(new_n12061_));
  AOI21  g11059(.A0(new_n9468_), .A1(new_n9540_), .B0(new_n9543_), .Y(new_n12062_));
  NOR2   g11060(.A(new_n12062_), .B(new_n12061_), .Y(new_n12063_));
  OAI22  g11061(.A0(new_n12063_), .A1(new_n12059_), .B0(new_n12056_), .B1(new_n9581_), .Y(new_n12064_));
  NAND2  g11062(.A(new_n9545_), .B(new_n9481_), .Y(new_n12065_));
  NAND2  g11063(.A(new_n12062_), .B(new_n12061_), .Y(new_n12066_));
  NAND2  g11064(.A(new_n12058_), .B(new_n12057_), .Y(new_n12067_));
  NAND4  g11065(.A(new_n12067_), .B(new_n12066_), .C(new_n12065_), .D(new_n9548_), .Y(new_n12068_));
  NAND2  g11066(.A(new_n12068_), .B(new_n12064_), .Y(new_n12069_));
  XOR2   g11067(.A(new_n12069_), .B(new_n12055_), .Y(new_n12070_));
  XOR2   g11068(.A(new_n12070_), .B(new_n12039_), .Y(new_n12071_));
  XOR2   g11069(.A(new_n12071_), .B(new_n12037_), .Y(new_n12072_));
  XOR2   g11070(.A(new_n12072_), .B(new_n12002_), .Y(new_n12073_));
  XOR2   g11071(.A(new_n12073_), .B(new_n12000_), .Y(new_n12074_));
  XOR2   g11072(.A(new_n12074_), .B(new_n11920_), .Y(new_n12075_));
  OAI21  g11073(.A0(new_n11131_), .A1(new_n10611_), .B0(new_n11142_), .Y(new_n12076_));
  OAI21  g11074(.A0(new_n11127_), .A1(new_n10606_), .B0(new_n10609_), .Y(new_n12077_));
  OAI22  g11075(.A0(new_n10583_), .A1(new_n10578_), .B0(new_n10518_), .B1(new_n10513_), .Y(new_n12078_));
  NOR2   g11076(.A(new_n10576_), .B(new_n10575_), .Y(new_n12079_));
  OAI21  g11077(.A0(new_n10548_), .A1(new_n10540_), .B0(new_n10549_), .Y(new_n12080_));
  AOI221 g11078(.A0(new_n12080_), .A1(new_n10559_), .C0(new_n10538_), .B0(new_n10536_), .B1(new_n10520_), .Y(new_n12081_));
  AOI21  g11079(.A0(new_n10549_), .A1(new_n10550_), .B0(new_n10548_), .Y(new_n12082_));
  OAI21  g11080(.A0(new_n10538_), .A1(new_n10564_), .B0(new_n10536_), .Y(new_n12083_));
  NOR2   g11081(.A(new_n12083_), .B(new_n12082_), .Y(new_n12084_));
  NAND2  g11082(.A(new_n10570_), .B(new_n10569_), .Y(new_n12085_));
  OAI21  g11083(.A0(new_n10562_), .A1(new_n10540_), .B0(new_n12085_), .Y(new_n12086_));
  XOR2   g11084(.A(new_n10433_), .B(new_n10431_), .Y(new_n12087_));
  NAND2  g11085(.A(new_n10537_), .B(new_n12087_), .Y(new_n12088_));
  XOR2   g11086(.A(new_n10537_), .B(new_n12087_), .Y(new_n12089_));
  AOI22  g11087(.A0(new_n12089_), .A1(new_n10520_), .B0(new_n10535_), .B1(new_n12088_), .Y(new_n12090_));
  NOR2   g11088(.A(new_n12090_), .B(new_n12086_), .Y(new_n12091_));
  OAI22  g11089(.A0(new_n12091_), .A1(new_n12084_), .B0(new_n12081_), .B1(new_n12079_), .Y(new_n12092_));
  NOR4   g11090(.A(new_n10564_), .B(new_n10562_), .C(new_n12085_), .D(new_n10540_), .Y(new_n12093_));
  OAI211 g11091(.A0(new_n10548_), .A1(new_n10540_), .B0(new_n12093_), .B1(new_n10558_), .Y(new_n12094_));
  OAI21  g11092(.A0(new_n10574_), .A1(new_n10566_), .B0(new_n10539_), .Y(new_n12095_));
  NAND2  g11093(.A(new_n12090_), .B(new_n12086_), .Y(new_n12096_));
  NAND2  g11094(.A(new_n12083_), .B(new_n12082_), .Y(new_n12097_));
  NAND4  g11095(.A(new_n12097_), .B(new_n12096_), .C(new_n12095_), .D(new_n12094_), .Y(new_n12098_));
  NAND2  g11096(.A(new_n12098_), .B(new_n12092_), .Y(new_n12099_));
  NAND2  g11097(.A(new_n10504_), .B(new_n10465_), .Y(new_n12100_));
  OAI21  g11098(.A0(new_n10492_), .A1(new_n10470_), .B0(new_n10598_), .Y(new_n12101_));
  AOI21  g11099(.A0(new_n10591_), .A1(new_n10446_), .B0(new_n10590_), .Y(new_n12102_));
  NAND2  g11100(.A(new_n12102_), .B(new_n12101_), .Y(new_n12103_));
  AOI21  g11101(.A0(new_n10479_), .A1(new_n10480_), .B0(new_n10478_), .Y(new_n12104_));
  OAI21  g11102(.A0(new_n10464_), .A1(new_n10494_), .B0(new_n10462_), .Y(new_n12105_));
  NAND2  g11103(.A(new_n12105_), .B(new_n12104_), .Y(new_n12106_));
  AOI22  g11104(.A0(new_n12106_), .A1(new_n12103_), .B0(new_n12100_), .B1(new_n10600_), .Y(new_n12107_));
  NOR2   g11105(.A(new_n10506_), .B(new_n10505_), .Y(new_n12108_));
  AOI21  g11106(.A0(new_n10593_), .A1(new_n10489_), .B0(new_n10592_), .Y(new_n12109_));
  NOR2   g11107(.A(new_n12105_), .B(new_n12104_), .Y(new_n12110_));
  NOR2   g11108(.A(new_n12102_), .B(new_n12101_), .Y(new_n12111_));
  NOR4   g11109(.A(new_n12111_), .B(new_n12110_), .C(new_n12109_), .D(new_n12108_), .Y(new_n12112_));
  NOR2   g11110(.A(new_n12112_), .B(new_n12107_), .Y(new_n12113_));
  XOR2   g11111(.A(new_n12113_), .B(new_n12099_), .Y(new_n12114_));
  XOR2   g11112(.A(new_n12114_), .B(new_n12078_), .Y(new_n12115_));
  NOR3   g11113(.A(new_n10339_), .B(new_n10321_), .C(new_n10311_), .Y(new_n12116_));
  OAI21  g11114(.A0(new_n12116_), .A1(new_n10217_), .B0(new_n10353_), .Y(new_n12117_));
  AOI21  g11115(.A0(new_n10201_), .A1(new_n10194_), .B0(new_n10159_), .Y(new_n12118_));
  AOI21  g11116(.A0(new_n10193_), .A1(new_n10199_), .B0(new_n10198_), .Y(new_n12119_));
  XOR2   g11117(.A(new_n10142_), .B(new_n10153_), .Y(new_n12120_));
  NOR2   g11118(.A(new_n10142_), .B(new_n10135_), .Y(new_n12121_));
  OAI22  g11119(.A0(new_n10157_), .A1(new_n12121_), .B0(new_n10148_), .B1(new_n12120_), .Y(new_n12122_));
  NOR2   g11120(.A(new_n12122_), .B(new_n12119_), .Y(new_n12123_));
  OAI21  g11121(.A0(new_n10200_), .A1(new_n10204_), .B0(new_n10343_), .Y(new_n12124_));
  AOI21  g11122(.A0(new_n10160_), .A1(new_n10143_), .B0(new_n10158_), .Y(new_n12125_));
  NOR2   g11123(.A(new_n12125_), .B(new_n12124_), .Y(new_n12126_));
  OAI22  g11124(.A0(new_n12126_), .A1(new_n12123_), .B0(new_n12118_), .B1(new_n10345_), .Y(new_n12127_));
  OAI211 g11125(.A0(new_n10158_), .A1(new_n10148_), .B0(new_n10212_), .B1(new_n10143_), .Y(new_n12128_));
  NAND2  g11126(.A(new_n12125_), .B(new_n12124_), .Y(new_n12129_));
  NAND2  g11127(.A(new_n12122_), .B(new_n12119_), .Y(new_n12130_));
  NAND4  g11128(.A(new_n12130_), .B(new_n12129_), .C(new_n12128_), .D(new_n10215_), .Y(new_n12131_));
  NAND2  g11129(.A(new_n12131_), .B(new_n12127_), .Y(new_n12132_));
  AOI21  g11130(.A0(new_n10317_), .A1(new_n10253_), .B0(new_n10350_), .Y(new_n12133_));
  NAND2  g11131(.A(new_n10308_), .B(new_n10307_), .Y(new_n12134_));
  OAI21  g11132(.A0(new_n10283_), .A1(new_n10296_), .B0(new_n12134_), .Y(new_n12135_));
  AOI21  g11133(.A0(new_n10240_), .A1(new_n10312_), .B0(new_n10315_), .Y(new_n12136_));
  NAND2  g11134(.A(new_n12136_), .B(new_n12135_), .Y(new_n12137_));
  AOI21  g11135(.A0(new_n10290_), .A1(new_n10278_), .B0(new_n10277_), .Y(new_n12138_));
  OAI21  g11136(.A0(new_n10297_), .A1(new_n10239_), .B0(new_n10252_), .Y(new_n12139_));
  NAND2  g11137(.A(new_n12139_), .B(new_n12138_), .Y(new_n12140_));
  AOI21  g11138(.A0(new_n12140_), .A1(new_n12137_), .B0(new_n12133_), .Y(new_n12141_));
  AOI21  g11139(.A0(new_n10330_), .A1(new_n10291_), .B0(new_n10316_), .Y(new_n12142_));
  NOR2   g11140(.A(new_n12139_), .B(new_n12138_), .Y(new_n12143_));
  NOR2   g11141(.A(new_n12136_), .B(new_n12135_), .Y(new_n12144_));
  NOR4   g11142(.A(new_n12144_), .B(new_n12143_), .C(new_n12142_), .D(new_n10350_), .Y(new_n12145_));
  NOR2   g11143(.A(new_n12145_), .B(new_n12141_), .Y(new_n12146_));
  XOR2   g11144(.A(new_n12146_), .B(new_n12132_), .Y(new_n12147_));
  XOR2   g11145(.A(new_n12147_), .B(new_n12117_), .Y(new_n12148_));
  XOR2   g11146(.A(new_n12148_), .B(new_n12115_), .Y(new_n12149_));
  XOR2   g11147(.A(new_n12149_), .B(new_n12077_), .Y(new_n12150_));
  AOI22  g11148(.A0(new_n11105_), .A1(new_n11071_), .B0(new_n10851_), .B1(new_n10833_), .Y(new_n12151_));
  NOR2   g11149(.A(new_n12151_), .B(new_n11120_), .Y(new_n12152_));
  NOR3   g11150(.A(new_n10773_), .B(new_n10715_), .C(new_n10705_), .Y(new_n12153_));
  OAI21  g11151(.A0(new_n12153_), .A1(new_n10832_), .B0(new_n10849_), .Y(new_n12154_));
  NOR2   g11152(.A(new_n10830_), .B(new_n10829_), .Y(new_n12155_));
  AOI21  g11153(.A0(new_n10839_), .A1(new_n10814_), .B0(new_n10838_), .Y(new_n12156_));
  AOI21  g11154(.A0(new_n10804_), .A1(new_n10805_), .B0(new_n10803_), .Y(new_n12157_));
  OAI21  g11155(.A0(new_n10793_), .A1(new_n10819_), .B0(new_n10791_), .Y(new_n12158_));
  NOR2   g11156(.A(new_n12158_), .B(new_n12157_), .Y(new_n12159_));
  NAND2  g11157(.A(new_n10824_), .B(new_n10823_), .Y(new_n12160_));
  OAI21  g11158(.A0(new_n10817_), .A1(new_n10795_), .B0(new_n12160_), .Y(new_n12161_));
  AOI21  g11159(.A0(new_n10837_), .A1(new_n10775_), .B0(new_n10836_), .Y(new_n12162_));
  NOR2   g11160(.A(new_n12162_), .B(new_n12161_), .Y(new_n12163_));
  OAI22  g11161(.A0(new_n12163_), .A1(new_n12159_), .B0(new_n12156_), .B1(new_n12155_), .Y(new_n12164_));
  NOR4   g11162(.A(new_n10819_), .B(new_n10817_), .C(new_n12160_), .D(new_n10795_), .Y(new_n12165_));
  OAI211 g11163(.A0(new_n10803_), .A1(new_n10795_), .B0(new_n12165_), .B1(new_n10813_), .Y(new_n12166_));
  NAND2  g11164(.A(new_n10828_), .B(new_n10794_), .Y(new_n12167_));
  NAND2  g11165(.A(new_n12162_), .B(new_n12161_), .Y(new_n12168_));
  NAND2  g11166(.A(new_n12158_), .B(new_n12157_), .Y(new_n12169_));
  NAND4  g11167(.A(new_n12169_), .B(new_n12168_), .C(new_n12167_), .D(new_n12166_), .Y(new_n12170_));
  NAND2  g11168(.A(new_n12170_), .B(new_n12164_), .Y(new_n12171_));
  AOI21  g11169(.A0(new_n10711_), .A1(new_n10647_), .B0(new_n10846_), .Y(new_n12172_));
  NAND2  g11170(.A(new_n10702_), .B(new_n10701_), .Y(new_n12173_));
  OAI21  g11171(.A0(new_n10677_), .A1(new_n10690_), .B0(new_n12173_), .Y(new_n12174_));
  AOI21  g11172(.A0(new_n10634_), .A1(new_n10706_), .B0(new_n10709_), .Y(new_n12175_));
  NAND2  g11173(.A(new_n12175_), .B(new_n12174_), .Y(new_n12176_));
  AOI21  g11174(.A0(new_n10684_), .A1(new_n10672_), .B0(new_n10671_), .Y(new_n12177_));
  OAI21  g11175(.A0(new_n10691_), .A1(new_n10633_), .B0(new_n10646_), .Y(new_n12178_));
  NAND2  g11176(.A(new_n12178_), .B(new_n12177_), .Y(new_n12179_));
  AOI21  g11177(.A0(new_n12179_), .A1(new_n12176_), .B0(new_n12172_), .Y(new_n12180_));
  AOI21  g11178(.A0(new_n10760_), .A1(new_n10685_), .B0(new_n10710_), .Y(new_n12181_));
  NOR2   g11179(.A(new_n12178_), .B(new_n12177_), .Y(new_n12182_));
  NOR2   g11180(.A(new_n12175_), .B(new_n12174_), .Y(new_n12183_));
  NOR4   g11181(.A(new_n12183_), .B(new_n12182_), .C(new_n12181_), .D(new_n10846_), .Y(new_n12184_));
  NOR2   g11182(.A(new_n12184_), .B(new_n12180_), .Y(new_n12185_));
  XOR2   g11183(.A(new_n12185_), .B(new_n12171_), .Y(new_n12186_));
  XOR2   g11184(.A(new_n12186_), .B(new_n12154_), .Y(new_n12187_));
  NOR3   g11185(.A(new_n11069_), .B(new_n11051_), .C(new_n11041_), .Y(new_n12188_));
  OAI21  g11186(.A0(new_n12188_), .A1(new_n10947_), .B0(new_n11086_), .Y(new_n12189_));
  NAND2  g11187(.A(new_n10940_), .B(new_n10939_), .Y(new_n12190_));
  NAND3  g11188(.A(new_n10943_), .B(new_n10916_), .C(new_n10929_), .Y(new_n12191_));
  AOI211 g11189(.A0(new_n10929_), .A1(new_n12190_), .B(new_n12191_), .C(new_n10941_), .Y(new_n12192_));
  AOI21  g11190(.A0(new_n10931_), .A1(new_n10924_), .B0(new_n10889_), .Y(new_n12193_));
  AOI21  g11191(.A0(new_n10923_), .A1(new_n10929_), .B0(new_n10928_), .Y(new_n12194_));
  OAI21  g11192(.A0(new_n10878_), .A1(new_n11072_), .B0(new_n11074_), .Y(new_n12195_));
  NOR2   g11193(.A(new_n12195_), .B(new_n12194_), .Y(new_n12196_));
  OAI21  g11194(.A0(new_n10930_), .A1(new_n10934_), .B0(new_n12190_), .Y(new_n12197_));
  AOI21  g11195(.A0(new_n10890_), .A1(new_n10873_), .B0(new_n10888_), .Y(new_n12198_));
  NOR2   g11196(.A(new_n12198_), .B(new_n12197_), .Y(new_n12199_));
  OAI22  g11197(.A0(new_n12199_), .A1(new_n12196_), .B0(new_n12193_), .B1(new_n12192_), .Y(new_n12200_));
  NAND2  g11198(.A(new_n10942_), .B(new_n11075_), .Y(new_n12201_));
  NAND2  g11199(.A(new_n12198_), .B(new_n12197_), .Y(new_n12202_));
  NAND2  g11200(.A(new_n12195_), .B(new_n12194_), .Y(new_n12203_));
  NAND4  g11201(.A(new_n12203_), .B(new_n12202_), .C(new_n12201_), .D(new_n10945_), .Y(new_n12204_));
  NAND2  g11202(.A(new_n12204_), .B(new_n12200_), .Y(new_n12205_));
  AOI21  g11203(.A0(new_n11060_), .A1(new_n11021_), .B0(new_n11046_), .Y(new_n12206_));
  AOI21  g11204(.A0(new_n11020_), .A1(new_n11008_), .B0(new_n11007_), .Y(new_n12207_));
  OAI21  g11205(.A0(new_n11027_), .A1(new_n10969_), .B0(new_n10982_), .Y(new_n12208_));
  NOR2   g11206(.A(new_n12208_), .B(new_n12207_), .Y(new_n12209_));
  NAND2  g11207(.A(new_n11038_), .B(new_n11037_), .Y(new_n12210_));
  OAI21  g11208(.A0(new_n11013_), .A1(new_n11026_), .B0(new_n12210_), .Y(new_n12211_));
  AOI21  g11209(.A0(new_n10970_), .A1(new_n11042_), .B0(new_n11045_), .Y(new_n12212_));
  NOR2   g11210(.A(new_n12212_), .B(new_n12211_), .Y(new_n12213_));
  OAI22  g11211(.A0(new_n12213_), .A1(new_n12209_), .B0(new_n12206_), .B1(new_n11083_), .Y(new_n12214_));
  NAND2  g11212(.A(new_n11047_), .B(new_n10983_), .Y(new_n12215_));
  NAND2  g11213(.A(new_n12212_), .B(new_n12211_), .Y(new_n12216_));
  NAND2  g11214(.A(new_n12208_), .B(new_n12207_), .Y(new_n12217_));
  NAND4  g11215(.A(new_n12217_), .B(new_n12216_), .C(new_n12215_), .D(new_n11050_), .Y(new_n12218_));
  NAND2  g11216(.A(new_n12218_), .B(new_n12214_), .Y(new_n12219_));
  XOR2   g11217(.A(new_n12219_), .B(new_n12205_), .Y(new_n12220_));
  XOR2   g11218(.A(new_n12220_), .B(new_n12189_), .Y(new_n12221_));
  XOR2   g11219(.A(new_n12221_), .B(new_n12187_), .Y(new_n12222_));
  XOR2   g11220(.A(new_n12222_), .B(new_n12152_), .Y(new_n12223_));
  XOR2   g11221(.A(new_n12223_), .B(new_n12150_), .Y(new_n12224_));
  XOR2   g11222(.A(new_n12224_), .B(new_n12076_), .Y(new_n12225_));
  XOR2   g11223(.A(new_n12225_), .B(new_n12075_), .Y(new_n12226_));
  XOR2   g11224(.A(new_n12226_), .B(new_n11919_), .Y(new_n12227_));
  XOR2   g11225(.A(new_n12227_), .B(new_n11918_), .Y(new_n12228_));
  XOR2   g11226(.A(new_n12228_), .B(new_n11609_), .Y(new_n12229_));
  XOR2   g11227(.A(new_n12229_), .B(new_n11608_), .Y(new_n12230_));
  XOR2   g11228(.A(new_n12230_), .B(new_n11219_), .Y(new_n12231_));
  NOR3   g11229(.A(new_n4165_), .B(new_n4164_), .C(new_n4161_), .Y(new_n12232_));
  AOI21  g11230(.A0(new_n4156_), .A1(new_n4145_), .B0(new_n4157_), .Y(new_n12233_));
  OAI21  g11231(.A0(new_n12233_), .A1(new_n12232_), .B0(new_n4763_), .Y(new_n12234_));
  NOR3   g11232(.A(new_n4157_), .B(new_n4164_), .C(new_n4161_), .Y(new_n12235_));
  AOI21  g11233(.A0(new_n4156_), .A1(new_n4145_), .B0(new_n4165_), .Y(new_n12236_));
  OAI21  g11234(.A0(new_n12236_), .A1(new_n12235_), .B0(new_n4755_), .Y(new_n12237_));
  NAND2  g11235(.A(new_n12237_), .B(new_n12234_), .Y(new_n12238_));
  AOI21  g11236(.A0(new_n2876_), .A1(new_n2866_), .B0(new_n3555_), .Y(new_n12239_));
  AOI21  g11237(.A0(new_n4768_), .A1(new_n12238_), .B0(new_n12239_), .Y(new_n12240_));
  OAI21  g11238(.A0(new_n12235_), .A1(new_n4763_), .B0(new_n4765_), .Y(new_n12241_));
  OAI21  g11239(.A0(new_n4752_), .A1(new_n4742_), .B0(new_n4761_), .Y(new_n12242_));
  OAI21  g11240(.A0(new_n4748_), .A1(new_n4732_), .B0(new_n4740_), .Y(new_n12243_));
  NOR2   g11241(.A(new_n4638_), .B(new_n4615_), .Y(new_n12244_));
  AOI21  g11242(.A0(new_n4649_), .A1(new_n4615_), .B0(new_n12244_), .Y(new_n12245_));
  NOR3   g11243(.A(new_n4725_), .B(new_n4713_), .C(new_n4696_), .Y(new_n12246_));
  OAI22  g11244(.A0(new_n12246_), .A1(new_n12245_), .B0(new_n4729_), .B1(new_n4714_), .Y(new_n12247_));
  XOR2   g11245(.A(new_n4635_), .B(new_n4644_), .Y(new_n12248_));
  NAND4  g11246(.A(new_n2911_), .B(new_n4629_), .C(new_n12248_), .D(new_n4616_), .Y(new_n12249_));
  AOI211 g11247(.A0(new_n4634_), .A1(new_n4616_), .B(new_n12249_), .C(new_n4642_), .Y(new_n12250_));
  OAI21  g11248(.A0(new_n4646_), .A1(new_n4639_), .B0(new_n12248_), .Y(new_n12251_));
  AOI221 g11249(.A0(new_n12251_), .A1(new_n4630_), .C0(new_n4611_), .B0(new_n4614_), .B1(new_n2911_), .Y(new_n12252_));
  AOI21  g11250(.A0(new_n12248_), .A1(new_n4616_), .B0(new_n4646_), .Y(new_n12253_));
  OAI21  g11251(.A0(new_n4611_), .A1(new_n4641_), .B0(new_n4614_), .Y(new_n12254_));
  NOR2   g11252(.A(new_n12254_), .B(new_n12253_), .Y(new_n12255_));
  OAI21  g11253(.A0(new_n4636_), .A1(new_n4639_), .B0(new_n4634_), .Y(new_n12256_));
  XOR2   g11254(.A(new_n4610_), .B(new_n4612_), .Y(new_n12257_));
  XOR2   g11255(.A(new_n2924_), .B(new_n2922_), .Y(new_n12258_));
  NAND2  g11256(.A(new_n12258_), .B(new_n4607_), .Y(new_n12259_));
  AOI22  g11257(.A0(new_n4613_), .A1(new_n12259_), .B0(new_n12257_), .B1(new_n2911_), .Y(new_n12260_));
  NOR2   g11258(.A(new_n12260_), .B(new_n12256_), .Y(new_n12261_));
  OAI22  g11259(.A0(new_n12261_), .A1(new_n12255_), .B0(new_n12252_), .B1(new_n12250_), .Y(new_n12262_));
  OAI21  g11260(.A0(new_n4637_), .A1(new_n4643_), .B0(new_n4615_), .Y(new_n12263_));
  NAND2  g11261(.A(new_n12260_), .B(new_n12256_), .Y(new_n12264_));
  NAND2  g11262(.A(new_n12254_), .B(new_n12253_), .Y(new_n12265_));
  NAND4  g11263(.A(new_n12265_), .B(new_n12264_), .C(new_n12263_), .D(new_n4648_), .Y(new_n12266_));
  NAND2  g11264(.A(new_n12266_), .B(new_n12262_), .Y(new_n12267_));
  OAI21  g11265(.A0(new_n4694_), .A1(new_n4717_), .B0(new_n4671_), .Y(new_n12268_));
  OAI21  g11266(.A0(new_n4693_), .A1(new_n4703_), .B0(new_n4691_), .Y(new_n12269_));
  AOI21  g11267(.A0(new_n4701_), .A1(new_n4652_), .B0(new_n4700_), .Y(new_n12270_));
  NAND2  g11268(.A(new_n12270_), .B(new_n12269_), .Y(new_n12271_));
  AOI21  g11269(.A0(new_n4707_), .A1(new_n4672_), .B0(new_n4706_), .Y(new_n12272_));
  OAI21  g11270(.A0(new_n4670_), .A1(new_n4697_), .B0(new_n4668_), .Y(new_n12273_));
  NAND2  g11271(.A(new_n12273_), .B(new_n12272_), .Y(new_n12274_));
  AOI22  g11272(.A0(new_n12274_), .A1(new_n12271_), .B0(new_n12268_), .B1(new_n4712_), .Y(new_n12275_));
  NOR2   g11273(.A(new_n4721_), .B(new_n4720_), .Y(new_n12276_));
  AOI21  g11274(.A0(new_n4708_), .A1(new_n4687_), .B0(new_n4702_), .Y(new_n12277_));
  NOR2   g11275(.A(new_n12273_), .B(new_n12272_), .Y(new_n12278_));
  NOR2   g11276(.A(new_n12270_), .B(new_n12269_), .Y(new_n12279_));
  NOR4   g11277(.A(new_n12279_), .B(new_n12278_), .C(new_n12277_), .D(new_n12276_), .Y(new_n12280_));
  NOR2   g11278(.A(new_n12280_), .B(new_n12275_), .Y(new_n12281_));
  XOR2   g11279(.A(new_n12281_), .B(new_n12267_), .Y(new_n12282_));
  XOR2   g11280(.A(new_n12282_), .B(new_n12247_), .Y(new_n12283_));
  OAI22  g11281(.A0(new_n4598_), .A1(new_n4594_), .B0(new_n4733_), .B1(new_n4587_), .Y(new_n12284_));
  XOR2   g11282(.A(new_n4508_), .B(new_n4517_), .Y(new_n12285_));
  NAND4  g11283(.A(new_n4468_), .B(new_n4501_), .C(new_n12285_), .D(new_n4488_), .Y(new_n12286_));
  AOI211 g11284(.A0(new_n4507_), .A1(new_n4488_), .B(new_n12286_), .C(new_n4515_), .Y(new_n12287_));
  OAI21  g11285(.A0(new_n4519_), .A1(new_n4512_), .B0(new_n12285_), .Y(new_n12288_));
  AOI221 g11286(.A0(new_n12288_), .A1(new_n4503_), .C0(new_n4486_), .B0(new_n4484_), .B1(new_n4468_), .Y(new_n12289_));
  OAI21  g11287(.A0(new_n4509_), .A1(new_n4512_), .B0(new_n4507_), .Y(new_n12290_));
  OAI21  g11288(.A0(new_n4486_), .A1(new_n4514_), .B0(new_n4484_), .Y(new_n12291_));
  XOR2   g11289(.A(new_n12291_), .B(new_n12290_), .Y(new_n12292_));
  OAI21  g11290(.A0(new_n12289_), .A1(new_n12287_), .B0(new_n12292_), .Y(new_n12293_));
  OAI21  g11291(.A0(new_n4510_), .A1(new_n4516_), .B0(new_n4487_), .Y(new_n12294_));
  XOR2   g11292(.A(new_n3045_), .B(new_n3043_), .Y(new_n12295_));
  NAND2  g11293(.A(new_n4485_), .B(new_n12295_), .Y(new_n12296_));
  XOR2   g11294(.A(new_n4485_), .B(new_n12295_), .Y(new_n12297_));
  AOI22  g11295(.A0(new_n12297_), .A1(new_n4468_), .B0(new_n4483_), .B1(new_n12296_), .Y(new_n12298_));
  NAND2  g11296(.A(new_n12298_), .B(new_n12290_), .Y(new_n12299_));
  AOI21  g11297(.A0(new_n12285_), .A1(new_n4488_), .B0(new_n4519_), .Y(new_n12300_));
  NAND2  g11298(.A(new_n12291_), .B(new_n12300_), .Y(new_n12301_));
  NAND4  g11299(.A(new_n12301_), .B(new_n12299_), .C(new_n12294_), .D(new_n4521_), .Y(new_n12302_));
  NAND2  g11300(.A(new_n12302_), .B(new_n12293_), .Y(new_n12303_));
  NOR4   g11301(.A(new_n4529_), .B(new_n4541_), .C(new_n4558_), .D(new_n4540_), .Y(new_n12304_));
  OAI211 g11302(.A0(new_n4582_), .A1(new_n4540_), .B0(new_n12304_), .B1(new_n4583_), .Y(new_n12305_));
  OAI21  g11303(.A0(new_n4559_), .A1(new_n4543_), .B0(new_n4576_), .Y(new_n12306_));
  OAI21  g11304(.A0(new_n4558_), .A1(new_n4540_), .B0(new_n4556_), .Y(new_n12307_));
  AOI21  g11305(.A0(new_n4534_), .A1(new_n4562_), .B0(new_n4533_), .Y(new_n12308_));
  NAND2  g11306(.A(new_n12308_), .B(new_n12307_), .Y(new_n12309_));
  AOI21  g11307(.A0(new_n4578_), .A1(new_n4544_), .B0(new_n4582_), .Y(new_n12310_));
  OAI21  g11308(.A0(new_n4575_), .A1(new_n4529_), .B0(new_n4574_), .Y(new_n12311_));
  NAND2  g11309(.A(new_n12311_), .B(new_n12310_), .Y(new_n12312_));
  AOI22  g11310(.A0(new_n12312_), .A1(new_n12309_), .B0(new_n12306_), .B1(new_n12305_), .Y(new_n12313_));
  OAI21  g11311(.A0(new_n4582_), .A1(new_n4540_), .B0(new_n4578_), .Y(new_n12314_));
  AOI21  g11312(.A0(new_n12314_), .A1(new_n4595_), .B0(new_n4535_), .Y(new_n12315_));
  OAI22  g11313(.A0(new_n12311_), .A1(new_n12310_), .B0(new_n4584_), .B1(new_n4580_), .Y(new_n12316_));
  AOI211 g11314(.A0(new_n12311_), .A1(new_n12310_), .B(new_n12316_), .C(new_n12315_), .Y(new_n12317_));
  NOR2   g11315(.A(new_n12317_), .B(new_n12313_), .Y(new_n12318_));
  XOR2   g11316(.A(new_n12318_), .B(new_n12303_), .Y(new_n12319_));
  XOR2   g11317(.A(new_n12319_), .B(new_n12284_), .Y(new_n12320_));
  XOR2   g11318(.A(new_n12320_), .B(new_n12283_), .Y(new_n12321_));
  XOR2   g11319(.A(new_n12321_), .B(new_n12243_), .Y(new_n12322_));
  OAI21  g11320(.A0(new_n4464_), .A1(new_n4452_), .B0(new_n4456_), .Y(new_n12323_));
  AOI21  g11321(.A0(new_n4223_), .A1(new_n4186_), .B0(new_n4211_), .Y(new_n12324_));
  OAI22  g11322(.A0(new_n4293_), .A1(new_n4291_), .B0(new_n12324_), .B1(new_n4224_), .Y(new_n12325_));
  NAND4  g11323(.A(new_n4236_), .B(new_n4260_), .C(new_n4285_), .D(new_n4247_), .Y(new_n12326_));
  AOI221 g11324(.A0(new_n4279_), .A1(new_n4240_), .C0(new_n12326_), .B0(new_n4268_), .B1(new_n4247_), .Y(new_n12327_));
  AOI21  g11325(.A0(new_n4286_), .A1(new_n4264_), .B0(new_n4280_), .Y(new_n12328_));
  AOI21  g11326(.A0(new_n4285_), .A1(new_n4247_), .B0(new_n4284_), .Y(new_n12329_));
  AOI211 g11327(.A0(new_n4279_), .A1(new_n4236_), .B(new_n12329_), .C(new_n4278_), .Y(new_n12330_));
  OAI21  g11328(.A0(new_n4270_), .A1(new_n4281_), .B0(new_n4268_), .Y(new_n12331_));
  AOI21  g11329(.A0(new_n4279_), .A1(new_n4236_), .B0(new_n4278_), .Y(new_n12332_));
  NOR2   g11330(.A(new_n12332_), .B(new_n12331_), .Y(new_n12333_));
  OAI22  g11331(.A0(new_n12333_), .A1(new_n12330_), .B0(new_n12328_), .B1(new_n12327_), .Y(new_n12334_));
  NAND2  g11332(.A(new_n4287_), .B(new_n4246_), .Y(new_n12335_));
  NAND2  g11333(.A(new_n12332_), .B(new_n12331_), .Y(new_n12336_));
  OAI21  g11334(.A0(new_n4245_), .A1(new_n4276_), .B0(new_n4240_), .Y(new_n12337_));
  NAND2  g11335(.A(new_n12337_), .B(new_n12329_), .Y(new_n12338_));
  NAND4  g11336(.A(new_n12338_), .B(new_n12336_), .C(new_n12335_), .D(new_n4289_), .Y(new_n12339_));
  NAND2  g11337(.A(new_n12339_), .B(new_n12334_), .Y(new_n12340_));
  NOR4   g11338(.A(new_n4214_), .B(new_n4213_), .C(new_n4208_), .D(new_n4212_), .Y(new_n12341_));
  OAI211 g11339(.A0(new_n4221_), .A1(new_n4212_), .B0(new_n12341_), .B1(new_n4201_), .Y(new_n12342_));
  OAI21  g11340(.A0(new_n4209_), .A1(new_n4216_), .B0(new_n4186_), .Y(new_n12343_));
  OAI21  g11341(.A0(new_n4208_), .A1(new_n4212_), .B0(new_n4206_), .Y(new_n12344_));
  AOI21  g11342(.A0(new_n4229_), .A1(new_n4167_), .B0(new_n4228_), .Y(new_n12345_));
  NAND2  g11343(.A(new_n12345_), .B(new_n12344_), .Y(new_n12346_));
  AOI21  g11344(.A0(new_n4218_), .A1(new_n4187_), .B0(new_n4221_), .Y(new_n12347_));
  OAI21  g11345(.A0(new_n4185_), .A1(new_n4214_), .B0(new_n4183_), .Y(new_n12348_));
  NAND2  g11346(.A(new_n12348_), .B(new_n12347_), .Y(new_n12349_));
  AOI22  g11347(.A0(new_n12349_), .A1(new_n12346_), .B0(new_n12343_), .B1(new_n12342_), .Y(new_n12350_));
  NOR2   g11348(.A(new_n4222_), .B(new_n4219_), .Y(new_n12351_));
  OAI21  g11349(.A0(new_n4221_), .A1(new_n4212_), .B0(new_n4218_), .Y(new_n12352_));
  AOI21  g11350(.A0(new_n12352_), .A1(new_n4202_), .B0(new_n4230_), .Y(new_n12353_));
  NOR2   g11351(.A(new_n12348_), .B(new_n12347_), .Y(new_n12354_));
  NOR2   g11352(.A(new_n12345_), .B(new_n12344_), .Y(new_n12355_));
  NOR4   g11353(.A(new_n12355_), .B(new_n12354_), .C(new_n12353_), .D(new_n12351_), .Y(new_n12356_));
  NOR2   g11354(.A(new_n12356_), .B(new_n12350_), .Y(new_n12357_));
  XOR2   g11355(.A(new_n12357_), .B(new_n12340_), .Y(new_n12358_));
  XOR2   g11356(.A(new_n12358_), .B(new_n12325_), .Y(new_n12359_));
  OAI22  g11357(.A0(new_n4423_), .A1(new_n4352_), .B0(new_n4420_), .B1(new_n4353_), .Y(new_n12360_));
  NAND4  g11358(.A(new_n4297_), .B(new_n4321_), .C(new_n4346_), .D(new_n4308_), .Y(new_n12361_));
  AOI221 g11359(.A0(new_n4340_), .A1(new_n4301_), .C0(new_n12361_), .B0(new_n4329_), .B1(new_n4308_), .Y(new_n12362_));
  AOI21  g11360(.A0(new_n4347_), .A1(new_n4325_), .B0(new_n4341_), .Y(new_n12363_));
  AOI21  g11361(.A0(new_n4346_), .A1(new_n4308_), .B0(new_n4345_), .Y(new_n12364_));
  AOI211 g11362(.A0(new_n4340_), .A1(new_n4297_), .B(new_n12364_), .C(new_n4339_), .Y(new_n12365_));
  OAI21  g11363(.A0(new_n4331_), .A1(new_n4342_), .B0(new_n4329_), .Y(new_n12366_));
  AOI21  g11364(.A0(new_n4340_), .A1(new_n4297_), .B0(new_n4339_), .Y(new_n12367_));
  NOR2   g11365(.A(new_n12367_), .B(new_n12366_), .Y(new_n12368_));
  OAI22  g11366(.A0(new_n12368_), .A1(new_n12365_), .B0(new_n12363_), .B1(new_n12362_), .Y(new_n12369_));
  NAND2  g11367(.A(new_n4348_), .B(new_n4307_), .Y(new_n12370_));
  NAND2  g11368(.A(new_n12367_), .B(new_n12366_), .Y(new_n12371_));
  OAI21  g11369(.A0(new_n4306_), .A1(new_n4337_), .B0(new_n4301_), .Y(new_n12372_));
  NAND2  g11370(.A(new_n12372_), .B(new_n12364_), .Y(new_n12373_));
  NAND4  g11371(.A(new_n12373_), .B(new_n12371_), .C(new_n12370_), .D(new_n4350_), .Y(new_n12374_));
  NAND2  g11372(.A(new_n12374_), .B(new_n12369_), .Y(new_n12375_));
  NOR4   g11373(.A(new_n4359_), .B(new_n4371_), .C(new_n4388_), .D(new_n4370_), .Y(new_n12376_));
  OAI211 g11374(.A0(new_n4411_), .A1(new_n4370_), .B0(new_n12376_), .B1(new_n4412_), .Y(new_n12377_));
  OAI21  g11375(.A0(new_n4389_), .A1(new_n4373_), .B0(new_n4405_), .Y(new_n12378_));
  OAI21  g11376(.A0(new_n4388_), .A1(new_n4370_), .B0(new_n4386_), .Y(new_n12379_));
  AOI21  g11377(.A0(new_n4364_), .A1(new_n4392_), .B0(new_n4363_), .Y(new_n12380_));
  NAND2  g11378(.A(new_n12380_), .B(new_n12379_), .Y(new_n12381_));
  AOI21  g11379(.A0(new_n4407_), .A1(new_n4374_), .B0(new_n4411_), .Y(new_n12382_));
  OAI21  g11380(.A0(new_n4404_), .A1(new_n4359_), .B0(new_n4403_), .Y(new_n12383_));
  NAND2  g11381(.A(new_n12383_), .B(new_n12382_), .Y(new_n12384_));
  AOI22  g11382(.A0(new_n12384_), .A1(new_n12381_), .B0(new_n12378_), .B1(new_n12377_), .Y(new_n12385_));
  NOR2   g11383(.A(new_n4431_), .B(new_n4365_), .Y(new_n12386_));
  NOR2   g11384(.A(new_n12383_), .B(new_n12382_), .Y(new_n12387_));
  NOR2   g11385(.A(new_n12380_), .B(new_n12379_), .Y(new_n12388_));
  NOR4   g11386(.A(new_n12388_), .B(new_n12387_), .C(new_n12386_), .D(new_n4432_), .Y(new_n12389_));
  NOR2   g11387(.A(new_n12389_), .B(new_n12385_), .Y(new_n12390_));
  XOR2   g11388(.A(new_n12390_), .B(new_n12375_), .Y(new_n12391_));
  XOR2   g11389(.A(new_n12391_), .B(new_n12360_), .Y(new_n12392_));
  XOR2   g11390(.A(new_n12392_), .B(new_n12359_), .Y(new_n12393_));
  XOR2   g11391(.A(new_n12393_), .B(new_n12323_), .Y(new_n12394_));
  XOR2   g11392(.A(new_n12394_), .B(new_n12322_), .Y(new_n12395_));
  XOR2   g11393(.A(new_n12395_), .B(new_n12242_), .Y(new_n12396_));
  OAI21  g11394(.A0(new_n4154_), .A1(new_n3843_), .B0(new_n4163_), .Y(new_n12397_));
  OAI21  g11395(.A0(new_n4150_), .A1(new_n3833_), .B0(new_n3841_), .Y(new_n12398_));
  NOR2   g11396(.A(new_n3740_), .B(new_n3716_), .Y(new_n12399_));
  AOI21  g11397(.A0(new_n3751_), .A1(new_n3716_), .B0(new_n12399_), .Y(new_n12400_));
  NOR3   g11398(.A(new_n3826_), .B(new_n3815_), .C(new_n3798_), .Y(new_n12401_));
  OAI22  g11399(.A0(new_n12401_), .A1(new_n12400_), .B0(new_n3830_), .B1(new_n3816_), .Y(new_n12402_));
  XOR2   g11400(.A(new_n3737_), .B(new_n3746_), .Y(new_n12403_));
  NAND4  g11401(.A(new_n3697_), .B(new_n3730_), .C(new_n12403_), .D(new_n3717_), .Y(new_n12404_));
  AOI211 g11402(.A0(new_n3736_), .A1(new_n3717_), .B(new_n12404_), .C(new_n3744_), .Y(new_n12405_));
  OAI21  g11403(.A0(new_n3748_), .A1(new_n3741_), .B0(new_n12403_), .Y(new_n12406_));
  AOI221 g11404(.A0(new_n12406_), .A1(new_n3732_), .C0(new_n3715_), .B0(new_n3713_), .B1(new_n3697_), .Y(new_n12407_));
  AOI21  g11405(.A0(new_n12403_), .A1(new_n3717_), .B0(new_n3748_), .Y(new_n12408_));
  OAI21  g11406(.A0(new_n3715_), .A1(new_n3743_), .B0(new_n3713_), .Y(new_n12409_));
  NOR2   g11407(.A(new_n12409_), .B(new_n12408_), .Y(new_n12410_));
  OAI21  g11408(.A0(new_n3738_), .A1(new_n3741_), .B0(new_n3736_), .Y(new_n12411_));
  XOR2   g11409(.A(new_n3537_), .B(new_n3535_), .Y(new_n12412_));
  NAND2  g11410(.A(new_n3714_), .B(new_n12412_), .Y(new_n12413_));
  XOR2   g11411(.A(new_n3714_), .B(new_n12412_), .Y(new_n12414_));
  AOI22  g11412(.A0(new_n12414_), .A1(new_n3697_), .B0(new_n3712_), .B1(new_n12413_), .Y(new_n12415_));
  NOR2   g11413(.A(new_n12415_), .B(new_n12411_), .Y(new_n12416_));
  OAI22  g11414(.A0(new_n12416_), .A1(new_n12410_), .B0(new_n12407_), .B1(new_n12405_), .Y(new_n12417_));
  OAI21  g11415(.A0(new_n3739_), .A1(new_n3745_), .B0(new_n3716_), .Y(new_n12418_));
  NAND2  g11416(.A(new_n12415_), .B(new_n12411_), .Y(new_n12419_));
  NAND2  g11417(.A(new_n12409_), .B(new_n12408_), .Y(new_n12420_));
  NAND4  g11418(.A(new_n12420_), .B(new_n12419_), .C(new_n12418_), .D(new_n3750_), .Y(new_n12421_));
  NAND2  g11419(.A(new_n12421_), .B(new_n12417_), .Y(new_n12422_));
  OAI21  g11420(.A0(new_n3796_), .A1(new_n3819_), .B0(new_n3773_), .Y(new_n12423_));
  OAI21  g11421(.A0(new_n3795_), .A1(new_n3805_), .B0(new_n3793_), .Y(new_n12424_));
  AOI21  g11422(.A0(new_n3803_), .A1(new_n3754_), .B0(new_n3802_), .Y(new_n12425_));
  NAND2  g11423(.A(new_n12425_), .B(new_n12424_), .Y(new_n12426_));
  AOI21  g11424(.A0(new_n3809_), .A1(new_n3774_), .B0(new_n3808_), .Y(new_n12427_));
  OAI21  g11425(.A0(new_n3772_), .A1(new_n3799_), .B0(new_n3770_), .Y(new_n12428_));
  NAND2  g11426(.A(new_n12428_), .B(new_n12427_), .Y(new_n12429_));
  AOI22  g11427(.A0(new_n12429_), .A1(new_n12426_), .B0(new_n12423_), .B1(new_n3814_), .Y(new_n12430_));
  NOR2   g11428(.A(new_n3823_), .B(new_n3822_), .Y(new_n12431_));
  AOI21  g11429(.A0(new_n3810_), .A1(new_n3789_), .B0(new_n3804_), .Y(new_n12432_));
  NOR2   g11430(.A(new_n12428_), .B(new_n12427_), .Y(new_n12433_));
  NOR2   g11431(.A(new_n12425_), .B(new_n12424_), .Y(new_n12434_));
  NOR4   g11432(.A(new_n12434_), .B(new_n12433_), .C(new_n12432_), .D(new_n12431_), .Y(new_n12435_));
  NOR2   g11433(.A(new_n12435_), .B(new_n12430_), .Y(new_n12436_));
  XOR2   g11434(.A(new_n12436_), .B(new_n12422_), .Y(new_n12437_));
  XOR2   g11435(.A(new_n12437_), .B(new_n12402_), .Y(new_n12438_));
  OAI22  g11436(.A0(new_n3688_), .A1(new_n3684_), .B0(new_n3834_), .B1(new_n3677_), .Y(new_n12439_));
  XOR2   g11437(.A(new_n3598_), .B(new_n3607_), .Y(new_n12440_));
  NAND4  g11438(.A(new_n3558_), .B(new_n3591_), .C(new_n12440_), .D(new_n3578_), .Y(new_n12441_));
  AOI211 g11439(.A0(new_n3597_), .A1(new_n3578_), .B(new_n12441_), .C(new_n3605_), .Y(new_n12442_));
  OAI21  g11440(.A0(new_n3609_), .A1(new_n3602_), .B0(new_n12440_), .Y(new_n12443_));
  AOI221 g11441(.A0(new_n12443_), .A1(new_n3593_), .C0(new_n3576_), .B0(new_n3574_), .B1(new_n3558_), .Y(new_n12444_));
  OAI21  g11442(.A0(new_n3599_), .A1(new_n3602_), .B0(new_n3597_), .Y(new_n12445_));
  OAI21  g11443(.A0(new_n3576_), .A1(new_n3604_), .B0(new_n3574_), .Y(new_n12446_));
  XOR2   g11444(.A(new_n12446_), .B(new_n12445_), .Y(new_n12447_));
  OAI21  g11445(.A0(new_n12444_), .A1(new_n12442_), .B0(new_n12447_), .Y(new_n12448_));
  OAI21  g11446(.A0(new_n3600_), .A1(new_n3606_), .B0(new_n3577_), .Y(new_n12449_));
  XOR2   g11447(.A(new_n3456_), .B(new_n3454_), .Y(new_n12450_));
  NAND2  g11448(.A(new_n3575_), .B(new_n12450_), .Y(new_n12451_));
  XOR2   g11449(.A(new_n3575_), .B(new_n12450_), .Y(new_n12452_));
  AOI22  g11450(.A0(new_n12452_), .A1(new_n3558_), .B0(new_n3573_), .B1(new_n12451_), .Y(new_n12453_));
  NAND2  g11451(.A(new_n12453_), .B(new_n12445_), .Y(new_n12454_));
  AOI21  g11452(.A0(new_n12440_), .A1(new_n3578_), .B0(new_n3609_), .Y(new_n12455_));
  NAND2  g11453(.A(new_n12446_), .B(new_n12455_), .Y(new_n12456_));
  NAND4  g11454(.A(new_n12456_), .B(new_n12454_), .C(new_n12449_), .D(new_n3611_), .Y(new_n12457_));
  NAND2  g11455(.A(new_n12457_), .B(new_n12448_), .Y(new_n12458_));
  NOR4   g11456(.A(new_n3619_), .B(new_n3631_), .C(new_n3648_), .D(new_n3630_), .Y(new_n12459_));
  OAI211 g11457(.A0(new_n3672_), .A1(new_n3630_), .B0(new_n12459_), .B1(new_n3673_), .Y(new_n12460_));
  OAI21  g11458(.A0(new_n3649_), .A1(new_n3633_), .B0(new_n3666_), .Y(new_n12461_));
  OAI21  g11459(.A0(new_n3648_), .A1(new_n3630_), .B0(new_n3646_), .Y(new_n12462_));
  AOI21  g11460(.A0(new_n3624_), .A1(new_n3652_), .B0(new_n3623_), .Y(new_n12463_));
  NAND2  g11461(.A(new_n12463_), .B(new_n12462_), .Y(new_n12464_));
  AOI21  g11462(.A0(new_n3668_), .A1(new_n3634_), .B0(new_n3672_), .Y(new_n12465_));
  OAI21  g11463(.A0(new_n3665_), .A1(new_n3619_), .B0(new_n3664_), .Y(new_n12466_));
  NAND2  g11464(.A(new_n12466_), .B(new_n12465_), .Y(new_n12467_));
  AOI22  g11465(.A0(new_n12467_), .A1(new_n12464_), .B0(new_n12461_), .B1(new_n12460_), .Y(new_n12468_));
  OAI21  g11466(.A0(new_n3672_), .A1(new_n3630_), .B0(new_n3668_), .Y(new_n12469_));
  AOI21  g11467(.A0(new_n12469_), .A1(new_n3685_), .B0(new_n3625_), .Y(new_n12470_));
  OAI22  g11468(.A0(new_n12466_), .A1(new_n12465_), .B0(new_n3674_), .B1(new_n3670_), .Y(new_n12471_));
  AOI211 g11469(.A0(new_n12466_), .A1(new_n12465_), .B(new_n12471_), .C(new_n12470_), .Y(new_n12472_));
  NOR2   g11470(.A(new_n12472_), .B(new_n12468_), .Y(new_n12473_));
  XOR2   g11471(.A(new_n12473_), .B(new_n12458_), .Y(new_n12474_));
  XOR2   g11472(.A(new_n12474_), .B(new_n12439_), .Y(new_n12475_));
  XOR2   g11473(.A(new_n12475_), .B(new_n12438_), .Y(new_n12476_));
  XOR2   g11474(.A(new_n12476_), .B(new_n12398_), .Y(new_n12477_));
  OAI21  g11475(.A0(new_n4141_), .A1(new_n4129_), .B0(new_n4133_), .Y(new_n12478_));
  AOI21  g11476(.A0(new_n3900_), .A1(new_n3863_), .B0(new_n3888_), .Y(new_n12479_));
  OAI22  g11477(.A0(new_n3970_), .A1(new_n3968_), .B0(new_n12479_), .B1(new_n3901_), .Y(new_n12480_));
  NAND4  g11478(.A(new_n3913_), .B(new_n3937_), .C(new_n3962_), .D(new_n3924_), .Y(new_n12481_));
  AOI221 g11479(.A0(new_n3956_), .A1(new_n3917_), .C0(new_n12481_), .B0(new_n3945_), .B1(new_n3924_), .Y(new_n12482_));
  AOI21  g11480(.A0(new_n3963_), .A1(new_n3941_), .B0(new_n3957_), .Y(new_n12483_));
  AOI21  g11481(.A0(new_n3962_), .A1(new_n3924_), .B0(new_n3961_), .Y(new_n12484_));
  AOI211 g11482(.A0(new_n3956_), .A1(new_n3913_), .B(new_n12484_), .C(new_n3955_), .Y(new_n12485_));
  OAI21  g11483(.A0(new_n3947_), .A1(new_n3958_), .B0(new_n3945_), .Y(new_n12486_));
  AOI21  g11484(.A0(new_n3956_), .A1(new_n3913_), .B0(new_n3955_), .Y(new_n12487_));
  NOR2   g11485(.A(new_n12487_), .B(new_n12486_), .Y(new_n12488_));
  OAI22  g11486(.A0(new_n12488_), .A1(new_n12485_), .B0(new_n12483_), .B1(new_n12482_), .Y(new_n12489_));
  NAND2  g11487(.A(new_n3964_), .B(new_n3923_), .Y(new_n12490_));
  NAND2  g11488(.A(new_n12487_), .B(new_n12486_), .Y(new_n12491_));
  OAI21  g11489(.A0(new_n3922_), .A1(new_n3953_), .B0(new_n3917_), .Y(new_n12492_));
  NAND2  g11490(.A(new_n12492_), .B(new_n12484_), .Y(new_n12493_));
  NAND4  g11491(.A(new_n12493_), .B(new_n12491_), .C(new_n12490_), .D(new_n3966_), .Y(new_n12494_));
  NAND2  g11492(.A(new_n12494_), .B(new_n12489_), .Y(new_n12495_));
  NOR4   g11493(.A(new_n3891_), .B(new_n3890_), .C(new_n3885_), .D(new_n3889_), .Y(new_n12496_));
  OAI211 g11494(.A0(new_n3898_), .A1(new_n3889_), .B0(new_n12496_), .B1(new_n3878_), .Y(new_n12497_));
  OAI21  g11495(.A0(new_n3886_), .A1(new_n3893_), .B0(new_n3863_), .Y(new_n12498_));
  OAI21  g11496(.A0(new_n3885_), .A1(new_n3889_), .B0(new_n3883_), .Y(new_n12499_));
  AOI21  g11497(.A0(new_n3906_), .A1(new_n3844_), .B0(new_n3905_), .Y(new_n12500_));
  NAND2  g11498(.A(new_n12500_), .B(new_n12499_), .Y(new_n12501_));
  AOI21  g11499(.A0(new_n3895_), .A1(new_n3864_), .B0(new_n3898_), .Y(new_n12502_));
  OAI21  g11500(.A0(new_n3862_), .A1(new_n3891_), .B0(new_n3860_), .Y(new_n12503_));
  NAND2  g11501(.A(new_n12503_), .B(new_n12502_), .Y(new_n12504_));
  AOI22  g11502(.A0(new_n12504_), .A1(new_n12501_), .B0(new_n12498_), .B1(new_n12497_), .Y(new_n12505_));
  NOR2   g11503(.A(new_n3899_), .B(new_n3896_), .Y(new_n12506_));
  OAI21  g11504(.A0(new_n3898_), .A1(new_n3889_), .B0(new_n3895_), .Y(new_n12507_));
  AOI21  g11505(.A0(new_n12507_), .A1(new_n3879_), .B0(new_n3907_), .Y(new_n12508_));
  NOR2   g11506(.A(new_n12503_), .B(new_n12502_), .Y(new_n12509_));
  NOR2   g11507(.A(new_n12500_), .B(new_n12499_), .Y(new_n12510_));
  NOR4   g11508(.A(new_n12510_), .B(new_n12509_), .C(new_n12508_), .D(new_n12506_), .Y(new_n12511_));
  NOR2   g11509(.A(new_n12511_), .B(new_n12505_), .Y(new_n12512_));
  XOR2   g11510(.A(new_n12512_), .B(new_n12495_), .Y(new_n12513_));
  XOR2   g11511(.A(new_n12513_), .B(new_n12480_), .Y(new_n12514_));
  OAI22  g11512(.A0(new_n4100_), .A1(new_n4029_), .B0(new_n4097_), .B1(new_n4030_), .Y(new_n12515_));
  NAND4  g11513(.A(new_n3974_), .B(new_n3998_), .C(new_n4023_), .D(new_n3985_), .Y(new_n12516_));
  AOI221 g11514(.A0(new_n4017_), .A1(new_n3978_), .C0(new_n12516_), .B0(new_n4006_), .B1(new_n3985_), .Y(new_n12517_));
  AOI21  g11515(.A0(new_n4024_), .A1(new_n4002_), .B0(new_n4018_), .Y(new_n12518_));
  AOI21  g11516(.A0(new_n4023_), .A1(new_n3985_), .B0(new_n4022_), .Y(new_n12519_));
  AOI211 g11517(.A0(new_n4017_), .A1(new_n3974_), .B(new_n12519_), .C(new_n4016_), .Y(new_n12520_));
  OAI21  g11518(.A0(new_n4008_), .A1(new_n4019_), .B0(new_n4006_), .Y(new_n12521_));
  AOI21  g11519(.A0(new_n4017_), .A1(new_n3974_), .B0(new_n4016_), .Y(new_n12522_));
  NOR2   g11520(.A(new_n12522_), .B(new_n12521_), .Y(new_n12523_));
  OAI22  g11521(.A0(new_n12523_), .A1(new_n12520_), .B0(new_n12518_), .B1(new_n12517_), .Y(new_n12524_));
  NAND2  g11522(.A(new_n4025_), .B(new_n3984_), .Y(new_n12525_));
  NAND2  g11523(.A(new_n12522_), .B(new_n12521_), .Y(new_n12526_));
  OAI21  g11524(.A0(new_n3983_), .A1(new_n4014_), .B0(new_n3978_), .Y(new_n12527_));
  NAND2  g11525(.A(new_n12527_), .B(new_n12519_), .Y(new_n12528_));
  NAND4  g11526(.A(new_n12528_), .B(new_n12526_), .C(new_n12525_), .D(new_n4027_), .Y(new_n12529_));
  NAND2  g11527(.A(new_n12529_), .B(new_n12524_), .Y(new_n12530_));
  NOR4   g11528(.A(new_n4036_), .B(new_n4048_), .C(new_n4065_), .D(new_n4047_), .Y(new_n12531_));
  OAI211 g11529(.A0(new_n4088_), .A1(new_n4047_), .B0(new_n12531_), .B1(new_n4089_), .Y(new_n12532_));
  OAI21  g11530(.A0(new_n4066_), .A1(new_n4050_), .B0(new_n4082_), .Y(new_n12533_));
  OAI21  g11531(.A0(new_n4065_), .A1(new_n4047_), .B0(new_n4063_), .Y(new_n12534_));
  AOI21  g11532(.A0(new_n4041_), .A1(new_n4069_), .B0(new_n4040_), .Y(new_n12535_));
  NAND2  g11533(.A(new_n12535_), .B(new_n12534_), .Y(new_n12536_));
  AOI21  g11534(.A0(new_n4084_), .A1(new_n4051_), .B0(new_n4088_), .Y(new_n12537_));
  OAI21  g11535(.A0(new_n4081_), .A1(new_n4036_), .B0(new_n4080_), .Y(new_n12538_));
  NAND2  g11536(.A(new_n12538_), .B(new_n12537_), .Y(new_n12539_));
  AOI22  g11537(.A0(new_n12539_), .A1(new_n12536_), .B0(new_n12533_), .B1(new_n12532_), .Y(new_n12540_));
  NOR2   g11538(.A(new_n4108_), .B(new_n4042_), .Y(new_n12541_));
  NOR2   g11539(.A(new_n12538_), .B(new_n12537_), .Y(new_n12542_));
  NOR2   g11540(.A(new_n12535_), .B(new_n12534_), .Y(new_n12543_));
  NOR4   g11541(.A(new_n12543_), .B(new_n12542_), .C(new_n12541_), .D(new_n4109_), .Y(new_n12544_));
  NOR2   g11542(.A(new_n12544_), .B(new_n12540_), .Y(new_n12545_));
  XOR2   g11543(.A(new_n12545_), .B(new_n12530_), .Y(new_n12546_));
  XOR2   g11544(.A(new_n12546_), .B(new_n12515_), .Y(new_n12547_));
  XOR2   g11545(.A(new_n12547_), .B(new_n12514_), .Y(new_n12548_));
  XOR2   g11546(.A(new_n12548_), .B(new_n12478_), .Y(new_n12549_));
  XOR2   g11547(.A(new_n12549_), .B(new_n12477_), .Y(new_n12550_));
  XOR2   g11548(.A(new_n12550_), .B(new_n12397_), .Y(new_n12551_));
  XOR2   g11549(.A(new_n12551_), .B(new_n12396_), .Y(new_n12552_));
  XOR2   g11550(.A(new_n12552_), .B(new_n12241_), .Y(new_n12553_));
  OAI21  g11551(.A0(new_n2874_), .A1(new_n1929_), .B0(new_n3553_), .Y(new_n12554_));
  OAI21  g11552(.A0(new_n2870_), .A1(new_n1925_), .B0(new_n1927_), .Y(new_n12555_));
  OAI21  g11553(.A0(new_n1913_), .A1(new_n1767_), .B0(new_n1923_), .Y(new_n12556_));
  NOR2   g11554(.A(new_n1674_), .B(new_n1650_), .Y(new_n12557_));
  AOI21  g11555(.A0(new_n1685_), .A1(new_n1650_), .B0(new_n12557_), .Y(new_n12558_));
  NOR3   g11556(.A(new_n1760_), .B(new_n1749_), .C(new_n1732_), .Y(new_n12559_));
  OAI22  g11557(.A0(new_n12559_), .A1(new_n12558_), .B0(new_n1764_), .B1(new_n1750_), .Y(new_n12560_));
  XOR2   g11558(.A(new_n1671_), .B(new_n1680_), .Y(new_n12561_));
  NAND4  g11559(.A(new_n1631_), .B(new_n1664_), .C(new_n12561_), .D(new_n1651_), .Y(new_n12562_));
  AOI211 g11560(.A0(new_n1670_), .A1(new_n1651_), .B(new_n12562_), .C(new_n1678_), .Y(new_n12563_));
  OAI21  g11561(.A0(new_n1682_), .A1(new_n1675_), .B0(new_n12561_), .Y(new_n12564_));
  AOI221 g11562(.A0(new_n12564_), .A1(new_n1666_), .C0(new_n1649_), .B0(new_n1647_), .B1(new_n1631_), .Y(new_n12565_));
  AOI21  g11563(.A0(new_n12561_), .A1(new_n1651_), .B0(new_n1682_), .Y(new_n12566_));
  OAI21  g11564(.A0(new_n1649_), .A1(new_n1677_), .B0(new_n1647_), .Y(new_n12567_));
  NOR2   g11565(.A(new_n12567_), .B(new_n12566_), .Y(new_n12568_));
  OAI21  g11566(.A0(new_n1672_), .A1(new_n1675_), .B0(new_n1670_), .Y(new_n12569_));
  XOR2   g11567(.A(new_n1615_), .B(new_n1613_), .Y(new_n12570_));
  NAND2  g11568(.A(new_n1648_), .B(new_n12570_), .Y(new_n12571_));
  XOR2   g11569(.A(new_n1648_), .B(new_n12570_), .Y(new_n12572_));
  AOI22  g11570(.A0(new_n12572_), .A1(new_n1631_), .B0(new_n1646_), .B1(new_n12571_), .Y(new_n12573_));
  NOR2   g11571(.A(new_n12573_), .B(new_n12569_), .Y(new_n12574_));
  OAI22  g11572(.A0(new_n12574_), .A1(new_n12568_), .B0(new_n12565_), .B1(new_n12563_), .Y(new_n12575_));
  OAI21  g11573(.A0(new_n1673_), .A1(new_n1679_), .B0(new_n1650_), .Y(new_n12576_));
  NAND2  g11574(.A(new_n12573_), .B(new_n12569_), .Y(new_n12577_));
  NAND2  g11575(.A(new_n12567_), .B(new_n12566_), .Y(new_n12578_));
  NAND4  g11576(.A(new_n12578_), .B(new_n12577_), .C(new_n12576_), .D(new_n1684_), .Y(new_n12579_));
  NAND2  g11577(.A(new_n12579_), .B(new_n12575_), .Y(new_n12580_));
  OAI21  g11578(.A0(new_n1730_), .A1(new_n1753_), .B0(new_n1707_), .Y(new_n12581_));
  OAI21  g11579(.A0(new_n1729_), .A1(new_n1739_), .B0(new_n1727_), .Y(new_n12582_));
  AOI21  g11580(.A0(new_n1737_), .A1(new_n1688_), .B0(new_n1736_), .Y(new_n12583_));
  NAND2  g11581(.A(new_n12583_), .B(new_n12582_), .Y(new_n12584_));
  AOI21  g11582(.A0(new_n1743_), .A1(new_n1708_), .B0(new_n1742_), .Y(new_n12585_));
  OAI21  g11583(.A0(new_n1706_), .A1(new_n1733_), .B0(new_n1704_), .Y(new_n12586_));
  NAND2  g11584(.A(new_n12586_), .B(new_n12585_), .Y(new_n12587_));
  AOI22  g11585(.A0(new_n12587_), .A1(new_n12584_), .B0(new_n12581_), .B1(new_n1748_), .Y(new_n12588_));
  NOR2   g11586(.A(new_n1757_), .B(new_n1756_), .Y(new_n12589_));
  AOI21  g11587(.A0(new_n1744_), .A1(new_n1723_), .B0(new_n1738_), .Y(new_n12590_));
  NOR2   g11588(.A(new_n12586_), .B(new_n12585_), .Y(new_n12591_));
  NOR2   g11589(.A(new_n12583_), .B(new_n12582_), .Y(new_n12592_));
  NOR4   g11590(.A(new_n12592_), .B(new_n12591_), .C(new_n12590_), .D(new_n12589_), .Y(new_n12593_));
  NOR2   g11591(.A(new_n12593_), .B(new_n12588_), .Y(new_n12594_));
  XOR2   g11592(.A(new_n12594_), .B(new_n12580_), .Y(new_n12595_));
  XOR2   g11593(.A(new_n12595_), .B(new_n12560_), .Y(new_n12596_));
  OAI22  g11594(.A0(new_n1898_), .A1(new_n1894_), .B0(new_n1904_), .B1(new_n1887_), .Y(new_n12597_));
  XOR2   g11595(.A(new_n1808_), .B(new_n1817_), .Y(new_n12598_));
  NAND4  g11596(.A(new_n1768_), .B(new_n1801_), .C(new_n12598_), .D(new_n1788_), .Y(new_n12599_));
  AOI211 g11597(.A0(new_n1807_), .A1(new_n1788_), .B(new_n12599_), .C(new_n1815_), .Y(new_n12600_));
  OAI21  g11598(.A0(new_n1819_), .A1(new_n1812_), .B0(new_n12598_), .Y(new_n12601_));
  AOI221 g11599(.A0(new_n12601_), .A1(new_n1803_), .C0(new_n1786_), .B0(new_n1784_), .B1(new_n1768_), .Y(new_n12602_));
  OAI21  g11600(.A0(new_n1809_), .A1(new_n1812_), .B0(new_n1807_), .Y(new_n12603_));
  OAI21  g11601(.A0(new_n1786_), .A1(new_n1814_), .B0(new_n1784_), .Y(new_n12604_));
  XOR2   g11602(.A(new_n12604_), .B(new_n12603_), .Y(new_n12605_));
  OAI21  g11603(.A0(new_n12602_), .A1(new_n12600_), .B0(new_n12605_), .Y(new_n12606_));
  OAI21  g11604(.A0(new_n1810_), .A1(new_n1816_), .B0(new_n1787_), .Y(new_n12607_));
  XOR2   g11605(.A(new_n1534_), .B(new_n1532_), .Y(new_n12608_));
  NAND2  g11606(.A(new_n1785_), .B(new_n12608_), .Y(new_n12609_));
  XOR2   g11607(.A(new_n1785_), .B(new_n12608_), .Y(new_n12610_));
  AOI22  g11608(.A0(new_n12610_), .A1(new_n1768_), .B0(new_n1783_), .B1(new_n12609_), .Y(new_n12611_));
  NAND2  g11609(.A(new_n12611_), .B(new_n12603_), .Y(new_n12612_));
  AOI21  g11610(.A0(new_n12598_), .A1(new_n1788_), .B0(new_n1819_), .Y(new_n12613_));
  NAND2  g11611(.A(new_n12604_), .B(new_n12613_), .Y(new_n12614_));
  NAND4  g11612(.A(new_n12614_), .B(new_n12612_), .C(new_n12607_), .D(new_n1821_), .Y(new_n12615_));
  NAND2  g11613(.A(new_n12615_), .B(new_n12606_), .Y(new_n12616_));
  NOR4   g11614(.A(new_n1829_), .B(new_n1841_), .C(new_n1858_), .D(new_n1840_), .Y(new_n12617_));
  OAI211 g11615(.A0(new_n1882_), .A1(new_n1840_), .B0(new_n12617_), .B1(new_n1883_), .Y(new_n12618_));
  OAI21  g11616(.A0(new_n1859_), .A1(new_n1843_), .B0(new_n1876_), .Y(new_n12619_));
  OAI21  g11617(.A0(new_n1858_), .A1(new_n1840_), .B0(new_n1856_), .Y(new_n12620_));
  AOI21  g11618(.A0(new_n1834_), .A1(new_n1862_), .B0(new_n1833_), .Y(new_n12621_));
  NAND2  g11619(.A(new_n12621_), .B(new_n12620_), .Y(new_n12622_));
  AOI21  g11620(.A0(new_n1878_), .A1(new_n1844_), .B0(new_n1882_), .Y(new_n12623_));
  OAI21  g11621(.A0(new_n1875_), .A1(new_n1829_), .B0(new_n1874_), .Y(new_n12624_));
  NAND2  g11622(.A(new_n12624_), .B(new_n12623_), .Y(new_n12625_));
  AOI22  g11623(.A0(new_n12625_), .A1(new_n12622_), .B0(new_n12619_), .B1(new_n12618_), .Y(new_n12626_));
  OAI21  g11624(.A0(new_n1882_), .A1(new_n1840_), .B0(new_n1878_), .Y(new_n12627_));
  AOI21  g11625(.A0(new_n12627_), .A1(new_n1895_), .B0(new_n1835_), .Y(new_n12628_));
  OAI22  g11626(.A0(new_n12624_), .A1(new_n12623_), .B0(new_n1884_), .B1(new_n1880_), .Y(new_n12629_));
  AOI211 g11627(.A0(new_n12624_), .A1(new_n12623_), .B(new_n12629_), .C(new_n12628_), .Y(new_n12630_));
  NOR2   g11628(.A(new_n12630_), .B(new_n12626_), .Y(new_n12631_));
  XOR2   g11629(.A(new_n12631_), .B(new_n12616_), .Y(new_n12632_));
  XOR2   g11630(.A(new_n12632_), .B(new_n12597_), .Y(new_n12633_));
  XOR2   g11631(.A(new_n12633_), .B(new_n12596_), .Y(new_n12634_));
  XOR2   g11632(.A(new_n12634_), .B(new_n12556_), .Y(new_n12635_));
  AOI21  g11633(.A0(new_n1452_), .A1(new_n1448_), .B0(new_n1454_), .Y(new_n12636_));
  NOR2   g11634(.A(new_n12636_), .B(new_n1455_), .Y(new_n12637_));
  OAI22  g11635(.A0(new_n1449_), .A1(new_n1080_), .B0(new_n1214_), .B1(new_n1209_), .Y(new_n12638_));
  NAND2  g11636(.A(new_n12638_), .B(new_n1217_), .Y(new_n12639_));
  NAND4  g11637(.A(new_n1156_), .B(new_n1180_), .C(new_n1197_), .D(new_n1167_), .Y(new_n12640_));
  AOI221 g11638(.A0(new_n1212_), .A1(new_n1160_), .C0(new_n12640_), .B0(new_n1188_), .B1(new_n1167_), .Y(new_n12641_));
  AOI21  g11639(.A0(new_n1198_), .A1(new_n1184_), .B0(new_n1213_), .Y(new_n12642_));
  AOI21  g11640(.A0(new_n1197_), .A1(new_n1167_), .B0(new_n1196_), .Y(new_n12643_));
  AOI211 g11641(.A0(new_n1212_), .A1(new_n1156_), .B(new_n12643_), .C(new_n1211_), .Y(new_n12644_));
  OAI21  g11642(.A0(new_n1190_), .A1(new_n1193_), .B0(new_n1188_), .Y(new_n12645_));
  AOI21  g11643(.A0(new_n1212_), .A1(new_n1156_), .B0(new_n1211_), .Y(new_n12646_));
  NOR2   g11644(.A(new_n12646_), .B(new_n12645_), .Y(new_n12647_));
  OAI22  g11645(.A0(new_n12647_), .A1(new_n12644_), .B0(new_n12642_), .B1(new_n12641_), .Y(new_n12648_));
  NAND2  g11646(.A(new_n1199_), .B(new_n1166_), .Y(new_n12649_));
  NAND2  g11647(.A(new_n12646_), .B(new_n12645_), .Y(new_n12650_));
  OAI21  g11648(.A0(new_n1165_), .A1(new_n1202_), .B0(new_n1160_), .Y(new_n12651_));
  NAND2  g11649(.A(new_n12651_), .B(new_n12643_), .Y(new_n12652_));
  NAND4  g11650(.A(new_n12652_), .B(new_n12650_), .C(new_n12649_), .D(new_n1204_), .Y(new_n12653_));
  NAND2  g11651(.A(new_n12653_), .B(new_n12648_), .Y(new_n12654_));
  NOR3   g11652(.A(new_n1095_), .B(new_n1094_), .C(new_n1077_), .Y(new_n12655_));
  OAI211 g11653(.A0(new_n1092_), .A1(new_n1090_), .B0(new_n12655_), .B1(new_n1060_), .Y(new_n12656_));
  OAI21  g11654(.A0(new_n1078_), .A1(new_n1145_), .B0(new_n1039_), .Y(new_n12657_));
  OAI21  g11655(.A0(new_n1092_), .A1(new_n1077_), .B0(new_n1075_), .Y(new_n12658_));
  OAI211 g11656(.A0(new_n1082_), .A1(new_n1024_), .B0(new_n12658_), .B1(new_n1038_), .Y(new_n12659_));
  AOI21  g11657(.A0(new_n1068_), .A1(new_n1091_), .B0(new_n1090_), .Y(new_n12660_));
  OAI21  g11658(.A0(new_n1082_), .A1(new_n1024_), .B0(new_n1038_), .Y(new_n12661_));
  NAND2  g11659(.A(new_n12661_), .B(new_n12660_), .Y(new_n12662_));
  AOI22  g11660(.A0(new_n12662_), .A1(new_n12659_), .B0(new_n12657_), .B1(new_n12656_), .Y(new_n12663_));
  AOI221 g11661(.A0(new_n1093_), .A1(new_n1069_), .C0(new_n1024_), .B0(new_n1038_), .B1(new_n1025_), .Y(new_n12664_));
  NOR2   g11662(.A(new_n12661_), .B(new_n12660_), .Y(new_n12665_));
  AOI21  g11663(.A0(new_n1025_), .A1(new_n1081_), .B0(new_n1084_), .Y(new_n12666_));
  NOR2   g11664(.A(new_n12666_), .B(new_n12658_), .Y(new_n12667_));
  NOR4   g11665(.A(new_n12667_), .B(new_n12665_), .C(new_n12664_), .D(new_n1097_), .Y(new_n12668_));
  NOR2   g11666(.A(new_n12668_), .B(new_n12663_), .Y(new_n12669_));
  XOR2   g11667(.A(new_n12669_), .B(new_n12654_), .Y(new_n12670_));
  XOR2   g11668(.A(new_n12670_), .B(new_n12639_), .Y(new_n12671_));
  OAI21  g11669(.A0(new_n1418_), .A1(new_n1344_), .B0(new_n1423_), .Y(new_n12672_));
  OAI22  g11670(.A0(new_n12672_), .A1(new_n1412_), .B0(new_n1432_), .B1(new_n1426_), .Y(new_n12673_));
  NAND2  g11671(.A(new_n12673_), .B(new_n1435_), .Y(new_n12674_));
  AOI221 g11672(.A0(new_n1430_), .A1(new_n1287_), .C0(new_n1241_), .B0(new_n1255_), .B1(new_n1242_), .Y(new_n12675_));
  AOI21  g11673(.A0(new_n1286_), .A1(new_n1299_), .B0(new_n1428_), .Y(new_n12676_));
  XOR2   g11674(.A(new_n1233_), .B(new_n1246_), .Y(new_n12677_));
  OAI21  g11675(.A0(new_n12677_), .A1(new_n1241_), .B0(new_n1255_), .Y(new_n12678_));
  NOR2   g11676(.A(new_n12678_), .B(new_n12676_), .Y(new_n12679_));
  OAI21  g11677(.A0(new_n1429_), .A1(new_n1295_), .B0(new_n1293_), .Y(new_n12680_));
  XOR2   g11678(.A(new_n1240_), .B(new_n1251_), .Y(new_n12681_));
  XOR2   g11679(.A(new_n1253_), .B(new_n1237_), .Y(new_n12682_));
  NAND2  g11680(.A(new_n12682_), .B(new_n1234_), .Y(new_n12683_));
  AOI22  g11681(.A0(new_n1254_), .A1(new_n12683_), .B0(new_n1242_), .B1(new_n12681_), .Y(new_n12684_));
  NOR2   g11682(.A(new_n12684_), .B(new_n12680_), .Y(new_n12685_));
  OAI22  g11683(.A0(new_n12685_), .A1(new_n12679_), .B0(new_n12675_), .B1(new_n1305_), .Y(new_n12686_));
  NOR3   g11684(.A(new_n1301_), .B(new_n1300_), .C(new_n1295_), .Y(new_n12687_));
  OAI211 g11685(.A0(new_n1429_), .A1(new_n1428_), .B0(new_n12687_), .B1(new_n1278_), .Y(new_n12688_));
  OAI21  g11686(.A0(new_n1296_), .A1(new_n1302_), .B0(new_n1256_), .Y(new_n12689_));
  NAND2  g11687(.A(new_n12684_), .B(new_n12680_), .Y(new_n12690_));
  NAND2  g11688(.A(new_n12678_), .B(new_n12676_), .Y(new_n12691_));
  NAND4  g11689(.A(new_n12691_), .B(new_n12690_), .C(new_n12689_), .D(new_n12688_), .Y(new_n12692_));
  NAND2  g11690(.A(new_n12692_), .B(new_n12686_), .Y(new_n12693_));
  AOI221 g11691(.A0(new_n1417_), .A1(new_n1410_), .C0(new_n1390_), .B0(new_n1392_), .B1(new_n1338_), .Y(new_n12694_));
  AOI21  g11692(.A0(new_n1365_), .A1(new_n1416_), .B0(new_n1415_), .Y(new_n12695_));
  OAI21  g11693(.A0(new_n1339_), .A1(new_n1390_), .B0(new_n1392_), .Y(new_n12696_));
  NOR2   g11694(.A(new_n12696_), .B(new_n12695_), .Y(new_n12697_));
  OAI21  g11695(.A0(new_n1398_), .A1(new_n1385_), .B0(new_n1383_), .Y(new_n12698_));
  NAND2  g11696(.A(new_n1338_), .B(new_n1329_), .Y(new_n12699_));
  AOI21  g11697(.A0(new_n12699_), .A1(new_n1392_), .B0(new_n12698_), .Y(new_n12700_));
  OAI22  g11698(.A0(new_n12700_), .A1(new_n12697_), .B0(new_n12694_), .B1(new_n1396_), .Y(new_n12701_));
  NOR3   g11699(.A(new_n1366_), .B(new_n1364_), .C(new_n1385_), .Y(new_n12702_));
  OAI211 g11700(.A0(new_n1398_), .A1(new_n1415_), .B0(new_n12702_), .B1(new_n1409_), .Y(new_n12703_));
  OAI21  g11701(.A0(new_n1386_), .A1(new_n1367_), .B0(new_n1393_), .Y(new_n12704_));
  OAI211 g11702(.A0(new_n1339_), .A1(new_n1390_), .B0(new_n12698_), .B1(new_n1392_), .Y(new_n12705_));
  NAND2  g11703(.A(new_n12696_), .B(new_n12695_), .Y(new_n12706_));
  NAND4  g11704(.A(new_n12706_), .B(new_n12705_), .C(new_n12704_), .D(new_n12703_), .Y(new_n12707_));
  NAND2  g11705(.A(new_n12707_), .B(new_n12701_), .Y(new_n12708_));
  XOR2   g11706(.A(new_n12708_), .B(new_n12693_), .Y(new_n12709_));
  XOR2   g11707(.A(new_n12709_), .B(new_n12674_), .Y(new_n12710_));
  XOR2   g11708(.A(new_n12710_), .B(new_n12671_), .Y(new_n12711_));
  XOR2   g11709(.A(new_n12711_), .B(new_n12637_), .Y(new_n12712_));
  XOR2   g11710(.A(new_n12712_), .B(new_n12635_), .Y(new_n12713_));
  XOR2   g11711(.A(new_n12713_), .B(new_n12555_), .Y(new_n12714_));
  OAI21  g11712(.A0(new_n2862_), .A1(new_n2849_), .B0(new_n2851_), .Y(new_n12715_));
  OAI21  g11713(.A0(new_n2369_), .A1(new_n2144_), .B0(new_n2847_), .Y(new_n12716_));
  NOR2   g11714(.A(new_n2005_), .B(new_n1965_), .Y(new_n12717_));
  AOI21  g11715(.A0(new_n2020_), .A1(new_n1965_), .B0(new_n12717_), .Y(new_n12718_));
  NOR3   g11716(.A(new_n2137_), .B(new_n2120_), .C(new_n2099_), .Y(new_n12719_));
  OAI22  g11717(.A0(new_n12719_), .A1(new_n12718_), .B0(new_n2141_), .B1(new_n2127_), .Y(new_n12720_));
  XOR2   g11718(.A(new_n2002_), .B(new_n2015_), .Y(new_n12721_));
  NAND4  g11719(.A(new_n1944_), .B(new_n1993_), .C(new_n12721_), .D(new_n1980_), .Y(new_n12722_));
  AOI211 g11720(.A0(new_n2001_), .A1(new_n1980_), .B(new_n12722_), .C(new_n2013_), .Y(new_n12723_));
  OAI21  g11721(.A0(new_n2017_), .A1(new_n2006_), .B0(new_n12721_), .Y(new_n12724_));
  AOI221 g11722(.A0(new_n12724_), .A1(new_n1995_), .C0(new_n1964_), .B0(new_n1962_), .B1(new_n1944_), .Y(new_n12725_));
  AOI21  g11723(.A0(new_n12721_), .A1(new_n1980_), .B0(new_n2017_), .Y(new_n12726_));
  OAI21  g11724(.A0(new_n1964_), .A1(new_n2010_), .B0(new_n1962_), .Y(new_n12727_));
  NOR2   g11725(.A(new_n12727_), .B(new_n12726_), .Y(new_n12728_));
  OAI21  g11726(.A0(new_n2003_), .A1(new_n2006_), .B0(new_n2001_), .Y(new_n12729_));
  XOR2   g11727(.A(new_n1949_), .B(new_n2012_), .Y(new_n12730_));
  NAND2  g11728(.A(new_n1963_), .B(new_n12730_), .Y(new_n12731_));
  XOR2   g11729(.A(new_n1963_), .B(new_n12730_), .Y(new_n12732_));
  AOI22  g11730(.A0(new_n12732_), .A1(new_n1944_), .B0(new_n1961_), .B1(new_n12731_), .Y(new_n12733_));
  NOR2   g11731(.A(new_n12733_), .B(new_n12729_), .Y(new_n12734_));
  OAI22  g11732(.A0(new_n12734_), .A1(new_n12728_), .B0(new_n12725_), .B1(new_n12723_), .Y(new_n12735_));
  OAI21  g11733(.A0(new_n2004_), .A1(new_n2014_), .B0(new_n1965_), .Y(new_n12736_));
  NAND2  g11734(.A(new_n12733_), .B(new_n12729_), .Y(new_n12737_));
  NAND2  g11735(.A(new_n12727_), .B(new_n12726_), .Y(new_n12738_));
  NAND4  g11736(.A(new_n12738_), .B(new_n12737_), .C(new_n12736_), .D(new_n2019_), .Y(new_n12739_));
  NAND2  g11737(.A(new_n12739_), .B(new_n12735_), .Y(new_n12740_));
  OAI21  g11738(.A0(new_n2097_), .A1(new_n2130_), .B0(new_n2058_), .Y(new_n12741_));
  OAI21  g11739(.A0(new_n2096_), .A1(new_n2108_), .B0(new_n2094_), .Y(new_n12742_));
  AOI21  g11740(.A0(new_n2106_), .A1(new_n2037_), .B0(new_n2105_), .Y(new_n12743_));
  NAND2  g11741(.A(new_n12743_), .B(new_n12742_), .Y(new_n12744_));
  AOI21  g11742(.A0(new_n2114_), .A1(new_n2073_), .B0(new_n2113_), .Y(new_n12745_));
  OAI21  g11743(.A0(new_n2057_), .A1(new_n2100_), .B0(new_n2055_), .Y(new_n12746_));
  NAND2  g11744(.A(new_n12746_), .B(new_n12745_), .Y(new_n12747_));
  AOI22  g11745(.A0(new_n12747_), .A1(new_n12744_), .B0(new_n12741_), .B1(new_n2119_), .Y(new_n12748_));
  NOR2   g11746(.A(new_n2134_), .B(new_n2133_), .Y(new_n12749_));
  AOI21  g11747(.A0(new_n2115_), .A1(new_n2088_), .B0(new_n2107_), .Y(new_n12750_));
  NOR2   g11748(.A(new_n12746_), .B(new_n12745_), .Y(new_n12751_));
  NOR2   g11749(.A(new_n12743_), .B(new_n12742_), .Y(new_n12752_));
  NOR4   g11750(.A(new_n12752_), .B(new_n12751_), .C(new_n12750_), .D(new_n12749_), .Y(new_n12753_));
  NOR2   g11751(.A(new_n12753_), .B(new_n12748_), .Y(new_n12754_));
  XOR2   g11752(.A(new_n12754_), .B(new_n12740_), .Y(new_n12755_));
  XOR2   g11753(.A(new_n12755_), .B(new_n12720_), .Y(new_n12756_));
  NOR3   g11754(.A(new_n2336_), .B(new_n2348_), .C(new_n2341_), .Y(new_n12757_));
  OAI21  g11755(.A0(new_n12757_), .A1(new_n2356_), .B0(new_n2358_), .Y(new_n12758_));
  NOR3   g11756(.A(new_n2220_), .B(new_n2214_), .C(new_n2222_), .Y(new_n12759_));
  OAI211 g11757(.A0(new_n2231_), .A1(new_n2230_), .B0(new_n12759_), .B1(new_n2226_), .Y(new_n12760_));
  OAI221 g11758(.A0(new_n2223_), .A1(new_n2221_), .C0(new_n2166_), .B0(new_n2176_), .B1(new_n2171_), .Y(new_n12761_));
  NAND2  g11759(.A(new_n12761_), .B(new_n12760_), .Y(new_n12762_));
  AOI21  g11760(.A0(new_n2219_), .A1(new_n2213_), .B0(new_n2230_), .Y(new_n12763_));
  NOR2   g11761(.A(new_n2170_), .B(new_n2217_), .Y(new_n12764_));
  XOR2   g11762(.A(new_n2165_), .B(new_n12764_), .Y(new_n12765_));
  NAND2  g11763(.A(new_n2174_), .B(new_n2161_), .Y(new_n12766_));
  OAI21  g11764(.A0(new_n2165_), .A1(new_n2157_), .B0(new_n12766_), .Y(new_n12767_));
  OAI21  g11765(.A0(new_n2171_), .A1(new_n12765_), .B0(new_n12767_), .Y(new_n12768_));
  NOR2   g11766(.A(new_n12768_), .B(new_n12763_), .Y(new_n12769_));
  OAI21  g11767(.A0(new_n2231_), .A1(new_n2222_), .B0(new_n2204_), .Y(new_n12770_));
  AOI21  g11768(.A0(new_n2218_), .A1(new_n2166_), .B0(new_n2176_), .Y(new_n12771_));
  NOR2   g11769(.A(new_n12771_), .B(new_n12770_), .Y(new_n12772_));
  OAI21  g11770(.A0(new_n12772_), .A1(new_n12769_), .B0(new_n12762_), .Y(new_n12773_));
  OAI211 g11771(.A0(new_n2171_), .A1(new_n12765_), .B0(new_n12770_), .B1(new_n12767_), .Y(new_n12774_));
  NAND2  g11772(.A(new_n12768_), .B(new_n12763_), .Y(new_n12775_));
  NAND4  g11773(.A(new_n12775_), .B(new_n12774_), .C(new_n12761_), .D(new_n12760_), .Y(new_n12776_));
  NAND2  g11774(.A(new_n12776_), .B(new_n12773_), .Y(new_n12777_));
  NOR3   g11775(.A(new_n2295_), .B(new_n2293_), .C(new_n2314_), .Y(new_n12778_));
  OAI211 g11776(.A0(new_n2327_), .A1(new_n2344_), .B0(new_n12778_), .B1(new_n2338_), .Y(new_n12779_));
  OAI21  g11777(.A0(new_n2315_), .A1(new_n2296_), .B0(new_n2322_), .Y(new_n12780_));
  OAI21  g11778(.A0(new_n2327_), .A1(new_n2314_), .B0(new_n2312_), .Y(new_n12781_));
  OAI211 g11779(.A0(new_n2268_), .A1(new_n2319_), .B0(new_n12781_), .B1(new_n2321_), .Y(new_n12782_));
  AOI21  g11780(.A0(new_n2294_), .A1(new_n2345_), .B0(new_n2344_), .Y(new_n12783_));
  OAI21  g11781(.A0(new_n2268_), .A1(new_n2319_), .B0(new_n2321_), .Y(new_n12784_));
  NAND2  g11782(.A(new_n12784_), .B(new_n12783_), .Y(new_n12785_));
  AOI22  g11783(.A0(new_n12785_), .A1(new_n12782_), .B0(new_n12780_), .B1(new_n12779_), .Y(new_n12786_));
  AOI221 g11784(.A0(new_n2346_), .A1(new_n2339_), .C0(new_n2319_), .B0(new_n2321_), .B1(new_n2267_), .Y(new_n12787_));
  NOR2   g11785(.A(new_n12784_), .B(new_n12783_), .Y(new_n12788_));
  NAND2  g11786(.A(new_n2267_), .B(new_n2258_), .Y(new_n12789_));
  AOI21  g11787(.A0(new_n12789_), .A1(new_n2321_), .B0(new_n12781_), .Y(new_n12790_));
  NOR4   g11788(.A(new_n12790_), .B(new_n12788_), .C(new_n12787_), .D(new_n2325_), .Y(new_n12791_));
  NOR2   g11789(.A(new_n12791_), .B(new_n12786_), .Y(new_n12792_));
  XOR2   g11790(.A(new_n12792_), .B(new_n12777_), .Y(new_n12793_));
  XOR2   g11791(.A(new_n12793_), .B(new_n12758_), .Y(new_n12794_));
  XOR2   g11792(.A(new_n12794_), .B(new_n12756_), .Y(new_n12795_));
  XOR2   g11793(.A(new_n12795_), .B(new_n12716_), .Y(new_n12796_));
  AOI21  g11794(.A0(new_n2822_), .A1(new_n2818_), .B0(new_n2824_), .Y(new_n12797_));
  NOR2   g11795(.A(new_n12797_), .B(new_n2825_), .Y(new_n12798_));
  OAI22  g11796(.A0(new_n2819_), .A1(new_n2450_), .B0(new_n2584_), .B1(new_n2579_), .Y(new_n12799_));
  NAND2  g11797(.A(new_n12799_), .B(new_n2587_), .Y(new_n12800_));
  NAND4  g11798(.A(new_n2526_), .B(new_n2550_), .C(new_n2567_), .D(new_n2537_), .Y(new_n12801_));
  AOI221 g11799(.A0(new_n2582_), .A1(new_n2530_), .C0(new_n12801_), .B0(new_n2558_), .B1(new_n2537_), .Y(new_n12802_));
  AOI21  g11800(.A0(new_n2568_), .A1(new_n2554_), .B0(new_n2583_), .Y(new_n12803_));
  AOI21  g11801(.A0(new_n2567_), .A1(new_n2537_), .B0(new_n2566_), .Y(new_n12804_));
  AOI211 g11802(.A0(new_n2582_), .A1(new_n2526_), .B(new_n12804_), .C(new_n2581_), .Y(new_n12805_));
  OAI21  g11803(.A0(new_n2560_), .A1(new_n2563_), .B0(new_n2558_), .Y(new_n12806_));
  AOI21  g11804(.A0(new_n2582_), .A1(new_n2526_), .B0(new_n2581_), .Y(new_n12807_));
  NOR2   g11805(.A(new_n12807_), .B(new_n12806_), .Y(new_n12808_));
  OAI22  g11806(.A0(new_n12808_), .A1(new_n12805_), .B0(new_n12803_), .B1(new_n12802_), .Y(new_n12809_));
  NAND2  g11807(.A(new_n2569_), .B(new_n2536_), .Y(new_n12810_));
  NAND2  g11808(.A(new_n12807_), .B(new_n12806_), .Y(new_n12811_));
  OAI21  g11809(.A0(new_n2535_), .A1(new_n2572_), .B0(new_n2530_), .Y(new_n12812_));
  NAND2  g11810(.A(new_n12812_), .B(new_n12804_), .Y(new_n12813_));
  NAND4  g11811(.A(new_n12813_), .B(new_n12811_), .C(new_n12810_), .D(new_n2574_), .Y(new_n12814_));
  NAND2  g11812(.A(new_n12814_), .B(new_n12809_), .Y(new_n12815_));
  NOR3   g11813(.A(new_n2465_), .B(new_n2464_), .C(new_n2447_), .Y(new_n12816_));
  OAI211 g11814(.A0(new_n2462_), .A1(new_n2460_), .B0(new_n12816_), .B1(new_n2430_), .Y(new_n12817_));
  OAI21  g11815(.A0(new_n2448_), .A1(new_n2515_), .B0(new_n2409_), .Y(new_n12818_));
  OAI21  g11816(.A0(new_n2462_), .A1(new_n2447_), .B0(new_n2445_), .Y(new_n12819_));
  OAI211 g11817(.A0(new_n2452_), .A1(new_n2394_), .B0(new_n12819_), .B1(new_n2408_), .Y(new_n12820_));
  AOI21  g11818(.A0(new_n2438_), .A1(new_n2461_), .B0(new_n2460_), .Y(new_n12821_));
  OAI21  g11819(.A0(new_n2452_), .A1(new_n2394_), .B0(new_n2408_), .Y(new_n12822_));
  NAND2  g11820(.A(new_n12822_), .B(new_n12821_), .Y(new_n12823_));
  AOI22  g11821(.A0(new_n12823_), .A1(new_n12820_), .B0(new_n12818_), .B1(new_n12817_), .Y(new_n12824_));
  AOI221 g11822(.A0(new_n2463_), .A1(new_n2439_), .C0(new_n2394_), .B0(new_n2408_), .B1(new_n2395_), .Y(new_n12825_));
  NOR2   g11823(.A(new_n12822_), .B(new_n12821_), .Y(new_n12826_));
  AOI21  g11824(.A0(new_n2395_), .A1(new_n2451_), .B0(new_n2454_), .Y(new_n12827_));
  NOR2   g11825(.A(new_n12827_), .B(new_n12819_), .Y(new_n12828_));
  NOR4   g11826(.A(new_n12828_), .B(new_n12826_), .C(new_n12825_), .D(new_n2467_), .Y(new_n12829_));
  NOR2   g11827(.A(new_n12829_), .B(new_n12824_), .Y(new_n12830_));
  XOR2   g11828(.A(new_n12830_), .B(new_n12815_), .Y(new_n12831_));
  XOR2   g11829(.A(new_n12831_), .B(new_n12800_), .Y(new_n12832_));
  OAI21  g11830(.A0(new_n2788_), .A1(new_n2714_), .B0(new_n2793_), .Y(new_n12833_));
  OAI22  g11831(.A0(new_n12833_), .A1(new_n2782_), .B0(new_n2802_), .B1(new_n2796_), .Y(new_n12834_));
  NAND2  g11832(.A(new_n12834_), .B(new_n2805_), .Y(new_n12835_));
  AOI221 g11833(.A0(new_n2800_), .A1(new_n2657_), .C0(new_n2611_), .B0(new_n2625_), .B1(new_n2612_), .Y(new_n12836_));
  AOI21  g11834(.A0(new_n2656_), .A1(new_n2669_), .B0(new_n2798_), .Y(new_n12837_));
  XOR2   g11835(.A(new_n2603_), .B(new_n2616_), .Y(new_n12838_));
  OAI21  g11836(.A0(new_n12838_), .A1(new_n2611_), .B0(new_n2625_), .Y(new_n12839_));
  NOR2   g11837(.A(new_n12839_), .B(new_n12837_), .Y(new_n12840_));
  OAI21  g11838(.A0(new_n2799_), .A1(new_n2665_), .B0(new_n2663_), .Y(new_n12841_));
  XOR2   g11839(.A(new_n2610_), .B(new_n2621_), .Y(new_n12842_));
  XOR2   g11840(.A(new_n2623_), .B(new_n2607_), .Y(new_n12843_));
  NAND2  g11841(.A(new_n12843_), .B(new_n2604_), .Y(new_n12844_));
  AOI22  g11842(.A0(new_n2624_), .A1(new_n12844_), .B0(new_n2612_), .B1(new_n12842_), .Y(new_n12845_));
  NOR2   g11843(.A(new_n12845_), .B(new_n12841_), .Y(new_n12846_));
  OAI22  g11844(.A0(new_n12846_), .A1(new_n12840_), .B0(new_n12836_), .B1(new_n2675_), .Y(new_n12847_));
  NOR3   g11845(.A(new_n2671_), .B(new_n2670_), .C(new_n2665_), .Y(new_n12848_));
  OAI211 g11846(.A0(new_n2799_), .A1(new_n2798_), .B0(new_n12848_), .B1(new_n2648_), .Y(new_n12849_));
  OAI21  g11847(.A0(new_n2666_), .A1(new_n2672_), .B0(new_n2626_), .Y(new_n12850_));
  NAND2  g11848(.A(new_n12845_), .B(new_n12841_), .Y(new_n12851_));
  NAND2  g11849(.A(new_n12839_), .B(new_n12837_), .Y(new_n12852_));
  NAND4  g11850(.A(new_n12852_), .B(new_n12851_), .C(new_n12850_), .D(new_n12849_), .Y(new_n12853_));
  NAND2  g11851(.A(new_n12853_), .B(new_n12847_), .Y(new_n12854_));
  AOI221 g11852(.A0(new_n2787_), .A1(new_n2780_), .C0(new_n2760_), .B0(new_n2762_), .B1(new_n2708_), .Y(new_n12855_));
  AOI21  g11853(.A0(new_n2735_), .A1(new_n2786_), .B0(new_n2785_), .Y(new_n12856_));
  OAI21  g11854(.A0(new_n2709_), .A1(new_n2760_), .B0(new_n2762_), .Y(new_n12857_));
  NOR2   g11855(.A(new_n12857_), .B(new_n12856_), .Y(new_n12858_));
  OAI21  g11856(.A0(new_n2768_), .A1(new_n2755_), .B0(new_n2753_), .Y(new_n12859_));
  NAND2  g11857(.A(new_n2708_), .B(new_n2699_), .Y(new_n12860_));
  AOI21  g11858(.A0(new_n12860_), .A1(new_n2762_), .B0(new_n12859_), .Y(new_n12861_));
  OAI22  g11859(.A0(new_n12861_), .A1(new_n12858_), .B0(new_n12855_), .B1(new_n2766_), .Y(new_n12862_));
  NOR3   g11860(.A(new_n2736_), .B(new_n2734_), .C(new_n2755_), .Y(new_n12863_));
  OAI211 g11861(.A0(new_n2768_), .A1(new_n2785_), .B0(new_n12863_), .B1(new_n2779_), .Y(new_n12864_));
  OAI21  g11862(.A0(new_n2756_), .A1(new_n2737_), .B0(new_n2763_), .Y(new_n12865_));
  OAI211 g11863(.A0(new_n2709_), .A1(new_n2760_), .B0(new_n12859_), .B1(new_n2762_), .Y(new_n12866_));
  NAND2  g11864(.A(new_n12857_), .B(new_n12856_), .Y(new_n12867_));
  NAND4  g11865(.A(new_n12867_), .B(new_n12866_), .C(new_n12865_), .D(new_n12864_), .Y(new_n12868_));
  NAND2  g11866(.A(new_n12868_), .B(new_n12862_), .Y(new_n12869_));
  XOR2   g11867(.A(new_n12869_), .B(new_n12854_), .Y(new_n12870_));
  XOR2   g11868(.A(new_n12870_), .B(new_n12835_), .Y(new_n12871_));
  XOR2   g11869(.A(new_n12871_), .B(new_n12832_), .Y(new_n12872_));
  XOR2   g11870(.A(new_n12872_), .B(new_n12798_), .Y(new_n12873_));
  XOR2   g11871(.A(new_n12873_), .B(new_n12796_), .Y(new_n12874_));
  XOR2   g11872(.A(new_n12874_), .B(new_n12715_), .Y(new_n12875_));
  XOR2   g11873(.A(new_n12875_), .B(new_n12714_), .Y(new_n12876_));
  XOR2   g11874(.A(new_n12876_), .B(new_n12554_), .Y(new_n12877_));
  XOR2   g11875(.A(new_n12877_), .B(new_n12553_), .Y(new_n12878_));
  XOR2   g11876(.A(new_n12878_), .B(new_n12240_), .Y(new_n12879_));
  NAND2  g11877(.A(new_n12879_), .B(new_n12231_), .Y(new_n12880_));
  AOI21  g11878(.A0(new_n11193_), .A1(new_n11178_), .B0(new_n11180_), .Y(new_n12881_));
  XOR2   g11879(.A(new_n12228_), .B(new_n12881_), .Y(new_n12882_));
  XOR2   g11880(.A(new_n12882_), .B(new_n11608_), .Y(new_n12883_));
  NOR2   g11881(.A(new_n12883_), .B(new_n11219_), .Y(new_n12884_));
  AOI21  g11882(.A0(new_n11181_), .A1(new_n11171_), .B0(new_n11196_), .Y(new_n12885_));
  AOI21  g11883(.A0(new_n11206_), .A1(new_n7058_), .B0(new_n12885_), .Y(new_n12886_));
  NOR3   g11884(.A(new_n3547_), .B(new_n3554_), .C(new_n3551_), .Y(new_n12887_));
  OAI21  g11885(.A0(new_n12887_), .A1(new_n4767_), .B0(new_n4769_), .Y(new_n12888_));
  XOR2   g11886(.A(new_n12878_), .B(new_n12888_), .Y(new_n12889_));
  OAI21  g11887(.A0(new_n12230_), .A1(new_n12886_), .B0(new_n12889_), .Y(new_n12890_));
  NOR2   g11888(.A(new_n12890_), .B(new_n12884_), .Y(new_n12891_));
  AOI21  g11889(.A0(new_n12880_), .A1(new_n11217_), .B0(new_n12891_), .Y(new_n12892_));
  NOR2   g11890(.A(new_n12882_), .B(new_n11608_), .Y(new_n12893_));
  NAND2  g11891(.A(new_n12882_), .B(new_n11608_), .Y(new_n12894_));
  OAI21  g11892(.A0(new_n12893_), .A1(new_n12886_), .B0(new_n12894_), .Y(new_n12895_));
  AOI21  g11893(.A0(new_n11154_), .A1(new_n10122_), .B0(new_n11168_), .Y(new_n12896_));
  XOR2   g11894(.A(new_n12226_), .B(new_n12896_), .Y(new_n12897_));
  NAND2  g11895(.A(new_n12897_), .B(new_n11918_), .Y(new_n12898_));
  NOR2   g11896(.A(new_n12897_), .B(new_n11918_), .Y(new_n12899_));
  AOI21  g11897(.A0(new_n12898_), .A1(new_n11609_), .B0(new_n12899_), .Y(new_n12900_));
  NOR2   g11898(.A(new_n12225_), .B(new_n12075_), .Y(new_n12901_));
  NAND2  g11899(.A(new_n12225_), .B(new_n12075_), .Y(new_n12902_));
  OAI21  g11900(.A0(new_n12901_), .A1(new_n12896_), .B0(new_n12902_), .Y(new_n12903_));
  AOI21  g11901(.A0(new_n11141_), .A1(new_n11130_), .B0(new_n11132_), .Y(new_n12904_));
  NOR2   g11902(.A(new_n12223_), .B(new_n12150_), .Y(new_n12905_));
  NAND2  g11903(.A(new_n12223_), .B(new_n12150_), .Y(new_n12906_));
  OAI21  g11904(.A0(new_n12905_), .A1(new_n12904_), .B0(new_n12906_), .Y(new_n12907_));
  OAI22  g11905(.A0(new_n12183_), .A1(new_n12182_), .B0(new_n12181_), .B1(new_n10846_), .Y(new_n12908_));
  NAND2  g11906(.A(new_n10711_), .B(new_n10647_), .Y(new_n12909_));
  NAND4  g11907(.A(new_n12179_), .B(new_n12176_), .C(new_n12909_), .D(new_n10714_), .Y(new_n12910_));
  NAND2  g11908(.A(new_n12910_), .B(new_n12908_), .Y(new_n12911_));
  XOR2   g11909(.A(new_n12911_), .B(new_n12171_), .Y(new_n12912_));
  XOR2   g11910(.A(new_n12912_), .B(new_n12154_), .Y(new_n12913_));
  OAI22  g11911(.A0(new_n12221_), .A1(new_n12913_), .B0(new_n12151_), .B1(new_n11120_), .Y(new_n12914_));
  NAND2  g11912(.A(new_n12221_), .B(new_n12913_), .Y(new_n12915_));
  NAND2  g11913(.A(new_n12915_), .B(new_n12914_), .Y(new_n12916_));
  NOR2   g11914(.A(new_n11077_), .B(new_n11075_), .Y(new_n12917_));
  OAI22  g11915(.A0(new_n11085_), .A1(new_n11041_), .B0(new_n10946_), .B1(new_n12917_), .Y(new_n12918_));
  AOI22  g11916(.A0(new_n12219_), .A1(new_n12205_), .B0(new_n12918_), .B1(new_n11086_), .Y(new_n12919_));
  AOI22  g11917(.A0(new_n12203_), .A1(new_n12202_), .B0(new_n12201_), .B1(new_n10945_), .Y(new_n12920_));
  NOR4   g11918(.A(new_n12199_), .B(new_n12196_), .C(new_n12193_), .D(new_n12192_), .Y(new_n12921_));
  AOI21  g11919(.A0(new_n11047_), .A1(new_n10983_), .B0(new_n11083_), .Y(new_n12922_));
  AOI21  g11920(.A0(new_n12217_), .A1(new_n12216_), .B0(new_n12922_), .Y(new_n12923_));
  NOR4   g11921(.A(new_n12213_), .B(new_n12209_), .C(new_n12206_), .D(new_n11083_), .Y(new_n12924_));
  NOR4   g11922(.A(new_n12924_), .B(new_n12923_), .C(new_n12921_), .D(new_n12920_), .Y(new_n12925_));
  AOI211 g11923(.A0(new_n11047_), .A1(new_n10983_), .B(new_n12207_), .C(new_n11083_), .Y(new_n12926_));
  OAI22  g11924(.A0(new_n12926_), .A1(new_n12208_), .B0(new_n12211_), .B1(new_n12922_), .Y(new_n12927_));
  NOR3   g11925(.A(new_n12194_), .B(new_n12193_), .C(new_n12192_), .Y(new_n12928_));
  OAI21  g11926(.A0(new_n12193_), .A1(new_n12192_), .B0(new_n12194_), .Y(new_n12929_));
  OAI21  g11927(.A0(new_n12928_), .A1(new_n12195_), .B0(new_n12929_), .Y(new_n12930_));
  XOR2   g11928(.A(new_n12930_), .B(new_n12927_), .Y(new_n12931_));
  OAI21  g11929(.A0(new_n12925_), .A1(new_n12919_), .B0(new_n12931_), .Y(new_n12932_));
  OAI22  g11930(.A0(new_n12924_), .A1(new_n12923_), .B0(new_n12921_), .B1(new_n12920_), .Y(new_n12933_));
  NAND2  g11931(.A(new_n12933_), .B(new_n12189_), .Y(new_n12934_));
  NAND3  g11932(.A(new_n12197_), .B(new_n12201_), .C(new_n10945_), .Y(new_n12935_));
  AOI21  g11933(.A0(new_n12201_), .A1(new_n10945_), .B0(new_n12197_), .Y(new_n12936_));
  AOI21  g11934(.A0(new_n12935_), .A1(new_n12198_), .B0(new_n12936_), .Y(new_n12937_));
  AOI21  g11935(.A0(new_n12937_), .A1(new_n12927_), .B0(new_n12925_), .Y(new_n12938_));
  OAI211 g11936(.A0(new_n12937_), .A1(new_n12927_), .B0(new_n12938_), .B1(new_n12934_), .Y(new_n12939_));
  NAND2  g11937(.A(new_n12939_), .B(new_n12932_), .Y(new_n12940_));
  AOI21  g11938(.A0(new_n12166_), .A1(new_n10828_), .B0(new_n10838_), .Y(new_n12941_));
  OAI22  g11939(.A0(new_n10848_), .A1(new_n10705_), .B0(new_n12941_), .B1(new_n10827_), .Y(new_n12942_));
  AOI22  g11940(.A0(new_n12911_), .A1(new_n12171_), .B0(new_n12942_), .B1(new_n10849_), .Y(new_n12943_));
  AOI22  g11941(.A0(new_n12169_), .A1(new_n12168_), .B0(new_n12167_), .B1(new_n12166_), .Y(new_n12944_));
  NOR4   g11942(.A(new_n12163_), .B(new_n12159_), .C(new_n12156_), .D(new_n12155_), .Y(new_n12945_));
  NOR4   g11943(.A(new_n12184_), .B(new_n12180_), .C(new_n12945_), .D(new_n12944_), .Y(new_n12946_));
  AOI211 g11944(.A0(new_n10711_), .A1(new_n10647_), .B(new_n12177_), .C(new_n10846_), .Y(new_n12947_));
  OAI22  g11945(.A0(new_n12947_), .A1(new_n12178_), .B0(new_n12174_), .B1(new_n12172_), .Y(new_n12948_));
  NOR3   g11946(.A(new_n12157_), .B(new_n12156_), .C(new_n12155_), .Y(new_n12949_));
  OAI21  g11947(.A0(new_n12156_), .A1(new_n12155_), .B0(new_n12157_), .Y(new_n12950_));
  OAI21  g11948(.A0(new_n12949_), .A1(new_n12158_), .B0(new_n12950_), .Y(new_n12951_));
  XOR2   g11949(.A(new_n12951_), .B(new_n12948_), .Y(new_n12952_));
  OAI21  g11950(.A0(new_n12946_), .A1(new_n12943_), .B0(new_n12952_), .Y(new_n12953_));
  OAI22  g11951(.A0(new_n12184_), .A1(new_n12180_), .B0(new_n12945_), .B1(new_n12944_), .Y(new_n12954_));
  NAND2  g11952(.A(new_n12954_), .B(new_n12154_), .Y(new_n12955_));
  NAND4  g11953(.A(new_n12910_), .B(new_n12908_), .C(new_n12170_), .D(new_n12164_), .Y(new_n12956_));
  OAI211 g11954(.A0(new_n12949_), .A1(new_n12158_), .B0(new_n12950_), .B1(new_n12948_), .Y(new_n12957_));
  NOR2   g11955(.A(new_n12947_), .B(new_n12178_), .Y(new_n12958_));
  NOR2   g11956(.A(new_n12174_), .B(new_n12172_), .Y(new_n12959_));
  NOR2   g11957(.A(new_n12959_), .B(new_n12958_), .Y(new_n12960_));
  NAND2  g11958(.A(new_n12951_), .B(new_n12960_), .Y(new_n12961_));
  NAND4  g11959(.A(new_n12961_), .B(new_n12957_), .C(new_n12956_), .D(new_n12955_), .Y(new_n12962_));
  NAND2  g11960(.A(new_n12962_), .B(new_n12953_), .Y(new_n12963_));
  XOR2   g11961(.A(new_n12963_), .B(new_n12940_), .Y(new_n12964_));
  XOR2   g11962(.A(new_n12964_), .B(new_n12916_), .Y(new_n12965_));
  NAND2  g11963(.A(new_n12148_), .B(new_n12115_), .Y(new_n12966_));
  NOR2   g11964(.A(new_n12148_), .B(new_n12115_), .Y(new_n12967_));
  AOI21  g11965(.A0(new_n12966_), .A1(new_n12077_), .B0(new_n12967_), .Y(new_n12968_));
  AOI22  g11966(.A0(new_n12130_), .A1(new_n12129_), .B0(new_n12128_), .B1(new_n10215_), .Y(new_n12969_));
  NOR4   g11967(.A(new_n12126_), .B(new_n12123_), .C(new_n12118_), .D(new_n10345_), .Y(new_n12970_));
  OAI22  g11968(.A0(new_n12145_), .A1(new_n12141_), .B0(new_n12970_), .B1(new_n12969_), .Y(new_n12971_));
  NOR4   g11969(.A(new_n12145_), .B(new_n12141_), .C(new_n12970_), .D(new_n12969_), .Y(new_n12972_));
  AOI21  g11970(.A0(new_n12971_), .A1(new_n12117_), .B0(new_n12972_), .Y(new_n12973_));
  AOI211 g11971(.A0(new_n10317_), .A1(new_n10253_), .B(new_n12138_), .C(new_n10350_), .Y(new_n12974_));
  OAI22  g11972(.A0(new_n12974_), .A1(new_n12139_), .B0(new_n12135_), .B1(new_n12133_), .Y(new_n12975_));
  NAND3  g11973(.A(new_n12124_), .B(new_n12128_), .C(new_n10215_), .Y(new_n12976_));
  AOI21  g11974(.A0(new_n12128_), .A1(new_n10215_), .B0(new_n12124_), .Y(new_n12977_));
  AOI21  g11975(.A0(new_n12976_), .A1(new_n12125_), .B0(new_n12977_), .Y(new_n12978_));
  XOR2   g11976(.A(new_n12978_), .B(new_n12975_), .Y(new_n12979_));
  NAND2  g11977(.A(new_n12971_), .B(new_n12117_), .Y(new_n12980_));
  AOI21  g11978(.A0(new_n12978_), .A1(new_n12975_), .B0(new_n12972_), .Y(new_n12981_));
  OAI211 g11979(.A0(new_n12978_), .A1(new_n12975_), .B0(new_n12981_), .B1(new_n12980_), .Y(new_n12982_));
  OAI21  g11980(.A0(new_n12979_), .A1(new_n12973_), .B0(new_n12982_), .Y(new_n12983_));
  AOI22  g11981(.A0(new_n12097_), .A1(new_n12096_), .B0(new_n12095_), .B1(new_n12094_), .Y(new_n12984_));
  NOR4   g11982(.A(new_n12091_), .B(new_n12084_), .C(new_n12081_), .D(new_n12079_), .Y(new_n12985_));
  OAI22  g11983(.A0(new_n12112_), .A1(new_n12107_), .B0(new_n12985_), .B1(new_n12984_), .Y(new_n12986_));
  NOR4   g11984(.A(new_n12112_), .B(new_n12107_), .C(new_n12985_), .D(new_n12984_), .Y(new_n12987_));
  AOI21  g11985(.A0(new_n12986_), .A1(new_n12078_), .B0(new_n12987_), .Y(new_n12988_));
  NOR3   g11986(.A(new_n12104_), .B(new_n12109_), .C(new_n12108_), .Y(new_n12989_));
  OAI21  g11987(.A0(new_n12109_), .A1(new_n12108_), .B0(new_n12104_), .Y(new_n12990_));
  OAI21  g11988(.A0(new_n12989_), .A1(new_n12105_), .B0(new_n12990_), .Y(new_n12991_));
  NAND3  g11989(.A(new_n12086_), .B(new_n12095_), .C(new_n12094_), .Y(new_n12992_));
  AOI21  g11990(.A0(new_n12095_), .A1(new_n12094_), .B0(new_n12086_), .Y(new_n12993_));
  AOI21  g11991(.A0(new_n12992_), .A1(new_n12090_), .B0(new_n12993_), .Y(new_n12994_));
  XOR2   g11992(.A(new_n12994_), .B(new_n12991_), .Y(new_n12995_));
  NOR2   g11993(.A(new_n12995_), .B(new_n12988_), .Y(new_n12996_));
  NAND3  g11994(.A(new_n12101_), .B(new_n12100_), .C(new_n10600_), .Y(new_n12997_));
  AOI21  g11995(.A0(new_n12100_), .A1(new_n10600_), .B0(new_n12101_), .Y(new_n12998_));
  AOI21  g11996(.A0(new_n12997_), .A1(new_n12102_), .B0(new_n12998_), .Y(new_n12999_));
  NOR3   g11997(.A(new_n12082_), .B(new_n12081_), .C(new_n12079_), .Y(new_n13000_));
  OAI21  g11998(.A0(new_n12081_), .A1(new_n12079_), .B0(new_n12082_), .Y(new_n13001_));
  OAI21  g11999(.A0(new_n13000_), .A1(new_n12083_), .B0(new_n13001_), .Y(new_n13002_));
  NAND4  g12000(.A(new_n12106_), .B(new_n12103_), .C(new_n12100_), .D(new_n10600_), .Y(new_n13003_));
  NAND3  g12001(.A(new_n13003_), .B(new_n12098_), .C(new_n12092_), .Y(new_n13004_));
  OAI22  g12002(.A0(new_n13002_), .A1(new_n12999_), .B0(new_n13004_), .B1(new_n12107_), .Y(new_n13005_));
  AOI221 g12003(.A0(new_n13002_), .A1(new_n12999_), .C0(new_n13005_), .B0(new_n12986_), .B1(new_n12078_), .Y(new_n13006_));
  NOR2   g12004(.A(new_n13006_), .B(new_n12996_), .Y(new_n13007_));
  XOR2   g12005(.A(new_n13007_), .B(new_n12983_), .Y(new_n13008_));
  XOR2   g12006(.A(new_n13008_), .B(new_n12968_), .Y(new_n13009_));
  XOR2   g12007(.A(new_n13009_), .B(new_n12965_), .Y(new_n13010_));
  XOR2   g12008(.A(new_n13010_), .B(new_n12907_), .Y(new_n13011_));
  AOI22  g12009(.A0(new_n10106_), .A1(new_n9914_), .B0(new_n10084_), .B1(new_n10078_), .Y(new_n13012_));
  NOR2   g12010(.A(new_n13012_), .B(new_n10116_), .Y(new_n13013_));
  XOR2   g12011(.A(new_n11999_), .B(new_n13013_), .Y(new_n13014_));
  OAI21  g12012(.A0(new_n9777_), .A1(new_n9602_), .B0(new_n9605_), .Y(new_n13015_));
  XOR2   g12013(.A(new_n12072_), .B(new_n13015_), .Y(new_n13016_));
  NAND2  g12014(.A(new_n13016_), .B(new_n13014_), .Y(new_n13017_));
  NOR2   g12015(.A(new_n13016_), .B(new_n13014_), .Y(new_n13018_));
  AOI21  g12016(.A0(new_n13017_), .A1(new_n11920_), .B0(new_n13018_), .Y(new_n13019_));
  OAI22  g12017(.A0(new_n12033_), .A1(new_n12032_), .B0(new_n12031_), .B1(new_n9344_), .Y(new_n13020_));
  NAND2  g12018(.A(new_n9209_), .B(new_n9145_), .Y(new_n13021_));
  NAND4  g12019(.A(new_n12029_), .B(new_n12026_), .C(new_n13021_), .D(new_n9212_), .Y(new_n13022_));
  NAND2  g12020(.A(new_n13022_), .B(new_n13020_), .Y(new_n13023_));
  XOR2   g12021(.A(new_n13023_), .B(new_n12021_), .Y(new_n13024_));
  XOR2   g12022(.A(new_n13024_), .B(new_n12004_), .Y(new_n13025_));
  OAI22  g12023(.A0(new_n12071_), .A1(new_n13025_), .B0(new_n12001_), .B1(new_n9778_), .Y(new_n13026_));
  NAND2  g12024(.A(new_n12071_), .B(new_n13025_), .Y(new_n13027_));
  NAND2  g12025(.A(new_n13027_), .B(new_n13026_), .Y(new_n13028_));
  NOR2   g12026(.A(new_n9575_), .B(new_n9573_), .Y(new_n13029_));
  OAI22  g12027(.A0(new_n9583_), .A1(new_n9539_), .B0(new_n9444_), .B1(new_n13029_), .Y(new_n13030_));
  AOI22  g12028(.A0(new_n12069_), .A1(new_n12055_), .B0(new_n13030_), .B1(new_n9584_), .Y(new_n13031_));
  AOI22  g12029(.A0(new_n12053_), .A1(new_n12052_), .B0(new_n12051_), .B1(new_n9443_), .Y(new_n13032_));
  NOR4   g12030(.A(new_n12049_), .B(new_n12046_), .C(new_n12043_), .D(new_n12042_), .Y(new_n13033_));
  AOI21  g12031(.A0(new_n9545_), .A1(new_n9481_), .B0(new_n9581_), .Y(new_n13034_));
  AOI21  g12032(.A0(new_n12067_), .A1(new_n12066_), .B0(new_n13034_), .Y(new_n13035_));
  NOR4   g12033(.A(new_n12063_), .B(new_n12059_), .C(new_n12056_), .D(new_n9581_), .Y(new_n13036_));
  NOR4   g12034(.A(new_n13036_), .B(new_n13035_), .C(new_n13033_), .D(new_n13032_), .Y(new_n13037_));
  AOI211 g12035(.A0(new_n9545_), .A1(new_n9481_), .B(new_n12057_), .C(new_n9581_), .Y(new_n13038_));
  OAI22  g12036(.A0(new_n13038_), .A1(new_n12058_), .B0(new_n12061_), .B1(new_n13034_), .Y(new_n13039_));
  NOR3   g12037(.A(new_n12044_), .B(new_n12043_), .C(new_n12042_), .Y(new_n13040_));
  OAI21  g12038(.A0(new_n12043_), .A1(new_n12042_), .B0(new_n12044_), .Y(new_n13041_));
  OAI21  g12039(.A0(new_n13040_), .A1(new_n12045_), .B0(new_n13041_), .Y(new_n13042_));
  XOR2   g12040(.A(new_n13042_), .B(new_n13039_), .Y(new_n13043_));
  OAI21  g12041(.A0(new_n13037_), .A1(new_n13031_), .B0(new_n13043_), .Y(new_n13044_));
  OAI22  g12042(.A0(new_n13036_), .A1(new_n13035_), .B0(new_n13033_), .B1(new_n13032_), .Y(new_n13045_));
  NAND2  g12043(.A(new_n13045_), .B(new_n12039_), .Y(new_n13046_));
  NAND3  g12044(.A(new_n12047_), .B(new_n12051_), .C(new_n9443_), .Y(new_n13047_));
  AOI21  g12045(.A0(new_n12051_), .A1(new_n9443_), .B0(new_n12047_), .Y(new_n13048_));
  AOI21  g12046(.A0(new_n13047_), .A1(new_n12048_), .B0(new_n13048_), .Y(new_n13049_));
  AOI21  g12047(.A0(new_n13049_), .A1(new_n13039_), .B0(new_n13037_), .Y(new_n13050_));
  OAI211 g12048(.A0(new_n13049_), .A1(new_n13039_), .B0(new_n13050_), .B1(new_n13046_), .Y(new_n13051_));
  NAND2  g12049(.A(new_n13051_), .B(new_n13044_), .Y(new_n13052_));
  AOI21  g12050(.A0(new_n12016_), .A1(new_n9326_), .B0(new_n9336_), .Y(new_n13053_));
  OAI22  g12051(.A0(new_n9346_), .A1(new_n9203_), .B0(new_n13053_), .B1(new_n9325_), .Y(new_n13054_));
  AOI22  g12052(.A0(new_n13023_), .A1(new_n12021_), .B0(new_n13054_), .B1(new_n9347_), .Y(new_n13055_));
  AOI22  g12053(.A0(new_n12019_), .A1(new_n12018_), .B0(new_n12017_), .B1(new_n12016_), .Y(new_n13056_));
  NOR4   g12054(.A(new_n12013_), .B(new_n12009_), .C(new_n12006_), .D(new_n12005_), .Y(new_n13057_));
  NOR4   g12055(.A(new_n12034_), .B(new_n12030_), .C(new_n13057_), .D(new_n13056_), .Y(new_n13058_));
  AOI211 g12056(.A0(new_n9209_), .A1(new_n9145_), .B(new_n12027_), .C(new_n9344_), .Y(new_n13059_));
  OAI22  g12057(.A0(new_n13059_), .A1(new_n12028_), .B0(new_n12024_), .B1(new_n12022_), .Y(new_n13060_));
  NOR3   g12058(.A(new_n12007_), .B(new_n12006_), .C(new_n12005_), .Y(new_n13061_));
  OAI21  g12059(.A0(new_n12006_), .A1(new_n12005_), .B0(new_n12007_), .Y(new_n13062_));
  OAI21  g12060(.A0(new_n13061_), .A1(new_n12008_), .B0(new_n13062_), .Y(new_n13063_));
  XOR2   g12061(.A(new_n13063_), .B(new_n13060_), .Y(new_n13064_));
  OAI21  g12062(.A0(new_n13058_), .A1(new_n13055_), .B0(new_n13064_), .Y(new_n13065_));
  OAI22  g12063(.A0(new_n12034_), .A1(new_n12030_), .B0(new_n13057_), .B1(new_n13056_), .Y(new_n13066_));
  NAND2  g12064(.A(new_n13066_), .B(new_n12004_), .Y(new_n13067_));
  NAND4  g12065(.A(new_n13022_), .B(new_n13020_), .C(new_n12020_), .D(new_n12014_), .Y(new_n13068_));
  OAI211 g12066(.A0(new_n13061_), .A1(new_n12008_), .B0(new_n13062_), .B1(new_n13060_), .Y(new_n13069_));
  NOR2   g12067(.A(new_n13059_), .B(new_n12028_), .Y(new_n13070_));
  NOR2   g12068(.A(new_n12024_), .B(new_n12022_), .Y(new_n13071_));
  NOR2   g12069(.A(new_n13071_), .B(new_n13070_), .Y(new_n13072_));
  NAND2  g12070(.A(new_n13063_), .B(new_n13072_), .Y(new_n13073_));
  NAND4  g12071(.A(new_n13073_), .B(new_n13069_), .C(new_n13068_), .D(new_n13067_), .Y(new_n13074_));
  NAND2  g12072(.A(new_n13074_), .B(new_n13065_), .Y(new_n13075_));
  XOR2   g12073(.A(new_n13075_), .B(new_n13052_), .Y(new_n13076_));
  XOR2   g12074(.A(new_n13076_), .B(new_n13028_), .Y(new_n13077_));
  AOI21  g12075(.A0(new_n10103_), .A1(new_n10081_), .B0(new_n10083_), .Y(new_n13078_));
  XOR2   g12076(.A(new_n11958_), .B(new_n13078_), .Y(new_n13079_));
  OAI22  g12077(.A0(new_n11994_), .A1(new_n11993_), .B0(new_n11992_), .B1(new_n11991_), .Y(new_n13080_));
  NAND2  g12078(.A(new_n9901_), .B(new_n9862_), .Y(new_n13081_));
  AOI22  g12079(.A0(new_n11985_), .A1(new_n11984_), .B0(new_n9926_), .B1(new_n9925_), .Y(new_n13082_));
  NAND3  g12080(.A(new_n13082_), .B(new_n11989_), .C(new_n13081_), .Y(new_n13083_));
  NAND2  g12081(.A(new_n13083_), .B(new_n13080_), .Y(new_n13084_));
  XOR2   g12082(.A(new_n13084_), .B(new_n11982_), .Y(new_n13085_));
  XOR2   g12083(.A(new_n13085_), .B(new_n11961_), .Y(new_n13086_));
  OAI22  g12084(.A0(new_n13086_), .A1(new_n13079_), .B0(new_n13012_), .B1(new_n10116_), .Y(new_n13087_));
  NAND2  g12085(.A(new_n13086_), .B(new_n13079_), .Y(new_n13088_));
  NAND2  g12086(.A(new_n13088_), .B(new_n13087_), .Y(new_n13089_));
  AOI22  g12087(.A0(new_n11980_), .A1(new_n11979_), .B0(new_n11978_), .B1(new_n11977_), .Y(new_n13090_));
  NOR4   g12088(.A(new_n11974_), .B(new_n11967_), .C(new_n11964_), .D(new_n11962_), .Y(new_n13091_));
  OAI22  g12089(.A0(new_n11995_), .A1(new_n11990_), .B0(new_n13091_), .B1(new_n13090_), .Y(new_n13092_));
  NOR4   g12090(.A(new_n11995_), .B(new_n11990_), .C(new_n13091_), .D(new_n13090_), .Y(new_n13093_));
  AOI21  g12091(.A0(new_n13092_), .A1(new_n11961_), .B0(new_n13093_), .Y(new_n13094_));
  AOI221 g12092(.A0(new_n9926_), .A1(new_n9925_), .C0(new_n11987_), .B0(new_n9901_), .B1(new_n9862_), .Y(new_n13095_));
  NOR2   g12093(.A(new_n13095_), .B(new_n11988_), .Y(new_n13096_));
  NOR2   g12094(.A(new_n11984_), .B(new_n11983_), .Y(new_n13097_));
  NOR2   g12095(.A(new_n13097_), .B(new_n13096_), .Y(new_n13098_));
  NOR3   g12096(.A(new_n11965_), .B(new_n11964_), .C(new_n11962_), .Y(new_n13099_));
  OAI21  g12097(.A0(new_n11964_), .A1(new_n11962_), .B0(new_n11965_), .Y(new_n13100_));
  OAI21  g12098(.A0(new_n13099_), .A1(new_n11966_), .B0(new_n13100_), .Y(new_n13101_));
  XOR2   g12099(.A(new_n13101_), .B(new_n13098_), .Y(new_n13102_));
  NAND2  g12100(.A(new_n13092_), .B(new_n11961_), .Y(new_n13103_));
  NAND4  g12101(.A(new_n13083_), .B(new_n13080_), .C(new_n11981_), .D(new_n11975_), .Y(new_n13104_));
  OAI22  g12102(.A0(new_n13095_), .A1(new_n11988_), .B0(new_n11984_), .B1(new_n11983_), .Y(new_n13105_));
  OAI211 g12103(.A0(new_n13099_), .A1(new_n11966_), .B0(new_n13100_), .B1(new_n13105_), .Y(new_n13106_));
  NAND2  g12104(.A(new_n13101_), .B(new_n13098_), .Y(new_n13107_));
  NAND4  g12105(.A(new_n13107_), .B(new_n13106_), .C(new_n13104_), .D(new_n13103_), .Y(new_n13108_));
  OAI21  g12106(.A0(new_n13102_), .A1(new_n13094_), .B0(new_n13108_), .Y(new_n13109_));
  AOI22  g12107(.A0(new_n11941_), .A1(new_n11940_), .B0(new_n11939_), .B1(new_n11938_), .Y(new_n13110_));
  NOR4   g12108(.A(new_n11935_), .B(new_n11928_), .C(new_n11925_), .D(new_n11923_), .Y(new_n13111_));
  OAI22  g12109(.A0(new_n11956_), .A1(new_n11951_), .B0(new_n13111_), .B1(new_n13110_), .Y(new_n13112_));
  NOR4   g12110(.A(new_n11956_), .B(new_n11951_), .C(new_n13111_), .D(new_n13110_), .Y(new_n13113_));
  AOI21  g12111(.A0(new_n13112_), .A1(new_n11922_), .B0(new_n13113_), .Y(new_n13114_));
  NOR3   g12112(.A(new_n11948_), .B(new_n11953_), .C(new_n11952_), .Y(new_n13115_));
  OAI21  g12113(.A0(new_n11953_), .A1(new_n11952_), .B0(new_n11948_), .Y(new_n13116_));
  OAI21  g12114(.A0(new_n13115_), .A1(new_n11949_), .B0(new_n13116_), .Y(new_n13117_));
  NAND3  g12115(.A(new_n11930_), .B(new_n11939_), .C(new_n11938_), .Y(new_n13118_));
  AOI21  g12116(.A0(new_n11939_), .A1(new_n11938_), .B0(new_n11930_), .Y(new_n13119_));
  AOI21  g12117(.A0(new_n13118_), .A1(new_n11934_), .B0(new_n13119_), .Y(new_n13120_));
  XOR2   g12118(.A(new_n13120_), .B(new_n13117_), .Y(new_n13121_));
  NAND2  g12119(.A(new_n13112_), .B(new_n11922_), .Y(new_n13122_));
  AOI21  g12120(.A0(new_n13120_), .A1(new_n13117_), .B0(new_n13113_), .Y(new_n13123_));
  OAI211 g12121(.A0(new_n13120_), .A1(new_n13117_), .B0(new_n13123_), .B1(new_n13122_), .Y(new_n13124_));
  OAI21  g12122(.A0(new_n13121_), .A1(new_n13114_), .B0(new_n13124_), .Y(new_n13125_));
  XOR2   g12123(.A(new_n13125_), .B(new_n13109_), .Y(new_n13126_));
  XOR2   g12124(.A(new_n13126_), .B(new_n13089_), .Y(new_n13127_));
  XOR2   g12125(.A(new_n13127_), .B(new_n13077_), .Y(new_n13128_));
  XOR2   g12126(.A(new_n13128_), .B(new_n13019_), .Y(new_n13129_));
  XOR2   g12127(.A(new_n13129_), .B(new_n13011_), .Y(new_n13130_));
  XOR2   g12128(.A(new_n13130_), .B(new_n12903_), .Y(new_n13131_));
  OAI21  g12129(.A0(new_n11175_), .A1(new_n9105_), .B0(new_n9107_), .Y(new_n13132_));
  AOI21  g12130(.A0(new_n9102_), .A1(new_n9093_), .B0(new_n9095_), .Y(new_n13133_));
  XOR2   g12131(.A(new_n11765_), .B(new_n13133_), .Y(new_n13134_));
  AOI21  g12132(.A0(new_n8402_), .A1(new_n8066_), .B0(new_n8068_), .Y(new_n13135_));
  XOR2   g12133(.A(new_n11915_), .B(new_n13135_), .Y(new_n13136_));
  NAND2  g12134(.A(new_n13136_), .B(new_n13134_), .Y(new_n13137_));
  NOR2   g12135(.A(new_n13136_), .B(new_n13134_), .Y(new_n13138_));
  AOI21  g12136(.A0(new_n13137_), .A1(new_n13132_), .B0(new_n13138_), .Y(new_n13139_));
  NOR2   g12137(.A(new_n11914_), .B(new_n11841_), .Y(new_n13140_));
  NAND2  g12138(.A(new_n11914_), .B(new_n11841_), .Y(new_n13141_));
  OAI21  g12139(.A0(new_n13140_), .A1(new_n13135_), .B0(new_n13141_), .Y(new_n13142_));
  OAI22  g12140(.A0(new_n11874_), .A1(new_n11873_), .B0(new_n11872_), .B1(new_n7782_), .Y(new_n13143_));
  NAND2  g12141(.A(new_n7647_), .B(new_n7583_), .Y(new_n13144_));
  NAND4  g12142(.A(new_n11870_), .B(new_n11867_), .C(new_n13144_), .D(new_n7650_), .Y(new_n13145_));
  NAND2  g12143(.A(new_n13145_), .B(new_n13143_), .Y(new_n13146_));
  XOR2   g12144(.A(new_n13146_), .B(new_n11862_), .Y(new_n13147_));
  XOR2   g12145(.A(new_n13147_), .B(new_n11845_), .Y(new_n13148_));
  OAI22  g12146(.A0(new_n11912_), .A1(new_n13148_), .B0(new_n11842_), .B1(new_n8056_), .Y(new_n13149_));
  NAND2  g12147(.A(new_n11912_), .B(new_n13148_), .Y(new_n13150_));
  NAND2  g12148(.A(new_n13150_), .B(new_n13149_), .Y(new_n13151_));
  NOR2   g12149(.A(new_n8013_), .B(new_n8011_), .Y(new_n13152_));
  OAI22  g12150(.A0(new_n8021_), .A1(new_n7977_), .B0(new_n7882_), .B1(new_n13152_), .Y(new_n13153_));
  AOI22  g12151(.A0(new_n11910_), .A1(new_n11896_), .B0(new_n13153_), .B1(new_n8022_), .Y(new_n13154_));
  AOI22  g12152(.A0(new_n11894_), .A1(new_n11893_), .B0(new_n11892_), .B1(new_n7881_), .Y(new_n13155_));
  NOR4   g12153(.A(new_n11890_), .B(new_n11887_), .C(new_n11884_), .D(new_n11883_), .Y(new_n13156_));
  AOI21  g12154(.A0(new_n7983_), .A1(new_n7919_), .B0(new_n8019_), .Y(new_n13157_));
  AOI21  g12155(.A0(new_n11908_), .A1(new_n11907_), .B0(new_n13157_), .Y(new_n13158_));
  NOR4   g12156(.A(new_n11904_), .B(new_n11900_), .C(new_n11897_), .D(new_n8019_), .Y(new_n13159_));
  NOR4   g12157(.A(new_n13159_), .B(new_n13158_), .C(new_n13156_), .D(new_n13155_), .Y(new_n13160_));
  AOI211 g12158(.A0(new_n7983_), .A1(new_n7919_), .B(new_n11898_), .C(new_n8019_), .Y(new_n13161_));
  OAI22  g12159(.A0(new_n13161_), .A1(new_n11899_), .B0(new_n11902_), .B1(new_n13157_), .Y(new_n13162_));
  NOR3   g12160(.A(new_n11885_), .B(new_n11884_), .C(new_n11883_), .Y(new_n13163_));
  OAI21  g12161(.A0(new_n11884_), .A1(new_n11883_), .B0(new_n11885_), .Y(new_n13164_));
  OAI21  g12162(.A0(new_n13163_), .A1(new_n11886_), .B0(new_n13164_), .Y(new_n13165_));
  XOR2   g12163(.A(new_n13165_), .B(new_n13162_), .Y(new_n13166_));
  OAI21  g12164(.A0(new_n13160_), .A1(new_n13154_), .B0(new_n13166_), .Y(new_n13167_));
  OAI22  g12165(.A0(new_n13159_), .A1(new_n13158_), .B0(new_n13156_), .B1(new_n13155_), .Y(new_n13168_));
  NAND2  g12166(.A(new_n13168_), .B(new_n11880_), .Y(new_n13169_));
  NAND3  g12167(.A(new_n11888_), .B(new_n11892_), .C(new_n7881_), .Y(new_n13170_));
  AOI21  g12168(.A0(new_n11892_), .A1(new_n7881_), .B0(new_n11888_), .Y(new_n13171_));
  AOI21  g12169(.A0(new_n13170_), .A1(new_n11889_), .B0(new_n13171_), .Y(new_n13172_));
  AOI21  g12170(.A0(new_n13172_), .A1(new_n13162_), .B0(new_n13160_), .Y(new_n13173_));
  OAI211 g12171(.A0(new_n13172_), .A1(new_n13162_), .B0(new_n13173_), .B1(new_n13169_), .Y(new_n13174_));
  NAND2  g12172(.A(new_n13174_), .B(new_n13167_), .Y(new_n13175_));
  AOI21  g12173(.A0(new_n11857_), .A1(new_n7764_), .B0(new_n7774_), .Y(new_n13176_));
  OAI22  g12174(.A0(new_n7784_), .A1(new_n7641_), .B0(new_n13176_), .B1(new_n7763_), .Y(new_n13177_));
  AOI22  g12175(.A0(new_n13146_), .A1(new_n11862_), .B0(new_n13177_), .B1(new_n7785_), .Y(new_n13178_));
  AOI22  g12176(.A0(new_n11860_), .A1(new_n11859_), .B0(new_n11858_), .B1(new_n11857_), .Y(new_n13179_));
  NOR4   g12177(.A(new_n11854_), .B(new_n11850_), .C(new_n11847_), .D(new_n11846_), .Y(new_n13180_));
  NOR4   g12178(.A(new_n11875_), .B(new_n11871_), .C(new_n13180_), .D(new_n13179_), .Y(new_n13181_));
  AOI211 g12179(.A0(new_n7647_), .A1(new_n7583_), .B(new_n11868_), .C(new_n7782_), .Y(new_n13182_));
  OAI22  g12180(.A0(new_n13182_), .A1(new_n11869_), .B0(new_n11865_), .B1(new_n11863_), .Y(new_n13183_));
  NOR3   g12181(.A(new_n11848_), .B(new_n11847_), .C(new_n11846_), .Y(new_n13184_));
  OAI21  g12182(.A0(new_n11847_), .A1(new_n11846_), .B0(new_n11848_), .Y(new_n13185_));
  OAI21  g12183(.A0(new_n13184_), .A1(new_n11849_), .B0(new_n13185_), .Y(new_n13186_));
  XOR2   g12184(.A(new_n13186_), .B(new_n13183_), .Y(new_n13187_));
  OAI21  g12185(.A0(new_n13181_), .A1(new_n13178_), .B0(new_n13187_), .Y(new_n13188_));
  OAI22  g12186(.A0(new_n11875_), .A1(new_n11871_), .B0(new_n13180_), .B1(new_n13179_), .Y(new_n13189_));
  NAND2  g12187(.A(new_n13189_), .B(new_n11845_), .Y(new_n13190_));
  NAND4  g12188(.A(new_n13145_), .B(new_n13143_), .C(new_n11861_), .D(new_n11855_), .Y(new_n13191_));
  OAI211 g12189(.A0(new_n13184_), .A1(new_n11849_), .B0(new_n13185_), .B1(new_n13183_), .Y(new_n13192_));
  NOR2   g12190(.A(new_n13182_), .B(new_n11869_), .Y(new_n13193_));
  NOR2   g12191(.A(new_n11865_), .B(new_n11863_), .Y(new_n13194_));
  NOR2   g12192(.A(new_n13194_), .B(new_n13193_), .Y(new_n13195_));
  NAND2  g12193(.A(new_n13186_), .B(new_n13195_), .Y(new_n13196_));
  NAND4  g12194(.A(new_n13196_), .B(new_n13192_), .C(new_n13191_), .D(new_n13190_), .Y(new_n13197_));
  NAND2  g12195(.A(new_n13197_), .B(new_n13188_), .Y(new_n13198_));
  XOR2   g12196(.A(new_n13198_), .B(new_n13175_), .Y(new_n13199_));
  XOR2   g12197(.A(new_n13199_), .B(new_n13151_), .Y(new_n13200_));
  NAND2  g12198(.A(new_n11839_), .B(new_n11806_), .Y(new_n13201_));
  NOR2   g12199(.A(new_n11839_), .B(new_n11806_), .Y(new_n13202_));
  AOI21  g12200(.A0(new_n13201_), .A1(new_n11768_), .B0(new_n13202_), .Y(new_n13203_));
  AOI22  g12201(.A0(new_n11821_), .A1(new_n11820_), .B0(new_n11819_), .B1(new_n7151_), .Y(new_n13204_));
  NOR4   g12202(.A(new_n11817_), .B(new_n11814_), .C(new_n11809_), .D(new_n7281_), .Y(new_n13205_));
  OAI22  g12203(.A0(new_n11836_), .A1(new_n11832_), .B0(new_n13205_), .B1(new_n13204_), .Y(new_n13206_));
  NOR4   g12204(.A(new_n11836_), .B(new_n11832_), .C(new_n13205_), .D(new_n13204_), .Y(new_n13207_));
  AOI21  g12205(.A0(new_n13206_), .A1(new_n11808_), .B0(new_n13207_), .Y(new_n13208_));
  AOI211 g12206(.A0(new_n7253_), .A1(new_n7189_), .B(new_n11829_), .C(new_n7286_), .Y(new_n13209_));
  OAI22  g12207(.A0(new_n13209_), .A1(new_n11830_), .B0(new_n11826_), .B1(new_n11824_), .Y(new_n13210_));
  NAND3  g12208(.A(new_n11815_), .B(new_n11819_), .C(new_n7151_), .Y(new_n13211_));
  AOI21  g12209(.A0(new_n11819_), .A1(new_n7151_), .B0(new_n11815_), .Y(new_n13212_));
  AOI21  g12210(.A0(new_n13211_), .A1(new_n11816_), .B0(new_n13212_), .Y(new_n13213_));
  XOR2   g12211(.A(new_n13213_), .B(new_n13210_), .Y(new_n13214_));
  NAND2  g12212(.A(new_n13206_), .B(new_n11808_), .Y(new_n13215_));
  AOI21  g12213(.A0(new_n13213_), .A1(new_n13210_), .B0(new_n13207_), .Y(new_n13216_));
  OAI211 g12214(.A0(new_n13213_), .A1(new_n13210_), .B0(new_n13216_), .B1(new_n13215_), .Y(new_n13217_));
  OAI21  g12215(.A0(new_n13214_), .A1(new_n13208_), .B0(new_n13217_), .Y(new_n13218_));
  AOI22  g12216(.A0(new_n11788_), .A1(new_n11787_), .B0(new_n11786_), .B1(new_n11785_), .Y(new_n13219_));
  NOR4   g12217(.A(new_n11782_), .B(new_n11775_), .C(new_n11772_), .D(new_n11770_), .Y(new_n13220_));
  OAI22  g12218(.A0(new_n11803_), .A1(new_n11798_), .B0(new_n13220_), .B1(new_n13219_), .Y(new_n13221_));
  NOR4   g12219(.A(new_n11803_), .B(new_n11798_), .C(new_n13220_), .D(new_n13219_), .Y(new_n13222_));
  AOI21  g12220(.A0(new_n13221_), .A1(new_n11769_), .B0(new_n13222_), .Y(new_n13223_));
  NOR3   g12221(.A(new_n11795_), .B(new_n11800_), .C(new_n11799_), .Y(new_n13224_));
  OAI21  g12222(.A0(new_n11800_), .A1(new_n11799_), .B0(new_n11795_), .Y(new_n13225_));
  OAI21  g12223(.A0(new_n13224_), .A1(new_n11796_), .B0(new_n13225_), .Y(new_n13226_));
  NAND3  g12224(.A(new_n11777_), .B(new_n11786_), .C(new_n11785_), .Y(new_n13227_));
  AOI21  g12225(.A0(new_n11786_), .A1(new_n11785_), .B0(new_n11777_), .Y(new_n13228_));
  AOI21  g12226(.A0(new_n13227_), .A1(new_n11781_), .B0(new_n13228_), .Y(new_n13229_));
  XOR2   g12227(.A(new_n13229_), .B(new_n13226_), .Y(new_n13230_));
  NOR2   g12228(.A(new_n13230_), .B(new_n13223_), .Y(new_n13231_));
  NAND3  g12229(.A(new_n11792_), .B(new_n11791_), .C(new_n7536_), .Y(new_n13232_));
  AOI21  g12230(.A0(new_n11791_), .A1(new_n7536_), .B0(new_n11792_), .Y(new_n13233_));
  AOI21  g12231(.A0(new_n13232_), .A1(new_n11793_), .B0(new_n13233_), .Y(new_n13234_));
  NOR3   g12232(.A(new_n11773_), .B(new_n11772_), .C(new_n11770_), .Y(new_n13235_));
  OAI21  g12233(.A0(new_n11772_), .A1(new_n11770_), .B0(new_n11773_), .Y(new_n13236_));
  OAI21  g12234(.A0(new_n13235_), .A1(new_n11774_), .B0(new_n13236_), .Y(new_n13237_));
  NAND4  g12235(.A(new_n11797_), .B(new_n11794_), .C(new_n11791_), .D(new_n7536_), .Y(new_n13238_));
  NAND3  g12236(.A(new_n13238_), .B(new_n11789_), .C(new_n11783_), .Y(new_n13239_));
  OAI22  g12237(.A0(new_n13237_), .A1(new_n13234_), .B0(new_n13239_), .B1(new_n11798_), .Y(new_n13240_));
  AOI221 g12238(.A0(new_n13237_), .A1(new_n13234_), .C0(new_n13240_), .B0(new_n13221_), .B1(new_n11769_), .Y(new_n13241_));
  NOR2   g12239(.A(new_n13241_), .B(new_n13231_), .Y(new_n13242_));
  XOR2   g12240(.A(new_n13242_), .B(new_n13218_), .Y(new_n13243_));
  XOR2   g12241(.A(new_n13243_), .B(new_n13203_), .Y(new_n13244_));
  XOR2   g12242(.A(new_n13244_), .B(new_n13200_), .Y(new_n13245_));
  XOR2   g12243(.A(new_n13245_), .B(new_n13142_), .Y(new_n13246_));
  AOI22  g12244(.A0(new_n9081_), .A1(new_n8889_), .B0(new_n9059_), .B1(new_n9053_), .Y(new_n13247_));
  NOR2   g12245(.A(new_n13247_), .B(new_n9091_), .Y(new_n13248_));
  XOR2   g12246(.A(new_n11690_), .B(new_n13248_), .Y(new_n13249_));
  AOI22  g12247(.A0(new_n8742_), .A1(new_n8696_), .B0(new_n8562_), .B1(new_n8539_), .Y(new_n13250_));
  NOR2   g12248(.A(new_n13250_), .B(new_n8753_), .Y(new_n13251_));
  XOR2   g12249(.A(new_n11763_), .B(new_n13251_), .Y(new_n13252_));
  NAND2  g12250(.A(new_n13252_), .B(new_n13249_), .Y(new_n13253_));
  NOR2   g12251(.A(new_n13252_), .B(new_n13249_), .Y(new_n13254_));
  AOI21  g12252(.A0(new_n13253_), .A1(new_n11611_), .B0(new_n13254_), .Y(new_n13255_));
  OAI22  g12253(.A0(new_n11723_), .A1(new_n11722_), .B0(new_n11721_), .B1(new_n11720_), .Y(new_n13256_));
  NAND2  g12254(.A(new_n8465_), .B(new_n8426_), .Y(new_n13257_));
  AOI22  g12255(.A0(new_n11714_), .A1(new_n11713_), .B0(new_n8558_), .B1(new_n8557_), .Y(new_n13258_));
  NAND3  g12256(.A(new_n13258_), .B(new_n11718_), .C(new_n13257_), .Y(new_n13259_));
  NAND2  g12257(.A(new_n13259_), .B(new_n13256_), .Y(new_n13260_));
  XOR2   g12258(.A(new_n13260_), .B(new_n11711_), .Y(new_n13261_));
  XOR2   g12259(.A(new_n13261_), .B(new_n11694_), .Y(new_n13262_));
  OAI22  g12260(.A0(new_n11758_), .A1(new_n11757_), .B0(new_n11756_), .B1(new_n11755_), .Y(new_n13263_));
  NAND2  g12261(.A(new_n8683_), .B(new_n8644_), .Y(new_n13264_));
  AOI22  g12262(.A0(new_n11749_), .A1(new_n11748_), .B0(new_n8715_), .B1(new_n8714_), .Y(new_n13265_));
  NAND3  g12263(.A(new_n13265_), .B(new_n11753_), .C(new_n13264_), .Y(new_n13266_));
  NAND2  g12264(.A(new_n13266_), .B(new_n13263_), .Y(new_n13267_));
  XOR2   g12265(.A(new_n13267_), .B(new_n11746_), .Y(new_n13268_));
  XOR2   g12266(.A(new_n13268_), .B(new_n11729_), .Y(new_n13269_));
  OAI22  g12267(.A0(new_n13269_), .A1(new_n13262_), .B0(new_n13250_), .B1(new_n8753_), .Y(new_n13270_));
  NAND2  g12268(.A(new_n13269_), .B(new_n13262_), .Y(new_n13271_));
  NAND2  g12269(.A(new_n13271_), .B(new_n13270_), .Y(new_n13272_));
  AOI21  g12270(.A0(new_n11741_), .A1(new_n8620_), .B0(new_n8701_), .Y(new_n13273_));
  OAI22  g12271(.A0(new_n8717_), .A1(new_n8682_), .B0(new_n13273_), .B1(new_n8619_), .Y(new_n13274_));
  AOI22  g12272(.A0(new_n13267_), .A1(new_n11746_), .B0(new_n13274_), .B1(new_n8730_), .Y(new_n13275_));
  AOI22  g12273(.A0(new_n11744_), .A1(new_n11743_), .B0(new_n11742_), .B1(new_n11741_), .Y(new_n13276_));
  NOR4   g12274(.A(new_n11738_), .B(new_n11734_), .C(new_n11731_), .D(new_n11730_), .Y(new_n13277_));
  NOR4   g12275(.A(new_n11759_), .B(new_n11754_), .C(new_n13277_), .D(new_n13276_), .Y(new_n13278_));
  AOI221 g12276(.A0(new_n8715_), .A1(new_n8714_), .C0(new_n11751_), .B0(new_n8683_), .B1(new_n8644_), .Y(new_n13279_));
  OAI22  g12277(.A0(new_n13279_), .A1(new_n11752_), .B0(new_n11748_), .B1(new_n11747_), .Y(new_n13280_));
  NOR3   g12278(.A(new_n11732_), .B(new_n11731_), .C(new_n11730_), .Y(new_n13281_));
  OAI21  g12279(.A0(new_n11731_), .A1(new_n11730_), .B0(new_n11732_), .Y(new_n13282_));
  OAI21  g12280(.A0(new_n13281_), .A1(new_n11733_), .B0(new_n13282_), .Y(new_n13283_));
  XOR2   g12281(.A(new_n13283_), .B(new_n13280_), .Y(new_n13284_));
  OAI21  g12282(.A0(new_n13278_), .A1(new_n13275_), .B0(new_n13284_), .Y(new_n13285_));
  OAI22  g12283(.A0(new_n11759_), .A1(new_n11754_), .B0(new_n13277_), .B1(new_n13276_), .Y(new_n13286_));
  NAND2  g12284(.A(new_n13286_), .B(new_n11729_), .Y(new_n13287_));
  NAND4  g12285(.A(new_n13266_), .B(new_n13263_), .C(new_n11745_), .D(new_n11739_), .Y(new_n13288_));
  OAI211 g12286(.A0(new_n13281_), .A1(new_n11733_), .B0(new_n13282_), .B1(new_n13280_), .Y(new_n13289_));
  NOR2   g12287(.A(new_n13279_), .B(new_n11752_), .Y(new_n13290_));
  NOR2   g12288(.A(new_n11748_), .B(new_n11747_), .Y(new_n13291_));
  NOR2   g12289(.A(new_n13291_), .B(new_n13290_), .Y(new_n13292_));
  NAND2  g12290(.A(new_n13283_), .B(new_n13292_), .Y(new_n13293_));
  NAND4  g12291(.A(new_n13293_), .B(new_n13289_), .C(new_n13288_), .D(new_n13287_), .Y(new_n13294_));
  NAND2  g12292(.A(new_n13294_), .B(new_n13285_), .Y(new_n13295_));
  OAI21  g12293(.A0(new_n8738_), .A1(new_n8464_), .B0(new_n8478_), .Y(new_n13296_));
  AOI21  g12294(.A0(new_n11706_), .A1(new_n8534_), .B0(new_n8544_), .Y(new_n13297_));
  OAI22  g12295(.A0(new_n8560_), .A1(new_n8464_), .B0(new_n13297_), .B1(new_n8533_), .Y(new_n13298_));
  AOI22  g12296(.A0(new_n13260_), .A1(new_n11711_), .B0(new_n13298_), .B1(new_n13296_), .Y(new_n13299_));
  AOI22  g12297(.A0(new_n11709_), .A1(new_n11708_), .B0(new_n11707_), .B1(new_n11706_), .Y(new_n13300_));
  NOR4   g12298(.A(new_n11703_), .B(new_n11699_), .C(new_n11696_), .D(new_n11695_), .Y(new_n13301_));
  NOR4   g12299(.A(new_n11724_), .B(new_n11719_), .C(new_n13301_), .D(new_n13300_), .Y(new_n13302_));
  AOI221 g12300(.A0(new_n8558_), .A1(new_n8557_), .C0(new_n11716_), .B0(new_n8465_), .B1(new_n8426_), .Y(new_n13303_));
  OAI22  g12301(.A0(new_n13303_), .A1(new_n11717_), .B0(new_n11713_), .B1(new_n11712_), .Y(new_n13304_));
  NOR3   g12302(.A(new_n11697_), .B(new_n11696_), .C(new_n11695_), .Y(new_n13305_));
  OAI21  g12303(.A0(new_n11696_), .A1(new_n11695_), .B0(new_n11697_), .Y(new_n13306_));
  OAI21  g12304(.A0(new_n13305_), .A1(new_n11698_), .B0(new_n13306_), .Y(new_n13307_));
  XOR2   g12305(.A(new_n13307_), .B(new_n13304_), .Y(new_n13308_));
  OAI21  g12306(.A0(new_n13302_), .A1(new_n13299_), .B0(new_n13308_), .Y(new_n13309_));
  OAI22  g12307(.A0(new_n11724_), .A1(new_n11719_), .B0(new_n13301_), .B1(new_n13300_), .Y(new_n13310_));
  NAND2  g12308(.A(new_n13310_), .B(new_n11694_), .Y(new_n13311_));
  NAND4  g12309(.A(new_n13259_), .B(new_n13256_), .C(new_n11710_), .D(new_n11704_), .Y(new_n13312_));
  OAI211 g12310(.A0(new_n13305_), .A1(new_n11698_), .B0(new_n13306_), .B1(new_n13304_), .Y(new_n13313_));
  NOR2   g12311(.A(new_n13303_), .B(new_n11717_), .Y(new_n13314_));
  NOR2   g12312(.A(new_n11713_), .B(new_n11712_), .Y(new_n13315_));
  NOR2   g12313(.A(new_n13315_), .B(new_n13314_), .Y(new_n13316_));
  NAND2  g12314(.A(new_n13307_), .B(new_n13316_), .Y(new_n13317_));
  NAND4  g12315(.A(new_n13317_), .B(new_n13313_), .C(new_n13312_), .D(new_n13311_), .Y(new_n13318_));
  NAND2  g12316(.A(new_n13318_), .B(new_n13309_), .Y(new_n13319_));
  XOR2   g12317(.A(new_n13319_), .B(new_n13295_), .Y(new_n13320_));
  XOR2   g12318(.A(new_n13320_), .B(new_n13272_), .Y(new_n13321_));
  AOI21  g12319(.A0(new_n9078_), .A1(new_n9056_), .B0(new_n9058_), .Y(new_n13322_));
  XOR2   g12320(.A(new_n11649_), .B(new_n13322_), .Y(new_n13323_));
  OAI22  g12321(.A0(new_n11685_), .A1(new_n11684_), .B0(new_n11683_), .B1(new_n11682_), .Y(new_n13324_));
  NAND2  g12322(.A(new_n8876_), .B(new_n8837_), .Y(new_n13325_));
  AOI22  g12323(.A0(new_n11676_), .A1(new_n11675_), .B0(new_n8901_), .B1(new_n8900_), .Y(new_n13326_));
  NAND3  g12324(.A(new_n13326_), .B(new_n11680_), .C(new_n13325_), .Y(new_n13327_));
  NAND2  g12325(.A(new_n13327_), .B(new_n13324_), .Y(new_n13328_));
  XOR2   g12326(.A(new_n13328_), .B(new_n11673_), .Y(new_n13329_));
  XOR2   g12327(.A(new_n13329_), .B(new_n11652_), .Y(new_n13330_));
  OAI22  g12328(.A0(new_n13330_), .A1(new_n13323_), .B0(new_n13247_), .B1(new_n9091_), .Y(new_n13331_));
  NAND2  g12329(.A(new_n13330_), .B(new_n13323_), .Y(new_n13332_));
  NAND2  g12330(.A(new_n13332_), .B(new_n13331_), .Y(new_n13333_));
  AOI22  g12331(.A0(new_n11671_), .A1(new_n11670_), .B0(new_n11669_), .B1(new_n11668_), .Y(new_n13334_));
  NOR4   g12332(.A(new_n11665_), .B(new_n11658_), .C(new_n11655_), .D(new_n11653_), .Y(new_n13335_));
  OAI22  g12333(.A0(new_n11686_), .A1(new_n11681_), .B0(new_n13335_), .B1(new_n13334_), .Y(new_n13336_));
  NOR4   g12334(.A(new_n11686_), .B(new_n11681_), .C(new_n13335_), .D(new_n13334_), .Y(new_n13337_));
  AOI21  g12335(.A0(new_n13336_), .A1(new_n11652_), .B0(new_n13337_), .Y(new_n13338_));
  AOI221 g12336(.A0(new_n8901_), .A1(new_n8900_), .C0(new_n11678_), .B0(new_n8876_), .B1(new_n8837_), .Y(new_n13339_));
  NOR2   g12337(.A(new_n13339_), .B(new_n11679_), .Y(new_n13340_));
  NOR2   g12338(.A(new_n11675_), .B(new_n11674_), .Y(new_n13341_));
  NOR2   g12339(.A(new_n13341_), .B(new_n13340_), .Y(new_n13342_));
  NOR3   g12340(.A(new_n11656_), .B(new_n11655_), .C(new_n11653_), .Y(new_n13343_));
  OAI21  g12341(.A0(new_n11655_), .A1(new_n11653_), .B0(new_n11656_), .Y(new_n13344_));
  OAI21  g12342(.A0(new_n13343_), .A1(new_n11657_), .B0(new_n13344_), .Y(new_n13345_));
  XOR2   g12343(.A(new_n13345_), .B(new_n13342_), .Y(new_n13346_));
  NAND2  g12344(.A(new_n13336_), .B(new_n11652_), .Y(new_n13347_));
  NAND4  g12345(.A(new_n13327_), .B(new_n13324_), .C(new_n11672_), .D(new_n11666_), .Y(new_n13348_));
  OAI22  g12346(.A0(new_n13339_), .A1(new_n11679_), .B0(new_n11675_), .B1(new_n11674_), .Y(new_n13349_));
  OAI211 g12347(.A0(new_n13343_), .A1(new_n11657_), .B0(new_n13344_), .B1(new_n13349_), .Y(new_n13350_));
  NAND2  g12348(.A(new_n13345_), .B(new_n13342_), .Y(new_n13351_));
  NAND4  g12349(.A(new_n13351_), .B(new_n13350_), .C(new_n13348_), .D(new_n13347_), .Y(new_n13352_));
  OAI21  g12350(.A0(new_n13346_), .A1(new_n13338_), .B0(new_n13352_), .Y(new_n13353_));
  AOI22  g12351(.A0(new_n11632_), .A1(new_n11631_), .B0(new_n11630_), .B1(new_n11629_), .Y(new_n13354_));
  NOR4   g12352(.A(new_n11626_), .B(new_n11619_), .C(new_n11616_), .D(new_n11614_), .Y(new_n13355_));
  OAI22  g12353(.A0(new_n11647_), .A1(new_n11642_), .B0(new_n13355_), .B1(new_n13354_), .Y(new_n13356_));
  NOR4   g12354(.A(new_n11647_), .B(new_n11642_), .C(new_n13355_), .D(new_n13354_), .Y(new_n13357_));
  AOI21  g12355(.A0(new_n13356_), .A1(new_n11613_), .B0(new_n13357_), .Y(new_n13358_));
  NOR3   g12356(.A(new_n11639_), .B(new_n11644_), .C(new_n11643_), .Y(new_n13359_));
  OAI21  g12357(.A0(new_n11644_), .A1(new_n11643_), .B0(new_n11639_), .Y(new_n13360_));
  OAI21  g12358(.A0(new_n13359_), .A1(new_n11640_), .B0(new_n13360_), .Y(new_n13361_));
  NAND3  g12359(.A(new_n11621_), .B(new_n11630_), .C(new_n11629_), .Y(new_n13362_));
  AOI21  g12360(.A0(new_n11630_), .A1(new_n11629_), .B0(new_n11621_), .Y(new_n13363_));
  AOI21  g12361(.A0(new_n13362_), .A1(new_n11625_), .B0(new_n13363_), .Y(new_n13364_));
  XOR2   g12362(.A(new_n13364_), .B(new_n13361_), .Y(new_n13365_));
  NAND2  g12363(.A(new_n13356_), .B(new_n11613_), .Y(new_n13366_));
  AOI21  g12364(.A0(new_n13364_), .A1(new_n13361_), .B0(new_n13357_), .Y(new_n13367_));
  OAI211 g12365(.A0(new_n13364_), .A1(new_n13361_), .B0(new_n13367_), .B1(new_n13366_), .Y(new_n13368_));
  OAI21  g12366(.A0(new_n13365_), .A1(new_n13358_), .B0(new_n13368_), .Y(new_n13369_));
  XOR2   g12367(.A(new_n13369_), .B(new_n13353_), .Y(new_n13370_));
  XOR2   g12368(.A(new_n13370_), .B(new_n13333_), .Y(new_n13371_));
  XOR2   g12369(.A(new_n13371_), .B(new_n13321_), .Y(new_n13372_));
  XOR2   g12370(.A(new_n13372_), .B(new_n13255_), .Y(new_n13373_));
  XOR2   g12371(.A(new_n13373_), .B(new_n13246_), .Y(new_n13374_));
  XOR2   g12372(.A(new_n13374_), .B(new_n13139_), .Y(new_n13375_));
  XOR2   g12373(.A(new_n13375_), .B(new_n13131_), .Y(new_n13376_));
  XOR2   g12374(.A(new_n13376_), .B(new_n12900_), .Y(new_n13377_));
  NOR2   g12375(.A(new_n11604_), .B(new_n11598_), .Y(new_n13378_));
  OAI21  g12376(.A0(new_n13378_), .A1(new_n11444_), .B0(new_n11597_), .Y(new_n13379_));
  OAI21  g12377(.A0(new_n7051_), .A1(new_n7037_), .B0(new_n7039_), .Y(new_n13380_));
  XOR2   g12378(.A(new_n11596_), .B(new_n13380_), .Y(new_n13381_));
  OAI21  g12379(.A0(new_n11604_), .A1(new_n11598_), .B0(new_n13381_), .Y(new_n13382_));
  NOR2   g12380(.A(new_n13382_), .B(new_n11444_), .Y(new_n13383_));
  AOI21  g12381(.A0(new_n13379_), .A1(new_n11220_), .B0(new_n13383_), .Y(new_n13384_));
  NAND2  g12382(.A(new_n11442_), .B(new_n11601_), .Y(new_n13385_));
  OAI21  g12383(.A0(new_n11363_), .A1(new_n11222_), .B0(new_n11436_), .Y(new_n13386_));
  NOR2   g12384(.A(new_n13386_), .B(new_n11599_), .Y(new_n13387_));
  AOI21  g12385(.A0(new_n13385_), .A1(new_n11598_), .B0(new_n13387_), .Y(new_n13388_));
  NOR2   g12386(.A(new_n11362_), .B(new_n11285_), .Y(new_n13389_));
  NAND2  g12387(.A(new_n11362_), .B(new_n11285_), .Y(new_n13390_));
  OAI21  g12388(.A0(new_n13389_), .A1(new_n11437_), .B0(new_n13390_), .Y(new_n13391_));
  AOI21  g12389(.A0(new_n6049_), .A1(new_n5796_), .B0(new_n5798_), .Y(new_n13392_));
  XOR2   g12390(.A(new_n11326_), .B(new_n13392_), .Y(new_n13393_));
  OAI22  g12391(.A0(new_n11360_), .A1(new_n13393_), .B0(new_n11286_), .B1(new_n6069_), .Y(new_n13394_));
  NAND2  g12392(.A(new_n11360_), .B(new_n13393_), .Y(new_n13395_));
  NAND2  g12393(.A(new_n13395_), .B(new_n13394_), .Y(new_n13396_));
  AOI22  g12394(.A0(new_n11342_), .A1(new_n11341_), .B0(new_n11340_), .B1(new_n5893_), .Y(new_n13397_));
  NOR4   g12395(.A(new_n11338_), .B(new_n11335_), .C(new_n11330_), .D(new_n6023_), .Y(new_n13398_));
  AOI21  g12396(.A0(new_n5995_), .A1(new_n5931_), .B0(new_n6028_), .Y(new_n13399_));
  AOI21  g12397(.A0(new_n11356_), .A1(new_n11355_), .B0(new_n13399_), .Y(new_n13400_));
  NOR4   g12398(.A(new_n11352_), .B(new_n11348_), .C(new_n11345_), .D(new_n6028_), .Y(new_n13401_));
  OAI22  g12399(.A0(new_n13401_), .A1(new_n13400_), .B0(new_n13398_), .B1(new_n13397_), .Y(new_n13402_));
  NOR4   g12400(.A(new_n13401_), .B(new_n13400_), .C(new_n13398_), .D(new_n13397_), .Y(new_n13403_));
  AOI21  g12401(.A0(new_n13402_), .A1(new_n11329_), .B0(new_n13403_), .Y(new_n13404_));
  AOI211 g12402(.A0(new_n5995_), .A1(new_n5931_), .B(new_n11346_), .C(new_n6028_), .Y(new_n13405_));
  OAI22  g12403(.A0(new_n13405_), .A1(new_n11347_), .B0(new_n11350_), .B1(new_n13399_), .Y(new_n13406_));
  NAND3  g12404(.A(new_n11336_), .B(new_n11340_), .C(new_n5893_), .Y(new_n13407_));
  AOI21  g12405(.A0(new_n11340_), .A1(new_n5893_), .B0(new_n11336_), .Y(new_n13408_));
  AOI21  g12406(.A0(new_n13407_), .A1(new_n11337_), .B0(new_n13408_), .Y(new_n13409_));
  XOR2   g12407(.A(new_n13409_), .B(new_n13406_), .Y(new_n13410_));
  NAND2  g12408(.A(new_n13402_), .B(new_n11329_), .Y(new_n13411_));
  AOI21  g12409(.A0(new_n13409_), .A1(new_n13406_), .B0(new_n13403_), .Y(new_n13412_));
  OAI211 g12410(.A0(new_n13409_), .A1(new_n13406_), .B0(new_n13412_), .B1(new_n13411_), .Y(new_n13413_));
  OAI21  g12411(.A0(new_n13410_), .A1(new_n13404_), .B0(new_n13413_), .Y(new_n13414_));
  AOI22  g12412(.A0(new_n11307_), .A1(new_n11306_), .B0(new_n11305_), .B1(new_n11304_), .Y(new_n13415_));
  NOR4   g12413(.A(new_n11301_), .B(new_n11294_), .C(new_n11291_), .D(new_n11289_), .Y(new_n13416_));
  OAI22  g12414(.A0(new_n11324_), .A1(new_n11318_), .B0(new_n13416_), .B1(new_n13415_), .Y(new_n13417_));
  NOR4   g12415(.A(new_n11324_), .B(new_n11318_), .C(new_n13416_), .D(new_n13415_), .Y(new_n13418_));
  AOI21  g12416(.A0(new_n13417_), .A1(new_n11288_), .B0(new_n13418_), .Y(new_n13419_));
  NOR3   g12417(.A(new_n11315_), .B(new_n11321_), .C(new_n11320_), .Y(new_n13420_));
  OAI21  g12418(.A0(new_n11321_), .A1(new_n11320_), .B0(new_n11315_), .Y(new_n13421_));
  OAI21  g12419(.A0(new_n13420_), .A1(new_n11316_), .B0(new_n13421_), .Y(new_n13422_));
  NAND3  g12420(.A(new_n11296_), .B(new_n11305_), .C(new_n11304_), .Y(new_n13423_));
  AOI21  g12421(.A0(new_n11305_), .A1(new_n11304_), .B0(new_n11296_), .Y(new_n13424_));
  AOI21  g12422(.A0(new_n13423_), .A1(new_n11300_), .B0(new_n13424_), .Y(new_n13425_));
  XOR2   g12423(.A(new_n13425_), .B(new_n13422_), .Y(new_n13426_));
  NAND2  g12424(.A(new_n13417_), .B(new_n11288_), .Y(new_n13427_));
  AOI21  g12425(.A0(new_n13425_), .A1(new_n13422_), .B0(new_n13418_), .Y(new_n13428_));
  OAI211 g12426(.A0(new_n13425_), .A1(new_n13422_), .B0(new_n13428_), .B1(new_n13427_), .Y(new_n13429_));
  OAI21  g12427(.A0(new_n13426_), .A1(new_n13419_), .B0(new_n13429_), .Y(new_n13430_));
  XOR2   g12428(.A(new_n13430_), .B(new_n13414_), .Y(new_n13431_));
  XOR2   g12429(.A(new_n13431_), .B(new_n13396_), .Y(new_n13432_));
  AOI21  g12430(.A0(new_n5398_), .A1(new_n5334_), .B0(new_n5434_), .Y(new_n13433_));
  AOI21  g12431(.A0(new_n11279_), .A1(new_n11278_), .B0(new_n13433_), .Y(new_n13434_));
  NOR4   g12432(.A(new_n11275_), .B(new_n11271_), .C(new_n11268_), .D(new_n5434_), .Y(new_n13435_));
  NOR2   g12433(.A(new_n13435_), .B(new_n13434_), .Y(new_n13436_));
  XOR2   g12434(.A(new_n13436_), .B(new_n11267_), .Y(new_n13437_));
  XOR2   g12435(.A(new_n13437_), .B(new_n11251_), .Y(new_n13438_));
  OAI22  g12436(.A0(new_n13438_), .A1(new_n11249_), .B0(new_n11223_), .B1(new_n6077_), .Y(new_n13439_));
  NAND2  g12437(.A(new_n13437_), .B(new_n11251_), .Y(new_n13440_));
  NOR3   g12438(.A(new_n5420_), .B(new_n5402_), .C(new_n5392_), .Y(new_n13441_));
  OAI21  g12439(.A0(new_n13441_), .A1(new_n5298_), .B0(new_n5437_), .Y(new_n13442_));
  AOI211 g12440(.A0(new_n11282_), .A1(new_n13442_), .B(new_n11248_), .C(new_n11244_), .Y(new_n13443_));
  NAND2  g12441(.A(new_n13443_), .B(new_n13440_), .Y(new_n13444_));
  NAND2  g12442(.A(new_n13444_), .B(new_n13439_), .Y(new_n13445_));
  AOI211 g12443(.A0(new_n5562_), .A1(new_n5519_), .B(new_n11240_), .C(new_n11239_), .Y(new_n13446_));
  AOI21  g12444(.A0(new_n13446_), .A1(new_n11225_), .B0(new_n11242_), .Y(new_n13447_));
  AOI22  g12445(.A0(new_n11235_), .A1(new_n11230_), .B0(new_n11225_), .B1(new_n5563_), .Y(new_n13448_));
  AOI21  g12446(.A0(new_n11232_), .A1(new_n11231_), .B0(new_n11229_), .Y(new_n13449_));
  OAI21  g12447(.A0(new_n13448_), .A1(new_n13447_), .B0(new_n13449_), .Y(new_n13450_));
  OAI211 g12448(.A0(new_n5550_), .A1(new_n5556_), .B0(new_n11235_), .B1(new_n11230_), .Y(new_n13451_));
  OAI21  g12449(.A0(new_n13451_), .A1(new_n11245_), .B0(new_n11237_), .Y(new_n13452_));
  OAI22  g12450(.A0(new_n11240_), .A1(new_n11239_), .B0(new_n11245_), .B1(new_n5557_), .Y(new_n13453_));
  INV    g12451(.A(new_n13449_), .Y(new_n13454_));
  NAND3  g12452(.A(new_n13454_), .B(new_n13453_), .C(new_n13452_), .Y(new_n13455_));
  NAND2  g12453(.A(new_n13455_), .B(new_n13450_), .Y(new_n13456_));
  NOR2   g12454(.A(new_n5428_), .B(new_n5426_), .Y(new_n13457_));
  OAI22  g12455(.A0(new_n5436_), .A1(new_n5392_), .B0(new_n5297_), .B1(new_n13457_), .Y(new_n13458_));
  AOI22  g12456(.A0(new_n11281_), .A1(new_n11267_), .B0(new_n13458_), .B1(new_n5437_), .Y(new_n13459_));
  AOI22  g12457(.A0(new_n11265_), .A1(new_n11264_), .B0(new_n11263_), .B1(new_n5296_), .Y(new_n13460_));
  NOR4   g12458(.A(new_n11261_), .B(new_n11258_), .C(new_n11255_), .D(new_n11254_), .Y(new_n13461_));
  NOR4   g12459(.A(new_n13435_), .B(new_n13434_), .C(new_n13461_), .D(new_n13460_), .Y(new_n13462_));
  AOI211 g12460(.A0(new_n5398_), .A1(new_n5334_), .B(new_n11269_), .C(new_n5434_), .Y(new_n13463_));
  OAI22  g12461(.A0(new_n13463_), .A1(new_n11270_), .B0(new_n11273_), .B1(new_n13433_), .Y(new_n13464_));
  NOR3   g12462(.A(new_n11256_), .B(new_n11255_), .C(new_n11254_), .Y(new_n13465_));
  OAI21  g12463(.A0(new_n11255_), .A1(new_n11254_), .B0(new_n11256_), .Y(new_n13466_));
  OAI21  g12464(.A0(new_n13465_), .A1(new_n11257_), .B0(new_n13466_), .Y(new_n13467_));
  XOR2   g12465(.A(new_n13467_), .B(new_n13464_), .Y(new_n13468_));
  OAI21  g12466(.A0(new_n13462_), .A1(new_n13459_), .B0(new_n13468_), .Y(new_n13469_));
  OAI22  g12467(.A0(new_n13435_), .A1(new_n13434_), .B0(new_n13461_), .B1(new_n13460_), .Y(new_n13470_));
  NAND2  g12468(.A(new_n13470_), .B(new_n13442_), .Y(new_n13471_));
  NAND3  g12469(.A(new_n11259_), .B(new_n11263_), .C(new_n5296_), .Y(new_n13472_));
  AOI21  g12470(.A0(new_n11263_), .A1(new_n5296_), .B0(new_n11259_), .Y(new_n13473_));
  AOI21  g12471(.A0(new_n13472_), .A1(new_n11260_), .B0(new_n13473_), .Y(new_n13474_));
  AOI21  g12472(.A0(new_n13474_), .A1(new_n13464_), .B0(new_n13462_), .Y(new_n13475_));
  OAI211 g12473(.A0(new_n13474_), .A1(new_n13464_), .B0(new_n13475_), .B1(new_n13471_), .Y(new_n13476_));
  NAND2  g12474(.A(new_n13476_), .B(new_n13469_), .Y(new_n13477_));
  XOR2   g12475(.A(new_n13477_), .B(new_n13456_), .Y(new_n13478_));
  XOR2   g12476(.A(new_n13478_), .B(new_n13445_), .Y(new_n13479_));
  XOR2   g12477(.A(new_n13479_), .B(new_n13432_), .Y(new_n13480_));
  NOR2   g12478(.A(new_n13480_), .B(new_n13391_), .Y(new_n13481_));
  XOR2   g12479(.A(new_n13480_), .B(new_n13391_), .Y(new_n13482_));
  OAI22  g12480(.A0(new_n11399_), .A1(new_n11398_), .B0(new_n11397_), .B1(new_n11396_), .Y(new_n13483_));
  NAND4  g12481(.A(new_n11394_), .B(new_n11391_), .C(new_n11388_), .D(new_n5176_), .Y(new_n13484_));
  NAND2  g12482(.A(new_n13484_), .B(new_n13483_), .Y(new_n13485_));
  XOR2   g12483(.A(new_n13485_), .B(new_n11387_), .Y(new_n13486_));
  XOR2   g12484(.A(new_n13486_), .B(new_n11369_), .Y(new_n13487_));
  OAI21  g12485(.A0(new_n5060_), .A1(new_n5065_), .B0(new_n5067_), .Y(new_n13488_));
  XOR2   g12486(.A(new_n11433_), .B(new_n13488_), .Y(new_n13489_));
  NOR2   g12487(.A(new_n13489_), .B(new_n13487_), .Y(new_n13490_));
  NAND2  g12488(.A(new_n13489_), .B(new_n13487_), .Y(new_n13491_));
  OAI21  g12489(.A0(new_n13490_), .A1(new_n11600_), .B0(new_n13491_), .Y(new_n13492_));
  AOI21  g12490(.A0(new_n11432_), .A1(new_n11417_), .B0(new_n11404_), .Y(new_n13493_));
  NOR2   g12491(.A(new_n11420_), .B(new_n11419_), .Y(new_n13494_));
  AOI21  g12492(.A0(new_n11430_), .A1(new_n11428_), .B0(new_n13494_), .Y(new_n13495_));
  NAND3  g12493(.A(new_n11431_), .B(new_n11416_), .C(new_n11412_), .Y(new_n13496_));
  NOR2   g12494(.A(new_n13496_), .B(new_n13495_), .Y(new_n13497_));
  NOR3   g12495(.A(new_n11421_), .B(new_n11420_), .C(new_n11419_), .Y(new_n13498_));
  OAI22  g12496(.A0(new_n13498_), .A1(new_n11429_), .B0(new_n11423_), .B1(new_n13494_), .Y(new_n13499_));
  AOI21  g12497(.A0(new_n4838_), .A1(new_n4835_), .B0(new_n4852_), .Y(new_n13500_));
  NOR3   g12498(.A(new_n13500_), .B(new_n11405_), .C(new_n4856_), .Y(new_n13501_));
  OAI21  g12499(.A0(new_n11405_), .A1(new_n4856_), .B0(new_n13500_), .Y(new_n13502_));
  OAI21  g12500(.A0(new_n13501_), .A1(new_n11410_), .B0(new_n13502_), .Y(new_n13503_));
  XOR2   g12501(.A(new_n13503_), .B(new_n13499_), .Y(new_n13504_));
  OAI21  g12502(.A0(new_n13497_), .A1(new_n13493_), .B0(new_n13504_), .Y(new_n13505_));
  NAND4  g12503(.A(new_n11431_), .B(new_n11426_), .C(new_n11416_), .D(new_n11412_), .Y(new_n13506_));
  NOR3   g12504(.A(new_n4839_), .B(new_n4836_), .C(new_n4841_), .Y(new_n13507_));
  OAI211 g12505(.A0(new_n4853_), .A1(new_n4852_), .B0(new_n13507_), .B1(new_n4845_), .Y(new_n13508_));
  NAND3  g12506(.A(new_n11406_), .B(new_n11413_), .C(new_n13508_), .Y(new_n13509_));
  AOI21  g12507(.A0(new_n11413_), .A1(new_n13508_), .B0(new_n11406_), .Y(new_n13510_));
  AOI21  g12508(.A0(new_n13509_), .A1(new_n11414_), .B0(new_n13510_), .Y(new_n13511_));
  NAND2  g12509(.A(new_n13511_), .B(new_n13499_), .Y(new_n13512_));
  NAND3  g12510(.A(new_n11423_), .B(new_n11427_), .C(new_n4947_), .Y(new_n13513_));
  AOI21  g12511(.A0(new_n11427_), .A1(new_n4947_), .B0(new_n11423_), .Y(new_n13514_));
  AOI21  g12512(.A0(new_n13513_), .A1(new_n11424_), .B0(new_n13514_), .Y(new_n13515_));
  NAND2  g12513(.A(new_n13503_), .B(new_n13515_), .Y(new_n13516_));
  NAND3  g12514(.A(new_n13516_), .B(new_n13512_), .C(new_n13506_), .Y(new_n13517_));
  OAI21  g12515(.A0(new_n13517_), .A1(new_n13493_), .B0(new_n13505_), .Y(new_n13518_));
  AOI22  g12516(.A0(new_n11385_), .A1(new_n11383_), .B0(new_n11382_), .B1(new_n5119_), .Y(new_n13519_));
  NOR4   g12517(.A(new_n11380_), .B(new_n11377_), .C(new_n11374_), .D(new_n11372_), .Y(new_n13520_));
  OAI22  g12518(.A0(new_n11400_), .A1(new_n11395_), .B0(new_n13520_), .B1(new_n13519_), .Y(new_n13521_));
  NOR4   g12519(.A(new_n11400_), .B(new_n11395_), .C(new_n13520_), .D(new_n13519_), .Y(new_n13522_));
  AOI21  g12520(.A0(new_n13521_), .A1(new_n11369_), .B0(new_n13522_), .Y(new_n13523_));
  NAND3  g12521(.A(new_n11389_), .B(new_n11388_), .C(new_n5176_), .Y(new_n13524_));
  AOI21  g12522(.A0(new_n11388_), .A1(new_n5176_), .B0(new_n11389_), .Y(new_n13525_));
  AOI21  g12523(.A0(new_n13524_), .A1(new_n11390_), .B0(new_n13525_), .Y(new_n13526_));
  NOR3   g12524(.A(new_n11376_), .B(new_n11374_), .C(new_n11372_), .Y(new_n13527_));
  OAI21  g12525(.A0(new_n11374_), .A1(new_n11372_), .B0(new_n11376_), .Y(new_n13528_));
  OAI21  g12526(.A0(new_n13527_), .A1(new_n11384_), .B0(new_n13528_), .Y(new_n13529_));
  XOR2   g12527(.A(new_n13529_), .B(new_n13526_), .Y(new_n13530_));
  NOR2   g12528(.A(new_n13530_), .B(new_n13523_), .Y(new_n13531_));
  NAND4  g12529(.A(new_n13484_), .B(new_n13483_), .C(new_n11386_), .D(new_n11381_), .Y(new_n13532_));
  OAI21  g12530(.A0(new_n13529_), .A1(new_n13526_), .B0(new_n13532_), .Y(new_n13533_));
  AOI221 g12531(.A0(new_n13529_), .A1(new_n13526_), .C0(new_n13533_), .B0(new_n13521_), .B1(new_n11369_), .Y(new_n13534_));
  NOR2   g12532(.A(new_n13534_), .B(new_n13531_), .Y(new_n13535_));
  XOR2   g12533(.A(new_n13535_), .B(new_n13518_), .Y(new_n13536_));
  XOR2   g12534(.A(new_n13536_), .B(new_n13492_), .Y(new_n13537_));
  OAI21  g12535(.A0(new_n6076_), .A1(new_n5565_), .B0(new_n5568_), .Y(new_n13538_));
  XOR2   g12536(.A(new_n11284_), .B(new_n13538_), .Y(new_n13539_));
  NAND2  g12537(.A(new_n11439_), .B(new_n13539_), .Y(new_n13540_));
  NOR2   g12538(.A(new_n11439_), .B(new_n13539_), .Y(new_n13541_));
  AOI21  g12539(.A0(new_n13540_), .A1(new_n11222_), .B0(new_n13541_), .Y(new_n13542_));
  NOR2   g12540(.A(new_n13401_), .B(new_n13400_), .Y(new_n13543_));
  XOR2   g12541(.A(new_n13543_), .B(new_n11344_), .Y(new_n13544_));
  XOR2   g12542(.A(new_n13544_), .B(new_n11329_), .Y(new_n13545_));
  NAND2  g12543(.A(new_n13545_), .B(new_n11327_), .Y(new_n13546_));
  NOR2   g12544(.A(new_n13545_), .B(new_n11327_), .Y(new_n13547_));
  AOI21  g12545(.A0(new_n13546_), .A1(new_n11438_), .B0(new_n13547_), .Y(new_n13548_));
  XOR2   g12546(.A(new_n13431_), .B(new_n13548_), .Y(new_n13549_));
  XOR2   g12547(.A(new_n13479_), .B(new_n13549_), .Y(new_n13550_));
  OAI21  g12548(.A0(new_n13550_), .A1(new_n13542_), .B0(new_n13537_), .Y(new_n13551_));
  OAI221 g12549(.A0(new_n13551_), .A1(new_n13481_), .C0(new_n13388_), .B0(new_n13537_), .B1(new_n13482_), .Y(new_n13552_));
  OAI22  g12550(.A0(new_n13551_), .A1(new_n13481_), .B0(new_n13537_), .B1(new_n13482_), .Y(new_n13553_));
  XOR2   g12551(.A(new_n13553_), .B(new_n13388_), .Y(new_n13554_));
  NOR2   g12552(.A(new_n11595_), .B(new_n11523_), .Y(new_n13555_));
  NAND2  g12553(.A(new_n11595_), .B(new_n11523_), .Y(new_n13556_));
  OAI21  g12554(.A0(new_n13555_), .A1(new_n11445_), .B0(new_n13556_), .Y(new_n13557_));
  AOI21  g12555(.A0(new_n6740_), .A1(new_n6731_), .B0(new_n6733_), .Y(new_n13558_));
  AOI21  g12556(.A0(new_n6577_), .A1(new_n6568_), .B0(new_n6729_), .Y(new_n13559_));
  XOR2   g12557(.A(new_n11559_), .B(new_n13559_), .Y(new_n13560_));
  AOI21  g12558(.A0(new_n6714_), .A1(new_n6633_), .B0(new_n6724_), .Y(new_n13561_));
  XOR2   g12559(.A(new_n11592_), .B(new_n13561_), .Y(new_n13562_));
  NOR2   g12560(.A(new_n13562_), .B(new_n13560_), .Y(new_n13563_));
  NAND2  g12561(.A(new_n13562_), .B(new_n13560_), .Y(new_n13564_));
  OAI21  g12562(.A0(new_n13563_), .A1(new_n13558_), .B0(new_n13564_), .Y(new_n13565_));
  OAI21  g12563(.A0(new_n6712_), .A1(new_n6707_), .B0(new_n6714_), .Y(new_n13566_));
  NAND2  g12564(.A(new_n11579_), .B(new_n11578_), .Y(new_n13567_));
  OAI21  g12565(.A0(new_n11589_), .A1(new_n11588_), .B0(new_n13567_), .Y(new_n13568_));
  NAND4  g12566(.A(new_n11585_), .B(new_n11582_), .C(new_n11579_), .D(new_n11578_), .Y(new_n13569_));
  AOI22  g12567(.A0(new_n13569_), .A1(new_n13568_), .B0(new_n11575_), .B1(new_n11570_), .Y(new_n13570_));
  AOI21  g12568(.A0(new_n13566_), .A1(new_n6715_), .B0(new_n13570_), .Y(new_n13571_));
  NOR2   g12569(.A(new_n11564_), .B(new_n11563_), .Y(new_n13572_));
  AOI21  g12570(.A0(new_n11574_), .A1(new_n11572_), .B0(new_n13572_), .Y(new_n13573_));
  NOR4   g12571(.A(new_n11569_), .B(new_n11566_), .C(new_n11564_), .D(new_n11563_), .Y(new_n13574_));
  NOR4   g12572(.A(new_n11590_), .B(new_n11586_), .C(new_n13574_), .D(new_n13573_), .Y(new_n13575_));
  NAND3  g12573(.A(new_n11580_), .B(new_n11579_), .C(new_n11578_), .Y(new_n13576_));
  AOI22  g12574(.A0(new_n13576_), .A1(new_n11581_), .B0(new_n11583_), .B1(new_n13567_), .Y(new_n13577_));
  NOR3   g12575(.A(new_n11565_), .B(new_n11564_), .C(new_n11563_), .Y(new_n13578_));
  OAI22  g12576(.A0(new_n13578_), .A1(new_n11573_), .B0(new_n11567_), .B1(new_n13572_), .Y(new_n13579_));
  NOR2   g12577(.A(new_n13579_), .B(new_n13577_), .Y(new_n13580_));
  NAND2  g12578(.A(new_n13576_), .B(new_n11581_), .Y(new_n13581_));
  NAND2  g12579(.A(new_n11583_), .B(new_n13567_), .Y(new_n13582_));
  NAND2  g12580(.A(new_n13582_), .B(new_n13581_), .Y(new_n13583_));
  NOR2   g12581(.A(new_n13578_), .B(new_n11573_), .Y(new_n13584_));
  NOR2   g12582(.A(new_n11567_), .B(new_n13572_), .Y(new_n13585_));
  NOR2   g12583(.A(new_n13585_), .B(new_n13584_), .Y(new_n13586_));
  NOR2   g12584(.A(new_n13586_), .B(new_n13583_), .Y(new_n13587_));
  OAI22  g12585(.A0(new_n13587_), .A1(new_n13580_), .B0(new_n13575_), .B1(new_n13571_), .Y(new_n13588_));
  NAND2  g12586(.A(new_n13579_), .B(new_n13577_), .Y(new_n13589_));
  NOR2   g12587(.A(new_n13580_), .B(new_n13575_), .Y(new_n13590_));
  OAI211 g12588(.A0(new_n13570_), .A1(new_n13561_), .B0(new_n13590_), .B1(new_n13589_), .Y(new_n13591_));
  NAND2  g12589(.A(new_n13591_), .B(new_n13588_), .Y(new_n13592_));
  OAI21  g12590(.A0(new_n6575_), .A1(new_n6570_), .B0(new_n6577_), .Y(new_n13593_));
  OAI22  g12591(.A0(new_n11556_), .A1(new_n11555_), .B0(new_n11554_), .B1(new_n11552_), .Y(new_n13594_));
  NAND4  g12592(.A(new_n11550_), .B(new_n11547_), .C(new_n11544_), .D(new_n11543_), .Y(new_n13595_));
  NAND2  g12593(.A(new_n13595_), .B(new_n13594_), .Y(new_n13596_));
  AOI22  g12594(.A0(new_n13596_), .A1(new_n11541_), .B0(new_n13593_), .B1(new_n6579_), .Y(new_n13597_));
  NOR2   g12595(.A(new_n11529_), .B(new_n11528_), .Y(new_n13598_));
  AOI21  g12596(.A0(new_n11539_), .A1(new_n11537_), .B0(new_n13598_), .Y(new_n13599_));
  NOR4   g12597(.A(new_n11534_), .B(new_n11531_), .C(new_n11529_), .D(new_n11528_), .Y(new_n13600_));
  NOR4   g12598(.A(new_n11557_), .B(new_n11551_), .C(new_n13600_), .D(new_n13599_), .Y(new_n13601_));
  NAND3  g12599(.A(new_n11545_), .B(new_n11544_), .C(new_n11543_), .Y(new_n13602_));
  AOI21  g12600(.A0(new_n11544_), .A1(new_n11543_), .B0(new_n11545_), .Y(new_n13603_));
  AOI21  g12601(.A0(new_n13602_), .A1(new_n11546_), .B0(new_n13603_), .Y(new_n13604_));
  NOR3   g12602(.A(new_n11530_), .B(new_n11529_), .C(new_n11528_), .Y(new_n13605_));
  OAI22  g12603(.A0(new_n13605_), .A1(new_n11538_), .B0(new_n11532_), .B1(new_n13598_), .Y(new_n13606_));
  NOR2   g12604(.A(new_n13606_), .B(new_n13604_), .Y(new_n13607_));
  NOR3   g12605(.A(new_n11548_), .B(new_n11554_), .C(new_n11552_), .Y(new_n13608_));
  OAI21  g12606(.A0(new_n11554_), .A1(new_n11552_), .B0(new_n11548_), .Y(new_n13609_));
  OAI21  g12607(.A0(new_n13608_), .A1(new_n11549_), .B0(new_n13609_), .Y(new_n13610_));
  NAND2  g12608(.A(new_n11532_), .B(new_n6565_), .Y(new_n13611_));
  OAI21  g12609(.A0(new_n13611_), .A1(new_n11529_), .B0(new_n11533_), .Y(new_n13612_));
  OAI21  g12610(.A0(new_n11529_), .A1(new_n11528_), .B0(new_n11530_), .Y(new_n13613_));
  AOI21  g12611(.A0(new_n13613_), .A1(new_n13612_), .B0(new_n13610_), .Y(new_n13614_));
  OAI22  g12612(.A0(new_n13614_), .A1(new_n13607_), .B0(new_n13601_), .B1(new_n13597_), .Y(new_n13615_));
  OAI21  g12613(.A0(new_n13600_), .A1(new_n13599_), .B0(new_n13596_), .Y(new_n13616_));
  NAND2  g12614(.A(new_n13616_), .B(new_n11526_), .Y(new_n13617_));
  NOR3   g12615(.A(new_n13614_), .B(new_n13607_), .C(new_n13601_), .Y(new_n13618_));
  NAND2  g12616(.A(new_n13618_), .B(new_n13617_), .Y(new_n13619_));
  NAND2  g12617(.A(new_n13619_), .B(new_n13615_), .Y(new_n13620_));
  XOR2   g12618(.A(new_n13620_), .B(new_n13592_), .Y(new_n13621_));
  XOR2   g12619(.A(new_n13621_), .B(new_n13565_), .Y(new_n13622_));
  AOI21  g12620(.A0(new_n7034_), .A1(new_n7030_), .B0(new_n7048_), .Y(new_n13623_));
  OAI22  g12621(.A0(new_n11482_), .A1(new_n11481_), .B0(new_n11480_), .B1(new_n11479_), .Y(new_n13624_));
  NAND4  g12622(.A(new_n11477_), .B(new_n11474_), .C(new_n11471_), .D(new_n6954_), .Y(new_n13625_));
  NAND2  g12623(.A(new_n13625_), .B(new_n13624_), .Y(new_n13626_));
  XOR2   g12624(.A(new_n13626_), .B(new_n11470_), .Y(new_n13627_));
  XOR2   g12625(.A(new_n13627_), .B(new_n11450_), .Y(new_n13628_));
  OAI22  g12626(.A0(new_n11517_), .A1(new_n11516_), .B0(new_n11515_), .B1(new_n11514_), .Y(new_n13629_));
  NAND4  g12627(.A(new_n11512_), .B(new_n11509_), .C(new_n11506_), .D(new_n6874_), .Y(new_n13630_));
  NAND2  g12628(.A(new_n13630_), .B(new_n13629_), .Y(new_n13631_));
  XOR2   g12629(.A(new_n13631_), .B(new_n11505_), .Y(new_n13632_));
  XOR2   g12630(.A(new_n13632_), .B(new_n11487_), .Y(new_n13633_));
  NOR2   g12631(.A(new_n13633_), .B(new_n13628_), .Y(new_n13634_));
  NAND2  g12632(.A(new_n13633_), .B(new_n13628_), .Y(new_n13635_));
  OAI21  g12633(.A0(new_n13634_), .A1(new_n13623_), .B0(new_n13635_), .Y(new_n13636_));
  AOI22  g12634(.A0(new_n11503_), .A1(new_n11502_), .B0(new_n11501_), .B1(new_n6800_), .Y(new_n13637_));
  NOR4   g12635(.A(new_n11499_), .B(new_n11493_), .C(new_n11490_), .D(new_n11489_), .Y(new_n13638_));
  OAI22  g12636(.A0(new_n11518_), .A1(new_n11513_), .B0(new_n13638_), .B1(new_n13637_), .Y(new_n13639_));
  NOR4   g12637(.A(new_n11518_), .B(new_n11513_), .C(new_n13638_), .D(new_n13637_), .Y(new_n13640_));
  AOI21  g12638(.A0(new_n13639_), .A1(new_n11487_), .B0(new_n13640_), .Y(new_n13641_));
  NOR3   g12639(.A(new_n11510_), .B(new_n11515_), .C(new_n11514_), .Y(new_n13642_));
  OAI21  g12640(.A0(new_n11515_), .A1(new_n11514_), .B0(new_n11510_), .Y(new_n13643_));
  OAI21  g12641(.A0(new_n13642_), .A1(new_n11511_), .B0(new_n13643_), .Y(new_n13644_));
  NAND3  g12642(.A(new_n11494_), .B(new_n11501_), .C(new_n6800_), .Y(new_n13645_));
  AOI21  g12643(.A0(new_n11501_), .A1(new_n6800_), .B0(new_n11494_), .Y(new_n13646_));
  AOI21  g12644(.A0(new_n13645_), .A1(new_n11498_), .B0(new_n13646_), .Y(new_n13647_));
  XOR2   g12645(.A(new_n13647_), .B(new_n13644_), .Y(new_n13648_));
  NAND2  g12646(.A(new_n13639_), .B(new_n11487_), .Y(new_n13649_));
  NOR2   g12647(.A(new_n13647_), .B(new_n13644_), .Y(new_n13650_));
  NAND4  g12648(.A(new_n13630_), .B(new_n13629_), .C(new_n11504_), .D(new_n11500_), .Y(new_n13651_));
  NAND3  g12649(.A(new_n11507_), .B(new_n11506_), .C(new_n6874_), .Y(new_n13652_));
  AOI21  g12650(.A0(new_n11506_), .A1(new_n6874_), .B0(new_n11507_), .Y(new_n13653_));
  AOI21  g12651(.A0(new_n13652_), .A1(new_n11508_), .B0(new_n13653_), .Y(new_n13654_));
  NOR3   g12652(.A(new_n11491_), .B(new_n11490_), .C(new_n11489_), .Y(new_n13655_));
  OAI21  g12653(.A0(new_n11490_), .A1(new_n11489_), .B0(new_n11491_), .Y(new_n13656_));
  OAI21  g12654(.A0(new_n13655_), .A1(new_n11492_), .B0(new_n13656_), .Y(new_n13657_));
  OAI21  g12655(.A0(new_n13657_), .A1(new_n13654_), .B0(new_n13651_), .Y(new_n13658_));
  NOR2   g12656(.A(new_n13658_), .B(new_n13650_), .Y(new_n13659_));
  NAND2  g12657(.A(new_n13659_), .B(new_n13649_), .Y(new_n13660_));
  OAI21  g12658(.A0(new_n13648_), .A1(new_n13641_), .B0(new_n13660_), .Y(new_n13661_));
  AOI22  g12659(.A0(new_n11468_), .A1(new_n11467_), .B0(new_n11466_), .B1(new_n7022_), .Y(new_n13662_));
  NOR4   g12660(.A(new_n11464_), .B(new_n11458_), .C(new_n11455_), .D(new_n11453_), .Y(new_n13663_));
  OAI22  g12661(.A0(new_n11483_), .A1(new_n11478_), .B0(new_n13663_), .B1(new_n13662_), .Y(new_n13664_));
  NOR4   g12662(.A(new_n11483_), .B(new_n11478_), .C(new_n13663_), .D(new_n13662_), .Y(new_n13665_));
  AOI21  g12663(.A0(new_n13664_), .A1(new_n11450_), .B0(new_n13665_), .Y(new_n13666_));
  NOR3   g12664(.A(new_n11475_), .B(new_n11480_), .C(new_n11479_), .Y(new_n13667_));
  OAI21  g12665(.A0(new_n11480_), .A1(new_n11479_), .B0(new_n11475_), .Y(new_n13668_));
  OAI21  g12666(.A0(new_n13667_), .A1(new_n11476_), .B0(new_n13668_), .Y(new_n13669_));
  NAND3  g12667(.A(new_n11459_), .B(new_n11466_), .C(new_n7022_), .Y(new_n13670_));
  AOI21  g12668(.A0(new_n11466_), .A1(new_n7022_), .B0(new_n11459_), .Y(new_n13671_));
  AOI21  g12669(.A0(new_n13670_), .A1(new_n11463_), .B0(new_n13671_), .Y(new_n13672_));
  XOR2   g12670(.A(new_n13672_), .B(new_n13669_), .Y(new_n13673_));
  NAND2  g12671(.A(new_n13664_), .B(new_n11450_), .Y(new_n13674_));
  NOR2   g12672(.A(new_n13672_), .B(new_n13669_), .Y(new_n13675_));
  NAND4  g12673(.A(new_n13625_), .B(new_n13624_), .C(new_n11469_), .D(new_n11465_), .Y(new_n13676_));
  NAND3  g12674(.A(new_n11472_), .B(new_n11471_), .C(new_n6954_), .Y(new_n13677_));
  AOI21  g12675(.A0(new_n11471_), .A1(new_n6954_), .B0(new_n11472_), .Y(new_n13678_));
  AOI21  g12676(.A0(new_n13677_), .A1(new_n11473_), .B0(new_n13678_), .Y(new_n13679_));
  NOR3   g12677(.A(new_n11456_), .B(new_n11455_), .C(new_n11453_), .Y(new_n13680_));
  OAI21  g12678(.A0(new_n11455_), .A1(new_n11453_), .B0(new_n11456_), .Y(new_n13681_));
  OAI21  g12679(.A0(new_n13680_), .A1(new_n11457_), .B0(new_n13681_), .Y(new_n13682_));
  OAI21  g12680(.A0(new_n13682_), .A1(new_n13679_), .B0(new_n13676_), .Y(new_n13683_));
  NOR2   g12681(.A(new_n13683_), .B(new_n13675_), .Y(new_n13684_));
  NAND2  g12682(.A(new_n13684_), .B(new_n13674_), .Y(new_n13685_));
  OAI21  g12683(.A0(new_n13673_), .A1(new_n13666_), .B0(new_n13685_), .Y(new_n13686_));
  XOR2   g12684(.A(new_n13686_), .B(new_n13661_), .Y(new_n13687_));
  XOR2   g12685(.A(new_n13687_), .B(new_n13636_), .Y(new_n13688_));
  XOR2   g12686(.A(new_n13688_), .B(new_n13622_), .Y(new_n13689_));
  XOR2   g12687(.A(new_n13689_), .B(new_n13557_), .Y(new_n13690_));
  NOR2   g12688(.A(new_n11603_), .B(new_n11436_), .Y(new_n13691_));
  OAI22  g12689(.A0(new_n13386_), .A1(new_n11599_), .B0(new_n13691_), .B1(new_n11221_), .Y(new_n13692_));
  AOI21  g12690(.A0(new_n13553_), .A1(new_n13692_), .B0(new_n13690_), .Y(new_n13693_));
  AOI22  g12691(.A0(new_n13693_), .A1(new_n13552_), .B0(new_n13690_), .B1(new_n13554_), .Y(new_n13694_));
  XOR2   g12692(.A(new_n13694_), .B(new_n13384_), .Y(new_n13695_));
  XOR2   g12693(.A(new_n13695_), .B(new_n13377_), .Y(new_n13696_));
  NOR2   g12694(.A(new_n13696_), .B(new_n12895_), .Y(new_n13697_));
  AOI21  g12695(.A0(new_n11202_), .A1(new_n7054_), .B0(new_n7056_), .Y(new_n13698_));
  XOR2   g12696(.A(new_n11607_), .B(new_n13698_), .Y(new_n13699_));
  NAND2  g12697(.A(new_n12229_), .B(new_n13699_), .Y(new_n13700_));
  NOR2   g12698(.A(new_n12229_), .B(new_n13699_), .Y(new_n13701_));
  AOI21  g12699(.A0(new_n13700_), .A1(new_n11219_), .B0(new_n13701_), .Y(new_n13702_));
  XOR2   g12700(.A(new_n11917_), .B(new_n13132_), .Y(new_n13703_));
  NOR2   g12701(.A(new_n12227_), .B(new_n13703_), .Y(new_n13704_));
  NAND2  g12702(.A(new_n12227_), .B(new_n13703_), .Y(new_n13705_));
  OAI21  g12703(.A0(new_n13704_), .A1(new_n12881_), .B0(new_n13705_), .Y(new_n13706_));
  XOR2   g12704(.A(new_n13376_), .B(new_n13706_), .Y(new_n13707_));
  XOR2   g12705(.A(new_n13695_), .B(new_n13707_), .Y(new_n13708_));
  XOR2   g12706(.A(new_n13708_), .B(new_n13702_), .Y(new_n13709_));
  AOI21  g12707(.A0(new_n4764_), .A1(new_n4755_), .B0(new_n12236_), .Y(new_n13710_));
  XOR2   g12708(.A(new_n12552_), .B(new_n13710_), .Y(new_n13711_));
  AOI21  g12709(.A0(new_n3552_), .A1(new_n2873_), .B0(new_n2875_), .Y(new_n13712_));
  XOR2   g12710(.A(new_n12876_), .B(new_n13712_), .Y(new_n13713_));
  NAND2  g12711(.A(new_n13713_), .B(new_n13711_), .Y(new_n13714_));
  NOR2   g12712(.A(new_n13713_), .B(new_n13711_), .Y(new_n13715_));
  AOI21  g12713(.A0(new_n13714_), .A1(new_n12888_), .B0(new_n13715_), .Y(new_n13716_));
  AOI21  g12714(.A0(new_n1926_), .A1(new_n1917_), .B0(new_n2871_), .Y(new_n13717_));
  XOR2   g12715(.A(new_n12713_), .B(new_n13717_), .Y(new_n13718_));
  AOI21  g12716(.A0(new_n2850_), .A1(new_n2372_), .B0(new_n2863_), .Y(new_n13719_));
  XOR2   g12717(.A(new_n12874_), .B(new_n13719_), .Y(new_n13720_));
  NAND2  g12718(.A(new_n13720_), .B(new_n13718_), .Y(new_n13721_));
  NOR2   g12719(.A(new_n13720_), .B(new_n13718_), .Y(new_n13722_));
  AOI21  g12720(.A0(new_n13721_), .A1(new_n12554_), .B0(new_n13722_), .Y(new_n13723_));
  NOR2   g12721(.A(new_n12873_), .B(new_n12796_), .Y(new_n13724_));
  NAND2  g12722(.A(new_n12873_), .B(new_n12796_), .Y(new_n13725_));
  OAI21  g12723(.A0(new_n13724_), .A1(new_n13719_), .B0(new_n13725_), .Y(new_n13726_));
  AOI21  g12724(.A0(new_n2586_), .A1(new_n2577_), .B0(new_n2821_), .Y(new_n13727_));
  XOR2   g12725(.A(new_n12831_), .B(new_n13727_), .Y(new_n13728_));
  OAI22  g12726(.A0(new_n12871_), .A1(new_n13728_), .B0(new_n12797_), .B1(new_n2825_), .Y(new_n13729_));
  NAND2  g12727(.A(new_n12871_), .B(new_n13728_), .Y(new_n13730_));
  NAND2  g12728(.A(new_n13730_), .B(new_n13729_), .Y(new_n13731_));
  AOI22  g12729(.A0(new_n12869_), .A1(new_n12854_), .B0(new_n12834_), .B1(new_n2805_), .Y(new_n13732_));
  AOI22  g12730(.A0(new_n12852_), .A1(new_n12851_), .B0(new_n12850_), .B1(new_n12849_), .Y(new_n13733_));
  NOR4   g12731(.A(new_n12846_), .B(new_n12840_), .C(new_n12836_), .D(new_n2675_), .Y(new_n13734_));
  AOI22  g12732(.A0(new_n12867_), .A1(new_n12866_), .B0(new_n12865_), .B1(new_n12864_), .Y(new_n13735_));
  NOR4   g12733(.A(new_n12861_), .B(new_n12858_), .C(new_n12855_), .D(new_n2766_), .Y(new_n13736_));
  NOR4   g12734(.A(new_n13736_), .B(new_n13735_), .C(new_n13734_), .D(new_n13733_), .Y(new_n13737_));
  NOR3   g12735(.A(new_n12856_), .B(new_n12855_), .C(new_n2766_), .Y(new_n13738_));
  OAI21  g12736(.A0(new_n12855_), .A1(new_n2766_), .B0(new_n12856_), .Y(new_n13739_));
  OAI21  g12737(.A0(new_n13738_), .A1(new_n12857_), .B0(new_n13739_), .Y(new_n13740_));
  NOR3   g12738(.A(new_n12837_), .B(new_n12836_), .C(new_n2675_), .Y(new_n13741_));
  OAI21  g12739(.A0(new_n12836_), .A1(new_n2675_), .B0(new_n12837_), .Y(new_n13742_));
  OAI21  g12740(.A0(new_n13741_), .A1(new_n12839_), .B0(new_n13742_), .Y(new_n13743_));
  XOR2   g12741(.A(new_n13743_), .B(new_n13740_), .Y(new_n13744_));
  OAI21  g12742(.A0(new_n13737_), .A1(new_n13732_), .B0(new_n13744_), .Y(new_n13745_));
  NAND3  g12743(.A(new_n12841_), .B(new_n12850_), .C(new_n12849_), .Y(new_n13746_));
  AOI21  g12744(.A0(new_n12850_), .A1(new_n12849_), .B0(new_n12841_), .Y(new_n13747_));
  AOI21  g12745(.A0(new_n13746_), .A1(new_n12845_), .B0(new_n13747_), .Y(new_n13748_));
  AOI21  g12746(.A0(new_n13748_), .A1(new_n13740_), .B0(new_n13737_), .Y(new_n13749_));
  OAI21  g12747(.A0(new_n13748_), .A1(new_n13740_), .B0(new_n13749_), .Y(new_n13750_));
  OAI21  g12748(.A0(new_n13750_), .A1(new_n13732_), .B0(new_n13745_), .Y(new_n13751_));
  NAND2  g12749(.A(new_n12818_), .B(new_n12817_), .Y(new_n13752_));
  OAI21  g12750(.A0(new_n12828_), .A1(new_n12826_), .B0(new_n13752_), .Y(new_n13753_));
  NAND4  g12751(.A(new_n12823_), .B(new_n12820_), .C(new_n12818_), .D(new_n12817_), .Y(new_n13754_));
  AOI22  g12752(.A0(new_n13754_), .A1(new_n13753_), .B0(new_n12814_), .B1(new_n12809_), .Y(new_n13755_));
  AOI21  g12753(.A0(new_n12799_), .A1(new_n2587_), .B0(new_n13755_), .Y(new_n13756_));
  NOR2   g12754(.A(new_n12803_), .B(new_n12802_), .Y(new_n13757_));
  AOI21  g12755(.A0(new_n12813_), .A1(new_n12811_), .B0(new_n13757_), .Y(new_n13758_));
  NOR4   g12756(.A(new_n12808_), .B(new_n12805_), .C(new_n12803_), .D(new_n12802_), .Y(new_n13759_));
  OAI22  g12757(.A0(new_n12829_), .A1(new_n12824_), .B0(new_n13759_), .B1(new_n13758_), .Y(new_n13760_));
  NOR4   g12758(.A(new_n12829_), .B(new_n12824_), .C(new_n13759_), .D(new_n13758_), .Y(new_n13761_));
  AOI21  g12759(.A0(new_n13760_), .A1(new_n12800_), .B0(new_n13761_), .Y(new_n13762_));
  NAND3  g12760(.A(new_n12819_), .B(new_n12818_), .C(new_n12817_), .Y(new_n13763_));
  AOI22  g12761(.A0(new_n13763_), .A1(new_n12827_), .B0(new_n12821_), .B1(new_n13752_), .Y(new_n13764_));
  NOR3   g12762(.A(new_n12804_), .B(new_n12803_), .C(new_n12802_), .Y(new_n13765_));
  OAI22  g12763(.A0(new_n13765_), .A1(new_n12812_), .B0(new_n12806_), .B1(new_n13757_), .Y(new_n13766_));
  XOR2   g12764(.A(new_n13766_), .B(new_n13764_), .Y(new_n13767_));
  NAND4  g12765(.A(new_n13754_), .B(new_n13753_), .C(new_n12814_), .D(new_n12809_), .Y(new_n13768_));
  NOR3   g12766(.A(new_n12821_), .B(new_n12825_), .C(new_n2467_), .Y(new_n13769_));
  OAI21  g12767(.A0(new_n12825_), .A1(new_n2467_), .B0(new_n12821_), .Y(new_n13770_));
  OAI21  g12768(.A0(new_n13769_), .A1(new_n12822_), .B0(new_n13770_), .Y(new_n13771_));
  OAI221 g12769(.A0(new_n13765_), .A1(new_n12812_), .C0(new_n13771_), .B0(new_n12806_), .B1(new_n13757_), .Y(new_n13772_));
  NAND2  g12770(.A(new_n13766_), .B(new_n13764_), .Y(new_n13773_));
  NAND3  g12771(.A(new_n13773_), .B(new_n13772_), .C(new_n13768_), .Y(new_n13774_));
  OAI22  g12772(.A0(new_n13774_), .A1(new_n13756_), .B0(new_n13767_), .B1(new_n13762_), .Y(new_n13775_));
  XOR2   g12773(.A(new_n13775_), .B(new_n13751_), .Y(new_n13776_));
  XOR2   g12774(.A(new_n13776_), .B(new_n13731_), .Y(new_n13777_));
  NAND2  g12775(.A(new_n12794_), .B(new_n12756_), .Y(new_n13778_));
  NOR2   g12776(.A(new_n12794_), .B(new_n12756_), .Y(new_n13779_));
  AOI21  g12777(.A0(new_n13778_), .A1(new_n12716_), .B0(new_n13779_), .Y(new_n13780_));
  AOI22  g12778(.A0(new_n12775_), .A1(new_n12774_), .B0(new_n12761_), .B1(new_n12760_), .Y(new_n13781_));
  AOI221 g12779(.A0(new_n2232_), .A1(new_n2228_), .C0(new_n12765_), .B0(new_n12767_), .B1(new_n2218_), .Y(new_n13782_));
  NOR4   g12780(.A(new_n12772_), .B(new_n12769_), .C(new_n13782_), .D(new_n2234_), .Y(new_n13783_));
  OAI22  g12781(.A0(new_n12790_), .A1(new_n12788_), .B0(new_n12787_), .B1(new_n2325_), .Y(new_n13784_));
  NAND4  g12782(.A(new_n12785_), .B(new_n12782_), .C(new_n12780_), .D(new_n12779_), .Y(new_n13785_));
  NAND2  g12783(.A(new_n13785_), .B(new_n13784_), .Y(new_n13786_));
  OAI21  g12784(.A0(new_n13783_), .A1(new_n13781_), .B0(new_n13786_), .Y(new_n13787_));
  NOR4   g12785(.A(new_n12791_), .B(new_n12786_), .C(new_n13783_), .D(new_n13781_), .Y(new_n13788_));
  AOI21  g12786(.A0(new_n13787_), .A1(new_n12758_), .B0(new_n13788_), .Y(new_n13789_));
  NOR3   g12787(.A(new_n12783_), .B(new_n12787_), .C(new_n2325_), .Y(new_n13790_));
  OAI21  g12788(.A0(new_n12787_), .A1(new_n2325_), .B0(new_n12783_), .Y(new_n13791_));
  OAI21  g12789(.A0(new_n13790_), .A1(new_n12784_), .B0(new_n13791_), .Y(new_n13792_));
  NAND3  g12790(.A(new_n12770_), .B(new_n12761_), .C(new_n12760_), .Y(new_n13793_));
  AOI22  g12791(.A0(new_n13793_), .A1(new_n12771_), .B0(new_n12763_), .B1(new_n12762_), .Y(new_n13794_));
  XOR2   g12792(.A(new_n13794_), .B(new_n13792_), .Y(new_n13795_));
  NAND2  g12793(.A(new_n13787_), .B(new_n12758_), .Y(new_n13796_));
  AOI21  g12794(.A0(new_n13794_), .A1(new_n13792_), .B0(new_n13788_), .Y(new_n13797_));
  OAI211 g12795(.A0(new_n13794_), .A1(new_n13792_), .B0(new_n13797_), .B1(new_n13796_), .Y(new_n13798_));
  OAI21  g12796(.A0(new_n13795_), .A1(new_n13789_), .B0(new_n13798_), .Y(new_n13799_));
  AOI22  g12797(.A0(new_n12738_), .A1(new_n12737_), .B0(new_n12736_), .B1(new_n2019_), .Y(new_n13800_));
  NOR4   g12798(.A(new_n12734_), .B(new_n12728_), .C(new_n12725_), .D(new_n12723_), .Y(new_n13801_));
  OAI22  g12799(.A0(new_n12753_), .A1(new_n12748_), .B0(new_n13801_), .B1(new_n13800_), .Y(new_n13802_));
  NOR4   g12800(.A(new_n12753_), .B(new_n12748_), .C(new_n13801_), .D(new_n13800_), .Y(new_n13803_));
  AOI21  g12801(.A0(new_n13802_), .A1(new_n12720_), .B0(new_n13803_), .Y(new_n13804_));
  NOR3   g12802(.A(new_n12745_), .B(new_n12750_), .C(new_n12749_), .Y(new_n13805_));
  OAI21  g12803(.A0(new_n12750_), .A1(new_n12749_), .B0(new_n12745_), .Y(new_n13806_));
  OAI21  g12804(.A0(new_n13805_), .A1(new_n12746_), .B0(new_n13806_), .Y(new_n13807_));
  NAND3  g12805(.A(new_n12729_), .B(new_n12736_), .C(new_n2019_), .Y(new_n13808_));
  AOI21  g12806(.A0(new_n12736_), .A1(new_n2019_), .B0(new_n12729_), .Y(new_n13809_));
  AOI21  g12807(.A0(new_n13808_), .A1(new_n12733_), .B0(new_n13809_), .Y(new_n13810_));
  XOR2   g12808(.A(new_n13810_), .B(new_n13807_), .Y(new_n13811_));
  NOR2   g12809(.A(new_n13811_), .B(new_n13804_), .Y(new_n13812_));
  NOR2   g12810(.A(new_n13810_), .B(new_n13807_), .Y(new_n13813_));
  OAI22  g12811(.A0(new_n12752_), .A1(new_n12751_), .B0(new_n12750_), .B1(new_n12749_), .Y(new_n13814_));
  NAND4  g12812(.A(new_n12747_), .B(new_n12744_), .C(new_n12741_), .D(new_n2119_), .Y(new_n13815_));
  NAND4  g12813(.A(new_n13815_), .B(new_n13814_), .C(new_n12739_), .D(new_n12735_), .Y(new_n13816_));
  NAND3  g12814(.A(new_n12742_), .B(new_n12741_), .C(new_n2119_), .Y(new_n13817_));
  AOI21  g12815(.A0(new_n12741_), .A1(new_n2119_), .B0(new_n12742_), .Y(new_n13818_));
  AOI21  g12816(.A0(new_n13817_), .A1(new_n12743_), .B0(new_n13818_), .Y(new_n13819_));
  NOR3   g12817(.A(new_n12726_), .B(new_n12725_), .C(new_n12723_), .Y(new_n13820_));
  OAI21  g12818(.A0(new_n12725_), .A1(new_n12723_), .B0(new_n12726_), .Y(new_n13821_));
  OAI21  g12819(.A0(new_n13820_), .A1(new_n12727_), .B0(new_n13821_), .Y(new_n13822_));
  OAI21  g12820(.A0(new_n13822_), .A1(new_n13819_), .B0(new_n13816_), .Y(new_n13823_));
  AOI211 g12821(.A0(new_n13802_), .A1(new_n12720_), .B(new_n13823_), .C(new_n13813_), .Y(new_n13824_));
  NOR2   g12822(.A(new_n13824_), .B(new_n13812_), .Y(new_n13825_));
  XOR2   g12823(.A(new_n13825_), .B(new_n13799_), .Y(new_n13826_));
  XOR2   g12824(.A(new_n13826_), .B(new_n13780_), .Y(new_n13827_));
  XOR2   g12825(.A(new_n13827_), .B(new_n13777_), .Y(new_n13828_));
  XOR2   g12826(.A(new_n13828_), .B(new_n13726_), .Y(new_n13829_));
  OAI21  g12827(.A0(new_n1761_), .A1(new_n1751_), .B0(new_n12558_), .Y(new_n13830_));
  NAND2  g12828(.A(new_n1766_), .B(new_n1687_), .Y(new_n13831_));
  AOI22  g12829(.A0(new_n1921_), .A1(new_n1906_), .B0(new_n13831_), .B1(new_n13830_), .Y(new_n13832_));
  NOR2   g12830(.A(new_n13832_), .B(new_n1915_), .Y(new_n13833_));
  XOR2   g12831(.A(new_n12634_), .B(new_n13833_), .Y(new_n13834_));
  OAI21  g12832(.A0(new_n1454_), .A1(new_n1219_), .B0(new_n1627_), .Y(new_n13835_));
  XOR2   g12833(.A(new_n12711_), .B(new_n13835_), .Y(new_n13836_));
  NAND2  g12834(.A(new_n13836_), .B(new_n13834_), .Y(new_n13837_));
  NOR2   g12835(.A(new_n13836_), .B(new_n13834_), .Y(new_n13838_));
  AOI21  g12836(.A0(new_n13837_), .A1(new_n12555_), .B0(new_n13838_), .Y(new_n13839_));
  AOI21  g12837(.A0(new_n1216_), .A1(new_n1207_), .B0(new_n1451_), .Y(new_n13840_));
  XOR2   g12838(.A(new_n12670_), .B(new_n13840_), .Y(new_n13841_));
  OAI22  g12839(.A0(new_n12710_), .A1(new_n13841_), .B0(new_n12636_), .B1(new_n1455_), .Y(new_n13842_));
  NAND2  g12840(.A(new_n12710_), .B(new_n13841_), .Y(new_n13843_));
  NAND2  g12841(.A(new_n13843_), .B(new_n13842_), .Y(new_n13844_));
  AOI22  g12842(.A0(new_n12708_), .A1(new_n12693_), .B0(new_n12673_), .B1(new_n1435_), .Y(new_n13845_));
  AOI22  g12843(.A0(new_n12691_), .A1(new_n12690_), .B0(new_n12689_), .B1(new_n12688_), .Y(new_n13846_));
  NOR4   g12844(.A(new_n12685_), .B(new_n12679_), .C(new_n12675_), .D(new_n1305_), .Y(new_n13847_));
  AOI22  g12845(.A0(new_n12706_), .A1(new_n12705_), .B0(new_n12704_), .B1(new_n12703_), .Y(new_n13848_));
  NOR4   g12846(.A(new_n12700_), .B(new_n12697_), .C(new_n12694_), .D(new_n1396_), .Y(new_n13849_));
  NOR4   g12847(.A(new_n13849_), .B(new_n13848_), .C(new_n13847_), .D(new_n13846_), .Y(new_n13850_));
  NOR3   g12848(.A(new_n12695_), .B(new_n12694_), .C(new_n1396_), .Y(new_n13851_));
  OAI21  g12849(.A0(new_n12694_), .A1(new_n1396_), .B0(new_n12695_), .Y(new_n13852_));
  OAI21  g12850(.A0(new_n13851_), .A1(new_n12696_), .B0(new_n13852_), .Y(new_n13853_));
  NOR3   g12851(.A(new_n12676_), .B(new_n12675_), .C(new_n1305_), .Y(new_n13854_));
  OAI21  g12852(.A0(new_n12675_), .A1(new_n1305_), .B0(new_n12676_), .Y(new_n13855_));
  OAI21  g12853(.A0(new_n13854_), .A1(new_n12678_), .B0(new_n13855_), .Y(new_n13856_));
  XOR2   g12854(.A(new_n13856_), .B(new_n13853_), .Y(new_n13857_));
  OAI21  g12855(.A0(new_n13850_), .A1(new_n13845_), .B0(new_n13857_), .Y(new_n13858_));
  NAND3  g12856(.A(new_n12680_), .B(new_n12689_), .C(new_n12688_), .Y(new_n13859_));
  AOI21  g12857(.A0(new_n12689_), .A1(new_n12688_), .B0(new_n12680_), .Y(new_n13860_));
  AOI21  g12858(.A0(new_n13859_), .A1(new_n12684_), .B0(new_n13860_), .Y(new_n13861_));
  AOI21  g12859(.A0(new_n13861_), .A1(new_n13853_), .B0(new_n13850_), .Y(new_n13862_));
  OAI21  g12860(.A0(new_n13861_), .A1(new_n13853_), .B0(new_n13862_), .Y(new_n13863_));
  OAI21  g12861(.A0(new_n13863_), .A1(new_n13845_), .B0(new_n13858_), .Y(new_n13864_));
  NAND2  g12862(.A(new_n12657_), .B(new_n12656_), .Y(new_n13865_));
  OAI21  g12863(.A0(new_n12667_), .A1(new_n12665_), .B0(new_n13865_), .Y(new_n13866_));
  NAND4  g12864(.A(new_n12662_), .B(new_n12659_), .C(new_n12657_), .D(new_n12656_), .Y(new_n13867_));
  AOI22  g12865(.A0(new_n13867_), .A1(new_n13866_), .B0(new_n12653_), .B1(new_n12648_), .Y(new_n13868_));
  AOI21  g12866(.A0(new_n12638_), .A1(new_n1217_), .B0(new_n13868_), .Y(new_n13869_));
  NOR2   g12867(.A(new_n12642_), .B(new_n12641_), .Y(new_n13870_));
  AOI21  g12868(.A0(new_n12652_), .A1(new_n12650_), .B0(new_n13870_), .Y(new_n13871_));
  NOR4   g12869(.A(new_n12647_), .B(new_n12644_), .C(new_n12642_), .D(new_n12641_), .Y(new_n13872_));
  OAI22  g12870(.A0(new_n12668_), .A1(new_n12663_), .B0(new_n13872_), .B1(new_n13871_), .Y(new_n13873_));
  NOR4   g12871(.A(new_n12668_), .B(new_n12663_), .C(new_n13872_), .D(new_n13871_), .Y(new_n13874_));
  AOI21  g12872(.A0(new_n13873_), .A1(new_n12639_), .B0(new_n13874_), .Y(new_n13875_));
  NAND3  g12873(.A(new_n12658_), .B(new_n12657_), .C(new_n12656_), .Y(new_n13876_));
  AOI22  g12874(.A0(new_n13876_), .A1(new_n12666_), .B0(new_n12660_), .B1(new_n13865_), .Y(new_n13877_));
  NOR3   g12875(.A(new_n12643_), .B(new_n12642_), .C(new_n12641_), .Y(new_n13878_));
  OAI22  g12876(.A0(new_n13878_), .A1(new_n12651_), .B0(new_n12645_), .B1(new_n13870_), .Y(new_n13879_));
  XOR2   g12877(.A(new_n13879_), .B(new_n13877_), .Y(new_n13880_));
  NAND4  g12878(.A(new_n13867_), .B(new_n13866_), .C(new_n12653_), .D(new_n12648_), .Y(new_n13881_));
  NOR3   g12879(.A(new_n12660_), .B(new_n12664_), .C(new_n1097_), .Y(new_n13882_));
  OAI21  g12880(.A0(new_n12664_), .A1(new_n1097_), .B0(new_n12660_), .Y(new_n13883_));
  OAI21  g12881(.A0(new_n13882_), .A1(new_n12661_), .B0(new_n13883_), .Y(new_n13884_));
  OAI221 g12882(.A0(new_n13878_), .A1(new_n12651_), .C0(new_n13884_), .B0(new_n12645_), .B1(new_n13870_), .Y(new_n13885_));
  NAND2  g12883(.A(new_n13879_), .B(new_n13877_), .Y(new_n13886_));
  NAND3  g12884(.A(new_n13886_), .B(new_n13885_), .C(new_n13881_), .Y(new_n13887_));
  OAI22  g12885(.A0(new_n13887_), .A1(new_n13869_), .B0(new_n13880_), .B1(new_n13875_), .Y(new_n13888_));
  XOR2   g12886(.A(new_n13888_), .B(new_n13864_), .Y(new_n13889_));
  XOR2   g12887(.A(new_n13889_), .B(new_n13844_), .Y(new_n13890_));
  NAND2  g12888(.A(new_n12633_), .B(new_n12596_), .Y(new_n13891_));
  OAI21  g12889(.A0(new_n13832_), .A1(new_n1915_), .B0(new_n13891_), .Y(new_n13892_));
  OAI22  g12890(.A0(new_n12592_), .A1(new_n12591_), .B0(new_n12590_), .B1(new_n12589_), .Y(new_n13893_));
  NAND4  g12891(.A(new_n12587_), .B(new_n12584_), .C(new_n12581_), .D(new_n1748_), .Y(new_n13894_));
  NAND2  g12892(.A(new_n13894_), .B(new_n13893_), .Y(new_n13895_));
  XOR2   g12893(.A(new_n13895_), .B(new_n12580_), .Y(new_n13896_));
  XOR2   g12894(.A(new_n13896_), .B(new_n12560_), .Y(new_n13897_));
  AOI21  g12895(.A0(new_n1907_), .A1(new_n1824_), .B0(new_n1899_), .Y(new_n13898_));
  XOR2   g12896(.A(new_n12632_), .B(new_n13898_), .Y(new_n13899_));
  NAND2  g12897(.A(new_n13899_), .B(new_n13897_), .Y(new_n13900_));
  NAND2  g12898(.A(new_n13900_), .B(new_n13892_), .Y(new_n13901_));
  OAI21  g12899(.A0(new_n12630_), .A1(new_n12626_), .B0(new_n12616_), .Y(new_n13902_));
  NAND4  g12900(.A(new_n12625_), .B(new_n12622_), .C(new_n12619_), .D(new_n12618_), .Y(new_n13903_));
  NAND3  g12901(.A(new_n13903_), .B(new_n12615_), .C(new_n12606_), .Y(new_n13904_));
  NOR2   g12902(.A(new_n13904_), .B(new_n12626_), .Y(new_n13905_));
  AOI21  g12903(.A0(new_n13902_), .A1(new_n12597_), .B0(new_n13905_), .Y(new_n13906_));
  NAND2  g12904(.A(new_n12619_), .B(new_n12618_), .Y(new_n13907_));
  NAND3  g12905(.A(new_n12620_), .B(new_n12619_), .C(new_n12618_), .Y(new_n13908_));
  AOI22  g12906(.A0(new_n13908_), .A1(new_n12621_), .B0(new_n12623_), .B1(new_n13907_), .Y(new_n13909_));
  NOR3   g12907(.A(new_n12613_), .B(new_n12602_), .C(new_n12600_), .Y(new_n13910_));
  OAI21  g12908(.A0(new_n12602_), .A1(new_n12600_), .B0(new_n12613_), .Y(new_n13911_));
  OAI21  g12909(.A0(new_n13910_), .A1(new_n12604_), .B0(new_n13911_), .Y(new_n13912_));
  XOR2   g12910(.A(new_n13912_), .B(new_n13909_), .Y(new_n13913_));
  NAND2  g12911(.A(new_n13902_), .B(new_n12597_), .Y(new_n13914_));
  NAND3  g12912(.A(new_n12603_), .B(new_n12607_), .C(new_n1821_), .Y(new_n13915_));
  AOI21  g12913(.A0(new_n12607_), .A1(new_n1821_), .B0(new_n12603_), .Y(new_n13916_));
  AOI21  g12914(.A0(new_n13915_), .A1(new_n12611_), .B0(new_n13916_), .Y(new_n13917_));
  AOI221 g12915(.A0(new_n13908_), .A1(new_n12621_), .C0(new_n13917_), .B0(new_n12623_), .B1(new_n13907_), .Y(new_n13918_));
  OAI22  g12916(.A0(new_n13912_), .A1(new_n13909_), .B0(new_n13904_), .B1(new_n12626_), .Y(new_n13919_));
  NOR2   g12917(.A(new_n13919_), .B(new_n13918_), .Y(new_n13920_));
  NAND2  g12918(.A(new_n13920_), .B(new_n13914_), .Y(new_n13921_));
  OAI21  g12919(.A0(new_n13913_), .A1(new_n13906_), .B0(new_n13921_), .Y(new_n13922_));
  AOI22  g12920(.A0(new_n12578_), .A1(new_n12577_), .B0(new_n12576_), .B1(new_n1684_), .Y(new_n13923_));
  NOR4   g12921(.A(new_n12574_), .B(new_n12568_), .C(new_n12565_), .D(new_n12563_), .Y(new_n13924_));
  OAI22  g12922(.A0(new_n12593_), .A1(new_n12588_), .B0(new_n13924_), .B1(new_n13923_), .Y(new_n13925_));
  NOR4   g12923(.A(new_n12593_), .B(new_n12588_), .C(new_n13924_), .D(new_n13923_), .Y(new_n13926_));
  AOI21  g12924(.A0(new_n13925_), .A1(new_n12560_), .B0(new_n13926_), .Y(new_n13927_));
  NOR3   g12925(.A(new_n12585_), .B(new_n12590_), .C(new_n12589_), .Y(new_n13928_));
  OAI21  g12926(.A0(new_n12590_), .A1(new_n12589_), .B0(new_n12585_), .Y(new_n13929_));
  OAI21  g12927(.A0(new_n13928_), .A1(new_n12586_), .B0(new_n13929_), .Y(new_n13930_));
  NAND3  g12928(.A(new_n12569_), .B(new_n12576_), .C(new_n1684_), .Y(new_n13931_));
  AOI21  g12929(.A0(new_n12576_), .A1(new_n1684_), .B0(new_n12569_), .Y(new_n13932_));
  AOI21  g12930(.A0(new_n13931_), .A1(new_n12573_), .B0(new_n13932_), .Y(new_n13933_));
  XOR2   g12931(.A(new_n13933_), .B(new_n13930_), .Y(new_n13934_));
  NAND2  g12932(.A(new_n13925_), .B(new_n12560_), .Y(new_n13935_));
  NOR2   g12933(.A(new_n13933_), .B(new_n13930_), .Y(new_n13936_));
  NAND4  g12934(.A(new_n13894_), .B(new_n13893_), .C(new_n12579_), .D(new_n12575_), .Y(new_n13937_));
  NAND3  g12935(.A(new_n12582_), .B(new_n12581_), .C(new_n1748_), .Y(new_n13938_));
  AOI21  g12936(.A0(new_n12581_), .A1(new_n1748_), .B0(new_n12582_), .Y(new_n13939_));
  AOI21  g12937(.A0(new_n13938_), .A1(new_n12583_), .B0(new_n13939_), .Y(new_n13940_));
  NOR3   g12938(.A(new_n12566_), .B(new_n12565_), .C(new_n12563_), .Y(new_n13941_));
  OAI21  g12939(.A0(new_n12565_), .A1(new_n12563_), .B0(new_n12566_), .Y(new_n13942_));
  OAI21  g12940(.A0(new_n13941_), .A1(new_n12567_), .B0(new_n13942_), .Y(new_n13943_));
  OAI21  g12941(.A0(new_n13943_), .A1(new_n13940_), .B0(new_n13937_), .Y(new_n13944_));
  NOR2   g12942(.A(new_n13944_), .B(new_n13936_), .Y(new_n13945_));
  NAND2  g12943(.A(new_n13945_), .B(new_n13935_), .Y(new_n13946_));
  OAI21  g12944(.A0(new_n13934_), .A1(new_n13927_), .B0(new_n13946_), .Y(new_n13947_));
  XOR2   g12945(.A(new_n13947_), .B(new_n13922_), .Y(new_n13948_));
  XOR2   g12946(.A(new_n13948_), .B(new_n13901_), .Y(new_n13949_));
  XOR2   g12947(.A(new_n13949_), .B(new_n13890_), .Y(new_n13950_));
  XOR2   g12948(.A(new_n13950_), .B(new_n13839_), .Y(new_n13951_));
  XOR2   g12949(.A(new_n13951_), .B(new_n13829_), .Y(new_n13952_));
  XOR2   g12950(.A(new_n13952_), .B(new_n13723_), .Y(new_n13953_));
  NOR2   g12951(.A(new_n12551_), .B(new_n12396_), .Y(new_n13954_));
  NAND2  g12952(.A(new_n12551_), .B(new_n12396_), .Y(new_n13955_));
  OAI21  g12953(.A0(new_n13954_), .A1(new_n13710_), .B0(new_n13955_), .Y(new_n13956_));
  OAI21  g12954(.A0(new_n3827_), .A1(new_n3817_), .B0(new_n12400_), .Y(new_n13957_));
  NAND2  g12955(.A(new_n3832_), .B(new_n3753_), .Y(new_n13958_));
  AOI22  g12956(.A0(new_n3839_), .A1(new_n3836_), .B0(new_n13958_), .B1(new_n13957_), .Y(new_n13959_));
  NOR2   g12957(.A(new_n13959_), .B(new_n4151_), .Y(new_n13960_));
  XOR2   g12958(.A(new_n12476_), .B(new_n13960_), .Y(new_n13961_));
  AOI22  g12959(.A0(new_n4131_), .A1(new_n4099_), .B0(new_n3972_), .B1(new_n3969_), .Y(new_n13962_));
  NOR2   g12960(.A(new_n13962_), .B(new_n4142_), .Y(new_n13963_));
  XOR2   g12961(.A(new_n12548_), .B(new_n13963_), .Y(new_n13964_));
  NAND2  g12962(.A(new_n13964_), .B(new_n13961_), .Y(new_n13965_));
  NOR2   g12963(.A(new_n13964_), .B(new_n13961_), .Y(new_n13966_));
  AOI21  g12964(.A0(new_n13965_), .A1(new_n12397_), .B0(new_n13966_), .Y(new_n13967_));
  AOI21  g12965(.A0(new_n4125_), .A1(new_n4123_), .B0(new_n3971_), .Y(new_n13968_));
  XOR2   g12966(.A(new_n12513_), .B(new_n13968_), .Y(new_n13969_));
  AOI21  g12967(.A0(new_n4114_), .A1(new_n4107_), .B0(new_n4101_), .Y(new_n13970_));
  XOR2   g12968(.A(new_n12546_), .B(new_n13970_), .Y(new_n13971_));
  OAI22  g12969(.A0(new_n13971_), .A1(new_n13969_), .B0(new_n13962_), .B1(new_n4142_), .Y(new_n13972_));
  NAND2  g12970(.A(new_n13971_), .B(new_n13969_), .Y(new_n13973_));
  NAND2  g12971(.A(new_n13973_), .B(new_n13972_), .Y(new_n13974_));
  OAI21  g12972(.A0(new_n4028_), .A1(new_n4011_), .B0(new_n4114_), .Y(new_n13975_));
  NAND2  g12973(.A(new_n12533_), .B(new_n12532_), .Y(new_n13976_));
  OAI21  g12974(.A0(new_n12543_), .A1(new_n12542_), .B0(new_n13976_), .Y(new_n13977_));
  NAND4  g12975(.A(new_n12539_), .B(new_n12536_), .C(new_n12533_), .D(new_n12532_), .Y(new_n13978_));
  AOI22  g12976(.A0(new_n13978_), .A1(new_n13977_), .B0(new_n12529_), .B1(new_n12524_), .Y(new_n13979_));
  AOI21  g12977(.A0(new_n13975_), .A1(new_n4115_), .B0(new_n13979_), .Y(new_n13980_));
  NOR2   g12978(.A(new_n12518_), .B(new_n12517_), .Y(new_n13981_));
  AOI21  g12979(.A0(new_n12528_), .A1(new_n12526_), .B0(new_n13981_), .Y(new_n13982_));
  NOR4   g12980(.A(new_n12523_), .B(new_n12520_), .C(new_n12518_), .D(new_n12517_), .Y(new_n13983_));
  NOR4   g12981(.A(new_n12544_), .B(new_n12540_), .C(new_n13983_), .D(new_n13982_), .Y(new_n13984_));
  NAND3  g12982(.A(new_n12534_), .B(new_n12533_), .C(new_n12532_), .Y(new_n13985_));
  AOI22  g12983(.A0(new_n13985_), .A1(new_n12535_), .B0(new_n12537_), .B1(new_n13976_), .Y(new_n13986_));
  NOR3   g12984(.A(new_n12519_), .B(new_n12518_), .C(new_n12517_), .Y(new_n13987_));
  OAI22  g12985(.A0(new_n13987_), .A1(new_n12527_), .B0(new_n12521_), .B1(new_n13981_), .Y(new_n13988_));
  NOR2   g12986(.A(new_n13988_), .B(new_n13986_), .Y(new_n13989_));
  NAND2  g12987(.A(new_n13985_), .B(new_n12535_), .Y(new_n13990_));
  NAND2  g12988(.A(new_n12537_), .B(new_n13976_), .Y(new_n13991_));
  NAND2  g12989(.A(new_n13991_), .B(new_n13990_), .Y(new_n13992_));
  NOR2   g12990(.A(new_n13987_), .B(new_n12527_), .Y(new_n13993_));
  NOR2   g12991(.A(new_n12521_), .B(new_n13981_), .Y(new_n13994_));
  NOR2   g12992(.A(new_n13994_), .B(new_n13993_), .Y(new_n13995_));
  NOR2   g12993(.A(new_n13995_), .B(new_n13992_), .Y(new_n13996_));
  OAI22  g12994(.A0(new_n13996_), .A1(new_n13989_), .B0(new_n13984_), .B1(new_n13980_), .Y(new_n13997_));
  NAND2  g12995(.A(new_n13988_), .B(new_n13986_), .Y(new_n13998_));
  NOR2   g12996(.A(new_n13989_), .B(new_n13984_), .Y(new_n13999_));
  OAI211 g12997(.A0(new_n13979_), .A1(new_n13970_), .B0(new_n13999_), .B1(new_n13998_), .Y(new_n14000_));
  NAND2  g12998(.A(new_n14000_), .B(new_n13997_), .Y(new_n14001_));
  OAI21  g12999(.A0(new_n3967_), .A1(new_n3950_), .B0(new_n4125_), .Y(new_n14002_));
  OAI22  g13000(.A0(new_n12510_), .A1(new_n12509_), .B0(new_n12508_), .B1(new_n12506_), .Y(new_n14003_));
  NAND4  g13001(.A(new_n12504_), .B(new_n12501_), .C(new_n12498_), .D(new_n12497_), .Y(new_n14004_));
  NAND2  g13002(.A(new_n14004_), .B(new_n14003_), .Y(new_n14005_));
  AOI22  g13003(.A0(new_n14005_), .A1(new_n12495_), .B0(new_n14002_), .B1(new_n4127_), .Y(new_n14006_));
  NOR2   g13004(.A(new_n12483_), .B(new_n12482_), .Y(new_n14007_));
  AOI21  g13005(.A0(new_n12493_), .A1(new_n12491_), .B0(new_n14007_), .Y(new_n14008_));
  NOR4   g13006(.A(new_n12488_), .B(new_n12485_), .C(new_n12483_), .D(new_n12482_), .Y(new_n14009_));
  NOR4   g13007(.A(new_n12511_), .B(new_n12505_), .C(new_n14009_), .D(new_n14008_), .Y(new_n14010_));
  NAND3  g13008(.A(new_n12499_), .B(new_n12498_), .C(new_n12497_), .Y(new_n14011_));
  AOI21  g13009(.A0(new_n12498_), .A1(new_n12497_), .B0(new_n12499_), .Y(new_n14012_));
  AOI21  g13010(.A0(new_n14011_), .A1(new_n12500_), .B0(new_n14012_), .Y(new_n14013_));
  NOR3   g13011(.A(new_n12484_), .B(new_n12483_), .C(new_n12482_), .Y(new_n14014_));
  OAI22  g13012(.A0(new_n14014_), .A1(new_n12492_), .B0(new_n12486_), .B1(new_n14007_), .Y(new_n14015_));
  NOR2   g13013(.A(new_n14015_), .B(new_n14013_), .Y(new_n14016_));
  NOR3   g13014(.A(new_n12502_), .B(new_n12508_), .C(new_n12506_), .Y(new_n14017_));
  OAI21  g13015(.A0(new_n12508_), .A1(new_n12506_), .B0(new_n12502_), .Y(new_n14018_));
  OAI21  g13016(.A0(new_n14017_), .A1(new_n12503_), .B0(new_n14018_), .Y(new_n14019_));
  NAND2  g13017(.A(new_n12486_), .B(new_n3966_), .Y(new_n14020_));
  OAI21  g13018(.A0(new_n14020_), .A1(new_n12483_), .B0(new_n12487_), .Y(new_n14021_));
  OAI21  g13019(.A0(new_n12483_), .A1(new_n12482_), .B0(new_n12484_), .Y(new_n14022_));
  AOI21  g13020(.A0(new_n14022_), .A1(new_n14021_), .B0(new_n14019_), .Y(new_n14023_));
  OAI22  g13021(.A0(new_n14023_), .A1(new_n14016_), .B0(new_n14010_), .B1(new_n14006_), .Y(new_n14024_));
  OAI21  g13022(.A0(new_n14009_), .A1(new_n14008_), .B0(new_n14005_), .Y(new_n14025_));
  NAND2  g13023(.A(new_n14025_), .B(new_n12480_), .Y(new_n14026_));
  NOR3   g13024(.A(new_n14023_), .B(new_n14016_), .C(new_n14010_), .Y(new_n14027_));
  NAND2  g13025(.A(new_n14027_), .B(new_n14026_), .Y(new_n14028_));
  NAND2  g13026(.A(new_n14028_), .B(new_n14024_), .Y(new_n14029_));
  XOR2   g13027(.A(new_n14029_), .B(new_n14001_), .Y(new_n14030_));
  XOR2   g13028(.A(new_n14030_), .B(new_n13974_), .Y(new_n14031_));
  NAND2  g13029(.A(new_n12475_), .B(new_n12438_), .Y(new_n14032_));
  OAI21  g13030(.A0(new_n13959_), .A1(new_n4151_), .B0(new_n14032_), .Y(new_n14033_));
  OAI22  g13031(.A0(new_n12434_), .A1(new_n12433_), .B0(new_n12432_), .B1(new_n12431_), .Y(new_n14034_));
  NAND4  g13032(.A(new_n12429_), .B(new_n12426_), .C(new_n12423_), .D(new_n3814_), .Y(new_n14035_));
  NAND2  g13033(.A(new_n14035_), .B(new_n14034_), .Y(new_n14036_));
  XOR2   g13034(.A(new_n14036_), .B(new_n12422_), .Y(new_n14037_));
  XOR2   g13035(.A(new_n14037_), .B(new_n12402_), .Y(new_n14038_));
  AOI21  g13036(.A0(new_n3837_), .A1(new_n3614_), .B0(new_n3689_), .Y(new_n14039_));
  XOR2   g13037(.A(new_n12474_), .B(new_n14039_), .Y(new_n14040_));
  NAND2  g13038(.A(new_n14040_), .B(new_n14038_), .Y(new_n14041_));
  NAND2  g13039(.A(new_n14041_), .B(new_n14033_), .Y(new_n14042_));
  OAI21  g13040(.A0(new_n12472_), .A1(new_n12468_), .B0(new_n12458_), .Y(new_n14043_));
  NAND4  g13041(.A(new_n12467_), .B(new_n12464_), .C(new_n12461_), .D(new_n12460_), .Y(new_n14044_));
  NAND3  g13042(.A(new_n14044_), .B(new_n12457_), .C(new_n12448_), .Y(new_n14045_));
  NOR2   g13043(.A(new_n14045_), .B(new_n12468_), .Y(new_n14046_));
  AOI21  g13044(.A0(new_n14043_), .A1(new_n12439_), .B0(new_n14046_), .Y(new_n14047_));
  NAND2  g13045(.A(new_n12461_), .B(new_n12460_), .Y(new_n14048_));
  NAND3  g13046(.A(new_n12462_), .B(new_n12461_), .C(new_n12460_), .Y(new_n14049_));
  AOI22  g13047(.A0(new_n14049_), .A1(new_n12463_), .B0(new_n12465_), .B1(new_n14048_), .Y(new_n14050_));
  NOR3   g13048(.A(new_n12455_), .B(new_n12444_), .C(new_n12442_), .Y(new_n14051_));
  OAI21  g13049(.A0(new_n12444_), .A1(new_n12442_), .B0(new_n12455_), .Y(new_n14052_));
  OAI21  g13050(.A0(new_n14051_), .A1(new_n12446_), .B0(new_n14052_), .Y(new_n14053_));
  XOR2   g13051(.A(new_n14053_), .B(new_n14050_), .Y(new_n14054_));
  NAND2  g13052(.A(new_n14043_), .B(new_n12439_), .Y(new_n14055_));
  NAND3  g13053(.A(new_n12445_), .B(new_n12449_), .C(new_n3611_), .Y(new_n14056_));
  AOI21  g13054(.A0(new_n12449_), .A1(new_n3611_), .B0(new_n12445_), .Y(new_n14057_));
  AOI21  g13055(.A0(new_n14056_), .A1(new_n12453_), .B0(new_n14057_), .Y(new_n14058_));
  AOI221 g13056(.A0(new_n14049_), .A1(new_n12463_), .C0(new_n14058_), .B0(new_n12465_), .B1(new_n14048_), .Y(new_n14059_));
  OAI22  g13057(.A0(new_n14053_), .A1(new_n14050_), .B0(new_n14045_), .B1(new_n12468_), .Y(new_n14060_));
  NOR2   g13058(.A(new_n14060_), .B(new_n14059_), .Y(new_n14061_));
  NAND2  g13059(.A(new_n14061_), .B(new_n14055_), .Y(new_n14062_));
  OAI21  g13060(.A0(new_n14054_), .A1(new_n14047_), .B0(new_n14062_), .Y(new_n14063_));
  AOI22  g13061(.A0(new_n12420_), .A1(new_n12419_), .B0(new_n12418_), .B1(new_n3750_), .Y(new_n14064_));
  NOR4   g13062(.A(new_n12416_), .B(new_n12410_), .C(new_n12407_), .D(new_n12405_), .Y(new_n14065_));
  OAI22  g13063(.A0(new_n12435_), .A1(new_n12430_), .B0(new_n14065_), .B1(new_n14064_), .Y(new_n14066_));
  NOR4   g13064(.A(new_n12435_), .B(new_n12430_), .C(new_n14065_), .D(new_n14064_), .Y(new_n14067_));
  AOI21  g13065(.A0(new_n14066_), .A1(new_n12402_), .B0(new_n14067_), .Y(new_n14068_));
  NOR3   g13066(.A(new_n12427_), .B(new_n12432_), .C(new_n12431_), .Y(new_n14069_));
  OAI21  g13067(.A0(new_n12432_), .A1(new_n12431_), .B0(new_n12427_), .Y(new_n14070_));
  OAI21  g13068(.A0(new_n14069_), .A1(new_n12428_), .B0(new_n14070_), .Y(new_n14071_));
  NAND3  g13069(.A(new_n12411_), .B(new_n12418_), .C(new_n3750_), .Y(new_n14072_));
  AOI21  g13070(.A0(new_n12418_), .A1(new_n3750_), .B0(new_n12411_), .Y(new_n14073_));
  AOI21  g13071(.A0(new_n14072_), .A1(new_n12415_), .B0(new_n14073_), .Y(new_n14074_));
  XOR2   g13072(.A(new_n14074_), .B(new_n14071_), .Y(new_n14075_));
  NAND2  g13073(.A(new_n14066_), .B(new_n12402_), .Y(new_n14076_));
  NOR2   g13074(.A(new_n14074_), .B(new_n14071_), .Y(new_n14077_));
  NAND4  g13075(.A(new_n14035_), .B(new_n14034_), .C(new_n12421_), .D(new_n12417_), .Y(new_n14078_));
  NAND3  g13076(.A(new_n12424_), .B(new_n12423_), .C(new_n3814_), .Y(new_n14079_));
  AOI21  g13077(.A0(new_n12423_), .A1(new_n3814_), .B0(new_n12424_), .Y(new_n14080_));
  AOI21  g13078(.A0(new_n14079_), .A1(new_n12425_), .B0(new_n14080_), .Y(new_n14081_));
  NOR3   g13079(.A(new_n12408_), .B(new_n12407_), .C(new_n12405_), .Y(new_n14082_));
  OAI21  g13080(.A0(new_n12407_), .A1(new_n12405_), .B0(new_n12408_), .Y(new_n14083_));
  OAI21  g13081(.A0(new_n14082_), .A1(new_n12409_), .B0(new_n14083_), .Y(new_n14084_));
  OAI21  g13082(.A0(new_n14084_), .A1(new_n14081_), .B0(new_n14078_), .Y(new_n14085_));
  NOR2   g13083(.A(new_n14085_), .B(new_n14077_), .Y(new_n14086_));
  NAND2  g13084(.A(new_n14086_), .B(new_n14076_), .Y(new_n14087_));
  OAI21  g13085(.A0(new_n14075_), .A1(new_n14068_), .B0(new_n14087_), .Y(new_n14088_));
  XOR2   g13086(.A(new_n14088_), .B(new_n14063_), .Y(new_n14089_));
  XOR2   g13087(.A(new_n14089_), .B(new_n14042_), .Y(new_n14090_));
  XOR2   g13088(.A(new_n14090_), .B(new_n14031_), .Y(new_n14091_));
  XOR2   g13089(.A(new_n14091_), .B(new_n13967_), .Y(new_n14092_));
  AOI21  g13090(.A0(new_n4760_), .A1(new_n4751_), .B0(new_n4753_), .Y(new_n14093_));
  NOR2   g13091(.A(new_n12394_), .B(new_n12322_), .Y(new_n14094_));
  NAND2  g13092(.A(new_n12394_), .B(new_n12322_), .Y(new_n14095_));
  OAI21  g13093(.A0(new_n14094_), .A1(new_n14093_), .B0(new_n14095_), .Y(new_n14096_));
  AOI22  g13094(.A0(new_n4454_), .A1(new_n4422_), .B0(new_n4295_), .B1(new_n4292_), .Y(new_n14097_));
  AOI21  g13095(.A0(new_n4448_), .A1(new_n4446_), .B0(new_n4294_), .Y(new_n14098_));
  XOR2   g13096(.A(new_n12358_), .B(new_n14098_), .Y(new_n14099_));
  AOI21  g13097(.A0(new_n4437_), .A1(new_n4430_), .B0(new_n4424_), .Y(new_n14100_));
  XOR2   g13098(.A(new_n12391_), .B(new_n14100_), .Y(new_n14101_));
  OAI22  g13099(.A0(new_n14101_), .A1(new_n14099_), .B0(new_n14097_), .B1(new_n4465_), .Y(new_n14102_));
  NAND2  g13100(.A(new_n14101_), .B(new_n14099_), .Y(new_n14103_));
  NAND2  g13101(.A(new_n14103_), .B(new_n14102_), .Y(new_n14104_));
  OAI21  g13102(.A0(new_n4351_), .A1(new_n4334_), .B0(new_n4437_), .Y(new_n14105_));
  NAND2  g13103(.A(new_n12378_), .B(new_n12377_), .Y(new_n14106_));
  OAI21  g13104(.A0(new_n12388_), .A1(new_n12387_), .B0(new_n14106_), .Y(new_n14107_));
  NAND4  g13105(.A(new_n12384_), .B(new_n12381_), .C(new_n12378_), .D(new_n12377_), .Y(new_n14108_));
  AOI22  g13106(.A0(new_n14108_), .A1(new_n14107_), .B0(new_n12374_), .B1(new_n12369_), .Y(new_n14109_));
  AOI21  g13107(.A0(new_n14105_), .A1(new_n4438_), .B0(new_n14109_), .Y(new_n14110_));
  NOR2   g13108(.A(new_n12363_), .B(new_n12362_), .Y(new_n14111_));
  AOI21  g13109(.A0(new_n12373_), .A1(new_n12371_), .B0(new_n14111_), .Y(new_n14112_));
  NOR4   g13110(.A(new_n12368_), .B(new_n12365_), .C(new_n12363_), .D(new_n12362_), .Y(new_n14113_));
  NOR4   g13111(.A(new_n12389_), .B(new_n12385_), .C(new_n14113_), .D(new_n14112_), .Y(new_n14114_));
  NAND3  g13112(.A(new_n12379_), .B(new_n12378_), .C(new_n12377_), .Y(new_n14115_));
  AOI22  g13113(.A0(new_n14115_), .A1(new_n12380_), .B0(new_n12382_), .B1(new_n14106_), .Y(new_n14116_));
  NOR3   g13114(.A(new_n12364_), .B(new_n12363_), .C(new_n12362_), .Y(new_n14117_));
  OAI22  g13115(.A0(new_n14117_), .A1(new_n12372_), .B0(new_n12366_), .B1(new_n14111_), .Y(new_n14118_));
  NOR2   g13116(.A(new_n14118_), .B(new_n14116_), .Y(new_n14119_));
  NAND2  g13117(.A(new_n14115_), .B(new_n12380_), .Y(new_n14120_));
  NAND2  g13118(.A(new_n12382_), .B(new_n14106_), .Y(new_n14121_));
  NAND2  g13119(.A(new_n14121_), .B(new_n14120_), .Y(new_n14122_));
  NOR2   g13120(.A(new_n14117_), .B(new_n12372_), .Y(new_n14123_));
  NOR2   g13121(.A(new_n12366_), .B(new_n14111_), .Y(new_n14124_));
  NOR2   g13122(.A(new_n14124_), .B(new_n14123_), .Y(new_n14125_));
  NOR2   g13123(.A(new_n14125_), .B(new_n14122_), .Y(new_n14126_));
  OAI22  g13124(.A0(new_n14126_), .A1(new_n14119_), .B0(new_n14114_), .B1(new_n14110_), .Y(new_n14127_));
  NAND2  g13125(.A(new_n14118_), .B(new_n14116_), .Y(new_n14128_));
  NOR2   g13126(.A(new_n14119_), .B(new_n14114_), .Y(new_n14129_));
  OAI211 g13127(.A0(new_n14109_), .A1(new_n14100_), .B0(new_n14129_), .B1(new_n14128_), .Y(new_n14130_));
  NAND2  g13128(.A(new_n14130_), .B(new_n14127_), .Y(new_n14131_));
  OAI21  g13129(.A0(new_n4290_), .A1(new_n4273_), .B0(new_n4448_), .Y(new_n14132_));
  OAI22  g13130(.A0(new_n12355_), .A1(new_n12354_), .B0(new_n12353_), .B1(new_n12351_), .Y(new_n14133_));
  NAND4  g13131(.A(new_n12349_), .B(new_n12346_), .C(new_n12343_), .D(new_n12342_), .Y(new_n14134_));
  NAND2  g13132(.A(new_n14134_), .B(new_n14133_), .Y(new_n14135_));
  AOI22  g13133(.A0(new_n14135_), .A1(new_n12340_), .B0(new_n14132_), .B1(new_n4450_), .Y(new_n14136_));
  NOR2   g13134(.A(new_n12328_), .B(new_n12327_), .Y(new_n14137_));
  AOI21  g13135(.A0(new_n12338_), .A1(new_n12336_), .B0(new_n14137_), .Y(new_n14138_));
  NOR4   g13136(.A(new_n12333_), .B(new_n12330_), .C(new_n12328_), .D(new_n12327_), .Y(new_n14139_));
  NOR4   g13137(.A(new_n12356_), .B(new_n12350_), .C(new_n14139_), .D(new_n14138_), .Y(new_n14140_));
  NAND3  g13138(.A(new_n12344_), .B(new_n12343_), .C(new_n12342_), .Y(new_n14141_));
  AOI21  g13139(.A0(new_n12343_), .A1(new_n12342_), .B0(new_n12344_), .Y(new_n14142_));
  AOI21  g13140(.A0(new_n14141_), .A1(new_n12345_), .B0(new_n14142_), .Y(new_n14143_));
  NOR3   g13141(.A(new_n12329_), .B(new_n12328_), .C(new_n12327_), .Y(new_n14144_));
  OAI22  g13142(.A0(new_n14144_), .A1(new_n12337_), .B0(new_n12331_), .B1(new_n14137_), .Y(new_n14145_));
  NOR2   g13143(.A(new_n14145_), .B(new_n14143_), .Y(new_n14146_));
  NOR3   g13144(.A(new_n12347_), .B(new_n12353_), .C(new_n12351_), .Y(new_n14147_));
  OAI21  g13145(.A0(new_n12353_), .A1(new_n12351_), .B0(new_n12347_), .Y(new_n14148_));
  OAI21  g13146(.A0(new_n14147_), .A1(new_n12348_), .B0(new_n14148_), .Y(new_n14149_));
  NAND2  g13147(.A(new_n12331_), .B(new_n4289_), .Y(new_n14150_));
  OAI21  g13148(.A0(new_n14150_), .A1(new_n12328_), .B0(new_n12332_), .Y(new_n14151_));
  OAI21  g13149(.A0(new_n12328_), .A1(new_n12327_), .B0(new_n12329_), .Y(new_n14152_));
  AOI21  g13150(.A0(new_n14152_), .A1(new_n14151_), .B0(new_n14149_), .Y(new_n14153_));
  OAI22  g13151(.A0(new_n14153_), .A1(new_n14146_), .B0(new_n14140_), .B1(new_n14136_), .Y(new_n14154_));
  OAI21  g13152(.A0(new_n14139_), .A1(new_n14138_), .B0(new_n14135_), .Y(new_n14155_));
  NAND2  g13153(.A(new_n14155_), .B(new_n12325_), .Y(new_n14156_));
  NOR3   g13154(.A(new_n14153_), .B(new_n14146_), .C(new_n14140_), .Y(new_n14157_));
  NAND2  g13155(.A(new_n14157_), .B(new_n14156_), .Y(new_n14158_));
  NAND2  g13156(.A(new_n14158_), .B(new_n14154_), .Y(new_n14159_));
  XOR2   g13157(.A(new_n14159_), .B(new_n14131_), .Y(new_n14160_));
  XOR2   g13158(.A(new_n14160_), .B(new_n14104_), .Y(new_n14161_));
  OAI21  g13159(.A0(new_n4726_), .A1(new_n4715_), .B0(new_n12245_), .Y(new_n14162_));
  NAND2  g13160(.A(new_n4731_), .B(new_n4651_), .Y(new_n14163_));
  AOI22  g13161(.A0(new_n4738_), .A1(new_n4735_), .B0(new_n14163_), .B1(new_n14162_), .Y(new_n14164_));
  NAND2  g13162(.A(new_n12320_), .B(new_n12283_), .Y(new_n14165_));
  OAI21  g13163(.A0(new_n14164_), .A1(new_n4749_), .B0(new_n14165_), .Y(new_n14166_));
  OAI22  g13164(.A0(new_n12279_), .A1(new_n12278_), .B0(new_n12277_), .B1(new_n12276_), .Y(new_n14167_));
  NAND4  g13165(.A(new_n12274_), .B(new_n12271_), .C(new_n12268_), .D(new_n4712_), .Y(new_n14168_));
  NAND2  g13166(.A(new_n14168_), .B(new_n14167_), .Y(new_n14169_));
  XOR2   g13167(.A(new_n14169_), .B(new_n12267_), .Y(new_n14170_));
  XOR2   g13168(.A(new_n14170_), .B(new_n12247_), .Y(new_n14171_));
  AOI21  g13169(.A0(new_n4736_), .A1(new_n4524_), .B0(new_n4599_), .Y(new_n14172_));
  XOR2   g13170(.A(new_n12319_), .B(new_n14172_), .Y(new_n14173_));
  NAND2  g13171(.A(new_n14173_), .B(new_n14171_), .Y(new_n14174_));
  NAND2  g13172(.A(new_n14174_), .B(new_n14166_), .Y(new_n14175_));
  OAI21  g13173(.A0(new_n12317_), .A1(new_n12313_), .B0(new_n12303_), .Y(new_n14176_));
  NAND4  g13174(.A(new_n12312_), .B(new_n12309_), .C(new_n12306_), .D(new_n12305_), .Y(new_n14177_));
  NAND3  g13175(.A(new_n14177_), .B(new_n12302_), .C(new_n12293_), .Y(new_n14178_));
  NOR2   g13176(.A(new_n14178_), .B(new_n12313_), .Y(new_n14179_));
  AOI21  g13177(.A0(new_n14176_), .A1(new_n12284_), .B0(new_n14179_), .Y(new_n14180_));
  NAND2  g13178(.A(new_n12306_), .B(new_n12305_), .Y(new_n14181_));
  NAND3  g13179(.A(new_n12307_), .B(new_n12306_), .C(new_n12305_), .Y(new_n14182_));
  AOI22  g13180(.A0(new_n14182_), .A1(new_n12308_), .B0(new_n12310_), .B1(new_n14181_), .Y(new_n14183_));
  NOR3   g13181(.A(new_n12300_), .B(new_n12289_), .C(new_n12287_), .Y(new_n14184_));
  OAI21  g13182(.A0(new_n12289_), .A1(new_n12287_), .B0(new_n12300_), .Y(new_n14185_));
  OAI21  g13183(.A0(new_n14184_), .A1(new_n12291_), .B0(new_n14185_), .Y(new_n14186_));
  XOR2   g13184(.A(new_n14186_), .B(new_n14183_), .Y(new_n14187_));
  NAND2  g13185(.A(new_n14176_), .B(new_n12284_), .Y(new_n14188_));
  NAND3  g13186(.A(new_n12290_), .B(new_n12294_), .C(new_n4521_), .Y(new_n14189_));
  AOI21  g13187(.A0(new_n12294_), .A1(new_n4521_), .B0(new_n12290_), .Y(new_n14190_));
  AOI21  g13188(.A0(new_n14189_), .A1(new_n12298_), .B0(new_n14190_), .Y(new_n14191_));
  AOI221 g13189(.A0(new_n14182_), .A1(new_n12308_), .C0(new_n14191_), .B0(new_n12310_), .B1(new_n14181_), .Y(new_n14192_));
  OAI22  g13190(.A0(new_n14186_), .A1(new_n14183_), .B0(new_n14178_), .B1(new_n12313_), .Y(new_n14193_));
  NOR2   g13191(.A(new_n14193_), .B(new_n14192_), .Y(new_n14194_));
  NAND2  g13192(.A(new_n14194_), .B(new_n14188_), .Y(new_n14195_));
  OAI21  g13193(.A0(new_n14187_), .A1(new_n14180_), .B0(new_n14195_), .Y(new_n14196_));
  AOI22  g13194(.A0(new_n12265_), .A1(new_n12264_), .B0(new_n12263_), .B1(new_n4648_), .Y(new_n14197_));
  NOR4   g13195(.A(new_n12261_), .B(new_n12255_), .C(new_n12252_), .D(new_n12250_), .Y(new_n14198_));
  OAI22  g13196(.A0(new_n12280_), .A1(new_n12275_), .B0(new_n14198_), .B1(new_n14197_), .Y(new_n14199_));
  NOR4   g13197(.A(new_n12280_), .B(new_n12275_), .C(new_n14198_), .D(new_n14197_), .Y(new_n14200_));
  AOI21  g13198(.A0(new_n14199_), .A1(new_n12247_), .B0(new_n14200_), .Y(new_n14201_));
  NOR3   g13199(.A(new_n12272_), .B(new_n12277_), .C(new_n12276_), .Y(new_n14202_));
  OAI21  g13200(.A0(new_n12277_), .A1(new_n12276_), .B0(new_n12272_), .Y(new_n14203_));
  OAI21  g13201(.A0(new_n14202_), .A1(new_n12273_), .B0(new_n14203_), .Y(new_n14204_));
  NAND3  g13202(.A(new_n12256_), .B(new_n12263_), .C(new_n4648_), .Y(new_n14205_));
  AOI21  g13203(.A0(new_n12263_), .A1(new_n4648_), .B0(new_n12256_), .Y(new_n14206_));
  AOI21  g13204(.A0(new_n14205_), .A1(new_n12260_), .B0(new_n14206_), .Y(new_n14207_));
  XOR2   g13205(.A(new_n14207_), .B(new_n14204_), .Y(new_n14208_));
  NAND2  g13206(.A(new_n14199_), .B(new_n12247_), .Y(new_n14209_));
  NAND4  g13207(.A(new_n14168_), .B(new_n14167_), .C(new_n12266_), .D(new_n12262_), .Y(new_n14210_));
  NAND2  g13208(.A(new_n14207_), .B(new_n14204_), .Y(new_n14211_));
  NOR3   g13209(.A(new_n12253_), .B(new_n12252_), .C(new_n12250_), .Y(new_n14212_));
  OAI21  g13210(.A0(new_n12252_), .A1(new_n12250_), .B0(new_n12253_), .Y(new_n14213_));
  OAI21  g13211(.A0(new_n14212_), .A1(new_n12254_), .B0(new_n14213_), .Y(new_n14214_));
  OAI211 g13212(.A0(new_n14202_), .A1(new_n12273_), .B0(new_n14214_), .B1(new_n14203_), .Y(new_n14215_));
  NAND4  g13213(.A(new_n14215_), .B(new_n14211_), .C(new_n14210_), .D(new_n14209_), .Y(new_n14216_));
  OAI21  g13214(.A0(new_n14208_), .A1(new_n14201_), .B0(new_n14216_), .Y(new_n14217_));
  XOR2   g13215(.A(new_n14217_), .B(new_n14196_), .Y(new_n14218_));
  XOR2   g13216(.A(new_n14218_), .B(new_n14175_), .Y(new_n14219_));
  XOR2   g13217(.A(new_n14219_), .B(new_n14161_), .Y(new_n14220_));
  XOR2   g13218(.A(new_n14220_), .B(new_n14096_), .Y(new_n14221_));
  XOR2   g13219(.A(new_n14221_), .B(new_n14092_), .Y(new_n14222_));
  XOR2   g13220(.A(new_n14222_), .B(new_n13956_), .Y(new_n14223_));
  XOR2   g13221(.A(new_n14223_), .B(new_n13953_), .Y(new_n14224_));
  XOR2   g13222(.A(new_n14224_), .B(new_n13716_), .Y(new_n14225_));
  NOR2   g13223(.A(new_n14225_), .B(new_n13709_), .Y(new_n14226_));
  OAI21  g13224(.A0(new_n13708_), .A1(new_n13702_), .B0(new_n14225_), .Y(new_n14227_));
  OAI22  g13225(.A0(new_n14227_), .A1(new_n13697_), .B0(new_n14226_), .B1(new_n12892_), .Y(new_n14228_));
  NOR2   g13226(.A(new_n11606_), .B(new_n13381_), .Y(new_n14229_));
  OAI22  g13227(.A0(new_n13382_), .A1(new_n11444_), .B0(new_n14229_), .B1(new_n13698_), .Y(new_n14230_));
  XOR2   g13228(.A(new_n13694_), .B(new_n14230_), .Y(new_n14231_));
  NAND2  g13229(.A(new_n14231_), .B(new_n13707_), .Y(new_n14232_));
  NOR2   g13230(.A(new_n14231_), .B(new_n13707_), .Y(new_n14233_));
  AOI21  g13231(.A0(new_n14232_), .A1(new_n12895_), .B0(new_n14233_), .Y(new_n14234_));
  XOR2   g13232(.A(new_n11522_), .B(new_n13623_), .Y(new_n14235_));
  XOR2   g13233(.A(new_n11594_), .B(new_n13558_), .Y(new_n14236_));
  NAND2  g13234(.A(new_n14236_), .B(new_n14235_), .Y(new_n14237_));
  NOR2   g13235(.A(new_n14236_), .B(new_n14235_), .Y(new_n14238_));
  AOI21  g13236(.A0(new_n14237_), .A1(new_n13380_), .B0(new_n14238_), .Y(new_n14239_));
  XOR2   g13237(.A(new_n13689_), .B(new_n14239_), .Y(new_n14240_));
  NAND2  g13238(.A(new_n14240_), .B(new_n13554_), .Y(new_n14241_));
  AOI21  g13239(.A0(new_n13553_), .A1(new_n13692_), .B0(new_n14240_), .Y(new_n14242_));
  AOI22  g13240(.A0(new_n14242_), .A1(new_n13552_), .B0(new_n14241_), .B1(new_n14230_), .Y(new_n14243_));
  XOR2   g13241(.A(new_n13480_), .B(new_n13542_), .Y(new_n14244_));
  NAND2  g13242(.A(new_n13537_), .B(new_n14244_), .Y(new_n14245_));
  NAND2  g13243(.A(new_n11434_), .B(new_n11403_), .Y(new_n14246_));
  NOR2   g13244(.A(new_n11434_), .B(new_n11403_), .Y(new_n14247_));
  AOI21  g13245(.A0(new_n14246_), .A1(new_n11365_), .B0(new_n14247_), .Y(new_n14248_));
  XOR2   g13246(.A(new_n13536_), .B(new_n14248_), .Y(new_n14249_));
  OAI21  g13247(.A0(new_n13550_), .A1(new_n13542_), .B0(new_n14249_), .Y(new_n14250_));
  NOR2   g13248(.A(new_n14250_), .B(new_n13481_), .Y(new_n14251_));
  AOI21  g13249(.A0(new_n14245_), .A1(new_n13692_), .B0(new_n14251_), .Y(new_n14252_));
  NOR2   g13250(.A(new_n13479_), .B(new_n13432_), .Y(new_n14253_));
  NAND2  g13251(.A(new_n13479_), .B(new_n13432_), .Y(new_n14254_));
  OAI21  g13252(.A0(new_n14253_), .A1(new_n13542_), .B0(new_n14254_), .Y(new_n14255_));
  NOR2   g13253(.A(new_n13477_), .B(new_n13456_), .Y(new_n14256_));
  AOI22  g13254(.A0(new_n13476_), .A1(new_n13469_), .B0(new_n13455_), .B1(new_n13450_), .Y(new_n14257_));
  AOI21  g13255(.A0(new_n13444_), .A1(new_n13439_), .B0(new_n14257_), .Y(new_n14258_));
  AOI21  g13256(.A0(new_n13453_), .A1(new_n13452_), .B0(new_n13454_), .Y(new_n14259_));
  AOI21  g13257(.A0(new_n13470_), .A1(new_n13442_), .B0(new_n13462_), .Y(new_n14260_));
  NOR2   g13258(.A(new_n13463_), .B(new_n11270_), .Y(new_n14261_));
  NOR2   g13259(.A(new_n11273_), .B(new_n13433_), .Y(new_n14262_));
  NOR2   g13260(.A(new_n14262_), .B(new_n14261_), .Y(new_n14263_));
  AOI21  g13261(.A0(new_n13474_), .A1(new_n14263_), .B0(new_n14260_), .Y(new_n14264_));
  NOR2   g13262(.A(new_n13474_), .B(new_n14263_), .Y(new_n14265_));
  NOR3   g13263(.A(new_n14265_), .B(new_n14264_), .C(new_n14259_), .Y(new_n14266_));
  OAI22  g13264(.A0(new_n13467_), .A1(new_n13464_), .B0(new_n13462_), .B1(new_n13459_), .Y(new_n14267_));
  NAND2  g13265(.A(new_n13467_), .B(new_n13464_), .Y(new_n14268_));
  AOI21  g13266(.A0(new_n14268_), .A1(new_n14267_), .B0(new_n13450_), .Y(new_n14269_));
  NOR2   g13267(.A(new_n14269_), .B(new_n14266_), .Y(new_n14270_));
  OAI21  g13268(.A0(new_n14258_), .A1(new_n14256_), .B0(new_n14270_), .Y(new_n14271_));
  OAI21  g13269(.A0(new_n11248_), .A1(new_n11244_), .B0(new_n11283_), .Y(new_n14272_));
  AOI22  g13270(.A0(new_n13443_), .A1(new_n13440_), .B0(new_n14272_), .B1(new_n13538_), .Y(new_n14273_));
  NAND4  g13271(.A(new_n13476_), .B(new_n13469_), .C(new_n13455_), .D(new_n13450_), .Y(new_n14274_));
  OAI221 g13272(.A0(new_n14269_), .A1(new_n14266_), .C0(new_n14274_), .B0(new_n14257_), .B1(new_n14273_), .Y(new_n14275_));
  NAND2  g13273(.A(new_n14275_), .B(new_n14271_), .Y(new_n14276_));
  AOI22  g13274(.A0(new_n13430_), .A1(new_n13414_), .B0(new_n13395_), .B1(new_n13394_), .Y(new_n14277_));
  NOR2   g13275(.A(new_n13410_), .B(new_n13404_), .Y(new_n14278_));
  NOR2   g13276(.A(new_n13409_), .B(new_n13406_), .Y(new_n14279_));
  NAND4  g13277(.A(new_n11357_), .B(new_n11353_), .C(new_n11343_), .D(new_n11339_), .Y(new_n14280_));
  NOR3   g13278(.A(new_n11331_), .B(new_n11330_), .C(new_n6023_), .Y(new_n14281_));
  OAI21  g13279(.A0(new_n11330_), .A1(new_n6023_), .B0(new_n11331_), .Y(new_n14282_));
  OAI211 g13280(.A0(new_n14281_), .A1(new_n11334_), .B0(new_n14282_), .B1(new_n13406_), .Y(new_n14283_));
  NAND2  g13281(.A(new_n14283_), .B(new_n14280_), .Y(new_n14284_));
  AOI211 g13282(.A0(new_n13402_), .A1(new_n11329_), .B(new_n14284_), .C(new_n14279_), .Y(new_n14285_));
  NOR2   g13283(.A(new_n13426_), .B(new_n13419_), .Y(new_n14286_));
  NAND3  g13284(.A(new_n11312_), .B(new_n11310_), .C(new_n5673_), .Y(new_n14287_));
  AOI21  g13285(.A0(new_n11310_), .A1(new_n5673_), .B0(new_n11312_), .Y(new_n14288_));
  AOI21  g13286(.A0(new_n14287_), .A1(new_n11313_), .B0(new_n14288_), .Y(new_n14289_));
  NOR3   g13287(.A(new_n11292_), .B(new_n11291_), .C(new_n11289_), .Y(new_n14290_));
  OAI21  g13288(.A0(new_n11291_), .A1(new_n11289_), .B0(new_n11292_), .Y(new_n14291_));
  OAI21  g13289(.A0(new_n14290_), .A1(new_n11293_), .B0(new_n14291_), .Y(new_n14292_));
  OAI22  g13290(.A0(new_n11323_), .A1(new_n11322_), .B0(new_n11321_), .B1(new_n11320_), .Y(new_n14293_));
  NAND4  g13291(.A(new_n11317_), .B(new_n11314_), .C(new_n11310_), .D(new_n5673_), .Y(new_n14294_));
  NAND4  g13292(.A(new_n14294_), .B(new_n14293_), .C(new_n11308_), .D(new_n11302_), .Y(new_n14295_));
  OAI21  g13293(.A0(new_n14292_), .A1(new_n14289_), .B0(new_n14295_), .Y(new_n14296_));
  AOI221 g13294(.A0(new_n14292_), .A1(new_n14289_), .C0(new_n14296_), .B0(new_n13417_), .B1(new_n11288_), .Y(new_n14297_));
  NOR4   g13295(.A(new_n14297_), .B(new_n14286_), .C(new_n14285_), .D(new_n14278_), .Y(new_n14298_));
  AOI211 g13296(.A0(new_n13407_), .A1(new_n11337_), .B(new_n13408_), .C(new_n13406_), .Y(new_n14299_));
  OAI21  g13297(.A0(new_n14281_), .A1(new_n11334_), .B0(new_n14282_), .Y(new_n14300_));
  NAND2  g13298(.A(new_n14300_), .B(new_n13406_), .Y(new_n14301_));
  OAI21  g13299(.A0(new_n14299_), .A1(new_n13404_), .B0(new_n14301_), .Y(new_n14302_));
  NOR2   g13300(.A(new_n14292_), .B(new_n13422_), .Y(new_n14303_));
  NAND2  g13301(.A(new_n14292_), .B(new_n13422_), .Y(new_n14304_));
  OAI21  g13302(.A0(new_n14303_), .A1(new_n13419_), .B0(new_n14304_), .Y(new_n14305_));
  XOR2   g13303(.A(new_n14305_), .B(new_n14302_), .Y(new_n14306_));
  OAI21  g13304(.A0(new_n14298_), .A1(new_n14277_), .B0(new_n14306_), .Y(new_n14307_));
  NAND2  g13305(.A(new_n14280_), .B(new_n13411_), .Y(new_n14308_));
  XOR2   g13306(.A(new_n14300_), .B(new_n13406_), .Y(new_n14309_));
  NAND2  g13307(.A(new_n14309_), .B(new_n14308_), .Y(new_n14310_));
  NAND2  g13308(.A(new_n14295_), .B(new_n13427_), .Y(new_n14311_));
  XOR2   g13309(.A(new_n14292_), .B(new_n13422_), .Y(new_n14312_));
  NAND2  g13310(.A(new_n14312_), .B(new_n14311_), .Y(new_n14313_));
  AOI22  g13311(.A0(new_n13429_), .A1(new_n14313_), .B0(new_n13413_), .B1(new_n14310_), .Y(new_n14314_));
  NOR2   g13312(.A(new_n14303_), .B(new_n13419_), .Y(new_n14315_));
  AOI21  g13313(.A0(new_n14292_), .A1(new_n13422_), .B0(new_n14315_), .Y(new_n14316_));
  AOI21  g13314(.A0(new_n14316_), .A1(new_n14302_), .B0(new_n14298_), .Y(new_n14317_));
  OAI221 g13315(.A0(new_n14316_), .A1(new_n14302_), .C0(new_n14317_), .B0(new_n14314_), .B1(new_n13548_), .Y(new_n14318_));
  NAND2  g13316(.A(new_n14318_), .B(new_n14307_), .Y(new_n14319_));
  XOR2   g13317(.A(new_n14319_), .B(new_n14276_), .Y(new_n14320_));
  NAND2  g13318(.A(new_n14320_), .B(new_n14255_), .Y(new_n14321_));
  XOR2   g13319(.A(new_n13478_), .B(new_n14273_), .Y(new_n14322_));
  NAND2  g13320(.A(new_n14322_), .B(new_n13549_), .Y(new_n14323_));
  NOR2   g13321(.A(new_n14322_), .B(new_n13549_), .Y(new_n14324_));
  AOI21  g13322(.A0(new_n14323_), .A1(new_n13391_), .B0(new_n14324_), .Y(new_n14325_));
  OAI21  g13323(.A0(new_n14257_), .A1(new_n14273_), .B0(new_n14274_), .Y(new_n14326_));
  NOR3   g13324(.A(new_n14270_), .B(new_n14258_), .C(new_n14256_), .Y(new_n14327_));
  AOI21  g13325(.A0(new_n14270_), .A1(new_n14326_), .B0(new_n14327_), .Y(new_n14328_));
  XOR2   g13326(.A(new_n14319_), .B(new_n14328_), .Y(new_n14329_));
  NAND2  g13327(.A(new_n14329_), .B(new_n14325_), .Y(new_n14330_));
  NOR4   g13328(.A(new_n11425_), .B(new_n11422_), .C(new_n11420_), .D(new_n11419_), .Y(new_n14331_));
  OAI21  g13329(.A0(new_n14331_), .A1(new_n13495_), .B0(new_n11417_), .Y(new_n14332_));
  NAND2  g13330(.A(new_n14332_), .B(new_n13488_), .Y(new_n14333_));
  AOI22  g13331(.A0(new_n13516_), .A1(new_n13512_), .B0(new_n13506_), .B1(new_n14333_), .Y(new_n14334_));
  NOR2   g13332(.A(new_n13517_), .B(new_n13493_), .Y(new_n14335_));
  NOR2   g13333(.A(new_n14335_), .B(new_n14334_), .Y(new_n14336_));
  NOR2   g13334(.A(new_n13535_), .B(new_n14336_), .Y(new_n14337_));
  NOR2   g13335(.A(new_n14337_), .B(new_n14248_), .Y(new_n14338_));
  OAI22  g13336(.A0(new_n13534_), .A1(new_n13531_), .B0(new_n14335_), .B1(new_n14334_), .Y(new_n14339_));
  NOR4   g13337(.A(new_n13534_), .B(new_n13531_), .C(new_n14335_), .D(new_n14334_), .Y(new_n14340_));
  AOI21  g13338(.A0(new_n14339_), .A1(new_n13492_), .B0(new_n14340_), .Y(new_n14341_));
  OAI22  g13339(.A0(new_n13503_), .A1(new_n13499_), .B0(new_n13497_), .B1(new_n13493_), .Y(new_n14342_));
  NAND2  g13340(.A(new_n13503_), .B(new_n13499_), .Y(new_n14343_));
  NAND2  g13341(.A(new_n14343_), .B(new_n14342_), .Y(new_n14344_));
  NOR3   g13342(.A(new_n11392_), .B(new_n11397_), .C(new_n11396_), .Y(new_n14345_));
  OAI21  g13343(.A0(new_n11397_), .A1(new_n11396_), .B0(new_n11392_), .Y(new_n14346_));
  OAI21  g13344(.A0(new_n14345_), .A1(new_n11393_), .B0(new_n14346_), .Y(new_n14347_));
  NOR2   g13345(.A(new_n13529_), .B(new_n14347_), .Y(new_n14348_));
  NAND2  g13346(.A(new_n13529_), .B(new_n14347_), .Y(new_n14349_));
  OAI21  g13347(.A0(new_n14348_), .A1(new_n13523_), .B0(new_n14349_), .Y(new_n14350_));
  INV    g13348(.A(new_n14350_), .Y(new_n14351_));
  XOR2   g13349(.A(new_n14351_), .B(new_n14344_), .Y(new_n14352_));
  AOI21  g13350(.A0(new_n14351_), .A1(new_n14344_), .B0(new_n14340_), .Y(new_n14353_));
  OAI21  g13351(.A0(new_n14351_), .A1(new_n14344_), .B0(new_n14353_), .Y(new_n14354_));
  OAI22  g13352(.A0(new_n14354_), .A1(new_n14338_), .B0(new_n14352_), .B1(new_n14341_), .Y(new_n14355_));
  NAND3  g13353(.A(new_n14355_), .B(new_n14330_), .C(new_n14321_), .Y(new_n14356_));
  NOR2   g13354(.A(new_n14352_), .B(new_n14341_), .Y(new_n14357_));
  NOR2   g13355(.A(new_n14354_), .B(new_n14338_), .Y(new_n14358_));
  NOR2   g13356(.A(new_n14358_), .B(new_n14357_), .Y(new_n14359_));
  XOR2   g13357(.A(new_n14329_), .B(new_n14255_), .Y(new_n14360_));
  NAND2  g13358(.A(new_n14360_), .B(new_n14359_), .Y(new_n14361_));
  AOI21  g13359(.A0(new_n14361_), .A1(new_n14356_), .B0(new_n14252_), .Y(new_n14362_));
  NAND2  g13360(.A(new_n11593_), .B(new_n11560_), .Y(new_n14363_));
  NOR2   g13361(.A(new_n11593_), .B(new_n11560_), .Y(new_n14364_));
  AOI21  g13362(.A0(new_n14363_), .A1(new_n11524_), .B0(new_n14364_), .Y(new_n14365_));
  XOR2   g13363(.A(new_n13621_), .B(new_n14365_), .Y(new_n14366_));
  NAND2  g13364(.A(new_n11521_), .B(new_n11486_), .Y(new_n14367_));
  NOR2   g13365(.A(new_n11521_), .B(new_n11486_), .Y(new_n14368_));
  AOI21  g13366(.A0(new_n14367_), .A1(new_n11446_), .B0(new_n14368_), .Y(new_n14369_));
  XOR2   g13367(.A(new_n13687_), .B(new_n14369_), .Y(new_n14370_));
  NAND2  g13368(.A(new_n14370_), .B(new_n14366_), .Y(new_n14371_));
  NOR2   g13369(.A(new_n14370_), .B(new_n14366_), .Y(new_n14372_));
  AOI21  g13370(.A0(new_n14371_), .A1(new_n13557_), .B0(new_n14372_), .Y(new_n14373_));
  NOR2   g13371(.A(new_n13648_), .B(new_n13641_), .Y(new_n14374_));
  AOI211 g13372(.A0(new_n13639_), .A1(new_n11487_), .B(new_n13658_), .C(new_n13650_), .Y(new_n14375_));
  NOR2   g13373(.A(new_n13673_), .B(new_n13666_), .Y(new_n14376_));
  AOI211 g13374(.A0(new_n13664_), .A1(new_n11450_), .B(new_n13683_), .C(new_n13675_), .Y(new_n14377_));
  OAI22  g13375(.A0(new_n14377_), .A1(new_n14376_), .B0(new_n14375_), .B1(new_n14374_), .Y(new_n14378_));
  NOR4   g13376(.A(new_n14377_), .B(new_n14376_), .C(new_n14375_), .D(new_n14374_), .Y(new_n14379_));
  AOI21  g13377(.A0(new_n14378_), .A1(new_n13636_), .B0(new_n14379_), .Y(new_n14380_));
  NOR2   g13378(.A(new_n13657_), .B(new_n13644_), .Y(new_n14381_));
  NAND2  g13379(.A(new_n13657_), .B(new_n13644_), .Y(new_n14382_));
  OAI21  g13380(.A0(new_n14381_), .A1(new_n13641_), .B0(new_n14382_), .Y(new_n14383_));
  NOR2   g13381(.A(new_n13682_), .B(new_n13669_), .Y(new_n14384_));
  NAND2  g13382(.A(new_n13682_), .B(new_n13669_), .Y(new_n14385_));
  OAI21  g13383(.A0(new_n14384_), .A1(new_n13666_), .B0(new_n14385_), .Y(new_n14386_));
  XOR2   g13384(.A(new_n14386_), .B(new_n14383_), .Y(new_n14387_));
  INV    g13385(.A(new_n14387_), .Y(new_n14388_));
  NAND2  g13386(.A(new_n13651_), .B(new_n13649_), .Y(new_n14389_));
  INV    g13387(.A(new_n13648_), .Y(new_n14390_));
  NAND2  g13388(.A(new_n14390_), .B(new_n14389_), .Y(new_n14391_));
  NAND2  g13389(.A(new_n13676_), .B(new_n13674_), .Y(new_n14392_));
  INV    g13390(.A(new_n13673_), .Y(new_n14393_));
  NAND2  g13391(.A(new_n14393_), .B(new_n14392_), .Y(new_n14394_));
  AOI22  g13392(.A0(new_n13685_), .A1(new_n14394_), .B0(new_n13660_), .B1(new_n14391_), .Y(new_n14395_));
  NOR2   g13393(.A(new_n14384_), .B(new_n13666_), .Y(new_n14396_));
  AOI21  g13394(.A0(new_n13682_), .A1(new_n13669_), .B0(new_n14396_), .Y(new_n14397_));
  AOI21  g13395(.A0(new_n14397_), .A1(new_n14383_), .B0(new_n14379_), .Y(new_n14398_));
  OAI221 g13396(.A0(new_n14397_), .A1(new_n14383_), .C0(new_n14398_), .B0(new_n14395_), .B1(new_n14369_), .Y(new_n14399_));
  OAI21  g13397(.A0(new_n14388_), .A1(new_n14380_), .B0(new_n14399_), .Y(new_n14400_));
  OAI22  g13398(.A0(new_n11590_), .A1(new_n11586_), .B0(new_n13574_), .B1(new_n13573_), .Y(new_n14401_));
  AOI21  g13399(.A0(new_n14401_), .A1(new_n11561_), .B0(new_n13575_), .Y(new_n14402_));
  NAND2  g13400(.A(new_n13586_), .B(new_n13583_), .Y(new_n14403_));
  AOI21  g13401(.A0(new_n13589_), .A1(new_n14403_), .B0(new_n14402_), .Y(new_n14404_));
  NOR4   g13402(.A(new_n13587_), .B(new_n13580_), .C(new_n13575_), .D(new_n13571_), .Y(new_n14405_));
  AOI21  g13403(.A0(new_n13616_), .A1(new_n11526_), .B0(new_n13601_), .Y(new_n14406_));
  OAI221 g13404(.A0(new_n13605_), .A1(new_n11538_), .C0(new_n13610_), .B0(new_n11532_), .B1(new_n13598_), .Y(new_n14407_));
  NAND2  g13405(.A(new_n13606_), .B(new_n13604_), .Y(new_n14408_));
  AOI21  g13406(.A0(new_n14408_), .A1(new_n14407_), .B0(new_n14406_), .Y(new_n14409_));
  NOR4   g13407(.A(new_n13614_), .B(new_n13607_), .C(new_n13601_), .D(new_n13597_), .Y(new_n14410_));
  OAI22  g13408(.A0(new_n14410_), .A1(new_n14409_), .B0(new_n14405_), .B1(new_n14404_), .Y(new_n14411_));
  NOR4   g13409(.A(new_n14410_), .B(new_n14409_), .C(new_n14405_), .D(new_n14404_), .Y(new_n14412_));
  AOI21  g13410(.A0(new_n14411_), .A1(new_n13565_), .B0(new_n14412_), .Y(new_n14413_));
  AOI221 g13411(.A0(new_n13576_), .A1(new_n11581_), .C0(new_n13579_), .B0(new_n11583_), .B1(new_n13567_), .Y(new_n14414_));
  NAND2  g13412(.A(new_n13579_), .B(new_n13583_), .Y(new_n14415_));
  OAI21  g13413(.A0(new_n14414_), .A1(new_n14402_), .B0(new_n14415_), .Y(new_n14416_));
  NOR2   g13414(.A(new_n13606_), .B(new_n13610_), .Y(new_n14417_));
  NAND2  g13415(.A(new_n13606_), .B(new_n13610_), .Y(new_n14418_));
  OAI21  g13416(.A0(new_n14417_), .A1(new_n14406_), .B0(new_n14418_), .Y(new_n14419_));
  XOR2   g13417(.A(new_n14419_), .B(new_n14416_), .Y(new_n14420_));
  INV    g13418(.A(new_n14420_), .Y(new_n14421_));
  AOI22  g13419(.A0(new_n13619_), .A1(new_n13615_), .B0(new_n13591_), .B1(new_n13588_), .Y(new_n14422_));
  NOR2   g13420(.A(new_n14417_), .B(new_n14406_), .Y(new_n14423_));
  AOI21  g13421(.A0(new_n13606_), .A1(new_n13610_), .B0(new_n14423_), .Y(new_n14424_));
  AOI21  g13422(.A0(new_n14424_), .A1(new_n14416_), .B0(new_n14412_), .Y(new_n14425_));
  OAI221 g13423(.A0(new_n14424_), .A1(new_n14416_), .C0(new_n14425_), .B0(new_n14422_), .B1(new_n14365_), .Y(new_n14426_));
  OAI21  g13424(.A0(new_n14421_), .A1(new_n14413_), .B0(new_n14426_), .Y(new_n14427_));
  XOR2   g13425(.A(new_n14427_), .B(new_n14400_), .Y(new_n14428_));
  XOR2   g13426(.A(new_n14428_), .B(new_n14373_), .Y(new_n14429_));
  NOR2   g13427(.A(new_n14249_), .B(new_n13482_), .Y(new_n14430_));
  OAI22  g13428(.A0(new_n14250_), .A1(new_n13481_), .B0(new_n14430_), .B1(new_n13388_), .Y(new_n14431_));
  NOR2   g13429(.A(new_n14329_), .B(new_n14325_), .Y(new_n14432_));
  OAI21  g13430(.A0(new_n14320_), .A1(new_n14255_), .B0(new_n14355_), .Y(new_n14433_));
  XOR2   g13431(.A(new_n14320_), .B(new_n14255_), .Y(new_n14434_));
  OAI22  g13432(.A0(new_n14434_), .A1(new_n14355_), .B0(new_n14433_), .B1(new_n14432_), .Y(new_n14435_));
  OAI21  g13433(.A0(new_n14435_), .A1(new_n14431_), .B0(new_n14429_), .Y(new_n14436_));
  XOR2   g13434(.A(new_n14435_), .B(new_n14431_), .Y(new_n14437_));
  OAI22  g13435(.A0(new_n14437_), .A1(new_n14429_), .B0(new_n14436_), .B1(new_n14362_), .Y(new_n14438_));
  XOR2   g13436(.A(new_n14438_), .B(new_n14243_), .Y(new_n14439_));
  NOR2   g13437(.A(new_n11916_), .B(new_n11766_), .Y(new_n14440_));
  NAND2  g13438(.A(new_n11916_), .B(new_n11766_), .Y(new_n14441_));
  OAI21  g13439(.A0(new_n14440_), .A1(new_n11610_), .B0(new_n14441_), .Y(new_n14442_));
  XOR2   g13440(.A(new_n13374_), .B(new_n14442_), .Y(new_n14443_));
  NAND2  g13441(.A(new_n14443_), .B(new_n13131_), .Y(new_n14444_));
  NOR2   g13442(.A(new_n14443_), .B(new_n13131_), .Y(new_n14445_));
  AOI21  g13443(.A0(new_n14444_), .A1(new_n13706_), .B0(new_n14445_), .Y(new_n14446_));
  NOR2   g13444(.A(new_n11764_), .B(new_n11691_), .Y(new_n14447_));
  NAND2  g13445(.A(new_n11764_), .B(new_n11691_), .Y(new_n14448_));
  OAI21  g13446(.A0(new_n14447_), .A1(new_n13133_), .B0(new_n14448_), .Y(new_n14449_));
  XOR2   g13447(.A(new_n13372_), .B(new_n14449_), .Y(new_n14450_));
  NOR2   g13448(.A(new_n14450_), .B(new_n13246_), .Y(new_n14451_));
  NAND2  g13449(.A(new_n14450_), .B(new_n13246_), .Y(new_n14452_));
  OAI21  g13450(.A0(new_n14451_), .A1(new_n13139_), .B0(new_n14452_), .Y(new_n14453_));
  NOR2   g13451(.A(new_n13371_), .B(new_n13321_), .Y(new_n14454_));
  NAND2  g13452(.A(new_n13371_), .B(new_n13321_), .Y(new_n14455_));
  OAI21  g13453(.A0(new_n14454_), .A1(new_n13255_), .B0(new_n14455_), .Y(new_n14456_));
  AOI22  g13454(.A0(new_n13369_), .A1(new_n13353_), .B0(new_n13332_), .B1(new_n13331_), .Y(new_n14457_));
  NOR2   g13455(.A(new_n13346_), .B(new_n13338_), .Y(new_n14458_));
  NAND2  g13456(.A(new_n13350_), .B(new_n13348_), .Y(new_n14459_));
  AOI221 g13457(.A0(new_n13345_), .A1(new_n13342_), .C0(new_n14459_), .B0(new_n13336_), .B1(new_n11652_), .Y(new_n14460_));
  NOR2   g13458(.A(new_n13365_), .B(new_n13358_), .Y(new_n14461_));
  NAND3  g13459(.A(new_n11636_), .B(new_n11635_), .C(new_n9074_), .Y(new_n14462_));
  AOI21  g13460(.A0(new_n11635_), .A1(new_n9074_), .B0(new_n11636_), .Y(new_n14463_));
  AOI21  g13461(.A0(new_n14462_), .A1(new_n11637_), .B0(new_n14463_), .Y(new_n14464_));
  NOR3   g13462(.A(new_n11617_), .B(new_n11616_), .C(new_n11614_), .Y(new_n14465_));
  OAI21  g13463(.A0(new_n11616_), .A1(new_n11614_), .B0(new_n11617_), .Y(new_n14466_));
  OAI21  g13464(.A0(new_n14465_), .A1(new_n11618_), .B0(new_n14466_), .Y(new_n14467_));
  OAI22  g13465(.A0(new_n11646_), .A1(new_n11645_), .B0(new_n11644_), .B1(new_n11643_), .Y(new_n14468_));
  NAND4  g13466(.A(new_n11641_), .B(new_n11638_), .C(new_n11635_), .D(new_n9074_), .Y(new_n14469_));
  NAND4  g13467(.A(new_n14469_), .B(new_n14468_), .C(new_n11633_), .D(new_n11627_), .Y(new_n14470_));
  OAI21  g13468(.A0(new_n14467_), .A1(new_n14464_), .B0(new_n14470_), .Y(new_n14471_));
  AOI221 g13469(.A0(new_n14467_), .A1(new_n14464_), .C0(new_n14471_), .B0(new_n13356_), .B1(new_n11613_), .Y(new_n14472_));
  NOR4   g13470(.A(new_n14472_), .B(new_n14461_), .C(new_n14460_), .D(new_n14458_), .Y(new_n14473_));
  NOR2   g13471(.A(new_n13345_), .B(new_n13349_), .Y(new_n14474_));
  NAND2  g13472(.A(new_n13345_), .B(new_n13349_), .Y(new_n14475_));
  OAI21  g13473(.A0(new_n14474_), .A1(new_n13338_), .B0(new_n14475_), .Y(new_n14476_));
  NOR2   g13474(.A(new_n14467_), .B(new_n13361_), .Y(new_n14477_));
  NAND2  g13475(.A(new_n14467_), .B(new_n13361_), .Y(new_n14478_));
  OAI21  g13476(.A0(new_n14477_), .A1(new_n13358_), .B0(new_n14478_), .Y(new_n14479_));
  XOR2   g13477(.A(new_n14479_), .B(new_n14476_), .Y(new_n14480_));
  OAI21  g13478(.A0(new_n14473_), .A1(new_n14457_), .B0(new_n14480_), .Y(new_n14481_));
  NAND2  g13479(.A(new_n11689_), .B(new_n11650_), .Y(new_n14482_));
  NOR2   g13480(.A(new_n11689_), .B(new_n11650_), .Y(new_n14483_));
  AOI21  g13481(.A0(new_n14482_), .A1(new_n11612_), .B0(new_n14483_), .Y(new_n14484_));
  NAND2  g13482(.A(new_n13348_), .B(new_n13347_), .Y(new_n14485_));
  XOR2   g13483(.A(new_n13345_), .B(new_n13349_), .Y(new_n14486_));
  NAND2  g13484(.A(new_n14486_), .B(new_n14485_), .Y(new_n14487_));
  NAND2  g13485(.A(new_n14470_), .B(new_n13366_), .Y(new_n14488_));
  XOR2   g13486(.A(new_n14467_), .B(new_n13361_), .Y(new_n14489_));
  NAND2  g13487(.A(new_n14489_), .B(new_n14488_), .Y(new_n14490_));
  AOI22  g13488(.A0(new_n13368_), .A1(new_n14490_), .B0(new_n13352_), .B1(new_n14487_), .Y(new_n14491_));
  NOR2   g13489(.A(new_n14477_), .B(new_n13358_), .Y(new_n14492_));
  AOI21  g13490(.A0(new_n14467_), .A1(new_n13361_), .B0(new_n14492_), .Y(new_n14493_));
  AOI21  g13491(.A0(new_n14493_), .A1(new_n14476_), .B0(new_n14473_), .Y(new_n14494_));
  OAI221 g13492(.A0(new_n14493_), .A1(new_n14476_), .C0(new_n14494_), .B0(new_n14491_), .B1(new_n14484_), .Y(new_n14495_));
  NAND2  g13493(.A(new_n14495_), .B(new_n14481_), .Y(new_n14496_));
  AOI22  g13494(.A0(new_n13318_), .A1(new_n13309_), .B0(new_n13294_), .B1(new_n13285_), .Y(new_n14497_));
  AOI21  g13495(.A0(new_n13271_), .A1(new_n13270_), .B0(new_n14497_), .Y(new_n14498_));
  AOI21  g13496(.A0(new_n13286_), .A1(new_n11729_), .B0(new_n13278_), .Y(new_n14499_));
  AOI21  g13497(.A0(new_n13293_), .A1(new_n13289_), .B0(new_n14499_), .Y(new_n14500_));
  NAND2  g13498(.A(new_n13289_), .B(new_n13288_), .Y(new_n14501_));
  AOI211 g13499(.A0(new_n13283_), .A1(new_n13292_), .B(new_n14501_), .C(new_n13275_), .Y(new_n14502_));
  AOI21  g13500(.A0(new_n13310_), .A1(new_n11694_), .B0(new_n13302_), .Y(new_n14503_));
  AOI21  g13501(.A0(new_n13317_), .A1(new_n13313_), .B0(new_n14503_), .Y(new_n14504_));
  NAND2  g13502(.A(new_n13313_), .B(new_n13312_), .Y(new_n14505_));
  AOI211 g13503(.A0(new_n13307_), .A1(new_n13316_), .B(new_n14505_), .C(new_n13299_), .Y(new_n14506_));
  NOR4   g13504(.A(new_n14506_), .B(new_n14504_), .C(new_n14502_), .D(new_n14500_), .Y(new_n14507_));
  NOR2   g13505(.A(new_n13283_), .B(new_n13280_), .Y(new_n14508_));
  NAND2  g13506(.A(new_n13283_), .B(new_n13280_), .Y(new_n14509_));
  OAI21  g13507(.A0(new_n14508_), .A1(new_n14499_), .B0(new_n14509_), .Y(new_n14510_));
  NOR2   g13508(.A(new_n13307_), .B(new_n13304_), .Y(new_n14511_));
  NAND2  g13509(.A(new_n13307_), .B(new_n13304_), .Y(new_n14512_));
  OAI21  g13510(.A0(new_n14511_), .A1(new_n14503_), .B0(new_n14512_), .Y(new_n14513_));
  XOR2   g13511(.A(new_n14513_), .B(new_n14510_), .Y(new_n14514_));
  OAI21  g13512(.A0(new_n14507_), .A1(new_n14498_), .B0(new_n14514_), .Y(new_n14515_));
  NAND2  g13513(.A(new_n11762_), .B(new_n11727_), .Y(new_n14516_));
  NOR2   g13514(.A(new_n11762_), .B(new_n11727_), .Y(new_n14517_));
  AOI21  g13515(.A0(new_n14516_), .A1(new_n11692_), .B0(new_n14517_), .Y(new_n14518_));
  NOR2   g13516(.A(new_n14511_), .B(new_n14503_), .Y(new_n14519_));
  AOI21  g13517(.A0(new_n13307_), .A1(new_n13304_), .B0(new_n14519_), .Y(new_n14520_));
  AOI21  g13518(.A0(new_n14520_), .A1(new_n14510_), .B0(new_n14507_), .Y(new_n14521_));
  OAI221 g13519(.A0(new_n14520_), .A1(new_n14510_), .C0(new_n14521_), .B0(new_n14497_), .B1(new_n14518_), .Y(new_n14522_));
  NAND2  g13520(.A(new_n14522_), .B(new_n14515_), .Y(new_n14523_));
  XOR2   g13521(.A(new_n14523_), .B(new_n14496_), .Y(new_n14524_));
  XOR2   g13522(.A(new_n14524_), .B(new_n14456_), .Y(new_n14525_));
  AOI22  g13523(.A0(new_n7543_), .A1(new_n7277_), .B0(new_n7521_), .B1(new_n7515_), .Y(new_n14526_));
  NOR2   g13524(.A(new_n14526_), .B(new_n8064_), .Y(new_n14527_));
  XOR2   g13525(.A(new_n11840_), .B(new_n14527_), .Y(new_n14528_));
  OAI21  g13526(.A0(new_n8055_), .A1(new_n8040_), .B0(new_n8043_), .Y(new_n14529_));
  XOR2   g13527(.A(new_n11913_), .B(new_n14529_), .Y(new_n14530_));
  NAND2  g13528(.A(new_n14530_), .B(new_n14528_), .Y(new_n14531_));
  NOR2   g13529(.A(new_n14530_), .B(new_n14528_), .Y(new_n14532_));
  AOI21  g13530(.A0(new_n14531_), .A1(new_n11767_), .B0(new_n14532_), .Y(new_n14533_));
  NOR2   g13531(.A(new_n13244_), .B(new_n13200_), .Y(new_n14534_));
  NAND2  g13532(.A(new_n13244_), .B(new_n13200_), .Y(new_n14535_));
  OAI21  g13533(.A0(new_n14534_), .A1(new_n14533_), .B0(new_n14535_), .Y(new_n14536_));
  AOI21  g13534(.A0(new_n7540_), .A1(new_n7518_), .B0(new_n7520_), .Y(new_n14537_));
  XOR2   g13535(.A(new_n11805_), .B(new_n14537_), .Y(new_n14538_));
  OAI22  g13536(.A0(new_n11835_), .A1(new_n11834_), .B0(new_n11833_), .B1(new_n7286_), .Y(new_n14539_));
  NAND2  g13537(.A(new_n7253_), .B(new_n7189_), .Y(new_n14540_));
  NAND4  g13538(.A(new_n11831_), .B(new_n11828_), .C(new_n14540_), .D(new_n7256_), .Y(new_n14541_));
  NAND2  g13539(.A(new_n14541_), .B(new_n14539_), .Y(new_n14542_));
  XOR2   g13540(.A(new_n14542_), .B(new_n11823_), .Y(new_n14543_));
  XOR2   g13541(.A(new_n14543_), .B(new_n11808_), .Y(new_n14544_));
  OAI22  g13542(.A0(new_n14544_), .A1(new_n14538_), .B0(new_n14526_), .B1(new_n8064_), .Y(new_n14545_));
  NAND2  g13543(.A(new_n14544_), .B(new_n14538_), .Y(new_n14546_));
  NAND2  g13544(.A(new_n13221_), .B(new_n11769_), .Y(new_n14547_));
  AOI21  g13545(.A0(new_n13229_), .A1(new_n13226_), .B0(new_n13222_), .Y(new_n14548_));
  OAI211 g13546(.A0(new_n13229_), .A1(new_n13226_), .B0(new_n14548_), .B1(new_n14547_), .Y(new_n14549_));
  OAI21  g13547(.A0(new_n13230_), .A1(new_n13223_), .B0(new_n14549_), .Y(new_n14550_));
  AOI22  g13548(.A0(new_n14550_), .A1(new_n13218_), .B0(new_n14546_), .B1(new_n14545_), .Y(new_n14551_));
  NOR2   g13549(.A(new_n13214_), .B(new_n13208_), .Y(new_n14552_));
  NOR2   g13550(.A(new_n13213_), .B(new_n13210_), .Y(new_n14553_));
  NAND4  g13551(.A(new_n14541_), .B(new_n14539_), .C(new_n11822_), .D(new_n11818_), .Y(new_n14554_));
  NOR3   g13552(.A(new_n11810_), .B(new_n11809_), .C(new_n7281_), .Y(new_n14555_));
  OAI21  g13553(.A0(new_n11809_), .A1(new_n7281_), .B0(new_n11810_), .Y(new_n14556_));
  OAI211 g13554(.A0(new_n14555_), .A1(new_n11813_), .B0(new_n14556_), .B1(new_n13210_), .Y(new_n14557_));
  NAND2  g13555(.A(new_n14557_), .B(new_n14554_), .Y(new_n14558_));
  AOI211 g13556(.A0(new_n13206_), .A1(new_n11808_), .B(new_n14558_), .C(new_n14553_), .Y(new_n14559_));
  NOR4   g13557(.A(new_n13241_), .B(new_n13231_), .C(new_n14559_), .D(new_n14552_), .Y(new_n14560_));
  AOI211 g13558(.A0(new_n13211_), .A1(new_n11816_), .B(new_n13212_), .C(new_n13210_), .Y(new_n14561_));
  OAI21  g13559(.A0(new_n14555_), .A1(new_n11813_), .B0(new_n14556_), .Y(new_n14562_));
  NAND2  g13560(.A(new_n14562_), .B(new_n13210_), .Y(new_n14563_));
  OAI21  g13561(.A0(new_n14561_), .A1(new_n13208_), .B0(new_n14563_), .Y(new_n14564_));
  NOR2   g13562(.A(new_n13237_), .B(new_n13226_), .Y(new_n14565_));
  NAND2  g13563(.A(new_n13237_), .B(new_n13226_), .Y(new_n14566_));
  OAI21  g13564(.A0(new_n14565_), .A1(new_n13223_), .B0(new_n14566_), .Y(new_n14567_));
  XOR2   g13565(.A(new_n14567_), .B(new_n14564_), .Y(new_n14568_));
  OAI21  g13566(.A0(new_n14560_), .A1(new_n14551_), .B0(new_n14568_), .Y(new_n14569_));
  NOR2   g13567(.A(new_n14559_), .B(new_n14552_), .Y(new_n14570_));
  NOR2   g13568(.A(new_n13242_), .B(new_n14570_), .Y(new_n14571_));
  NOR2   g13569(.A(new_n14565_), .B(new_n13223_), .Y(new_n14572_));
  AOI21  g13570(.A0(new_n13237_), .A1(new_n13226_), .B0(new_n14572_), .Y(new_n14573_));
  AOI21  g13571(.A0(new_n14573_), .A1(new_n14564_), .B0(new_n14560_), .Y(new_n14574_));
  OAI221 g13572(.A0(new_n14573_), .A1(new_n14564_), .C0(new_n14574_), .B0(new_n14571_), .B1(new_n13203_), .Y(new_n14575_));
  NAND2  g13573(.A(new_n14575_), .B(new_n14569_), .Y(new_n14576_));
  AOI22  g13574(.A0(new_n13197_), .A1(new_n13188_), .B0(new_n13174_), .B1(new_n13167_), .Y(new_n14577_));
  AOI21  g13575(.A0(new_n13150_), .A1(new_n13149_), .B0(new_n14577_), .Y(new_n14578_));
  AOI21  g13576(.A0(new_n13168_), .A1(new_n11880_), .B0(new_n13160_), .Y(new_n14579_));
  XOR2   g13577(.A(new_n13172_), .B(new_n13162_), .Y(new_n14580_));
  NOR2   g13578(.A(new_n14580_), .B(new_n14579_), .Y(new_n14581_));
  NOR2   g13579(.A(new_n13172_), .B(new_n13162_), .Y(new_n14582_));
  NAND4  g13580(.A(new_n11909_), .B(new_n11905_), .C(new_n11895_), .D(new_n11891_), .Y(new_n14583_));
  OAI211 g13581(.A0(new_n13163_), .A1(new_n11886_), .B0(new_n13164_), .B1(new_n13162_), .Y(new_n14584_));
  NAND2  g13582(.A(new_n14584_), .B(new_n14583_), .Y(new_n14585_));
  NOR3   g13583(.A(new_n14585_), .B(new_n14582_), .C(new_n13154_), .Y(new_n14586_));
  AOI21  g13584(.A0(new_n13189_), .A1(new_n11845_), .B0(new_n13181_), .Y(new_n14587_));
  AOI21  g13585(.A0(new_n13196_), .A1(new_n13192_), .B0(new_n14587_), .Y(new_n14588_));
  NAND2  g13586(.A(new_n13192_), .B(new_n13191_), .Y(new_n14589_));
  AOI211 g13587(.A0(new_n13186_), .A1(new_n13195_), .B(new_n14589_), .C(new_n13178_), .Y(new_n14590_));
  NOR4   g13588(.A(new_n14590_), .B(new_n14588_), .C(new_n14586_), .D(new_n14581_), .Y(new_n14591_));
  AOI211 g13589(.A0(new_n13170_), .A1(new_n11889_), .B(new_n13171_), .C(new_n13162_), .Y(new_n14592_));
  NAND2  g13590(.A(new_n13165_), .B(new_n13162_), .Y(new_n14593_));
  OAI21  g13591(.A0(new_n14592_), .A1(new_n14579_), .B0(new_n14593_), .Y(new_n14594_));
  NOR2   g13592(.A(new_n13186_), .B(new_n13183_), .Y(new_n14595_));
  NAND2  g13593(.A(new_n13186_), .B(new_n13183_), .Y(new_n14596_));
  OAI21  g13594(.A0(new_n14595_), .A1(new_n14587_), .B0(new_n14596_), .Y(new_n14597_));
  XOR2   g13595(.A(new_n14597_), .B(new_n14594_), .Y(new_n14598_));
  OAI21  g13596(.A0(new_n14591_), .A1(new_n14578_), .B0(new_n14598_), .Y(new_n14599_));
  NOR2   g13597(.A(new_n13159_), .B(new_n13158_), .Y(new_n14600_));
  XOR2   g13598(.A(new_n14600_), .B(new_n11896_), .Y(new_n14601_));
  XOR2   g13599(.A(new_n14601_), .B(new_n11880_), .Y(new_n14602_));
  NAND2  g13600(.A(new_n14602_), .B(new_n11878_), .Y(new_n14603_));
  NOR2   g13601(.A(new_n14602_), .B(new_n11878_), .Y(new_n14604_));
  AOI21  g13602(.A0(new_n14603_), .A1(new_n14529_), .B0(new_n14604_), .Y(new_n14605_));
  NOR2   g13603(.A(new_n14595_), .B(new_n14587_), .Y(new_n14606_));
  AOI21  g13604(.A0(new_n13186_), .A1(new_n13183_), .B0(new_n14606_), .Y(new_n14607_));
  AOI21  g13605(.A0(new_n14607_), .A1(new_n14594_), .B0(new_n14591_), .Y(new_n14608_));
  OAI221 g13606(.A0(new_n14607_), .A1(new_n14594_), .C0(new_n14608_), .B0(new_n14577_), .B1(new_n14605_), .Y(new_n14609_));
  NAND2  g13607(.A(new_n14609_), .B(new_n14599_), .Y(new_n14610_));
  XOR2   g13608(.A(new_n14610_), .B(new_n14576_), .Y(new_n14611_));
  XOR2   g13609(.A(new_n14611_), .B(new_n14536_), .Y(new_n14612_));
  XOR2   g13610(.A(new_n14612_), .B(new_n14525_), .Y(new_n14613_));
  XOR2   g13611(.A(new_n14613_), .B(new_n14453_), .Y(new_n14614_));
  AOI22  g13612(.A0(new_n10607_), .A1(new_n10341_), .B0(new_n10585_), .B1(new_n10579_), .Y(new_n14615_));
  NOR2   g13613(.A(new_n14615_), .B(new_n11128_), .Y(new_n14616_));
  XOR2   g13614(.A(new_n12149_), .B(new_n14616_), .Y(new_n14617_));
  OAI21  g13615(.A0(new_n11119_), .A1(new_n11104_), .B0(new_n11107_), .Y(new_n14618_));
  XOR2   g13616(.A(new_n12222_), .B(new_n14618_), .Y(new_n14619_));
  NAND2  g13617(.A(new_n14619_), .B(new_n14617_), .Y(new_n14620_));
  NOR2   g13618(.A(new_n14619_), .B(new_n14617_), .Y(new_n14621_));
  AOI21  g13619(.A0(new_n14620_), .A1(new_n12076_), .B0(new_n14621_), .Y(new_n14622_));
  XOR2   g13620(.A(new_n13010_), .B(new_n14622_), .Y(new_n14623_));
  NAND2  g13621(.A(new_n13129_), .B(new_n14623_), .Y(new_n14624_));
  NOR2   g13622(.A(new_n13129_), .B(new_n14623_), .Y(new_n14625_));
  AOI21  g13623(.A0(new_n14624_), .A1(new_n12903_), .B0(new_n14625_), .Y(new_n14626_));
  NOR2   g13624(.A(new_n13127_), .B(new_n13077_), .Y(new_n14627_));
  NAND2  g13625(.A(new_n13127_), .B(new_n13077_), .Y(new_n14628_));
  OAI21  g13626(.A0(new_n14627_), .A1(new_n13019_), .B0(new_n14628_), .Y(new_n14629_));
  AOI22  g13627(.A0(new_n13125_), .A1(new_n13109_), .B0(new_n13088_), .B1(new_n13087_), .Y(new_n14630_));
  NOR2   g13628(.A(new_n13102_), .B(new_n13094_), .Y(new_n14631_));
  NAND2  g13629(.A(new_n13106_), .B(new_n13104_), .Y(new_n14632_));
  AOI221 g13630(.A0(new_n13101_), .A1(new_n13098_), .C0(new_n14632_), .B0(new_n13092_), .B1(new_n11961_), .Y(new_n14633_));
  NOR2   g13631(.A(new_n13121_), .B(new_n13114_), .Y(new_n14634_));
  NAND3  g13632(.A(new_n11945_), .B(new_n11944_), .C(new_n10099_), .Y(new_n14635_));
  AOI21  g13633(.A0(new_n11944_), .A1(new_n10099_), .B0(new_n11945_), .Y(new_n14636_));
  AOI21  g13634(.A0(new_n14635_), .A1(new_n11946_), .B0(new_n14636_), .Y(new_n14637_));
  NOR3   g13635(.A(new_n11926_), .B(new_n11925_), .C(new_n11923_), .Y(new_n14638_));
  OAI21  g13636(.A0(new_n11925_), .A1(new_n11923_), .B0(new_n11926_), .Y(new_n14639_));
  OAI21  g13637(.A0(new_n14638_), .A1(new_n11927_), .B0(new_n14639_), .Y(new_n14640_));
  OAI22  g13638(.A0(new_n11955_), .A1(new_n11954_), .B0(new_n11953_), .B1(new_n11952_), .Y(new_n14641_));
  NAND4  g13639(.A(new_n11950_), .B(new_n11947_), .C(new_n11944_), .D(new_n10099_), .Y(new_n14642_));
  NAND4  g13640(.A(new_n14642_), .B(new_n14641_), .C(new_n11942_), .D(new_n11936_), .Y(new_n14643_));
  OAI21  g13641(.A0(new_n14640_), .A1(new_n14637_), .B0(new_n14643_), .Y(new_n14644_));
  AOI221 g13642(.A0(new_n14640_), .A1(new_n14637_), .C0(new_n14644_), .B0(new_n13112_), .B1(new_n11922_), .Y(new_n14645_));
  NOR4   g13643(.A(new_n14645_), .B(new_n14634_), .C(new_n14633_), .D(new_n14631_), .Y(new_n14646_));
  NOR2   g13644(.A(new_n13101_), .B(new_n13105_), .Y(new_n14647_));
  NAND2  g13645(.A(new_n13101_), .B(new_n13105_), .Y(new_n14648_));
  OAI21  g13646(.A0(new_n14647_), .A1(new_n13094_), .B0(new_n14648_), .Y(new_n14649_));
  NOR2   g13647(.A(new_n14640_), .B(new_n13117_), .Y(new_n14650_));
  NAND2  g13648(.A(new_n14640_), .B(new_n13117_), .Y(new_n14651_));
  OAI21  g13649(.A0(new_n14650_), .A1(new_n13114_), .B0(new_n14651_), .Y(new_n14652_));
  XOR2   g13650(.A(new_n14652_), .B(new_n14649_), .Y(new_n14653_));
  OAI21  g13651(.A0(new_n14646_), .A1(new_n14630_), .B0(new_n14653_), .Y(new_n14654_));
  NAND2  g13652(.A(new_n11998_), .B(new_n11959_), .Y(new_n14655_));
  NOR2   g13653(.A(new_n11998_), .B(new_n11959_), .Y(new_n14656_));
  AOI21  g13654(.A0(new_n14655_), .A1(new_n11921_), .B0(new_n14656_), .Y(new_n14657_));
  NAND2  g13655(.A(new_n13104_), .B(new_n13103_), .Y(new_n14658_));
  XOR2   g13656(.A(new_n13101_), .B(new_n13105_), .Y(new_n14659_));
  NAND2  g13657(.A(new_n14659_), .B(new_n14658_), .Y(new_n14660_));
  NAND2  g13658(.A(new_n14643_), .B(new_n13122_), .Y(new_n14661_));
  XOR2   g13659(.A(new_n14640_), .B(new_n13117_), .Y(new_n14662_));
  NAND2  g13660(.A(new_n14662_), .B(new_n14661_), .Y(new_n14663_));
  AOI22  g13661(.A0(new_n13124_), .A1(new_n14663_), .B0(new_n13108_), .B1(new_n14660_), .Y(new_n14664_));
  NOR2   g13662(.A(new_n14650_), .B(new_n13114_), .Y(new_n14665_));
  AOI21  g13663(.A0(new_n14640_), .A1(new_n13117_), .B0(new_n14665_), .Y(new_n14666_));
  AOI21  g13664(.A0(new_n14666_), .A1(new_n14649_), .B0(new_n14646_), .Y(new_n14667_));
  OAI221 g13665(.A0(new_n14666_), .A1(new_n14649_), .C0(new_n14667_), .B0(new_n14664_), .B1(new_n14657_), .Y(new_n14668_));
  NAND2  g13666(.A(new_n14668_), .B(new_n14654_), .Y(new_n14669_));
  AOI22  g13667(.A0(new_n13074_), .A1(new_n13065_), .B0(new_n13051_), .B1(new_n13044_), .Y(new_n14670_));
  AOI21  g13668(.A0(new_n13027_), .A1(new_n13026_), .B0(new_n14670_), .Y(new_n14671_));
  AOI21  g13669(.A0(new_n13045_), .A1(new_n12039_), .B0(new_n13037_), .Y(new_n14672_));
  XOR2   g13670(.A(new_n13049_), .B(new_n13039_), .Y(new_n14673_));
  NOR2   g13671(.A(new_n14673_), .B(new_n14672_), .Y(new_n14674_));
  NOR2   g13672(.A(new_n13049_), .B(new_n13039_), .Y(new_n14675_));
  NAND4  g13673(.A(new_n12068_), .B(new_n12064_), .C(new_n12054_), .D(new_n12050_), .Y(new_n14676_));
  OAI211 g13674(.A0(new_n13040_), .A1(new_n12045_), .B0(new_n13041_), .B1(new_n13039_), .Y(new_n14677_));
  NAND2  g13675(.A(new_n14677_), .B(new_n14676_), .Y(new_n14678_));
  NOR3   g13676(.A(new_n14678_), .B(new_n14675_), .C(new_n13031_), .Y(new_n14679_));
  AOI21  g13677(.A0(new_n13066_), .A1(new_n12004_), .B0(new_n13058_), .Y(new_n14680_));
  AOI21  g13678(.A0(new_n13073_), .A1(new_n13069_), .B0(new_n14680_), .Y(new_n14681_));
  NAND2  g13679(.A(new_n13069_), .B(new_n13068_), .Y(new_n14682_));
  AOI211 g13680(.A0(new_n13063_), .A1(new_n13072_), .B(new_n14682_), .C(new_n13055_), .Y(new_n14683_));
  NOR4   g13681(.A(new_n14683_), .B(new_n14681_), .C(new_n14679_), .D(new_n14674_), .Y(new_n14684_));
  AOI211 g13682(.A0(new_n13047_), .A1(new_n12048_), .B(new_n13048_), .C(new_n13039_), .Y(new_n14685_));
  NAND2  g13683(.A(new_n13042_), .B(new_n13039_), .Y(new_n14686_));
  OAI21  g13684(.A0(new_n14685_), .A1(new_n14672_), .B0(new_n14686_), .Y(new_n14687_));
  NOR2   g13685(.A(new_n13063_), .B(new_n13060_), .Y(new_n14688_));
  NAND2  g13686(.A(new_n13063_), .B(new_n13060_), .Y(new_n14689_));
  OAI21  g13687(.A0(new_n14688_), .A1(new_n14680_), .B0(new_n14689_), .Y(new_n14690_));
  XOR2   g13688(.A(new_n14690_), .B(new_n14687_), .Y(new_n14691_));
  OAI21  g13689(.A0(new_n14684_), .A1(new_n14671_), .B0(new_n14691_), .Y(new_n14692_));
  NOR2   g13690(.A(new_n13036_), .B(new_n13035_), .Y(new_n14693_));
  XOR2   g13691(.A(new_n14693_), .B(new_n12055_), .Y(new_n14694_));
  XOR2   g13692(.A(new_n14694_), .B(new_n12039_), .Y(new_n14695_));
  NAND2  g13693(.A(new_n14695_), .B(new_n12037_), .Y(new_n14696_));
  NOR2   g13694(.A(new_n14695_), .B(new_n12037_), .Y(new_n14697_));
  AOI21  g13695(.A0(new_n14696_), .A1(new_n13015_), .B0(new_n14697_), .Y(new_n14698_));
  NOR2   g13696(.A(new_n14688_), .B(new_n14680_), .Y(new_n14699_));
  AOI21  g13697(.A0(new_n13063_), .A1(new_n13060_), .B0(new_n14699_), .Y(new_n14700_));
  AOI21  g13698(.A0(new_n14700_), .A1(new_n14687_), .B0(new_n14684_), .Y(new_n14701_));
  OAI221 g13699(.A0(new_n14700_), .A1(new_n14687_), .C0(new_n14701_), .B0(new_n14670_), .B1(new_n14698_), .Y(new_n14702_));
  NAND2  g13700(.A(new_n14702_), .B(new_n14692_), .Y(new_n14703_));
  XOR2   g13701(.A(new_n14703_), .B(new_n14669_), .Y(new_n14704_));
  XOR2   g13702(.A(new_n14704_), .B(new_n14629_), .Y(new_n14705_));
  NOR2   g13703(.A(new_n13009_), .B(new_n12965_), .Y(new_n14706_));
  NAND2  g13704(.A(new_n13009_), .B(new_n12965_), .Y(new_n14707_));
  OAI21  g13705(.A0(new_n14706_), .A1(new_n14622_), .B0(new_n14707_), .Y(new_n14708_));
  AOI21  g13706(.A0(new_n10604_), .A1(new_n10582_), .B0(new_n10584_), .Y(new_n14709_));
  XOR2   g13707(.A(new_n12114_), .B(new_n14709_), .Y(new_n14710_));
  OAI22  g13708(.A0(new_n12144_), .A1(new_n12143_), .B0(new_n12142_), .B1(new_n10350_), .Y(new_n14711_));
  NAND2  g13709(.A(new_n10317_), .B(new_n10253_), .Y(new_n14712_));
  NAND4  g13710(.A(new_n12140_), .B(new_n12137_), .C(new_n14712_), .D(new_n10320_), .Y(new_n14713_));
  NAND2  g13711(.A(new_n14713_), .B(new_n14711_), .Y(new_n14714_));
  XOR2   g13712(.A(new_n14714_), .B(new_n12132_), .Y(new_n14715_));
  XOR2   g13713(.A(new_n14715_), .B(new_n12117_), .Y(new_n14716_));
  OAI22  g13714(.A0(new_n14716_), .A1(new_n14710_), .B0(new_n14615_), .B1(new_n11128_), .Y(new_n14717_));
  NAND2  g13715(.A(new_n14716_), .B(new_n14710_), .Y(new_n14718_));
  NAND2  g13716(.A(new_n12986_), .B(new_n12078_), .Y(new_n14719_));
  AOI21  g13717(.A0(new_n12994_), .A1(new_n12991_), .B0(new_n12987_), .Y(new_n14720_));
  OAI211 g13718(.A0(new_n12994_), .A1(new_n12991_), .B0(new_n14720_), .B1(new_n14719_), .Y(new_n14721_));
  OAI21  g13719(.A0(new_n12995_), .A1(new_n12988_), .B0(new_n14721_), .Y(new_n14722_));
  AOI22  g13720(.A0(new_n14722_), .A1(new_n12983_), .B0(new_n14718_), .B1(new_n14717_), .Y(new_n14723_));
  NOR2   g13721(.A(new_n12979_), .B(new_n12973_), .Y(new_n14724_));
  NOR2   g13722(.A(new_n12978_), .B(new_n12975_), .Y(new_n14725_));
  NAND4  g13723(.A(new_n14713_), .B(new_n14711_), .C(new_n12131_), .D(new_n12127_), .Y(new_n14726_));
  NOR3   g13724(.A(new_n12119_), .B(new_n12118_), .C(new_n10345_), .Y(new_n14727_));
  OAI21  g13725(.A0(new_n12118_), .A1(new_n10345_), .B0(new_n12119_), .Y(new_n14728_));
  OAI211 g13726(.A0(new_n14727_), .A1(new_n12122_), .B0(new_n14728_), .B1(new_n12975_), .Y(new_n14729_));
  NAND2  g13727(.A(new_n14729_), .B(new_n14726_), .Y(new_n14730_));
  AOI211 g13728(.A0(new_n12971_), .A1(new_n12117_), .B(new_n14730_), .C(new_n14725_), .Y(new_n14731_));
  NOR4   g13729(.A(new_n13006_), .B(new_n12996_), .C(new_n14731_), .D(new_n14724_), .Y(new_n14732_));
  AOI211 g13730(.A0(new_n12976_), .A1(new_n12125_), .B(new_n12977_), .C(new_n12975_), .Y(new_n14733_));
  OAI21  g13731(.A0(new_n14727_), .A1(new_n12122_), .B0(new_n14728_), .Y(new_n14734_));
  NAND2  g13732(.A(new_n14734_), .B(new_n12975_), .Y(new_n14735_));
  OAI21  g13733(.A0(new_n14733_), .A1(new_n12973_), .B0(new_n14735_), .Y(new_n14736_));
  NOR2   g13734(.A(new_n13002_), .B(new_n12991_), .Y(new_n14737_));
  NAND2  g13735(.A(new_n13002_), .B(new_n12991_), .Y(new_n14738_));
  OAI21  g13736(.A0(new_n14737_), .A1(new_n12988_), .B0(new_n14738_), .Y(new_n14739_));
  XOR2   g13737(.A(new_n14739_), .B(new_n14736_), .Y(new_n14740_));
  OAI21  g13738(.A0(new_n14732_), .A1(new_n14723_), .B0(new_n14740_), .Y(new_n14741_));
  NOR2   g13739(.A(new_n14731_), .B(new_n14724_), .Y(new_n14742_));
  NOR2   g13740(.A(new_n13007_), .B(new_n14742_), .Y(new_n14743_));
  NOR2   g13741(.A(new_n14737_), .B(new_n12988_), .Y(new_n14744_));
  AOI21  g13742(.A0(new_n13002_), .A1(new_n12991_), .B0(new_n14744_), .Y(new_n14745_));
  AOI21  g13743(.A0(new_n14745_), .A1(new_n14736_), .B0(new_n14732_), .Y(new_n14746_));
  OAI221 g13744(.A0(new_n14745_), .A1(new_n14736_), .C0(new_n14746_), .B0(new_n14743_), .B1(new_n12968_), .Y(new_n14747_));
  NAND2  g13745(.A(new_n14747_), .B(new_n14741_), .Y(new_n14748_));
  AOI22  g13746(.A0(new_n12962_), .A1(new_n12953_), .B0(new_n12939_), .B1(new_n12932_), .Y(new_n14749_));
  AOI21  g13747(.A0(new_n12915_), .A1(new_n12914_), .B0(new_n14749_), .Y(new_n14750_));
  AOI21  g13748(.A0(new_n12933_), .A1(new_n12189_), .B0(new_n12925_), .Y(new_n14751_));
  XOR2   g13749(.A(new_n12937_), .B(new_n12927_), .Y(new_n14752_));
  NOR2   g13750(.A(new_n14752_), .B(new_n14751_), .Y(new_n14753_));
  NOR2   g13751(.A(new_n12937_), .B(new_n12927_), .Y(new_n14754_));
  NAND4  g13752(.A(new_n12218_), .B(new_n12214_), .C(new_n12204_), .D(new_n12200_), .Y(new_n14755_));
  OAI211 g13753(.A0(new_n12928_), .A1(new_n12195_), .B0(new_n12929_), .B1(new_n12927_), .Y(new_n14756_));
  NAND2  g13754(.A(new_n14756_), .B(new_n14755_), .Y(new_n14757_));
  NOR3   g13755(.A(new_n14757_), .B(new_n14754_), .C(new_n12919_), .Y(new_n14758_));
  AOI21  g13756(.A0(new_n12954_), .A1(new_n12154_), .B0(new_n12946_), .Y(new_n14759_));
  AOI21  g13757(.A0(new_n12961_), .A1(new_n12957_), .B0(new_n14759_), .Y(new_n14760_));
  NAND2  g13758(.A(new_n12957_), .B(new_n12956_), .Y(new_n14761_));
  AOI211 g13759(.A0(new_n12951_), .A1(new_n12960_), .B(new_n14761_), .C(new_n12943_), .Y(new_n14762_));
  NOR4   g13760(.A(new_n14762_), .B(new_n14760_), .C(new_n14758_), .D(new_n14753_), .Y(new_n14763_));
  AOI211 g13761(.A0(new_n12935_), .A1(new_n12198_), .B(new_n12936_), .C(new_n12927_), .Y(new_n14764_));
  NAND2  g13762(.A(new_n12930_), .B(new_n12927_), .Y(new_n14765_));
  OAI21  g13763(.A0(new_n14764_), .A1(new_n14751_), .B0(new_n14765_), .Y(new_n14766_));
  NOR2   g13764(.A(new_n12951_), .B(new_n12948_), .Y(new_n14767_));
  NAND2  g13765(.A(new_n12951_), .B(new_n12948_), .Y(new_n14768_));
  OAI21  g13766(.A0(new_n14767_), .A1(new_n14759_), .B0(new_n14768_), .Y(new_n14769_));
  XOR2   g13767(.A(new_n14769_), .B(new_n14766_), .Y(new_n14770_));
  OAI21  g13768(.A0(new_n14763_), .A1(new_n14750_), .B0(new_n14770_), .Y(new_n14771_));
  NOR2   g13769(.A(new_n12924_), .B(new_n12923_), .Y(new_n14772_));
  XOR2   g13770(.A(new_n14772_), .B(new_n12205_), .Y(new_n14773_));
  XOR2   g13771(.A(new_n14773_), .B(new_n12189_), .Y(new_n14774_));
  NAND2  g13772(.A(new_n14774_), .B(new_n12187_), .Y(new_n14775_));
  NOR2   g13773(.A(new_n14774_), .B(new_n12187_), .Y(new_n14776_));
  AOI21  g13774(.A0(new_n14775_), .A1(new_n14618_), .B0(new_n14776_), .Y(new_n14777_));
  NOR2   g13775(.A(new_n14767_), .B(new_n14759_), .Y(new_n14778_));
  AOI21  g13776(.A0(new_n12951_), .A1(new_n12948_), .B0(new_n14778_), .Y(new_n14779_));
  AOI21  g13777(.A0(new_n14779_), .A1(new_n14766_), .B0(new_n14763_), .Y(new_n14780_));
  OAI221 g13778(.A0(new_n14779_), .A1(new_n14766_), .C0(new_n14780_), .B0(new_n14749_), .B1(new_n14777_), .Y(new_n14781_));
  NAND2  g13779(.A(new_n14781_), .B(new_n14771_), .Y(new_n14782_));
  XOR2   g13780(.A(new_n14782_), .B(new_n14748_), .Y(new_n14783_));
  XOR2   g13781(.A(new_n14783_), .B(new_n14708_), .Y(new_n14784_));
  XOR2   g13782(.A(new_n14784_), .B(new_n14705_), .Y(new_n14785_));
  XOR2   g13783(.A(new_n14785_), .B(new_n14626_), .Y(new_n14786_));
  XOR2   g13784(.A(new_n14786_), .B(new_n14614_), .Y(new_n14787_));
  XOR2   g13785(.A(new_n14787_), .B(new_n14446_), .Y(new_n14788_));
  XOR2   g13786(.A(new_n14788_), .B(new_n14439_), .Y(new_n14789_));
  NAND2  g13787(.A(new_n14789_), .B(new_n14234_), .Y(new_n14790_));
  NOR2   g13788(.A(new_n13695_), .B(new_n13377_), .Y(new_n14791_));
  NAND2  g13789(.A(new_n13695_), .B(new_n13377_), .Y(new_n14792_));
  OAI21  g13790(.A0(new_n14791_), .A1(new_n13702_), .B0(new_n14792_), .Y(new_n14793_));
  XOR2   g13791(.A(new_n14789_), .B(new_n14793_), .Y(new_n14794_));
  NOR2   g13792(.A(new_n12877_), .B(new_n12553_), .Y(new_n14795_));
  NAND2  g13793(.A(new_n12877_), .B(new_n12553_), .Y(new_n14796_));
  OAI21  g13794(.A0(new_n14795_), .A1(new_n12240_), .B0(new_n14796_), .Y(new_n14797_));
  NOR2   g13795(.A(new_n12875_), .B(new_n12714_), .Y(new_n14798_));
  NAND2  g13796(.A(new_n12875_), .B(new_n12714_), .Y(new_n14799_));
  OAI21  g13797(.A0(new_n14798_), .A1(new_n13712_), .B0(new_n14799_), .Y(new_n14800_));
  XOR2   g13798(.A(new_n13952_), .B(new_n14800_), .Y(new_n14801_));
  NAND2  g13799(.A(new_n14223_), .B(new_n14801_), .Y(new_n14802_));
  NOR2   g13800(.A(new_n14223_), .B(new_n14801_), .Y(new_n14803_));
  AOI21  g13801(.A0(new_n14802_), .A1(new_n14797_), .B0(new_n14803_), .Y(new_n14804_));
  NOR2   g13802(.A(new_n14164_), .B(new_n4749_), .Y(new_n14805_));
  XOR2   g13803(.A(new_n12321_), .B(new_n14805_), .Y(new_n14806_));
  NOR2   g13804(.A(new_n14097_), .B(new_n4465_), .Y(new_n14807_));
  XOR2   g13805(.A(new_n12393_), .B(new_n14807_), .Y(new_n14808_));
  NAND2  g13806(.A(new_n14808_), .B(new_n14806_), .Y(new_n14809_));
  NOR2   g13807(.A(new_n14808_), .B(new_n14806_), .Y(new_n14810_));
  AOI21  g13808(.A0(new_n14809_), .A1(new_n12242_), .B0(new_n14810_), .Y(new_n14811_));
  XOR2   g13809(.A(new_n14220_), .B(new_n14811_), .Y(new_n14812_));
  NAND2  g13810(.A(new_n14812_), .B(new_n14092_), .Y(new_n14813_));
  NOR2   g13811(.A(new_n14812_), .B(new_n14092_), .Y(new_n14814_));
  AOI21  g13812(.A0(new_n14813_), .A1(new_n13956_), .B0(new_n14814_), .Y(new_n14815_));
  NOR2   g13813(.A(new_n14219_), .B(new_n14161_), .Y(new_n14816_));
  NAND2  g13814(.A(new_n14219_), .B(new_n14161_), .Y(new_n14817_));
  OAI21  g13815(.A0(new_n14816_), .A1(new_n14811_), .B0(new_n14817_), .Y(new_n14818_));
  AOI22  g13816(.A0(new_n14217_), .A1(new_n14196_), .B0(new_n14174_), .B1(new_n14166_), .Y(new_n14819_));
  NOR2   g13817(.A(new_n14187_), .B(new_n14180_), .Y(new_n14820_));
  AOI211 g13818(.A0(new_n14176_), .A1(new_n12284_), .B(new_n14193_), .C(new_n14192_), .Y(new_n14821_));
  NOR2   g13819(.A(new_n14208_), .B(new_n14201_), .Y(new_n14822_));
  NAND3  g13820(.A(new_n14215_), .B(new_n14211_), .C(new_n14210_), .Y(new_n14823_));
  AOI21  g13821(.A0(new_n14199_), .A1(new_n12247_), .B0(new_n14823_), .Y(new_n14824_));
  NOR4   g13822(.A(new_n14824_), .B(new_n14822_), .C(new_n14821_), .D(new_n14820_), .Y(new_n14825_));
  AOI221 g13823(.A0(new_n14182_), .A1(new_n12308_), .C0(new_n14186_), .B0(new_n12310_), .B1(new_n14181_), .Y(new_n14826_));
  INV    g13824(.A(new_n14183_), .Y(new_n14827_));
  NAND2  g13825(.A(new_n14186_), .B(new_n14827_), .Y(new_n14828_));
  OAI21  g13826(.A0(new_n14826_), .A1(new_n14180_), .B0(new_n14828_), .Y(new_n14829_));
  NOR2   g13827(.A(new_n14214_), .B(new_n14204_), .Y(new_n14830_));
  NAND2  g13828(.A(new_n14214_), .B(new_n14204_), .Y(new_n14831_));
  OAI21  g13829(.A0(new_n14830_), .A1(new_n14201_), .B0(new_n14831_), .Y(new_n14832_));
  XOR2   g13830(.A(new_n14832_), .B(new_n14829_), .Y(new_n14833_));
  OAI21  g13831(.A0(new_n14825_), .A1(new_n14819_), .B0(new_n14833_), .Y(new_n14834_));
  NOR2   g13832(.A(new_n12320_), .B(new_n12283_), .Y(new_n14835_));
  AOI21  g13833(.A0(new_n14165_), .A1(new_n12243_), .B0(new_n14835_), .Y(new_n14836_));
  OAI21  g13834(.A0(new_n14178_), .A1(new_n12313_), .B0(new_n14188_), .Y(new_n14837_));
  INV    g13835(.A(new_n14187_), .Y(new_n14838_));
  NAND2  g13836(.A(new_n14838_), .B(new_n14837_), .Y(new_n14839_));
  NAND2  g13837(.A(new_n14210_), .B(new_n14209_), .Y(new_n14840_));
  INV    g13838(.A(new_n14208_), .Y(new_n14841_));
  NAND2  g13839(.A(new_n14841_), .B(new_n14840_), .Y(new_n14842_));
  AOI22  g13840(.A0(new_n14216_), .A1(new_n14842_), .B0(new_n14195_), .B1(new_n14839_), .Y(new_n14843_));
  NOR2   g13841(.A(new_n14830_), .B(new_n14201_), .Y(new_n14844_));
  AOI21  g13842(.A0(new_n14214_), .A1(new_n14204_), .B0(new_n14844_), .Y(new_n14845_));
  AOI21  g13843(.A0(new_n14845_), .A1(new_n14829_), .B0(new_n14825_), .Y(new_n14846_));
  OAI221 g13844(.A0(new_n14845_), .A1(new_n14829_), .C0(new_n14846_), .B0(new_n14843_), .B1(new_n14836_), .Y(new_n14847_));
  NAND2  g13845(.A(new_n14847_), .B(new_n14834_), .Y(new_n14848_));
  AOI22  g13846(.A0(new_n14158_), .A1(new_n14154_), .B0(new_n14130_), .B1(new_n14127_), .Y(new_n14849_));
  AOI21  g13847(.A0(new_n14103_), .A1(new_n14102_), .B0(new_n14849_), .Y(new_n14850_));
  OAI22  g13848(.A0(new_n12389_), .A1(new_n12385_), .B0(new_n14113_), .B1(new_n14112_), .Y(new_n14851_));
  AOI21  g13849(.A0(new_n14851_), .A1(new_n12360_), .B0(new_n14114_), .Y(new_n14852_));
  NAND2  g13850(.A(new_n14125_), .B(new_n14122_), .Y(new_n14853_));
  AOI21  g13851(.A0(new_n14128_), .A1(new_n14853_), .B0(new_n14852_), .Y(new_n14854_));
  NOR4   g13852(.A(new_n14126_), .B(new_n14119_), .C(new_n14114_), .D(new_n14110_), .Y(new_n14855_));
  AOI21  g13853(.A0(new_n14155_), .A1(new_n12325_), .B0(new_n14140_), .Y(new_n14856_));
  OAI221 g13854(.A0(new_n14144_), .A1(new_n12337_), .C0(new_n14149_), .B0(new_n12331_), .B1(new_n14137_), .Y(new_n14857_));
  NAND2  g13855(.A(new_n14145_), .B(new_n14143_), .Y(new_n14858_));
  AOI21  g13856(.A0(new_n14858_), .A1(new_n14857_), .B0(new_n14856_), .Y(new_n14859_));
  NOR4   g13857(.A(new_n14153_), .B(new_n14146_), .C(new_n14140_), .D(new_n14136_), .Y(new_n14860_));
  NOR4   g13858(.A(new_n14860_), .B(new_n14859_), .C(new_n14855_), .D(new_n14854_), .Y(new_n14861_));
  AOI221 g13859(.A0(new_n14115_), .A1(new_n12380_), .C0(new_n14118_), .B0(new_n12382_), .B1(new_n14106_), .Y(new_n14862_));
  NAND2  g13860(.A(new_n14118_), .B(new_n14122_), .Y(new_n14863_));
  OAI21  g13861(.A0(new_n14862_), .A1(new_n14852_), .B0(new_n14863_), .Y(new_n14864_));
  NOR2   g13862(.A(new_n14145_), .B(new_n14149_), .Y(new_n14865_));
  NAND2  g13863(.A(new_n14145_), .B(new_n14149_), .Y(new_n14866_));
  OAI21  g13864(.A0(new_n14865_), .A1(new_n14856_), .B0(new_n14866_), .Y(new_n14867_));
  XOR2   g13865(.A(new_n14867_), .B(new_n14864_), .Y(new_n14868_));
  OAI21  g13866(.A0(new_n14861_), .A1(new_n14850_), .B0(new_n14868_), .Y(new_n14869_));
  NAND2  g13867(.A(new_n12392_), .B(new_n12359_), .Y(new_n14870_));
  NOR2   g13868(.A(new_n12392_), .B(new_n12359_), .Y(new_n14871_));
  AOI21  g13869(.A0(new_n14870_), .A1(new_n12323_), .B0(new_n14871_), .Y(new_n14872_));
  NOR2   g13870(.A(new_n14865_), .B(new_n14856_), .Y(new_n14873_));
  AOI21  g13871(.A0(new_n14145_), .A1(new_n14149_), .B0(new_n14873_), .Y(new_n14874_));
  AOI21  g13872(.A0(new_n14874_), .A1(new_n14864_), .B0(new_n14861_), .Y(new_n14875_));
  OAI221 g13873(.A0(new_n14874_), .A1(new_n14864_), .C0(new_n14875_), .B0(new_n14849_), .B1(new_n14872_), .Y(new_n14876_));
  NAND2  g13874(.A(new_n14876_), .B(new_n14869_), .Y(new_n14877_));
  XOR2   g13875(.A(new_n14877_), .B(new_n14848_), .Y(new_n14878_));
  XOR2   g13876(.A(new_n14878_), .B(new_n14818_), .Y(new_n14879_));
  NOR2   g13877(.A(new_n14090_), .B(new_n14031_), .Y(new_n14880_));
  NAND2  g13878(.A(new_n14090_), .B(new_n14031_), .Y(new_n14881_));
  OAI21  g13879(.A0(new_n14880_), .A1(new_n13967_), .B0(new_n14881_), .Y(new_n14882_));
  AOI22  g13880(.A0(new_n14088_), .A1(new_n14063_), .B0(new_n14041_), .B1(new_n14033_), .Y(new_n14883_));
  NOR2   g13881(.A(new_n14054_), .B(new_n14047_), .Y(new_n14884_));
  AOI211 g13882(.A0(new_n14043_), .A1(new_n12439_), .B(new_n14060_), .C(new_n14059_), .Y(new_n14885_));
  NOR2   g13883(.A(new_n14075_), .B(new_n14068_), .Y(new_n14886_));
  AOI211 g13884(.A0(new_n14066_), .A1(new_n12402_), .B(new_n14085_), .C(new_n14077_), .Y(new_n14887_));
  NOR4   g13885(.A(new_n14887_), .B(new_n14886_), .C(new_n14885_), .D(new_n14884_), .Y(new_n14888_));
  AOI221 g13886(.A0(new_n14049_), .A1(new_n12463_), .C0(new_n14053_), .B0(new_n12465_), .B1(new_n14048_), .Y(new_n14889_));
  INV    g13887(.A(new_n14050_), .Y(new_n14890_));
  NAND2  g13888(.A(new_n14053_), .B(new_n14890_), .Y(new_n14891_));
  OAI21  g13889(.A0(new_n14889_), .A1(new_n14047_), .B0(new_n14891_), .Y(new_n14892_));
  NOR2   g13890(.A(new_n14084_), .B(new_n14071_), .Y(new_n14893_));
  NAND2  g13891(.A(new_n14084_), .B(new_n14071_), .Y(new_n14894_));
  OAI21  g13892(.A0(new_n14893_), .A1(new_n14068_), .B0(new_n14894_), .Y(new_n14895_));
  XOR2   g13893(.A(new_n14895_), .B(new_n14892_), .Y(new_n14896_));
  OAI21  g13894(.A0(new_n14888_), .A1(new_n14883_), .B0(new_n14896_), .Y(new_n14897_));
  NOR2   g13895(.A(new_n12475_), .B(new_n12438_), .Y(new_n14898_));
  AOI21  g13896(.A0(new_n14032_), .A1(new_n12398_), .B0(new_n14898_), .Y(new_n14899_));
  OAI21  g13897(.A0(new_n14045_), .A1(new_n12468_), .B0(new_n14055_), .Y(new_n14900_));
  INV    g13898(.A(new_n14054_), .Y(new_n14901_));
  NAND2  g13899(.A(new_n14901_), .B(new_n14900_), .Y(new_n14902_));
  NAND2  g13900(.A(new_n14078_), .B(new_n14076_), .Y(new_n14903_));
  INV    g13901(.A(new_n14075_), .Y(new_n14904_));
  NAND2  g13902(.A(new_n14904_), .B(new_n14903_), .Y(new_n14905_));
  AOI22  g13903(.A0(new_n14087_), .A1(new_n14905_), .B0(new_n14062_), .B1(new_n14902_), .Y(new_n14906_));
  NOR2   g13904(.A(new_n14893_), .B(new_n14068_), .Y(new_n14907_));
  AOI21  g13905(.A0(new_n14084_), .A1(new_n14071_), .B0(new_n14907_), .Y(new_n14908_));
  AOI21  g13906(.A0(new_n14908_), .A1(new_n14892_), .B0(new_n14888_), .Y(new_n14909_));
  OAI221 g13907(.A0(new_n14908_), .A1(new_n14892_), .C0(new_n14909_), .B0(new_n14906_), .B1(new_n14899_), .Y(new_n14910_));
  NAND2  g13908(.A(new_n14910_), .B(new_n14897_), .Y(new_n14911_));
  AOI22  g13909(.A0(new_n14028_), .A1(new_n14024_), .B0(new_n14000_), .B1(new_n13997_), .Y(new_n14912_));
  AOI21  g13910(.A0(new_n13973_), .A1(new_n13972_), .B0(new_n14912_), .Y(new_n14913_));
  OAI22  g13911(.A0(new_n12544_), .A1(new_n12540_), .B0(new_n13983_), .B1(new_n13982_), .Y(new_n14914_));
  AOI21  g13912(.A0(new_n14914_), .A1(new_n12515_), .B0(new_n13984_), .Y(new_n14915_));
  NAND2  g13913(.A(new_n13995_), .B(new_n13992_), .Y(new_n14916_));
  AOI21  g13914(.A0(new_n13998_), .A1(new_n14916_), .B0(new_n14915_), .Y(new_n14917_));
  NOR4   g13915(.A(new_n13996_), .B(new_n13989_), .C(new_n13984_), .D(new_n13980_), .Y(new_n14918_));
  AOI21  g13916(.A0(new_n14025_), .A1(new_n12480_), .B0(new_n14010_), .Y(new_n14919_));
  OAI221 g13917(.A0(new_n14014_), .A1(new_n12492_), .C0(new_n14019_), .B0(new_n12486_), .B1(new_n14007_), .Y(new_n14920_));
  NAND2  g13918(.A(new_n14015_), .B(new_n14013_), .Y(new_n14921_));
  AOI21  g13919(.A0(new_n14921_), .A1(new_n14920_), .B0(new_n14919_), .Y(new_n14922_));
  NOR4   g13920(.A(new_n14023_), .B(new_n14016_), .C(new_n14010_), .D(new_n14006_), .Y(new_n14923_));
  NOR4   g13921(.A(new_n14923_), .B(new_n14922_), .C(new_n14918_), .D(new_n14917_), .Y(new_n14924_));
  AOI221 g13922(.A0(new_n13985_), .A1(new_n12535_), .C0(new_n13988_), .B0(new_n12537_), .B1(new_n13976_), .Y(new_n14925_));
  NAND2  g13923(.A(new_n13988_), .B(new_n13992_), .Y(new_n14926_));
  OAI21  g13924(.A0(new_n14925_), .A1(new_n14915_), .B0(new_n14926_), .Y(new_n14927_));
  NOR2   g13925(.A(new_n14015_), .B(new_n14019_), .Y(new_n14928_));
  NAND2  g13926(.A(new_n14015_), .B(new_n14019_), .Y(new_n14929_));
  OAI21  g13927(.A0(new_n14928_), .A1(new_n14919_), .B0(new_n14929_), .Y(new_n14930_));
  XOR2   g13928(.A(new_n14930_), .B(new_n14927_), .Y(new_n14931_));
  OAI21  g13929(.A0(new_n14924_), .A1(new_n14913_), .B0(new_n14931_), .Y(new_n14932_));
  NAND2  g13930(.A(new_n12547_), .B(new_n12514_), .Y(new_n14933_));
  NOR2   g13931(.A(new_n12547_), .B(new_n12514_), .Y(new_n14934_));
  AOI21  g13932(.A0(new_n14933_), .A1(new_n12478_), .B0(new_n14934_), .Y(new_n14935_));
  NOR2   g13933(.A(new_n14928_), .B(new_n14919_), .Y(new_n14936_));
  AOI21  g13934(.A0(new_n14015_), .A1(new_n14019_), .B0(new_n14936_), .Y(new_n14937_));
  AOI21  g13935(.A0(new_n14937_), .A1(new_n14927_), .B0(new_n14924_), .Y(new_n14938_));
  OAI221 g13936(.A0(new_n14937_), .A1(new_n14927_), .C0(new_n14938_), .B0(new_n14912_), .B1(new_n14935_), .Y(new_n14939_));
  NAND2  g13937(.A(new_n14939_), .B(new_n14932_), .Y(new_n14940_));
  XOR2   g13938(.A(new_n14940_), .B(new_n14911_), .Y(new_n14941_));
  XOR2   g13939(.A(new_n14941_), .B(new_n14882_), .Y(new_n14942_));
  XOR2   g13940(.A(new_n14942_), .B(new_n14879_), .Y(new_n14943_));
  XOR2   g13941(.A(new_n14943_), .B(new_n14815_), .Y(new_n14944_));
  OAI21  g13942(.A0(new_n2138_), .A1(new_n2128_), .B0(new_n12718_), .Y(new_n14945_));
  NAND2  g13943(.A(new_n2143_), .B(new_n2022_), .Y(new_n14946_));
  AOI21  g13944(.A0(new_n14946_), .A1(new_n14945_), .B0(new_n2369_), .Y(new_n14947_));
  NOR2   g13945(.A(new_n14947_), .B(new_n2370_), .Y(new_n14948_));
  XOR2   g13946(.A(new_n12795_), .B(new_n14948_), .Y(new_n14949_));
  OAI21  g13947(.A0(new_n2824_), .A1(new_n2589_), .B0(new_n2836_), .Y(new_n14950_));
  XOR2   g13948(.A(new_n12872_), .B(new_n14950_), .Y(new_n14951_));
  NAND2  g13949(.A(new_n14951_), .B(new_n14949_), .Y(new_n14952_));
  NOR2   g13950(.A(new_n14951_), .B(new_n14949_), .Y(new_n14953_));
  AOI21  g13951(.A0(new_n14952_), .A1(new_n12715_), .B0(new_n14953_), .Y(new_n14954_));
  XOR2   g13952(.A(new_n13828_), .B(new_n14954_), .Y(new_n14955_));
  NAND2  g13953(.A(new_n13951_), .B(new_n14955_), .Y(new_n14956_));
  NOR2   g13954(.A(new_n13951_), .B(new_n14955_), .Y(new_n14957_));
  AOI21  g13955(.A0(new_n14956_), .A1(new_n14800_), .B0(new_n14957_), .Y(new_n14958_));
  NOR2   g13956(.A(new_n13949_), .B(new_n13890_), .Y(new_n14959_));
  NAND2  g13957(.A(new_n13949_), .B(new_n13890_), .Y(new_n14960_));
  OAI21  g13958(.A0(new_n14959_), .A1(new_n13839_), .B0(new_n14960_), .Y(new_n14961_));
  AOI22  g13959(.A0(new_n13947_), .A1(new_n13922_), .B0(new_n13900_), .B1(new_n13892_), .Y(new_n14962_));
  NOR2   g13960(.A(new_n13913_), .B(new_n13906_), .Y(new_n14963_));
  AOI211 g13961(.A0(new_n13902_), .A1(new_n12597_), .B(new_n13919_), .C(new_n13918_), .Y(new_n14964_));
  NOR2   g13962(.A(new_n13934_), .B(new_n13927_), .Y(new_n14965_));
  AOI211 g13963(.A0(new_n13925_), .A1(new_n12560_), .B(new_n13944_), .C(new_n13936_), .Y(new_n14966_));
  NOR4   g13964(.A(new_n14966_), .B(new_n14965_), .C(new_n14964_), .D(new_n14963_), .Y(new_n14967_));
  AOI221 g13965(.A0(new_n13908_), .A1(new_n12621_), .C0(new_n13912_), .B0(new_n12623_), .B1(new_n13907_), .Y(new_n14968_));
  INV    g13966(.A(new_n13909_), .Y(new_n14969_));
  NAND2  g13967(.A(new_n13912_), .B(new_n14969_), .Y(new_n14970_));
  OAI21  g13968(.A0(new_n14968_), .A1(new_n13906_), .B0(new_n14970_), .Y(new_n14971_));
  NOR2   g13969(.A(new_n13943_), .B(new_n13930_), .Y(new_n14972_));
  NAND2  g13970(.A(new_n13943_), .B(new_n13930_), .Y(new_n14973_));
  OAI21  g13971(.A0(new_n14972_), .A1(new_n13927_), .B0(new_n14973_), .Y(new_n14974_));
  XOR2   g13972(.A(new_n14974_), .B(new_n14971_), .Y(new_n14975_));
  OAI21  g13973(.A0(new_n14967_), .A1(new_n14962_), .B0(new_n14975_), .Y(new_n14976_));
  NOR2   g13974(.A(new_n12633_), .B(new_n12596_), .Y(new_n14977_));
  AOI21  g13975(.A0(new_n13891_), .A1(new_n12556_), .B0(new_n14977_), .Y(new_n14978_));
  OAI21  g13976(.A0(new_n13904_), .A1(new_n12626_), .B0(new_n13914_), .Y(new_n14979_));
  INV    g13977(.A(new_n13913_), .Y(new_n14980_));
  NAND2  g13978(.A(new_n14980_), .B(new_n14979_), .Y(new_n14981_));
  NAND2  g13979(.A(new_n13937_), .B(new_n13935_), .Y(new_n14982_));
  INV    g13980(.A(new_n13934_), .Y(new_n14983_));
  NAND2  g13981(.A(new_n14983_), .B(new_n14982_), .Y(new_n14984_));
  AOI22  g13982(.A0(new_n13946_), .A1(new_n14984_), .B0(new_n13921_), .B1(new_n14981_), .Y(new_n14985_));
  NOR2   g13983(.A(new_n14972_), .B(new_n13927_), .Y(new_n14986_));
  AOI21  g13984(.A0(new_n13943_), .A1(new_n13930_), .B0(new_n14986_), .Y(new_n14987_));
  AOI21  g13985(.A0(new_n14987_), .A1(new_n14971_), .B0(new_n14967_), .Y(new_n14988_));
  OAI221 g13986(.A0(new_n14987_), .A1(new_n14971_), .C0(new_n14988_), .B0(new_n14985_), .B1(new_n14978_), .Y(new_n14989_));
  NAND2  g13987(.A(new_n14989_), .B(new_n14976_), .Y(new_n14990_));
  OAI22  g13988(.A0(new_n13849_), .A1(new_n13848_), .B0(new_n13847_), .B1(new_n13846_), .Y(new_n14991_));
  NAND2  g13989(.A(new_n14991_), .B(new_n12674_), .Y(new_n14992_));
  OAI211 g13990(.A0(new_n13861_), .A1(new_n13853_), .B0(new_n13862_), .B1(new_n14992_), .Y(new_n14993_));
  XOR2   g13991(.A(new_n13879_), .B(new_n13884_), .Y(new_n14994_));
  OAI21  g13992(.A0(new_n13874_), .A1(new_n13869_), .B0(new_n14994_), .Y(new_n14995_));
  NAND2  g13993(.A(new_n13873_), .B(new_n12639_), .Y(new_n14996_));
  NAND4  g13994(.A(new_n13886_), .B(new_n13885_), .C(new_n13881_), .D(new_n14996_), .Y(new_n14997_));
  AOI22  g13995(.A0(new_n14997_), .A1(new_n14995_), .B0(new_n14993_), .B1(new_n13858_), .Y(new_n14998_));
  AOI21  g13996(.A0(new_n13843_), .A1(new_n13842_), .B0(new_n14998_), .Y(new_n14999_));
  NOR2   g13997(.A(new_n13880_), .B(new_n13875_), .Y(new_n15000_));
  OAI221 g13998(.A0(new_n13887_), .A1(new_n13869_), .C0(new_n13858_), .B0(new_n13863_), .B1(new_n13845_), .Y(new_n15001_));
  NOR2   g13999(.A(new_n15001_), .B(new_n15000_), .Y(new_n15002_));
  NOR2   g14000(.A(new_n13850_), .B(new_n13845_), .Y(new_n15003_));
  NOR2   g14001(.A(new_n13856_), .B(new_n13853_), .Y(new_n15004_));
  NAND2  g14002(.A(new_n13856_), .B(new_n13853_), .Y(new_n15005_));
  OAI21  g14003(.A0(new_n15004_), .A1(new_n15003_), .B0(new_n15005_), .Y(new_n15006_));
  NOR2   g14004(.A(new_n13879_), .B(new_n13884_), .Y(new_n15007_));
  NAND2  g14005(.A(new_n13879_), .B(new_n13884_), .Y(new_n15008_));
  OAI21  g14006(.A0(new_n15007_), .A1(new_n13875_), .B0(new_n15008_), .Y(new_n15009_));
  XOR2   g14007(.A(new_n15009_), .B(new_n15006_), .Y(new_n15010_));
  OAI21  g14008(.A0(new_n15002_), .A1(new_n14999_), .B0(new_n15010_), .Y(new_n15011_));
  NOR2   g14009(.A(new_n13849_), .B(new_n13848_), .Y(new_n15012_));
  XOR2   g14010(.A(new_n15012_), .B(new_n12693_), .Y(new_n15013_));
  XOR2   g14011(.A(new_n15013_), .B(new_n12674_), .Y(new_n15014_));
  NAND2  g14012(.A(new_n15014_), .B(new_n12671_), .Y(new_n15015_));
  NOR2   g14013(.A(new_n15014_), .B(new_n12671_), .Y(new_n15016_));
  AOI21  g14014(.A0(new_n15015_), .A1(new_n13835_), .B0(new_n15016_), .Y(new_n15017_));
  NOR2   g14015(.A(new_n15007_), .B(new_n13875_), .Y(new_n15018_));
  AOI21  g14016(.A0(new_n13879_), .A1(new_n13884_), .B0(new_n15018_), .Y(new_n15019_));
  AOI21  g14017(.A0(new_n15019_), .A1(new_n15006_), .B0(new_n15002_), .Y(new_n15020_));
  OAI221 g14018(.A0(new_n15019_), .A1(new_n15006_), .C0(new_n15020_), .B0(new_n14998_), .B1(new_n15017_), .Y(new_n15021_));
  NAND2  g14019(.A(new_n15021_), .B(new_n15011_), .Y(new_n15022_));
  XOR2   g14020(.A(new_n15022_), .B(new_n14990_), .Y(new_n15023_));
  XOR2   g14021(.A(new_n15023_), .B(new_n14961_), .Y(new_n15024_));
  NOR2   g14022(.A(new_n13827_), .B(new_n13777_), .Y(new_n15025_));
  NAND2  g14023(.A(new_n13827_), .B(new_n13777_), .Y(new_n15026_));
  OAI21  g14024(.A0(new_n15025_), .A1(new_n14954_), .B0(new_n15026_), .Y(new_n15027_));
  NAND2  g14025(.A(new_n13815_), .B(new_n13814_), .Y(new_n15028_));
  XOR2   g14026(.A(new_n15028_), .B(new_n12740_), .Y(new_n15029_));
  XOR2   g14027(.A(new_n15029_), .B(new_n12720_), .Y(new_n15030_));
  XOR2   g14028(.A(new_n13786_), .B(new_n12777_), .Y(new_n15031_));
  XOR2   g14029(.A(new_n15031_), .B(new_n12758_), .Y(new_n15032_));
  OAI22  g14030(.A0(new_n15032_), .A1(new_n15030_), .B0(new_n14947_), .B1(new_n2370_), .Y(new_n15033_));
  NAND2  g14031(.A(new_n15032_), .B(new_n15030_), .Y(new_n15034_));
  NAND2  g14032(.A(new_n13802_), .B(new_n12720_), .Y(new_n15035_));
  NOR2   g14033(.A(new_n13823_), .B(new_n13813_), .Y(new_n15036_));
  NAND2  g14034(.A(new_n15036_), .B(new_n15035_), .Y(new_n15037_));
  OAI21  g14035(.A0(new_n13811_), .A1(new_n13804_), .B0(new_n15037_), .Y(new_n15038_));
  AOI22  g14036(.A0(new_n15038_), .A1(new_n13799_), .B0(new_n15034_), .B1(new_n15033_), .Y(new_n15039_));
  NOR2   g14037(.A(new_n13795_), .B(new_n13789_), .Y(new_n15040_));
  NOR2   g14038(.A(new_n13794_), .B(new_n13792_), .Y(new_n15041_));
  NAND4  g14039(.A(new_n13785_), .B(new_n13784_), .C(new_n12776_), .D(new_n12773_), .Y(new_n15042_));
  NAND2  g14040(.A(new_n13794_), .B(new_n13792_), .Y(new_n15043_));
  NAND2  g14041(.A(new_n15043_), .B(new_n15042_), .Y(new_n15044_));
  AOI211 g14042(.A0(new_n13787_), .A1(new_n12758_), .B(new_n15044_), .C(new_n15041_), .Y(new_n15045_));
  NOR4   g14043(.A(new_n13824_), .B(new_n13812_), .C(new_n15045_), .D(new_n15040_), .Y(new_n15046_));
  AOI221 g14044(.A0(new_n13793_), .A1(new_n12771_), .C0(new_n13792_), .B0(new_n12763_), .B1(new_n12762_), .Y(new_n15047_));
  INV    g14045(.A(new_n13794_), .Y(new_n15048_));
  NAND2  g14046(.A(new_n15048_), .B(new_n13792_), .Y(new_n15049_));
  OAI21  g14047(.A0(new_n15047_), .A1(new_n13789_), .B0(new_n15049_), .Y(new_n15050_));
  NOR2   g14048(.A(new_n13822_), .B(new_n13807_), .Y(new_n15051_));
  NAND2  g14049(.A(new_n13822_), .B(new_n13807_), .Y(new_n15052_));
  OAI21  g14050(.A0(new_n15051_), .A1(new_n13804_), .B0(new_n15052_), .Y(new_n15053_));
  XOR2   g14051(.A(new_n15053_), .B(new_n15050_), .Y(new_n15054_));
  OAI21  g14052(.A0(new_n15046_), .A1(new_n15039_), .B0(new_n15054_), .Y(new_n15055_));
  NOR2   g14053(.A(new_n15045_), .B(new_n15040_), .Y(new_n15056_));
  NOR2   g14054(.A(new_n13825_), .B(new_n15056_), .Y(new_n15057_));
  NOR2   g14055(.A(new_n15051_), .B(new_n13804_), .Y(new_n15058_));
  AOI21  g14056(.A0(new_n13822_), .A1(new_n13807_), .B0(new_n15058_), .Y(new_n15059_));
  AOI21  g14057(.A0(new_n15059_), .A1(new_n15050_), .B0(new_n15046_), .Y(new_n15060_));
  OAI221 g14058(.A0(new_n15059_), .A1(new_n15050_), .C0(new_n15060_), .B0(new_n15057_), .B1(new_n13780_), .Y(new_n15061_));
  NAND2  g14059(.A(new_n15061_), .B(new_n15055_), .Y(new_n15062_));
  OAI22  g14060(.A0(new_n13736_), .A1(new_n13735_), .B0(new_n13734_), .B1(new_n13733_), .Y(new_n15063_));
  NAND2  g14061(.A(new_n15063_), .B(new_n12835_), .Y(new_n15064_));
  OAI211 g14062(.A0(new_n13748_), .A1(new_n13740_), .B0(new_n13749_), .B1(new_n15064_), .Y(new_n15065_));
  XOR2   g14063(.A(new_n13766_), .B(new_n13771_), .Y(new_n15066_));
  OAI21  g14064(.A0(new_n13761_), .A1(new_n13756_), .B0(new_n15066_), .Y(new_n15067_));
  NAND2  g14065(.A(new_n13760_), .B(new_n12800_), .Y(new_n15068_));
  NAND4  g14066(.A(new_n13773_), .B(new_n13772_), .C(new_n13768_), .D(new_n15068_), .Y(new_n15069_));
  AOI22  g14067(.A0(new_n15069_), .A1(new_n15067_), .B0(new_n15065_), .B1(new_n13745_), .Y(new_n15070_));
  AOI21  g14068(.A0(new_n13730_), .A1(new_n13729_), .B0(new_n15070_), .Y(new_n15071_));
  NOR2   g14069(.A(new_n13767_), .B(new_n13762_), .Y(new_n15072_));
  OAI221 g14070(.A0(new_n13774_), .A1(new_n13756_), .C0(new_n13745_), .B0(new_n13750_), .B1(new_n13732_), .Y(new_n15073_));
  NOR2   g14071(.A(new_n15073_), .B(new_n15072_), .Y(new_n15074_));
  NOR2   g14072(.A(new_n13737_), .B(new_n13732_), .Y(new_n15075_));
  NOR2   g14073(.A(new_n13743_), .B(new_n13740_), .Y(new_n15076_));
  NAND2  g14074(.A(new_n13743_), .B(new_n13740_), .Y(new_n15077_));
  OAI21  g14075(.A0(new_n15076_), .A1(new_n15075_), .B0(new_n15077_), .Y(new_n15078_));
  NOR2   g14076(.A(new_n13766_), .B(new_n13771_), .Y(new_n15079_));
  NAND2  g14077(.A(new_n13766_), .B(new_n13771_), .Y(new_n15080_));
  OAI21  g14078(.A0(new_n15079_), .A1(new_n13762_), .B0(new_n15080_), .Y(new_n15081_));
  XOR2   g14079(.A(new_n15081_), .B(new_n15078_), .Y(new_n15082_));
  OAI21  g14080(.A0(new_n15074_), .A1(new_n15071_), .B0(new_n15082_), .Y(new_n15083_));
  NOR2   g14081(.A(new_n13736_), .B(new_n13735_), .Y(new_n15084_));
  XOR2   g14082(.A(new_n15084_), .B(new_n12854_), .Y(new_n15085_));
  XOR2   g14083(.A(new_n15085_), .B(new_n12835_), .Y(new_n15086_));
  NAND2  g14084(.A(new_n15086_), .B(new_n12832_), .Y(new_n15087_));
  NOR2   g14085(.A(new_n15086_), .B(new_n12832_), .Y(new_n15088_));
  AOI21  g14086(.A0(new_n15087_), .A1(new_n14950_), .B0(new_n15088_), .Y(new_n15089_));
  NOR2   g14087(.A(new_n15079_), .B(new_n13762_), .Y(new_n15090_));
  AOI21  g14088(.A0(new_n13766_), .A1(new_n13771_), .B0(new_n15090_), .Y(new_n15091_));
  AOI21  g14089(.A0(new_n15091_), .A1(new_n15078_), .B0(new_n15074_), .Y(new_n15092_));
  OAI221 g14090(.A0(new_n15091_), .A1(new_n15078_), .C0(new_n15092_), .B0(new_n15070_), .B1(new_n15089_), .Y(new_n15093_));
  NAND2  g14091(.A(new_n15093_), .B(new_n15083_), .Y(new_n15094_));
  XOR2   g14092(.A(new_n15094_), .B(new_n15062_), .Y(new_n15095_));
  XOR2   g14093(.A(new_n15095_), .B(new_n15027_), .Y(new_n15096_));
  XOR2   g14094(.A(new_n15096_), .B(new_n15024_), .Y(new_n15097_));
  XOR2   g14095(.A(new_n15097_), .B(new_n14958_), .Y(new_n15098_));
  XOR2   g14096(.A(new_n15098_), .B(new_n14944_), .Y(new_n15099_));
  XOR2   g14097(.A(new_n15099_), .B(new_n14804_), .Y(new_n15100_));
  NAND2  g14098(.A(new_n15100_), .B(new_n14794_), .Y(new_n15101_));
  NAND2  g14099(.A(new_n13553_), .B(new_n13692_), .Y(new_n15102_));
  AOI21  g14100(.A0(new_n13552_), .A1(new_n15102_), .B0(new_n13690_), .Y(new_n15103_));
  NAND2  g14101(.A(new_n14242_), .B(new_n13552_), .Y(new_n15104_));
  OAI21  g14102(.A0(new_n15103_), .A1(new_n13384_), .B0(new_n15104_), .Y(new_n15105_));
  XOR2   g14103(.A(new_n14438_), .B(new_n15105_), .Y(new_n15106_));
  XOR2   g14104(.A(new_n14788_), .B(new_n15106_), .Y(new_n15107_));
  AOI21  g14105(.A0(new_n15107_), .A1(new_n14793_), .B0(new_n15100_), .Y(new_n15108_));
  AOI22  g14106(.A0(new_n15108_), .A1(new_n14790_), .B0(new_n15101_), .B1(new_n14228_), .Y(new_n15109_));
  NOR2   g14107(.A(new_n14788_), .B(new_n15106_), .Y(new_n15110_));
  NAND2  g14108(.A(new_n14788_), .B(new_n15106_), .Y(new_n15111_));
  OAI21  g14109(.A0(new_n15110_), .A1(new_n14234_), .B0(new_n15111_), .Y(new_n15112_));
  AOI21  g14110(.A0(new_n11150_), .A1(new_n10118_), .B0(new_n10120_), .Y(new_n15113_));
  XOR2   g14111(.A(new_n12074_), .B(new_n15113_), .Y(new_n15114_));
  XOR2   g14112(.A(new_n12224_), .B(new_n12904_), .Y(new_n15115_));
  NAND2  g14113(.A(new_n15115_), .B(new_n15114_), .Y(new_n15116_));
  NOR2   g14114(.A(new_n15115_), .B(new_n15114_), .Y(new_n15117_));
  AOI21  g14115(.A0(new_n15116_), .A1(new_n11919_), .B0(new_n15117_), .Y(new_n15118_));
  XOR2   g14116(.A(new_n13130_), .B(new_n15118_), .Y(new_n15119_));
  NOR2   g14117(.A(new_n13375_), .B(new_n15119_), .Y(new_n15120_));
  NAND2  g14118(.A(new_n13375_), .B(new_n15119_), .Y(new_n15121_));
  OAI21  g14119(.A0(new_n15120_), .A1(new_n12900_), .B0(new_n15121_), .Y(new_n15122_));
  XOR2   g14120(.A(new_n13245_), .B(new_n14533_), .Y(new_n15123_));
  NAND2  g14121(.A(new_n13373_), .B(new_n15123_), .Y(new_n15124_));
  NOR2   g14122(.A(new_n13373_), .B(new_n15123_), .Y(new_n15125_));
  AOI21  g14123(.A0(new_n15124_), .A1(new_n14442_), .B0(new_n15125_), .Y(new_n15126_));
  XOR2   g14124(.A(new_n14613_), .B(new_n15126_), .Y(new_n15127_));
  NAND2  g14125(.A(new_n14786_), .B(new_n15127_), .Y(new_n15128_));
  NOR2   g14126(.A(new_n14786_), .B(new_n15127_), .Y(new_n15129_));
  AOI21  g14127(.A0(new_n15128_), .A1(new_n15122_), .B0(new_n15129_), .Y(new_n15130_));
  NOR2   g14128(.A(new_n14784_), .B(new_n14705_), .Y(new_n15131_));
  NAND2  g14129(.A(new_n14784_), .B(new_n14705_), .Y(new_n15132_));
  OAI21  g14130(.A0(new_n15131_), .A1(new_n14626_), .B0(new_n15132_), .Y(new_n15133_));
  XOR2   g14131(.A(new_n12964_), .B(new_n14777_), .Y(new_n15134_));
  NAND2  g14132(.A(new_n14718_), .B(new_n14717_), .Y(new_n15135_));
  XOR2   g14133(.A(new_n13008_), .B(new_n15135_), .Y(new_n15136_));
  NAND2  g14134(.A(new_n15136_), .B(new_n15134_), .Y(new_n15137_));
  NOR2   g14135(.A(new_n15136_), .B(new_n15134_), .Y(new_n15138_));
  AOI21  g14136(.A0(new_n15137_), .A1(new_n12907_), .B0(new_n15138_), .Y(new_n15139_));
  AOI22  g14137(.A0(new_n14781_), .A1(new_n14771_), .B0(new_n14747_), .B1(new_n14741_), .Y(new_n15140_));
  NOR2   g14138(.A(new_n15140_), .B(new_n15139_), .Y(new_n15141_));
  NAND2  g14139(.A(new_n14782_), .B(new_n14748_), .Y(new_n15142_));
  NAND4  g14140(.A(new_n12962_), .B(new_n12953_), .C(new_n12939_), .D(new_n12932_), .Y(new_n15143_));
  OAI21  g14141(.A0(new_n14749_), .A1(new_n14777_), .B0(new_n15143_), .Y(new_n15144_));
  NAND3  g14142(.A(new_n14781_), .B(new_n14747_), .C(new_n14741_), .Y(new_n15145_));
  AOI21  g14143(.A0(new_n14770_), .A1(new_n15144_), .B0(new_n15145_), .Y(new_n15146_));
  AOI21  g14144(.A0(new_n15142_), .A1(new_n14708_), .B0(new_n15146_), .Y(new_n15147_));
  AOI22  g14145(.A0(new_n12951_), .A1(new_n12948_), .B0(new_n12930_), .B1(new_n12927_), .Y(new_n15148_));
  OAI221 g14146(.A0(new_n14767_), .A1(new_n14759_), .C0(new_n15148_), .B0(new_n14764_), .B1(new_n14751_), .Y(new_n15149_));
  AOI22  g14147(.A0(new_n15149_), .A1(new_n15144_), .B0(new_n14769_), .B1(new_n14766_), .Y(new_n15150_));
  AOI22  g14148(.A0(new_n13002_), .A1(new_n12991_), .B0(new_n14734_), .B1(new_n12975_), .Y(new_n15151_));
  OAI221 g14149(.A0(new_n14737_), .A1(new_n12988_), .C0(new_n15151_), .B0(new_n14733_), .B1(new_n12973_), .Y(new_n15152_));
  OAI21  g14150(.A0(new_n14732_), .A1(new_n14723_), .B0(new_n15152_), .Y(new_n15153_));
  NAND2  g14151(.A(new_n14739_), .B(new_n14736_), .Y(new_n15154_));
  NAND2  g14152(.A(new_n15154_), .B(new_n15153_), .Y(new_n15155_));
  XOR2   g14153(.A(new_n15155_), .B(new_n15150_), .Y(new_n15156_));
  NAND4  g14154(.A(new_n14781_), .B(new_n14771_), .C(new_n14747_), .D(new_n14741_), .Y(new_n15157_));
  OAI21  g14155(.A0(new_n14763_), .A1(new_n14750_), .B0(new_n15149_), .Y(new_n15158_));
  NAND2  g14156(.A(new_n14769_), .B(new_n14766_), .Y(new_n15159_));
  NAND2  g14157(.A(new_n15159_), .B(new_n15158_), .Y(new_n15160_));
  OAI211 g14158(.A0(new_n12979_), .A1(new_n12973_), .B0(new_n14721_), .B1(new_n12982_), .Y(new_n15161_));
  OAI22  g14159(.A0(new_n15161_), .A1(new_n12996_), .B0(new_n14743_), .B1(new_n12968_), .Y(new_n15162_));
  AOI22  g14160(.A0(new_n15152_), .A1(new_n15162_), .B0(new_n14739_), .B1(new_n14736_), .Y(new_n15163_));
  NAND2  g14161(.A(new_n15163_), .B(new_n15160_), .Y(new_n15164_));
  NAND2  g14162(.A(new_n15155_), .B(new_n15150_), .Y(new_n15165_));
  NAND3  g14163(.A(new_n15165_), .B(new_n15164_), .C(new_n15157_), .Y(new_n15166_));
  OAI22  g14164(.A0(new_n15166_), .A1(new_n15141_), .B0(new_n15156_), .B1(new_n15147_), .Y(new_n15167_));
  NOR2   g14165(.A(new_n12073_), .B(new_n12000_), .Y(new_n15168_));
  NAND2  g14166(.A(new_n12073_), .B(new_n12000_), .Y(new_n15169_));
  OAI21  g14167(.A0(new_n15168_), .A1(new_n15113_), .B0(new_n15169_), .Y(new_n15170_));
  XOR2   g14168(.A(new_n13076_), .B(new_n14698_), .Y(new_n15171_));
  XOR2   g14169(.A(new_n13126_), .B(new_n14657_), .Y(new_n15172_));
  NAND2  g14170(.A(new_n15172_), .B(new_n15171_), .Y(new_n15173_));
  NOR2   g14171(.A(new_n15172_), .B(new_n15171_), .Y(new_n15174_));
  AOI21  g14172(.A0(new_n15173_), .A1(new_n15170_), .B0(new_n15174_), .Y(new_n15175_));
  AOI22  g14173(.A0(new_n14702_), .A1(new_n14692_), .B0(new_n14668_), .B1(new_n14654_), .Y(new_n15176_));
  NOR2   g14174(.A(new_n15176_), .B(new_n15175_), .Y(new_n15177_));
  NAND2  g14175(.A(new_n14703_), .B(new_n14669_), .Y(new_n15178_));
  NAND4  g14176(.A(new_n13074_), .B(new_n13065_), .C(new_n13051_), .D(new_n13044_), .Y(new_n15179_));
  OAI21  g14177(.A0(new_n14670_), .A1(new_n14698_), .B0(new_n15179_), .Y(new_n15180_));
  NAND3  g14178(.A(new_n14702_), .B(new_n14668_), .C(new_n14654_), .Y(new_n15181_));
  AOI21  g14179(.A0(new_n14691_), .A1(new_n15180_), .B0(new_n15181_), .Y(new_n15182_));
  AOI21  g14180(.A0(new_n15178_), .A1(new_n14629_), .B0(new_n15182_), .Y(new_n15183_));
  AOI22  g14181(.A0(new_n13063_), .A1(new_n13060_), .B0(new_n13042_), .B1(new_n13039_), .Y(new_n15184_));
  OAI221 g14182(.A0(new_n14688_), .A1(new_n14680_), .C0(new_n15184_), .B0(new_n14685_), .B1(new_n14672_), .Y(new_n15185_));
  AOI22  g14183(.A0(new_n15185_), .A1(new_n15180_), .B0(new_n14690_), .B1(new_n14687_), .Y(new_n15186_));
  AOI22  g14184(.A0(new_n14640_), .A1(new_n13117_), .B0(new_n13101_), .B1(new_n13105_), .Y(new_n15187_));
  OAI221 g14185(.A0(new_n14650_), .A1(new_n13114_), .C0(new_n15187_), .B0(new_n14647_), .B1(new_n13094_), .Y(new_n15188_));
  OAI21  g14186(.A0(new_n14646_), .A1(new_n14630_), .B0(new_n15188_), .Y(new_n15189_));
  NAND2  g14187(.A(new_n14652_), .B(new_n14649_), .Y(new_n15190_));
  NAND2  g14188(.A(new_n15190_), .B(new_n15189_), .Y(new_n15191_));
  XOR2   g14189(.A(new_n15191_), .B(new_n15186_), .Y(new_n15192_));
  NAND4  g14190(.A(new_n14702_), .B(new_n14692_), .C(new_n14668_), .D(new_n14654_), .Y(new_n15193_));
  OAI21  g14191(.A0(new_n14684_), .A1(new_n14671_), .B0(new_n15185_), .Y(new_n15194_));
  NAND2  g14192(.A(new_n14690_), .B(new_n14687_), .Y(new_n15195_));
  NAND2  g14193(.A(new_n15195_), .B(new_n15194_), .Y(new_n15196_));
  NAND4  g14194(.A(new_n13124_), .B(new_n14663_), .C(new_n13108_), .D(new_n14660_), .Y(new_n15197_));
  OAI21  g14195(.A0(new_n14664_), .A1(new_n14657_), .B0(new_n15197_), .Y(new_n15198_));
  AOI22  g14196(.A0(new_n15188_), .A1(new_n15198_), .B0(new_n14652_), .B1(new_n14649_), .Y(new_n15199_));
  NAND2  g14197(.A(new_n15199_), .B(new_n15196_), .Y(new_n15200_));
  NAND2  g14198(.A(new_n15191_), .B(new_n15186_), .Y(new_n15201_));
  NAND3  g14199(.A(new_n15201_), .B(new_n15200_), .C(new_n15193_), .Y(new_n15202_));
  OAI22  g14200(.A0(new_n15202_), .A1(new_n15177_), .B0(new_n15192_), .B1(new_n15183_), .Y(new_n15203_));
  XOR2   g14201(.A(new_n15203_), .B(new_n15167_), .Y(new_n15204_));
  XOR2   g14202(.A(new_n15204_), .B(new_n15133_), .Y(new_n15205_));
  NOR2   g14203(.A(new_n14612_), .B(new_n14525_), .Y(new_n15206_));
  NAND2  g14204(.A(new_n14612_), .B(new_n14525_), .Y(new_n15207_));
  OAI21  g14205(.A0(new_n15206_), .A1(new_n15126_), .B0(new_n15207_), .Y(new_n15208_));
  XOR2   g14206(.A(new_n13199_), .B(new_n14605_), .Y(new_n15209_));
  NAND2  g14207(.A(new_n14546_), .B(new_n14545_), .Y(new_n15210_));
  XOR2   g14208(.A(new_n13243_), .B(new_n15210_), .Y(new_n15211_));
  NAND2  g14209(.A(new_n15211_), .B(new_n15209_), .Y(new_n15212_));
  NOR2   g14210(.A(new_n15211_), .B(new_n15209_), .Y(new_n15213_));
  AOI21  g14211(.A0(new_n15212_), .A1(new_n13142_), .B0(new_n15213_), .Y(new_n15214_));
  AOI22  g14212(.A0(new_n14609_), .A1(new_n14599_), .B0(new_n14575_), .B1(new_n14569_), .Y(new_n15215_));
  NOR2   g14213(.A(new_n15215_), .B(new_n15214_), .Y(new_n15216_));
  NAND2  g14214(.A(new_n14610_), .B(new_n14576_), .Y(new_n15217_));
  NAND4  g14215(.A(new_n13197_), .B(new_n13188_), .C(new_n13174_), .D(new_n13167_), .Y(new_n15218_));
  OAI21  g14216(.A0(new_n14577_), .A1(new_n14605_), .B0(new_n15218_), .Y(new_n15219_));
  NAND3  g14217(.A(new_n14609_), .B(new_n14575_), .C(new_n14569_), .Y(new_n15220_));
  AOI21  g14218(.A0(new_n14598_), .A1(new_n15219_), .B0(new_n15220_), .Y(new_n15221_));
  AOI21  g14219(.A0(new_n15217_), .A1(new_n14536_), .B0(new_n15221_), .Y(new_n15222_));
  AOI22  g14220(.A0(new_n13186_), .A1(new_n13183_), .B0(new_n13165_), .B1(new_n13162_), .Y(new_n15223_));
  OAI221 g14221(.A0(new_n14595_), .A1(new_n14587_), .C0(new_n15223_), .B0(new_n14592_), .B1(new_n14579_), .Y(new_n15224_));
  AOI22  g14222(.A0(new_n15224_), .A1(new_n15219_), .B0(new_n14597_), .B1(new_n14594_), .Y(new_n15225_));
  AOI22  g14223(.A0(new_n13237_), .A1(new_n13226_), .B0(new_n14562_), .B1(new_n13210_), .Y(new_n15226_));
  OAI221 g14224(.A0(new_n14565_), .A1(new_n13223_), .C0(new_n15226_), .B0(new_n14561_), .B1(new_n13208_), .Y(new_n15227_));
  OAI21  g14225(.A0(new_n14560_), .A1(new_n14551_), .B0(new_n15227_), .Y(new_n15228_));
  NAND2  g14226(.A(new_n14567_), .B(new_n14564_), .Y(new_n15229_));
  NAND2  g14227(.A(new_n15229_), .B(new_n15228_), .Y(new_n15230_));
  XOR2   g14228(.A(new_n15230_), .B(new_n15225_), .Y(new_n15231_));
  NAND4  g14229(.A(new_n14609_), .B(new_n14599_), .C(new_n14575_), .D(new_n14569_), .Y(new_n15232_));
  OAI21  g14230(.A0(new_n14591_), .A1(new_n14578_), .B0(new_n15224_), .Y(new_n15233_));
  NAND2  g14231(.A(new_n14597_), .B(new_n14594_), .Y(new_n15234_));
  NAND2  g14232(.A(new_n15234_), .B(new_n15233_), .Y(new_n15235_));
  OAI211 g14233(.A0(new_n13214_), .A1(new_n13208_), .B0(new_n14549_), .B1(new_n13217_), .Y(new_n15236_));
  OAI22  g14234(.A0(new_n15236_), .A1(new_n13231_), .B0(new_n14571_), .B1(new_n13203_), .Y(new_n15237_));
  AOI22  g14235(.A0(new_n15227_), .A1(new_n15237_), .B0(new_n14567_), .B1(new_n14564_), .Y(new_n15238_));
  NAND2  g14236(.A(new_n15238_), .B(new_n15235_), .Y(new_n15239_));
  NAND2  g14237(.A(new_n15230_), .B(new_n15225_), .Y(new_n15240_));
  NAND3  g14238(.A(new_n15240_), .B(new_n15239_), .C(new_n15232_), .Y(new_n15241_));
  OAI22  g14239(.A0(new_n15241_), .A1(new_n15216_), .B0(new_n15231_), .B1(new_n15222_), .Y(new_n15242_));
  XOR2   g14240(.A(new_n13320_), .B(new_n14518_), .Y(new_n15243_));
  XOR2   g14241(.A(new_n13370_), .B(new_n14484_), .Y(new_n15244_));
  NAND2  g14242(.A(new_n15244_), .B(new_n15243_), .Y(new_n15245_));
  NOR2   g14243(.A(new_n15244_), .B(new_n15243_), .Y(new_n15246_));
  AOI21  g14244(.A0(new_n15245_), .A1(new_n14449_), .B0(new_n15246_), .Y(new_n15247_));
  AOI22  g14245(.A0(new_n14522_), .A1(new_n14515_), .B0(new_n14495_), .B1(new_n14481_), .Y(new_n15248_));
  NOR2   g14246(.A(new_n15248_), .B(new_n15247_), .Y(new_n15249_));
  NAND2  g14247(.A(new_n14523_), .B(new_n14496_), .Y(new_n15250_));
  NAND4  g14248(.A(new_n13318_), .B(new_n13309_), .C(new_n13294_), .D(new_n13285_), .Y(new_n15251_));
  OAI21  g14249(.A0(new_n14497_), .A1(new_n14518_), .B0(new_n15251_), .Y(new_n15252_));
  NAND3  g14250(.A(new_n14522_), .B(new_n14495_), .C(new_n14481_), .Y(new_n15253_));
  AOI21  g14251(.A0(new_n14514_), .A1(new_n15252_), .B0(new_n15253_), .Y(new_n15254_));
  AOI21  g14252(.A0(new_n15250_), .A1(new_n14456_), .B0(new_n15254_), .Y(new_n15255_));
  AOI22  g14253(.A0(new_n13307_), .A1(new_n13304_), .B0(new_n13283_), .B1(new_n13280_), .Y(new_n15256_));
  OAI221 g14254(.A0(new_n14511_), .A1(new_n14503_), .C0(new_n15256_), .B0(new_n14508_), .B1(new_n14499_), .Y(new_n15257_));
  AOI22  g14255(.A0(new_n15257_), .A1(new_n15252_), .B0(new_n14513_), .B1(new_n14510_), .Y(new_n15258_));
  AOI22  g14256(.A0(new_n14467_), .A1(new_n13361_), .B0(new_n13345_), .B1(new_n13349_), .Y(new_n15259_));
  OAI221 g14257(.A0(new_n14477_), .A1(new_n13358_), .C0(new_n15259_), .B0(new_n14474_), .B1(new_n13338_), .Y(new_n15260_));
  OAI21  g14258(.A0(new_n14473_), .A1(new_n14457_), .B0(new_n15260_), .Y(new_n15261_));
  NAND2  g14259(.A(new_n14479_), .B(new_n14476_), .Y(new_n15262_));
  NAND2  g14260(.A(new_n15262_), .B(new_n15261_), .Y(new_n15263_));
  XOR2   g14261(.A(new_n15263_), .B(new_n15258_), .Y(new_n15264_));
  NAND4  g14262(.A(new_n14522_), .B(new_n14515_), .C(new_n14495_), .D(new_n14481_), .Y(new_n15265_));
  OAI21  g14263(.A0(new_n14507_), .A1(new_n14498_), .B0(new_n15257_), .Y(new_n15266_));
  NAND2  g14264(.A(new_n14513_), .B(new_n14510_), .Y(new_n15267_));
  NAND2  g14265(.A(new_n15267_), .B(new_n15266_), .Y(new_n15268_));
  NAND4  g14266(.A(new_n13368_), .B(new_n14490_), .C(new_n13352_), .D(new_n14487_), .Y(new_n15269_));
  OAI21  g14267(.A0(new_n14491_), .A1(new_n14484_), .B0(new_n15269_), .Y(new_n15270_));
  AOI22  g14268(.A0(new_n15260_), .A1(new_n15270_), .B0(new_n14479_), .B1(new_n14476_), .Y(new_n15271_));
  NAND2  g14269(.A(new_n15271_), .B(new_n15268_), .Y(new_n15272_));
  NAND2  g14270(.A(new_n15263_), .B(new_n15258_), .Y(new_n15273_));
  NAND3  g14271(.A(new_n15273_), .B(new_n15272_), .C(new_n15265_), .Y(new_n15274_));
  OAI22  g14272(.A0(new_n15274_), .A1(new_n15249_), .B0(new_n15264_), .B1(new_n15255_), .Y(new_n15275_));
  XOR2   g14273(.A(new_n15275_), .B(new_n15242_), .Y(new_n15276_));
  XOR2   g14274(.A(new_n15276_), .B(new_n15208_), .Y(new_n15277_));
  XOR2   g14275(.A(new_n15277_), .B(new_n15205_), .Y(new_n15278_));
  XOR2   g14276(.A(new_n15278_), .B(new_n15130_), .Y(new_n15279_));
  NOR2   g14277(.A(new_n14435_), .B(new_n14431_), .Y(new_n15280_));
  OAI21  g14278(.A0(new_n15280_), .A1(new_n14362_), .B0(new_n14429_), .Y(new_n15281_));
  NOR2   g14279(.A(new_n13688_), .B(new_n13622_), .Y(new_n15282_));
  NAND2  g14280(.A(new_n13688_), .B(new_n13622_), .Y(new_n15283_));
  OAI21  g14281(.A0(new_n15282_), .A1(new_n14239_), .B0(new_n15283_), .Y(new_n15284_));
  XOR2   g14282(.A(new_n14428_), .B(new_n15284_), .Y(new_n15285_));
  OAI21  g14283(.A0(new_n14435_), .A1(new_n14431_), .B0(new_n15285_), .Y(new_n15286_));
  NOR2   g14284(.A(new_n15286_), .B(new_n14362_), .Y(new_n15287_));
  AOI21  g14285(.A0(new_n15281_), .A1(new_n15105_), .B0(new_n15287_), .Y(new_n15288_));
  INV    g14286(.A(new_n14340_), .Y(new_n15289_));
  OAI21  g14287(.A0(new_n14337_), .A1(new_n14248_), .B0(new_n15289_), .Y(new_n15290_));
  AOI22  g14288(.A0(new_n13529_), .A1(new_n14347_), .B0(new_n13503_), .B1(new_n13499_), .Y(new_n15291_));
  OAI211 g14289(.A0(new_n14348_), .A1(new_n13523_), .B0(new_n15291_), .B1(new_n14342_), .Y(new_n15292_));
  NAND2  g14290(.A(new_n15292_), .B(new_n15290_), .Y(new_n15293_));
  NAND2  g14291(.A(new_n14350_), .B(new_n14344_), .Y(new_n15294_));
  NAND2  g14292(.A(new_n15294_), .B(new_n15293_), .Y(new_n15295_));
  AOI22  g14293(.A0(new_n14318_), .A1(new_n14307_), .B0(new_n14275_), .B1(new_n14271_), .Y(new_n15296_));
  NOR2   g14294(.A(new_n15296_), .B(new_n14325_), .Y(new_n15297_));
  NAND2  g14295(.A(new_n14319_), .B(new_n14276_), .Y(new_n15298_));
  NAND4  g14296(.A(new_n13429_), .B(new_n14313_), .C(new_n13413_), .D(new_n14310_), .Y(new_n15299_));
  OAI21  g14297(.A0(new_n14314_), .A1(new_n13548_), .B0(new_n15299_), .Y(new_n15300_));
  NAND3  g14298(.A(new_n14318_), .B(new_n14275_), .C(new_n14271_), .Y(new_n15301_));
  AOI21  g14299(.A0(new_n14306_), .A1(new_n15300_), .B0(new_n15301_), .Y(new_n15302_));
  AOI21  g14300(.A0(new_n15298_), .A1(new_n14255_), .B0(new_n15302_), .Y(new_n15303_));
  AOI22  g14301(.A0(new_n14292_), .A1(new_n13422_), .B0(new_n14300_), .B1(new_n13406_), .Y(new_n15304_));
  OAI221 g14302(.A0(new_n14303_), .A1(new_n13419_), .C0(new_n15304_), .B0(new_n14299_), .B1(new_n13404_), .Y(new_n15305_));
  AOI22  g14303(.A0(new_n15305_), .A1(new_n15300_), .B0(new_n14305_), .B1(new_n14302_), .Y(new_n15306_));
  OAI21  g14304(.A0(new_n14265_), .A1(new_n14264_), .B0(new_n14259_), .Y(new_n15307_));
  NAND3  g14305(.A(new_n14268_), .B(new_n14267_), .C(new_n13450_), .Y(new_n15308_));
  OAI21  g14306(.A0(new_n14258_), .A1(new_n14256_), .B0(new_n15308_), .Y(new_n15309_));
  NAND2  g14307(.A(new_n15309_), .B(new_n15307_), .Y(new_n15310_));
  XOR2   g14308(.A(new_n15310_), .B(new_n15306_), .Y(new_n15311_));
  NAND4  g14309(.A(new_n14318_), .B(new_n14307_), .C(new_n14275_), .D(new_n14271_), .Y(new_n15312_));
  OAI21  g14310(.A0(new_n14298_), .A1(new_n14277_), .B0(new_n15305_), .Y(new_n15313_));
  NAND2  g14311(.A(new_n14305_), .B(new_n14302_), .Y(new_n15314_));
  NAND2  g14312(.A(new_n15314_), .B(new_n15313_), .Y(new_n15315_));
  AOI21  g14313(.A0(new_n15308_), .A1(new_n14326_), .B0(new_n14269_), .Y(new_n15316_));
  NAND2  g14314(.A(new_n15316_), .B(new_n15315_), .Y(new_n15317_));
  NAND2  g14315(.A(new_n15310_), .B(new_n15306_), .Y(new_n15318_));
  NAND3  g14316(.A(new_n15318_), .B(new_n15317_), .C(new_n15312_), .Y(new_n15319_));
  OAI22  g14317(.A0(new_n15319_), .A1(new_n15297_), .B0(new_n15311_), .B1(new_n15303_), .Y(new_n15320_));
  NOR2   g14318(.A(new_n14434_), .B(new_n14359_), .Y(new_n15321_));
  NAND3  g14319(.A(new_n14359_), .B(new_n14330_), .C(new_n14321_), .Y(new_n15322_));
  AOI22  g14320(.A0(new_n15292_), .A1(new_n15290_), .B0(new_n14350_), .B1(new_n14344_), .Y(new_n15323_));
  OAI221 g14321(.A0(new_n15319_), .A1(new_n15297_), .C0(new_n15323_), .B0(new_n15311_), .B1(new_n15303_), .Y(new_n15324_));
  OAI211 g14322(.A0(new_n15321_), .A1(new_n14252_), .B0(new_n15324_), .B1(new_n15322_), .Y(new_n15325_));
  AOI21  g14323(.A0(new_n15320_), .A1(new_n15295_), .B0(new_n15325_), .Y(new_n15326_));
  OAI21  g14324(.A0(new_n15321_), .A1(new_n14252_), .B0(new_n15322_), .Y(new_n15327_));
  NAND2  g14325(.A(new_n15320_), .B(new_n15295_), .Y(new_n15328_));
  OAI21  g14326(.A0(new_n15296_), .A1(new_n14325_), .B0(new_n15312_), .Y(new_n15329_));
  XOR2   g14327(.A(new_n15310_), .B(new_n15315_), .Y(new_n15330_));
  OAI21  g14328(.A0(new_n15310_), .A1(new_n15306_), .B0(new_n15312_), .Y(new_n15331_));
  AOI221 g14329(.A0(new_n15310_), .A1(new_n15306_), .C0(new_n15331_), .B0(new_n15298_), .B1(new_n14255_), .Y(new_n15332_));
  AOI21  g14330(.A0(new_n15330_), .A1(new_n15329_), .B0(new_n15332_), .Y(new_n15333_));
  OAI21  g14331(.A0(new_n15333_), .A1(new_n15323_), .B0(new_n15324_), .Y(new_n15334_));
  NAND2  g14332(.A(new_n14360_), .B(new_n14355_), .Y(new_n15335_));
  NOR2   g14333(.A(new_n14320_), .B(new_n14255_), .Y(new_n15336_));
  NOR3   g14334(.A(new_n14355_), .B(new_n15336_), .C(new_n14432_), .Y(new_n15337_));
  AOI211 g14335(.A0(new_n15330_), .A1(new_n15329_), .B(new_n15295_), .C(new_n15332_), .Y(new_n15338_));
  AOI211 g14336(.A0(new_n15335_), .A1(new_n14431_), .B(new_n15338_), .C(new_n15337_), .Y(new_n15339_));
  AOI22  g14337(.A0(new_n15339_), .A1(new_n15328_), .B0(new_n15334_), .B1(new_n15327_), .Y(new_n15340_));
  NAND4  g14338(.A(new_n13685_), .B(new_n14394_), .C(new_n13660_), .D(new_n14391_), .Y(new_n15341_));
  OAI21  g14339(.A0(new_n14395_), .A1(new_n14369_), .B0(new_n15341_), .Y(new_n15342_));
  NAND2  g14340(.A(new_n14387_), .B(new_n15342_), .Y(new_n15343_));
  NAND4  g14341(.A(new_n13619_), .B(new_n13615_), .C(new_n13591_), .D(new_n13588_), .Y(new_n15344_));
  OAI21  g14342(.A0(new_n14422_), .A1(new_n14365_), .B0(new_n15344_), .Y(new_n15345_));
  NAND2  g14343(.A(new_n14420_), .B(new_n15345_), .Y(new_n15346_));
  AOI22  g14344(.A0(new_n14426_), .A1(new_n15346_), .B0(new_n14399_), .B1(new_n15343_), .Y(new_n15347_));
  NOR2   g14345(.A(new_n15347_), .B(new_n14373_), .Y(new_n15348_));
  NAND2  g14346(.A(new_n14427_), .B(new_n14400_), .Y(new_n15349_));
  OAI211 g14347(.A0(new_n14388_), .A1(new_n14380_), .B0(new_n14426_), .B1(new_n14399_), .Y(new_n15350_));
  AOI21  g14348(.A0(new_n14420_), .A1(new_n15345_), .B0(new_n15350_), .Y(new_n15351_));
  AOI21  g14349(.A0(new_n15349_), .A1(new_n15284_), .B0(new_n15351_), .Y(new_n15352_));
  AOI22  g14350(.A0(new_n13606_), .A1(new_n13610_), .B0(new_n13579_), .B1(new_n13583_), .Y(new_n15353_));
  OAI221 g14351(.A0(new_n14417_), .A1(new_n14406_), .C0(new_n15353_), .B0(new_n14414_), .B1(new_n14402_), .Y(new_n15354_));
  AOI22  g14352(.A0(new_n15354_), .A1(new_n15345_), .B0(new_n14419_), .B1(new_n14416_), .Y(new_n15355_));
  AOI22  g14353(.A0(new_n13682_), .A1(new_n13669_), .B0(new_n13657_), .B1(new_n13644_), .Y(new_n15356_));
  OAI221 g14354(.A0(new_n14384_), .A1(new_n13666_), .C0(new_n15356_), .B0(new_n14381_), .B1(new_n13641_), .Y(new_n15357_));
  INV    g14355(.A(new_n15357_), .Y(new_n15358_));
  NAND2  g14356(.A(new_n14386_), .B(new_n14383_), .Y(new_n15359_));
  OAI21  g14357(.A0(new_n15358_), .A1(new_n14380_), .B0(new_n15359_), .Y(new_n15360_));
  XOR2   g14358(.A(new_n15360_), .B(new_n15355_), .Y(new_n15361_));
  NAND4  g14359(.A(new_n14426_), .B(new_n15346_), .C(new_n14399_), .D(new_n15343_), .Y(new_n15362_));
  INV    g14360(.A(new_n15354_), .Y(new_n15363_));
  NAND2  g14361(.A(new_n14419_), .B(new_n14416_), .Y(new_n15364_));
  OAI21  g14362(.A0(new_n15363_), .A1(new_n14413_), .B0(new_n15364_), .Y(new_n15365_));
  OAI211 g14363(.A0(new_n15358_), .A1(new_n14380_), .B0(new_n15359_), .B1(new_n15365_), .Y(new_n15366_));
  NAND2  g14364(.A(new_n15360_), .B(new_n15355_), .Y(new_n15367_));
  NAND3  g14365(.A(new_n15367_), .B(new_n15366_), .C(new_n15362_), .Y(new_n15368_));
  OAI22  g14366(.A0(new_n15368_), .A1(new_n15348_), .B0(new_n15361_), .B1(new_n15352_), .Y(new_n15369_));
  AOI21  g14367(.A0(new_n15335_), .A1(new_n14431_), .B0(new_n15337_), .Y(new_n15370_));
  AOI21  g14368(.A0(new_n15320_), .A1(new_n15295_), .B0(new_n15338_), .Y(new_n15371_));
  OAI21  g14369(.A0(new_n15371_), .A1(new_n15370_), .B0(new_n15369_), .Y(new_n15372_));
  OAI22  g14370(.A0(new_n15372_), .A1(new_n15326_), .B0(new_n15369_), .B1(new_n15340_), .Y(new_n15373_));
  XOR2   g14371(.A(new_n15373_), .B(new_n15288_), .Y(new_n15374_));
  XOR2   g14372(.A(new_n15374_), .B(new_n15279_), .Y(new_n15375_));
  NOR2   g14373(.A(new_n15375_), .B(new_n15112_), .Y(new_n15376_));
  XOR2   g14374(.A(new_n14787_), .B(new_n15122_), .Y(new_n15377_));
  NAND2  g14375(.A(new_n15377_), .B(new_n14439_), .Y(new_n15378_));
  NOR2   g14376(.A(new_n15377_), .B(new_n14439_), .Y(new_n15379_));
  AOI21  g14377(.A0(new_n15378_), .A1(new_n14793_), .B0(new_n15379_), .Y(new_n15380_));
  XOR2   g14378(.A(new_n13128_), .B(new_n15170_), .Y(new_n15381_));
  NOR2   g14379(.A(new_n15381_), .B(new_n13011_), .Y(new_n15382_));
  NAND2  g14380(.A(new_n15381_), .B(new_n13011_), .Y(new_n15383_));
  OAI21  g14381(.A0(new_n15382_), .A1(new_n15118_), .B0(new_n15383_), .Y(new_n15384_));
  XOR2   g14382(.A(new_n14785_), .B(new_n15384_), .Y(new_n15385_));
  NOR2   g14383(.A(new_n15385_), .B(new_n14614_), .Y(new_n15386_));
  NAND2  g14384(.A(new_n15385_), .B(new_n14614_), .Y(new_n15387_));
  OAI21  g14385(.A0(new_n15386_), .A1(new_n14446_), .B0(new_n15387_), .Y(new_n15388_));
  XOR2   g14386(.A(new_n15278_), .B(new_n15388_), .Y(new_n15389_));
  XOR2   g14387(.A(new_n15374_), .B(new_n15389_), .Y(new_n15390_));
  XOR2   g14388(.A(new_n15390_), .B(new_n15380_), .Y(new_n15391_));
  XOR2   g14389(.A(new_n12395_), .B(new_n14093_), .Y(new_n15392_));
  AOI21  g14390(.A0(new_n4162_), .A1(new_n4153_), .B0(new_n4155_), .Y(new_n15393_));
  XOR2   g14391(.A(new_n12550_), .B(new_n15393_), .Y(new_n15394_));
  NAND2  g14392(.A(new_n15394_), .B(new_n15392_), .Y(new_n15395_));
  NOR2   g14393(.A(new_n15394_), .B(new_n15392_), .Y(new_n15396_));
  AOI21  g14394(.A0(new_n15395_), .A1(new_n12241_), .B0(new_n15396_), .Y(new_n15397_));
  NOR2   g14395(.A(new_n12549_), .B(new_n12477_), .Y(new_n15398_));
  NAND2  g14396(.A(new_n12549_), .B(new_n12477_), .Y(new_n15399_));
  OAI21  g14397(.A0(new_n15398_), .A1(new_n15393_), .B0(new_n15399_), .Y(new_n15400_));
  XOR2   g14398(.A(new_n14091_), .B(new_n15400_), .Y(new_n15401_));
  NOR2   g14399(.A(new_n14221_), .B(new_n15401_), .Y(new_n15402_));
  NAND2  g14400(.A(new_n14221_), .B(new_n15401_), .Y(new_n15403_));
  OAI21  g14401(.A0(new_n15402_), .A1(new_n15397_), .B0(new_n15403_), .Y(new_n15404_));
  XOR2   g14402(.A(new_n14943_), .B(new_n15404_), .Y(new_n15405_));
  NOR2   g14403(.A(new_n12712_), .B(new_n12635_), .Y(new_n15406_));
  NAND2  g14404(.A(new_n12712_), .B(new_n12635_), .Y(new_n15407_));
  OAI21  g14405(.A0(new_n15406_), .A1(new_n13717_), .B0(new_n15407_), .Y(new_n15408_));
  XOR2   g14406(.A(new_n13950_), .B(new_n15408_), .Y(new_n15409_));
  NOR2   g14407(.A(new_n15409_), .B(new_n13829_), .Y(new_n15410_));
  NAND2  g14408(.A(new_n15409_), .B(new_n13829_), .Y(new_n15411_));
  OAI21  g14409(.A0(new_n15410_), .A1(new_n13723_), .B0(new_n15411_), .Y(new_n15412_));
  XOR2   g14410(.A(new_n15097_), .B(new_n15412_), .Y(new_n15413_));
  NOR2   g14411(.A(new_n15413_), .B(new_n15405_), .Y(new_n15414_));
  NAND2  g14412(.A(new_n15413_), .B(new_n15405_), .Y(new_n15415_));
  OAI21  g14413(.A0(new_n15414_), .A1(new_n14804_), .B0(new_n15415_), .Y(new_n15416_));
  NOR2   g14414(.A(new_n15096_), .B(new_n15024_), .Y(new_n15417_));
  NAND2  g14415(.A(new_n15096_), .B(new_n15024_), .Y(new_n15418_));
  OAI21  g14416(.A0(new_n15417_), .A1(new_n14958_), .B0(new_n15418_), .Y(new_n15419_));
  XOR2   g14417(.A(new_n13776_), .B(new_n15089_), .Y(new_n15420_));
  NAND2  g14418(.A(new_n15034_), .B(new_n15033_), .Y(new_n15421_));
  XOR2   g14419(.A(new_n13826_), .B(new_n15421_), .Y(new_n15422_));
  NAND2  g14420(.A(new_n15422_), .B(new_n15420_), .Y(new_n15423_));
  NOR2   g14421(.A(new_n15422_), .B(new_n15420_), .Y(new_n15424_));
  AOI21  g14422(.A0(new_n15423_), .A1(new_n13726_), .B0(new_n15424_), .Y(new_n15425_));
  AOI22  g14423(.A0(new_n15093_), .A1(new_n15083_), .B0(new_n15061_), .B1(new_n15055_), .Y(new_n15426_));
  NOR2   g14424(.A(new_n15426_), .B(new_n15425_), .Y(new_n15427_));
  NAND2  g14425(.A(new_n15094_), .B(new_n15062_), .Y(new_n15428_));
  OAI22  g14426(.A0(new_n15073_), .A1(new_n15072_), .B0(new_n15070_), .B1(new_n15089_), .Y(new_n15429_));
  NAND3  g14427(.A(new_n15093_), .B(new_n15061_), .C(new_n15055_), .Y(new_n15430_));
  AOI21  g14428(.A0(new_n15082_), .A1(new_n15429_), .B0(new_n15430_), .Y(new_n15431_));
  AOI21  g14429(.A0(new_n15428_), .A1(new_n15027_), .B0(new_n15431_), .Y(new_n15432_));
  AOI22  g14430(.A0(new_n13766_), .A1(new_n13771_), .B0(new_n13743_), .B1(new_n13740_), .Y(new_n15433_));
  OAI221 g14431(.A0(new_n15079_), .A1(new_n13762_), .C0(new_n15433_), .B0(new_n15076_), .B1(new_n15075_), .Y(new_n15434_));
  AOI22  g14432(.A0(new_n15434_), .A1(new_n15429_), .B0(new_n15081_), .B1(new_n15078_), .Y(new_n15435_));
  AOI22  g14433(.A0(new_n13822_), .A1(new_n13807_), .B0(new_n15048_), .B1(new_n13792_), .Y(new_n15436_));
  OAI221 g14434(.A0(new_n15051_), .A1(new_n13804_), .C0(new_n15436_), .B0(new_n15047_), .B1(new_n13789_), .Y(new_n15437_));
  OAI21  g14435(.A0(new_n15046_), .A1(new_n15039_), .B0(new_n15437_), .Y(new_n15438_));
  NAND2  g14436(.A(new_n15053_), .B(new_n15050_), .Y(new_n15439_));
  NAND2  g14437(.A(new_n15439_), .B(new_n15438_), .Y(new_n15440_));
  XOR2   g14438(.A(new_n15440_), .B(new_n15435_), .Y(new_n15441_));
  NAND4  g14439(.A(new_n15093_), .B(new_n15083_), .C(new_n15061_), .D(new_n15055_), .Y(new_n15442_));
  OAI21  g14440(.A0(new_n15074_), .A1(new_n15071_), .B0(new_n15434_), .Y(new_n15443_));
  NAND2  g14441(.A(new_n15081_), .B(new_n15078_), .Y(new_n15444_));
  NAND2  g14442(.A(new_n15444_), .B(new_n15443_), .Y(new_n15445_));
  OAI211 g14443(.A0(new_n13795_), .A1(new_n13789_), .B0(new_n15037_), .B1(new_n13798_), .Y(new_n15446_));
  OAI22  g14444(.A0(new_n15446_), .A1(new_n13812_), .B0(new_n15057_), .B1(new_n13780_), .Y(new_n15447_));
  AOI22  g14445(.A0(new_n15437_), .A1(new_n15447_), .B0(new_n15053_), .B1(new_n15050_), .Y(new_n15448_));
  NAND2  g14446(.A(new_n15448_), .B(new_n15445_), .Y(new_n15449_));
  NAND2  g14447(.A(new_n15440_), .B(new_n15435_), .Y(new_n15450_));
  NAND3  g14448(.A(new_n15450_), .B(new_n15449_), .C(new_n15442_), .Y(new_n15451_));
  OAI22  g14449(.A0(new_n15451_), .A1(new_n15427_), .B0(new_n15441_), .B1(new_n15432_), .Y(new_n15452_));
  XOR2   g14450(.A(new_n13889_), .B(new_n15017_), .Y(new_n15453_));
  XOR2   g14451(.A(new_n13948_), .B(new_n14978_), .Y(new_n15454_));
  NAND2  g14452(.A(new_n15454_), .B(new_n15453_), .Y(new_n15455_));
  NOR2   g14453(.A(new_n15454_), .B(new_n15453_), .Y(new_n15456_));
  AOI21  g14454(.A0(new_n15455_), .A1(new_n15408_), .B0(new_n15456_), .Y(new_n15457_));
  AOI22  g14455(.A0(new_n15021_), .A1(new_n15011_), .B0(new_n14989_), .B1(new_n14976_), .Y(new_n15458_));
  NOR2   g14456(.A(new_n15458_), .B(new_n15457_), .Y(new_n15459_));
  NAND2  g14457(.A(new_n15022_), .B(new_n14990_), .Y(new_n15460_));
  OAI22  g14458(.A0(new_n15001_), .A1(new_n15000_), .B0(new_n14998_), .B1(new_n15017_), .Y(new_n15461_));
  NAND3  g14459(.A(new_n15021_), .B(new_n14989_), .C(new_n14976_), .Y(new_n15462_));
  AOI21  g14460(.A0(new_n15010_), .A1(new_n15461_), .B0(new_n15462_), .Y(new_n15463_));
  AOI21  g14461(.A0(new_n15460_), .A1(new_n14961_), .B0(new_n15463_), .Y(new_n15464_));
  AOI22  g14462(.A0(new_n13879_), .A1(new_n13884_), .B0(new_n13856_), .B1(new_n13853_), .Y(new_n15465_));
  OAI221 g14463(.A0(new_n15007_), .A1(new_n13875_), .C0(new_n15465_), .B0(new_n15004_), .B1(new_n15003_), .Y(new_n15466_));
  AOI22  g14464(.A0(new_n15466_), .A1(new_n15461_), .B0(new_n15009_), .B1(new_n15006_), .Y(new_n15467_));
  AOI22  g14465(.A0(new_n13943_), .A1(new_n13930_), .B0(new_n13912_), .B1(new_n14969_), .Y(new_n15468_));
  OAI221 g14466(.A0(new_n14972_), .A1(new_n13927_), .C0(new_n15468_), .B0(new_n14968_), .B1(new_n13906_), .Y(new_n15469_));
  OAI21  g14467(.A0(new_n14967_), .A1(new_n14962_), .B0(new_n15469_), .Y(new_n15470_));
  NAND2  g14468(.A(new_n14974_), .B(new_n14971_), .Y(new_n15471_));
  NAND2  g14469(.A(new_n15471_), .B(new_n15470_), .Y(new_n15472_));
  XOR2   g14470(.A(new_n15472_), .B(new_n15467_), .Y(new_n15473_));
  NAND4  g14471(.A(new_n15021_), .B(new_n15011_), .C(new_n14989_), .D(new_n14976_), .Y(new_n15474_));
  OAI21  g14472(.A0(new_n15002_), .A1(new_n14999_), .B0(new_n15466_), .Y(new_n15475_));
  NAND2  g14473(.A(new_n15009_), .B(new_n15006_), .Y(new_n15476_));
  NAND2  g14474(.A(new_n15476_), .B(new_n15475_), .Y(new_n15477_));
  NAND4  g14475(.A(new_n13946_), .B(new_n14984_), .C(new_n13921_), .D(new_n14981_), .Y(new_n15478_));
  OAI21  g14476(.A0(new_n14985_), .A1(new_n14978_), .B0(new_n15478_), .Y(new_n15479_));
  AOI22  g14477(.A0(new_n15469_), .A1(new_n15479_), .B0(new_n14974_), .B1(new_n14971_), .Y(new_n15480_));
  NAND2  g14478(.A(new_n15480_), .B(new_n15477_), .Y(new_n15481_));
  NAND2  g14479(.A(new_n15472_), .B(new_n15467_), .Y(new_n15482_));
  NAND3  g14480(.A(new_n15482_), .B(new_n15481_), .C(new_n15474_), .Y(new_n15483_));
  OAI22  g14481(.A0(new_n15483_), .A1(new_n15459_), .B0(new_n15473_), .B1(new_n15464_), .Y(new_n15484_));
  XOR2   g14482(.A(new_n15484_), .B(new_n15452_), .Y(new_n15485_));
  XOR2   g14483(.A(new_n15485_), .B(new_n15419_), .Y(new_n15486_));
  NOR2   g14484(.A(new_n14942_), .B(new_n14879_), .Y(new_n15487_));
  NAND2  g14485(.A(new_n14942_), .B(new_n14879_), .Y(new_n15488_));
  OAI21  g14486(.A0(new_n15487_), .A1(new_n14815_), .B0(new_n15488_), .Y(new_n15489_));
  XOR2   g14487(.A(new_n14030_), .B(new_n14935_), .Y(new_n15490_));
  XOR2   g14488(.A(new_n14089_), .B(new_n14899_), .Y(new_n15491_));
  NAND2  g14489(.A(new_n15491_), .B(new_n15490_), .Y(new_n15492_));
  NOR2   g14490(.A(new_n15491_), .B(new_n15490_), .Y(new_n15493_));
  AOI21  g14491(.A0(new_n15492_), .A1(new_n15400_), .B0(new_n15493_), .Y(new_n15494_));
  AOI22  g14492(.A0(new_n14939_), .A1(new_n14932_), .B0(new_n14910_), .B1(new_n14897_), .Y(new_n15495_));
  NOR2   g14493(.A(new_n15495_), .B(new_n15494_), .Y(new_n15496_));
  NAND2  g14494(.A(new_n14940_), .B(new_n14911_), .Y(new_n15497_));
  NAND4  g14495(.A(new_n14028_), .B(new_n14024_), .C(new_n14000_), .D(new_n13997_), .Y(new_n15498_));
  OAI21  g14496(.A0(new_n14912_), .A1(new_n14935_), .B0(new_n15498_), .Y(new_n15499_));
  NAND3  g14497(.A(new_n14939_), .B(new_n14910_), .C(new_n14897_), .Y(new_n15500_));
  AOI21  g14498(.A0(new_n14931_), .A1(new_n15499_), .B0(new_n15500_), .Y(new_n15501_));
  AOI21  g14499(.A0(new_n15497_), .A1(new_n14882_), .B0(new_n15501_), .Y(new_n15502_));
  AOI22  g14500(.A0(new_n14015_), .A1(new_n14019_), .B0(new_n13988_), .B1(new_n13992_), .Y(new_n15503_));
  OAI221 g14501(.A0(new_n14928_), .A1(new_n14919_), .C0(new_n15503_), .B0(new_n14925_), .B1(new_n14915_), .Y(new_n15504_));
  AOI22  g14502(.A0(new_n15504_), .A1(new_n15499_), .B0(new_n14930_), .B1(new_n14927_), .Y(new_n15505_));
  AOI22  g14503(.A0(new_n14084_), .A1(new_n14071_), .B0(new_n14053_), .B1(new_n14890_), .Y(new_n15506_));
  OAI221 g14504(.A0(new_n14893_), .A1(new_n14068_), .C0(new_n15506_), .B0(new_n14889_), .B1(new_n14047_), .Y(new_n15507_));
  OAI21  g14505(.A0(new_n14888_), .A1(new_n14883_), .B0(new_n15507_), .Y(new_n15508_));
  NAND2  g14506(.A(new_n14895_), .B(new_n14892_), .Y(new_n15509_));
  NAND2  g14507(.A(new_n15509_), .B(new_n15508_), .Y(new_n15510_));
  XOR2   g14508(.A(new_n15510_), .B(new_n15505_), .Y(new_n15511_));
  NAND4  g14509(.A(new_n14939_), .B(new_n14932_), .C(new_n14910_), .D(new_n14897_), .Y(new_n15512_));
  OAI21  g14510(.A0(new_n14924_), .A1(new_n14913_), .B0(new_n15504_), .Y(new_n15513_));
  NAND2  g14511(.A(new_n14930_), .B(new_n14927_), .Y(new_n15514_));
  NAND2  g14512(.A(new_n15514_), .B(new_n15513_), .Y(new_n15515_));
  NAND4  g14513(.A(new_n14087_), .B(new_n14905_), .C(new_n14062_), .D(new_n14902_), .Y(new_n15516_));
  OAI21  g14514(.A0(new_n14906_), .A1(new_n14899_), .B0(new_n15516_), .Y(new_n15517_));
  AOI22  g14515(.A0(new_n15507_), .A1(new_n15517_), .B0(new_n14895_), .B1(new_n14892_), .Y(new_n15518_));
  NAND2  g14516(.A(new_n15518_), .B(new_n15515_), .Y(new_n15519_));
  NAND2  g14517(.A(new_n15510_), .B(new_n15505_), .Y(new_n15520_));
  NAND3  g14518(.A(new_n15520_), .B(new_n15519_), .C(new_n15512_), .Y(new_n15521_));
  OAI22  g14519(.A0(new_n15521_), .A1(new_n15496_), .B0(new_n15511_), .B1(new_n15502_), .Y(new_n15522_));
  XOR2   g14520(.A(new_n14160_), .B(new_n14872_), .Y(new_n15523_));
  XOR2   g14521(.A(new_n14218_), .B(new_n14836_), .Y(new_n15524_));
  NAND2  g14522(.A(new_n15524_), .B(new_n15523_), .Y(new_n15525_));
  NOR2   g14523(.A(new_n15524_), .B(new_n15523_), .Y(new_n15526_));
  AOI21  g14524(.A0(new_n15525_), .A1(new_n14096_), .B0(new_n15526_), .Y(new_n15527_));
  AOI22  g14525(.A0(new_n14876_), .A1(new_n14869_), .B0(new_n14847_), .B1(new_n14834_), .Y(new_n15528_));
  NOR2   g14526(.A(new_n15528_), .B(new_n15527_), .Y(new_n15529_));
  NAND2  g14527(.A(new_n14877_), .B(new_n14848_), .Y(new_n15530_));
  NAND4  g14528(.A(new_n14158_), .B(new_n14154_), .C(new_n14130_), .D(new_n14127_), .Y(new_n15531_));
  OAI21  g14529(.A0(new_n14849_), .A1(new_n14872_), .B0(new_n15531_), .Y(new_n15532_));
  NAND3  g14530(.A(new_n14876_), .B(new_n14847_), .C(new_n14834_), .Y(new_n15533_));
  AOI21  g14531(.A0(new_n14868_), .A1(new_n15532_), .B0(new_n15533_), .Y(new_n15534_));
  AOI21  g14532(.A0(new_n15530_), .A1(new_n14818_), .B0(new_n15534_), .Y(new_n15535_));
  AOI22  g14533(.A0(new_n14145_), .A1(new_n14149_), .B0(new_n14118_), .B1(new_n14122_), .Y(new_n15536_));
  OAI221 g14534(.A0(new_n14865_), .A1(new_n14856_), .C0(new_n15536_), .B0(new_n14862_), .B1(new_n14852_), .Y(new_n15537_));
  AOI22  g14535(.A0(new_n15537_), .A1(new_n15532_), .B0(new_n14867_), .B1(new_n14864_), .Y(new_n15538_));
  AOI22  g14536(.A0(new_n14214_), .A1(new_n14204_), .B0(new_n14186_), .B1(new_n14827_), .Y(new_n15539_));
  OAI221 g14537(.A0(new_n14830_), .A1(new_n14201_), .C0(new_n15539_), .B0(new_n14826_), .B1(new_n14180_), .Y(new_n15540_));
  OAI21  g14538(.A0(new_n14825_), .A1(new_n14819_), .B0(new_n15540_), .Y(new_n15541_));
  NAND2  g14539(.A(new_n14832_), .B(new_n14829_), .Y(new_n15542_));
  NAND2  g14540(.A(new_n15542_), .B(new_n15541_), .Y(new_n15543_));
  XOR2   g14541(.A(new_n15543_), .B(new_n15538_), .Y(new_n15544_));
  NAND4  g14542(.A(new_n14876_), .B(new_n14869_), .C(new_n14847_), .D(new_n14834_), .Y(new_n15545_));
  OAI21  g14543(.A0(new_n14861_), .A1(new_n14850_), .B0(new_n15537_), .Y(new_n15546_));
  NAND2  g14544(.A(new_n14867_), .B(new_n14864_), .Y(new_n15547_));
  NAND2  g14545(.A(new_n15547_), .B(new_n15546_), .Y(new_n15548_));
  NAND4  g14546(.A(new_n14216_), .B(new_n14842_), .C(new_n14195_), .D(new_n14839_), .Y(new_n15549_));
  OAI21  g14547(.A0(new_n14843_), .A1(new_n14836_), .B0(new_n15549_), .Y(new_n15550_));
  AOI22  g14548(.A0(new_n15540_), .A1(new_n15550_), .B0(new_n14832_), .B1(new_n14829_), .Y(new_n15551_));
  NAND2  g14549(.A(new_n15551_), .B(new_n15548_), .Y(new_n15552_));
  NAND2  g14550(.A(new_n15543_), .B(new_n15538_), .Y(new_n15553_));
  NAND3  g14551(.A(new_n15553_), .B(new_n15552_), .C(new_n15545_), .Y(new_n15554_));
  OAI22  g14552(.A0(new_n15554_), .A1(new_n15529_), .B0(new_n15544_), .B1(new_n15535_), .Y(new_n15555_));
  XOR2   g14553(.A(new_n15555_), .B(new_n15522_), .Y(new_n15556_));
  XOR2   g14554(.A(new_n15556_), .B(new_n15489_), .Y(new_n15557_));
  XOR2   g14555(.A(new_n15557_), .B(new_n15486_), .Y(new_n15558_));
  XOR2   g14556(.A(new_n15558_), .B(new_n15416_), .Y(new_n15559_));
  NOR2   g14557(.A(new_n15559_), .B(new_n15391_), .Y(new_n15560_));
  OAI21  g14558(.A0(new_n15390_), .A1(new_n15380_), .B0(new_n15559_), .Y(new_n15561_));
  OAI22  g14559(.A0(new_n15561_), .A1(new_n15376_), .B0(new_n15560_), .B1(new_n15109_), .Y(new_n15562_));
  NAND2  g14560(.A(new_n15374_), .B(new_n15279_), .Y(new_n15563_));
  NOR2   g14561(.A(new_n15374_), .B(new_n15279_), .Y(new_n15564_));
  AOI21  g14562(.A0(new_n15563_), .A1(new_n15112_), .B0(new_n15564_), .Y(new_n15565_));
  NOR2   g14563(.A(new_n14437_), .B(new_n15285_), .Y(new_n15566_));
  OAI22  g14564(.A0(new_n15286_), .A1(new_n14362_), .B0(new_n15566_), .B1(new_n14243_), .Y(new_n15567_));
  NAND2  g14565(.A(new_n15339_), .B(new_n15328_), .Y(new_n15568_));
  NOR2   g14566(.A(new_n15371_), .B(new_n15370_), .Y(new_n15569_));
  OAI21  g14567(.A0(new_n15326_), .A1(new_n15569_), .B0(new_n15369_), .Y(new_n15570_));
  AOI21  g14568(.A0(new_n15334_), .A1(new_n15327_), .B0(new_n15369_), .Y(new_n15571_));
  AOI22  g14569(.A0(new_n15571_), .A1(new_n15568_), .B0(new_n15570_), .B1(new_n15567_), .Y(new_n15572_));
  OAI21  g14570(.A0(new_n15347_), .A1(new_n14373_), .B0(new_n15362_), .Y(new_n15573_));
  AOI22  g14571(.A0(new_n14419_), .A1(new_n14416_), .B0(new_n14386_), .B1(new_n14383_), .Y(new_n15574_));
  OAI221 g14572(.A0(new_n15358_), .A1(new_n14380_), .C0(new_n15574_), .B0(new_n15363_), .B1(new_n14413_), .Y(new_n15575_));
  NAND2  g14573(.A(new_n15575_), .B(new_n15573_), .Y(new_n15576_));
  NAND2  g14574(.A(new_n15360_), .B(new_n15365_), .Y(new_n15577_));
  NAND2  g14575(.A(new_n15577_), .B(new_n15576_), .Y(new_n15578_));
  NAND2  g14576(.A(new_n15320_), .B(new_n15323_), .Y(new_n15579_));
  AOI211 g14577(.A0(new_n15330_), .A1(new_n15329_), .B(new_n15323_), .C(new_n15332_), .Y(new_n15580_));
  AOI21  g14578(.A0(new_n15579_), .A1(new_n15327_), .B0(new_n15580_), .Y(new_n15581_));
  NAND2  g14579(.A(new_n15314_), .B(new_n15307_), .Y(new_n15582_));
  AOI221 g14580(.A0(new_n15305_), .A1(new_n15300_), .C0(new_n15582_), .B0(new_n15308_), .B1(new_n14326_), .Y(new_n15583_));
  OAI22  g14581(.A0(new_n15583_), .A1(new_n15303_), .B0(new_n15316_), .B1(new_n15306_), .Y(new_n15584_));
  NOR2   g14582(.A(new_n15333_), .B(new_n15295_), .Y(new_n15585_));
  OAI221 g14583(.A0(new_n15319_), .A1(new_n15297_), .C0(new_n15295_), .B0(new_n15311_), .B1(new_n15303_), .Y(new_n15586_));
  OAI211 g14584(.A0(new_n15585_), .A1(new_n15370_), .B0(new_n15584_), .B1(new_n15586_), .Y(new_n15587_));
  OAI21  g14585(.A0(new_n15584_), .A1(new_n15581_), .B0(new_n15587_), .Y(new_n15588_));
  OAI21  g14586(.A0(new_n15585_), .A1(new_n15370_), .B0(new_n15586_), .Y(new_n15589_));
  NAND4  g14587(.A(new_n15309_), .B(new_n15314_), .C(new_n15313_), .D(new_n15307_), .Y(new_n15590_));
  AOI22  g14588(.A0(new_n15590_), .A1(new_n15329_), .B0(new_n15310_), .B1(new_n15315_), .Y(new_n15591_));
  AOI211 g14589(.A0(new_n15579_), .A1(new_n15327_), .B(new_n15591_), .C(new_n15580_), .Y(new_n15592_));
  AOI211 g14590(.A0(new_n15591_), .A1(new_n15589_), .B(new_n15592_), .C(new_n15578_), .Y(new_n15593_));
  AOI21  g14591(.A0(new_n15588_), .A1(new_n15578_), .B0(new_n15593_), .Y(new_n15594_));
  XOR2   g14592(.A(new_n15594_), .B(new_n15572_), .Y(new_n15595_));
  NOR2   g14593(.A(new_n15277_), .B(new_n15205_), .Y(new_n15596_));
  NAND2  g14594(.A(new_n15277_), .B(new_n15205_), .Y(new_n15597_));
  OAI21  g14595(.A0(new_n15596_), .A1(new_n15130_), .B0(new_n15597_), .Y(new_n15598_));
  NAND2  g14596(.A(new_n15275_), .B(new_n15242_), .Y(new_n15599_));
  NAND2  g14597(.A(new_n15599_), .B(new_n15208_), .Y(new_n15600_));
  XOR2   g14598(.A(new_n14524_), .B(new_n15247_), .Y(new_n15601_));
  XOR2   g14599(.A(new_n14611_), .B(new_n15214_), .Y(new_n15602_));
  NAND2  g14600(.A(new_n15602_), .B(new_n15601_), .Y(new_n15603_));
  NOR2   g14601(.A(new_n15602_), .B(new_n15601_), .Y(new_n15604_));
  AOI21  g14602(.A0(new_n15603_), .A1(new_n14453_), .B0(new_n15604_), .Y(new_n15605_));
  OAI21  g14603(.A0(new_n15215_), .A1(new_n15214_), .B0(new_n15232_), .Y(new_n15606_));
  XOR2   g14604(.A(new_n15230_), .B(new_n15235_), .Y(new_n15607_));
  OAI21  g14605(.A0(new_n15230_), .A1(new_n15225_), .B0(new_n15232_), .Y(new_n15608_));
  AOI221 g14606(.A0(new_n15230_), .A1(new_n15225_), .C0(new_n15608_), .B0(new_n15217_), .B1(new_n14536_), .Y(new_n15609_));
  AOI21  g14607(.A0(new_n15607_), .A1(new_n15606_), .B0(new_n15609_), .Y(new_n15610_));
  OAI21  g14608(.A0(new_n15248_), .A1(new_n15247_), .B0(new_n15265_), .Y(new_n15611_));
  XOR2   g14609(.A(new_n15263_), .B(new_n15268_), .Y(new_n15612_));
  OAI21  g14610(.A0(new_n15263_), .A1(new_n15258_), .B0(new_n15265_), .Y(new_n15613_));
  AOI221 g14611(.A0(new_n15263_), .A1(new_n15258_), .C0(new_n15613_), .B0(new_n15250_), .B1(new_n14456_), .Y(new_n15614_));
  AOI21  g14612(.A0(new_n15612_), .A1(new_n15611_), .B0(new_n15614_), .Y(new_n15615_));
  NOR2   g14613(.A(new_n15615_), .B(new_n15610_), .Y(new_n15616_));
  AOI211 g14614(.A0(new_n15607_), .A1(new_n15606_), .B(new_n15614_), .C(new_n15609_), .Y(new_n15617_));
  OAI21  g14615(.A0(new_n15264_), .A1(new_n15255_), .B0(new_n15617_), .Y(new_n15618_));
  OAI21  g14616(.A0(new_n15616_), .A1(new_n15605_), .B0(new_n15618_), .Y(new_n15619_));
  NAND4  g14617(.A(new_n15229_), .B(new_n15228_), .C(new_n15234_), .D(new_n15233_), .Y(new_n15620_));
  INV    g14618(.A(new_n15620_), .Y(new_n15621_));
  OAI22  g14619(.A0(new_n15621_), .A1(new_n15222_), .B0(new_n15238_), .B1(new_n15225_), .Y(new_n15622_));
  NAND4  g14620(.A(new_n15262_), .B(new_n15261_), .C(new_n15267_), .D(new_n15266_), .Y(new_n15623_));
  INV    g14621(.A(new_n15623_), .Y(new_n15624_));
  OAI22  g14622(.A0(new_n15624_), .A1(new_n15255_), .B0(new_n15271_), .B1(new_n15258_), .Y(new_n15625_));
  XOR2   g14623(.A(new_n15625_), .B(new_n15622_), .Y(new_n15626_));
  OAI22  g14624(.A0(new_n15274_), .A1(new_n15249_), .B0(new_n15241_), .B1(new_n15216_), .Y(new_n15627_));
  AOI221 g14625(.A0(new_n15612_), .A1(new_n15611_), .C0(new_n15627_), .B0(new_n15607_), .B1(new_n15606_), .Y(new_n15628_));
  AOI22  g14626(.A0(new_n15620_), .A1(new_n15606_), .B0(new_n15230_), .B1(new_n15235_), .Y(new_n15629_));
  NOR2   g14627(.A(new_n15625_), .B(new_n15629_), .Y(new_n15630_));
  AOI22  g14628(.A0(new_n15623_), .A1(new_n15611_), .B0(new_n15263_), .B1(new_n15268_), .Y(new_n15631_));
  NOR2   g14629(.A(new_n15631_), .B(new_n15622_), .Y(new_n15632_));
  NOR3   g14630(.A(new_n15632_), .B(new_n15630_), .C(new_n15628_), .Y(new_n15633_));
  AOI22  g14631(.A0(new_n15633_), .A1(new_n15600_), .B0(new_n15626_), .B1(new_n15619_), .Y(new_n15634_));
  NAND2  g14632(.A(new_n15203_), .B(new_n15167_), .Y(new_n15635_));
  NAND2  g14633(.A(new_n15635_), .B(new_n15133_), .Y(new_n15636_));
  XOR2   g14634(.A(new_n14704_), .B(new_n15175_), .Y(new_n15637_));
  XOR2   g14635(.A(new_n14783_), .B(new_n15139_), .Y(new_n15638_));
  NAND2  g14636(.A(new_n15638_), .B(new_n15637_), .Y(new_n15639_));
  NOR2   g14637(.A(new_n15638_), .B(new_n15637_), .Y(new_n15640_));
  AOI21  g14638(.A0(new_n15639_), .A1(new_n15384_), .B0(new_n15640_), .Y(new_n15641_));
  OAI21  g14639(.A0(new_n15140_), .A1(new_n15139_), .B0(new_n15157_), .Y(new_n15642_));
  XOR2   g14640(.A(new_n15155_), .B(new_n15160_), .Y(new_n15643_));
  OAI21  g14641(.A0(new_n15155_), .A1(new_n15150_), .B0(new_n15157_), .Y(new_n15644_));
  AOI221 g14642(.A0(new_n15155_), .A1(new_n15150_), .C0(new_n15644_), .B0(new_n15142_), .B1(new_n14708_), .Y(new_n15645_));
  AOI21  g14643(.A0(new_n15643_), .A1(new_n15642_), .B0(new_n15645_), .Y(new_n15646_));
  OAI21  g14644(.A0(new_n15176_), .A1(new_n15175_), .B0(new_n15193_), .Y(new_n15647_));
  XOR2   g14645(.A(new_n15191_), .B(new_n15196_), .Y(new_n15648_));
  OAI21  g14646(.A0(new_n15191_), .A1(new_n15186_), .B0(new_n15193_), .Y(new_n15649_));
  AOI221 g14647(.A0(new_n15191_), .A1(new_n15186_), .C0(new_n15649_), .B0(new_n15178_), .B1(new_n14629_), .Y(new_n15650_));
  AOI21  g14648(.A0(new_n15648_), .A1(new_n15647_), .B0(new_n15650_), .Y(new_n15651_));
  NOR2   g14649(.A(new_n15651_), .B(new_n15646_), .Y(new_n15652_));
  AOI211 g14650(.A0(new_n15643_), .A1(new_n15642_), .B(new_n15650_), .C(new_n15645_), .Y(new_n15653_));
  OAI21  g14651(.A0(new_n15192_), .A1(new_n15183_), .B0(new_n15653_), .Y(new_n15654_));
  OAI21  g14652(.A0(new_n15652_), .A1(new_n15641_), .B0(new_n15654_), .Y(new_n15655_));
  NAND4  g14653(.A(new_n15154_), .B(new_n15153_), .C(new_n15159_), .D(new_n15158_), .Y(new_n15656_));
  INV    g14654(.A(new_n15656_), .Y(new_n15657_));
  OAI22  g14655(.A0(new_n15657_), .A1(new_n15147_), .B0(new_n15163_), .B1(new_n15150_), .Y(new_n15658_));
  NAND4  g14656(.A(new_n15190_), .B(new_n15189_), .C(new_n15195_), .D(new_n15194_), .Y(new_n15659_));
  INV    g14657(.A(new_n15659_), .Y(new_n15660_));
  OAI22  g14658(.A0(new_n15660_), .A1(new_n15183_), .B0(new_n15199_), .B1(new_n15186_), .Y(new_n15661_));
  XOR2   g14659(.A(new_n15661_), .B(new_n15658_), .Y(new_n15662_));
  OAI22  g14660(.A0(new_n15202_), .A1(new_n15177_), .B0(new_n15166_), .B1(new_n15141_), .Y(new_n15663_));
  AOI221 g14661(.A0(new_n15648_), .A1(new_n15647_), .C0(new_n15663_), .B0(new_n15643_), .B1(new_n15642_), .Y(new_n15664_));
  AOI22  g14662(.A0(new_n15656_), .A1(new_n15642_), .B0(new_n15155_), .B1(new_n15160_), .Y(new_n15665_));
  NOR2   g14663(.A(new_n15661_), .B(new_n15665_), .Y(new_n15666_));
  AOI22  g14664(.A0(new_n15659_), .A1(new_n15647_), .B0(new_n15191_), .B1(new_n15196_), .Y(new_n15667_));
  NOR2   g14665(.A(new_n15667_), .B(new_n15658_), .Y(new_n15668_));
  NOR3   g14666(.A(new_n15668_), .B(new_n15666_), .C(new_n15664_), .Y(new_n15669_));
  AOI22  g14667(.A0(new_n15669_), .A1(new_n15636_), .B0(new_n15662_), .B1(new_n15655_), .Y(new_n15670_));
  XOR2   g14668(.A(new_n15670_), .B(new_n15634_), .Y(new_n15671_));
  XOR2   g14669(.A(new_n15671_), .B(new_n15598_), .Y(new_n15672_));
  XOR2   g14670(.A(new_n15672_), .B(new_n15595_), .Y(new_n15673_));
  NAND2  g14671(.A(new_n15673_), .B(new_n15565_), .Y(new_n15674_));
  XOR2   g14672(.A(new_n15373_), .B(new_n15567_), .Y(new_n15675_));
  NOR2   g14673(.A(new_n15675_), .B(new_n15389_), .Y(new_n15676_));
  NAND2  g14674(.A(new_n15675_), .B(new_n15389_), .Y(new_n15677_));
  OAI21  g14675(.A0(new_n15676_), .A1(new_n15380_), .B0(new_n15677_), .Y(new_n15678_));
  XOR2   g14676(.A(new_n15673_), .B(new_n15678_), .Y(new_n15679_));
  XOR2   g14677(.A(new_n15023_), .B(new_n15457_), .Y(new_n15680_));
  XOR2   g14678(.A(new_n15095_), .B(new_n15425_), .Y(new_n15681_));
  NAND2  g14679(.A(new_n15681_), .B(new_n15680_), .Y(new_n15682_));
  NOR2   g14680(.A(new_n15681_), .B(new_n15680_), .Y(new_n15683_));
  AOI21  g14681(.A0(new_n15682_), .A1(new_n15412_), .B0(new_n15683_), .Y(new_n15684_));
  XOR2   g14682(.A(new_n15485_), .B(new_n15684_), .Y(new_n15685_));
  XOR2   g14683(.A(new_n14878_), .B(new_n15527_), .Y(new_n15686_));
  XOR2   g14684(.A(new_n14941_), .B(new_n15494_), .Y(new_n15687_));
  NAND2  g14685(.A(new_n15687_), .B(new_n15686_), .Y(new_n15688_));
  NOR2   g14686(.A(new_n15687_), .B(new_n15686_), .Y(new_n15689_));
  AOI21  g14687(.A0(new_n15688_), .A1(new_n15404_), .B0(new_n15689_), .Y(new_n15690_));
  XOR2   g14688(.A(new_n15556_), .B(new_n15690_), .Y(new_n15691_));
  NAND2  g14689(.A(new_n15691_), .B(new_n15685_), .Y(new_n15692_));
  NOR2   g14690(.A(new_n15691_), .B(new_n15685_), .Y(new_n15693_));
  AOI21  g14691(.A0(new_n15692_), .A1(new_n15416_), .B0(new_n15693_), .Y(new_n15694_));
  NAND2  g14692(.A(new_n15555_), .B(new_n15522_), .Y(new_n15695_));
  NAND2  g14693(.A(new_n15695_), .B(new_n15489_), .Y(new_n15696_));
  OAI21  g14694(.A0(new_n15495_), .A1(new_n15494_), .B0(new_n15512_), .Y(new_n15697_));
  XOR2   g14695(.A(new_n15510_), .B(new_n15515_), .Y(new_n15698_));
  OAI21  g14696(.A0(new_n15510_), .A1(new_n15505_), .B0(new_n15512_), .Y(new_n15699_));
  AOI221 g14697(.A0(new_n15510_), .A1(new_n15505_), .C0(new_n15699_), .B0(new_n15497_), .B1(new_n14882_), .Y(new_n15700_));
  AOI21  g14698(.A0(new_n15698_), .A1(new_n15697_), .B0(new_n15700_), .Y(new_n15701_));
  OAI21  g14699(.A0(new_n15528_), .A1(new_n15527_), .B0(new_n15545_), .Y(new_n15702_));
  XOR2   g14700(.A(new_n15543_), .B(new_n15548_), .Y(new_n15703_));
  OAI21  g14701(.A0(new_n15543_), .A1(new_n15538_), .B0(new_n15545_), .Y(new_n15704_));
  AOI221 g14702(.A0(new_n15543_), .A1(new_n15538_), .C0(new_n15704_), .B0(new_n15530_), .B1(new_n14818_), .Y(new_n15705_));
  AOI21  g14703(.A0(new_n15703_), .A1(new_n15702_), .B0(new_n15705_), .Y(new_n15706_));
  NOR2   g14704(.A(new_n15706_), .B(new_n15701_), .Y(new_n15707_));
  AOI211 g14705(.A0(new_n15698_), .A1(new_n15697_), .B(new_n15705_), .C(new_n15700_), .Y(new_n15708_));
  OAI21  g14706(.A0(new_n15544_), .A1(new_n15535_), .B0(new_n15708_), .Y(new_n15709_));
  OAI21  g14707(.A0(new_n15707_), .A1(new_n15690_), .B0(new_n15709_), .Y(new_n15710_));
  NAND4  g14708(.A(new_n15509_), .B(new_n15508_), .C(new_n15514_), .D(new_n15513_), .Y(new_n15711_));
  INV    g14709(.A(new_n15711_), .Y(new_n15712_));
  OAI22  g14710(.A0(new_n15712_), .A1(new_n15502_), .B0(new_n15518_), .B1(new_n15505_), .Y(new_n15713_));
  NAND4  g14711(.A(new_n15542_), .B(new_n15541_), .C(new_n15547_), .D(new_n15546_), .Y(new_n15714_));
  INV    g14712(.A(new_n15714_), .Y(new_n15715_));
  OAI22  g14713(.A0(new_n15715_), .A1(new_n15535_), .B0(new_n15551_), .B1(new_n15538_), .Y(new_n15716_));
  XOR2   g14714(.A(new_n15716_), .B(new_n15713_), .Y(new_n15717_));
  OAI22  g14715(.A0(new_n15554_), .A1(new_n15529_), .B0(new_n15521_), .B1(new_n15496_), .Y(new_n15718_));
  AOI221 g14716(.A0(new_n15703_), .A1(new_n15702_), .C0(new_n15718_), .B0(new_n15698_), .B1(new_n15697_), .Y(new_n15719_));
  AOI22  g14717(.A0(new_n15711_), .A1(new_n15697_), .B0(new_n15510_), .B1(new_n15515_), .Y(new_n15720_));
  NOR2   g14718(.A(new_n15716_), .B(new_n15720_), .Y(new_n15721_));
  AOI22  g14719(.A0(new_n15714_), .A1(new_n15702_), .B0(new_n15543_), .B1(new_n15548_), .Y(new_n15722_));
  NOR2   g14720(.A(new_n15722_), .B(new_n15713_), .Y(new_n15723_));
  NOR3   g14721(.A(new_n15723_), .B(new_n15721_), .C(new_n15719_), .Y(new_n15724_));
  AOI22  g14722(.A0(new_n15724_), .A1(new_n15696_), .B0(new_n15717_), .B1(new_n15710_), .Y(new_n15725_));
  NAND2  g14723(.A(new_n15484_), .B(new_n15452_), .Y(new_n15726_));
  NAND2  g14724(.A(new_n15726_), .B(new_n15419_), .Y(new_n15727_));
  OAI21  g14725(.A0(new_n15426_), .A1(new_n15425_), .B0(new_n15442_), .Y(new_n15728_));
  XOR2   g14726(.A(new_n15440_), .B(new_n15445_), .Y(new_n15729_));
  OAI21  g14727(.A0(new_n15440_), .A1(new_n15435_), .B0(new_n15442_), .Y(new_n15730_));
  AOI221 g14728(.A0(new_n15440_), .A1(new_n15435_), .C0(new_n15730_), .B0(new_n15428_), .B1(new_n15027_), .Y(new_n15731_));
  AOI21  g14729(.A0(new_n15729_), .A1(new_n15728_), .B0(new_n15731_), .Y(new_n15732_));
  OAI21  g14730(.A0(new_n15458_), .A1(new_n15457_), .B0(new_n15474_), .Y(new_n15733_));
  XOR2   g14731(.A(new_n15472_), .B(new_n15477_), .Y(new_n15734_));
  OAI21  g14732(.A0(new_n15472_), .A1(new_n15467_), .B0(new_n15474_), .Y(new_n15735_));
  AOI221 g14733(.A0(new_n15472_), .A1(new_n15467_), .C0(new_n15735_), .B0(new_n15460_), .B1(new_n14961_), .Y(new_n15736_));
  AOI21  g14734(.A0(new_n15734_), .A1(new_n15733_), .B0(new_n15736_), .Y(new_n15737_));
  NOR2   g14735(.A(new_n15737_), .B(new_n15732_), .Y(new_n15738_));
  AOI211 g14736(.A0(new_n15729_), .A1(new_n15728_), .B(new_n15736_), .C(new_n15731_), .Y(new_n15739_));
  OAI21  g14737(.A0(new_n15473_), .A1(new_n15464_), .B0(new_n15739_), .Y(new_n15740_));
  OAI21  g14738(.A0(new_n15738_), .A1(new_n15684_), .B0(new_n15740_), .Y(new_n15741_));
  NAND4  g14739(.A(new_n15439_), .B(new_n15438_), .C(new_n15444_), .D(new_n15443_), .Y(new_n15742_));
  INV    g14740(.A(new_n15742_), .Y(new_n15743_));
  OAI22  g14741(.A0(new_n15743_), .A1(new_n15432_), .B0(new_n15448_), .B1(new_n15435_), .Y(new_n15744_));
  NAND4  g14742(.A(new_n15471_), .B(new_n15470_), .C(new_n15476_), .D(new_n15475_), .Y(new_n15745_));
  INV    g14743(.A(new_n15745_), .Y(new_n15746_));
  OAI22  g14744(.A0(new_n15746_), .A1(new_n15464_), .B0(new_n15480_), .B1(new_n15467_), .Y(new_n15747_));
  XOR2   g14745(.A(new_n15747_), .B(new_n15744_), .Y(new_n15748_));
  OAI22  g14746(.A0(new_n15483_), .A1(new_n15459_), .B0(new_n15451_), .B1(new_n15427_), .Y(new_n15749_));
  AOI221 g14747(.A0(new_n15734_), .A1(new_n15733_), .C0(new_n15749_), .B0(new_n15729_), .B1(new_n15728_), .Y(new_n15750_));
  AOI22  g14748(.A0(new_n15742_), .A1(new_n15728_), .B0(new_n15440_), .B1(new_n15445_), .Y(new_n15751_));
  NOR2   g14749(.A(new_n15747_), .B(new_n15751_), .Y(new_n15752_));
  AOI22  g14750(.A0(new_n15745_), .A1(new_n15733_), .B0(new_n15472_), .B1(new_n15477_), .Y(new_n15753_));
  NOR2   g14751(.A(new_n15753_), .B(new_n15744_), .Y(new_n15754_));
  NOR3   g14752(.A(new_n15754_), .B(new_n15752_), .C(new_n15750_), .Y(new_n15755_));
  AOI22  g14753(.A0(new_n15755_), .A1(new_n15727_), .B0(new_n15748_), .B1(new_n15741_), .Y(new_n15756_));
  XOR2   g14754(.A(new_n15756_), .B(new_n15725_), .Y(new_n15757_));
  XOR2   g14755(.A(new_n15757_), .B(new_n15694_), .Y(new_n15758_));
  NAND2  g14756(.A(new_n15758_), .B(new_n15679_), .Y(new_n15759_));
  XOR2   g14757(.A(new_n15204_), .B(new_n15641_), .Y(new_n15760_));
  XOR2   g14758(.A(new_n15276_), .B(new_n15605_), .Y(new_n15761_));
  NAND2  g14759(.A(new_n15761_), .B(new_n15760_), .Y(new_n15762_));
  NOR2   g14760(.A(new_n15761_), .B(new_n15760_), .Y(new_n15763_));
  AOI21  g14761(.A0(new_n15762_), .A1(new_n15388_), .B0(new_n15763_), .Y(new_n15764_));
  XOR2   g14762(.A(new_n15671_), .B(new_n15764_), .Y(new_n15765_));
  XOR2   g14763(.A(new_n15765_), .B(new_n15595_), .Y(new_n15766_));
  AOI21  g14764(.A0(new_n15766_), .A1(new_n15678_), .B0(new_n15758_), .Y(new_n15767_));
  AOI22  g14765(.A0(new_n15767_), .A1(new_n15674_), .B0(new_n15759_), .B1(new_n15562_), .Y(new_n15768_));
  NOR2   g14766(.A(new_n15361_), .B(new_n15352_), .Y(new_n15769_));
  NOR2   g14767(.A(new_n15368_), .B(new_n15348_), .Y(new_n15770_));
  NOR2   g14768(.A(new_n15770_), .B(new_n15769_), .Y(new_n15771_));
  NOR2   g14769(.A(new_n15771_), .B(new_n15340_), .Y(new_n15772_));
  NAND2  g14770(.A(new_n15571_), .B(new_n15568_), .Y(new_n15773_));
  OAI21  g14771(.A0(new_n15772_), .A1(new_n15288_), .B0(new_n15773_), .Y(new_n15774_));
  XOR2   g14772(.A(new_n15594_), .B(new_n15774_), .Y(new_n15775_));
  NOR2   g14773(.A(new_n15672_), .B(new_n15775_), .Y(new_n15776_));
  NAND2  g14774(.A(new_n15672_), .B(new_n15775_), .Y(new_n15777_));
  OAI21  g14775(.A0(new_n15776_), .A1(new_n15565_), .B0(new_n15777_), .Y(new_n15778_));
  NAND2  g14776(.A(new_n15588_), .B(new_n15578_), .Y(new_n15779_));
  OAI21  g14777(.A0(new_n15593_), .A1(new_n15572_), .B0(new_n15779_), .Y(new_n15780_));
  NOR2   g14778(.A(new_n15591_), .B(new_n15581_), .Y(new_n15781_));
  AOI22  g14779(.A0(new_n15575_), .A1(new_n15573_), .B0(new_n15360_), .B1(new_n15365_), .Y(new_n15782_));
  AOI21  g14780(.A0(new_n15591_), .A1(new_n15589_), .B0(new_n15592_), .Y(new_n15783_));
  NOR2   g14781(.A(new_n15783_), .B(new_n15782_), .Y(new_n15784_));
  OAI211 g14782(.A0(new_n15584_), .A1(new_n15581_), .B0(new_n15587_), .B1(new_n15782_), .Y(new_n15785_));
  AOI211 g14783(.A0(new_n15785_), .A1(new_n15774_), .B(new_n15781_), .C(new_n15784_), .Y(new_n15786_));
  AOI21  g14784(.A0(new_n15781_), .A1(new_n15780_), .B0(new_n15786_), .Y(new_n15787_));
  AOI21  g14785(.A0(new_n15599_), .A1(new_n15208_), .B0(new_n15628_), .Y(new_n15788_));
  XOR2   g14786(.A(new_n15625_), .B(new_n15629_), .Y(new_n15789_));
  NOR2   g14787(.A(new_n15789_), .B(new_n15788_), .Y(new_n15790_));
  NOR2   g14788(.A(new_n15616_), .B(new_n15605_), .Y(new_n15791_));
  NOR4   g14789(.A(new_n15632_), .B(new_n15630_), .C(new_n15628_), .D(new_n15791_), .Y(new_n15792_));
  AOI21  g14790(.A0(new_n15635_), .A1(new_n15133_), .B0(new_n15664_), .Y(new_n15793_));
  XOR2   g14791(.A(new_n15661_), .B(new_n15665_), .Y(new_n15794_));
  NOR2   g14792(.A(new_n15794_), .B(new_n15793_), .Y(new_n15795_));
  NOR2   g14793(.A(new_n15652_), .B(new_n15641_), .Y(new_n15796_));
  NOR4   g14794(.A(new_n15668_), .B(new_n15666_), .C(new_n15664_), .D(new_n15796_), .Y(new_n15797_));
  OAI22  g14795(.A0(new_n15797_), .A1(new_n15795_), .B0(new_n15792_), .B1(new_n15790_), .Y(new_n15798_));
  NOR4   g14796(.A(new_n15797_), .B(new_n15795_), .C(new_n15792_), .D(new_n15790_), .Y(new_n15799_));
  AOI21  g14797(.A0(new_n15798_), .A1(new_n15598_), .B0(new_n15799_), .Y(new_n15800_));
  AOI22  g14798(.A0(new_n15191_), .A1(new_n15196_), .B0(new_n15155_), .B1(new_n15160_), .Y(new_n15801_));
  OAI221 g14799(.A0(new_n15660_), .A1(new_n15183_), .C0(new_n15801_), .B0(new_n15657_), .B1(new_n15147_), .Y(new_n15802_));
  INV    g14800(.A(new_n15802_), .Y(new_n15803_));
  OAI22  g14801(.A0(new_n15803_), .A1(new_n15793_), .B0(new_n15667_), .B1(new_n15665_), .Y(new_n15804_));
  AOI22  g14802(.A0(new_n15263_), .A1(new_n15268_), .B0(new_n15230_), .B1(new_n15235_), .Y(new_n15805_));
  OAI221 g14803(.A0(new_n15624_), .A1(new_n15255_), .C0(new_n15805_), .B0(new_n15621_), .B1(new_n15222_), .Y(new_n15806_));
  AOI22  g14804(.A0(new_n15806_), .A1(new_n15619_), .B0(new_n15625_), .B1(new_n15622_), .Y(new_n15807_));
  XOR2   g14805(.A(new_n15807_), .B(new_n15804_), .Y(new_n15808_));
  NOR2   g14806(.A(new_n15808_), .B(new_n15800_), .Y(new_n15809_));
  NAND2  g14807(.A(new_n15798_), .B(new_n15598_), .Y(new_n15810_));
  NOR2   g14808(.A(new_n15670_), .B(new_n15634_), .Y(new_n15811_));
  AOI22  g14809(.A0(new_n15669_), .A1(new_n15636_), .B0(new_n15633_), .B1(new_n15600_), .Y(new_n15812_));
  OAI221 g14810(.A0(new_n15794_), .A1(new_n15793_), .C0(new_n15812_), .B0(new_n15789_), .B1(new_n15788_), .Y(new_n15813_));
  OAI21  g14811(.A0(new_n15811_), .A1(new_n15764_), .B0(new_n15813_), .Y(new_n15814_));
  INV    g14812(.A(new_n15806_), .Y(new_n15815_));
  OAI22  g14813(.A0(new_n15815_), .A1(new_n15788_), .B0(new_n15631_), .B1(new_n15629_), .Y(new_n15816_));
  XOR2   g14814(.A(new_n15816_), .B(new_n15804_), .Y(new_n15817_));
  AOI22  g14815(.A0(new_n15802_), .A1(new_n15655_), .B0(new_n15661_), .B1(new_n15658_), .Y(new_n15818_));
  NOR2   g14816(.A(new_n15816_), .B(new_n15818_), .Y(new_n15819_));
  NOR2   g14817(.A(new_n15807_), .B(new_n15804_), .Y(new_n15820_));
  NOR3   g14818(.A(new_n15820_), .B(new_n15819_), .C(new_n15799_), .Y(new_n15821_));
  AOI22  g14819(.A0(new_n15821_), .A1(new_n15810_), .B0(new_n15817_), .B1(new_n15814_), .Y(new_n15822_));
  AOI21  g14820(.A0(new_n15785_), .A1(new_n15774_), .B0(new_n15784_), .Y(new_n15823_));
  NAND2  g14821(.A(new_n15584_), .B(new_n15589_), .Y(new_n15824_));
  OAI211 g14822(.A0(new_n15593_), .A1(new_n15572_), .B0(new_n15824_), .B1(new_n15779_), .Y(new_n15825_));
  NOR2   g14823(.A(new_n15811_), .B(new_n15764_), .Y(new_n15826_));
  NAND2  g14824(.A(new_n15807_), .B(new_n15804_), .Y(new_n15827_));
  NAND2  g14825(.A(new_n15816_), .B(new_n15818_), .Y(new_n15828_));
  NAND3  g14826(.A(new_n15828_), .B(new_n15827_), .C(new_n15813_), .Y(new_n15829_));
  OAI221 g14827(.A0(new_n15829_), .A1(new_n15826_), .C0(new_n15825_), .B0(new_n15824_), .B1(new_n15823_), .Y(new_n15830_));
  OAI22  g14828(.A0(new_n15830_), .A1(new_n15809_), .B0(new_n15822_), .B1(new_n15787_), .Y(new_n15831_));
  XOR2   g14829(.A(new_n15831_), .B(new_n15778_), .Y(new_n15832_));
  NOR2   g14830(.A(new_n15756_), .B(new_n15725_), .Y(new_n15833_));
  NAND2  g14831(.A(new_n15717_), .B(new_n15710_), .Y(new_n15834_));
  NAND2  g14832(.A(new_n15748_), .B(new_n15741_), .Y(new_n15835_));
  AOI22  g14833(.A0(new_n15755_), .A1(new_n15727_), .B0(new_n15724_), .B1(new_n15696_), .Y(new_n15836_));
  NAND3  g14834(.A(new_n15836_), .B(new_n15835_), .C(new_n15834_), .Y(new_n15837_));
  OAI21  g14835(.A0(new_n15833_), .A1(new_n15694_), .B0(new_n15837_), .Y(new_n15838_));
  AOI22  g14836(.A0(new_n15472_), .A1(new_n15477_), .B0(new_n15440_), .B1(new_n15445_), .Y(new_n15839_));
  OAI221 g14837(.A0(new_n15746_), .A1(new_n15464_), .C0(new_n15839_), .B0(new_n15743_), .B1(new_n15432_), .Y(new_n15840_));
  AOI22  g14838(.A0(new_n15840_), .A1(new_n15741_), .B0(new_n15747_), .B1(new_n15744_), .Y(new_n15841_));
  AOI22  g14839(.A0(new_n15543_), .A1(new_n15548_), .B0(new_n15510_), .B1(new_n15515_), .Y(new_n15842_));
  OAI221 g14840(.A0(new_n15715_), .A1(new_n15535_), .C0(new_n15842_), .B0(new_n15712_), .B1(new_n15502_), .Y(new_n15843_));
  AOI22  g14841(.A0(new_n15843_), .A1(new_n15710_), .B0(new_n15716_), .B1(new_n15713_), .Y(new_n15844_));
  XOR2   g14842(.A(new_n15844_), .B(new_n15841_), .Y(new_n15845_));
  NAND2  g14843(.A(new_n15845_), .B(new_n15838_), .Y(new_n15846_));
  XOR2   g14844(.A(new_n14222_), .B(new_n15397_), .Y(new_n15847_));
  NOR2   g14845(.A(new_n15847_), .B(new_n13953_), .Y(new_n15848_));
  NAND2  g14846(.A(new_n15847_), .B(new_n13953_), .Y(new_n15849_));
  OAI21  g14847(.A0(new_n15848_), .A1(new_n13716_), .B0(new_n15849_), .Y(new_n15850_));
  NAND2  g14848(.A(new_n15098_), .B(new_n14944_), .Y(new_n15851_));
  NOR2   g14849(.A(new_n15098_), .B(new_n14944_), .Y(new_n15852_));
  AOI21  g14850(.A0(new_n15851_), .A1(new_n15850_), .B0(new_n15852_), .Y(new_n15853_));
  NOR2   g14851(.A(new_n15557_), .B(new_n15486_), .Y(new_n15854_));
  NAND2  g14852(.A(new_n15557_), .B(new_n15486_), .Y(new_n15855_));
  OAI21  g14853(.A0(new_n15854_), .A1(new_n15853_), .B0(new_n15855_), .Y(new_n15856_));
  OAI21  g14854(.A0(new_n15756_), .A1(new_n15725_), .B0(new_n15856_), .Y(new_n15857_));
  NOR2   g14855(.A(new_n15707_), .B(new_n15690_), .Y(new_n15858_));
  NAND2  g14856(.A(new_n15722_), .B(new_n15713_), .Y(new_n15859_));
  NAND2  g14857(.A(new_n15716_), .B(new_n15720_), .Y(new_n15860_));
  NAND3  g14858(.A(new_n15860_), .B(new_n15859_), .C(new_n15709_), .Y(new_n15861_));
  NOR2   g14859(.A(new_n15738_), .B(new_n15684_), .Y(new_n15862_));
  NAND2  g14860(.A(new_n15753_), .B(new_n15744_), .Y(new_n15863_));
  NAND2  g14861(.A(new_n15747_), .B(new_n15751_), .Y(new_n15864_));
  NAND3  g14862(.A(new_n15864_), .B(new_n15863_), .C(new_n15740_), .Y(new_n15865_));
  OAI22  g14863(.A0(new_n15865_), .A1(new_n15862_), .B0(new_n15861_), .B1(new_n15858_), .Y(new_n15866_));
  AOI221 g14864(.A0(new_n15748_), .A1(new_n15741_), .C0(new_n15866_), .B0(new_n15717_), .B1(new_n15710_), .Y(new_n15867_));
  AOI21  g14865(.A0(new_n15695_), .A1(new_n15489_), .B0(new_n15719_), .Y(new_n15868_));
  INV    g14866(.A(new_n15843_), .Y(new_n15869_));
  OAI22  g14867(.A0(new_n15869_), .A1(new_n15868_), .B0(new_n15722_), .B1(new_n15720_), .Y(new_n15870_));
  NOR2   g14868(.A(new_n15870_), .B(new_n15841_), .Y(new_n15871_));
  AOI21  g14869(.A0(new_n15726_), .A1(new_n15419_), .B0(new_n15750_), .Y(new_n15872_));
  INV    g14870(.A(new_n15840_), .Y(new_n15873_));
  OAI22  g14871(.A0(new_n15873_), .A1(new_n15872_), .B0(new_n15753_), .B1(new_n15751_), .Y(new_n15874_));
  NOR2   g14872(.A(new_n15844_), .B(new_n15874_), .Y(new_n15875_));
  NOR3   g14873(.A(new_n15875_), .B(new_n15871_), .C(new_n15867_), .Y(new_n15876_));
  NAND2  g14874(.A(new_n15876_), .B(new_n15857_), .Y(new_n15877_));
  NAND2  g14875(.A(new_n15877_), .B(new_n15846_), .Y(new_n15878_));
  AOI21  g14876(.A0(new_n15878_), .A1(new_n15832_), .B0(new_n15768_), .Y(new_n15879_));
  NAND2  g14877(.A(new_n15765_), .B(new_n15595_), .Y(new_n15880_));
  NOR2   g14878(.A(new_n15765_), .B(new_n15595_), .Y(new_n15881_));
  AOI21  g14879(.A0(new_n15880_), .A1(new_n15678_), .B0(new_n15881_), .Y(new_n15882_));
  AOI22  g14880(.A0(new_n15876_), .A1(new_n15857_), .B0(new_n15845_), .B1(new_n15838_), .Y(new_n15883_));
  OAI21  g14881(.A0(new_n15831_), .A1(new_n15882_), .B0(new_n15883_), .Y(new_n15884_));
  AOI21  g14882(.A0(new_n15831_), .A1(new_n15882_), .B0(new_n15884_), .Y(new_n15885_));
  NAND2  g14883(.A(new_n15817_), .B(new_n15814_), .Y(new_n15886_));
  AOI221 g14884(.A0(new_n15821_), .A1(new_n15810_), .C0(new_n15786_), .B0(new_n15781_), .B1(new_n15780_), .Y(new_n15887_));
  NAND2  g14885(.A(new_n15887_), .B(new_n15886_), .Y(new_n15888_));
  OAI21  g14886(.A0(new_n15822_), .A1(new_n15787_), .B0(new_n15778_), .Y(new_n15889_));
  NAND2  g14887(.A(new_n15781_), .B(new_n15780_), .Y(new_n15890_));
  AOI22  g14888(.A0(new_n15661_), .A1(new_n15658_), .B0(new_n15625_), .B1(new_n15622_), .Y(new_n15891_));
  OAI221 g14889(.A0(new_n15815_), .A1(new_n15788_), .C0(new_n15891_), .B0(new_n15803_), .B1(new_n15793_), .Y(new_n15892_));
  NAND2  g14890(.A(new_n15892_), .B(new_n15814_), .Y(new_n15893_));
  OAI211 g14891(.A0(new_n15807_), .A1(new_n15818_), .B0(new_n15893_), .B1(new_n15890_), .Y(new_n15894_));
  NOR2   g14892(.A(new_n15807_), .B(new_n15818_), .Y(new_n15895_));
  AOI21  g14893(.A0(new_n15892_), .A1(new_n15814_), .B0(new_n15895_), .Y(new_n15896_));
  OAI21  g14894(.A0(new_n15896_), .A1(new_n15890_), .B0(new_n15894_), .Y(new_n15897_));
  AOI21  g14895(.A0(new_n15889_), .A1(new_n15888_), .B0(new_n15897_), .Y(new_n15898_));
  NOR2   g14896(.A(new_n15830_), .B(new_n15809_), .Y(new_n15899_));
  OAI21  g14897(.A0(new_n15824_), .A1(new_n15823_), .B0(new_n15825_), .Y(new_n15900_));
  OAI22  g14898(.A0(new_n15829_), .A1(new_n15826_), .B0(new_n15808_), .B1(new_n15800_), .Y(new_n15901_));
  AOI21  g14899(.A0(new_n15901_), .A1(new_n15900_), .B0(new_n15882_), .Y(new_n15902_));
  AOI221 g14900(.A0(new_n15892_), .A1(new_n15814_), .C0(new_n15895_), .B0(new_n15781_), .B1(new_n15780_), .Y(new_n15903_));
  NOR2   g14901(.A(new_n15896_), .B(new_n15890_), .Y(new_n15904_));
  NOR2   g14902(.A(new_n15904_), .B(new_n15903_), .Y(new_n15905_));
  NOR3   g14903(.A(new_n15905_), .B(new_n15902_), .C(new_n15899_), .Y(new_n15906_));
  AOI22  g14904(.A0(new_n15747_), .A1(new_n15744_), .B0(new_n15716_), .B1(new_n15713_), .Y(new_n15907_));
  OAI221 g14905(.A0(new_n15869_), .A1(new_n15868_), .C0(new_n15907_), .B0(new_n15873_), .B1(new_n15872_), .Y(new_n15908_));
  AOI22  g14906(.A0(new_n15908_), .A1(new_n15838_), .B0(new_n15870_), .B1(new_n15874_), .Y(new_n15909_));
  OAI21  g14907(.A0(new_n15906_), .A1(new_n15898_), .B0(new_n15909_), .Y(new_n15910_));
  OAI21  g14908(.A0(new_n15885_), .A1(new_n15879_), .B0(new_n15910_), .Y(new_n15911_));
  NAND2  g14909(.A(new_n4767_), .B(new_n3557_), .Y(new_n15912_));
  OAI21  g14910(.A0(new_n12239_), .A1(new_n12887_), .B0(new_n12238_), .Y(new_n15913_));
  NAND2  g14911(.A(new_n15913_), .B(new_n15912_), .Y(new_n15914_));
  NOR3   g14912(.A(new_n11196_), .B(new_n11195_), .C(new_n11192_), .Y(new_n15915_));
  AOI21  g14913(.A0(new_n11181_), .A1(new_n11171_), .B0(new_n11188_), .Y(new_n15916_));
  OAI21  g14914(.A0(new_n15916_), .A1(new_n15915_), .B0(new_n11205_), .Y(new_n15917_));
  OAI21  g14915(.A0(new_n12885_), .A1(new_n11218_), .B0(new_n7058_), .Y(new_n15918_));
  INV    g14916(.A(new_n11214_), .Y(new_n15919_));
  NAND3  g14917(.A(new_n15919_), .B(new_n15918_), .C(new_n15917_), .Y(new_n15920_));
  AOI21  g14918(.A0(new_n15918_), .A1(new_n15917_), .B0(new_n15919_), .Y(new_n15921_));
  AOI21  g14919(.A0(new_n15920_), .A1(new_n15914_), .B0(new_n15921_), .Y(new_n15922_));
  XOR2   g14920(.A(new_n12883_), .B(new_n11219_), .Y(new_n15923_));
  NOR2   g14921(.A(new_n12889_), .B(new_n15923_), .Y(new_n15924_));
  OAI22  g14922(.A0(new_n12890_), .A1(new_n12884_), .B0(new_n15924_), .B1(new_n15922_), .Y(new_n15925_));
  NOR2   g14923(.A(new_n13708_), .B(new_n13702_), .Y(new_n15926_));
  XOR2   g14924(.A(new_n14224_), .B(new_n14797_), .Y(new_n15927_));
  OAI21  g14925(.A0(new_n13697_), .A1(new_n15926_), .B0(new_n15927_), .Y(new_n15928_));
  NOR2   g14926(.A(new_n14227_), .B(new_n13697_), .Y(new_n15929_));
  AOI21  g14927(.A0(new_n15928_), .A1(new_n15925_), .B0(new_n15929_), .Y(new_n15930_));
  NAND2  g14928(.A(new_n15107_), .B(new_n14793_), .Y(new_n15931_));
  XOR2   g14929(.A(new_n15099_), .B(new_n15850_), .Y(new_n15932_));
  AOI21  g14930(.A0(new_n14790_), .A1(new_n15931_), .B0(new_n15932_), .Y(new_n15933_));
  NAND2  g14931(.A(new_n15108_), .B(new_n14790_), .Y(new_n15934_));
  OAI21  g14932(.A0(new_n15933_), .A1(new_n15930_), .B0(new_n15934_), .Y(new_n15935_));
  NOR2   g14933(.A(new_n15390_), .B(new_n15380_), .Y(new_n15936_));
  XOR2   g14934(.A(new_n15558_), .B(new_n15853_), .Y(new_n15937_));
  OAI21  g14935(.A0(new_n15376_), .A1(new_n15936_), .B0(new_n15937_), .Y(new_n15938_));
  NOR2   g14936(.A(new_n15561_), .B(new_n15376_), .Y(new_n15939_));
  AOI21  g14937(.A0(new_n15938_), .A1(new_n15935_), .B0(new_n15939_), .Y(new_n15940_));
  NAND2  g14938(.A(new_n15766_), .B(new_n15678_), .Y(new_n15941_));
  XOR2   g14939(.A(new_n15757_), .B(new_n15856_), .Y(new_n15942_));
  AOI21  g14940(.A0(new_n15674_), .A1(new_n15941_), .B0(new_n15942_), .Y(new_n15943_));
  NAND2  g14941(.A(new_n15767_), .B(new_n15674_), .Y(new_n15944_));
  OAI21  g14942(.A0(new_n15943_), .A1(new_n15940_), .B0(new_n15944_), .Y(new_n15945_));
  NAND2  g14943(.A(new_n15878_), .B(new_n15832_), .Y(new_n15946_));
  AOI21  g14944(.A0(new_n15946_), .A1(new_n15945_), .B0(new_n15885_), .Y(new_n15947_));
  OAI21  g14945(.A0(new_n15902_), .A1(new_n15899_), .B0(new_n15905_), .Y(new_n15948_));
  NAND3  g14946(.A(new_n15897_), .B(new_n15889_), .C(new_n15888_), .Y(new_n15949_));
  INV    g14947(.A(new_n15909_), .Y(new_n15950_));
  AOI21  g14948(.A0(new_n15949_), .A1(new_n15948_), .B0(new_n15950_), .Y(new_n15951_));
  NAND3  g14949(.A(new_n15950_), .B(new_n15949_), .C(new_n15948_), .Y(new_n15952_));
  OAI21  g14950(.A0(new_n15951_), .A1(new_n15947_), .B0(new_n15952_), .Y(new_n15953_));
  AOI21  g14951(.A0(new_n15889_), .A1(new_n15888_), .B0(new_n15903_), .Y(new_n15954_));
  NOR2   g14952(.A(new_n15954_), .B(new_n15904_), .Y(new_n15955_));
  NOR3   g14953(.A(new_n15909_), .B(new_n15906_), .C(new_n15898_), .Y(new_n15956_));
  NOR2   g14954(.A(new_n15955_), .B(new_n15956_), .Y(new_n15957_));
  AOI22  g14955(.A0(new_n15957_), .A1(new_n15911_), .B0(new_n15955_), .B1(new_n15953_), .Y(new_n15958_));
  NAND2  g14956(.A(new_n12230_), .B(new_n12886_), .Y(new_n15959_));
  AOI21  g14957(.A0(new_n12883_), .A1(new_n11219_), .B0(new_n12889_), .Y(new_n15960_));
  AOI22  g14958(.A0(new_n15960_), .A1(new_n15959_), .B0(new_n12889_), .B1(new_n12231_), .Y(new_n15961_));
  INV    g14959(.A(\A[1000] ), .Y(new_n15962_));
  NOR3   g14960(.A(new_n11212_), .B(new_n11211_), .C(new_n11209_), .Y(new_n15963_));
  INV    g14961(.A(new_n15963_), .Y(new_n15964_));
  OAI21  g14962(.A0(new_n11212_), .A1(new_n11211_), .B0(new_n11209_), .Y(new_n15965_));
  AOI21  g14963(.A0(new_n15965_), .A1(new_n15964_), .B0(new_n15962_), .Y(new_n15966_));
  OAI21  g14964(.A0(new_n15961_), .A1(new_n15922_), .B0(new_n15966_), .Y(new_n15967_));
  NOR3   g14965(.A(new_n15919_), .B(new_n11208_), .C(new_n11198_), .Y(new_n15968_));
  AOI21  g14966(.A0(new_n15918_), .A1(new_n15917_), .B0(new_n11214_), .Y(new_n15969_));
  OAI21  g14967(.A0(new_n15969_), .A1(new_n15968_), .B0(new_n4771_), .Y(new_n15970_));
  OAI21  g14968(.A0(new_n15921_), .A1(new_n11215_), .B0(new_n15914_), .Y(new_n15971_));
  AOI221 g14969(.A0(new_n15971_), .A1(new_n15970_), .C0(new_n15967_), .B0(new_n15961_), .B1(new_n15922_), .Y(new_n15972_));
  OAI21  g14970(.A0(new_n13708_), .A1(new_n13702_), .B0(new_n15927_), .Y(new_n15973_));
  OAI22  g14971(.A0(new_n15973_), .A1(new_n13697_), .B0(new_n15927_), .B1(new_n13709_), .Y(new_n15974_));
  XOR2   g14972(.A(new_n15974_), .B(new_n15925_), .Y(new_n15975_));
  NAND2  g14973(.A(new_n15975_), .B(new_n15972_), .Y(new_n15976_));
  AOI21  g14974(.A0(new_n15107_), .A1(new_n14793_), .B0(new_n15932_), .Y(new_n15977_));
  AOI22  g14975(.A0(new_n15977_), .A1(new_n14790_), .B0(new_n15932_), .B1(new_n14794_), .Y(new_n15978_));
  XOR2   g14976(.A(new_n15978_), .B(new_n14228_), .Y(new_n15979_));
  NOR2   g14977(.A(new_n15979_), .B(new_n15976_), .Y(new_n15980_));
  OAI21  g14978(.A0(new_n15390_), .A1(new_n15380_), .B0(new_n15937_), .Y(new_n15981_));
  OAI22  g14979(.A0(new_n15981_), .A1(new_n15376_), .B0(new_n15937_), .B1(new_n15391_), .Y(new_n15982_));
  XOR2   g14980(.A(new_n15982_), .B(new_n15935_), .Y(new_n15983_));
  NAND2  g14981(.A(new_n15983_), .B(new_n15980_), .Y(new_n15984_));
  AOI21  g14982(.A0(new_n15766_), .A1(new_n15678_), .B0(new_n15942_), .Y(new_n15985_));
  AOI22  g14983(.A0(new_n15985_), .A1(new_n15674_), .B0(new_n15942_), .B1(new_n15679_), .Y(new_n15986_));
  XOR2   g14984(.A(new_n15986_), .B(new_n15562_), .Y(new_n15987_));
  NOR2   g14985(.A(new_n15987_), .B(new_n15984_), .Y(new_n15988_));
  NAND2  g14986(.A(new_n15831_), .B(new_n15882_), .Y(new_n15989_));
  AOI22  g14987(.A0(new_n15887_), .A1(new_n15886_), .B0(new_n15901_), .B1(new_n15900_), .Y(new_n15990_));
  AOI21  g14988(.A0(new_n15990_), .A1(new_n15778_), .B0(new_n15883_), .Y(new_n15991_));
  AOI22  g14989(.A0(new_n15991_), .A1(new_n15989_), .B0(new_n15883_), .B1(new_n15832_), .Y(new_n15992_));
  XOR2   g14990(.A(new_n15992_), .B(new_n15768_), .Y(new_n15993_));
  NAND2  g14991(.A(new_n15993_), .B(new_n15988_), .Y(new_n15994_));
  AOI21  g14992(.A0(new_n15949_), .A1(new_n15948_), .B0(new_n15909_), .Y(new_n15995_));
  NOR3   g14993(.A(new_n15950_), .B(new_n15906_), .C(new_n15898_), .Y(new_n15996_));
  NOR4   g14994(.A(new_n15996_), .B(new_n15995_), .C(new_n15885_), .D(new_n15879_), .Y(new_n15997_));
  OAI21  g14995(.A0(new_n15906_), .A1(new_n15898_), .B0(new_n15950_), .Y(new_n15998_));
  NAND3  g14996(.A(new_n15909_), .B(new_n15949_), .C(new_n15948_), .Y(new_n15999_));
  AOI21  g14997(.A0(new_n15999_), .A1(new_n15998_), .B0(new_n15947_), .Y(new_n16000_));
  NOR3   g14998(.A(new_n16000_), .B(new_n15997_), .C(new_n15994_), .Y(new_n16001_));
  XOR2   g14999(.A(new_n16001_), .B(new_n15958_), .Y(new_n16002_));
  NOR2   g15000(.A(new_n16000_), .B(new_n15997_), .Y(new_n16003_));
  AOI22  g15001(.A0(new_n15971_), .A1(new_n15970_), .B0(new_n15961_), .B1(new_n15922_), .Y(new_n16004_));
  OAI211 g15002(.A0(new_n15961_), .A1(new_n15922_), .B0(new_n16004_), .B1(new_n15966_), .Y(new_n16005_));
  XOR2   g15003(.A(new_n15961_), .B(new_n15922_), .Y(new_n16006_));
  INV    g15004(.A(new_n15966_), .Y(new_n16007_));
  AOI21  g15005(.A0(new_n15971_), .A1(new_n15970_), .B0(new_n16007_), .Y(new_n16008_));
  OAI21  g15006(.A0(new_n16008_), .A1(new_n16006_), .B0(new_n16005_), .Y(new_n16009_));
  NOR2   g15007(.A(new_n15969_), .B(new_n15968_), .Y(new_n16010_));
  NOR2   g15008(.A(new_n16010_), .B(new_n15914_), .Y(new_n16011_));
  AOI21  g15009(.A0(new_n11216_), .A1(new_n15920_), .B0(new_n4771_), .Y(new_n16012_));
  NOR3   g15010(.A(new_n16012_), .B(new_n16011_), .C(new_n16007_), .Y(new_n16013_));
  AOI21  g15011(.A0(new_n15971_), .A1(new_n15970_), .B0(new_n15966_), .Y(new_n16014_));
  NOR2   g15012(.A(new_n16014_), .B(new_n16013_), .Y(new_n16015_));
  NAND2  g15013(.A(new_n16015_), .B(new_n16009_), .Y(new_n16016_));
  XOR2   g15014(.A(new_n15975_), .B(new_n15972_), .Y(new_n16017_));
  NAND2  g15015(.A(new_n16017_), .B(new_n16016_), .Y(new_n16018_));
  XOR2   g15016(.A(new_n15978_), .B(new_n15930_), .Y(new_n16019_));
  XOR2   g15017(.A(new_n16019_), .B(new_n15976_), .Y(new_n16020_));
  NAND2  g15018(.A(new_n16020_), .B(new_n16018_), .Y(new_n16021_));
  XOR2   g15019(.A(new_n15983_), .B(new_n15980_), .Y(new_n16022_));
  NAND2  g15020(.A(new_n16022_), .B(new_n16021_), .Y(new_n16023_));
  XOR2   g15021(.A(new_n15986_), .B(new_n15940_), .Y(new_n16024_));
  XOR2   g15022(.A(new_n16024_), .B(new_n15984_), .Y(new_n16025_));
  NOR2   g15023(.A(new_n16025_), .B(new_n16023_), .Y(new_n16026_));
  XOR2   g15024(.A(new_n15982_), .B(new_n15109_), .Y(new_n16027_));
  NOR3   g15025(.A(new_n16027_), .B(new_n15979_), .C(new_n15976_), .Y(new_n16028_));
  NAND2  g15026(.A(new_n16024_), .B(new_n16028_), .Y(new_n16029_));
  XOR2   g15027(.A(new_n15992_), .B(new_n15945_), .Y(new_n16030_));
  NAND2  g15028(.A(new_n16030_), .B(new_n16029_), .Y(new_n16031_));
  NAND4  g15029(.A(new_n16031_), .B(new_n16026_), .C(new_n16003_), .D(new_n15994_), .Y(new_n16032_));
  NOR2   g15030(.A(new_n16032_), .B(new_n16002_), .Y(new_n16033_));
  AOI21  g15031(.A0(new_n15952_), .A1(new_n15911_), .B0(new_n15955_), .Y(new_n16034_));
  OAI21  g15032(.A0(new_n15902_), .A1(new_n15899_), .B0(new_n15894_), .Y(new_n16035_));
  OAI21  g15033(.A0(new_n15896_), .A1(new_n15890_), .B0(new_n16035_), .Y(new_n16036_));
  INV    g15034(.A(new_n16001_), .Y(new_n16037_));
  AOI211 g15035(.A0(new_n16036_), .A1(new_n15953_), .B(new_n16037_), .C(new_n15958_), .Y(new_n16038_));
  NAND3  g15036(.A(new_n15993_), .B(new_n15988_), .C(new_n16036_), .Y(new_n16039_));
  NOR3   g15037(.A(new_n16039_), .B(new_n16000_), .C(new_n15997_), .Y(new_n16040_));
  NAND2  g15038(.A(new_n16040_), .B(new_n15953_), .Y(new_n16041_));
  NOR2   g15039(.A(new_n16041_), .B(new_n15958_), .Y(new_n16042_));
  NOR4   g15040(.A(new_n16042_), .B(new_n16038_), .C(new_n16034_), .D(new_n16033_), .Y(new_n16043_));
  INV    g15041(.A(new_n16002_), .Y(new_n16044_));
  XOR2   g15042(.A(new_n16003_), .B(new_n15994_), .Y(new_n16045_));
  XOR2   g15043(.A(new_n16030_), .B(new_n16029_), .Y(new_n16046_));
  XOR2   g15044(.A(new_n16024_), .B(new_n16028_), .Y(new_n16047_));
  NAND3  g15045(.A(new_n16047_), .B(new_n16022_), .C(new_n16021_), .Y(new_n16048_));
  XOR2   g15046(.A(new_n16046_), .B(new_n16048_), .Y(new_n16049_));
  XOR2   g15047(.A(new_n16017_), .B(new_n16016_), .Y(new_n16050_));
  INV    g15048(.A(new_n15965_), .Y(new_n16051_));
  NOR2   g15049(.A(new_n16051_), .B(new_n15963_), .Y(new_n16052_));
  NAND2  g15050(.A(new_n15964_), .B(\A[1000] ), .Y(new_n16053_));
  OAI22  g15051(.A0(new_n16053_), .A1(new_n16051_), .B0(new_n16052_), .B1(\A[1000] ), .Y(new_n16054_));
  INV    g15052(.A(new_n16054_), .Y(new_n16055_));
  NOR2   g15053(.A(new_n16012_), .B(new_n16011_), .Y(new_n16056_));
  NAND3  g15054(.A(new_n15971_), .B(new_n15970_), .C(new_n15966_), .Y(new_n16057_));
  OAI21  g15055(.A0(new_n16056_), .A1(new_n15966_), .B0(new_n16057_), .Y(new_n16058_));
  OAI221 g15056(.A0(new_n16054_), .A1(new_n16058_), .C0(new_n16005_), .B0(new_n16008_), .B1(new_n16006_), .Y(new_n16059_));
  XOR2   g15057(.A(new_n16015_), .B(new_n16009_), .Y(new_n16060_));
  OAI21  g15058(.A0(new_n16060_), .A1(new_n16055_), .B0(new_n16059_), .Y(new_n16061_));
  OAI21  g15059(.A0(new_n16061_), .A1(new_n16050_), .B0(new_n16017_), .Y(new_n16062_));
  NAND2  g15060(.A(new_n16061_), .B(new_n16050_), .Y(new_n16063_));
  AOI22  g15061(.A0(new_n16063_), .A1(new_n16062_), .B0(new_n16017_), .B1(new_n16016_), .Y(new_n16064_));
  NOR2   g15062(.A(new_n16020_), .B(new_n16018_), .Y(new_n16065_));
  OAI211 g15063(.A0(new_n16065_), .A1(new_n16064_), .B0(new_n16022_), .B1(new_n16021_), .Y(new_n16066_));
  NAND2  g15064(.A(new_n16047_), .B(new_n16023_), .Y(new_n16067_));
  AOI21  g15065(.A0(new_n16067_), .A1(new_n16066_), .B0(new_n16049_), .Y(new_n16068_));
  NAND3  g15066(.A(new_n16067_), .B(new_n16066_), .C(new_n16049_), .Y(new_n16069_));
  AOI211 g15067(.A0(new_n16069_), .A1(new_n16046_), .B(new_n16068_), .C(new_n16032_), .Y(new_n16070_));
  NAND4  g15068(.A(new_n16046_), .B(new_n16047_), .C(new_n16022_), .D(new_n16021_), .Y(new_n16071_));
  NOR3   g15069(.A(new_n16045_), .B(new_n16071_), .C(new_n16002_), .Y(new_n16073_));
  OAI21  g15070(.A0(new_n16070_), .A1(new_n16045_), .B0(new_n16073_), .Y(new_n16074_));
  AOI211 g15071(.A0(new_n16070_), .A1(new_n16002_), .B(new_n16045_), .C(new_n16071_), .Y(new_n16075_));
  AOI21  g15072(.A0(new_n16074_), .A1(new_n16044_), .B0(new_n16075_), .Y(new_n16076_));
  NOR4   g15073(.A(new_n16038_), .B(new_n16034_), .C(new_n16032_), .D(new_n16002_), .Y(new_n16077_));
  OAI21  g15074(.A0(new_n16077_), .A1(new_n16076_), .B0(new_n16043_), .Y(maj));
endmodule


