//Converted to Combinational , Module name: s1488 , Timestamp: 2018-12-03T15:51:02.584905 
module s1488 ( CLR, v6, v5, v4, v3, v2, v1, v0, v12, v11, v10, v9, v8, v7, v13_D_20, v13_D_21, v13_D_16, v13_D_22, v13_D_19, v13_D_18, v13_D_11, v13_D_23, v13_D_6, v13_D_15, v13_D_9, v13_D_10, v13_D_8, v13_D_24, v13_D_14, v13_D_7, v13_D_17, v13_D_12, v13_D_13, n55, n60, n65, n70, n75, n80 );
input CLR, v6, v5, v4, v3, v2, v1, v0, v12, v11, v10, v9, v8, v7;
output v13_D_20, v13_D_21, v13_D_16, v13_D_22, v13_D_19, v13_D_18, v13_D_11, v13_D_23, v13_D_6, v13_D_15, v13_D_9, v13_D_10, v13_D_8, v13_D_24, v13_D_14, v13_D_7, v13_D_17, v13_D_12, v13_D_13, n55, n60, n65, n70, n75, n80;
wire n45, n46, n47, n48, n49, n50, n51, n53, n54, n55_1, n56, n57, n58, n60_1, n61, n62, n63, n64, n65_1, n66, n68, n69, n70_1, n71, n72, n73, n74, n75_1, n76, n78, n79, n80_1, n81, n82, n83, n84, n85, n86, n87, n88, n90, n91, n92, n93, n94, n95, n96, n97, n98, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n115, n116, n117, n118, n119, n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n139, n140, n141, n142, n143, n144, n146, n147, n148, n149, n150, n151, n152, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n208, n209, n210, n211, n212, n213, n214, n215, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n241, n242, n243, n244, n245, n246, n247, n248, n249, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416;
INVX1    g000(.A(v7), .Y(n45));
NAND3X1  g001(.A(n45), .B(v10), .C(v3), .Y(n46));
NAND2X1  g002(.A(v11), .B(v12), .Y(n47));
INVX1    g003(.A(v6), .Y(n48));
NOR2X1   g004(.A(v1), .B(n48), .Y(n49));
AND2X1   g005(.A(v8), .B(v9), .Y(n50));
INVX1    g006(.A(n50), .Y(n51));
NOR4X1   g007(.A(n49), .B(n47), .C(n46), .D(n51), .Y(v13_D_20));
OR2X1    g008(.A(v8), .B(v9), .Y(n53));
NAND2X1  g009(.A(v4), .B(v5), .Y(n54));
NOR3X1   g010(.A(n54), .B(n53), .C(v11), .Y(n55_1));
AOI21X1  g011(.A0(n50), .A1(v2), .B0(n55_1), .Y(n56));
NOR2X1   g012(.A(v10), .B(v12), .Y(n57));
INVX1    g013(.A(n57), .Y(n58));
NOR3X1   g014(.A(n58), .B(n56), .C(v7), .Y(v13_D_21));
AND2X1   g015(.A(v3), .B(v6), .Y(n60_1));
NOR2X1   g016(.A(v11), .B(v12), .Y(n61));
NAND4X1  g017(.A(n60_1), .B(n45), .C(v9), .D(n61), .Y(n62));
INVX1    g018(.A(v9), .Y(n63));
AND2X1   g019(.A(v11), .B(v12), .Y(n64));
NAND4X1  g020(.A(v7), .B(n63), .C(v2), .D(n64), .Y(n65_1));
NAND2X1  g021(.A(v8), .B(v10), .Y(n66));
AOI21X1  g022(.A0(n65_1), .A1(n62), .B0(n66), .Y(v13_D_16));
INVX1    g023(.A(v10), .Y(n68));
NOR3X1   g024(.A(n68), .B(v11), .C(v12), .Y(n69));
INVX1    g025(.A(n69), .Y(n70_1));
NAND3X1  g026(.A(v7), .B(v8), .C(v9), .Y(n71));
INVX1    g027(.A(v8), .Y(n72));
NOR4X1   g028(.A(v11), .B(v12), .C(v2), .D(n72), .Y(n73));
NOR2X1   g029(.A(v8), .B(n63), .Y(n74));
AOI21X1  g030(.A0(n74), .A1(v12), .B0(n73), .Y(n75_1));
OR2X1    g031(.A(v7), .B(v10), .Y(n76));
OAI22X1  g032(.A0(n75_1), .A1(n76), .B0(n71), .B1(n70_1), .Y(v13_D_22));
AND2X1   g033(.A(v10), .B(v2), .Y(n78));
AND2X1   g034(.A(v7), .B(v8), .Y(n79));
NAND4X1  g035(.A(n78), .B(n64), .C(n63), .D(n79), .Y(n80_1));
NOR4X1   g036(.A(n68), .B(v12), .C(n48), .D(n51), .Y(n81));
INVX1    g037(.A(v12), .Y(n82));
NOR2X1   g038(.A(v9), .B(v10), .Y(n83));
INVX1    g039(.A(n83), .Y(n84));
NOR4X1   g040(.A(v8), .B(n82), .C(v6), .D(n84), .Y(n85));
INVX1    g041(.A(v3), .Y(n86));
NOR3X1   g042(.A(v7), .B(v11), .C(n86), .Y(n87));
OAI21X1  g043(.A0(n85), .A1(n81), .B0(n87), .Y(n88));
NAND2X1  g044(.A(n88), .B(n80_1), .Y(v13_D_19));
AND2X1   g045(.A(v4), .B(v5), .Y(n90));
NOR2X1   g046(.A(v10), .B(v11), .Y(n91));
NAND4X1  g047(.A(n90), .B(n72), .C(n63), .D(n91), .Y(n92));
NOR3X1   g048(.A(n53), .B(n68), .C(v0), .Y(n93));
NOR3X1   g049(.A(n72), .B(n63), .C(v2), .Y(n94));
OR2X1    g050(.A(v4), .B(v5), .Y(n95));
AND2X1   g051(.A(n95), .B(v11), .Y(n96));
OAI21X1  g052(.A0(n94), .A1(n93), .B0(n96), .Y(n97));
OR2X1    g053(.A(v7), .B(v12), .Y(n98));
AOI21X1  g054(.A0(n97), .A1(n92), .B0(n98), .Y(v13_D_18));
MX2X1    g055(.A(v10), .B(v0), .S0(v11), .Y(n100));
NOR2X1   g056(.A(n100), .B(v9), .Y(n101));
NOR2X1   g057(.A(n101), .B(v8), .Y(n102));
INVX1    g058(.A(v2), .Y(n103));
INVX1    g059(.A(v11), .Y(n104));
MX2X1    g060(.A(n103), .B(n60_1), .S0(n104), .Y(n105));
NOR2X1   g061(.A(n105), .B(n72), .Y(n106));
AOI21X1  g062(.A0(v8), .A1(n104), .B0(n54), .Y(n107));
NOR4X1   g063(.A(n106), .B(n102), .C(v12), .D(n107), .Y(n108));
NOR2X1   g064(.A(n104), .B(v12), .Y(n109));
NOR2X1   g065(.A(v8), .B(v10), .Y(n110));
OR2X1    g066(.A(v10), .B(v11), .Y(n111));
AOI21X1  g067(.A0(n111), .A1(v9), .B0(n72), .Y(n112));
AOI21X1  g068(.A0(n110), .A1(n109), .B0(n112), .Y(n113));
OAI21X1  g069(.A0(n108), .A1(v7), .B0(n113), .Y(v13_D_11));
NAND4X1  g070(.A(v10), .B(v11), .C(v12), .D(v9), .Y(n115));
INVX1    g071(.A(v0), .Y(n116));
NOR4X1   g072(.A(n104), .B(v12), .C(n116), .D(n68), .Y(n117));
NOR3X1   g073(.A(n111), .B(n82), .C(n48), .Y(n118));
OAI21X1  g074(.A0(n118), .A1(n117), .B0(n63), .Y(n119));
NOR2X1   g075(.A(v7), .B(v8), .Y(n120));
INVX1    g076(.A(n120), .Y(n121));
AOI21X1  g077(.A0(n119), .A1(n115), .B0(n121), .Y(v13_D_23));
AND2X1   g078(.A(v9), .B(v12), .Y(n123));
NOR2X1   g079(.A(n45), .B(v10), .Y(n124));
MX2X1    g080(.A(n111), .B(n124), .S0(n82), .Y(n125));
AOI22X1  g081(.A0(n123), .A1(n91), .B0(n63), .B1(n125), .Y(n126));
OR2X1    g082(.A(n78), .B(v11), .Y(n127));
OAI21X1  g083(.A0(n63), .A1(v2), .B0(v11), .Y(n128));
AOI21X1  g084(.A0(n128), .A1(n127), .B0(n72), .Y(n129));
INVX1    g085(.A(v5), .Y(n130));
OAI21X1  g086(.A0(v4), .A1(n130), .B0(n68), .Y(n131));
AOI21X1  g087(.A0(n131), .A1(n82), .B0(v11), .Y(n132));
INVX1    g088(.A(n110), .Y(n133));
AOI21X1  g089(.A0(n133), .A1(n109), .B0(n63), .Y(n134));
NAND2X1  g090(.A(v10), .B(v12), .Y(n135));
INVX1    g091(.A(n135), .Y(n136));
NOR4X1   g092(.A(n134), .B(n132), .C(n129), .D(n136), .Y(n137));
OAI22X1  g093(.A0(n126), .A1(n72), .B0(v7), .B1(n137), .Y(v13_D_6));
INVX1    g094(.A(v4), .Y(n139));
INVX1    g095(.A(n53), .Y(n140));
NOR4X1   g096(.A(n63), .B(n104), .C(v2), .D(n72), .Y(n141));
NAND2X1  g097(.A(v10), .B(v11), .Y(n142));
OAI21X1  g098(.A0(n142), .A1(v0), .B0(n111), .Y(n143));
AOI21X1  g099(.A0(n143), .A1(n140), .B0(n141), .Y(n144));
NOR4X1   g100(.A(n98), .B(n139), .C(v5), .D(n144), .Y(v13_D_15));
INVX1    g101(.A(n79), .Y(n146));
OAI22X1  g102(.A0(n91), .A1(n146), .B0(v8), .B1(n142), .Y(n147));
NAND2X1  g103(.A(n147), .B(v9), .Y(n148));
NAND2X1  g104(.A(v11), .B(v0), .Y(n149));
NAND2X1  g105(.A(v8), .B(n103), .Y(n150));
OAI22X1  g106(.A0(n149), .A1(v8), .B0(v9), .B1(n150), .Y(n151));
NAND3X1  g107(.A(n151), .B(n45), .C(v10), .Y(n152));
AOI21X1  g108(.A0(n152), .A1(n148), .B0(v12), .Y(v13_D_9));
NAND2X1  g109(.A(n63), .B(v12), .Y(n154));
NOR2X1   g110(.A(v7), .B(v2), .Y(n155));
OR2X1    g111(.A(n83), .B(v12), .Y(n156));
OAI22X1  g112(.A0(n155), .A1(n156), .B0(n154), .B1(n68), .Y(n157));
AOI21X1  g113(.A0(n135), .A1(n63), .B0(n57), .Y(n158));
NOR3X1   g114(.A(n158), .B(n45), .C(v11), .Y(n159));
AOI21X1  g115(.A0(n157), .A1(v11), .B0(n159), .Y(n160));
AOI22X1  g116(.A0(n78), .A1(n104), .B0(n72), .B1(n100), .Y(n161));
NOR3X1   g117(.A(n161), .B(v7), .C(v9), .Y(n162));
XOR2X1   g118(.A(v9), .B(v10), .Y(n163));
NAND2X1  g119(.A(n72), .B(v11), .Y(n164));
AOI22X1  g120(.A0(n50), .A1(v11), .B0(n63), .B1(n120), .Y(n165));
OAI22X1  g121(.A0(n164), .A1(n163), .B0(n54), .B1(n165), .Y(n166));
OAI21X1  g122(.A0(n166), .A1(n162), .B0(n82), .Y(n167));
OAI21X1  g123(.A0(n160), .A1(n72), .B0(n167), .Y(v13_D_10));
OAI21X1  g124(.A0(v12), .A1(v0), .B0(v11), .Y(n169));
AND2X1   g125(.A(n169), .B(n63), .Y(n170));
AOI21X1  g126(.A0(n170), .A1(n70_1), .B0(v8), .Y(n171));
NOR2X1   g127(.A(n68), .B(v12), .Y(n172));
INVX1    g128(.A(n78), .Y(n173));
OAI22X1  g129(.A0(n172), .A1(n72), .B0(v12), .B1(n173), .Y(n174));
AND2X1   g130(.A(n174), .B(n104), .Y(n175));
AOI21X1  g131(.A0(n63), .A1(v11), .B0(v12), .Y(n176));
NOR2X1   g132(.A(n176), .B(v10), .Y(n177));
NOR2X1   g133(.A(v4), .B(n130), .Y(n178));
AOI22X1  g134(.A0(v9), .A1(n103), .B0(v11), .B1(n72), .Y(n179));
OAI22X1  g135(.A0(n178), .A1(n179), .B0(n109), .B1(n63), .Y(n180));
NOR4X1   g136(.A(n177), .B(n175), .C(n171), .D(n180), .Y(n181));
MX2X1    g137(.A(v12), .B(n104), .S0(v9), .Y(n182));
NOR2X1   g138(.A(n72), .B(v10), .Y(n183));
NAND2X1  g139(.A(v11), .B(n82), .Y(n184));
AOI21X1  g140(.A0(n47), .A1(n63), .B0(n61), .Y(n185));
OAI22X1  g141(.A0(n133), .A1(n184), .B0(n66), .B1(n185), .Y(n186));
AOI22X1  g142(.A0(n183), .A1(n182), .B0(v7), .B1(n186), .Y(n187));
OAI21X1  g143(.A0(n181), .A1(v7), .B0(n187), .Y(v13_D_8));
AND2X1   g144(.A(n60_1), .B(n50), .Y(n189));
OR2X1    g145(.A(n135), .B(v11), .Y(n190));
AOI21X1  g146(.A0(n61), .A1(n130), .B0(n64), .Y(n191));
OAI21X1  g147(.A0(n191), .A1(v10), .B0(n190), .Y(n192));
AOI22X1  g148(.A0(n189), .A1(n69), .B0(n140), .B1(n192), .Y(n193));
NAND4X1  g149(.A(v10), .B(v11), .C(n130), .D(n120), .Y(n194));
NAND4X1  g150(.A(v8), .B(n68), .C(n103), .D(v7), .Y(n195));
OR2X1    g151(.A(v9), .B(v12), .Y(n196));
OR2X1    g152(.A(n196), .B(v0), .Y(n197));
AOI21X1  g153(.A0(n195), .A1(n194), .B0(n197), .Y(n198));
NOR4X1   g154(.A(v9), .B(n68), .C(n82), .D(n45), .Y(n199));
NOR4X1   g155(.A(n63), .B(v12), .C(v5), .D(n124), .Y(n200));
NOR2X1   g156(.A(n200), .B(n199), .Y(n201));
XOR2X1   g157(.A(n50), .B(v10), .Y(n202));
NOR2X1   g158(.A(n45), .B(v12), .Y(n203));
INVX1    g159(.A(n203), .Y(n204));
OAI22X1  g160(.A0(n202), .A1(n204), .B0(n201), .B1(n150), .Y(n205));
AOI21X1  g161(.A0(n205), .A1(v11), .B0(n198), .Y(n206));
OAI21X1  g162(.A0(n193), .A1(v7), .B0(n206), .Y(v13_D_24));
AOI21X1  g163(.A0(v10), .A1(n116), .B0(n104), .Y(n208));
OR2X1    g164(.A(n208), .B(v9), .Y(n209));
AOI22X1  g165(.A0(v10), .A1(n104), .B0(v2), .B1(v8), .Y(n210));
NAND4X1  g166(.A(n95), .B(n54), .C(n82), .D(n210), .Y(n211));
AOI21X1  g167(.A0(n209), .A1(n72), .B0(n211), .Y(n212));
NOR2X1   g168(.A(v9), .B(n68), .Y(n213));
OAI21X1  g169(.A0(n213), .A1(n104), .B0(n72), .Y(n214));
AOI21X1  g170(.A0(n214), .A1(n203), .B0(n112), .Y(n215));
OAI21X1  g171(.A0(n212), .A1(v7), .B0(n215), .Y(v13_D_14));
NOR2X1   g172(.A(n72), .B(v11), .Y(n217));
INVX1    g173(.A(n217), .Y(n218));
INVX1    g174(.A(n154), .Y(n219));
AOI22X1  g175(.A0(n84), .A1(n82), .B0(n68), .B1(n219), .Y(n220));
OR4X1    g176(.A(n63), .B(n104), .C(v12), .D(n183), .Y(n221));
OAI21X1  g177(.A0(n220), .A1(n218), .B0(n221), .Y(n222));
OAI21X1  g178(.A0(n47), .A1(v10), .B0(n70_1), .Y(n223));
AOI22X1  g179(.A0(n78), .A1(n61), .B0(n72), .B1(n223), .Y(n224));
AOI21X1  g180(.A0(n139), .A1(v5), .B0(v12), .Y(n225));
OAI21X1  g181(.A0(n141), .A1(n93), .B0(n225), .Y(n226));
OAI21X1  g182(.A0(n224), .A1(v9), .B0(n226), .Y(n227));
MX2X1    g183(.A(n222), .B(n227), .S0(n45), .Y(v13_D_7));
OR4X1    g184(.A(n121), .B(n111), .C(n54), .D(n196), .Y(n229));
AND2X1   g185(.A(v8), .B(v11), .Y(n230));
INVX1    g186(.A(n230), .Y(n231));
AND2X1   g187(.A(v9), .B(v11), .Y(n232));
MX2X1    g188(.A(n116), .B(n63), .S0(n104), .Y(n233));
AOI21X1  g189(.A0(n233), .A1(n45), .B0(n232), .Y(n234));
OAI22X1  g190(.A0(n231), .A1(n83), .B0(n68), .B1(n234), .Y(n235));
INVX1    g191(.A(n142), .Y(n236));
AOI21X1  g192(.A0(n236), .A1(n63), .B0(n82), .Y(n237));
OAI22X1  g193(.A0(n184), .A1(v10), .B0(n72), .B1(n237), .Y(n238));
AOI22X1  g194(.A0(n235), .A1(n82), .B0(v7), .B1(n238), .Y(n239));
OAI21X1  g195(.A0(n239), .A1(n103), .B0(n229), .Y(v13_D_17));
NAND2X1  g196(.A(v9), .B(v10), .Y(n241));
NOR3X1   g197(.A(n241), .B(n104), .C(v12), .Y(n242));
AOI22X1  g198(.A0(n68), .A1(n90), .B0(v11), .B1(v0), .Y(n243));
OAI21X1  g199(.A0(n243), .A1(v12), .B0(n190), .Y(n244));
AOI21X1  g200(.A0(n244), .A1(n63), .B0(n242), .Y(n245));
OAI22X1  g201(.A0(n184), .A1(n84), .B0(v7), .B1(n245), .Y(n246));
NOR2X1   g202(.A(v12), .B(n103), .Y(n247));
AOI22X1  g203(.A0(n219), .A1(v10), .B0(n84), .B1(n247), .Y(n248));
OAI21X1  g204(.A0(n248), .A1(n104), .B0(n204), .Y(n249));
MX2X1    g205(.A(n246), .B(n249), .S0(v8), .Y(v13_D_12));
MX2X1    g206(.A(v11), .B(n47), .S0(n68), .Y(n251));
OAI21X1  g207(.A0(n251), .A1(v8), .B0(n70_1), .Y(n252));
NOR3X1   g208(.A(n208), .B(v8), .C(v9), .Y(n253));
OAI21X1  g209(.A0(n253), .A1(n141), .B0(n90), .Y(n254));
NAND3X1  g210(.A(n230), .B(n84), .C(v2), .Y(n255));
AOI21X1  g211(.A0(n255), .A1(n254), .B0(v12), .Y(n256));
AOI21X1  g212(.A0(n252), .A1(n63), .B0(n256), .Y(n257));
NAND4X1  g213(.A(v11), .B(n82), .C(v1), .D(v9), .Y(n258));
INVX1    g214(.A(v1), .Y(n259));
OAI21X1  g215(.A0(n72), .A1(n104), .B0(n98), .Y(n260));
AOI22X1  g216(.A0(n64), .A1(v8), .B0(n259), .B1(n260), .Y(n261));
OAI21X1  g217(.A0(n261), .A1(v9), .B0(n258), .Y(n262));
AOI22X1  g218(.A0(n69), .A1(v9), .B0(n47), .B1(n83), .Y(n263));
OAI22X1  g219(.A0(n133), .A1(n184), .B0(n72), .B1(n263), .Y(n264));
AOI22X1  g220(.A0(n262), .A1(v10), .B0(v7), .B1(n264), .Y(n265));
OAI21X1  g221(.A0(n257), .A1(v7), .B0(n265), .Y(v13_D_13));
INVX1    g222(.A(CLR), .Y(n267));
NAND4X1  g223(.A(n68), .B(v11), .C(n82), .D(v9), .Y(n268));
AOI21X1  g224(.A0(n54), .A1(n103), .B0(n184), .Y(n269));
OAI21X1  g225(.A0(n269), .A1(n63), .B0(v10), .Y(n270));
AOI21X1  g226(.A0(n270), .A1(n268), .B0(n72), .Y(n271));
NOR3X1   g227(.A(v9), .B(v11), .C(v12), .Y(n272));
NAND4X1  g228(.A(n259), .B(v3), .C(v6), .D(v8), .Y(n273));
OAI22X1  g229(.A0(n196), .A1(n54), .B0(n47), .B1(n273), .Y(n274));
AOI21X1  g230(.A0(n274), .A1(n116), .B0(n272), .Y(n275));
NAND4X1  g231(.A(n63), .B(v12), .C(v6), .D(n91), .Y(n276));
OAI21X1  g232(.A0(n142), .A1(n63), .B0(n276), .Y(n277));
NAND4X1  g233(.A(v10), .B(v11), .C(v0), .D(v8), .Y(n278));
OAI22X1  g234(.A0(n111), .A1(n53), .B0(n49), .B1(n278), .Y(n279));
AND2X1   g235(.A(v12), .B(v3), .Y(n280));
AOI22X1  g236(.A0(n279), .A1(n280), .B0(n277), .B1(n72), .Y(n281));
OAI21X1  g237(.A0(n275), .A1(n68), .B0(n281), .Y(n282));
OAI21X1  g238(.A0(n282), .A1(n271), .B0(n45), .Y(n283));
AOI22X1  g239(.A0(n109), .A1(n72), .B0(n217), .B1(n196), .Y(n284));
OAI22X1  g240(.A0(n241), .A1(n184), .B0(v10), .B1(n284), .Y(n285));
NOR3X1   g241(.A(n142), .B(n72), .C(v9), .Y(n286));
NOR3X1   g242(.A(n98), .B(n259), .C(n48), .Y(n287));
NOR3X1   g243(.A(n111), .B(v8), .C(n63), .Y(n288));
AOI21X1  g244(.A0(n288), .A1(n287), .B0(n286), .Y(n289));
OAI22X1  g245(.A0(n196), .A1(n66), .B0(v2), .B1(n289), .Y(n290));
AOI21X1  g246(.A0(n285), .A1(v7), .B0(n290), .Y(n291));
AOI21X1  g247(.A0(n291), .A1(n283), .B0(n267), .Y(n55));
MX2X1    g248(.A(v10), .B(n90), .S0(v9), .Y(n293));
NAND3X1  g249(.A(n293), .B(n82), .C(n103), .Y(n294));
NAND3X1  g250(.A(v0), .B(n259), .C(v6), .Y(n295));
AND2X1   g251(.A(n123), .B(v3), .Y(n296));
OAI21X1  g252(.A0(v9), .A1(v3), .B0(n109), .Y(n297));
AOI22X1  g253(.A0(n296), .A1(n295), .B0(n68), .B1(n297), .Y(n298));
AOI21X1  g254(.A0(n298), .A1(n294), .B0(n72), .Y(n299));
NAND3X1  g255(.A(v9), .B(n68), .C(n259), .Y(n300));
OAI21X1  g256(.A0(n142), .A1(v9), .B0(n300), .Y(n301));
NAND3X1  g257(.A(n301), .B(n72), .C(n82), .Y(n302));
NAND2X1  g258(.A(n72), .B(v9), .Y(n303));
OAI22X1  g259(.A0(n303), .A1(n58), .B0(v11), .B1(n154), .Y(n304));
NOR2X1   g260(.A(n251), .B(n63), .Y(n305));
AOI21X1  g261(.A0(n304), .A1(n48), .B0(n305), .Y(n306));
NAND3X1  g262(.A(n306), .B(n302), .C(n190), .Y(n307));
OAI21X1  g263(.A0(n307), .A1(n299), .B0(n45), .Y(n308));
NAND4X1  g264(.A(n64), .B(n63), .C(v10), .D(n79), .Y(n309));
NAND3X1  g265(.A(n57), .B(n45), .C(v9), .Y(n310));
AOI21X1  g266(.A0(n310), .A1(n309), .B0(n103), .Y(n311));
AOI22X1  g267(.A0(n110), .A1(v11), .B0(n217), .B1(n213), .Y(n312));
AOI22X1  g268(.A0(n74), .A1(n109), .B0(n217), .B1(v12), .Y(n313));
OAI22X1  g269(.A0(n312), .A1(n204), .B0(v10), .B1(n313), .Y(n314));
NOR2X1   g270(.A(n314), .B(n311), .Y(n315));
AOI21X1  g271(.A0(n315), .A1(n308), .B0(n267), .Y(n60));
NOR2X1   g272(.A(n47), .B(n86), .Y(n317));
AOI22X1  g273(.A0(n295), .A1(n317), .B0(n61), .B1(n48), .Y(n318));
OR2X1    g274(.A(n318), .B(n63), .Y(n319));
AOI21X1  g275(.A0(n90), .A1(n47), .B0(v10), .Y(n320));
OAI21X1  g276(.A0(n247), .A1(v11), .B0(v10), .Y(n321));
AOI21X1  g277(.A0(n321), .A1(n63), .B0(n320), .Y(n322));
AOI21X1  g278(.A0(n322), .A1(n319), .B0(n72), .Y(n323));
NOR2X1   g279(.A(n54), .B(v12), .Y(n324));
MX2X1    g280(.A(n68), .B(n50), .S0(n82), .Y(n325));
AOI22X1  g281(.A0(n324), .A1(n83), .B0(n86), .B1(n325), .Y(n326));
NOR2X1   g282(.A(v8), .B(n82), .Y(n327));
AOI21X1  g283(.A0(n104), .A1(v6), .B0(v9), .Y(n328));
OAI22X1  g284(.A0(n142), .A1(v9), .B0(v10), .B1(n328), .Y(n329));
MX2X1    g285(.A(v8), .B(n74), .S0(v10), .Y(n330));
AOI22X1  g286(.A0(n329), .A1(n327), .B0(n247), .B1(n330), .Y(n331));
OAI21X1  g287(.A0(n326), .A1(v11), .B0(n331), .Y(n332));
OAI21X1  g288(.A0(n332), .A1(n323), .B0(n45), .Y(n333));
NAND3X1  g289(.A(n63), .B(v10), .C(v12), .Y(n334));
OAI21X1  g290(.A0(n219), .A1(v10), .B0(n334), .Y(n335));
AOI22X1  g291(.A0(n232), .A1(n203), .B0(n217), .B1(n335), .Y(n336));
AOI21X1  g292(.A0(n336), .A1(n333), .B0(n267), .Y(n65));
NAND4X1  g293(.A(v10), .B(n104), .C(n82), .D(n63), .Y(n338));
AOI21X1  g294(.A0(v12), .A1(v1), .B0(v9), .Y(n339));
NOR3X1   g295(.A(n339), .B(n72), .C(n104), .Y(n340));
NOR4X1   g296(.A(n63), .B(v11), .C(v12), .D(v8), .Y(n341));
OAI21X1  g297(.A0(n341), .A1(n340), .B0(n68), .Y(n342));
AOI21X1  g298(.A0(n342), .A1(n338), .B0(n103), .Y(n343));
INVX1    g299(.A(n61), .Y(n344));
OAI22X1  g300(.A0(n303), .A1(n344), .B0(n47), .B1(n150), .Y(n345));
AOI22X1  g301(.A0(n272), .A1(n90), .B0(n259), .B1(n345), .Y(n346));
NAND4X1  g302(.A(v9), .B(n82), .C(n48), .D(n91), .Y(n347));
NAND2X1  g303(.A(v11), .B(n116), .Y(n348));
AOI22X1  g304(.A0(n172), .A1(n348), .B0(n64), .B1(n68), .Y(n349));
OAI21X1  g305(.A0(n349), .A1(v9), .B0(n347), .Y(n350));
NOR3X1   g306(.A(n196), .B(v8), .C(n68), .Y(n351));
NOR4X1   g307(.A(n63), .B(v10), .C(n104), .D(n72), .Y(n352));
OAI21X1  g308(.A0(n352), .A1(n351), .B0(n54), .Y(n353));
NOR3X1   g309(.A(n111), .B(v12), .C(n86), .Y(n354));
AND2X1   g310(.A(n142), .B(n123), .Y(n355));
OAI21X1  g311(.A0(n355), .A1(n354), .B0(v8), .Y(n356));
NAND4X1  g312(.A(v10), .B(n104), .C(v12), .D(v9), .Y(n357));
NAND3X1  g313(.A(n357), .B(n356), .C(n353), .Y(n358));
AOI21X1  g314(.A0(n350), .A1(n72), .B0(n358), .Y(n359));
OAI21X1  g315(.A0(n346), .A1(v10), .B0(n359), .Y(n360));
OAI21X1  g316(.A0(n360), .A1(n343), .B0(n45), .Y(n361));
NOR4X1   g317(.A(v8), .B(n82), .C(v6), .D(v7), .Y(n362));
NOR2X1   g318(.A(n72), .B(v12), .Y(n363));
OAI21X1  g319(.A0(n363), .A1(n362), .B0(n86), .Y(n364));
OAI21X1  g320(.A0(n218), .A1(v12), .B0(n364), .Y(n365));
MX2X1    g321(.A(v10), .B(n173), .S0(v11), .Y(n366));
AOI22X1  g322(.A0(n111), .A1(n82), .B0(n63), .B1(n366), .Y(n367));
OAI22X1  g323(.A0(n213), .A1(n184), .B0(n72), .B1(n367), .Y(n368));
AOI22X1  g324(.A0(n365), .A1(n83), .B0(v7), .B1(n368), .Y(n369));
AOI21X1  g325(.A0(n369), .A1(n361), .B0(n267), .Y(n70));
NOR2X1   g326(.A(n68), .B(v11), .Y(n371));
OR2X1    g327(.A(v3), .B(v6), .Y(n372));
AOI21X1  g328(.A0(n372), .A1(n104), .B0(v10), .Y(n373));
OAI21X1  g329(.A0(n373), .A1(n371), .B0(v12), .Y(n374));
AOI22X1  g330(.A0(n143), .A1(n324), .B0(n70_1), .B1(v9), .Y(n375));
AOI21X1  g331(.A0(n375), .A1(n374), .B0(v8), .Y(n376));
NOR3X1   g332(.A(n47), .B(v10), .C(v1), .Y(n377));
OAI21X1  g333(.A0(n135), .A1(v3), .B0(n63), .Y(n378));
AOI21X1  g334(.A0(n378), .A1(n72), .B0(n377), .Y(n379));
AOI22X1  g335(.A0(n83), .A1(n363), .B0(n64), .B1(v9), .Y(n380));
OAI21X1  g336(.A0(n379), .A1(n103), .B0(n380), .Y(n381));
OAI21X1  g337(.A0(n381), .A1(n376), .B0(n45), .Y(n382));
MX2X1    g338(.A(n63), .B(v8), .S0(n68), .Y(n383));
AOI21X1  g339(.A0(n63), .A1(v12), .B0(n104), .Y(n384));
MX2X1    g340(.A(n184), .B(n384), .S0(n68), .Y(n385));
OAI22X1  g341(.A0(n383), .A1(n184), .B0(n72), .B1(n385), .Y(n386));
OAI22X1  g342(.A0(n184), .A1(n68), .B0(n45), .B1(n154), .Y(n387));
NAND3X1  g343(.A(n90), .B(v8), .C(n82), .Y(n388));
NAND3X1  g344(.A(n68), .B(v12), .C(v1), .Y(n389));
NAND2X1  g345(.A(n389), .B(n388), .Y(n390));
NOR2X1   g346(.A(v7), .B(n104), .Y(n391));
AOI22X1  g347(.A0(n390), .A1(n391), .B0(n387), .B1(v8), .Y(n392));
AOI22X1  g348(.A0(n63), .A1(v12), .B0(v3), .B1(n57), .Y(n393));
OAI22X1  g349(.A0(n392), .A1(v2), .B0(n218), .B1(n393), .Y(n394));
AOI21X1  g350(.A0(n386), .A1(v7), .B0(n394), .Y(n395));
AOI21X1  g351(.A0(n395), .A1(n382), .B0(n267), .Y(n75));
NOR3X1   g352(.A(v8), .B(v11), .C(v12), .Y(n397));
AOI21X1  g353(.A0(n64), .A1(v6), .B0(n397), .Y(n398));
OR2X1    g354(.A(n398), .B(v1), .Y(n399));
OAI21X1  g355(.A0(n72), .A1(v11), .B0(v10), .Y(n400));
OR2X1    g356(.A(n397), .B(n64), .Y(n401));
AOI22X1  g357(.A0(n400), .A1(v12), .B0(n86), .B1(n401), .Y(n402));
AOI21X1  g358(.A0(n402), .A1(n399), .B0(n63), .Y(n403));
NOR3X1   g359(.A(v9), .B(n68), .C(v0), .Y(n404));
NAND3X1  g360(.A(n404), .B(n109), .C(n90), .Y(n405));
AOI21X1  g361(.A0(v10), .A1(n82), .B0(n104), .Y(n406));
AOI21X1  g362(.A0(n68), .A1(v6), .B0(n344), .Y(n407));
OAI21X1  g363(.A0(n407), .A1(n406), .B0(v9), .Y(n408));
AOI21X1  g364(.A0(n408), .A1(n405), .B0(v8), .Y(n409));
OAI21X1  g365(.A0(n409), .A1(n403), .B0(n45), .Y(n410));
OAI22X1  g366(.A0(n236), .A1(n154), .B0(n111), .B1(n63), .Y(n411));
NOR2X1   g367(.A(v8), .B(v11), .Y(n412));
AOI21X1  g368(.A0(n230), .A1(n90), .B0(n412), .Y(n413));
NAND3X1  g369(.A(n45), .B(v9), .C(n82), .Y(n414));
OAI22X1  g370(.A0(n413), .A1(n414), .B0(n154), .B1(n146), .Y(n415));
AOI22X1  g371(.A0(n411), .A1(n79), .B0(n103), .B1(n415), .Y(n416));
AOI21X1  g372(.A0(n416), .A1(n410), .B0(n267), .Y(n80));
endmodule
