//Converted to Combinational , Module name: s386 , Timestamp: 2018-12-03T15:51:01.495559 
module s386 ( v6, v5, v4, v3, v2, v1, v0, v12, v11, v10, v9, v8, v7, v13_D_12, v13_D_11, v13_D_10, v13_D_9, v13_D_8, v13_D_7, v13_D_6, n29, n34, n39, n44, n49, n54 );
input v6, v5, v4, v3, v2, v1, v0, v12, v11, v10, v9, v8, v7;
output v13_D_12, v13_D_11, v13_D_10, v13_D_9, v13_D_8, v13_D_7, v13_D_6, n29, n34, n39, n44, n49, n54;
wire n32, n33, n34_1, n35, n36, n37, n38, n40, n41, n42, n43, n44_1, n45, n46, n47, n48, n49_1, n50, n51, n52, n54_1, n55, n56, n58, n59, n60, n61, n62, n64, n65, n67, n68, n69, n70, n71, n72, n74, n75, n76, n77, n78, n79, n80, n81, n83, n84, n85, n86, n87, n89, n90, n91, n92, n94, n95, n96, n97, n98, n99, n101, n102, n103, n104, n105, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n118;
INVX1    g00(.A(v0), .Y(n32));
INVX1    g01(.A(v12), .Y(n33));
INVX1    g02(.A(v7), .Y(n34_1));
NAND4X1  g03(.A(n33), .B(n32), .C(v5), .D(n34_1), .Y(n35));
INVX1    g04(.A(v11), .Y(n36));
INVX1    g05(.A(v8), .Y(n37));
NAND4X1  g06(.A(v9), .B(v10), .C(n36), .D(n37), .Y(n38));
NOR2X1   g07(.A(n38), .B(n35), .Y(v13_D_12));
INVX1    g08(.A(v10), .Y(n40));
NOR2X1   g09(.A(n40), .B(v11), .Y(n41));
NOR3X1   g10(.A(v11), .B(v3), .C(v4), .Y(n42));
AOI21X1  g11(.A0(v7), .A1(v11), .B0(n42), .Y(n43));
NAND2X1  g12(.A(v8), .B(n33), .Y(n44_1));
NOR2X1   g13(.A(v7), .B(v8), .Y(n45));
OAI21X1  g14(.A0(n45), .A1(n33), .B0(v1), .Y(n46));
OAI21X1  g15(.A0(n44_1), .A1(n43), .B0(n46), .Y(n47));
OR2X1    g16(.A(v7), .B(v8), .Y(n48));
NOR3X1   g17(.A(n48), .B(v12), .C(n32), .Y(n49_1));
AOI22X1  g18(.A0(n47), .A1(n40), .B0(n41), .B1(n49_1), .Y(n50));
OAI22X1  g19(.A0(v8), .A1(v7), .B0(v9), .B1(v12), .Y(n51));
NAND3X1  g20(.A(n51), .B(n40), .C(n32), .Y(n52));
OAI21X1  g21(.A0(n50), .A1(v9), .B0(n52), .Y(v13_D_11));
INVX1    g22(.A(v9), .Y(n54_1));
AOI21X1  g23(.A0(v0), .A1(v5), .B0(n40), .Y(n55));
NAND4X1  g24(.A(n36), .B(n33), .C(v1), .D(n34_1), .Y(n56));
NOR4X1   g25(.A(n55), .B(v8), .C(n54_1), .D(n56), .Y(v13_D_10));
INVX1    g26(.A(v3), .Y(n58));
NOR2X1   g27(.A(v10), .B(v1), .Y(n59));
NAND4X1  g28(.A(v8), .B(n58), .C(v4), .D(n59), .Y(n60));
NAND3X1  g29(.A(n37), .B(v10), .C(v0), .Y(n61));
OR4X1    g30(.A(v9), .B(v11), .C(v12), .D(v7), .Y(n62));
AOI21X1  g31(.A0(n61), .A1(n60), .B0(n62), .Y(v13_D_9));
OR4X1    g32(.A(v11), .B(n32), .C(v6), .D(v7), .Y(n64));
NAND4X1  g33(.A(n54_1), .B(v10), .C(n33), .D(n37), .Y(n65));
NOR2X1   g34(.A(n65), .B(n64), .Y(v13_D_8));
NOR4X1   g35(.A(v11), .B(v3), .C(v4), .D(n37), .Y(n67));
INVX1    g36(.A(n67), .Y(n68));
NAND3X1  g37(.A(v7), .B(n37), .C(v11), .Y(n69));
INVX1    g38(.A(v1), .Y(n70));
NOR2X1   g39(.A(v9), .B(v10), .Y(n71));
NAND4X1  g40(.A(n33), .B(v0), .C(n70), .D(n71), .Y(n72));
AOI21X1  g41(.A0(n69), .A1(n68), .B0(n72), .Y(v13_D_7));
NAND4X1  g42(.A(v11), .B(v12), .C(v5), .D(n45), .Y(n74));
OR2X1    g43(.A(v11), .B(v12), .Y(n75));
INVX1    g44(.A(n75), .Y(n76));
INVX1    g45(.A(v2), .Y(n77));
AOI22X1  g46(.A0(v8), .A1(n58), .B0(n77), .B1(n34_1), .Y(n78));
AND2X1   g47(.A(v7), .B(v4), .Y(n79));
OAI21X1  g48(.A0(n79), .A1(n78), .B0(n76), .Y(n80));
NAND3X1  g49(.A(n71), .B(v0), .C(n70), .Y(n81));
AOI21X1  g50(.A0(n80), .A1(n74), .B0(n81), .Y(v13_D_6));
NAND4X1  g51(.A(v8), .B(v11), .C(n33), .D(v7), .Y(n83));
NAND2X1  g52(.A(v11), .B(v12), .Y(n84));
NOR2X1   g53(.A(n84), .B(v8), .Y(n85));
NOR4X1   g54(.A(n37), .B(n77), .C(n58), .D(n75), .Y(n86));
OAI21X1  g55(.A0(n86), .A1(n85), .B0(n34_1), .Y(n87));
AOI21X1  g56(.A0(n87), .A1(n83), .B0(n81), .Y(n29));
OAI21X1  g57(.A0(n67), .A1(v7), .B0(n33), .Y(n89));
OR2X1    g58(.A(v7), .B(v5), .Y(n90));
OAI22X1  g59(.A0(n84), .A1(n90), .B0(n75), .B1(n77), .Y(n91));
NAND2X1  g60(.A(n91), .B(n37), .Y(n92));
AOI21X1  g61(.A0(n92), .A1(n89), .B0(n81), .Y(n34));
NOR4X1   g62(.A(v8), .B(n40), .C(v11), .D(n90), .Y(n94));
OR2X1    g63(.A(n94), .B(n71), .Y(n95));
AOI22X1  g64(.A0(n71), .A1(n32), .B0(v1), .B1(n95), .Y(n96));
OAI21X1  g65(.A0(v11), .A1(v12), .B0(v10), .Y(n97));
OAI21X1  g66(.A0(v9), .A1(n70), .B0(v0), .Y(n98));
NAND3X1  g67(.A(n98), .B(n97), .C(n45), .Y(n99));
OAI21X1  g68(.A0(n96), .A1(v12), .B0(n99), .Y(n39));
OAI22X1  g69(.A0(v9), .A1(v10), .B0(n32), .B1(n75), .Y(n101));
AOI22X1  g70(.A0(n71), .A1(n33), .B0(n45), .B1(n101), .Y(n102));
OR4X1    g71(.A(v11), .B(v12), .C(v5), .D(n54_1), .Y(n103));
AOI21X1  g72(.A0(n103), .A1(v10), .B0(n48), .Y(n104));
AOI21X1  g73(.A0(n71), .A1(n33), .B0(n104), .Y(n105));
OAI22X1  g74(.A0(n102), .A1(n70), .B0(v0), .B1(n105), .Y(n44));
MX2X1    g75(.A(v2), .B(v11), .S0(v7), .Y(n107));
NOR3X1   g76(.A(n107), .B(n37), .C(n58), .Y(n108));
AOI21X1  g77(.A0(n37), .A1(v2), .B0(v7), .Y(n109));
NAND2X1  g78(.A(n36), .B(v4), .Y(n110));
NAND4X1  g79(.A(n37), .B(v11), .C(v5), .D(v7), .Y(n111));
OAI21X1  g80(.A0(n110), .A1(n109), .B0(n111), .Y(n112));
OAI21X1  g81(.A0(n112), .A1(n108), .B0(n33), .Y(n113));
NOR3X1   g82(.A(v8), .B(v11), .C(n33), .Y(n114));
NOR3X1   g83(.A(n37), .B(n36), .C(v12), .Y(n115));
OAI21X1  g84(.A0(n115), .A1(n114), .B0(n34_1), .Y(n116));
AOI21X1  g85(.A0(n116), .A1(n113), .B0(n81), .Y(n49));
OAI21X1  g86(.A0(n34_1), .A1(n37), .B0(v11), .Y(n118));
AOI21X1  g87(.A0(n118), .A1(n68), .B0(n72), .Y(n54));
endmodule
