// Benchmark "b06_C" written by ABC on Wed Aug 05 14:38:19 2020

module b06_C ( 
    EQL, ACKOUT_REG_SCAN_IN, CONT_EQL, STATE_REG_2__SCAN_IN,
    STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, CC_MUX_REG_2__SCAN_IN,
    CC_MUX_REG_1__SCAN_IN, USCITE_REG_2__SCAN_IN, USCITE_REG_1__SCAN_IN,
    ENABLE_COUNT_REG_SCAN_IN,
    U57, U56, U55, U59, U58, U61, U60, U62, U62  );
  input  EQL, ACKOUT_REG_SCAN_IN, CONT_EQL, STATE_REG_2__SCAN_IN,
    STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, CC_MUX_REG_2__SCAN_IN,
    CC_MUX_REG_1__SCAN_IN, USCITE_REG_2__SCAN_IN, USCITE_REG_1__SCAN_IN,
    ENABLE_COUNT_REG_SCAN_IN;
  output U57, U56, U55, U59, U58, U61, U60, U62, U62;
  wire n26, n27, n28, n29, n30, n32, n33, n34, n35, n36, n37, n39, n40, n42,
    n44, n45, n46, n49, n51, n52;
  NOR2X1  g00(.A(STATE_REG_0__SCAN_IN), .B(STATE_REG_1__SCAN_IN), .Y(n26));
  OAI21X1 g01(.A0(n26), .A1(EQL), .B0(STATE_REG_2__SCAN_IN), .Y(n27));
  INVX1   g02(.A(STATE_REG_2__SCAN_IN), .Y(n28));
  INVX1   g03(.A(STATE_REG_1__SCAN_IN), .Y(n29));
  NAND3X1 g04(.A(STATE_REG_0__SCAN_IN), .B(n29), .C(n28), .Y(n30));
  OAI21X1 g05(.A0(n30), .A1(EQL), .B0(n27), .Y(U57));
  NAND2X1 g06(.A(STATE_REG_1__SCAN_IN), .B(EQL), .Y(n32));
  NAND3X1 g07(.A(STATE_REG_0__SCAN_IN), .B(n28), .C(EQL), .Y(n33));
  INVX1   g08(.A(EQL), .Y(n34));
  NAND3X1 g09(.A(n26), .B(STATE_REG_2__SCAN_IN), .C(n34), .Y(n35));
  INVX1   g10(.A(STATE_REG_0__SCAN_IN), .Y(n36));
  NAND3X1 g11(.A(n36), .B(STATE_REG_1__SCAN_IN), .C(n28), .Y(n37));
  NAND4X1 g12(.A(n35), .B(n33), .C(n32), .D(n37), .Y(U56));
  NOR3X1  g13(.A(STATE_REG_0__SCAN_IN), .B(STATE_REG_1__SCAN_IN), .C(STATE_REG_2__SCAN_IN), .Y(n39));
  AOI21X1 g14(.A0(STATE_REG_0__SCAN_IN), .A1(STATE_REG_1__SCAN_IN), .B0(n39), .Y(n40));
  OAI21X1 g15(.A0(n26), .A1(EQL), .B0(n40), .Y(U55));
  NAND3X1 g16(.A(n36), .B(STATE_REG_1__SCAN_IN), .C(EQL), .Y(n42));
  NAND3X1 g17(.A(n42), .B(n30), .C(n27), .Y(U59));
  NAND2X1 g18(.A(n36), .B(n28), .Y(n44));
  OAI21X1 g19(.A0(STATE_REG_0__SCAN_IN), .A1(n34), .B0(STATE_REG_1__SCAN_IN), .Y(n45));
  AOI22X1 g20(.A0(n29), .A1(EQL), .B0(STATE_REG_2__SCAN_IN), .B1(STATE_REG_0__SCAN_IN), .Y(n46));
  NAND3X1 g21(.A(n46), .B(n45), .C(n44), .Y(U58));
  OAI21X1 g22(.A0(n32), .A1(n28), .B0(n35), .Y(U61));
  AOI21X1 g23(.A0(STATE_REG_1__SCAN_IN), .A1(STATE_REG_2__SCAN_IN), .B0(n34), .Y(n49));
  NAND2X1 g24(.A(n49), .B(n40), .Y(U60));
  NOR3X1  g25(.A(n36), .B(n29), .C(n28), .Y(n51));
  NAND4X1 g26(.A(STATE_REG_1__SCAN_IN), .B(n28), .C(n34), .D(n36), .Y(n52));
  OAI21X1 g27(.A0(n51), .A1(CONT_EQL), .B0(n52), .Y(U62));
endmodule


