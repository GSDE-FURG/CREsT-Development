// Benchmark "b10_C" written by ABC on Wed Aug 05 14:39:43 2020

module b10_C ( 
    R_BUTTON, G_BUTTON, KEY, START, TEST, RTS, RTR, VOTO0_REG_SCAN_IN,
    V_IN_3_, V_IN_2_, V_IN_1_, V_IN_0_, STATO_REG_3__SCAN_IN,
    STATO_REG_2__SCAN_IN, STATO_REG_1__SCAN_IN, STATO_REG_0__SCAN_IN,
    V_OUT_REG_3__SCAN_IN, V_OUT_REG_2__SCAN_IN, V_OUT_REG_1__SCAN_IN,
    V_OUT_REG_0__SCAN_IN, SIGN_REG_3__SCAN_IN, VOTO1_REG_SCAN_IN,
    CTR_REG_SCAN_IN, VOTO3_REG_SCAN_IN, LAST_R_REG_SCAN_IN,
    CTS_REG_SCAN_IN, VOTO2_REG_SCAN_IN, LAST_G_REG_SCAN_IN,
    U212, U211, U210, U233, U234, U235, U236, U237, U209, U238, U208, U239,
    U240, U207, U241, U242, U243  );
  input  R_BUTTON, G_BUTTON, KEY, START, TEST, RTS, RTR,
    VOTO0_REG_SCAN_IN, V_IN_3_, V_IN_2_, V_IN_1_, V_IN_0_,
    STATO_REG_3__SCAN_IN, STATO_REG_2__SCAN_IN, STATO_REG_1__SCAN_IN,
    STATO_REG_0__SCAN_IN, V_OUT_REG_3__SCAN_IN, V_OUT_REG_2__SCAN_IN,
    V_OUT_REG_1__SCAN_IN, V_OUT_REG_0__SCAN_IN, SIGN_REG_3__SCAN_IN,
    VOTO1_REG_SCAN_IN, CTR_REG_SCAN_IN, VOTO3_REG_SCAN_IN,
    LAST_R_REG_SCAN_IN, CTS_REG_SCAN_IN, VOTO2_REG_SCAN_IN,
    LAST_G_REG_SCAN_IN;
  output U212, U211, U210, U233, U234, U235, U236, U237, U209, U238, U208,
    U239, U240, U207, U241, U242, U243;
  wire n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
    n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
    n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n92, n93,
    n94, n95, n96, n97, n98, n99, n101, n102, n103, n104, n106, n107, n108,
    n109, n111, n113, n115, n117, n119, n120, n122, n123, n124, n125, n126,
    n127, n128, n129, n130, n131, n132, n133, n134, n136, n140, n142, n143,
    n144, n145, n146, n147, n148, n149, n151, n152, n153, n154, n156, n157,
    n158, n159, n160, n161, n163, n164, n165, n166, n167, n168, n170, n172,
    n173, n174, n175, n176, n177, n178;
  INVX1   g000(.A(STATO_REG_3__SCAN_IN), .Y(n51));
  NOR2X1  g001(.A(STATO_REG_1__SCAN_IN), .B(RTR), .Y(n52));
  INVX1   g002(.A(STATO_REG_1__SCAN_IN), .Y(n53));
  INVX1   g003(.A(STATO_REG_0__SCAN_IN), .Y(n54));
  OAI21X1 g004(.A0(n53), .A1(STATO_REG_2__SCAN_IN), .B0(n54), .Y(n55));
  NAND4X1 g005(.A(V_IN_1_), .B(V_IN_2_), .C(V_IN_3_), .D(V_IN_0_), .Y(n56));
  AOI21X1 g006(.A0(n56), .A1(STATO_REG_0__SCAN_IN), .B0(n51), .Y(n57));
  OAI21X1 g007(.A0(n55), .A1(n52), .B0(n57), .Y(n58));
  INVX1   g008(.A(RTS), .Y(n59));
  NOR2X1  g009(.A(STATO_REG_2__SCAN_IN), .B(STATO_REG_3__SCAN_IN), .Y(n60));
  NAND2X1 g010(.A(n60), .B(n54), .Y(n61));
  NAND3X1 g011(.A(n54), .B(STATO_REG_1__SCAN_IN), .C(STATO_REG_2__SCAN_IN), .Y(n62));
  OAI22X1 g012(.A0(n61), .A1(STATO_REG_1__SCAN_IN), .B0(n59), .B1(n62), .Y(n63));
  INVX1   g013(.A(START), .Y(n64));
  NOR4X1  g014(.A(STATO_REG_2__SCAN_IN), .B(STATO_REG_3__SCAN_IN), .C(n64), .D(n54), .Y(n65));
  INVX1   g015(.A(RTR), .Y(n66));
  NAND4X1 g016(.A(STATO_REG_1__SCAN_IN), .B(STATO_REG_2__SCAN_IN), .C(n66), .D(STATO_REG_0__SCAN_IN), .Y(n67));
  NAND4X1 g017(.A(n53), .B(STATO_REG_2__SCAN_IN), .C(n59), .D(STATO_REG_0__SCAN_IN), .Y(n68));
  INVX1   g018(.A(STATO_REG_2__SCAN_IN), .Y(n69));
  NAND4X1 g019(.A(n69), .B(n51), .C(n64), .D(STATO_REG_1__SCAN_IN), .Y(n70));
  NAND4X1 g020(.A(n53), .B(STATO_REG_2__SCAN_IN), .C(RTR), .D(n54), .Y(n71));
  NAND4X1 g021(.A(n70), .B(n68), .C(n67), .D(n71), .Y(n72));
  NOR3X1  g022(.A(n72), .B(n65), .C(n63), .Y(n73));
  AOI21X1 g023(.A0(n73), .A1(n58), .B0(STATO_REG_0__SCAN_IN), .Y(n74));
  NOR3X1  g024(.A(STATO_REG_0__SCAN_IN), .B(STATO_REG_2__SCAN_IN), .C(STATO_REG_3__SCAN_IN), .Y(n75));
  NOR3X1  g025(.A(STATO_REG_0__SCAN_IN), .B(n53), .C(n69), .Y(n76));
  AOI22X1 g026(.A0(n75), .A1(n53), .B0(RTS), .B1(n76), .Y(n77));
  NAND3X1 g027(.A(n60), .B(STATO_REG_0__SCAN_IN), .C(START), .Y(n78));
  NOR4X1  g028(.A(n53), .B(n69), .C(RTR), .D(n54), .Y(n79));
  NOR4X1  g029(.A(STATO_REG_1__SCAN_IN), .B(n69), .C(RTS), .D(n54), .Y(n80));
  NOR4X1  g030(.A(STATO_REG_2__SCAN_IN), .B(STATO_REG_3__SCAN_IN), .C(START), .D(n53), .Y(n81));
  NOR4X1  g031(.A(STATO_REG_1__SCAN_IN), .B(n69), .C(n66), .D(STATO_REG_0__SCAN_IN), .Y(n82));
  NOR4X1  g032(.A(n81), .B(n80), .C(n79), .D(n82), .Y(n83));
  NAND4X1 g033(.A(n78), .B(n77), .C(n58), .D(n83), .Y(n84));
  NAND2X1 g034(.A(n54), .B(STATO_REG_2__SCAN_IN), .Y(n85));
  INVX1   g035(.A(VOTO0_REG_SCAN_IN), .Y(n86));
  INVX1   g036(.A(VOTO3_REG_SCAN_IN), .Y(n87));
  NAND4X1 g037(.A(n87), .B(VOTO1_REG_SCAN_IN), .C(n86), .D(VOTO2_REG_SCAN_IN), .Y(n88));
  OAI22X1 g038(.A0(n85), .A1(n88), .B0(n61), .B1(TEST), .Y(n89));
  NAND3X1 g039(.A(n89), .B(n84), .C(n53), .Y(n90));
  OAI21X1 g040(.A0(n74), .A1(n51), .B0(n90), .Y(U212));
  NAND2X1 g041(.A(STATO_REG_0__SCAN_IN), .B(n53), .Y(n92));
  INVX1   g042(.A(VOTO1_REG_SCAN_IN), .Y(n93));
  INVX1   g043(.A(VOTO2_REG_SCAN_IN), .Y(n94));
  NOR4X1  g044(.A(VOTO3_REG_SCAN_IN), .B(n93), .C(VOTO0_REG_SCAN_IN), .D(n94), .Y(n95));
  OAI21X1 g045(.A0(n95), .A1(STATO_REG_0__SCAN_IN), .B0(n92), .Y(n96));
  AOI21X1 g046(.A0(n73), .A1(n58), .B0(n96), .Y(n97));
  XOR2X1  g047(.A(STATO_REG_0__SCAN_IN), .B(STATO_REG_3__SCAN_IN), .Y(n98));
  AOI21X1 g048(.A0(n98), .A1(STATO_REG_1__SCAN_IN), .B0(n76), .Y(n99));
  OAI21X1 g049(.A0(n97), .A1(n69), .B0(n99), .Y(U211));
  AOI21X1 g050(.A0(STATO_REG_1__SCAN_IN), .A1(n51), .B0(n54), .Y(n101));
  NAND3X1 g051(.A(n54), .B(STATO_REG_1__SCAN_IN), .C(n51), .Y(n102));
  NAND2X1 g052(.A(n102), .B(n62), .Y(n103));
  AOI21X1 g053(.A0(n101), .A1(n84), .B0(n103), .Y(n104));
  OAI21X1 g054(.A0(n84), .A1(n53), .B0(n104), .Y(U210));
  NOR2X1  g055(.A(STATO_REG_0__SCAN_IN), .B(STATO_REG_1__SCAN_IN), .Y(n106));
  OAI21X1 g056(.A0(n88), .A1(STATO_REG_3__SCAN_IN), .B0(n106), .Y(n107));
  NAND3X1 g057(.A(n107), .B(n62), .C(n61), .Y(n108));
  NAND2X1 g058(.A(n108), .B(n84), .Y(n109));
  OAI21X1 g059(.A0(n84), .A1(n54), .B0(n109), .Y(U233));
  NAND2X1 g060(.A(n71), .B(V_OUT_REG_3__SCAN_IN), .Y(n111));
  OAI21X1 g061(.A0(n71), .A1(n87), .B0(n111), .Y(U234));
  NAND2X1 g062(.A(n71), .B(V_OUT_REG_2__SCAN_IN), .Y(n113));
  OAI21X1 g063(.A0(n71), .A1(n94), .B0(n113), .Y(U235));
  NAND2X1 g064(.A(n71), .B(V_OUT_REG_1__SCAN_IN), .Y(n115));
  OAI21X1 g065(.A0(n71), .A1(n93), .B0(n115), .Y(U236));
  NAND2X1 g066(.A(n71), .B(V_OUT_REG_0__SCAN_IN), .Y(n117));
  OAI21X1 g067(.A0(n71), .A1(n86), .B0(n117), .Y(U237));
  INVX1   g068(.A(SIGN_REG_3__SCAN_IN), .Y(n119));
  NOR3X1  g069(.A(n61), .B(STATO_REG_1__SCAN_IN), .C(TEST), .Y(n120));
  OAI22X1 g070(.A0(n119), .A1(n120), .B0(n54), .B1(n51), .Y(U209));
  NAND4X1 g071(.A(n53), .B(n69), .C(STATO_REG_3__SCAN_IN), .D(STATO_REG_0__SCAN_IN), .Y(n122));
  OAI21X1 g072(.A0(n62), .A1(STATO_REG_3__SCAN_IN), .B0(n122), .Y(n123));
  INVX1   g073(.A(KEY), .Y(n124));
  NOR4X1  g074(.A(n53), .B(STATO_REG_2__SCAN_IN), .C(n124), .D(VOTO1_REG_SCAN_IN), .Y(n125));
  AOI21X1 g075(.A0(n123), .A1(V_IN_1_), .B0(n125), .Y(n126));
  NOR4X1  g076(.A(STATO_REG_1__SCAN_IN), .B(STATO_REG_2__SCAN_IN), .C(n51), .D(n54), .Y(n127));
  NOR4X1  g077(.A(STATO_REG_1__SCAN_IN), .B(STATO_REG_2__SCAN_IN), .C(n64), .D(n54), .Y(n128));
  INVX1   g078(.A(LAST_G_REG_SCAN_IN), .Y(n129));
  NAND4X1 g079(.A(n129), .B(START), .C(G_BUTTON), .D(n75), .Y(n130));
  NAND3X1 g080(.A(n75), .B(START), .C(n124), .Y(n131));
  NAND2X1 g081(.A(n131), .B(n130), .Y(n132));
  NOR4X1  g082(.A(n128), .B(n127), .C(n63), .D(n132), .Y(n133));
  NAND2X1 g083(.A(n133), .B(VOTO1_REG_SCAN_IN), .Y(n134));
  OAI21X1 g084(.A0(n133), .A1(n126), .B0(n134), .Y(U238));
  XOR2X1  g085(.A(STATO_REG_1__SCAN_IN), .B(n69), .Y(n136));
  NAND2X1 g086(.A(n77), .B(CTR_REG_SCAN_IN), .Y(n140));
  NAND2X1 g087(.A(n140), .B(n68), .Y(U208));
  XOR2X1  g088(.A(VOTO2_REG_SCAN_IN), .B(VOTO0_REG_SCAN_IN), .Y(n142));
  XOR2X1  g089(.A(n142), .B(n93), .Y(n143));
  NOR3X1  g090(.A(n143), .B(n54), .C(n53), .Y(n144));
  AOI21X1 g091(.A0(n123), .A1(V_IN_3_), .B0(n144), .Y(n145));
  AOI22X1 g092(.A0(STATO_REG_1__SCAN_IN), .A1(STATO_REG_0__SCAN_IN), .B0(START), .B1(n124), .Y(n146));
  NOR3X1  g093(.A(n146), .B(STATO_REG_2__SCAN_IN), .C(STATO_REG_3__SCAN_IN), .Y(n147));
  NOR4X1  g094(.A(n128), .B(n127), .C(n63), .D(n147), .Y(n148));
  NAND2X1 g095(.A(n148), .B(VOTO3_REG_SCAN_IN), .Y(n149));
  OAI21X1 g096(.A0(n148), .A1(n145), .B0(n149), .Y(U239));
  INVX1   g097(.A(LAST_R_REG_SCAN_IN), .Y(n151));
  NOR4X1  g098(.A(n53), .B(n64), .C(n124), .D(n61), .Y(n152));
  NOR4X1  g099(.A(STATO_REG_2__SCAN_IN), .B(STATO_REG_3__SCAN_IN), .C(n64), .D(STATO_REG_0__SCAN_IN), .Y(n153));
  NAND4X1 g100(.A(STATO_REG_1__SCAN_IN), .B(KEY), .C(R_BUTTON), .D(n153), .Y(n154));
  OAI21X1 g101(.A0(n152), .A1(n151), .B0(n154), .Y(U240));
  OAI21X1 g102(.A0(STATO_REG_0__SCAN_IN), .A1(STATO_REG_3__SCAN_IN), .B0(RTR), .Y(n156));
  OAI21X1 g103(.A0(STATO_REG_0__SCAN_IN), .A1(n53), .B0(n156), .Y(n157));
  OAI21X1 g104(.A0(n92), .A1(n51), .B0(n136), .Y(n158));
  OAI21X1 g105(.A0(n158), .A1(n157), .B0(CTS_REG_SCAN_IN), .Y(n159));
  NAND4X1 g106(.A(STATO_REG_0__SCAN_IN), .B(n53), .C(RTR), .D(n60), .Y(n160));
  NAND4X1 g107(.A(n53), .B(STATO_REG_2__SCAN_IN), .C(STATO_REG_3__SCAN_IN), .D(n54), .Y(n161));
  NAND4X1 g108(.A(n160), .B(n159), .C(n71), .D(n161), .Y(U207));
  NOR4X1  g109(.A(n53), .B(STATO_REG_2__SCAN_IN), .C(n124), .D(VOTO2_REG_SCAN_IN), .Y(n163));
  AOI21X1 g110(.A0(n123), .A1(V_IN_2_), .B0(n163), .Y(n164));
  NAND4X1 g111(.A(n151), .B(START), .C(R_BUTTON), .D(n75), .Y(n165));
  NAND2X1 g112(.A(n165), .B(n131), .Y(n166));
  NOR4X1  g113(.A(n128), .B(n127), .C(n63), .D(n166), .Y(n167));
  NAND2X1 g114(.A(n167), .B(VOTO2_REG_SCAN_IN), .Y(n168));
  OAI21X1 g115(.A0(n167), .A1(n164), .B0(n168), .Y(U241));
  NAND4X1 g116(.A(STATO_REG_1__SCAN_IN), .B(KEY), .C(G_BUTTON), .D(n153), .Y(n170));
  OAI21X1 g117(.A0(n152), .A1(n129), .B0(n170), .Y(U242));
  OAI22X1 g118(.A0(SIGN_REG_3__SCAN_IN), .A1(n51), .B0(n124), .B1(n61), .Y(n172));
  AOI22X1 g119(.A0(n123), .A1(V_IN_0_), .B0(STATO_REG_1__SCAN_IN), .B1(n172), .Y(n173));
  NAND2X1 g120(.A(n60), .B(START), .Y(n174));
  NAND3X1 g121(.A(n98), .B(STATO_REG_1__SCAN_IN), .C(n69), .Y(n175));
  NAND2X1 g122(.A(n175), .B(n174), .Y(n176));
  NOR3X1  g123(.A(n176), .B(n127), .C(n63), .Y(n177));
  NAND2X1 g124(.A(n177), .B(VOTO0_REG_SCAN_IN), .Y(n178));
  OAI21X1 g125(.A0(n177), .A1(n173), .B0(n178), .Y(U243));
endmodule


