//Converted to Combinational (Partial output: g31793) , Module name: s38584_g31793 , Timestamp: 2018-12-03T15:51:18.280857 
module s38584_g31793 ( g35, g5471, g5817, g5124, g6163, g3817, g3115, g6509, g3466, g4427, g4420, g31793 );
input g35, g5471, g5817, g5124, g6163, g3817, g3115, g6509, g3466, g4427, g4420;
output g31793;
wire n4777, n4763, n4768, n4772, n4773, n4774, n4776, n4762, n4745, n4751_1, n4758, n4740, n4764, n4767, n4769, n4771, n4746_1, n4737, n4738, n4739, n4753, n4620, n4756_1, n4752, n4775_1, n4736_1, n4748, n4749, n4759, n4761_1, n4744, n4750, n4747, n4757, n4755, n4760, n4765, n4766_1, n4741_1, n4770_1, n4743, n4742, n4754;
NAND4X1  g0158(.A(n4772), .B(n4768), .C(n4763), .D(n4777), .Y(g31793));
OAI21X1  g0157(.A0(n4776), .A1(n4774), .B0(n4773), .Y(n4777));
NOR4X1   g0143(.A(n4758), .B(n4751_1), .C(n4745), .D(n4762), .Y(n4763));
OAI21X1  g0148(.A0(n4767), .A1(n4764), .B0(n4740), .Y(n4768));
OAI21X1  g0152(.A0(n4771), .A1(n4769), .B0(n4740), .Y(n4772));
NOR4X1   g0153(.A(n4739), .B(n4738), .C(n4737), .D(n4746_1), .Y(n4773));
NOR4X1   g0154(.A(n4752), .B(n4756_1), .C(n4620), .D(n4753), .Y(n4774));
NOR4X1   g0156(.A(n4749), .B(n4748), .C(n4736_1), .D(n4775_1), .Y(n4776));
NOR2X1   g0142(.A(n4761_1), .B(n4759), .Y(n4762));
INVX1    g0125(.A(n4744), .Y(n4745));
NOR4X1   g0131(.A(n4747), .B(n4746_1), .C(n4739), .D(n4750), .Y(n4751_1));
NOR4X1   g0138(.A(n4755), .B(n4753), .C(n4752), .D(n4757), .Y(n4758));
NOR4X1   g0120(.A(n4738), .B(n4737), .C(n4736_1), .D(n4739), .Y(n4740));
NOR4X1   g0144(.A(n4748), .B(n4752), .C(n4746_1), .D(n4760), .Y(n4764));
NOR4X1   g0147(.A(n4766_1), .B(n4765), .C(n4746_1), .D(n4753), .Y(n4767));
NOR3X1   g0149(.A(n4753), .B(n4752), .C(n4741_1), .Y(n4769));
NOR4X1   g0151(.A(n4770_1), .B(n4752), .C(n4746_1), .D(n4749), .Y(n4771));
INVX1    g0126(.A(n4741_1), .Y(n4746_1));
AND2X1   g0117(.A(g5471), .B(g35), .Y(n4737));
AND2X1   g0118(.A(g5817), .B(g35), .Y(n4738));
AND2X1   g0119(.A(g5124), .B(g35), .Y(n4739));
INVX1    g0133(.A(n4743), .Y(n4753));
INVX1    g0000(.A(g35), .Y(n4620));
INVX1    g0136(.A(g6163), .Y(n4756_1));
INVX1    g0132(.A(n4742), .Y(n4752));
NAND2X1  g0155(.A(n4766_1), .B(n4765), .Y(n4775_1));
AND2X1   g0116(.A(g6163), .B(g35), .Y(n4736_1));
AND2X1   g0128(.A(g3817), .B(g35), .Y(n4748));
AND2X1   g0129(.A(g3115), .B(g35), .Y(n4749));
OR4X1    g0139(.A(n4738), .B(n4737), .C(n4736_1), .D(n4748), .Y(n4759));
NAND4X1  g0141(.A(n4742), .B(n4741_1), .C(n4739), .D(n4760), .Y(n4761_1));
NAND4X1  g0124(.A(n4742), .B(n4741_1), .C(n4740), .D(n4743), .Y(n4744));
OR4X1    g0130(.A(n4748), .B(n4738), .C(n4736_1), .D(n4749), .Y(n4750));
NAND2X1  g0127(.A(n4742), .B(n4737), .Y(n4747));
NAND3X1  g0137(.A(n4756_1), .B(g5817), .C(g35), .Y(n4757));
OR2X1    g0135(.A(n4754), .B(n4737), .Y(n4755));
INVX1    g0140(.A(n4749), .Y(n4760));
AND2X1   g0145(.A(g6509), .B(g35), .Y(n4765));
NAND2X1  g0146(.A(g3466), .B(g35), .Y(n4766_1));
OAI21X1  g0121(.A0(g4420), .A1(g4427), .B0(g35), .Y(n4741_1));
INVX1    g0150(.A(n4748), .Y(n4770_1));
OAI21X1  g0123(.A0(g3115), .A1(g3817), .B0(g35), .Y(n4743));
OAI21X1  g0122(.A0(g6509), .A1(g3466), .B0(g35), .Y(n4742));
OR2X1    g0134(.A(n4746_1), .B(n4739), .Y(n4754));

endmodule
