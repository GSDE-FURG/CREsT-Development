//Converted to Combinational (Partial output: n65) , Module name: s1494_n65 , Timestamp: 2018-12-03T15:51:02.656860 
module s1494_n65 ( v1, CLR, v7, v11, v12, v10, v8, v9, v6, v3, v5, v4, v2, v0, n65 );
input v1, CLR, v7, v11, v12, v10, v8, v9, v6, v3, v5, v4, v2, v0;
output n65;
wire n267, n334, n339, n68, n324, n333, n338, n94, n336, n93, n320, n323, n332, n327, n337, n70_1, n335, n191, n318, n319, n322, n45, n321, n331, n192, n328, n330, n326, n119, n116, n325, n190, n107, n293, n104, n67, n100, n96, n62, n329, n140, n178, n47, n86, n83, n103, n84;
AOI21X1  g294(.A0(n339), .A1(n334), .B0(n267), .Y(n65));
INVX1    g221(.A(CLR), .Y(n267));
OAI21X1  g288(.A0(n333), .A1(n324), .B0(n68), .Y(n334));
AOI21X1  g293(.A0(n336), .A1(n94), .B0(n338), .Y(n339));
INVX1    g023(.A(v7), .Y(n68));
AOI21X1  g278(.A0(n323), .A1(n320), .B0(n93), .Y(n324));
OAI21X1  g287(.A0(n327), .A1(v11), .B0(n332), .Y(n333));
NOR4X1   g292(.A(n68), .B(n70_1), .C(v12), .D(n337), .Y(n338));
NOR2X1   g049(.A(n93), .B(v11), .Y(n94));
OAI21X1  g290(.A0(n191), .A1(v10), .B0(n335), .Y(n336));
INVX1    g048(.A(v8), .Y(n93));
OAI21X1  g274(.A0(n319), .A1(n318), .B0(v9), .Y(n320));
AOI22X1  g277(.A0(n321), .A1(n45), .B0(n70_1), .B1(n322), .Y(n323));
AOI22X1  g286(.A0(n330), .A1(n328), .B0(n192), .B1(n331), .Y(n332));
AOI22X1  g281(.A0(n325), .A1(n116), .B0(n119), .B1(n326), .Y(n327));
AOI21X1  g291(.A0(v8), .A1(n45), .B0(v11), .Y(n337));
INVX1    g025(.A(v9), .Y(n70_1));
NAND3X1  g289(.A(n70_1), .B(v10), .C(v12), .Y(n335));
INVX1    g145(.A(n190), .Y(n191));
NOR3X1   g272(.A(n293), .B(n107), .C(n119), .Y(n318));
NOR3X1   g273(.A(v11), .B(v12), .C(v6), .Y(n319));
OAI21X1  g276(.A0(n192), .A1(v11), .B0(n104), .Y(n322));
INVX1    g000(.A(v10), .Y(n45));
MX2X1    g275(.A(v11), .B(n100), .S0(n67), .Y(n321));
MX2X1    g285(.A(v8), .B(n96), .S0(v10), .Y(n331));
NOR2X1   g146(.A(v12), .B(n62), .Y(n192));
NOR2X1   g282(.A(v8), .B(n67), .Y(n328));
OAI22X1  g284(.A0(n140), .A1(v9), .B0(v10), .B1(n329), .Y(n330));
MX2X1    g280(.A(n47), .B(n178), .S0(v12), .Y(n326));
INVX1    g073(.A(v3), .Y(n119));
NOR2X1   g071(.A(v9), .B(v10), .Y(n116));
NOR2X1   g279(.A(n100), .B(v12), .Y(n325));
NAND2X1  g144(.A(n70_1), .B(v12), .Y(n190));
NAND2X1  g062(.A(v11), .B(v12), .Y(n107));
NOR3X1   g247(.A(n83), .B(v1), .C(n86), .Y(n293));
INVX1    g059(.A(n103), .Y(n104));
INVX1    g022(.A(v12), .Y(n67));
NAND2X1  g055(.A(v4), .B(v5), .Y(n100));
NOR2X1   g051(.A(v8), .B(n70_1), .Y(n96));
INVX1    g017(.A(v2), .Y(n62));
AOI21X1  g283(.A0(n84), .A1(v6), .B0(v9), .Y(n329));
NAND2X1  g094(.A(v10), .B(v11), .Y(n140));
NOR2X1   g132(.A(v8), .B(v10), .Y(n178));
AND2X1   g002(.A(v8), .B(v9), .Y(n47));
INVX1    g041(.A(v6), .Y(n86));
INVX1    g038(.A(v0), .Y(n83));
NOR2X1   g058(.A(v10), .B(v12), .Y(n103));
INVX1    g039(.A(v11), .Y(n84));

endmodule
