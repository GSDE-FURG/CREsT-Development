//Converted to Combinational (Partial output: n2982) , Module name: s38417_n2982 , Timestamp: 2018-12-03T15:51:12.739128 
module s38417_n2982 ( g823, g876, g785, g826, g873, g879, g853, g869, g999, g1001, g1000, g1090, g1089, g1091, g1005, g1007, g1006, g857, g856, g858, g1002, g1004, g1003, g963, g1088, g1092, g909, g915, g912, g882, g888, g885, g918, g924, g921, g897, g894, g900, g906, g903, g891, g945, g951, g948, g936, g942, g939, g954, g960, g957, g927, g933, g930, g809, g801, g797, g805, g813, g845, g844, g846, g793, g789, g1009, g1008, g1010, g842, g841, g843, g860, g859, g861, g851, g850, g852, g863, g862, g864, g848, g847, g849, g836, g835, g837, g833, g832, g834, g839, g838, g840, g818, g817, g819, g830, g829, g831, g821, g820, g822, n2982 );
input g823, g876, g785, g826, g873, g879, g853, g869, g999, g1001, g1000, g1090, g1089, g1091, g1005, g1007, g1006, g857, g856, g858, g1002, g1004, g1003, g963, g1088, g1092, g909, g915, g912, g882, g888, g885, g918, g924, g921, g897, g894, g900, g906, g903, g891, g945, g951, g948, g936, g942, g939, g954, g960, g957, g927, g933, g930, g809, g801, g797, g805, g813, g845, g844, g846, g793, g789, g1009, g1008, g1010, g842, g841, g843, g860, g859, g861, g851, g850, g852, g863, g862, g864, g848, g847, g849, g836, g835, g837, g833, g832, g834, g839, g838, g840, g818, g817, g819, g830, g829, g831, g821, g820, g822;
output n2982;
wire n6611, n6606, n6610_1, n6608, n6605_1, n3496, n6609, n6604, n6501, n6607, n6577, n6580, n6587_1, n6590, n6592_1, n6603, n6600_1, n6499_1, n6500, n6483, n6558, n6576, n6579_1, n6586, n6570, n6583_1, n6589, n6564_1, n6591, n6602, n6596_1, n6601, n6594, n6599, n6451, n6468, n6482, n6442, n6520, n6557, n6575, n6567, n6571, n6578, n6585, n6568, n6569_1, n6581, n6582, n6588, n6560, n6563, n6492, n6505, n6538, n6595, n6533, n6546, n6529_1, n6542, n6593, n6598, n6450, n6439_1, n6446, n6467, n6455, n6459_1, n6463, n6481, n6469_1, n6473, n6477, n6440, n6441, n6512, n6515, n6519_1, n6549_1, n6552, n6556, n6574_1, n6565, n6566, n6584, n6559_1, n6562, n6561, n6484_1, n6485, n6503, n6504_1, n6536, n6537, n6508, n6494_1, n6495, n6507, n6531, n6532, n6544_1, n6545, n6521, n6522, n6540, n6541, n6597, n3442, n6449_1, n6412, n6438, n6406, n6445, n6466, n3460, n6454_1, n3469, n6458, n3451, n6462, n6480, n3433, n6464_1, n6465, n3478, n6472, n3487, n6476, n6401, n6404_1, n6403, n6498, n6511, n6513, n6514_1, n6516, n6517, n6518, n6535, n6548, n6550, n6551, n6553, n6554_1, n6555, n6572, n6573, n6447, n6448, n6410, n6411, n6436, n6437, n6402, n6405, n6443, n6444_1, n6452, n6453, n6456, n6457, n6460, n6461, n6478, n6479_1, n6470, n6471, n6474_1, n6475, n6487, n6493, n6497, n6502, n6506, n6510, n6509_1, n6524_1, n6530, n6534_1, n6539_1, n6543, n6547, n6486, n6488, n6491, n6496, n6523, n6525, n6528, n6490, n6489_1, n6527, n6526;
MX2X1    g1570(.A(g876), .B(n6611), .S0(g823), .Y(n2982));
MX2X1    g1568(.A(n6608), .B(n6610_1), .S0(n6606), .Y(n6611));
INVX1    g1563(.A(n6605_1), .Y(n6606));
AOI21X1  g1567(.A0(n6604), .A1(n6609), .B0(n3496), .Y(n6610_1));
XOR2X1   g1565(.A(n6607), .B(n6501), .Y(n6608));
NOR4X1   g1562(.A(n6587_1), .B(n6580), .C(n6577), .D(n6604), .Y(n6605_1));
INVX1    g1323(.A(g785), .Y(n3496));
NOR3X1   g1566(.A(n6587_1), .B(n6580), .C(n6577), .Y(n6609));
AOI22X1  g1561(.A0(n6600_1), .A1(n6603), .B0(n6592_1), .B1(n6590), .Y(n6604));
NAND2X1  g1458(.A(n6500), .B(n6499_1), .Y(n6501));
NAND2X1  g1564(.A(n6592_1), .B(n6590), .Y(n6607));
NOR3X1   g1534(.A(n6576), .B(n6558), .C(n6483), .Y(n6577));
NOR2X1   g1537(.A(n6579_1), .B(n6483), .Y(n6580));
OAI22X1  g1544(.A0(n6583_1), .A1(n6483), .B0(n6570), .B1(n6586), .Y(n6587_1));
INVX1    g1547(.A(n6589), .Y(n6590));
NAND3X1  g1549(.A(n6570), .B(n6591), .C(n6564_1), .Y(n6592_1));
OR4X1    g1560(.A(n6601), .B(n6596_1), .C(n6592_1), .D(n6602), .Y(n6603));
OR2X1    g1557(.A(n6599), .B(n6594), .Y(n6600_1));
NAND2X1  g1456(.A(g873), .B(g826), .Y(n6499_1));
AOI22X1  g1457(.A0(g876), .A1(g823), .B0(g853), .B1(g879), .Y(n6500));
NAND3X1  g1440(.A(n6482), .B(n6468), .C(n6451), .Y(n6483));
AOI21X1  g1515(.A0(n6557), .A1(n6520), .B0(n6442), .Y(n6558));
NAND4X1  g1533(.A(n6571), .B(n6567), .C(n6564_1), .D(n6575), .Y(n6576));
NAND2X1  g1536(.A(n6578), .B(n6575), .Y(n6579_1));
INVX1    g1543(.A(n6585), .Y(n6586));
NOR2X1   g1527(.A(n6569_1), .B(n6568), .Y(n6570));
NOR2X1   g1540(.A(n6582), .B(n6581), .Y(n6583_1));
NOR3X1   g1546(.A(n6569_1), .B(n6568), .C(n6588), .Y(n6589));
NOR2X1   g1521(.A(n6563), .B(n6560), .Y(n6564_1));
INVX1    g1548(.A(n6567), .Y(n6591));
NAND3X1  g1559(.A(n6538), .B(n6505), .C(n6492), .Y(n6602));
OR4X1    g1553(.A(n6546), .B(n6533), .C(n6501), .D(n6595), .Y(n6596_1));
NAND2X1  g1558(.A(n6542), .B(n6529_1), .Y(n6601));
NOR3X1   g1551(.A(n6571), .B(n6567), .C(n6593), .Y(n6594));
OR2X1    g1556(.A(n6598), .B(n6596_1), .Y(n6599));
NOR4X1   g1408(.A(n6446), .B(n6442), .C(n6439_1), .D(n6450), .Y(n6451));
NOR4X1   g1425(.A(n6463), .B(n6459_1), .C(n6455), .D(n6467), .Y(n6468));
NOR4X1   g1439(.A(n6477), .B(n6473), .C(n6469_1), .D(n6481), .Y(n6482));
OAI21X1  g1399(.A0(n6441), .A1(n6440), .B0(g869), .Y(n6442));
NOR3X1   g1477(.A(n6519_1), .B(n6515), .C(n6512), .Y(n6520));
NOR3X1   g1514(.A(n6556), .B(n6552), .C(n6549_1), .Y(n6557));
INVX1    g1532(.A(n6574_1), .Y(n6575));
NOR2X1   g1524(.A(n6566), .B(n6565), .Y(n6567));
INVX1    g1528(.A(n6570), .Y(n6571));
NOR4X1   g1535(.A(n6566), .B(n6565), .C(n6564_1), .D(n6570), .Y(n6578));
NOR3X1   g1542(.A(n6441), .B(n6440), .C(n6584), .Y(n6585));
NOR2X1   g1525(.A(g999), .B(n6559_1), .Y(n6568));
OAI22X1  g1526(.A0(g1000), .A1(n6561), .B0(n6562), .B1(g1001), .Y(n6569_1));
NOR2X1   g1538(.A(g1090), .B(n6559_1), .Y(n6581));
OAI22X1  g1539(.A0(g1091), .A1(n6561), .B0(n6562), .B1(g1089), .Y(n6582));
OR4X1    g1545(.A(n6565), .B(n6563), .C(n6560), .D(n6566), .Y(n6588));
NOR2X1   g1517(.A(g1005), .B(n6559_1), .Y(n6560));
OAI22X1  g1520(.A0(g1006), .A1(n6561), .B0(n6562), .B1(g1007), .Y(n6563));
NAND2X1  g1449(.A(n6485), .B(n6484_1), .Y(n6492));
NAND2X1  g1462(.A(n6504_1), .B(n6503), .Y(n6505));
NAND2X1  g1495(.A(n6537), .B(n6536), .Y(n6538));
NAND4X1  g1552(.A(n6507), .B(n6495), .C(n6494_1), .D(n6508), .Y(n6595));
NAND2X1  g1490(.A(n6532), .B(n6531), .Y(n6533));
NAND2X1  g1503(.A(n6545), .B(n6544_1), .Y(n6546));
NAND2X1  g1486(.A(n6522), .B(n6521), .Y(n6529_1));
NAND2X1  g1499(.A(n6541), .B(n6540), .Y(n6542));
INVX1    g1550(.A(n6564_1), .Y(n6593));
OR4X1    g1555(.A(n6542), .B(n6538), .C(n6529_1), .D(n6597), .Y(n6598));
XOR2X1   g1407(.A(n6449_1), .B(n3442), .Y(n6450));
AND2X1   g1396(.A(n6438), .B(n6412), .Y(n6439_1));
XOR2X1   g1403(.A(n6445), .B(n6406), .Y(n6446));
OAI21X1  g1424(.A0(n6438), .A1(n6412), .B0(n6466), .Y(n6467));
XOR2X1   g1412(.A(n6454_1), .B(n3460), .Y(n6455));
XOR2X1   g1416(.A(n6458), .B(n3469), .Y(n6459_1));
XOR2X1   g1420(.A(n6462), .B(n3451), .Y(n6463));
XOR2X1   g1438(.A(n6480), .B(n3496), .Y(n6481));
NOR3X1   g1426(.A(n6465), .B(n6464_1), .C(n3433), .Y(n6469_1));
XOR2X1   g1430(.A(n6472), .B(n3478), .Y(n6473));
XOR2X1   g1434(.A(n6476), .B(n3487), .Y(n6477));
NOR2X1   g1397(.A(g857), .B(n6401), .Y(n6440));
OAI22X1  g1398(.A0(g858), .A1(n6403), .B0(n6404_1), .B1(g856), .Y(n6441));
NOR2X1   g1469(.A(n6511), .B(n6498), .Y(n6512));
NOR2X1   g1472(.A(n6514_1), .B(n6513), .Y(n6515));
NOR3X1   g1476(.A(n6518), .B(n6517), .C(n6516), .Y(n6519_1));
NOR2X1   g1506(.A(n6548), .B(n6535), .Y(n6549_1));
NOR2X1   g1509(.A(n6551), .B(n6550), .Y(n6552));
NOR3X1   g1513(.A(n6555), .B(n6554_1), .C(n6553), .Y(n6556));
NOR2X1   g1531(.A(n6573), .B(n6572), .Y(n6574_1));
NOR2X1   g1522(.A(g1002), .B(n6559_1), .Y(n6565));
OAI22X1  g1523(.A0(g1003), .A1(n6561), .B0(n6562), .B1(g1004), .Y(n6566));
INVX1    g1541(.A(g869), .Y(n6584));
INVX1    g1516(.A(g963), .Y(n6559_1));
INVX1    g1519(.A(g1088), .Y(n6562));
INVX1    g1518(.A(g1092), .Y(n6561));
NAND2X1  g1441(.A(g909), .B(g826), .Y(n6484_1));
AOI22X1  g1442(.A0(g912), .A1(g823), .B0(g853), .B1(g915), .Y(n6485));
NAND2X1  g1460(.A(g882), .B(g826), .Y(n6503));
AOI22X1  g1461(.A0(g885), .A1(g823), .B0(g853), .B1(g888), .Y(n6504_1));
NAND2X1  g1493(.A(g918), .B(g826), .Y(n6536));
AOI22X1  g1494(.A0(g921), .A1(g823), .B0(g853), .B1(g924), .Y(n6537));
AOI22X1  g1465(.A0(g894), .A1(g823), .B0(g853), .B1(g897), .Y(n6508));
NAND2X1  g1451(.A(g900), .B(g826), .Y(n6494_1));
AOI22X1  g1452(.A0(g903), .A1(g823), .B0(g853), .B1(g906), .Y(n6495));
NAND2X1  g1464(.A(g891), .B(g826), .Y(n6507));
NAND2X1  g1488(.A(g945), .B(g826), .Y(n6531));
AOI22X1  g1489(.A0(g948), .A1(g823), .B0(g853), .B1(g951), .Y(n6532));
NAND2X1  g1501(.A(g936), .B(g826), .Y(n6544_1));
AOI22X1  g1502(.A0(g939), .A1(g823), .B0(g853), .B1(g942), .Y(n6545));
NAND2X1  g1478(.A(g954), .B(g826), .Y(n6521));
AOI22X1  g1479(.A0(g957), .A1(g823), .B0(g853), .B1(g960), .Y(n6522));
NAND2X1  g1497(.A(g927), .B(g826), .Y(n6540));
AOI22X1  g1498(.A0(g930), .A1(g823), .B0(g853), .B1(g933), .Y(n6541));
NAND4X1  g1554(.A(n6503), .B(n6485), .C(n6484_1), .D(n6504_1), .Y(n6597));
INVX1    g1350(.A(g809), .Y(n3442));
NOR2X1   g1406(.A(n6448), .B(n6447), .Y(n6449_1));
NOR2X1   g1369(.A(n6411), .B(n6410), .Y(n6412));
OR2X1    g1395(.A(n6437), .B(n6436), .Y(n6438));
NOR2X1   g1363(.A(n6405), .B(n6402), .Y(n6406));
NOR2X1   g1402(.A(n6444_1), .B(n6443), .Y(n6445));
OAI21X1  g1423(.A0(n6465), .A1(n6464_1), .B0(n3433), .Y(n6466));
INVX1    g1342(.A(g801), .Y(n3460));
NOR2X1   g1411(.A(n6453), .B(n6452), .Y(n6454_1));
INVX1    g1338(.A(g797), .Y(n3469));
NOR2X1   g1415(.A(n6457), .B(n6456), .Y(n6458));
INVX1    g1346(.A(g805), .Y(n3451));
NOR2X1   g1419(.A(n6461), .B(n6460), .Y(n6462));
NOR2X1   g1437(.A(n6479_1), .B(n6478), .Y(n6480));
INVX1    g1354(.A(g813), .Y(n3433));
NOR2X1   g1421(.A(g845), .B(n6401), .Y(n6464_1));
OAI22X1  g1422(.A0(g846), .A1(n6403), .B0(n6404_1), .B1(g844), .Y(n6465));
INVX1    g1334(.A(g793), .Y(n3478));
NOR2X1   g1429(.A(n6471), .B(n6470), .Y(n6472));
INVX1    g1330(.A(g789), .Y(n3487));
NOR2X1   g1433(.A(n6475), .B(n6474_1), .Y(n6476));
INVX1    g1358(.A(g826), .Y(n6401));
INVX1    g1361(.A(g853), .Y(n6404_1));
INVX1    g1360(.A(g823), .Y(n6403));
NOR3X1   g1455(.A(n6497), .B(n6493), .C(n6487), .Y(n6498));
OAI21X1  g1468(.A0(n6510), .A1(n6506), .B0(n6502), .Y(n6511));
NOR2X1   g1470(.A(n6510), .B(n6497), .Y(n6513));
OAI22X1  g1471(.A0(n6502), .A1(n6506), .B0(n6493), .B1(n6487), .Y(n6514_1));
XOR2X1   g1473(.A(n6509_1), .B(n3460), .Y(n6516));
NOR2X1   g1474(.A(n6502), .B(n6497), .Y(n6517));
NOR3X1   g1475(.A(n6506), .B(n6493), .C(n6487), .Y(n6518));
NOR3X1   g1492(.A(n6534_1), .B(n6530), .C(n6524_1), .Y(n6535));
OAI21X1  g1505(.A0(n6547), .A1(n6543), .B0(n6539_1), .Y(n6548));
NOR2X1   g1507(.A(n6547), .B(n6534_1), .Y(n6550));
OAI22X1  g1508(.A0(n6539_1), .A1(n6543), .B0(n6530), .B1(n6524_1), .Y(n6551));
XOR2X1   g1510(.A(n6546), .B(n3451), .Y(n6553));
NOR2X1   g1511(.A(n6539_1), .B(n6534_1), .Y(n6554_1));
NOR3X1   g1512(.A(n6543), .B(n6530), .C(n6524_1), .Y(n6555));
NOR2X1   g1529(.A(g1009), .B(n6559_1), .Y(n6572));
OAI22X1  g1530(.A0(g1010), .A1(n6561), .B0(n6562), .B1(g1008), .Y(n6573));
NOR2X1   g1404(.A(g842), .B(n6401), .Y(n6447));
OAI22X1  g1405(.A0(g843), .A1(n6403), .B0(n6404_1), .B1(g841), .Y(n6448));
NOR2X1   g1367(.A(g860), .B(n6401), .Y(n6410));
OAI22X1  g1368(.A0(g861), .A1(n6403), .B0(n6404_1), .B1(g859), .Y(n6411));
NOR2X1   g1393(.A(g851), .B(n6401), .Y(n6436));
OAI22X1  g1394(.A0(g852), .A1(n6403), .B0(n6404_1), .B1(g850), .Y(n6437));
NOR2X1   g1359(.A(g863), .B(n6401), .Y(n6402));
OAI22X1  g1362(.A0(g864), .A1(n6403), .B0(n6404_1), .B1(g862), .Y(n6405));
NOR2X1   g1400(.A(g848), .B(n6401), .Y(n6443));
OAI22X1  g1401(.A0(g849), .A1(n6403), .B0(n6404_1), .B1(g847), .Y(n6444_1));
NOR2X1   g1409(.A(g836), .B(n6401), .Y(n6452));
OAI22X1  g1410(.A0(g837), .A1(n6403), .B0(n6404_1), .B1(g835), .Y(n6453));
NOR2X1   g1413(.A(g833), .B(n6401), .Y(n6456));
OAI22X1  g1414(.A0(g834), .A1(n6403), .B0(n6404_1), .B1(g832), .Y(n6457));
NOR2X1   g1417(.A(g839), .B(n6401), .Y(n6460));
OAI22X1  g1418(.A0(g840), .A1(n6403), .B0(n6404_1), .B1(g838), .Y(n6461));
NOR2X1   g1435(.A(g818), .B(n6401), .Y(n6478));
OAI22X1  g1436(.A0(g819), .A1(n6403), .B0(n6404_1), .B1(g817), .Y(n6479_1));
NOR2X1   g1427(.A(g830), .B(n6401), .Y(n6470));
OAI22X1  g1428(.A0(g831), .A1(n6403), .B0(n6404_1), .B1(g829), .Y(n6471));
NOR2X1   g1431(.A(g821), .B(n6401), .Y(n6474_1));
OAI22X1  g1432(.A0(g822), .A1(n6403), .B0(n6404_1), .B1(g820), .Y(n6475));
NOR3X1   g1444(.A(n6486), .B(n6405), .C(n6402), .Y(n6487));
AOI21X1  g1450(.A0(n6491), .A1(n6488), .B0(n6492), .Y(n6493));
XOR2X1   g1454(.A(n6496), .B(g809), .Y(n6497));
XOR2X1   g1459(.A(n6501), .B(g785), .Y(n6502));
XOR2X1   g1463(.A(n6505), .B(g793), .Y(n6506));
XOR2X1   g1467(.A(n6509_1), .B(g801), .Y(n6510));
NAND2X1  g1466(.A(n6508), .B(n6507), .Y(n6509_1));
NOR3X1   g1481(.A(n6523), .B(n6411), .C(n6410), .Y(n6524_1));
AOI21X1  g1487(.A0(n6528), .A1(n6525), .B0(n6529_1), .Y(n6530));
XOR2X1   g1491(.A(n6533), .B(g813), .Y(n6534_1));
XOR2X1   g1496(.A(n6538), .B(g789), .Y(n6539_1));
XOR2X1   g1500(.A(n6542), .B(g797), .Y(n6543));
XOR2X1   g1504(.A(n6546), .B(g805), .Y(n6547));
AND2X1   g1443(.A(n6485), .B(n6484_1), .Y(n6486));
OR2X1    g1445(.A(g863), .B(n6401), .Y(n6488));
AOI22X1  g1448(.A0(n6489_1), .A1(g823), .B0(g853), .B1(n6490), .Y(n6491));
NAND2X1  g1453(.A(n6495), .B(n6494_1), .Y(n6496));
AND2X1   g1480(.A(n6522), .B(n6521), .Y(n6523));
OR2X1    g1482(.A(g860), .B(n6401), .Y(n6525));
AOI22X1  g1485(.A0(n6526), .A1(g823), .B0(g853), .B1(n6527), .Y(n6528));
INVX1    g1447(.A(g862), .Y(n6490));
INVX1    g1446(.A(g864), .Y(n6489_1));
INVX1    g1484(.A(g859), .Y(n6527));
INVX1    g1483(.A(g861), .Y(n6526));

endmodule
