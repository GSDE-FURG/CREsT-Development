// Benchmark "b22_C" written by ABC on Wed Aug 05 14:45:14 2020

module b22_C ( 
    P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
    SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_, SI_17_,
    SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_, SI_8_,
    SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
    P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
    P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
    P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
    P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
    P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
    P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
    P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
    P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
    P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
    P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN,
    P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN,
    P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN,
    P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN,
    P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN,
    P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
    P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
    P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
    P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
    P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
    P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
    P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
    P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
    P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
    P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
    P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
    P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
    P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
    P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
    P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
    P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
    P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN,
    P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
    P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN,
    P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN,
    P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
    P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
    P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
    P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
    P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
    P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
    P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
    P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
    P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
    P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
    P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
    P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
    P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
    P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
    P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
    P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
    P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
    P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
    P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
    P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
    P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
    P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
    P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
    P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
    P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
    P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
    P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
    P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
    P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
    P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
    P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
    P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
    P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
    P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
    P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
    P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
    P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
    P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
    P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
    P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
    P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
    P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
    P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
    P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
    P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
    P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
    P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
    P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
    P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
    P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
    P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
    P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
    P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
    P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
    P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
    P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
    P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
    P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
    P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
    P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
    P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
    P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
    P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
    P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
    P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
    P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
    P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
    P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
    P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
    P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
    P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
    P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
    P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
    P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
    P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
    P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
    P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
    P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
    P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
    P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
    P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
    P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
    P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
    P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
    P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
    P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
    P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
    P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
    P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
    P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
    P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
    P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
    P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
    P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
    P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
    P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
    P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
    P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
    P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
    P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
    P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
    P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
    P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
    P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
    P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
    P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
    P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
    P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
    P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
    P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
    P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
    P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
    P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
    P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
    P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
    P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
    P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
    P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
    P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
    P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
    P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
    P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
    P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
    P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
    P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
    P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
    P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
    P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
    P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
    P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
    P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
    P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
    P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
    P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
    P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
    P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
    P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
    P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
    P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
    P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
    P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
    P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
    P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
    P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
    P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
    P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
    P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
    P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
    P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
    P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
    P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
    P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
    P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
    P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
    P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
    P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
    P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
    P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
    P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
    P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
    P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
    P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
    P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
    P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
    P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
    P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
    P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
    P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
    P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
    P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
    P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
    P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
    P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
    P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
    P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
    P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
    P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
    P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
    P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
    P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
    P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
    P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
    P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
    P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
    P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
    P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
    P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
    P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
    P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
    P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
    P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
    P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
    P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
    P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
    P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
    P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
    P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
    P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
    P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN,
    P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN,
    P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN,
    P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN,
    P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN,
    P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN,
    P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN,
    P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN,
    P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN,
    P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN,
    P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN,
    P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN,
    P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN,
    P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN,
    P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN,
    P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN,
    P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN,
    P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN,
    P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN,
    P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN,
    P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN,
    P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN,
    P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN,
    P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN,
    P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN,
    P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN,
    P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN,
    P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN,
    P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN,
    P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN,
    P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN,
    P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN,
    P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
    P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN,
    P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
    P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
    P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
    P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
    P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
    P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
    P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
    P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
    P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
    P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
    P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
    P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
    P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN,
    P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
    P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN,
    P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN,
    P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN,
    P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN,
    P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN,
    P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN,
    P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN,
    P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN,
    P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN,
    P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN,
    P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN,
    P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN,
    P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN,
    P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
    P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN,
    P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
    P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
    P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
    P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
    P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
    P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
    P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
    P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
    P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
    P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
    P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
    P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
    P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
    P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
    P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
    P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
    P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN,
    SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
    SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
    SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
    SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
    U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
    P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
    P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
    P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
    P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
    P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
    P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
    P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
    P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
    P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
    P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
    P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
    P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
    P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
    P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
    P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
    P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
    P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
    P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
    P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
    P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
    P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
    P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
    P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
    P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
    P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
    P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
    P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
    P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
    P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
    P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
    P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
    P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
    P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
    P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
    P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
    P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
    P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
    P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
    P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
    P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
    P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
    P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
    P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
    P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
    P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
    P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
    P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
    P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
    P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
    P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
    P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
    P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
    P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
    P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
    P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
    P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
    P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
    P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
    P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
    P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
    P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
    P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
    P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
    P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
    P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
    P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
    P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
    P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
    P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
    P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
    P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
    P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
    P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
    P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
    P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
    P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
    P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
    P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
    P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
    P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
    P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
    P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
    P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
    P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
    P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
    P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
    P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
    P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
    P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
    P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
    P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
    P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
    P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
    P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
    P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
    P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
    P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
    P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
    P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
    P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
    P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
    P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
    P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
    P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
    P3_U3897  );
  input  P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_,
    SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
    SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
    SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
    P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
    P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
    P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
    P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
    P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
    P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
    P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
    P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
    P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
    P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN,
    P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN,
    P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN,
    P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN,
    P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN,
    P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
    P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
    P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
    P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
    P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
    P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
    P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
    P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
    P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
    P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
    P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
    P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
    P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
    P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
    P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
    P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
    P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN,
    P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
    P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN,
    P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN,
    P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN,
    P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN,
    P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN,
    P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN,
    P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN,
    P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN,
    P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN,
    P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN,
    P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN,
    P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN,
    P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN,
    P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN,
    P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN,
    P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN,
    P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN,
    P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN,
    P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN,
    P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN,
    P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN,
    P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN,
    P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN,
    P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
    P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
    P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
    P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
    P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
    P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
    P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
    P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
    P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
    P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
    P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
    P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
    P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
    P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
    P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
    P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
    P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
    P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
    P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
    P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
    P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
    P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
    P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
    P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
    P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
    P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
    P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
    P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
    P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
    P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
    P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
    P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
    P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
    P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
    P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
    P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
    P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
    P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
    P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
    P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
    P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
    P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
    P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
    P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
    P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
    P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
    P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
    P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
    P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
    P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
    P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
    P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
    P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
    P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
    P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
    P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
    P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
    P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
    P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
    P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
    P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
    P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
    P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
    P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
    P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
    P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
    P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
    P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
    P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
    P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
    P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
    P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
    P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
    P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
    P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
    P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
    P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
    P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
    P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
    P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
    P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
    P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
    P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
    P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
    P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
    P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
    P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
    P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
    P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
    P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
    P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
    P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
    P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
    P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
    P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
    P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
    P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
    P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
    P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
    P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
    P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
    P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
    P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
    P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
    P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
    P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
    P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
    P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
    P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
    P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
    P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
    P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
    P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
    P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
    P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
    P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
    P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
    P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
    P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
    P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
    P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
    P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
    P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
    P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
    P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
    P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
    P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
    P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
    P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
    P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
    P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
    P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
    P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
    P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
    P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
    P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
    P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
    P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
    P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
    P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
    P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
    P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
    P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
    P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
    P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
    P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
    P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
    P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
    P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
    P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
    P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
    P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
    P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
    P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
    P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
    P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
    P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
    P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
    P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
    P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
    P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
    P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
    P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
    P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
    P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
    P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
    P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
    P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
    P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
    P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
    P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
    P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
    P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
    P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
    P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
    P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
    P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
    P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN,
    P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN,
    P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN,
    P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN,
    P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN,
    P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN,
    P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN,
    P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN,
    P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN,
    P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN,
    P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN,
    P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN,
    P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN,
    P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN,
    P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN,
    P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN,
    P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN,
    P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN,
    P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN,
    P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN,
    P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN,
    P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN,
    P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN,
    P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN,
    P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN,
    P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN,
    P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN,
    P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN,
    P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN,
    P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN,
    P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN,
    P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN,
    P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
    P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN,
    P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
    P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
    P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
    P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
    P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
    P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
    P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
    P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
    P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
    P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
    P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
    P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
    P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN,
    P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
    P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN,
    P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN,
    P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN,
    P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN,
    P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN,
    P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN,
    P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN,
    P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN,
    P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN,
    P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN,
    P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN,
    P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN,
    P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN,
    P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
    P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN,
    P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
    P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
    P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
    P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
    P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
    P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
    P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
    P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
    P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
    P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
    P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
    P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
    P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
    P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
    P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
    P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
    P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
    SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
    SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
    SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
    U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
    P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
    P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
    P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
    P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
    P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
    P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
    P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
    P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
    P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
    P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
    P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
    P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
    P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
    P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
    P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
    P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
    P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
    P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
    P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
    P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
    P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
    P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
    P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
    P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
    P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
    P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
    P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
    P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
    P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
    P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
    P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
    P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
    P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
    P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
    P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
    P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
    P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
    P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
    P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
    P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
    P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
    P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
    P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
    P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
    P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
    P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
    P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
    P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
    P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
    P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
    P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
    P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
    P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
    P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
    P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
    P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
    P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
    P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
    P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
    P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
    P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
    P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
    P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
    P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
    P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
    P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
    P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
    P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
    P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
    P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
    P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
    P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
    P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
    P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
    P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
    P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
    P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
    P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
    P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
    P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
    P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
    P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
    P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
    P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
    P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
    P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
    P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
    P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
    P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
    P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
    P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
    P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
    P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
    P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
    P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
    P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
    P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
    P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
    P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
    P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
    P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
    P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
    P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
    P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
    P3_U3897;
  wire n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
    n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
    n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
    n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
    n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
    n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
    n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
    n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
    n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
    n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
    n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
    n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
    n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
    n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
    n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
    n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
    n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
    n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
    n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
    n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
    n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1733, n1735,
    n1737, n1739, n1740, n1742, n1744, n1745, n1747, n1748, n1750, n1751,
    n1753, n1754, n1756, n1757, n1759, n1761, n1763, n1765, n1767, n1769,
    n1771, n1773, n1774, n1775, n1776, n1779, n1780, n1782, n1783, n1785,
    n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
    n1796, n1797, n1798, n1799, n1800, n1801, n1803, n1804, n1806, n1807,
    n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
    n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
    n1828, n1829, n1830, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
    n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1848, n1849,
    n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
    n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
    n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
    n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
    n1891, n1892, n1893, n1894, n1895, n1896, n1898, n1899, n1900, n1901,
    n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
    n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
    n1922, n1923, n1924, n1925, n1927, n1928, n1929, n1930, n1931, n1932,
    n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
    n1943, n1944, n1945, n1946, n1947, n1948, n1950, n1951, n1952, n1953,
    n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
    n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1974,
    n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
    n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
    n1995, n1996, n1997, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
    n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
    n2016, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
    n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
    n2037, n2038, n2039, n2040, n2041, n2043, n2044, n2045, n2046, n2047,
    n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
    n2058, n2059, n2060, n2061, n2062, n2063, n2065, n2066, n2067, n2068,
    n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
    n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2088, n2089,
    n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
    n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2109, n2110,
    n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
    n2121, n2122, n2123, n2124, n2125, n2126, n2128, n2129, n2130, n2131,
    n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
    n2142, n2143, n2144, n2145, n2146, n2148, n2149, n2150, n2151, n2152,
    n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
    n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
    n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2181, n2182, n2183,
    n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
    n2194, n2195, n2196, n2197, n2199, n2200, n2201, n2202, n2203, n2204,
    n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
    n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
    n2225, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
    n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
    n2246, n2247, n2248, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
    n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
    n2267, n2268, n2269, n2270, n2271, n2272, n2274, n2275, n2276, n2277,
    n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
    n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
    n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
    n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2319,
    n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
    n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2338, n2339, n2340,
    n2341, n2342, n2343, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
    n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
    n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2371, n2372,
    n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
    n2383, n2384, n2385, n2386, n2387, n2389, n2390, n2391, n2392, n2393,
    n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
    n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
    n2414, n2415, n2416, n2417, n2418, n2419, n2421, n2422, n2423, n2424,
    n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
    n2435, n2436, n2437, n2438, n2439, n2441, n2442, n2443, n2444, n2445,
    n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
    n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2466,
    n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
    n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
    n2487, n2488, n2489, n2490, n2492, n2493, n2494, n2495, n2496, n2497,
    n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
    n2508, n2509, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
    n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
    n2529, n2530, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
    n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
    n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
    n2560, n2561, n2562, n2564, n2565, n2566, n2568, n2570, n2572, n2574,
    n2576, n2578, n2580, n2582, n2584, n2586, n2588, n2590, n2592, n2594,
    n2596, n2598, n2600, n2602, n2604, n2606, n2608, n2610, n2612, n2614,
    n2616, n2618, n2620, n2622, n2624, n2626, n2628, n2629, n2630, n2631,
    n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
    n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
    n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
    n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
    n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
    n2682, n2683, n2684, n2685, n2686, n2687, n2691, n2692, n2693, n2694,
    n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
    n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2713, n2714, n2715,
    n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
    n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
    n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
    n2746, n2747, n2748, n2749, n2751, n2752, n2753, n2754, n2755, n2756,
    n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
    n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
    n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
    n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
    n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2806, n2807,
    n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
    n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
    n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
    n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
    n2848, n2849, n2850, n2851, n2852, n2854, n2855, n2856, n2857, n2858,
    n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
    n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
    n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
    n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
    n2899, n2900, n2901, n2902, n2903, n2905, n2906, n2907, n2908, n2909,
    n2910, n2911, n2912, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
    n2921, n2922, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
    n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
    n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
    n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
    n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
    n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
    n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
    n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3003,
    n3004, n3005, n3006, n3007, n3008, n3010, n3011, n3012, n3013, n3014,
    n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
    n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
    n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
    n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
    n3055, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
    n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
    n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
    n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
    n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
    n3106, n3107, n3108, n3109, n3111, n3112, n3113, n3114, n3115, n3116,
    n3117, n3118, n3119, n3120, n3121, n3123, n3124, n3125, n3126, n3127,
    n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
    n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
    n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
    n3158, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
    n3169, n3170, n3171, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
    n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
    n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
    n3200, n3201, n3202, n3203, n3204, n3206, n3207, n3208, n3209, n3210,
    n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3221, n3222,
    n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
    n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
    n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3252, n3253,
    n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
    n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3274,
    n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
    n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
    n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
    n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
    n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
    n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
    n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
    n3347, n3348, n3349, n3350, n3351, n3353, n3354, n3355, n3356, n3357,
    n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
    n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
    n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
    n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
    n3398, n3399, n3400, n3401, n3402, n3403, n3405, n3406, n3407, n3408,
    n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
    n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
    n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
    n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3448, n3449,
    n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
    n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
    n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
    n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3489, n3490,
    n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
    n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
    n3511, n3512, n3513, n3514, n3515, n3517, n3518, n3519, n3520, n3521,
    n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
    n3532, n3533, n3534, n3535, n3536, n3537, n3539, n3540, n3541, n3542,
    n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3554,
    n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
    n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
    n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3585,
    n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
    n3596, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
    n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
    n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3626, n3627,
    n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
    n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3648,
    n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
    n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
    n3669, n3670, n3671, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
    n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
    n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
    n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
    n3710, n3711, n3712, n3713, n3715, n3716, n3717, n3718, n3719, n3720,
    n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
    n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
    n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
    n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3761,
    n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
    n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
    n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
    n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3802, n3803, n3804,
    n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
    n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
    n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
    n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3845,
    n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857,
    n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867,
    n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877,
    n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3887, n3888,
    n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
    n3899, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
    n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
    n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
    n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
    n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
    n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
    n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
    n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3980, n3981,
    n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3991, n3992,
    n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
    n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
    n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
    n4023, n4024, n4025, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
    n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4042, n4043, n4044,
    n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
    n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
    n4065, n4066, n4067, n4068, n4069, n4071, n4072, n4073, n4074, n4075,
    n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
    n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
    n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
    n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
    n4116, n4117, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
    n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
    n4137, n4138, n4140, n4141, n4142, n4143, n4144, n4145, n4147, n4148,
    n4149, n4151, n4153, n4155, n4157, n4159, n4161, n4163, n4165, n4167,
    n4169, n4171, n4173, n4175, n4177, n4179, n4181, n4183, n4185, n4187,
    n4189, n4191, n4193, n4195, n4197, n4199, n4201, n4203, n4205, n4207,
    n4209, n4211, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
    n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
    n4231, n4232, n4233, n4235, n4236, n4237, n4238, n4239, n4241, n4242,
    n4243, n4244, n4245, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
    n4254, n4255, n4256, n4257, n4258, n4260, n4261, n4262, n4263, n4264,
    n4265, n4266, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4276,
    n4277, n4278, n4279, n4280, n4281, n4282, n4284, n4285, n4286, n4287,
    n4288, n4289, n4290, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
    n4300, n4301, n4302, n4303, n4304, n4305, n4307, n4308, n4309, n4310,
    n4311, n4312, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
    n4322, n4324, n4325, n4326, n4327, n4328, n4329, n4331, n4332, n4333,
    n4334, n4335, n4336, n4337, n4339, n4340, n4341, n4342, n4343, n4344,
    n4346, n4347, n4348, n4349, n4350, n4352, n4353, n4354, n4355, n4356,
    n4357, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4368,
    n4369, n4370, n4371, n4372, n4373, n4375, n4376, n4377, n4378, n4379,
    n4380, n4381, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4391,
    n4392, n4393, n4394, n4395, n4396, n4397, n4399, n4400, n4401, n4402,
    n4403, n4404, n4405, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
    n4414, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4425,
    n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4434, n4435, n4436,
    n4437, n4438, n4439, n4440, n4441, n4442, n4444, n4445, n4446, n4447,
    n4448, n4449, n4450, n4451, n4453, n4454, n4455, n4456, n4457, n4458,
    n4459, n4460, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
    n4471, n4472, n4473, n4474, n4476, n4477, n4478, n4479, n4480, n4481,
    n4482, n4483, n4484, n4486, n4487, n4488, n4489, n4491, n4492, n4493,
    n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
    n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
    n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
    n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
    n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
    n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
    n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
    n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
    n4574, n4575, n4576, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
    n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
    n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
    n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
    n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
    n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
    n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
    n4646, n4647, n4648, n4649, n4650, n4651, n4654, n4657, n4658, n4659,
    n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
    n4671, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
    n4682, n4683, n4684, n4685, n4686, n4688, n4689, n4690, n4691, n4692,
    n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
    n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4711, n4712, n4713,
    n4714, n4715, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
    n4725, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
    n4736, n4737, n4738, n4740, n4741, n4742, n4743, n4744, n4745, n4746,
    n4747, n4748, n4749, n4750, n4751, n4753, n4754, n4755, n4756, n4757,
    n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
    n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
    n4778, n4779, n4780, n4781, n4783, n4784, n4785, n4786, n4787, n4789,
    n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4799, n4801,
    n4802, n4803, n4804, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
    n4813, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
    n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
    n4834, n4835, n4836, n4837, n4838, n4840, n4842, n4843, n4844, n4845,
    n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4856, n4857,
    n4858, n4860, n4861, n4862, n4864, n4865, n4866, n4867, n4868, n4869,
    n4870, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
    n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
    n4891, n4892, n4893, n4894, n4896, n4897, n4898, n4899, n4900, n4901,
    n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
    n4912, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
    n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
    n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
    n4943, n4944, n4945, n4946, n4947, n4948, n4950, n4952, n4953, n4954,
    n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
    n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
    n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
    n4985, n4986, n4988, n4989, n4990, n4992, n4993, n4994, n4995, n4996,
    n4997, n4998, n4999, n5000, n5002, n5003, n5004, n5005, n5006, n5007,
    n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5017, n5018,
    n5020, n5021, n5022, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
    n5031, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
    n5042, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5053,
    n5055, n5057, n5059, n5061, n5063, n5065, n5067, n5069, n5070, n5072,
    n5074, n5076, n5077, n5079, n5080, n5082, n5084, n5086, n5088, n5090,
    n5092, n5094, n5096, n5098, n5100, n5102, n5104, n5106, n5108, n5110,
    n5112, n5114, n5116, n5117, n5118, n5119, n5121, n5122, n5123, n5124,
    n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
    n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
    n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
    n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
    n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
    n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
    n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
    n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
    n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
    n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
    n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
    n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
    n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
    n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
    n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
    n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
    n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
    n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
    n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
    n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
    n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
    n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
    n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
    n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
    n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
    n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
    n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
    n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
    n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
    n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
    n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
    n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
    n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
    n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
    n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
    n5477, n5478, n5480, n5481, n5484, n5487, n5490, n5491, n5492, n5493,
    n5494, n5495, n5496, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
    n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
    n5515, n5516, n5517, n5518, n5520, n5521, n5522, n5523, n5524, n5525,
    n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
    n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
    n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
    n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
    n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
    n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
    n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
    n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
    n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
    n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
    n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
    n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
    n5646, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656,
    n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666,
    n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676,
    n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686,
    n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696,
    n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706,
    n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716,
    n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726,
    n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
    n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
    n5747, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5758, n5759,
    n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5769, n5770, n5771,
    n5772, n5773, n5774, n5775, n5777, n5778, n5780, n5781, n5782, n5783,
    n5784, n5785, n5786, n5788, n5789, n5791, n5792, n5793, n5794, n5795,
    n5796, n5797, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806,
    n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
    n5818, n5819, n5820, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
    n5829, n5830, n5831, n5832, n5833, n5835, n5836, n5837, n5838, n5839,
    n5840, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5851,
    n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5861, n5862,
    n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5871, n5872, n5873,
    n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
    n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
    n5896, n5897, n5899, n5900, n5901, n5902, n5903, n5904, n5906, n5908,
    n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5917, n5919, n5920,
    n5921, n5922, n5923, n5924, n5925, n5927, n5928, n5929, n5930, n5931,
    n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5940, n5941, n5942,
    n5943, n5944, n5945, n5946, n5947, n5949, n5950, n5951, n5952, n5953,
    n5954, n5955, n5956, n5957, n5959, n5960, n5961, n5962, n5963, n5964,
    n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
    n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
    n5985, n5987, n5988, n5989, n5991, n5992, n5993, n5994, n5995, n5996,
    n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
    n6008, n6009, n6010, n6011, n6012, n6014, n6015, n6016, n6017, n6018,
    n6019, n6020, n6021, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
    n6030, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6040, n6041,
    n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6050, n6051, n6052,
    n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
    n6064, n6065, n6067, n6068, n6070, n6071, n6072, n6073, n6074, n6075,
    n6077, n6078, n6079, n6080, n6081, n6082, n6084, n6085, n6086, n6087,
    n6088, n6089, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
    n6099, n6100, n6102, n6103, n6104, n6105, n6106, n6107, n6109, n6110,
    n6111, n6112, n6113, n6114, n6115, n6117, n6118, n6119, n6120, n6121,
    n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6132, n6133,
    n6134, n6135, n6136, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
    n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6155, n6156,
    n6157, n6158, n6159, n6160, n6162, n6163, n6164, n6165, n6166, n6168,
    n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6177, n6178, n6179,
    n6180, n6181, n6182, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
    n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6201,
    n6202, n6203, n6204, n6205, n6206, n6208, n6209, n6210, n6211, n6212,
    n6213, n6214, n6215, n6216, n6217, n6219, n6220, n6221, n6222, n6223,
    n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6234, n6235,
    n6236, n6237, n6238, n6239, n6240, n6242, n6243, n6244, n6245, n6246,
    n6247, n6248, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257,
    n6259, n6260, n6261, n6262, n6263, n6264, n6266, n6267, n6268, n6269,
    n6270, n6271, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
    n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
    n6291, n6292, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6302,
    n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6312, n6313,
    n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
    n6324, n6325, n6327, n6328, n6329, n6330, n6331, n6332, n6334, n6335,
    n6336, n6337, n6338, n6340, n6341, n6342, n6343, n6344, n6345, n6346,
    n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356,
    n6357, n6358, n6359, n6361, n6362, n6363, n6365, n6367, n6369, n6371,
    n6373, n6375, n6377, n6379, n6381, n6383, n6385, n6387, n6389, n6391,
    n6393, n6395, n6397, n6399, n6401, n6403, n6405, n6407, n6409, n6411,
    n6413, n6415, n6417, n6419, n6421, n6423, n6425, n6426, n6427, n6428,
    n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
    n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
    n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
    n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
    n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6479, n6480, n6481,
    n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
    n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
    n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6512,
    n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
    n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
    n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
    n6543, n6544, n6545, n6546, n6547, n6549, n6550, n6551, n6552, n6553,
    n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
    n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
    n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
    n6584, n6585, n6586, n6587, n6589, n6590, n6591, n6592, n6593, n6594,
    n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
    n6605, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
    n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
    n6626, n6627, n6628, n6629, n6630, n6631, n6633, n6634, n6635, n6636,
    n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
    n6647, n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657,
    n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
    n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677,
    n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687,
    n6688, n6689, n6690, n6692, n6699, n6700, n6701, n6702, n6703, n6704,
    n6705, n6706, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716,
    n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726,
    n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736,
    n6737, n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747,
    n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757,
    n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767,
    n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777,
    n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787,
    n6788, n6789, n6790, n6791, n6793, n6794, n6795, n6796, n6797, n6798,
    n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
    n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
    n6820, n6821, n6822, n6823, n6830, n6831, n6832, n6833, n6834, n6835,
    n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
    n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856,
    n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866,
    n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876,
    n6877, n6878, n6879, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
    n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
    n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
    n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
    n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6934, n6935,
    n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
    n6946, n6947, n6948, n6949, n6950, n6952, n6953, n6954, n6955, n6956,
    n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
    n6967, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977,
    n6978, n6979, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
    n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n7000, n7001,
    n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
    n7012, n7013, n7014, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
    n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
    n7033, n7034, n7035, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
    n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
    n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067,
    n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077,
    n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
    n7089, n7090, n7091, n7092, n7096, n7097, n7098, n7099, n7100, n7101,
    n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7111, n7112,
    n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
    n7123, n7124, n7125, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
    n7134, n7135, n7136, n7137, n7138, n7139, n7144, n7145, n7146, n7147,
    n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
    n7158, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
    n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
    n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
    n7189, n7190, n7191, n7192, n7193, n7194, n7199, n7200, n7201, n7202,
    n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
    n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
    n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
    n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7245,
    n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
    n7256, n7257, n7258, n7259, n7261, n7262, n7263, n7264, n7265, n7266,
    n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276,
    n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286,
    n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7295, n7296, n7297,
    n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307,
    n7308, n7309, n7310, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
    n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
    n7329, n7330, n7331, n7333, n7334, n7335, n7336, n7338, n7341, n7342,
    n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
    n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
    n7363, n7364, n7365, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
    n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7384,
    n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
    n7395, n7396, n7397, n7398, n7399, n7400, n7403, n7405, n7406, n7407,
    n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417,
    n7418, n7419, n7421, n7422, n7423, n7424, n7425, n7426, n7428, n7429,
    n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
    n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7448, n7449, n7452,
    n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
    n7463, n7464, n7465, n7466, n7467, n7469, n7470, n7471, n7472, n7473,
    n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
    n7484, n7485, n7486, n7487, n7489, n7490, n7491, n7492, n7493, n7494,
    n7495, n7497, n7498, n7499, n7500, n7502, n7503, n7504, n7505, n7506,
    n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7517,
    n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
    n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
    n7540, n7541, n7542, n7543, n7544, n7545, n7548, n7549, n7550, n7551,
    n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561,
    n7562, n7563, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
    n7573, n7574, n7575, n7576, n7577, n7579, n7580, n7581, n7582, n7583,
    n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
    n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
    n7604, n7605, n7606, n7608, n7609, n7611, n7612, n7613, n7614, n7615,
    n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
    n7626, n7627, n7628, n7629, n7630, n7631, n7633, n7634, n7635, n7636,
    n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646,
    n7647, n7648, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657,
    n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667,
    n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677,
    n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
    n7689, n7690, n7691, n7692, n7694, n7695, n7696, n7698, n7699, n7700,
    n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710,
    n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720,
    n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
    n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
    n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
    n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
    n7762, n7763, n7764, n7765, n7766, n7768, n7769, n7770, n7771, n7772,
    n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
    n7783, n7784, n7785, n7787, n7788, n7789, n7790, n7791, n7795, n7796,
    n7797, n7798, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
    n7808, n7809, n7810, n7811, n7812, n7815, n7816, n7817, n7818, n7819,
    n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
    n7830, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
    n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
    n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
    n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
    n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
    n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
    n7891, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901,
    n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911,
    n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
    n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931,
    n7932, n7933, n7934, n7935, n7936, n7937, n7939, n7940, n7941, n7942,
    n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
    n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
    n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7972, n7973,
    n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7983, n7984,
    n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7995,
    n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8005, n8006,
    n8007, n8009, n8011, n8013, n8015, n8017, n8019, n8021, n8023, n8025,
    n8027, n8029, n8031, n8033, n8035, n8037, n8039, n8041, n8043, n8045,
    n8047, n8049, n8051, n8053, n8055, n8057, n8059, n8061, n8063, n8065,
    n8067, n8069, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
    n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8089,
    n8090, n8091, n8093, n8094, n8095, n8096, n8097, n8098, n8100, n8101,
    n8102, n8103, n8104, n8106, n8107, n8108, n8109, n8110, n8111, n8113,
    n8114, n8115, n8116, n8117, n8118, n8120, n8121, n8122, n8123, n8125,
    n8126, n8127, n8128, n8129, n8130, n8131, n8133, n8134, n8135, n8136,
    n8137, n8138, n8139, n8140, n8141, n8143, n8144, n8145, n8146, n8147,
    n8149, n8150, n8151, n8152, n8153, n8154, n8156, n8157, n8158, n8159,
    n8160, n8161, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8171,
    n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8180, n8181, n8182,
    n8183, n8184, n8185, n8186, n8188, n8189, n8190, n8191, n8192, n8193,
    n8195, n8196, n8197, n8198, n8199, n8200, n8202, n8203, n8204, n8205,
    n8206, n8207, n8208, n8210, n8211, n8212, n8213, n8214, n8215, n8216,
    n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8226, n8228, n8229,
    n8230, n8231, n8232, n8234, n8236, n8237, n8238, n8239, n8240, n8241,
    n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8253,
    n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8263, n8264,
    n8265, n8266, n8267, n8268, n8269, n8271, n8272, n8273, n8274, n8275,
    n8276, n8277, n8278, n8280, n8281, n8282, n8283, n8284, n8285, n8286,
    n8287, n8288, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8298,
    n8300, n8301, n8302, n8303, n8304, n8305, n8307, n8308, n8309, n8310,
    n8311, n8312, n8313, n8314, n8316, n8317, n8318, n8319, n8320, n8321,
    n8322, n8324, n8325, n8326, n8327, n8328, n8329, n8331, n8332, n8333,
    n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
    n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
    n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
    n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
    n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
    n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
    n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
    n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
    n8415, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
    n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
    n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
    n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
    n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
    n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
    n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
    n8486, n8487, n8490, n8491, n8492, n8493, n8495, n8496, n8497, n8498,
    n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
    n8509, n8510, n8511, n8512, n8513, n8515, n8516, n8517, n8518, n8519,
    n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
    n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540,
    n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550,
    n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8559, n8561, n8562,
    n8563, n8564, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
    n8574, n8575, n8576, n8577, n8579, n8580, n8581, n8582, n8583, n8584,
    n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
    n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
    n8606, n8607, n8608, n8609, n8610, n8612, n8613, n8614, n8615, n8616,
    n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626,
    n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636,
    n8637, n8638, n8639, n8640, n8641, n8643, n8645, n8646, n8647, n8648,
    n8649, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
    n8660, n8661, n8663, n8664, n8665, n8667, n8668, n8669, n8670, n8671,
    n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8681, n8682,
    n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
    n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
    n8703, n8704, n8705, n8706, n8707, n8708, n8710, n8711, n8713, n8714,
    n8715, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
    n8726, n8727, n8729, n8730, n8731, n8733, n8734, n8735, n8737, n8738,
    n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8747, n8748, n8749,
    n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
    n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
    n8770, n8771, n8772, n8774, n8775, n8776, n8779, n8780, n8781, n8782,
    n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
    n8793, n8794, n8795, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
    n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
    n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
    n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
    n8834, n8836, n8837, n8839, n8840, n8841, n8843, n8844, n8845, n8846,
    n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8856, n8857,
    n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867,
    n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8876, n8877, n8878,
    n8880, n8881, n8882, n8883, n8885, n8886, n8887, n8888, n8889, n8890,
    n8891, n8892, n8893, n8894, n8895, n8896, n8898, n8899, n8900, n8901,
    n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911,
    n8912, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
    n8923, n8924, n8925, n8926, n8927, n8928, n8930, n8932, n8934, n8936,
    n8938, n8940, n8942, n8944, n8946, n8948, n8950, n8952, n8954, n8956,
    n8958, n8960, n8962, n8964, n8966, n8968, n8970, n8972, n8974, n8976,
    n8978, n8980, n8982, n8984, n8986, n8988, n8990, n8991, n8993, n8994,
    n8996, n8997, n8998, n8999, n9000, n9001, n9004, n9005, n9006, n9007,
    n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017,
    n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027,
    n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037,
    n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047,
    n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057,
    n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067,
    n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077,
    n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087,
    n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097,
    n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107,
    n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117,
    n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127,
    n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137,
    n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
    n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
    n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
    n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
    n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
    n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
    n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
    n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
    n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
    n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
    n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
    n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257,
    n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267,
    n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277,
    n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287,
    n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297,
    n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307,
    n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
    n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327,
    n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337,
    n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347,
    n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357,
    n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
    n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377,
    n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387,
    n9388, n9389, n9390, n9391, n9395, n9396, n9397, n9398, n9401, n9403,
    n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
    n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
    n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9432, n9434, n9435,
    n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
    n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
    n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
    n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
    n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
    n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
    n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
    n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
    n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
    n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
    n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
    n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9556,
    n9557, n9558, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567,
    n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577,
    n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587,
    n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597,
    n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607,
    n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617,
    n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627,
    n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637,
    n9638, n9639, n9640, n9641, n9644, n9646, n9647, n9648, n9650, n9651,
    n9652, n9653, n9654, n9655, n9656, n9657, n9659, n9660, n9661, n9662,
    n9663, n9664, n9665, n9666, n9668, n9669, n9670, n9671, n9672, n9673,
    n9674, n9675, n9676, n9677, n9678, n9679, n9681, n9682, n9683, n9684,
    n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9695,
    n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9704, n9705, n9706,
    n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
    n9717, n9718, n9720, n9721, n9722, n9724, n9725, n9726, n9727, n9728,
    n9729, n9730, n9731, n9733, n9734, n9735, n9737, n9738, n9739, n9740,
    n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9750, n9751, n9752,
    n9753, n9754, n9755, n9756, n9757, n9759, n9761, n9762, n9763, n9764,
    n9765, n9766, n9767, n9768, n9770, n9771, n9772, n9773, n9774, n9775,
    n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9784, n9785, n9786,
    n9787, n9788, n9789, n9790, n9791, n9793, n9795, n9796, n9797, n9798,
    n9799, n9800, n9801, n9803, n9805, n9806, n9807, n9808, n9809, n9810,
    n9811, n9812, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
    n9822, n9823, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
    n9833, n9834, n9835, n9836, n9837, n9839, n9840, n9841, n9842, n9843,
    n9844, n9845, n9846, n9847, n9849, n9850, n9851, n9852, n9853, n9854,
    n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9863, n9864, n9865,
    n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
    n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
    n9886, n9887, n9888, n9890, n9892, n9893, n9894, n9895, n9896, n9897,
    n9898, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
    n9909, n9910, n9911, n9912, n9913, n9914, n9916, n9917, n9918, n9919,
    n9920, n9921, n9922, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
    n9931, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9942,
    n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9952, n9953,
    n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
    n9964, n9966, n9967, n9968, n9970, n9971, n9972, n9973, n9975, n9976,
    n9977, n9978, n9979, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
    n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
    n9999, n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
    n10009, n10010, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
    n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
    n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
    n10038, n10039, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
    n10048, n10049, n10050, n10051, n10052, n10053, n10055, n10056, n10057,
    n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
    n10067, n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
    n10077, n10078, n10079, n10080, n10081, n10083, n10084, n10085, n10086,
    n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
    n10096, n10097, n10098, n10099, n10101, n10102, n10103, n10104, n10105,
    n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10114, n10115,
    n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
    n10125, n10126, n10127, n10129, n10130, n10131, n10132, n10133, n10134,
    n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
    n10144, n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
    n10154, n10155, n10156, n10157, n10158, n10160, n10161, n10162, n10163,
    n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
    n10173, n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182,
    n10183, n10184, n10185, n10187, n10188, n10189, n10190, n10191, n10192,
    n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
    n10202, n10203, n10204, n10205, n10206, n10207, n10209, n10210, n10211,
    n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10221,
    n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
    n10231, n10232, n10233, n10234, n10236, n10237, n10238, n10239, n10240,
    n10241, n10242, n10243, n10244, n10245, n10246, n10248, n10249, n10250,
    n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
    n10260, n10261, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
    n10270, n10271, n10272, n10273, n10275, n10276, n10277, n10278, n10279,
    n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
    n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
    n10299, n10300, n10301, n10302, n10304, n10305, n10306, n10307, n10308,
    n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
    n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
    n10328, n10329, n10330, n10332, n10333, n10334, n10335, n10336, n10337,
    n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
    n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356,
    n10357, n10358, n10359, n10361, n10362, n10363, n10364, n10365, n10366,
    n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
    n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
    n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
    n10394, n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
    n10404, n10405, n10406, n10407, n10408, n10409, n10411, n10412, n10413,
    n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422,
    n10423, n10424, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
    n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
    n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
    n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459, n10460,
    n10461, n10463, n10464, n10465, n10467, n10469, n10471, n10473, n10475,
    n10477, n10479, n10481, n10483, n10485, n10487, n10489, n10491, n10493,
    n10495, n10497, n10499, n10501, n10503, n10505, n10507, n10509, n10511,
    n10513, n10515, n10517, n10519, n10521, n10523, n10525, n10527, n10528,
    n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
    n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
    n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
    n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564,
    n10565, n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573,
    n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582,
    n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
    n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
    n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
    n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
    n10619, n10620, n10622, n10623, n10624, n10625, n10626, n10627, n10628,
    n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637,
    n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646,
    n10647, n10648, n10649, n10650, n10652, n10653, n10654, n10655, n10656,
    n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
    n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
    n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
    n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692,
    n10693, n10694, n10695, n10697, n10698, n10699, n10700, n10701, n10702,
    n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
    n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
    n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
    n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
    n10739, n10740, n10741, n10742, n10744, n10745, n10746, n10747, n10748,
    n10749, n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757,
    n10758, n10759, n10760, n10761, n10762, n10764, n10765, n10766, n10767,
    n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
    n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
    n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,
    n10795, n10796, n10797, n10799, n10800, n10801, n10802, n10803, n10804,
    n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814,
    n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
    n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
    n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
    n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10850, n10851,
    n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859, n10860,
    n10861, n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869,
    n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878,
    n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
    n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
    n10897, n10898, n10899, n10900, n10901, n10903, n10904, n10905, n10906,
    n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
    n10916, n10917, n10918, n10919, n10920, n10921, n10923, n10924, n10925,
    n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934,
    n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
    n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10952, n10953,
    n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,
    n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971,
    n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980,
    n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989,
    n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998,
    n10999, n11000, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
    n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11018,
    n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
    n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036,
    n11037, n11038, n11039, n11040, n11042, n11043, n11044, n11045, n11046,
    n11047, n11048, n11049, n11050, n11051, n11052, n11054, n11055, n11056,
    n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
    n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
    n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
    n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11092, n11093,
    n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102,
    n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
    n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
    n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
    n11130, n11131, n11132, n11133, n11134, n11135, n11137, n11138, n11139,
    n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148,
    n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157,
    n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
    n11167, n11168, n11169, n11170, n11171, n11172, n11180, n11181, n11182,
    n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
    n11192, n11193, n11194, n11195, n11197, n11198, n11199, n11200, n11201,
    n11202, n11203, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
    n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220,
    n11221, n11222, n11223, n11224, n11225, n11229, n11230, n11231, n11232,
    n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
    n11242, n11243, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
    n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260,
    n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269,
    n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278,
    n11279, n11280, n11281, n11282, n11286, n11287, n11288, n11289, n11290,
    n11291, n11292, n11293, n11294, n11295, n11296, n11298, n11299, n11300,
    n11301, n11302, n11303, n11305, n11306, n11307, n11308, n11309, n11310,
    n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
    n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
    n11330, n11331, n11332, n11333, n11334, n11335, n11337, n11338, n11339,
    n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348,
    n11349, n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
    n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
    n11368, n11369, n11370, n11371, n11372, n11373, n11375, n11376, n11377,
    n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
    n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
    n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404,
    n11405, n11406, n11407, n11408, n11409, n11410, n11414, n11415, n11416,
    n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
    n11426, n11427, n11428, n11430, n11431, n11432, n11433, n11434, n11435,
    n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444,
    n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454,
    n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
    n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
    n11473, n11474, n11475, n11476, n11477, n11479, n11480, n11481, n11482,
    n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
    n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11501,
    n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
    n11514, n11515, n11516, n11517, n11518, n11519, n11521, n11522, n11523,
    n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532,
    n11533, n11534, n11535, n11536, n11537, n11540, n11541, n11542, n11543,
    n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
    n11556, n11557, n11558, n11560, n11561, n11562, n11563, n11564, n11565,
    n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574,
    n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
    n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
    n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
    n11602, n11603, n11604, n11605, n11607, n11608, n11609, n11610, n11611,
    n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620,
    n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
    n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
    n11642, n11643, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
    n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660,
    n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669,
    n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11680,
    n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
    n11690, n11691, n11692, n11693, n11694, n11695, n11697, n11698, n11699,
    n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708,
    n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717,
    n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
    n11729, n11730, n11731, n11732, n11733, n11734, n11736, n11737, n11738,
    n11739, n11740, n11741, n11742, n11745, n11746, n11747, n11749, n11750,
    n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
    n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
    n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
    n11778, n11779, n11780, n11781, n11782, n11784, n11785, n11786, n11787,
    n11788, n11789, n11790, n11791, n11793, n11794, n11796, n11797, n11798,
    n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
    n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
    n11817, n11818, n11820, n11821, n11822, n11824, n11825, n11830, n11831,
    n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
    n11841, n11842, n11843, n11844, n11845, n11846, n11850, n11851, n11852,
    n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861,
    n11862, n11863, n11864, n11865, n11866, n11867, n11869, n11870, n11871,
    n11872, n11873, n11874, n11875, n11876, n11877, n11880, n11881, n11882,
    n11883, n11884, n11885, n11887, n11888, n11889, n11890, n11891, n11892,
    n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901,
    n11902, n11903, n11904, n11905, n11906, n11908, n11909, n11910, n11911,
    n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
    n11921, n11922, n11923, n11924, n11925, n11927, n11928, n11929, n11930,
    n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
    n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948,
    n11949, n11950, n11951, n11952, n11953, n11954, n11956, n11957, n11958,
    n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
    n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11979,
    n11980, n11981, n11982, n11985, n11986, n11987, n11988, n11989, n11990,
    n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
    n12000, n12001, n12002, n12003, n12004, n12005, n12007, n12008, n12009,
    n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
    n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12029,
    n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038,
    n12040, n12042, n12043, n12045, n12047, n12049, n12051, n12053, n12055,
    n12057, n12059, n12061, n12063, n12065, n12067, n12069, n12071, n12073,
    n12075, n12077, n12079, n12081, n12083, n12085, n12087, n12089, n12091,
    n12093, n12095, n12097, n12099, n12101, n12103, n12104, n12105, n12106,
    n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
    n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124,
    n12125, n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12135,
    n12136, n12137, n12138, n12139, n12141, n12142, n12143, n12144, n12145,
    n12147, n12148, n12149, n12150, n12151, n12152, n12154, n12155, n12156,
    n12157, n12158, n12159, n12161, n12162, n12163, n12164, n12165, n12166,
    n12168, n12169, n12170, n12171, n12173, n12174, n12175, n12176, n12177,
    n12178, n12180, n12181, n12182, n12183, n12184, n12186, n12187, n12188,
    n12189, n12190, n12191, n12193, n12194, n12195, n12196, n12197, n12198,
    n12200, n12201, n12202, n12203, n12204, n12206, n12207, n12208, n12209,
    n12210, n12212, n12213, n12214, n12215, n12216, n12217, n12219, n12220,
    n12221, n12222, n12223, n12224, n12225, n12227, n12228, n12229, n12230,
    n12231, n12233, n12234, n12235, n12236, n12237, n12239, n12240, n12241,
    n12242, n12243, n12245, n12246, n12247, n12248, n12250, n12251, n12252,
    n12253, n12254, n12255, n12257, n12258, n12259, n12260, n12261, n12262,
    n12263, n12265, n12266, n12267, n12268, n12269, n12271, n12272, n12273,
    n12274, n12275, n12276, n12277, n12279, n12280, n12281, n12282, n12283,
    n12284, n12285, n12287, n12288, n12289, n12290, n12291, n12292, n12294,
    n12295, n12296, n12297, n12298, n12299, n12301, n12302, n12303, n12304,
    n12305, n12306, n12308, n12309, n12310, n12311, n12312, n12313, n12315,
    n12316, n12317, n12318, n12319, n12321, n12322, n12323, n12324, n12326,
    n12327, n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
    n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
    n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
    n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
    n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371, n12372,
    n12373, n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381,
    n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390,
    n12391, n12392, n12393, n12400, n12401, n12402, n12403, n12404, n12405,
    n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414,
    n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
    n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
    n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
    n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,
    n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459,
    n12460, n12461, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
    n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
    n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
    n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
    n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507, n12508,
    n12509, n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517,
    n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526,
    n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
    n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
    n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
    n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
    n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
    n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579, n12580,
    n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589,
    n12590, n12591, n12592, n12593, n12594, n12596, n12597, n12598, n12599,
    n12600, n12601, n12602, n12603, n12605, n12606, n12607, n12608, n12609,
    n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618,
    n12619, n12620, n12622, n12623, n12624, n12625, n12626, n12627, n12628,
    n12629, n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637,
    n12638, n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
    n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
    n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12665, n12666,
    n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
    n12676, n12677, n12678, n12679, n12681, n12682, n12683, n12684, n12685,
    n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694,
    n12695, n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
    n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12714,
    n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723,
    n12724, n12725, n12726, n12727, n12728, n12730, n12731, n12732, n12733,
    n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742,
    n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12751, n12752,
    n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
    n12762, n12763, n12764, n12765, n12767, n12768, n12769, n12770, n12771,
    n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779, n12780,
    n12781, n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790,
    n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
    n12800, n12801, n12802, n12803, n12805, n12806, n12807, n12808, n12809,
    n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
    n12819, n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828,
    n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837,
    n12838, n12839, n12840, n12842, n12843, n12844, n12845, n12846, n12847,
    n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
    n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,
    n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12875, n12876,
    n12877, n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885,
    n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894,
    n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12903, n12904,
    n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
    n12914, n12915, n12916, n12918, n12919, n12920, n12921, n12922, n12923,
    n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931, n12932,
    n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942,
    n12943, n12944, n12945, n12947, n12949, n12951, n12953, n12955, n12957,
    n12959, n12961, n12963, n12965, n12967, n12969, n12971, n12973, n12975,
    n12977, n12979, n12981, n12983, n12985, n12987, n12989, n12991, n12993,
    n12995, n12997, n12999, n13001, n13003, n13005, n13007, n13008, n13010,
    n13013, n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021,
    n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030,
    n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
    n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
    n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
    n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
    n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075,
    n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084,
    n13085, n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093,
    n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102,
    n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
    n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
    n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
    n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
    n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147,
    n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155, n13156,
    n13157, n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165,
    n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174,
    n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
    n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
    n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
    n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
    n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219,
    n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227, n13228,
    n13229, n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237,
    n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246,
    n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
    n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
    n13265, n13266, n13267, n13269, n13270, n13271, n13272, n13273, n13274,
    n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
    n13284, n13285, n13286, n13287, n13290, n13291, n13294, n13295, n13297,
    n13298, n13300, n13301, n13302, n13303, n13305, n13306, n13307, n13309,
    n13311, n13312, n13314, n13317, n13318, n13319, n13320, n13321, n13322,
    n13324, n13325, n13326, n13327, n13329, n13330, n13331, n13332, n13333,
    n13334, n13335, n13337, n13338, n13340, n13343, n13344, n13345, n13346,
    n13348, n13349, n13350, n13351, n13352, n13353, n13355, n13356, n13357,
    n13358, n13359, n13360, n13361, n13363, n13365, n13366, n13367, n13368,
    n13370, n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13380,
    n13381, n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389,
    n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13401,
    n13402, n13405, n13406, n13407, n13408, n13409, n13410, n13411, n13412,
    n13413, n13415, n13416, n13419, n13420, n13421, n13422, n13423, n13424,
    n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
    n13434, n13435, n13436, n13437, n13439, n13440, n13441, n13442, n13443,
    n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451, n13452,
    n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461,
    n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470,
    n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
    n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
    n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
    n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
    n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515,
    n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524,
    n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533,
    n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542,
    n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
    n13553, n13554, n13555, n13557, n13558, n13559, n13560, n13561, n13562,
    n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571,
    n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580,
    n13581, n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589,
    n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598,
    n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
    n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
    n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
    n13626, n13627, n13630, n13631, n13632, n13633, n13634, n13635, n13637,
    n13638, n13639, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
    n13648, n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
    n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667,
    n13668, n13669, n13670, n13672, n13673, n13674, n13675, n13676, n13677,
    n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686,
    n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13696, n13697,
    n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
    n13707, n13708, n13709, n13710, n13712, n13713, n13714, n13715, n13717,
    n13718, n13719, n13720, n13721, n13722, n13723, n13725, n13727, n13728,
    n13729, n13730, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
    n13739, n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13749,
    n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758,
    n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
    n13769, n13770, n13771, n13772, n13774, n13775, n13776, n13777, n13778,
    n13779, n13780, n13781, n13783, n13785, n13786, n13787, n13788, n13789,
    n13790, n13791, n13792, n13794, n13795, n13797, n13798, n13799, n13800,
    n13801, n13802, n13803, n13805, n13806, n13808, n13809, n13810, n13811,
    n13812, n13813, n13814, n13816, n13817, n13818, n13819, n13820, n13821,
    n13822, n13823, n13824, n13825, n13826, n13827, n13829, n13830, n13831,
    n13832, n13833, n13834, n13835, n13836, n13837, n13839, n13840, n13841,
    n13842, n13843, n13844, n13845, n13846, n13847, n13849, n13850, n13851,
    n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859, n13860,
    n13861, n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869,
    n13870, n13871, n13872, n13873, n13874, n13875, n13877, n13879, n13880,
    n13881, n13882, n13883, n13884, n13885, n13886, n13888, n13889, n13890,
    n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899,
    n13901, n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13910,
    n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13919, n13920,
    n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
    n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939,
    n13941, n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949,
    n13950, n13951, n13952, n13953, n13955, n13956;
  INVX1   g00000(.A(P2_ADDR_REG_18__SCAN_IN), .Y(n1524));
  INVX1   g00001(.A(P2_ADDR_REG_17__SCAN_IN), .Y(n1525));
  INVX1   g00002(.A(P1_ADDR_REG_16__SCAN_IN), .Y(n1526));
  NOR2X1  g00003(.A(P3_ADDR_REG_16__SCAN_IN), .B(n1526), .Y(n1527));
  INVX1   g00004(.A(P1_ADDR_REG_15__SCAN_IN), .Y(n1528));
  NOR2X1  g00005(.A(P3_ADDR_REG_15__SCAN_IN), .B(n1528), .Y(n1529));
  INVX1   g00006(.A(P3_ADDR_REG_15__SCAN_IN), .Y(n1530));
  NOR2X1  g00007(.A(n1530), .B(P1_ADDR_REG_15__SCAN_IN), .Y(n1531));
  INVX1   g00008(.A(n1531), .Y(n1532));
  INVX1   g00009(.A(P1_ADDR_REG_14__SCAN_IN), .Y(n1533));
  NOR2X1  g00010(.A(P3_ADDR_REG_14__SCAN_IN), .B(n1533), .Y(n1534));
  INVX1   g00011(.A(n1534), .Y(n1535));
  INVX1   g00012(.A(P3_ADDR_REG_14__SCAN_IN), .Y(n1536));
  NOR2X1  g00013(.A(n1536), .B(P1_ADDR_REG_14__SCAN_IN), .Y(n1537));
  INVX1   g00014(.A(P1_ADDR_REG_13__SCAN_IN), .Y(n1538));
  NOR2X1  g00015(.A(P3_ADDR_REG_13__SCAN_IN), .B(n1538), .Y(n1539));
  INVX1   g00016(.A(P3_ADDR_REG_13__SCAN_IN), .Y(n1540));
  NOR2X1  g00017(.A(n1540), .B(P1_ADDR_REG_13__SCAN_IN), .Y(n1541));
  INVX1   g00018(.A(n1541), .Y(n1542));
  INVX1   g00019(.A(P1_ADDR_REG_12__SCAN_IN), .Y(n1543));
  INVX1   g00020(.A(P3_ADDR_REG_12__SCAN_IN), .Y(n1544));
  INVX1   g00021(.A(P1_ADDR_REG_11__SCAN_IN), .Y(n1545));
  NOR2X1  g00022(.A(P3_ADDR_REG_11__SCAN_IN), .B(n1545), .Y(n1546));
  INVX1   g00023(.A(P1_ADDR_REG_10__SCAN_IN), .Y(n1547));
  NOR2X1  g00024(.A(P3_ADDR_REG_10__SCAN_IN), .B(n1547), .Y(n1548));
  NAND2X1 g00025(.A(P3_ADDR_REG_10__SCAN_IN), .B(n1547), .Y(n1549));
  INVX1   g00026(.A(P1_ADDR_REG_9__SCAN_IN), .Y(n1550));
  NOR2X1  g00027(.A(n1550), .B(P3_ADDR_REG_9__SCAN_IN), .Y(n1551));
  INVX1   g00028(.A(P3_ADDR_REG_9__SCAN_IN), .Y(n1552));
  NOR2X1  g00029(.A(P1_ADDR_REG_9__SCAN_IN), .B(n1552), .Y(n1553));
  INVX1   g00030(.A(n1553), .Y(n1554));
  INVX1   g00031(.A(P1_ADDR_REG_8__SCAN_IN), .Y(n1555));
  INVX1   g00032(.A(P3_ADDR_REG_8__SCAN_IN), .Y(n1556));
  INVX1   g00033(.A(P1_ADDR_REG_7__SCAN_IN), .Y(n1557));
  NOR2X1  g00034(.A(n1557), .B(P3_ADDR_REG_7__SCAN_IN), .Y(n1558));
  INVX1   g00035(.A(P3_ADDR_REG_6__SCAN_IN), .Y(n1559));
  INVX1   g00036(.A(P1_ADDR_REG_6__SCAN_IN), .Y(n1560));
  INVX1   g00037(.A(P3_ADDR_REG_5__SCAN_IN), .Y(n1561));
  NOR2X1  g00038(.A(P1_ADDR_REG_5__SCAN_IN), .B(n1561), .Y(n1562));
  INVX1   g00039(.A(P1_ADDR_REG_4__SCAN_IN), .Y(n1563));
  NOR2X1  g00040(.A(n1563), .B(P3_ADDR_REG_4__SCAN_IN), .Y(n1564));
  INVX1   g00041(.A(n1564), .Y(n1565));
  INVX1   g00042(.A(P3_ADDR_REG_4__SCAN_IN), .Y(n1566));
  NOR2X1  g00043(.A(P1_ADDR_REG_4__SCAN_IN), .B(n1566), .Y(n1567));
  INVX1   g00044(.A(P1_ADDR_REG_3__SCAN_IN), .Y(n1568));
  NOR2X1  g00045(.A(n1568), .B(P3_ADDR_REG_3__SCAN_IN), .Y(n1569));
  INVX1   g00046(.A(P3_ADDR_REG_3__SCAN_IN), .Y(n1570));
  NOR2X1  g00047(.A(P1_ADDR_REG_3__SCAN_IN), .B(n1570), .Y(n1571));
  INVX1   g00048(.A(n1571), .Y(n1572));
  INVX1   g00049(.A(P3_ADDR_REG_2__SCAN_IN), .Y(n1573));
  NAND2X1 g00050(.A(P1_ADDR_REG_2__SCAN_IN), .B(n1573), .Y(n1574));
  NOR2X1  g00051(.A(P1_ADDR_REG_2__SCAN_IN), .B(n1573), .Y(n1575));
  INVX1   g00052(.A(P1_ADDR_REG_0__SCAN_IN), .Y(n1576));
  NAND2X1 g00053(.A(n1576), .B(P3_ADDR_REG_0__SCAN_IN), .Y(n1577));
  INVX1   g00054(.A(P1_ADDR_REG_1__SCAN_IN), .Y(n1578));
  INVX1   g00055(.A(P3_ADDR_REG_0__SCAN_IN), .Y(n1579));
  NOR2X1  g00056(.A(P1_ADDR_REG_0__SCAN_IN), .B(n1579), .Y(n1580));
  AOI21X1 g00057(.A0(n1580), .A1(n1578), .B0(P3_ADDR_REG_1__SCAN_IN), .Y(n1581));
  AOI21X1 g00058(.A0(n1577), .A1(P1_ADDR_REG_1__SCAN_IN), .B0(n1581), .Y(n1582));
  OAI21X1 g00059(.A0(n1582), .A1(n1575), .B0(n1574), .Y(n1583));
  AOI21X1 g00060(.A0(n1583), .A1(n1572), .B0(n1569), .Y(n1584));
  OAI21X1 g00061(.A0(n1584), .A1(n1567), .B0(n1565), .Y(n1585));
  INVX1   g00062(.A(n1585), .Y(n1586));
  NOR2X1  g00063(.A(n1586), .B(n1562), .Y(n1587));
  AOI21X1 g00064(.A0(P1_ADDR_REG_5__SCAN_IN), .A1(n1561), .B0(n1587), .Y(n1588));
  AOI21X1 g00065(.A0(n1560), .A1(P3_ADDR_REG_6__SCAN_IN), .B0(n1588), .Y(n1589));
  AOI21X1 g00066(.A0(P1_ADDR_REG_6__SCAN_IN), .A1(n1559), .B0(n1589), .Y(n1590));
  AOI21X1 g00067(.A0(n1557), .A1(P3_ADDR_REG_7__SCAN_IN), .B0(n1590), .Y(n1591));
  OAI22X1 g00068(.A0(n1558), .A1(n1591), .B0(P1_ADDR_REG_8__SCAN_IN), .B1(n1556), .Y(n1592));
  OAI21X1 g00069(.A0(n1555), .A1(P3_ADDR_REG_8__SCAN_IN), .B0(n1592), .Y(n1593));
  AOI21X1 g00070(.A0(n1593), .A1(n1554), .B0(n1551), .Y(n1594));
  INVX1   g00071(.A(n1594), .Y(n1595));
  AOI21X1 g00072(.A0(n1595), .A1(n1549), .B0(n1548), .Y(n1596));
  AOI21X1 g00073(.A0(P3_ADDR_REG_11__SCAN_IN), .A1(n1545), .B0(n1596), .Y(n1597));
  OAI22X1 g00074(.A0(n1546), .A1(n1597), .B0(n1544), .B1(P1_ADDR_REG_12__SCAN_IN), .Y(n1598));
  OAI21X1 g00075(.A0(P3_ADDR_REG_12__SCAN_IN), .A1(n1543), .B0(n1598), .Y(n1599));
  AOI21X1 g00076(.A0(n1599), .A1(n1542), .B0(n1539), .Y(n1600));
  OAI21X1 g00077(.A0(n1600), .A1(n1537), .B0(n1535), .Y(n1601));
  AOI21X1 g00078(.A0(n1601), .A1(n1532), .B0(n1529), .Y(n1602));
  AOI21X1 g00079(.A0(P3_ADDR_REG_16__SCAN_IN), .A1(n1526), .B0(n1602), .Y(n1603));
  NOR2X1  g00080(.A(n1603), .B(n1527), .Y(n1604));
  INVX1   g00081(.A(P1_ADDR_REG_17__SCAN_IN), .Y(n1605));
  XOR2X1  g00082(.A(P3_ADDR_REG_17__SCAN_IN), .B(n1605), .Y(n1606));
  XOR2X1  g00083(.A(n1606), .B(n1604), .Y(n1607));
  NOR2X1  g00084(.A(n1607), .B(n1525), .Y(n1608));
  NAND2X1 g00085(.A(n1607), .B(n1525), .Y(n1609));
  INVX1   g00086(.A(P2_ADDR_REG_16__SCAN_IN), .Y(n1610));
  XOR2X1  g00087(.A(P3_ADDR_REG_16__SCAN_IN), .B(n1526), .Y(n1611));
  XOR2X1  g00088(.A(n1611), .B(n1602), .Y(n1612));
  NOR2X1  g00089(.A(n1612), .B(n1610), .Y(n1613));
  INVX1   g00090(.A(n1613), .Y(n1614));
  NAND2X1 g00091(.A(n1612), .B(n1610), .Y(n1615));
  INVX1   g00092(.A(n1615), .Y(n1616));
  INVX1   g00093(.A(P2_ADDR_REG_15__SCAN_IN), .Y(n1617));
  INVX1   g00094(.A(P2_ADDR_REG_12__SCAN_IN), .Y(n1618));
  NOR2X1  g00095(.A(n1597), .B(n1546), .Y(n1619));
  XOR2X1  g00096(.A(P3_ADDR_REG_12__SCAN_IN), .B(n1543), .Y(n1620));
  XOR2X1  g00097(.A(n1620), .B(n1619), .Y(n1621));
  NOR2X1  g00098(.A(n1621), .B(n1618), .Y(n1622));
  XOR2X1  g00099(.A(P3_ADDR_REG_11__SCAN_IN), .B(n1545), .Y(n1623));
  XOR2X1  g00100(.A(n1623), .B(n1596), .Y(n1624));
  INVX1   g00101(.A(n1624), .Y(n1625));
  NAND2X1 g00102(.A(n1625), .B(P2_ADDR_REG_11__SCAN_IN), .Y(n1626));
  XOR2X1  g00103(.A(P1_ADDR_REG_9__SCAN_IN), .B(n1552), .Y(n1627));
  XOR2X1  g00104(.A(n1627), .B(n1593), .Y(n1628));
  NAND2X1 g00105(.A(n1628), .B(P2_ADDR_REG_9__SCAN_IN), .Y(n1629));
  NOR2X1  g00106(.A(n1628), .B(P2_ADDR_REG_9__SCAN_IN), .Y(n1630));
  INVX1   g00107(.A(P2_ADDR_REG_8__SCAN_IN), .Y(n1631));
  INVX1   g00108(.A(P2_ADDR_REG_7__SCAN_IN), .Y(n1632));
  INVX1   g00109(.A(P3_ADDR_REG_7__SCAN_IN), .Y(n1633));
  XOR2X1  g00110(.A(P1_ADDR_REG_7__SCAN_IN), .B(n1633), .Y(n1634));
  XOR2X1  g00111(.A(n1634), .B(n1590), .Y(n1635));
  NOR2X1  g00112(.A(n1635), .B(n1632), .Y(n1636));
  INVX1   g00113(.A(P2_ADDR_REG_6__SCAN_IN), .Y(n1637));
  XOR2X1  g00114(.A(P1_ADDR_REG_6__SCAN_IN), .B(n1559), .Y(n1638));
  XOR2X1  g00115(.A(n1638), .B(n1588), .Y(n1639));
  NOR2X1  g00116(.A(n1639), .B(n1637), .Y(n1640));
  INVX1   g00117(.A(P2_ADDR_REG_5__SCAN_IN), .Y(n1641));
  INVX1   g00118(.A(P2_ADDR_REG_4__SCAN_IN), .Y(n1642));
  XOR2X1  g00119(.A(P1_ADDR_REG_4__SCAN_IN), .B(n1566), .Y(n1643));
  XOR2X1  g00120(.A(n1643), .B(n1584), .Y(n1644));
  NOR2X1  g00121(.A(n1644), .B(n1642), .Y(n1645));
  INVX1   g00122(.A(P2_ADDR_REG_3__SCAN_IN), .Y(n1646));
  INVX1   g00123(.A(P2_ADDR_REG_2__SCAN_IN), .Y(n1647));
  XOR2X1  g00124(.A(P1_ADDR_REG_2__SCAN_IN), .B(n1573), .Y(n1648));
  XOR2X1  g00125(.A(n1648), .B(n1582), .Y(n1649));
  NOR2X1  g00126(.A(n1649), .B(n1647), .Y(n1650));
  XOR2X1  g00127(.A(n1578), .B(P3_ADDR_REG_1__SCAN_IN), .Y(n1651));
  XOR2X1  g00128(.A(n1651), .B(n1577), .Y(n1652));
  XOR2X1  g00129(.A(P1_ADDR_REG_0__SCAN_IN), .B(P3_ADDR_REG_0__SCAN_IN), .Y(n1653));
  NAND2X1 g00130(.A(n1653), .B(P2_ADDR_REG_0__SCAN_IN), .Y(n1654));
  INVX1   g00131(.A(n1654), .Y(n1655));
  INVX1   g00132(.A(P2_ADDR_REG_1__SCAN_IN), .Y(n1656));
  XOR2X1  g00133(.A(n1651), .B(n1580), .Y(n1657));
  AOI21X1 g00134(.A0(n1654), .A1(n1657), .B0(n1656), .Y(n1658));
  AOI21X1 g00135(.A0(n1655), .A1(n1652), .B0(n1658), .Y(n1659));
  AOI21X1 g00136(.A0(n1649), .A1(n1647), .B0(n1659), .Y(n1660));
  NOR2X1  g00137(.A(n1660), .B(n1650), .Y(n1661));
  NOR2X1  g00138(.A(n1661), .B(n1646), .Y(n1662));
  XOR2X1  g00139(.A(P1_ADDR_REG_3__SCAN_IN), .B(n1570), .Y(n1663));
  XOR2X1  g00140(.A(n1663), .B(n1583), .Y(n1664));
  NAND2X1 g00141(.A(n1661), .B(n1646), .Y(n1665));
  AOI21X1 g00142(.A0(n1665), .A1(n1664), .B0(n1662), .Y(n1666));
  AOI21X1 g00143(.A0(n1644), .A1(n1642), .B0(n1666), .Y(n1667));
  NOR2X1  g00144(.A(n1667), .B(n1645), .Y(n1668));
  NOR2X1  g00145(.A(n1668), .B(n1641), .Y(n1669));
  XOR2X1  g00146(.A(P1_ADDR_REG_5__SCAN_IN), .B(n1561), .Y(n1670));
  XOR2X1  g00147(.A(n1670), .B(n1585), .Y(n1671));
  NAND2X1 g00148(.A(n1668), .B(n1641), .Y(n1672));
  AOI21X1 g00149(.A0(n1672), .A1(n1671), .B0(n1669), .Y(n1673));
  AOI21X1 g00150(.A0(n1639), .A1(n1637), .B0(n1673), .Y(n1674));
  NOR2X1  g00151(.A(n1674), .B(n1640), .Y(n1675));
  AOI21X1 g00152(.A0(n1635), .A1(n1632), .B0(n1675), .Y(n1676));
  NOR2X1  g00153(.A(n1676), .B(n1636), .Y(n1677));
  NOR2X1  g00154(.A(n1677), .B(n1631), .Y(n1678));
  AOI21X1 g00155(.A0(P1_ADDR_REG_7__SCAN_IN), .A1(n1633), .B0(n1591), .Y(n1679));
  XOR2X1  g00156(.A(P1_ADDR_REG_8__SCAN_IN), .B(P3_ADDR_REG_8__SCAN_IN), .Y(n1680));
  XOR2X1  g00157(.A(n1680), .B(n1679), .Y(n1681));
  NAND2X1 g00158(.A(n1677), .B(n1631), .Y(n1682));
  AOI21X1 g00159(.A0(n1682), .A1(n1681), .B0(n1678), .Y(n1683));
  OAI21X1 g00160(.A0(n1683), .A1(n1630), .B0(n1629), .Y(n1684));
  NAND2X1 g00161(.A(n1684), .B(P2_ADDR_REG_10__SCAN_IN), .Y(n1685));
  XOR2X1  g00162(.A(P3_ADDR_REG_10__SCAN_IN), .B(n1547), .Y(n1686));
  XOR2X1  g00163(.A(n1686), .B(n1594), .Y(n1687));
  NOR2X1  g00164(.A(n1684), .B(P2_ADDR_REG_10__SCAN_IN), .Y(n1688));
  OAI21X1 g00165(.A0(n1688), .A1(n1687), .B0(n1685), .Y(n1689));
  OAI21X1 g00166(.A0(n1625), .A1(P2_ADDR_REG_11__SCAN_IN), .B0(n1689), .Y(n1690));
  AOI22X1 g00167(.A0(n1626), .A1(n1690), .B0(n1621), .B1(n1618), .Y(n1691));
  OAI21X1 g00168(.A0(n1691), .A1(n1622), .B0(P2_ADDR_REG_13__SCAN_IN), .Y(n1692));
  XOR2X1  g00169(.A(P3_ADDR_REG_13__SCAN_IN), .B(n1538), .Y(n1693));
  XOR2X1  g00170(.A(n1693), .B(n1599), .Y(n1694));
  INVX1   g00171(.A(n1694), .Y(n1695));
  NOR3X1  g00172(.A(n1691), .B(n1622), .C(P2_ADDR_REG_13__SCAN_IN), .Y(n1696));
  OAI21X1 g00173(.A0(n1696), .A1(n1695), .B0(n1692), .Y(n1697));
  NAND2X1 g00174(.A(n1697), .B(P2_ADDR_REG_14__SCAN_IN), .Y(n1698));
  XOR2X1  g00175(.A(P3_ADDR_REG_14__SCAN_IN), .B(n1533), .Y(n1699));
  XOR2X1  g00176(.A(n1699), .B(n1600), .Y(n1700));
  INVX1   g00177(.A(n1700), .Y(n1701));
  OAI21X1 g00178(.A0(n1697), .A1(P2_ADDR_REG_14__SCAN_IN), .B0(n1701), .Y(n1702));
  AOI21X1 g00179(.A0(n1702), .A1(n1698), .B0(n1617), .Y(n1703));
  XOR2X1  g00180(.A(P3_ADDR_REG_15__SCAN_IN), .B(n1528), .Y(n1704));
  XOR2X1  g00181(.A(n1704), .B(n1601), .Y(n1705));
  NAND3X1 g00182(.A(n1702), .B(n1698), .C(n1617), .Y(n1706));
  AOI21X1 g00183(.A0(n1706), .A1(n1705), .B0(n1703), .Y(n1707));
  OAI21X1 g00184(.A0(n1707), .A1(n1616), .B0(n1614), .Y(n1708));
  AOI21X1 g00185(.A0(n1708), .A1(n1609), .B0(n1608), .Y(n1709));
  INVX1   g00186(.A(P3_ADDR_REG_17__SCAN_IN), .Y(n1710));
  AOI21X1 g00187(.A0(P3_ADDR_REG_17__SCAN_IN), .A1(n1605), .B0(n1604), .Y(n1711));
  AOI21X1 g00188(.A0(n1710), .A1(P1_ADDR_REG_17__SCAN_IN), .B0(n1711), .Y(n1712));
  INVX1   g00189(.A(P1_ADDR_REG_18__SCAN_IN), .Y(n1713));
  XOR2X1  g00190(.A(P3_ADDR_REG_18__SCAN_IN), .B(n1713), .Y(n1714));
  XOR2X1  g00191(.A(n1714), .B(n1712), .Y(n1715));
  OAI21X1 g00192(.A0(n1709), .A1(n1524), .B0(n1715), .Y(n1716));
  OAI21X1 g00193(.A0(P3_ADDR_REG_18__SCAN_IN), .A1(n1713), .B0(n1712), .Y(n1717));
  INVX1   g00194(.A(P1_ADDR_REG_19__SCAN_IN), .Y(n1718));
  XOR2X1  g00195(.A(P3_ADDR_REG_19__SCAN_IN), .B(n1718), .Y(n1719));
  AOI21X1 g00196(.A0(P3_ADDR_REG_18__SCAN_IN), .A1(n1713), .B0(n1719), .Y(n1720));
  AOI21X1 g00197(.A0(P3_ADDR_REG_18__SCAN_IN), .A1(n1713), .B0(n1712), .Y(n1721));
  OAI21X1 g00198(.A0(P3_ADDR_REG_18__SCAN_IN), .A1(n1713), .B0(n1719), .Y(n1722));
  NOR2X1  g00199(.A(n1722), .B(n1721), .Y(n1723));
  AOI21X1 g00200(.A0(n1720), .A1(n1717), .B0(n1723), .Y(n1724));
  XOR2X1  g00201(.A(n1724), .B(P2_ADDR_REG_19__SCAN_IN), .Y(n1725));
  AOI21X1 g00202(.A0(n1709), .A1(n1524), .B0(n1725), .Y(n1726));
  NOR2X1  g00203(.A(n1709), .B(n1524), .Y(n1727));
  INVX1   g00204(.A(P2_ADDR_REG_19__SCAN_IN), .Y(n1728));
  XOR2X1  g00205(.A(n1724), .B(n1728), .Y(n1729));
  AOI21X1 g00206(.A0(n1709), .A1(n1524), .B0(n1715), .Y(n1730));
  NOR3X1  g00207(.A(n1730), .B(n1729), .C(n1727), .Y(n1731));
  AOI21X1 g00208(.A0(n1726), .A1(n1716), .B0(n1731), .Y(SUB_1596_U4));
  XOR2X1  g00209(.A(n1709), .B(P2_ADDR_REG_18__SCAN_IN), .Y(n1733));
  XOR2X1  g00210(.A(n1733), .B(n1715), .Y(SUB_1596_U62));
  XOR2X1  g00211(.A(n1607), .B(n1525), .Y(n1735));
  XOR2X1  g00212(.A(n1735), .B(n1708), .Y(SUB_1596_U63));
  XOR2X1  g00213(.A(n1612), .B(P2_ADDR_REG_16__SCAN_IN), .Y(n1737));
  XOR2X1  g00214(.A(n1737), .B(n1707), .Y(SUB_1596_U64));
  NAND2X1 g00215(.A(n1702), .B(n1698), .Y(n1739));
  XOR2X1  g00216(.A(n1739), .B(P2_ADDR_REG_15__SCAN_IN), .Y(n1740));
  XOR2X1  g00217(.A(n1740), .B(n1705), .Y(SUB_1596_U65));
  XOR2X1  g00218(.A(n1697), .B(P2_ADDR_REG_14__SCAN_IN), .Y(n1742));
  XOR2X1  g00219(.A(n1742), .B(n1701), .Y(SUB_1596_U66));
  NOR2X1  g00220(.A(n1691), .B(n1622), .Y(n1744));
  XOR2X1  g00221(.A(n1744), .B(P2_ADDR_REG_13__SCAN_IN), .Y(n1745));
  XOR2X1  g00222(.A(n1745), .B(n1695), .Y(SUB_1596_U67));
  NAND2X1 g00223(.A(n1690), .B(n1626), .Y(n1747));
  XOR2X1  g00224(.A(n1621), .B(n1618), .Y(n1748));
  XOR2X1  g00225(.A(n1748), .B(n1747), .Y(SUB_1596_U68));
  INVX1   g00226(.A(P2_ADDR_REG_11__SCAN_IN), .Y(n1750));
  XOR2X1  g00227(.A(n1624), .B(n1750), .Y(n1751));
  XOR2X1  g00228(.A(n1751), .B(n1689), .Y(SUB_1596_U69));
  INVX1   g00229(.A(P2_ADDR_REG_10__SCAN_IN), .Y(n1753));
  XOR2X1  g00230(.A(n1684), .B(n1753), .Y(n1754));
  XOR2X1  g00231(.A(n1754), .B(n1687), .Y(SUB_1596_U70));
  INVX1   g00232(.A(P2_ADDR_REG_9__SCAN_IN), .Y(n1756));
  XOR2X1  g00233(.A(n1628), .B(n1756), .Y(n1757));
  XOR2X1  g00234(.A(n1757), .B(n1683), .Y(SUB_1596_U54));
  XOR2X1  g00235(.A(n1677), .B(n1631), .Y(n1759));
  XOR2X1  g00236(.A(n1759), .B(n1681), .Y(SUB_1596_U55));
  XOR2X1  g00237(.A(n1635), .B(P2_ADDR_REG_7__SCAN_IN), .Y(n1761));
  XOR2X1  g00238(.A(n1761), .B(n1675), .Y(SUB_1596_U56));
  XOR2X1  g00239(.A(n1639), .B(P2_ADDR_REG_6__SCAN_IN), .Y(n1763));
  XOR2X1  g00240(.A(n1763), .B(n1673), .Y(SUB_1596_U57));
  XOR2X1  g00241(.A(n1668), .B(n1641), .Y(n1765));
  XOR2X1  g00242(.A(n1765), .B(n1671), .Y(SUB_1596_U58));
  XOR2X1  g00243(.A(n1644), .B(P2_ADDR_REG_4__SCAN_IN), .Y(n1767));
  XOR2X1  g00244(.A(n1767), .B(n1666), .Y(SUB_1596_U59));
  XOR2X1  g00245(.A(n1661), .B(n1646), .Y(n1769));
  XOR2X1  g00246(.A(n1769), .B(n1664), .Y(SUB_1596_U60));
  XOR2X1  g00247(.A(n1649), .B(P2_ADDR_REG_2__SCAN_IN), .Y(n1771));
  XOR2X1  g00248(.A(n1771), .B(n1659), .Y(SUB_1596_U61));
  NAND3X1 g00249(.A(n1655), .B(n1652), .C(P2_ADDR_REG_1__SCAN_IN), .Y(n1773));
  XOR2X1  g00250(.A(n1654), .B(n1656), .Y(n1774));
  NAND2X1 g00251(.A(n1774), .B(n1657), .Y(n1775));
  NAND3X1 g00252(.A(n1654), .B(n1652), .C(n1656), .Y(n1776));
  NAND3X1 g00253(.A(n1776), .B(n1775), .C(n1773), .Y(SUB_1596_U5));
  XOR2X1  g00254(.A(n1653), .B(P2_ADDR_REG_0__SCAN_IN), .Y(SUB_1596_U53));
  INVX1   g00255(.A(P3_RD_REG_SCAN_IN), .Y(n1779));
  XOR2X1  g00256(.A(P2_RD_REG_SCAN_IN), .B(P1_RD_REG_SCAN_IN), .Y(n1780));
  NAND2X1 g00257(.A(n1780), .B(n1779), .Y(U29));
  INVX1   g00258(.A(P3_WR_REG_SCAN_IN), .Y(n1782));
  XOR2X1  g00259(.A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .Y(n1783));
  NAND2X1 g00260(.A(n1783), .B(n1782), .Y(U28));
  NOR2X1  g00261(.A(P2_ADDR_REG_19__SCAN_IN), .B(P1_RD_REG_SCAN_IN), .Y(n1785));
  NAND3X1 g00262(.A(n1785), .B(P3_ADDR_REG_19__SCAN_IN), .C(n1718), .Y(n1786));
  INVX1   g00263(.A(P2_RD_REG_SCAN_IN), .Y(n1787));
  INVX1   g00264(.A(P3_ADDR_REG_19__SCAN_IN), .Y(n1788));
  NAND4X1 g00265(.A(n1787), .B(P2_ADDR_REG_19__SCAN_IN), .C(P1_ADDR_REG_19__SCAN_IN), .D(n1788), .Y(n1789));
  NAND2X1 g00266(.A(n1789), .B(n1786), .Y(n1790));
  INVX1   g00267(.A(P2_DATAO_REG_0__SCAN_IN), .Y(n1791));
  NOR4X1  g00268(.A(P2_ADDR_REG_19__SCAN_IN), .B(P1_RD_REG_SCAN_IN), .C(P1_ADDR_REG_19__SCAN_IN), .D(n1788), .Y(n1792));
  NOR4X1  g00269(.A(P2_RD_REG_SCAN_IN), .B(n1728), .C(n1718), .D(P3_ADDR_REG_19__SCAN_IN), .Y(n1793));
  NOR3X1  g00270(.A(n1793), .B(n1792), .C(n1791), .Y(n1794));
  INVX1   g00271(.A(SI_0_), .Y(n1795));
  INVX1   g00272(.A(P1_DATAO_REG_0__SCAN_IN), .Y(n1796));
  NOR3X1  g00273(.A(n1793), .B(n1792), .C(n1796), .Y(n1797));
  AOI21X1 g00274(.A0(n1789), .A1(n1786), .B0(n1791), .Y(n1798));
  NOR2X1  g00275(.A(n1798), .B(n1797), .Y(n1799));
  XOR2X1  g00276(.A(n1799), .B(n1795), .Y(n1800));
  AOI21X1 g00277(.A0(n1800), .A1(n1790), .B0(n1794), .Y(n1801));
  INVX1   g00278(.A(P1_STATE_REG_SCAN_IN), .Y(P1_U3086));
  NOR2X1  g00279(.A(P1_U3086), .B(P1_IR_REG_31__SCAN_IN), .Y(n1803));
  OAI21X1 g00280(.A0(n1803), .A1(P1_STATE_REG_SCAN_IN), .B0(P1_IR_REG_0__SCAN_IN), .Y(n1804));
  OAI21X1 g00281(.A0(n1801), .A1(P1_STATE_REG_SCAN_IN), .B0(n1804), .Y(P1_U3355));
  INVX1   g00282(.A(P2_DATAO_REG_1__SCAN_IN), .Y(n1806));
  NOR3X1  g00283(.A(n1793), .B(n1792), .C(n1806), .Y(n1807));
  INVX1   g00284(.A(P1_DATAO_REG_1__SCAN_IN), .Y(n1808));
  NOR3X1  g00285(.A(n1793), .B(n1792), .C(n1808), .Y(n1809));
  AOI21X1 g00286(.A0(n1789), .A1(n1786), .B0(n1806), .Y(n1810));
  NOR2X1  g00287(.A(n1810), .B(n1809), .Y(n1811));
  NAND3X1 g00288(.A(n1789), .B(n1786), .C(P1_DATAO_REG_0__SCAN_IN), .Y(n1812));
  OAI21X1 g00289(.A0(n1793), .A1(n1792), .B0(P2_DATAO_REG_0__SCAN_IN), .Y(n1813));
  AOI21X1 g00290(.A0(n1813), .A1(n1812), .B0(n1795), .Y(n1814));
  XOR2X1  g00291(.A(n1814), .B(n1811), .Y(n1815));
  NAND3X1 g00292(.A(n1789), .B(n1786), .C(P1_DATAO_REG_1__SCAN_IN), .Y(n1816));
  OAI21X1 g00293(.A0(n1793), .A1(n1792), .B0(P2_DATAO_REG_1__SCAN_IN), .Y(n1817));
  NAND2X1 g00294(.A(n1817), .B(n1816), .Y(n1818));
  OAI21X1 g00295(.A0(n1798), .A1(n1797), .B0(SI_0_), .Y(n1819));
  NAND2X1 g00296(.A(SI_0_), .B(SI_1_), .Y(n1820));
  AOI21X1 g00297(.A0(n1813), .A1(n1812), .B0(n1820), .Y(n1821));
  INVX1   g00298(.A(SI_1_), .Y(n1822));
  NOR3X1  g00299(.A(n1810), .B(n1809), .C(n1822), .Y(n1823));
  AOI22X1 g00300(.A0(n1821), .A1(n1818), .B0(n1819), .B1(n1823), .Y(n1824));
  OAI21X1 g00301(.A0(n1815), .A1(SI_1_), .B0(n1824), .Y(n1825));
  AOI21X1 g00302(.A0(n1825), .A1(n1790), .B0(n1807), .Y(n1826));
  INVX1   g00303(.A(P1_IR_REG_31__SCAN_IN), .Y(n1827));
  NOR2X1  g00304(.A(P1_U3086), .B(n1827), .Y(n1828));
  XOR2X1  g00305(.A(P1_IR_REG_1__SCAN_IN), .B(P1_IR_REG_0__SCAN_IN), .Y(n1829));
  AOI22X1 g00306(.A0(n1828), .A1(n1829), .B0(n1803), .B1(P1_IR_REG_1__SCAN_IN), .Y(n1830));
  OAI21X1 g00307(.A0(n1826), .A1(P1_STATE_REG_SCAN_IN), .B0(n1830), .Y(P1_U3354));
  INVX1   g00308(.A(P2_DATAO_REG_2__SCAN_IN), .Y(n1832));
  NOR3X1  g00309(.A(n1793), .B(n1792), .C(n1832), .Y(n1833));
  NOR2X1  g00310(.A(n1819), .B(n1811), .Y(n1834));
  OAI22X1 g00311(.A0(n1811), .A1(n1822), .B0(n1799), .B1(n1820), .Y(n1835));
  NOR2X1  g00312(.A(n1835), .B(n1834), .Y(n1836));
  NOR2X1  g00313(.A(n1793), .B(n1792), .Y(n1837));
  AOI21X1 g00314(.A0(n1789), .A1(n1786), .B0(n1832), .Y(n1838));
  AOI21X1 g00315(.A0(n1837), .A1(P1_DATAO_REG_2__SCAN_IN), .B0(n1838), .Y(n1839));
  XOR2X1  g00316(.A(n1839), .B(SI_2_), .Y(n1840));
  XOR2X1  g00317(.A(n1840), .B(n1836), .Y(n1841));
  AOI21X1 g00318(.A0(n1841), .A1(n1790), .B0(n1833), .Y(n1842));
  INVX1   g00319(.A(P1_IR_REG_2__SCAN_IN), .Y(n1843));
  NOR2X1  g00320(.A(P1_IR_REG_1__SCAN_IN), .B(P1_IR_REG_0__SCAN_IN), .Y(n1844));
  XOR2X1  g00321(.A(n1844), .B(n1843), .Y(n1845));
  AOI22X1 g00322(.A0(n1828), .A1(n1845), .B0(n1803), .B1(P1_IR_REG_2__SCAN_IN), .Y(n1846));
  OAI21X1 g00323(.A0(n1842), .A1(P1_STATE_REG_SCAN_IN), .B0(n1846), .Y(P1_U3353));
  INVX1   g00324(.A(P2_DATAO_REG_3__SCAN_IN), .Y(n1848));
  NOR3X1  g00325(.A(n1793), .B(n1792), .C(n1848), .Y(n1849));
  INVX1   g00326(.A(SI_2_), .Y(n1850));
  NAND2X1 g00327(.A(n1839), .B(n1850), .Y(n1851));
  NAND2X1 g00328(.A(n1851), .B(n1834), .Y(n1852));
  NAND3X1 g00329(.A(n1851), .B(n1814), .C(SI_1_), .Y(n1853));
  INVX1   g00330(.A(P1_DATAO_REG_2__SCAN_IN), .Y(n1854));
  OAI21X1 g00331(.A0(n1793), .A1(n1792), .B0(P2_DATAO_REG_2__SCAN_IN), .Y(n1855));
  OAI21X1 g00332(.A0(n1790), .A1(n1854), .B0(n1855), .Y(n1856));
  NAND2X1 g00333(.A(n1856), .B(SI_2_), .Y(n1857));
  NAND3X1 g00334(.A(n1851), .B(n1818), .C(SI_1_), .Y(n1858));
  NAND4X1 g00335(.A(n1857), .B(n1853), .C(n1852), .D(n1858), .Y(n1859));
  AOI21X1 g00336(.A0(n1789), .A1(n1786), .B0(n1848), .Y(n1860));
  AOI21X1 g00337(.A0(n1837), .A1(P1_DATAO_REG_3__SCAN_IN), .B0(n1860), .Y(n1861));
  XOR2X1  g00338(.A(n1861), .B(SI_3_), .Y(n1862));
  INVX1   g00339(.A(n1862), .Y(n1863));
  XOR2X1  g00340(.A(n1863), .B(n1859), .Y(n1864));
  AOI21X1 g00341(.A0(n1864), .A1(n1790), .B0(n1849), .Y(n1865));
  INVX1   g00342(.A(P1_IR_REG_3__SCAN_IN), .Y(n1866));
  NOR3X1  g00343(.A(P1_IR_REG_2__SCAN_IN), .B(P1_IR_REG_1__SCAN_IN), .C(P1_IR_REG_0__SCAN_IN), .Y(n1867));
  XOR2X1  g00344(.A(n1867), .B(n1866), .Y(n1868));
  AOI22X1 g00345(.A0(n1828), .A1(n1868), .B0(n1803), .B1(P1_IR_REG_3__SCAN_IN), .Y(n1869));
  OAI21X1 g00346(.A0(n1865), .A1(P1_STATE_REG_SCAN_IN), .B0(n1869), .Y(P1_U3352));
  INVX1   g00347(.A(P2_DATAO_REG_4__SCAN_IN), .Y(n1871));
  NOR3X1  g00348(.A(n1793), .B(n1792), .C(n1871), .Y(n1872));
  NAND2X1 g00349(.A(n1814), .B(n1818), .Y(n1873));
  AOI21X1 g00350(.A0(n1818), .A1(SI_1_), .B0(n1821), .Y(n1874));
  INVX1   g00351(.A(P1_DATAO_REG_3__SCAN_IN), .Y(n1875));
  OAI21X1 g00352(.A0(n1793), .A1(n1792), .B0(P2_DATAO_REG_3__SCAN_IN), .Y(n1876));
  OAI21X1 g00353(.A0(n1790), .A1(n1875), .B0(n1876), .Y(n1877));
  OAI22X1 g00354(.A0(n1856), .A1(SI_2_), .B0(SI_3_), .B1(n1877), .Y(n1878));
  AOI21X1 g00355(.A0(n1874), .A1(n1873), .B0(n1878), .Y(n1879));
  NOR2X1  g00356(.A(n1877), .B(SI_3_), .Y(n1880));
  NAND2X1 g00357(.A(n1877), .B(SI_3_), .Y(n1881));
  OAI21X1 g00358(.A0(n1880), .A1(n1857), .B0(n1881), .Y(n1882));
  NOR2X1  g00359(.A(n1882), .B(n1879), .Y(n1883));
  INVX1   g00360(.A(P1_DATAO_REG_4__SCAN_IN), .Y(n1884));
  NOR3X1  g00361(.A(n1793), .B(n1792), .C(n1884), .Y(n1885));
  AOI21X1 g00362(.A0(n1789), .A1(n1786), .B0(n1871), .Y(n1886));
  NOR2X1  g00363(.A(n1886), .B(n1885), .Y(n1887));
  XOR2X1  g00364(.A(n1887), .B(SI_4_), .Y(n1888));
  XOR2X1  g00365(.A(n1888), .B(n1883), .Y(n1889));
  AOI21X1 g00366(.A0(n1889), .A1(n1790), .B0(n1872), .Y(n1890));
  INVX1   g00367(.A(P1_IR_REG_4__SCAN_IN), .Y(n1891));
  NOR4X1  g00368(.A(P1_IR_REG_2__SCAN_IN), .B(P1_IR_REG_1__SCAN_IN), .C(P1_IR_REG_0__SCAN_IN), .D(P1_IR_REG_3__SCAN_IN), .Y(n1892));
  NAND3X1 g00369(.A(n1867), .B(n1891), .C(n1866), .Y(n1893));
  OAI21X1 g00370(.A0(n1892), .A1(n1891), .B0(n1893), .Y(n1894));
  NOR3X1  g00371(.A(n1894), .B(P1_U3086), .C(n1827), .Y(n1895));
  AOI21X1 g00372(.A0(n1803), .A1(P1_IR_REG_4__SCAN_IN), .B0(n1895), .Y(n1896));
  OAI21X1 g00373(.A0(n1890), .A1(P1_STATE_REG_SCAN_IN), .B0(n1896), .Y(P1_U3351));
  INVX1   g00374(.A(P2_DATAO_REG_5__SCAN_IN), .Y(n1898));
  NOR3X1  g00375(.A(n1793), .B(n1792), .C(n1898), .Y(n1899));
  OAI21X1 g00376(.A0(n1886), .A1(n1885), .B0(SI_4_), .Y(n1900));
  INVX1   g00377(.A(SI_4_), .Y(n1901));
  NAND2X1 g00378(.A(n1887), .B(n1901), .Y(n1902));
  OAI21X1 g00379(.A0(n1882), .A1(n1879), .B0(n1902), .Y(n1903));
  INVX1   g00380(.A(P1_DATAO_REG_5__SCAN_IN), .Y(n1904));
  NOR3X1  g00381(.A(n1793), .B(n1792), .C(n1904), .Y(n1905));
  AOI21X1 g00382(.A0(n1789), .A1(n1786), .B0(n1898), .Y(n1906));
  NOR2X1  g00383(.A(n1906), .B(n1905), .Y(n1907));
  XOR2X1  g00384(.A(n1907), .B(SI_5_), .Y(n1908));
  INVX1   g00385(.A(n1908), .Y(n1909));
  NAND3X1 g00386(.A(n1909), .B(n1903), .C(n1900), .Y(n1910));
  INVX1   g00387(.A(n1900), .Y(n1911));
  INVX1   g00388(.A(SI_3_), .Y(n1912));
  AOI22X1 g00389(.A0(n1839), .A1(n1850), .B0(n1912), .B1(n1861), .Y(n1913));
  OAI21X1 g00390(.A0(n1835), .A1(n1834), .B0(n1913), .Y(n1914));
  NOR2X1  g00391(.A(n1839), .B(n1850), .Y(n1915));
  NAND2X1 g00392(.A(n1861), .B(n1912), .Y(n1916));
  NOR2X1  g00393(.A(n1861), .B(n1912), .Y(n1917));
  AOI21X1 g00394(.A0(n1916), .A1(n1915), .B0(n1917), .Y(n1918));
  NOR3X1  g00395(.A(n1886), .B(n1885), .C(SI_4_), .Y(n1919));
  AOI21X1 g00396(.A0(n1918), .A1(n1914), .B0(n1919), .Y(n1920));
  OAI21X1 g00397(.A0(n1920), .A1(n1911), .B0(n1908), .Y(n1921));
  AOI21X1 g00398(.A0(n1921), .A1(n1910), .B0(n1837), .Y(n1922));
  OAI21X1 g00399(.A0(n1922), .A1(n1899), .B0(P1_U3086), .Y(n1923));
  XOR2X1  g00400(.A(n1893), .B(P1_IR_REG_5__SCAN_IN), .Y(n1924));
  AOI22X1 g00401(.A0(n1828), .A1(n1924), .B0(n1803), .B1(P1_IR_REG_5__SCAN_IN), .Y(n1925));
  NAND2X1 g00402(.A(n1925), .B(n1923), .Y(P1_U3350));
  INVX1   g00403(.A(P2_DATAO_REG_6__SCAN_IN), .Y(n1927));
  NOR3X1  g00404(.A(n1793), .B(n1792), .C(n1927), .Y(n1928));
  NAND2X1 g00405(.A(n1918), .B(n1914), .Y(n1929));
  NOR3X1  g00406(.A(n1906), .B(n1905), .C(SI_5_), .Y(n1930));
  OAI21X1 g00407(.A0(n1906), .A1(n1905), .B0(SI_5_), .Y(n1931));
  OAI21X1 g00408(.A0(n1930), .A1(n1900), .B0(n1931), .Y(n1932));
  NOR2X1  g00409(.A(n1930), .B(n1919), .Y(n1933));
  AOI21X1 g00410(.A0(n1933), .A1(n1929), .B0(n1932), .Y(n1934));
  INVX1   g00411(.A(P1_DATAO_REG_6__SCAN_IN), .Y(n1935));
  NOR3X1  g00412(.A(n1793), .B(n1792), .C(n1935), .Y(n1936));
  AOI21X1 g00413(.A0(n1789), .A1(n1786), .B0(n1927), .Y(n1937));
  NOR2X1  g00414(.A(n1937), .B(n1936), .Y(n1938));
  XOR2X1  g00415(.A(n1938), .B(SI_6_), .Y(n1939));
  XOR2X1  g00416(.A(n1939), .B(n1934), .Y(n1940));
  AOI21X1 g00417(.A0(n1940), .A1(n1790), .B0(n1928), .Y(n1941));
  INVX1   g00418(.A(P1_IR_REG_5__SCAN_IN), .Y(n1942));
  NAND4X1 g00419(.A(n1942), .B(n1891), .C(n1866), .D(n1867), .Y(n1943));
  INVX1   g00420(.A(P1_IR_REG_6__SCAN_IN), .Y(n1944));
  NAND2X1 g00421(.A(n1944), .B(n1942), .Y(n1945));
  NOR2X1  g00422(.A(n1945), .B(n1893), .Y(n1946));
  AOI21X1 g00423(.A0(n1943), .A1(P1_IR_REG_6__SCAN_IN), .B0(n1946), .Y(n1947));
  AOI22X1 g00424(.A0(n1828), .A1(n1947), .B0(n1803), .B1(P1_IR_REG_6__SCAN_IN), .Y(n1948));
  OAI21X1 g00425(.A0(n1941), .A1(P1_STATE_REG_SCAN_IN), .B0(n1948), .Y(P1_U3349));
  INVX1   g00426(.A(P2_DATAO_REG_7__SCAN_IN), .Y(n1950));
  NOR3X1  g00427(.A(n1793), .B(n1792), .C(n1950), .Y(n1951));
  NOR3X1  g00428(.A(n1937), .B(n1936), .C(SI_6_), .Y(n1952));
  NOR3X1  g00429(.A(n1952), .B(n1930), .C(n1919), .Y(n1953));
  OAI21X1 g00430(.A0(n1882), .A1(n1879), .B0(n1953), .Y(n1954));
  INVX1   g00431(.A(SI_6_), .Y(n1955));
  NAND3X1 g00432(.A(n1789), .B(n1786), .C(P1_DATAO_REG_6__SCAN_IN), .Y(n1956));
  OAI21X1 g00433(.A0(n1793), .A1(n1792), .B0(P2_DATAO_REG_6__SCAN_IN), .Y(n1957));
  NAND3X1 g00434(.A(n1957), .B(n1956), .C(n1955), .Y(n1958));
  AOI21X1 g00435(.A0(n1957), .A1(n1956), .B0(n1955), .Y(n1959));
  AOI21X1 g00436(.A0(n1958), .A1(n1932), .B0(n1959), .Y(n1960));
  NAND2X1 g00437(.A(n1960), .B(n1954), .Y(n1961));
  INVX1   g00438(.A(SI_7_), .Y(n1962));
  INVX1   g00439(.A(P1_DATAO_REG_7__SCAN_IN), .Y(n1963));
  NOR3X1  g00440(.A(n1793), .B(n1792), .C(n1963), .Y(n1964));
  AOI21X1 g00441(.A0(n1789), .A1(n1786), .B0(n1950), .Y(n1965));
  NOR2X1  g00442(.A(n1965), .B(n1964), .Y(n1966));
  XOR2X1  g00443(.A(n1966), .B(n1962), .Y(n1967));
  XOR2X1  g00444(.A(n1967), .B(n1961), .Y(n1968));
  AOI21X1 g00445(.A0(n1968), .A1(n1790), .B0(n1951), .Y(n1969));
  INVX1   g00446(.A(P1_IR_REG_7__SCAN_IN), .Y(n1970));
  XOR2X1  g00447(.A(n1946), .B(n1970), .Y(n1971));
  AOI22X1 g00448(.A0(n1828), .A1(n1971), .B0(n1803), .B1(P1_IR_REG_7__SCAN_IN), .Y(n1972));
  OAI21X1 g00449(.A0(n1969), .A1(P1_STATE_REG_SCAN_IN), .B0(n1972), .Y(P1_U3348));
  INVX1   g00450(.A(P2_DATAO_REG_8__SCAN_IN), .Y(n1974));
  NOR3X1  g00451(.A(n1793), .B(n1792), .C(n1974), .Y(n1975));
  NAND2X1 g00452(.A(n1958), .B(n1933), .Y(n1976));
  AOI21X1 g00453(.A0(n1918), .A1(n1914), .B0(n1976), .Y(n1977));
  NAND2X1 g00454(.A(n1958), .B(n1932), .Y(n1978));
  OAI21X1 g00455(.A0(n1938), .A1(n1955), .B0(n1978), .Y(n1979));
  NAND3X1 g00456(.A(n1789), .B(n1786), .C(P1_DATAO_REG_7__SCAN_IN), .Y(n1980));
  OAI21X1 g00457(.A0(n1793), .A1(n1792), .B0(P2_DATAO_REG_7__SCAN_IN), .Y(n1981));
  NAND2X1 g00458(.A(n1981), .B(n1980), .Y(n1982));
  OAI22X1 g00459(.A0(n1979), .A1(n1977), .B0(SI_7_), .B1(n1982), .Y(n1983));
  OAI21X1 g00460(.A0(n1966), .A1(n1962), .B0(n1983), .Y(n1984));
  INVX1   g00461(.A(SI_8_), .Y(n1985));
  AOI21X1 g00462(.A0(n1789), .A1(n1786), .B0(n1974), .Y(n1986));
  AOI21X1 g00463(.A0(n1837), .A1(P1_DATAO_REG_8__SCAN_IN), .B0(n1986), .Y(n1987));
  XOR2X1  g00464(.A(n1987), .B(n1985), .Y(n1988));
  XOR2X1  g00465(.A(n1988), .B(n1984), .Y(n1989));
  AOI21X1 g00466(.A0(n1989), .A1(n1790), .B0(n1975), .Y(n1990));
  INVX1   g00467(.A(P1_IR_REG_8__SCAN_IN), .Y(n1991));
  AOI21X1 g00468(.A0(n1946), .A1(n1970), .B0(n1991), .Y(n1992));
  NOR4X1  g00469(.A(P1_IR_REG_5__SCAN_IN), .B(P1_IR_REG_4__SCAN_IN), .C(P1_IR_REG_3__SCAN_IN), .D(P1_IR_REG_6__SCAN_IN), .Y(n1993));
  NAND4X1 g00470(.A(n1867), .B(n1991), .C(n1970), .D(n1993), .Y(n1994));
  INVX1   g00471(.A(n1994), .Y(n1995));
  NOR2X1  g00472(.A(n1995), .B(n1992), .Y(n1996));
  AOI22X1 g00473(.A0(n1828), .A1(n1996), .B0(n1803), .B1(P1_IR_REG_8__SCAN_IN), .Y(n1997));
  OAI21X1 g00474(.A0(n1990), .A1(P1_STATE_REG_SCAN_IN), .B0(n1997), .Y(P1_U3347));
  INVX1   g00475(.A(P2_DATAO_REG_9__SCAN_IN), .Y(n1999));
  NOR3X1  g00476(.A(n1793), .B(n1792), .C(n1999), .Y(n2000));
  AOI21X1 g00477(.A0(n1981), .A1(n1980), .B0(n1962), .Y(n2001));
  NAND3X1 g00478(.A(n1789), .B(n1786), .C(P1_DATAO_REG_8__SCAN_IN), .Y(n2002));
  OAI21X1 g00479(.A0(n1793), .A1(n1792), .B0(P2_DATAO_REG_8__SCAN_IN), .Y(n2003));
  NAND3X1 g00480(.A(n2003), .B(n2002), .C(n1985), .Y(n2004));
  AOI21X1 g00481(.A0(n2003), .A1(n2002), .B0(n1985), .Y(n2005));
  AOI21X1 g00482(.A0(n2004), .A1(n2001), .B0(n2005), .Y(n2006));
  INVX1   g00483(.A(n2006), .Y(n2007));
  AOI22X1 g00484(.A0(n1966), .A1(n1962), .B0(n1985), .B1(n1987), .Y(n2008));
  AOI21X1 g00485(.A0(n2008), .A1(n1961), .B0(n2007), .Y(n2009));
  AOI21X1 g00486(.A0(n1789), .A1(n1786), .B0(n1999), .Y(n2010));
  AOI21X1 g00487(.A0(n1837), .A1(P1_DATAO_REG_9__SCAN_IN), .B0(n2010), .Y(n2011));
  XOR2X1  g00488(.A(n2011), .B(SI_9_), .Y(n2012));
  XOR2X1  g00489(.A(n2012), .B(n2009), .Y(n2013));
  AOI21X1 g00490(.A0(n2013), .A1(n1790), .B0(n2000), .Y(n2014));
  XOR2X1  g00491(.A(n1994), .B(P1_IR_REG_9__SCAN_IN), .Y(n2015));
  AOI22X1 g00492(.A0(n1828), .A1(n2015), .B0(n1803), .B1(P1_IR_REG_9__SCAN_IN), .Y(n2016));
  OAI21X1 g00493(.A0(n2014), .A1(P1_STATE_REG_SCAN_IN), .B0(n2016), .Y(P1_U3346));
  INVX1   g00494(.A(P2_DATAO_REG_10__SCAN_IN), .Y(n2018));
  NOR3X1  g00495(.A(n1793), .B(n1792), .C(n2018), .Y(n2019));
  INVX1   g00496(.A(P1_DATAO_REG_9__SCAN_IN), .Y(n2020));
  OAI21X1 g00497(.A0(n1793), .A1(n1792), .B0(P2_DATAO_REG_9__SCAN_IN), .Y(n2021));
  OAI21X1 g00498(.A0(n1790), .A1(n2020), .B0(n2021), .Y(n2022));
  NOR2X1  g00499(.A(n2022), .B(SI_9_), .Y(n2023));
  NAND2X1 g00500(.A(n2022), .B(SI_9_), .Y(n2024));
  OAI21X1 g00501(.A0(n2023), .A1(n2006), .B0(n2024), .Y(n2025));
  OAI21X1 g00502(.A0(n1982), .A1(SI_7_), .B0(n2004), .Y(n2026));
  NOR2X1  g00503(.A(n2023), .B(n2026), .Y(n2027));
  AOI21X1 g00504(.A0(n2027), .A1(n1961), .B0(n2025), .Y(n2028));
  AOI21X1 g00505(.A0(n1789), .A1(n1786), .B0(n2018), .Y(n2029));
  AOI21X1 g00506(.A0(n1837), .A1(P1_DATAO_REG_10__SCAN_IN), .B0(n2029), .Y(n2030));
  XOR2X1  g00507(.A(n2030), .B(SI_10_), .Y(n2031));
  XOR2X1  g00508(.A(n2031), .B(n2028), .Y(n2032));
  AOI21X1 g00509(.A0(n2032), .A1(n1790), .B0(n2019), .Y(n2033));
  INVX1   g00510(.A(P1_IR_REG_9__SCAN_IN), .Y(n2034));
  INVX1   g00511(.A(P1_IR_REG_10__SCAN_IN), .Y(n2035));
  AOI21X1 g00512(.A0(n1995), .A1(n2034), .B0(n2035), .Y(n2036));
  NOR2X1  g00513(.A(P1_IR_REG_10__SCAN_IN), .B(P1_IR_REG_9__SCAN_IN), .Y(n2037));
  INVX1   g00514(.A(n2037), .Y(n2038));
  NOR2X1  g00515(.A(n2038), .B(n1994), .Y(n2039));
  NOR2X1  g00516(.A(n2039), .B(n2036), .Y(n2040));
  AOI22X1 g00517(.A0(n1828), .A1(n2040), .B0(n1803), .B1(P1_IR_REG_10__SCAN_IN), .Y(n2041));
  OAI21X1 g00518(.A0(n2033), .A1(P1_STATE_REG_SCAN_IN), .B0(n2041), .Y(P1_U3345));
  INVX1   g00519(.A(P2_DATAO_REG_11__SCAN_IN), .Y(n2043));
  NOR3X1  g00520(.A(n1793), .B(n1792), .C(n2043), .Y(n2044));
  INVX1   g00521(.A(P1_DATAO_REG_10__SCAN_IN), .Y(n2045));
  NOR3X1  g00522(.A(n1793), .B(n1792), .C(n2045), .Y(n2046));
  NOR3X1  g00523(.A(n2029), .B(n2046), .C(SI_10_), .Y(n2047));
  NOR3X1  g00524(.A(n2047), .B(n2023), .C(n2026), .Y(n2048));
  OAI21X1 g00525(.A0(n1979), .A1(n1977), .B0(n2048), .Y(n2049));
  INVX1   g00526(.A(n2047), .Y(n2050));
  INVX1   g00527(.A(SI_10_), .Y(n2051));
  NOR2X1  g00528(.A(n2030), .B(n2051), .Y(n2052));
  AOI21X1 g00529(.A0(n2050), .A1(n2025), .B0(n2052), .Y(n2053));
  NAND2X1 g00530(.A(n2053), .B(n2049), .Y(n2054));
  NAND3X1 g00531(.A(n1789), .B(n1786), .C(P1_DATAO_REG_11__SCAN_IN), .Y(n2055));
  OAI21X1 g00532(.A0(n1793), .A1(n1792), .B0(P2_DATAO_REG_11__SCAN_IN), .Y(n2056));
  NAND2X1 g00533(.A(n2056), .B(n2055), .Y(n2057));
  XOR2X1  g00534(.A(n2057), .B(SI_11_), .Y(n2058));
  XOR2X1  g00535(.A(n2058), .B(n2054), .Y(n2059));
  AOI21X1 g00536(.A0(n2059), .A1(n1790), .B0(n2044), .Y(n2060));
  INVX1   g00537(.A(P1_IR_REG_11__SCAN_IN), .Y(n2061));
  XOR2X1  g00538(.A(n2039), .B(n2061), .Y(n2062));
  AOI22X1 g00539(.A0(n1828), .A1(n2062), .B0(n1803), .B1(P1_IR_REG_11__SCAN_IN), .Y(n2063));
  OAI21X1 g00540(.A0(n2060), .A1(P1_STATE_REG_SCAN_IN), .B0(n2063), .Y(P1_U3344));
  INVX1   g00541(.A(P2_DATAO_REG_12__SCAN_IN), .Y(n2065));
  NOR3X1  g00542(.A(n1793), .B(n1792), .C(n2065), .Y(n2066));
  INVX1   g00543(.A(SI_11_), .Y(n2067));
  INVX1   g00544(.A(n2057), .Y(n2068));
  NAND2X1 g00545(.A(n2050), .B(n2027), .Y(n2069));
  AOI21X1 g00546(.A0(n1960), .A1(n1954), .B0(n2069), .Y(n2070));
  NAND2X1 g00547(.A(n2050), .B(n2025), .Y(n2071));
  OAI21X1 g00548(.A0(n2030), .A1(n2051), .B0(n2071), .Y(n2072));
  OAI22X1 g00549(.A0(n2072), .A1(n2070), .B0(SI_11_), .B1(n2057), .Y(n2073));
  OAI21X1 g00550(.A0(n2068), .A1(n2067), .B0(n2073), .Y(n2074));
  INVX1   g00551(.A(SI_12_), .Y(n2075));
  OAI21X1 g00552(.A0(n1793), .A1(n1792), .B0(P2_DATAO_REG_12__SCAN_IN), .Y(n2076));
  INVX1   g00553(.A(n2076), .Y(n2077));
  AOI21X1 g00554(.A0(n1837), .A1(P1_DATAO_REG_12__SCAN_IN), .B0(n2077), .Y(n2078));
  XOR2X1  g00555(.A(n2078), .B(n2075), .Y(n2079));
  XOR2X1  g00556(.A(n2079), .B(n2074), .Y(n2080));
  AOI21X1 g00557(.A0(n2080), .A1(n1790), .B0(n2066), .Y(n2081));
  INVX1   g00558(.A(P1_IR_REG_12__SCAN_IN), .Y(n2082));
  AOI21X1 g00559(.A0(n2039), .A1(n2061), .B0(n2082), .Y(n2083));
  NOR4X1  g00560(.A(n1994), .B(P1_IR_REG_12__SCAN_IN), .C(P1_IR_REG_11__SCAN_IN), .D(n2038), .Y(n2084));
  NOR2X1  g00561(.A(n2084), .B(n2083), .Y(n2085));
  AOI22X1 g00562(.A0(n1828), .A1(n2085), .B0(n1803), .B1(P1_IR_REG_12__SCAN_IN), .Y(n2086));
  OAI21X1 g00563(.A0(n2081), .A1(P1_STATE_REG_SCAN_IN), .B0(n2086), .Y(P1_U3343));
  INVX1   g00564(.A(P2_DATAO_REG_13__SCAN_IN), .Y(n2088));
  NOR3X1  g00565(.A(n1793), .B(n1792), .C(n2088), .Y(n2089));
  AOI21X1 g00566(.A0(n2056), .A1(n2055), .B0(n2067), .Y(n2090));
  NAND3X1 g00567(.A(n1789), .B(n1786), .C(P1_DATAO_REG_12__SCAN_IN), .Y(n2091));
  NAND3X1 g00568(.A(n2076), .B(n2091), .C(n2075), .Y(n2092));
  AOI21X1 g00569(.A0(n2076), .A1(n2091), .B0(n2075), .Y(n2093));
  AOI21X1 g00570(.A0(n2092), .A1(n2090), .B0(n2093), .Y(n2094));
  OAI21X1 g00571(.A0(n2057), .A1(SI_11_), .B0(n2092), .Y(n2095));
  INVX1   g00572(.A(n2095), .Y(n2096));
  OAI21X1 g00573(.A0(n2072), .A1(n2070), .B0(n2096), .Y(n2097));
  NAND2X1 g00574(.A(n2097), .B(n2094), .Y(n2098));
  INVX1   g00575(.A(P1_DATAO_REG_13__SCAN_IN), .Y(n2099));
  OAI21X1 g00576(.A0(n1793), .A1(n1792), .B0(P2_DATAO_REG_13__SCAN_IN), .Y(n2100));
  OAI21X1 g00577(.A0(n1790), .A1(n2099), .B0(n2100), .Y(n2101));
  XOR2X1  g00578(.A(n2101), .B(SI_13_), .Y(n2102));
  XOR2X1  g00579(.A(n2102), .B(n2098), .Y(n2103));
  AOI21X1 g00580(.A0(n2103), .A1(n1790), .B0(n2089), .Y(n2104));
  INVX1   g00581(.A(P1_IR_REG_13__SCAN_IN), .Y(n2105));
  XOR2X1  g00582(.A(n2084), .B(n2105), .Y(n2106));
  AOI22X1 g00583(.A0(n1828), .A1(n2106), .B0(n1803), .B1(P1_IR_REG_13__SCAN_IN), .Y(n2107));
  OAI21X1 g00584(.A0(n2104), .A1(P1_STATE_REG_SCAN_IN), .B0(n2107), .Y(P1_U3342));
  INVX1   g00585(.A(P2_DATAO_REG_14__SCAN_IN), .Y(n2109));
  NOR3X1  g00586(.A(n1793), .B(n1792), .C(n2109), .Y(n2110));
  NOR2X1  g00587(.A(n2101), .B(SI_13_), .Y(n2111));
  NAND2X1 g00588(.A(n2101), .B(SI_13_), .Y(n2112));
  OAI21X1 g00589(.A0(n2111), .A1(n2094), .B0(n2112), .Y(n2113));
  NOR2X1  g00590(.A(n2111), .B(n2095), .Y(n2114));
  AOI21X1 g00591(.A0(n2114), .A1(n2054), .B0(n2113), .Y(n2115));
  AOI21X1 g00592(.A0(n1789), .A1(n1786), .B0(n2109), .Y(n2116));
  AOI21X1 g00593(.A0(n1837), .A1(P1_DATAO_REG_14__SCAN_IN), .B0(n2116), .Y(n2117));
  XOR2X1  g00594(.A(n2117), .B(SI_14_), .Y(n2118));
  XOR2X1  g00595(.A(n2118), .B(n2115), .Y(n2119));
  AOI21X1 g00596(.A0(n2119), .A1(n1790), .B0(n2110), .Y(n2120));
  INVX1   g00597(.A(P1_IR_REG_14__SCAN_IN), .Y(n2121));
  AOI21X1 g00598(.A0(n2084), .A1(n2105), .B0(n2121), .Y(n2122));
  INVX1   g00599(.A(n2084), .Y(n2123));
  NOR3X1  g00600(.A(n2123), .B(P1_IR_REG_14__SCAN_IN), .C(P1_IR_REG_13__SCAN_IN), .Y(n2124));
  NOR2X1  g00601(.A(n2124), .B(n2122), .Y(n2125));
  AOI22X1 g00602(.A0(n1828), .A1(n2125), .B0(n1803), .B1(P1_IR_REG_14__SCAN_IN), .Y(n2126));
  OAI21X1 g00603(.A0(n2120), .A1(P1_STATE_REG_SCAN_IN), .B0(n2126), .Y(P1_U3341));
  INVX1   g00604(.A(P2_DATAO_REG_15__SCAN_IN), .Y(n2128));
  NOR3X1  g00605(.A(n1793), .B(n1792), .C(n2128), .Y(n2129));
  INVX1   g00606(.A(SI_14_), .Y(n2130));
  INVX1   g00607(.A(P1_DATAO_REG_14__SCAN_IN), .Y(n2131));
  NOR3X1  g00608(.A(n1793), .B(n1792), .C(n2131), .Y(n2132));
  NOR3X1  g00609(.A(n2116), .B(n2132), .C(SI_14_), .Y(n2133));
  INVX1   g00610(.A(n2133), .Y(n2134));
  NAND2X1 g00611(.A(n2134), .B(n2113), .Y(n2135));
  OAI21X1 g00612(.A0(n2117), .A1(n2130), .B0(n2135), .Y(n2136));
  NOR3X1  g00613(.A(n2133), .B(n2111), .C(n2095), .Y(n2137));
  AOI21X1 g00614(.A0(n2137), .A1(n2054), .B0(n2136), .Y(n2138));
  AOI21X1 g00615(.A0(n1789), .A1(n1786), .B0(n2128), .Y(n2139));
  AOI21X1 g00616(.A0(n1837), .A1(P1_DATAO_REG_15__SCAN_IN), .B0(n2139), .Y(n2140));
  XOR2X1  g00617(.A(n2140), .B(SI_15_), .Y(n2141));
  XOR2X1  g00618(.A(n2141), .B(n2138), .Y(n2142));
  AOI21X1 g00619(.A0(n2142), .A1(n1790), .B0(n2129), .Y(n2143));
  INVX1   g00620(.A(P1_IR_REG_15__SCAN_IN), .Y(n2144));
  XOR2X1  g00621(.A(n2124), .B(n2144), .Y(n2145));
  AOI22X1 g00622(.A0(n1828), .A1(n2145), .B0(n1803), .B1(P1_IR_REG_15__SCAN_IN), .Y(n2146));
  OAI21X1 g00623(.A0(n2143), .A1(P1_STATE_REG_SCAN_IN), .B0(n2146), .Y(P1_U3340));
  INVX1   g00624(.A(P2_DATAO_REG_16__SCAN_IN), .Y(n2148));
  NOR3X1  g00625(.A(n1793), .B(n1792), .C(n2148), .Y(n2149));
  INVX1   g00626(.A(SI_15_), .Y(n2150));
  NAND2X1 g00627(.A(n2140), .B(n2150), .Y(n2151));
  NAND2X1 g00628(.A(n2151), .B(n2137), .Y(n2152));
  AOI21X1 g00629(.A0(n2053), .A1(n2049), .B0(n2152), .Y(n2153));
  NOR2X1  g00630(.A(n2117), .B(n2130), .Y(n2154));
  AOI21X1 g00631(.A0(n2134), .A1(n2113), .B0(n2154), .Y(n2155));
  INVX1   g00632(.A(n2151), .Y(n2156));
  NOR2X1  g00633(.A(n2140), .B(n2150), .Y(n2157));
  INVX1   g00634(.A(n2157), .Y(n2158));
  OAI21X1 g00635(.A0(n2156), .A1(n2155), .B0(n2158), .Y(n2159));
  NOR2X1  g00636(.A(n2159), .B(n2153), .Y(n2160));
  AOI21X1 g00637(.A0(n1789), .A1(n1786), .B0(n2148), .Y(n2161));
  AOI21X1 g00638(.A0(n1837), .A1(P1_DATAO_REG_16__SCAN_IN), .B0(n2161), .Y(n2162));
  XOR2X1  g00639(.A(n2162), .B(SI_16_), .Y(n2163));
  XOR2X1  g00640(.A(n2163), .B(n2160), .Y(n2164));
  AOI21X1 g00641(.A0(n2164), .A1(n1790), .B0(n2149), .Y(n2165));
  INVX1   g00642(.A(P1_IR_REG_16__SCAN_IN), .Y(n2166));
  NOR4X1  g00643(.A(P1_IR_REG_15__SCAN_IN), .B(P1_IR_REG_14__SCAN_IN), .C(P1_IR_REG_13__SCAN_IN), .D(n2123), .Y(n2167));
  NOR4X1  g00644(.A(P1_IR_REG_12__SCAN_IN), .B(P1_IR_REG_11__SCAN_IN), .C(P1_IR_REG_10__SCAN_IN), .D(P1_IR_REG_13__SCAN_IN), .Y(n2168));
  NAND2X1 g00645(.A(n2168), .B(n2121), .Y(n2169));
  NOR2X1  g00646(.A(P1_IR_REG_16__SCAN_IN), .B(P1_IR_REG_15__SCAN_IN), .Y(n2170));
  NAND3X1 g00647(.A(n2170), .B(n1844), .C(n1942), .Y(n2171));
  NAND4X1 g00648(.A(n1991), .B(n1970), .C(n1944), .D(n2034), .Y(n2172));
  NOR2X1  g00649(.A(P1_IR_REG_3__SCAN_IN), .B(P1_IR_REG_2__SCAN_IN), .Y(n2173));
  NAND2X1 g00650(.A(n2173), .B(n1891), .Y(n2174));
  NOR4X1  g00651(.A(n2172), .B(n2171), .C(n2169), .D(n2174), .Y(n2175));
  INVX1   g00652(.A(n2175), .Y(n2176));
  OAI21X1 g00653(.A0(n2167), .A1(n2166), .B0(n2176), .Y(n2177));
  INVX1   g00654(.A(n2177), .Y(n2178));
  AOI22X1 g00655(.A0(n1828), .A1(n2178), .B0(n1803), .B1(P1_IR_REG_16__SCAN_IN), .Y(n2179));
  OAI21X1 g00656(.A0(n2165), .A1(P1_STATE_REG_SCAN_IN), .B0(n2179), .Y(P1_U3339));
  INVX1   g00657(.A(P2_DATAO_REG_17__SCAN_IN), .Y(n2181));
  NOR3X1  g00658(.A(n1793), .B(n1792), .C(n2181), .Y(n2182));
  INVX1   g00659(.A(SI_16_), .Y(n2183));
  NOR2X1  g00660(.A(n2162), .B(n2183), .Y(n2184));
  NOR4X1  g00661(.A(n2133), .B(n2111), .C(n2095), .D(n2156), .Y(n2185));
  OAI21X1 g00662(.A0(n2072), .A1(n2070), .B0(n2185), .Y(n2186));
  AOI21X1 g00663(.A0(n2151), .A1(n2136), .B0(n2157), .Y(n2187));
  AOI22X1 g00664(.A0(n2187), .A1(n2186), .B0(n2183), .B1(n2162), .Y(n2188));
  NOR2X1  g00665(.A(n2188), .B(n2184), .Y(n2189));
  AOI21X1 g00666(.A0(n1789), .A1(n1786), .B0(n2181), .Y(n2190));
  AOI21X1 g00667(.A0(n1837), .A1(P1_DATAO_REG_17__SCAN_IN), .B0(n2190), .Y(n2191));
  XOR2X1  g00668(.A(n2191), .B(SI_17_), .Y(n2192));
  XOR2X1  g00669(.A(n2192), .B(n2189), .Y(n2193));
  AOI21X1 g00670(.A0(n2193), .A1(n1790), .B0(n2182), .Y(n2194));
  INVX1   g00671(.A(P1_IR_REG_17__SCAN_IN), .Y(n2195));
  XOR2X1  g00672(.A(n2175), .B(n2195), .Y(n2196));
  AOI22X1 g00673(.A0(n1828), .A1(n2196), .B0(n1803), .B1(P1_IR_REG_17__SCAN_IN), .Y(n2197));
  OAI21X1 g00674(.A0(n2194), .A1(P1_STATE_REG_SCAN_IN), .B0(n2197), .Y(P1_U3338));
  INVX1   g00675(.A(P2_DATAO_REG_18__SCAN_IN), .Y(n2199));
  NOR3X1  g00676(.A(n1793), .B(n1792), .C(n2199), .Y(n2200));
  INVX1   g00677(.A(SI_17_), .Y(n2201));
  NOR2X1  g00678(.A(n2191), .B(n2201), .Y(n2202));
  INVX1   g00679(.A(n2184), .Y(n2203));
  NAND2X1 g00680(.A(n2162), .B(n2183), .Y(n2204));
  OAI21X1 g00681(.A0(n2159), .A1(n2153), .B0(n2204), .Y(n2205));
  AOI22X1 g00682(.A0(n2205), .A1(n2203), .B0(n2201), .B1(n2191), .Y(n2206));
  NOR2X1  g00683(.A(n2206), .B(n2202), .Y(n2207));
  AOI21X1 g00684(.A0(n1789), .A1(n1786), .B0(n2199), .Y(n2208));
  AOI21X1 g00685(.A0(n1837), .A1(P1_DATAO_REG_18__SCAN_IN), .B0(n2208), .Y(n2209));
  XOR2X1  g00686(.A(n2209), .B(SI_18_), .Y(n2210));
  XOR2X1  g00687(.A(n2210), .B(n2207), .Y(n2211));
  AOI21X1 g00688(.A0(n2211), .A1(n1790), .B0(n2200), .Y(n2212));
  OAI21X1 g00689(.A0(n2176), .A1(P1_IR_REG_17__SCAN_IN), .B0(P1_IR_REG_18__SCAN_IN), .Y(n2213));
  NOR3X1  g00690(.A(P1_IR_REG_12__SCAN_IN), .B(P1_IR_REG_11__SCAN_IN), .C(P1_IR_REG_10__SCAN_IN), .Y(n2214));
  NAND2X1 g00691(.A(n2214), .B(n2105), .Y(n2215));
  NOR2X1  g00692(.A(n2215), .B(P1_IR_REG_14__SCAN_IN), .Y(n2216));
  NOR4X1  g00693(.A(P1_IR_REG_17__SCAN_IN), .B(P1_IR_REG_5__SCAN_IN), .C(P1_IR_REG_1__SCAN_IN), .D(P1_IR_REG_18__SCAN_IN), .Y(n2217));
  NAND2X1 g00694(.A(n2217), .B(n2170), .Y(n2218));
  INVX1   g00695(.A(P1_IR_REG_0__SCAN_IN), .Y(n2219));
  NAND4X1 g00696(.A(n1866), .B(n1843), .C(n2219), .D(n1891), .Y(n2220));
  NOR3X1  g00697(.A(n2220), .B(n2218), .C(n2172), .Y(n2221));
  NAND2X1 g00698(.A(n2221), .B(n2216), .Y(n2222));
  NAND2X1 g00699(.A(n2222), .B(n2213), .Y(n2223));
  INVX1   g00700(.A(n2223), .Y(n2224));
  AOI22X1 g00701(.A0(n1828), .A1(n2224), .B0(n1803), .B1(P1_IR_REG_18__SCAN_IN), .Y(n2225));
  OAI21X1 g00702(.A0(n2212), .A1(P1_STATE_REG_SCAN_IN), .B0(n2225), .Y(P1_U3337));
  INVX1   g00703(.A(P2_DATAO_REG_19__SCAN_IN), .Y(n2227));
  NOR3X1  g00704(.A(n1793), .B(n1792), .C(n2227), .Y(n2228));
  INVX1   g00705(.A(SI_18_), .Y(n2229));
  NOR2X1  g00706(.A(n2209), .B(n2229), .Y(n2230));
  INVX1   g00707(.A(n2202), .Y(n2231));
  INVX1   g00708(.A(n2191), .Y(n2232));
  OAI22X1 g00709(.A0(n2188), .A1(n2184), .B0(SI_17_), .B1(n2232), .Y(n2233));
  AOI22X1 g00710(.A0(n2233), .A1(n2231), .B0(n2229), .B1(n2209), .Y(n2234));
  NOR2X1  g00711(.A(n2234), .B(n2230), .Y(n2235));
  AOI21X1 g00712(.A0(n1789), .A1(n1786), .B0(n2227), .Y(n2236));
  AOI21X1 g00713(.A0(n1837), .A1(P1_DATAO_REG_19__SCAN_IN), .B0(n2236), .Y(n2237));
  XOR2X1  g00714(.A(n2237), .B(SI_19_), .Y(n2238));
  XOR2X1  g00715(.A(n2238), .B(n2235), .Y(n2239));
  AOI21X1 g00716(.A0(n2239), .A1(n1790), .B0(n2228), .Y(n2240));
  NOR2X1  g00717(.A(P1_IR_REG_6__SCAN_IN), .B(P1_IR_REG_5__SCAN_IN), .Y(n2241));
  NOR3X1  g00718(.A(P1_IR_REG_9__SCAN_IN), .B(P1_IR_REG_8__SCAN_IN), .C(P1_IR_REG_7__SCAN_IN), .Y(n2242));
  NAND2X1 g00719(.A(n2242), .B(n2241), .Y(n2243));
  NOR4X1  g00720(.A(P1_IR_REG_18__SCAN_IN), .B(P1_IR_REG_16__SCAN_IN), .C(P1_IR_REG_4__SCAN_IN), .D(P1_IR_REG_19__SCAN_IN), .Y(n2244));
  NAND4X1 g00721(.A(n1892), .B(n2195), .C(n2144), .D(n2244), .Y(n2245));
  NOR3X1  g00722(.A(n2245), .B(n2243), .C(n2169), .Y(n2246));
  AOI21X1 g00723(.A0(n2222), .A1(P1_IR_REG_19__SCAN_IN), .B0(n2246), .Y(n2247));
  AOI22X1 g00724(.A0(n1828), .A1(n2247), .B0(n1803), .B1(P1_IR_REG_19__SCAN_IN), .Y(n2248));
  OAI21X1 g00725(.A0(n2240), .A1(P1_STATE_REG_SCAN_IN), .B0(n2248), .Y(P1_U3336));
  INVX1   g00726(.A(P2_DATAO_REG_20__SCAN_IN), .Y(n2250));
  NOR3X1  g00727(.A(n1793), .B(n1792), .C(n2250), .Y(n2251));
  INVX1   g00728(.A(SI_19_), .Y(n2252));
  NOR2X1  g00729(.A(n2237), .B(n2252), .Y(n2253));
  INVX1   g00730(.A(n2253), .Y(n2254));
  INVX1   g00731(.A(n2237), .Y(n2255));
  OAI22X1 g00732(.A0(n2234), .A1(n2230), .B0(SI_19_), .B1(n2255), .Y(n2256));
  NAND2X1 g00733(.A(n2256), .B(n2254), .Y(n2257));
  AOI21X1 g00734(.A0(n1789), .A1(n1786), .B0(n2250), .Y(n2258));
  AOI21X1 g00735(.A0(n1837), .A1(P1_DATAO_REG_20__SCAN_IN), .B0(n2258), .Y(n2259));
  XOR2X1  g00736(.A(n2259), .B(SI_20_), .Y(n2260));
  XOR2X1  g00737(.A(n2260), .B(n2257), .Y(n2261));
  NOR2X1  g00738(.A(n2261), .B(n1837), .Y(n2262));
  NOR2X1  g00739(.A(n2262), .B(n2251), .Y(n2263));
  NOR2X1  g00740(.A(n2245), .B(n2243), .Y(n2264));
  NAND2X1 g00741(.A(n2264), .B(n2216), .Y(n2265));
  NAND4X1 g00742(.A(n2144), .B(n2121), .C(n2105), .D(n2214), .Y(n2266));
  NOR2X1  g00743(.A(P1_IR_REG_19__SCAN_IN), .B(P1_IR_REG_16__SCAN_IN), .Y(n2267));
  NOR3X1  g00744(.A(P1_IR_REG_18__SCAN_IN), .B(P1_IR_REG_17__SCAN_IN), .C(P1_IR_REG_1__SCAN_IN), .Y(n2268));
  NAND4X1 g00745(.A(n2267), .B(n2242), .C(n2241), .D(n2268), .Y(n2269));
  NOR4X1  g00746(.A(n2266), .B(n2220), .C(P1_IR_REG_20__SCAN_IN), .D(n2269), .Y(n2270));
  AOI21X1 g00747(.A0(n2265), .A1(P1_IR_REG_20__SCAN_IN), .B0(n2270), .Y(n2271));
  AOI22X1 g00748(.A0(n1828), .A1(n2271), .B0(n1803), .B1(P1_IR_REG_20__SCAN_IN), .Y(n2272));
  OAI21X1 g00749(.A0(n2263), .A1(P1_STATE_REG_SCAN_IN), .B0(n2272), .Y(P1_U3335));
  INVX1   g00750(.A(P2_DATAO_REG_21__SCAN_IN), .Y(n2274));
  NOR3X1  g00751(.A(n1793), .B(n1792), .C(n2274), .Y(n2275));
  INVX1   g00752(.A(SI_20_), .Y(n2276));
  NOR2X1  g00753(.A(n2259), .B(n2276), .Y(n2277));
  AOI22X1 g00754(.A0(n2256), .A1(n2254), .B0(n2276), .B1(n2259), .Y(n2278));
  NOR2X1  g00755(.A(n2278), .B(n2277), .Y(n2279));
  AOI21X1 g00756(.A0(n1789), .A1(n1786), .B0(n2274), .Y(n2280));
  AOI21X1 g00757(.A0(n1837), .A1(P1_DATAO_REG_21__SCAN_IN), .B0(n2280), .Y(n2281));
  XOR2X1  g00758(.A(n2281), .B(SI_21_), .Y(n2282));
  XOR2X1  g00759(.A(n2282), .B(n2279), .Y(n2283));
  AOI21X1 g00760(.A0(n2283), .A1(n1790), .B0(n2275), .Y(n2284));
  INVX1   g00761(.A(P1_IR_REG_21__SCAN_IN), .Y(n2285));
  XOR2X1  g00762(.A(n2270), .B(n2285), .Y(n2286));
  AOI22X1 g00763(.A0(n1828), .A1(n2286), .B0(n1803), .B1(P1_IR_REG_21__SCAN_IN), .Y(n2287));
  OAI21X1 g00764(.A0(n2284), .A1(P1_STATE_REG_SCAN_IN), .B0(n2287), .Y(P1_U3334));
  INVX1   g00765(.A(P2_DATAO_REG_22__SCAN_IN), .Y(n2289));
  NOR3X1  g00766(.A(n1793), .B(n1792), .C(n2289), .Y(n2290));
  INVX1   g00767(.A(SI_21_), .Y(n2291));
  NOR2X1  g00768(.A(n2281), .B(n2291), .Y(n2292));
  INVX1   g00769(.A(n2277), .Y(n2293));
  INVX1   g00770(.A(n2230), .Y(n2294));
  INVX1   g00771(.A(n2209), .Y(n2295));
  OAI22X1 g00772(.A0(n2206), .A1(n2202), .B0(SI_18_), .B1(n2295), .Y(n2296));
  AOI22X1 g00773(.A0(n2296), .A1(n2294), .B0(n2252), .B1(n2237), .Y(n2297));
  INVX1   g00774(.A(n2259), .Y(n2298));
  OAI22X1 g00775(.A0(n2297), .A1(n2253), .B0(SI_20_), .B1(n2298), .Y(n2299));
  AOI22X1 g00776(.A0(n2299), .A1(n2293), .B0(n2291), .B1(n2281), .Y(n2300));
  NOR2X1  g00777(.A(n2300), .B(n2292), .Y(n2301));
  AOI21X1 g00778(.A0(n1789), .A1(n1786), .B0(n2289), .Y(n2302));
  AOI21X1 g00779(.A0(n1837), .A1(P1_DATAO_REG_22__SCAN_IN), .B0(n2302), .Y(n2303));
  XOR2X1  g00780(.A(n2303), .B(SI_22_), .Y(n2304));
  XOR2X1  g00781(.A(n2304), .B(n2301), .Y(n2305));
  AOI21X1 g00782(.A0(n2305), .A1(n1790), .B0(n2290), .Y(n2306));
  INVX1   g00783(.A(P1_IR_REG_22__SCAN_IN), .Y(n2307));
  NOR3X1  g00784(.A(P1_IR_REG_21__SCAN_IN), .B(P1_IR_REG_20__SCAN_IN), .C(P1_IR_REG_0__SCAN_IN), .Y(n2308));
  NAND3X1 g00785(.A(n2308), .B(n2173), .C(n1891), .Y(n2309));
  NOR3X1  g00786(.A(n2309), .B(n2269), .C(n2266), .Y(n2310));
  NOR2X1  g00787(.A(n2310), .B(n2307), .Y(n2311));
  INVX1   g00788(.A(P1_IR_REG_19__SCAN_IN), .Y(n2312));
  INVX1   g00789(.A(P1_IR_REG_20__SCAN_IN), .Y(n2313));
  NAND4X1 g00790(.A(n2285), .B(n2313), .C(n2312), .D(n2307), .Y(n2314));
  NOR3X1  g00791(.A(n2314), .B(P1_IR_REG_18__SCAN_IN), .C(P1_IR_REG_17__SCAN_IN), .Y(n2315));
  AOI21X1 g00792(.A0(n2315), .A1(n2175), .B0(n2311), .Y(n2316));
  AOI22X1 g00793(.A0(n1828), .A1(n2316), .B0(n1803), .B1(P1_IR_REG_22__SCAN_IN), .Y(n2317));
  OAI21X1 g00794(.A0(n2306), .A1(P1_STATE_REG_SCAN_IN), .B0(n2317), .Y(P1_U3333));
  INVX1   g00795(.A(P2_DATAO_REG_23__SCAN_IN), .Y(n2319));
  NOR3X1  g00796(.A(n1793), .B(n1792), .C(n2319), .Y(n2320));
  INVX1   g00797(.A(SI_22_), .Y(n2321));
  NOR2X1  g00798(.A(n2303), .B(n2321), .Y(n2322));
  INVX1   g00799(.A(n2292), .Y(n2323));
  INVX1   g00800(.A(n2281), .Y(n2324));
  OAI22X1 g00801(.A0(n2278), .A1(n2277), .B0(SI_21_), .B1(n2324), .Y(n2325));
  AOI22X1 g00802(.A0(n2325), .A1(n2323), .B0(n2321), .B1(n2303), .Y(n2326));
  NOR2X1  g00803(.A(n2326), .B(n2322), .Y(n2327));
  AOI21X1 g00804(.A0(n1789), .A1(n1786), .B0(n2319), .Y(n2328));
  AOI21X1 g00805(.A0(n1837), .A1(P1_DATAO_REG_23__SCAN_IN), .B0(n2328), .Y(n2329));
  XOR2X1  g00806(.A(n2329), .B(SI_23_), .Y(n2330));
  XOR2X1  g00807(.A(n2330), .B(n2327), .Y(n2331));
  AOI21X1 g00808(.A0(n2331), .A1(n1790), .B0(n2320), .Y(n2332));
  NAND2X1 g00809(.A(n2315), .B(n2175), .Y(n2333));
  INVX1   g00810(.A(P1_IR_REG_18__SCAN_IN), .Y(n2334));
  NOR3X1  g00811(.A(P1_IR_REG_22__SCAN_IN), .B(P1_IR_REG_21__SCAN_IN), .C(P1_IR_REG_20__SCAN_IN), .Y(n2335));
  NAND4X1 g00812(.A(n2312), .B(n2334), .C(n2166), .D(n2335), .Y(n2336));
  NAND3X1 g00813(.A(n2242), .B(n2241), .C(n1891), .Y(n2338));
  INVX1   g00814(.A(P1_IR_REG_23__SCAN_IN), .Y(n2339));
  NAND4X1 g00815(.A(n1844), .B(n2339), .C(n2195), .D(n2173), .Y(n2340));
  NOR4X1  g00816(.A(n2338), .B(n2336), .C(n2266), .D(n2340), .Y(n2341));
  AOI21X1 g00817(.A0(n2333), .A1(P1_IR_REG_23__SCAN_IN), .B0(n2341), .Y(n2342));
  AOI22X1 g00818(.A0(n1828), .A1(n2342), .B0(n1803), .B1(P1_IR_REG_23__SCAN_IN), .Y(n2343));
  OAI21X1 g00819(.A0(n2332), .A1(P1_STATE_REG_SCAN_IN), .B0(n2343), .Y(P1_U3332));
  INVX1   g00820(.A(P2_DATAO_REG_24__SCAN_IN), .Y(n2345));
  NOR3X1  g00821(.A(n1793), .B(n1792), .C(n2345), .Y(n2346));
  INVX1   g00822(.A(SI_23_), .Y(n2347));
  NOR2X1  g00823(.A(n2329), .B(n2347), .Y(n2348));
  INVX1   g00824(.A(n2322), .Y(n2349));
  INVX1   g00825(.A(n2303), .Y(n2350));
  OAI22X1 g00826(.A0(n2300), .A1(n2292), .B0(SI_22_), .B1(n2350), .Y(n2351));
  AOI22X1 g00827(.A0(n2351), .A1(n2349), .B0(n2347), .B1(n2329), .Y(n2352));
  NOR2X1  g00828(.A(n2352), .B(n2348), .Y(n2353));
  AOI21X1 g00829(.A0(n1789), .A1(n1786), .B0(n2345), .Y(n2354));
  AOI21X1 g00830(.A0(n1837), .A1(P1_DATAO_REG_24__SCAN_IN), .B0(n2354), .Y(n2355));
  XOR2X1  g00831(.A(n2355), .B(SI_24_), .Y(n2356));
  XOR2X1  g00832(.A(n2356), .B(n2353), .Y(n2357));
  AOI21X1 g00833(.A0(n2357), .A1(n1790), .B0(n2346), .Y(n2358));
  INVX1   g00834(.A(P1_IR_REG_24__SCAN_IN), .Y(n2359));
  NOR2X1  g00835(.A(n2341), .B(n2359), .Y(n2360));
  NOR3X1  g00836(.A(P1_IR_REG_16__SCAN_IN), .B(P1_IR_REG_15__SCAN_IN), .C(P1_IR_REG_14__SCAN_IN), .Y(n2361));
  NOR4X1  g00837(.A(P1_IR_REG_19__SCAN_IN), .B(P1_IR_REG_18__SCAN_IN), .C(P1_IR_REG_17__SCAN_IN), .D(P1_IR_REG_20__SCAN_IN), .Y(n2362));
  NAND4X1 g00838(.A(n2361), .B(n2168), .C(n1844), .D(n2362), .Y(n2363));
  NOR3X1  g00839(.A(P1_IR_REG_23__SCAN_IN), .B(P1_IR_REG_22__SCAN_IN), .C(P1_IR_REG_21__SCAN_IN), .Y(n2364));
  NOR3X1  g00840(.A(P1_IR_REG_24__SCAN_IN), .B(P1_IR_REG_3__SCAN_IN), .C(P1_IR_REG_2__SCAN_IN), .Y(n2365));
  NAND2X1 g00841(.A(n2365), .B(n2364), .Y(n2366));
  NOR3X1  g00842(.A(n2366), .B(n2363), .C(n2338), .Y(n2367));
  NOR2X1  g00843(.A(n2367), .B(n2360), .Y(n2368));
  AOI22X1 g00844(.A0(n1828), .A1(n2368), .B0(n1803), .B1(P1_IR_REG_24__SCAN_IN), .Y(n2369));
  OAI21X1 g00845(.A0(n2358), .A1(P1_STATE_REG_SCAN_IN), .B0(n2369), .Y(P1_U3331));
  INVX1   g00846(.A(P2_DATAO_REG_25__SCAN_IN), .Y(n2371));
  NOR3X1  g00847(.A(n1793), .B(n1792), .C(n2371), .Y(n2372));
  INVX1   g00848(.A(SI_24_), .Y(n2373));
  NOR2X1  g00849(.A(n2355), .B(n2373), .Y(n2374));
  INVX1   g00850(.A(n2348), .Y(n2375));
  INVX1   g00851(.A(n2329), .Y(n2376));
  OAI22X1 g00852(.A0(n2326), .A1(n2322), .B0(SI_23_), .B1(n2376), .Y(n2377));
  AOI22X1 g00853(.A0(n2377), .A1(n2375), .B0(n2373), .B1(n2355), .Y(n2378));
  NOR2X1  g00854(.A(n2378), .B(n2374), .Y(n2379));
  AOI21X1 g00855(.A0(n1789), .A1(n1786), .B0(n2371), .Y(n2380));
  AOI21X1 g00856(.A0(n1837), .A1(P1_DATAO_REG_25__SCAN_IN), .B0(n2380), .Y(n2381));
  XOR2X1  g00857(.A(n2381), .B(SI_25_), .Y(n2382));
  XOR2X1  g00858(.A(n2382), .B(n2379), .Y(n2383));
  AOI21X1 g00859(.A0(n2383), .A1(n1790), .B0(n2372), .Y(n2384));
  INVX1   g00860(.A(P1_IR_REG_25__SCAN_IN), .Y(n2385));
  XOR2X1  g00861(.A(n2367), .B(n2385), .Y(n2386));
  AOI22X1 g00862(.A0(n1828), .A1(n2386), .B0(n1803), .B1(P1_IR_REG_25__SCAN_IN), .Y(n2387));
  OAI21X1 g00863(.A0(n2384), .A1(P1_STATE_REG_SCAN_IN), .B0(n2387), .Y(P1_U3330));
  INVX1   g00864(.A(P2_DATAO_REG_26__SCAN_IN), .Y(n2389));
  NOR3X1  g00865(.A(n1793), .B(n1792), .C(n2389), .Y(n2390));
  INVX1   g00866(.A(SI_25_), .Y(n2391));
  NOR2X1  g00867(.A(n2381), .B(n2391), .Y(n2392));
  INVX1   g00868(.A(n2392), .Y(n2393));
  INVX1   g00869(.A(n2381), .Y(n2394));
  OAI22X1 g00870(.A0(n2378), .A1(n2374), .B0(SI_25_), .B1(n2394), .Y(n2395));
  AOI21X1 g00871(.A0(n1789), .A1(n1786), .B0(n2389), .Y(n2396));
  AOI21X1 g00872(.A0(n1837), .A1(P1_DATAO_REG_26__SCAN_IN), .B0(n2396), .Y(n2397));
  XOR2X1  g00873(.A(n2397), .B(SI_26_), .Y(n2398));
  INVX1   g00874(.A(n2398), .Y(n2399));
  NAND3X1 g00875(.A(n2399), .B(n2395), .C(n2393), .Y(n2400));
  INVX1   g00876(.A(n2374), .Y(n2401));
  INVX1   g00877(.A(n2355), .Y(n2402));
  OAI22X1 g00878(.A0(n2352), .A1(n2348), .B0(SI_24_), .B1(n2402), .Y(n2403));
  AOI22X1 g00879(.A0(n2403), .A1(n2401), .B0(n2391), .B1(n2381), .Y(n2404));
  OAI21X1 g00880(.A0(n2404), .A1(n2392), .B0(n2398), .Y(n2405));
  AOI21X1 g00881(.A0(n2405), .A1(n2400), .B0(n1837), .Y(n2406));
  OAI21X1 g00882(.A0(n2406), .A1(n2390), .B0(P1_U3086), .Y(n2407));
  INVX1   g00883(.A(P1_IR_REG_26__SCAN_IN), .Y(n2408));
  NAND4X1 g00884(.A(n2173), .B(n2385), .C(n2359), .D(n2364), .Y(n2409));
  NOR3X1  g00885(.A(n2409), .B(n2363), .C(n2338), .Y(n2410));
  NOR2X1  g00886(.A(n2410), .B(n2408), .Y(n2411));
  NOR4X1  g00887(.A(P1_IR_REG_18__SCAN_IN), .B(P1_IR_REG_17__SCAN_IN), .C(P1_IR_REG_1__SCAN_IN), .D(P1_IR_REG_19__SCAN_IN), .Y(n2412));
  NAND4X1 g00888(.A(n2361), .B(n2308), .C(n2168), .D(n2412), .Y(n2413));
  NOR4X1  g00889(.A(P1_IR_REG_24__SCAN_IN), .B(P1_IR_REG_23__SCAN_IN), .C(P1_IR_REG_22__SCAN_IN), .D(P1_IR_REG_25__SCAN_IN), .Y(n2414));
  NOR3X1  g00890(.A(P1_IR_REG_26__SCAN_IN), .B(P1_IR_REG_3__SCAN_IN), .C(P1_IR_REG_2__SCAN_IN), .Y(n2415));
  NAND2X1 g00891(.A(n2415), .B(n2414), .Y(n2416));
  NOR3X1  g00892(.A(n2416), .B(n2413), .C(n2338), .Y(n2417));
  NOR2X1  g00893(.A(n2417), .B(n2411), .Y(n2418));
  AOI22X1 g00894(.A0(n1828), .A1(n2418), .B0(n1803), .B1(P1_IR_REG_26__SCAN_IN), .Y(n2419));
  NAND2X1 g00895(.A(n2419), .B(n2407), .Y(P1_U3329));
  INVX1   g00896(.A(P2_DATAO_REG_27__SCAN_IN), .Y(n2421));
  NOR3X1  g00897(.A(n1793), .B(n1792), .C(n2421), .Y(n2422));
  INVX1   g00898(.A(SI_26_), .Y(n2423));
  NOR2X1  g00899(.A(n2397), .B(n2423), .Y(n2424));
  INVX1   g00900(.A(n2424), .Y(n2425));
  INVX1   g00901(.A(n2397), .Y(n2426));
  OAI22X1 g00902(.A0(n2404), .A1(n2392), .B0(SI_26_), .B1(n2426), .Y(n2427));
  AOI21X1 g00903(.A0(n1789), .A1(n1786), .B0(n2421), .Y(n2428));
  AOI21X1 g00904(.A0(n1837), .A1(P1_DATAO_REG_27__SCAN_IN), .B0(n2428), .Y(n2429));
  XOR2X1  g00905(.A(n2429), .B(SI_27_), .Y(n2430));
  INVX1   g00906(.A(n2430), .Y(n2431));
  NAND3X1 g00907(.A(n2431), .B(n2427), .C(n2425), .Y(n2432));
  AOI22X1 g00908(.A0(n2395), .A1(n2393), .B0(n2423), .B1(n2397), .Y(n2433));
  OAI21X1 g00909(.A0(n2433), .A1(n2424), .B0(n2430), .Y(n2434));
  AOI21X1 g00910(.A0(n2434), .A1(n2432), .B0(n1837), .Y(n2435));
  OAI21X1 g00911(.A0(n2435), .A1(n2422), .B0(P1_U3086), .Y(n2436));
  INVX1   g00912(.A(P1_IR_REG_27__SCAN_IN), .Y(n2437));
  XOR2X1  g00913(.A(n2417), .B(n2437), .Y(n2438));
  AOI22X1 g00914(.A0(n1828), .A1(n2438), .B0(n1803), .B1(P1_IR_REG_27__SCAN_IN), .Y(n2439));
  NAND2X1 g00915(.A(n2439), .B(n2436), .Y(P1_U3328));
  INVX1   g00916(.A(P2_DATAO_REG_28__SCAN_IN), .Y(n2441));
  NOR3X1  g00917(.A(n1793), .B(n1792), .C(n2441), .Y(n2442));
  INVX1   g00918(.A(SI_27_), .Y(n2443));
  NOR2X1  g00919(.A(n2429), .B(n2443), .Y(n2444));
  AOI22X1 g00920(.A0(n2427), .A1(n2425), .B0(n2443), .B1(n2429), .Y(n2445));
  NOR2X1  g00921(.A(n2445), .B(n2444), .Y(n2446));
  AOI21X1 g00922(.A0(n1789), .A1(n1786), .B0(n2441), .Y(n2447));
  AOI21X1 g00923(.A0(n1837), .A1(P1_DATAO_REG_28__SCAN_IN), .B0(n2447), .Y(n2448));
  XOR2X1  g00924(.A(n2448), .B(SI_28_), .Y(n2449));
  XOR2X1  g00925(.A(n2449), .B(n2446), .Y(n2450));
  AOI21X1 g00926(.A0(n2450), .A1(n1790), .B0(n2442), .Y(n2451));
  INVX1   g00927(.A(P1_IR_REG_28__SCAN_IN), .Y(n2452));
  NAND2X1 g00928(.A(n2242), .B(n1993), .Y(n2453));
  NAND4X1 g00929(.A(n2437), .B(n2408), .C(n1843), .D(n2414), .Y(n2454));
  NOR3X1  g00930(.A(n2454), .B(n2453), .C(n2413), .Y(n2455));
  NOR2X1  g00931(.A(n2455), .B(n2452), .Y(n2456));
  NOR3X1  g00932(.A(P1_IR_REG_19__SCAN_IN), .B(P1_IR_REG_18__SCAN_IN), .C(P1_IR_REG_17__SCAN_IN), .Y(n2457));
  NAND4X1 g00933(.A(n2361), .B(n2335), .C(n1844), .D(n2457), .Y(n2458));
  NOR4X1  g00934(.A(P1_IR_REG_25__SCAN_IN), .B(P1_IR_REG_24__SCAN_IN), .C(P1_IR_REG_23__SCAN_IN), .D(P1_IR_REG_26__SCAN_IN), .Y(n2459));
  NOR3X1  g00935(.A(P1_IR_REG_28__SCAN_IN), .B(P1_IR_REG_27__SCAN_IN), .C(P1_IR_REG_2__SCAN_IN), .Y(n2460));
  NAND4X1 g00936(.A(n2459), .B(n2242), .C(n1993), .D(n2460), .Y(n2461));
  NOR3X1  g00937(.A(n2461), .B(n2458), .C(n2215), .Y(n2462));
  NOR4X1  g00938(.A(n2456), .B(P1_U3086), .C(n1827), .D(n2462), .Y(n2463));
  AOI21X1 g00939(.A0(n1803), .A1(P1_IR_REG_28__SCAN_IN), .B0(n2463), .Y(n2464));
  OAI21X1 g00940(.A0(n2451), .A1(P1_STATE_REG_SCAN_IN), .B0(n2464), .Y(P1_U3327));
  INVX1   g00941(.A(P2_DATAO_REG_29__SCAN_IN), .Y(n2466));
  NOR3X1  g00942(.A(n1793), .B(n1792), .C(n2466), .Y(n2467));
  INVX1   g00943(.A(SI_28_), .Y(n2468));
  NOR2X1  g00944(.A(n2448), .B(n2468), .Y(n2469));
  INVX1   g00945(.A(n2469), .Y(n2470));
  INVX1   g00946(.A(n2448), .Y(n2471));
  OAI22X1 g00947(.A0(n2445), .A1(n2444), .B0(SI_28_), .B1(n2471), .Y(n2472));
  AOI21X1 g00948(.A0(n1789), .A1(n1786), .B0(n2466), .Y(n2473));
  AOI21X1 g00949(.A0(n1837), .A1(P1_DATAO_REG_29__SCAN_IN), .B0(n2473), .Y(n2474));
  XOR2X1  g00950(.A(n2474), .B(SI_29_), .Y(n2475));
  INVX1   g00951(.A(n2475), .Y(n2476));
  NAND3X1 g00952(.A(n2476), .B(n2472), .C(n2470), .Y(n2477));
  INVX1   g00953(.A(n2444), .Y(n2478));
  INVX1   g00954(.A(n2429), .Y(n2479));
  OAI22X1 g00955(.A0(n2433), .A1(n2424), .B0(SI_27_), .B1(n2479), .Y(n2480));
  AOI22X1 g00956(.A0(n2480), .A1(n2478), .B0(n2468), .B1(n2448), .Y(n2481));
  OAI21X1 g00957(.A0(n2481), .A1(n2469), .B0(n2475), .Y(n2482));
  AOI21X1 g00958(.A0(n2482), .A1(n2477), .B0(n1837), .Y(n2483));
  OAI21X1 g00959(.A0(n2483), .A1(n2467), .B0(P1_U3086), .Y(n2484));
  INVX1   g00960(.A(P1_IR_REG_29__SCAN_IN), .Y(n2485));
  NOR2X1  g00961(.A(n2462), .B(n2485), .Y(n2486));
  NAND3X1 g00962(.A(n2460), .B(n2459), .C(n2485), .Y(n2487));
  NOR4X1  g00963(.A(n2458), .B(n2453), .C(n2215), .D(n2487), .Y(n2488));
  NOR4X1  g00964(.A(n2486), .B(P1_U3086), .C(n1827), .D(n2488), .Y(n2489));
  AOI21X1 g00965(.A0(n1803), .A1(P1_IR_REG_29__SCAN_IN), .B0(n2489), .Y(n2490));
  NAND2X1 g00966(.A(n2490), .B(n2484), .Y(P1_U3326));
  INVX1   g00967(.A(P2_DATAO_REG_30__SCAN_IN), .Y(n2492));
  NOR3X1  g00968(.A(n1793), .B(n1792), .C(n2492), .Y(n2493));
  INVX1   g00969(.A(n2493), .Y(n2494));
  INVX1   g00970(.A(SI_29_), .Y(n2495));
  NOR2X1  g00971(.A(n2474), .B(n2495), .Y(n2496));
  INVX1   g00972(.A(n2496), .Y(n2497));
  NAND2X1 g00973(.A(n2474), .B(n2495), .Y(n2498));
  OAI21X1 g00974(.A0(n2481), .A1(n2469), .B0(n2498), .Y(n2499));
  NAND2X1 g00975(.A(n2499), .B(n2497), .Y(n2500));
  AOI21X1 g00976(.A0(n1789), .A1(n1786), .B0(n2492), .Y(n2501));
  AOI21X1 g00977(.A0(n1837), .A1(P1_DATAO_REG_30__SCAN_IN), .B0(n2501), .Y(n2502));
  XOR2X1  g00978(.A(n2502), .B(SI_30_), .Y(n2503));
  XOR2X1  g00979(.A(n2503), .B(n2500), .Y(n2504));
  OAI21X1 g00980(.A0(n2504), .A1(n1837), .B0(n2494), .Y(n2505));
  INVX1   g00981(.A(n2505), .Y(n2506));
  INVX1   g00982(.A(P1_IR_REG_30__SCAN_IN), .Y(n2507));
  XOR2X1  g00983(.A(n2488), .B(n2507), .Y(n2508));
  AOI22X1 g00984(.A0(n1828), .A1(n2508), .B0(n1803), .B1(P1_IR_REG_30__SCAN_IN), .Y(n2509));
  OAI21X1 g00985(.A0(n2506), .A1(P1_STATE_REG_SCAN_IN), .B0(n2509), .Y(P1_U3325));
  INVX1   g00986(.A(P2_DATAO_REG_31__SCAN_IN), .Y(n2511));
  NOR3X1  g00987(.A(n1793), .B(n1792), .C(n2511), .Y(n2512));
  INVX1   g00988(.A(SI_30_), .Y(n2513));
  AOI21X1 g00989(.A0(n1789), .A1(n1786), .B0(n2511), .Y(n2514));
  AOI21X1 g00990(.A0(n1837), .A1(P1_DATAO_REG_31__SCAN_IN), .B0(n2514), .Y(n2515));
  XOR2X1  g00991(.A(n2515), .B(SI_31_), .Y(n2516));
  AOI21X1 g00992(.A0(n2502), .A1(n2513), .B0(n2516), .Y(n2517));
  INVX1   g00993(.A(n2517), .Y(n2518));
  AOI21X1 g00994(.A0(n2499), .A1(n2497), .B0(n2518), .Y(n2519));
  AOI22X1 g00995(.A0(n2472), .A1(n2470), .B0(n2495), .B1(n2474), .Y(n2520));
  INVX1   g00996(.A(n2516), .Y(n2521));
  NOR2X1  g00997(.A(n2502), .B(n2513), .Y(n2522));
  NOR4X1  g00998(.A(n2521), .B(n2520), .C(n2496), .D(n2522), .Y(n2523));
  NAND3X1 g00999(.A(n2516), .B(n2502), .C(n2513), .Y(n2524));
  INVX1   g01000(.A(n2524), .Y(n2525));
  AOI21X1 g01001(.A0(n2522), .A1(n2521), .B0(n2525), .Y(n2526));
  INVX1   g01002(.A(n2526), .Y(n2527));
  NOR4X1  g01003(.A(n2523), .B(n2519), .C(n1837), .D(n2527), .Y(n2528));
  OAI21X1 g01004(.A0(n2528), .A1(n2512), .B0(P1_U3086), .Y(n2529));
  NAND4X1 g01005(.A(P1_STATE_REG_SCAN_IN), .B(P1_IR_REG_31__SCAN_IN), .C(n2507), .D(n2488), .Y(n2530));
  NAND2X1 g01006(.A(n2530), .B(n2529), .Y(P1_U3324));
  NOR2X1  g01007(.A(P1_IR_REG_31__SCAN_IN), .B(n2408), .Y(n2532));
  AOI21X1 g01008(.A0(n2418), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2532), .Y(n2533));
  NOR2X1  g01009(.A(P1_IR_REG_31__SCAN_IN), .B(n2385), .Y(n2534));
  AOI21X1 g01010(.A0(n2386), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2534), .Y(n2535));
  NOR2X1  g01011(.A(P1_IR_REG_31__SCAN_IN), .B(n2359), .Y(n2536));
  AOI21X1 g01012(.A0(n2368), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2536), .Y(n2537));
  NOR3X1  g01013(.A(n2537), .B(n2535), .C(n2533), .Y(n2538));
  NAND2X1 g01014(.A(n2342), .B(P1_IR_REG_31__SCAN_IN), .Y(n2539));
  OAI21X1 g01015(.A0(P1_IR_REG_31__SCAN_IN), .A1(n2339), .B0(n2539), .Y(n2540));
  INVX1   g01016(.A(P1_B_REG_SCAN_IN), .Y(n2541));
  NAND2X1 g01017(.A(n2386), .B(P1_IR_REG_31__SCAN_IN), .Y(n2542));
  OAI21X1 g01018(.A0(P1_IR_REG_31__SCAN_IN), .A1(n2385), .B0(n2542), .Y(n2543));
  NAND3X1 g01019(.A(n2034), .B(n1991), .C(n1970), .Y(n2544));
  NOR3X1  g01020(.A(n2544), .B(n1945), .C(P1_IR_REG_4__SCAN_IN), .Y(n2545));
  NAND3X1 g01021(.A(n2365), .B(n2364), .C(n2545), .Y(n2546));
  OAI22X1 g01022(.A0(n2363), .A1(n2546), .B0(n2341), .B1(n2359), .Y(n2547));
  INVX1   g01023(.A(n2536), .Y(n2548));
  OAI21X1 g01024(.A0(n2547), .A1(n1827), .B0(n2548), .Y(n2549));
  NOR4X1  g01025(.A(n2543), .B(n2533), .C(n2541), .D(n2549), .Y(n2550));
  NAND3X1 g01026(.A(n2415), .B(n2414), .C(n2545), .Y(n2551));
  OAI22X1 g01027(.A0(n2413), .A1(n2551), .B0(n2410), .B1(n2408), .Y(n2552));
  INVX1   g01028(.A(n2532), .Y(n2553));
  OAI21X1 g01029(.A0(n2552), .A1(n1827), .B0(n2553), .Y(n2554));
  OAI21X1 g01030(.A0(n2537), .A1(P1_B_REG_SCAN_IN), .B0(n2554), .Y(n2555));
  NOR2X1  g01031(.A(n2555), .B(n2550), .Y(n2556));
  NOR4X1  g01032(.A(n2540), .B(n2538), .C(P1_U3086), .D(n2556), .Y(n2557));
  OAI21X1 g01033(.A0(n2543), .A1(n2533), .B0(n2537), .Y(n2558));
  NAND2X1 g01034(.A(n2558), .B(n2557), .Y(n2559));
  NOR3X1  g01035(.A(n2540), .B(n2538), .C(P1_U3086), .Y(n2560));
  INVX1   g01036(.A(n2560), .Y(n2561));
  OAI21X1 g01037(.A0(n2556), .A1(n2561), .B0(P1_D_REG_0__SCAN_IN), .Y(n2562));
  NAND2X1 g01038(.A(n2562), .B(n2559), .Y(P1_U3445));
  INVX1   g01039(.A(P1_D_REG_1__SCAN_IN), .Y(n2564));
  NAND2X1 g01040(.A(n2535), .B(n2533), .Y(n2565));
  NAND2X1 g01041(.A(n2565), .B(n2557), .Y(n2566));
  OAI21X1 g01042(.A0(n2557), .A1(n2564), .B0(n2566), .Y(P1_U3446));
  INVX1   g01043(.A(P1_D_REG_2__SCAN_IN), .Y(n2568));
  NOR2X1  g01044(.A(n2557), .B(n2568), .Y(P1_U3323));
  INVX1   g01045(.A(P1_D_REG_3__SCAN_IN), .Y(n2570));
  NOR2X1  g01046(.A(n2557), .B(n2570), .Y(P1_U3322));
  INVX1   g01047(.A(P1_D_REG_4__SCAN_IN), .Y(n2572));
  NOR2X1  g01048(.A(n2557), .B(n2572), .Y(P1_U3321));
  INVX1   g01049(.A(P1_D_REG_5__SCAN_IN), .Y(n2574));
  NOR2X1  g01050(.A(n2557), .B(n2574), .Y(P1_U3320));
  INVX1   g01051(.A(P1_D_REG_6__SCAN_IN), .Y(n2576));
  NOR2X1  g01052(.A(n2557), .B(n2576), .Y(P1_U3319));
  INVX1   g01053(.A(P1_D_REG_7__SCAN_IN), .Y(n2578));
  NOR2X1  g01054(.A(n2557), .B(n2578), .Y(P1_U3318));
  INVX1   g01055(.A(P1_D_REG_8__SCAN_IN), .Y(n2580));
  NOR2X1  g01056(.A(n2557), .B(n2580), .Y(P1_U3317));
  INVX1   g01057(.A(P1_D_REG_9__SCAN_IN), .Y(n2582));
  NOR2X1  g01058(.A(n2557), .B(n2582), .Y(P1_U3316));
  INVX1   g01059(.A(P1_D_REG_10__SCAN_IN), .Y(n2584));
  NOR2X1  g01060(.A(n2557), .B(n2584), .Y(P1_U3315));
  INVX1   g01061(.A(P1_D_REG_11__SCAN_IN), .Y(n2586));
  NOR2X1  g01062(.A(n2557), .B(n2586), .Y(P1_U3314));
  INVX1   g01063(.A(P1_D_REG_12__SCAN_IN), .Y(n2588));
  NOR2X1  g01064(.A(n2557), .B(n2588), .Y(P1_U3313));
  INVX1   g01065(.A(P1_D_REG_13__SCAN_IN), .Y(n2590));
  NOR2X1  g01066(.A(n2557), .B(n2590), .Y(P1_U3312));
  INVX1   g01067(.A(P1_D_REG_14__SCAN_IN), .Y(n2592));
  NOR2X1  g01068(.A(n2557), .B(n2592), .Y(P1_U3311));
  INVX1   g01069(.A(P1_D_REG_15__SCAN_IN), .Y(n2594));
  NOR2X1  g01070(.A(n2557), .B(n2594), .Y(P1_U3310));
  INVX1   g01071(.A(P1_D_REG_16__SCAN_IN), .Y(n2596));
  NOR2X1  g01072(.A(n2557), .B(n2596), .Y(P1_U3309));
  INVX1   g01073(.A(P1_D_REG_17__SCAN_IN), .Y(n2598));
  NOR2X1  g01074(.A(n2557), .B(n2598), .Y(P1_U3308));
  INVX1   g01075(.A(P1_D_REG_18__SCAN_IN), .Y(n2600));
  NOR2X1  g01076(.A(n2557), .B(n2600), .Y(P1_U3307));
  INVX1   g01077(.A(P1_D_REG_19__SCAN_IN), .Y(n2602));
  NOR2X1  g01078(.A(n2557), .B(n2602), .Y(P1_U3306));
  INVX1   g01079(.A(P1_D_REG_20__SCAN_IN), .Y(n2604));
  NOR2X1  g01080(.A(n2557), .B(n2604), .Y(P1_U3305));
  INVX1   g01081(.A(P1_D_REG_21__SCAN_IN), .Y(n2606));
  NOR2X1  g01082(.A(n2557), .B(n2606), .Y(P1_U3304));
  INVX1   g01083(.A(P1_D_REG_22__SCAN_IN), .Y(n2608));
  NOR2X1  g01084(.A(n2557), .B(n2608), .Y(P1_U3303));
  INVX1   g01085(.A(P1_D_REG_23__SCAN_IN), .Y(n2610));
  NOR2X1  g01086(.A(n2557), .B(n2610), .Y(P1_U3302));
  INVX1   g01087(.A(P1_D_REG_24__SCAN_IN), .Y(n2612));
  NOR2X1  g01088(.A(n2557), .B(n2612), .Y(P1_U3301));
  INVX1   g01089(.A(P1_D_REG_25__SCAN_IN), .Y(n2614));
  NOR2X1  g01090(.A(n2557), .B(n2614), .Y(P1_U3300));
  INVX1   g01091(.A(P1_D_REG_26__SCAN_IN), .Y(n2616));
  NOR2X1  g01092(.A(n2557), .B(n2616), .Y(P1_U3299));
  INVX1   g01093(.A(P1_D_REG_27__SCAN_IN), .Y(n2618));
  NOR2X1  g01094(.A(n2557), .B(n2618), .Y(P1_U3298));
  INVX1   g01095(.A(P1_D_REG_28__SCAN_IN), .Y(n2620));
  NOR2X1  g01096(.A(n2557), .B(n2620), .Y(P1_U3297));
  INVX1   g01097(.A(P1_D_REG_29__SCAN_IN), .Y(n2622));
  NOR2X1  g01098(.A(n2557), .B(n2622), .Y(P1_U3296));
  INVX1   g01099(.A(P1_D_REG_30__SCAN_IN), .Y(n2624));
  NOR2X1  g01100(.A(n2557), .B(n2624), .Y(P1_U3295));
  INVX1   g01101(.A(P1_D_REG_31__SCAN_IN), .Y(n2626));
  NOR2X1  g01102(.A(n2557), .B(n2626), .Y(P1_U3294));
  OAI21X1 g01103(.A0(P1_D_REG_7__SCAN_IN), .A1(P1_D_REG_3__SCAN_IN), .B0(n2556), .Y(n2628));
  OAI21X1 g01104(.A0(P1_D_REG_9__SCAN_IN), .A1(P1_D_REG_8__SCAN_IN), .B0(n2556), .Y(n2629));
  OAI21X1 g01105(.A0(P1_D_REG_10__SCAN_IN), .A1(P1_D_REG_5__SCAN_IN), .B0(n2556), .Y(n2630));
  OAI21X1 g01106(.A0(P1_D_REG_6__SCAN_IN), .A1(P1_D_REG_4__SCAN_IN), .B0(n2556), .Y(n2631));
  NAND4X1 g01107(.A(n2630), .B(n2629), .C(n2628), .D(n2631), .Y(n2632));
  OAI21X1 g01108(.A0(P1_D_REG_28__SCAN_IN), .A1(P1_D_REG_27__SCAN_IN), .B0(n2556), .Y(n2633));
  OAI21X1 g01109(.A0(P1_D_REG_26__SCAN_IN), .A1(P1_D_REG_25__SCAN_IN), .B0(n2556), .Y(n2634));
  OAI21X1 g01110(.A0(P1_D_REG_31__SCAN_IN), .A1(P1_D_REG_30__SCAN_IN), .B0(n2556), .Y(n2635));
  OAI21X1 g01111(.A0(P1_D_REG_29__SCAN_IN), .A1(P1_D_REG_2__SCAN_IN), .B0(n2556), .Y(n2636));
  NAND4X1 g01112(.A(n2635), .B(n2634), .C(n2633), .D(n2636), .Y(n2637));
  OAI21X1 g01113(.A0(P1_D_REG_21__SCAN_IN), .A1(P1_D_REG_20__SCAN_IN), .B0(n2556), .Y(n2638));
  OAI21X1 g01114(.A0(P1_D_REG_19__SCAN_IN), .A1(P1_D_REG_18__SCAN_IN), .B0(n2556), .Y(n2639));
  OAI21X1 g01115(.A0(P1_D_REG_23__SCAN_IN), .A1(P1_D_REG_22__SCAN_IN), .B0(n2556), .Y(n2640));
  NAND3X1 g01116(.A(n2640), .B(n2639), .C(n2638), .Y(n2641));
  OAI21X1 g01117(.A0(P1_D_REG_14__SCAN_IN), .A1(P1_D_REG_12__SCAN_IN), .B0(n2556), .Y(n2642));
  OAI21X1 g01118(.A0(P1_D_REG_13__SCAN_IN), .A1(P1_D_REG_11__SCAN_IN), .B0(n2556), .Y(n2643));
  OAI21X1 g01119(.A0(P1_D_REG_24__SCAN_IN), .A1(P1_D_REG_16__SCAN_IN), .B0(n2556), .Y(n2644));
  OAI21X1 g01120(.A0(P1_D_REG_17__SCAN_IN), .A1(P1_D_REG_15__SCAN_IN), .B0(n2556), .Y(n2645));
  NAND4X1 g01121(.A(n2644), .B(n2643), .C(n2642), .D(n2645), .Y(n2646));
  NOR4X1  g01122(.A(n2641), .B(n2637), .C(n2632), .D(n2646), .Y(n2647));
  INVX1   g01123(.A(n2647), .Y(n2648));
  AOI21X1 g01124(.A0(n2535), .A1(n2533), .B0(n2556), .Y(n2649));
  AOI21X1 g01125(.A0(n2556), .A1(P1_D_REG_1__SCAN_IN), .B0(n2649), .Y(n2650));
  OAI21X1 g01126(.A0(n2310), .A1(n2307), .B0(n2333), .Y(n2651));
  NOR2X1  g01127(.A(P1_IR_REG_31__SCAN_IN), .B(n2307), .Y(n2652));
  INVX1   g01128(.A(n2652), .Y(n2653));
  OAI21X1 g01129(.A0(n2651), .A1(n1827), .B0(n2653), .Y(n2654));
  NOR2X1  g01130(.A(P1_IR_REG_31__SCAN_IN), .B(n2313), .Y(n2655));
  AOI21X1 g01131(.A0(n2271), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2655), .Y(n2656));
  NOR2X1  g01132(.A(P1_IR_REG_31__SCAN_IN), .B(n2285), .Y(n2657));
  AOI21X1 g01133(.A0(n2286), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2657), .Y(n2658));
  AOI21X1 g01134(.A0(n2658), .A1(n2656), .B0(n2654), .Y(n2659));
  AOI21X1 g01135(.A0(n2316), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2652), .Y(n2660));
  NOR4X1  g01136(.A(P1_IR_REG_3__SCAN_IN), .B(P1_IR_REG_2__SCAN_IN), .C(P1_IR_REG_0__SCAN_IN), .D(P1_IR_REG_4__SCAN_IN), .Y(n2661));
  NOR3X1  g01137(.A(P1_IR_REG_15__SCAN_IN), .B(P1_IR_REG_14__SCAN_IN), .C(P1_IR_REG_13__SCAN_IN), .Y(n2662));
  NAND4X1 g01138(.A(n2661), .B(n2214), .C(n2313), .D(n2662), .Y(n2663));
  OAI22X1 g01139(.A0(n2663), .A1(n2269), .B0(n2246), .B1(n2313), .Y(n2664));
  INVX1   g01140(.A(n2655), .Y(n2665));
  OAI21X1 g01141(.A0(n2664), .A1(n1827), .B0(n2665), .Y(n2666));
  NAND2X1 g01142(.A(n2286), .B(P1_IR_REG_31__SCAN_IN), .Y(n2667));
  OAI21X1 g01143(.A0(P1_IR_REG_31__SCAN_IN), .A1(n2285), .B0(n2667), .Y(n2668));
  NOR4X1  g01144(.A(n2218), .B(n2172), .C(n2169), .D(n2220), .Y(n2669));
  OAI21X1 g01145(.A0(n2669), .A1(n2312), .B0(n2265), .Y(n2670));
  NOR2X1  g01146(.A(P1_IR_REG_31__SCAN_IN), .B(n2312), .Y(n2671));
  INVX1   g01147(.A(n2671), .Y(n2672));
  OAI21X1 g01148(.A0(n2670), .A1(n1827), .B0(n2672), .Y(n2673));
  OAI22X1 g01149(.A0(n2668), .A1(n2660), .B0(n2666), .B1(n2673), .Y(n2674));
  OAI21X1 g01150(.A0(n2674), .A1(n2659), .B0(n2650), .Y(n2675));
  NOR2X1  g01151(.A(n2675), .B(n2648), .Y(n2676));
  AOI21X1 g01152(.A0(n2537), .A1(n2533), .B0(n2556), .Y(n2677));
  AOI21X1 g01153(.A0(n2556), .A1(P1_D_REG_0__SCAN_IN), .B0(n2677), .Y(n2678));
  NAND3X1 g01154(.A(n2678), .B(n2676), .C(n2560), .Y(n2679));
  NAND2X1 g01155(.A(n2438), .B(P1_IR_REG_31__SCAN_IN), .Y(n2680));
  OAI21X1 g01156(.A0(P1_IR_REG_31__SCAN_IN), .A1(n2437), .B0(n2680), .Y(n2681));
  NOR3X1  g01157(.A(n2462), .B(n2456), .C(n1827), .Y(n2682));
  NOR2X1  g01158(.A(P1_IR_REG_31__SCAN_IN), .B(n2452), .Y(n2683));
  NOR3X1  g01159(.A(n2683), .B(n2682), .C(n2681), .Y(n2684));
  NOR2X1  g01160(.A(P1_IR_REG_31__SCAN_IN), .B(n2437), .Y(n2685));
  AOI21X1 g01161(.A0(n2438), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2685), .Y(n2686));
  NOR2X1  g01162(.A(n2683), .B(n2682), .Y(n2687));
  INVX1   g01163(.A(n2219), .Y(n2691));
  NAND3X1 g01164(.A(n2691), .B(n2687), .C(n2686), .Y(n2692));
  OAI21X1 g01165(.A0(n2684), .A1(n1801), .B0(n2692), .Y(n2693));
  INVX1   g01166(.A(P1_REG0_REG_0__SCAN_IN), .Y(n2694));
  XOR2X1  g01167(.A(n2488), .B(P1_IR_REG_30__SCAN_IN), .Y(n2695));
  NOR2X1  g01168(.A(P1_IR_REG_31__SCAN_IN), .B(n2507), .Y(n2696));
  INVX1   g01169(.A(n2696), .Y(n2697));
  OAI21X1 g01170(.A0(n2695), .A1(n1827), .B0(n2697), .Y(n2698));
  NOR3X1  g01171(.A(n2488), .B(n2486), .C(n1827), .Y(n2699));
  NOR2X1  g01172(.A(P1_IR_REG_31__SCAN_IN), .B(n2485), .Y(n2700));
  NOR4X1  g01173(.A(n2699), .B(n2698), .C(n2694), .D(n2700), .Y(n2701));
  INVX1   g01174(.A(P1_REG2_REG_0__SCAN_IN), .Y(n2702));
  AOI21X1 g01175(.A0(n2508), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2696), .Y(n2703));
  NOR4X1  g01176(.A(n2699), .B(n2703), .C(n2702), .D(n2700), .Y(n2704));
  INVX1   g01177(.A(P1_REG1_REG_0__SCAN_IN), .Y(n2705));
  INVX1   g01178(.A(P1_REG3_REG_0__SCAN_IN), .Y(n2706));
  OAI21X1 g01179(.A0(n2700), .A1(n2699), .B0(n2703), .Y(n2707));
  OAI21X1 g01180(.A0(n2700), .A1(n2699), .B0(n2698), .Y(n2708));
  OAI22X1 g01181(.A0(n2707), .A1(n2705), .B0(n2706), .B1(n2708), .Y(n2709));
  NOR3X1  g01182(.A(n2709), .B(n2704), .C(n2701), .Y(n2710));
  XOR2X1  g01183(.A(n2710), .B(n2693), .Y(n2711));
  AOI21X1 g01184(.A0(n2247), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2671), .Y(n2713));
  NOR3X1  g01185(.A(n2713), .B(n2666), .C(n2660), .Y(n2714));
  NOR3X1  g01186(.A(n2713), .B(n2658), .C(n2656), .Y(n2715));
  INVX1   g01187(.A(n2715), .Y(n2716));
  NAND3X1 g01188(.A(n2713), .B(n2666), .C(n2654), .Y(n2717));
  AOI21X1 g01189(.A0(n2717), .A1(n2716), .B0(n2711), .Y(n2718));
  AOI21X1 g01190(.A0(n2714), .A1(n5490), .B0(n2718), .Y(n2719));
  NOR3X1  g01191(.A(n2713), .B(n2656), .C(n2660), .Y(n2720));
  NOR3X1  g01192(.A(n2673), .B(n2658), .C(n2656), .Y(n2721));
  OAI21X1 g01193(.A0(n2721), .A1(n2720), .B0(n5490), .Y(n2722));
  NAND4X1 g01194(.A(n2668), .B(n2656), .C(n2660), .D(n2713), .Y(n2723));
  INVX1   g01195(.A(n2723), .Y(n2724));
  NOR4X1  g01196(.A(n2668), .B(n2666), .C(n2660), .D(n2673), .Y(n2725));
  OAI21X1 g01197(.A0(n2725), .A1(n2724), .B0(n5490), .Y(n2726));
  NAND3X1 g01198(.A(n2726), .B(n2722), .C(n2719), .Y(n2727));
  NAND3X1 g01199(.A(n2673), .B(n2656), .C(n2660), .Y(n2728));
  NOR4X1  g01200(.A(n2682), .B(n2658), .C(n2660), .D(n2683), .Y(n2729));
  NOR3X1  g01201(.A(n2700), .B(n2699), .C(n2698), .Y(n2730));
  NOR3X1  g01202(.A(n2700), .B(n2699), .C(n2703), .Y(n2731));
  AOI22X1 g01203(.A0(n2730), .A1(P1_REG0_REG_1__SCAN_IN), .B0(P1_REG2_REG_1__SCAN_IN), .B1(n2731), .Y(n2732));
  NOR2X1  g01204(.A(n2700), .B(n2699), .Y(n2733));
  NOR2X1  g01205(.A(n2733), .B(n2698), .Y(n2734));
  NOR2X1  g01206(.A(n2733), .B(n2703), .Y(n2735));
  AOI22X1 g01207(.A0(n2734), .A1(P1_REG1_REG_1__SCAN_IN), .B0(P1_REG3_REG_1__SCAN_IN), .B1(n2735), .Y(n2736));
  NAND2X1 g01208(.A(n2736), .B(n2732), .Y(n2737));
  AOI21X1 g01209(.A0(n2687), .A1(n2686), .B0(n1801), .Y(n2738));
  AOI21X1 g01210(.A0(n2691), .A1(n2684), .B0(n2738), .Y(n2739));
  NOR3X1  g01211(.A(n2668), .B(n2666), .C(n2654), .Y(n2740));
  INVX1   g01212(.A(n2740), .Y(n2741));
  NOR3X1  g01213(.A(n2713), .B(n2668), .C(n2654), .Y(n2742));
  NOR3X1  g01214(.A(n2673), .B(n2668), .C(n2654), .Y(n2743));
  AOI21X1 g01215(.A0(n2743), .A1(n2666), .B0(n2742), .Y(n2744));
  AOI21X1 g01216(.A0(n2744), .A1(n2741), .B0(n2739), .Y(n2745));
  AOI21X1 g01217(.A0(n2737), .A1(n2729), .B0(n2745), .Y(n2746));
  OAI21X1 g01218(.A0(n2728), .A1(n2711), .B0(n2746), .Y(n2747));
  NOR2X1  g01219(.A(n2747), .B(n2727), .Y(n2748));
  NAND2X1 g01220(.A(n2679), .B(P1_REG0_REG_0__SCAN_IN), .Y(n2749));
  OAI21X1 g01221(.A0(n2748), .A1(n2679), .B0(n2749), .Y(P1_U3459));
  NOR3X1  g01222(.A(n2673), .B(n2656), .C(n2660), .Y(n2751));
  INVX1   g01223(.A(P1_IR_REG_1__SCAN_IN), .Y(n2752));
  NOR2X1  g01224(.A(P1_IR_REG_31__SCAN_IN), .B(n2752), .Y(n2753));
  AOI21X1 g01225(.A0(n1829), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2753), .Y(n2754));
  INVX1   g01226(.A(n2754), .Y(n2755));
  NAND3X1 g01227(.A(n2755), .B(n2687), .C(n2686), .Y(n2756));
  OAI21X1 g01228(.A0(n2684), .A1(n1826), .B0(n2756), .Y(n2757));
  XOR2X1  g01229(.A(n2757), .B(n2737), .Y(n2758));
  NOR2X1  g01230(.A(n2704), .B(n2701), .Y(n2759));
  NOR2X1  g01231(.A(n2458), .B(n2215), .Y(n2760));
  NOR2X1  g01232(.A(n2487), .B(n2453), .Y(n2761));
  NAND2X1 g01233(.A(n2761), .B(n2760), .Y(n2762));
  OAI21X1 g01234(.A0(n2462), .A1(n2485), .B0(n2762), .Y(n2763));
  INVX1   g01235(.A(n2700), .Y(n2764));
  OAI21X1 g01236(.A0(n2763), .A1(n1827), .B0(n2764), .Y(n2765));
  NAND3X1 g01237(.A(n2765), .B(n2703), .C(P1_REG1_REG_0__SCAN_IN), .Y(n2766));
  NAND3X1 g01238(.A(n2765), .B(n2698), .C(P1_REG3_REG_0__SCAN_IN), .Y(n2767));
  NAND3X1 g01239(.A(n2767), .B(n2766), .C(n2759), .Y(n2768));
  NAND2X1 g01240(.A(n2768), .B(n2693), .Y(n2769));
  XOR2X1  g01241(.A(n2769), .B(n2758), .Y(n2770));
  INVX1   g01242(.A(n2770), .Y(n2771));
  OAI21X1 g01243(.A0(n2725), .A1(n2751), .B0(n2771), .Y(n2772));
  NOR2X1  g01244(.A(n2768), .B(n2739), .Y(n2773));
  INVX1   g01245(.A(P1_REG2_REG_1__SCAN_IN), .Y(n2774));
  NAND2X1 g01246(.A(n2733), .B(n2698), .Y(n2775));
  NAND2X1 g01247(.A(n2730), .B(P1_REG0_REG_1__SCAN_IN), .Y(n2776));
  OAI21X1 g01248(.A0(n2775), .A1(n2774), .B0(n2776), .Y(n2777));
  INVX1   g01249(.A(P1_REG1_REG_1__SCAN_IN), .Y(n2778));
  INVX1   g01250(.A(P1_REG3_REG_1__SCAN_IN), .Y(n2779));
  OAI22X1 g01251(.A0(n2707), .A1(n2778), .B0(n2779), .B1(n2708), .Y(n2780));
  NOR2X1  g01252(.A(n2780), .B(n2777), .Y(n2781));
  XOR2X1  g01253(.A(n2757), .B(n2781), .Y(n2782));
  XOR2X1  g01254(.A(n2782), .B(n2773), .Y(n2783));
  INVX1   g01255(.A(n2783), .Y(n2784));
  AOI22X1 g01256(.A0(n2771), .A1(n2724), .B0(n2715), .B1(n2784), .Y(n2785));
  NOR3X1  g01257(.A(n2687), .B(n2658), .C(n2660), .Y(n2786));
  AOI22X1 g01258(.A0(n2784), .A1(n2721), .B0(n2768), .B1(n2786), .Y(n2787));
  OAI21X1 g01259(.A0(n2720), .A1(n2714), .B0(n2784), .Y(n2788));
  NAND4X1 g01260(.A(n2787), .B(n2785), .C(n2772), .D(n2788), .Y(n2789));
  XOR2X1  g01261(.A(n2757), .B(n2693), .Y(n2790));
  INVX1   g01262(.A(n2729), .Y(n2791));
  INVX1   g01263(.A(n2757), .Y(n2792));
  INVX1   g01264(.A(P1_REG2_REG_2__SCAN_IN), .Y(n2793));
  NAND2X1 g01265(.A(n2730), .B(P1_REG0_REG_2__SCAN_IN), .Y(n2794));
  OAI21X1 g01266(.A0(n2775), .A1(n2793), .B0(n2794), .Y(n2795));
  INVX1   g01267(.A(P1_REG1_REG_2__SCAN_IN), .Y(n2796));
  INVX1   g01268(.A(P1_REG3_REG_2__SCAN_IN), .Y(n2797));
  OAI22X1 g01269(.A0(n2707), .A1(n2796), .B0(n2797), .B1(n2708), .Y(n2798));
  NOR2X1  g01270(.A(n2798), .B(n2795), .Y(n2799));
  OAI22X1 g01271(.A0(n2792), .A1(n2744), .B0(n2791), .B1(n2799), .Y(n2800));
  AOI21X1 g01272(.A0(n2790), .A1(n2740), .B0(n2800), .Y(n2801));
  OAI21X1 g01273(.A0(n2770), .A1(n2728), .B0(n2801), .Y(n2802));
  NOR2X1  g01274(.A(n2802), .B(n2789), .Y(n2803));
  NAND2X1 g01275(.A(n2679), .B(P1_REG0_REG_1__SCAN_IN), .Y(n2804));
  OAI21X1 g01276(.A0(n2803), .A1(n2679), .B0(n2804), .Y(P1_U3462));
  INVX1   g01277(.A(n1833), .Y(n2806));
  NAND2X1 g01278(.A(n1874), .B(n1873), .Y(n2807));
  XOR2X1  g01279(.A(n1840), .B(n2807), .Y(n2808));
  OAI21X1 g01280(.A0(n2808), .A1(n1837), .B0(n2806), .Y(n2809));
  NAND2X1 g01281(.A(n2687), .B(n2686), .Y(n2810));
  NOR2X1  g01282(.A(P1_IR_REG_31__SCAN_IN), .B(n1843), .Y(n2811));
  AOI21X1 g01283(.A0(n1845), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2811), .Y(n2812));
  NOR4X1  g01284(.A(n2683), .B(n2682), .C(n2681), .D(n2812), .Y(n2813));
  AOI21X1 g01285(.A0(n2810), .A1(n2809), .B0(n2813), .Y(n2814));
  NOR2X1  g01286(.A(n2814), .B(n2799), .Y(n2815));
  NAND2X1 g01287(.A(n2814), .B(n2799), .Y(n2816));
  INVX1   g01288(.A(n2816), .Y(n2817));
  NOR2X1  g01289(.A(n2792), .B(n2781), .Y(n2818));
  AOI21X1 g01290(.A0(n2792), .A1(n2781), .B0(n2769), .Y(n2819));
  NOR2X1  g01291(.A(n2819), .B(n2818), .Y(n2820));
  NOR3X1  g01292(.A(n2820), .B(n2817), .C(n2815), .Y(n2821));
  AOI22X1 g01293(.A0(n2730), .A1(P1_REG0_REG_2__SCAN_IN), .B0(P1_REG2_REG_2__SCAN_IN), .B1(n2731), .Y(n2822));
  AOI22X1 g01294(.A0(n2734), .A1(P1_REG1_REG_2__SCAN_IN), .B0(P1_REG3_REG_2__SCAN_IN), .B1(n2735), .Y(n2823));
  NAND2X1 g01295(.A(n2823), .B(n2822), .Y(n2824));
  INVX1   g01296(.A(n2812), .Y(n2825));
  NAND3X1 g01297(.A(n2825), .B(n2687), .C(n2686), .Y(n2826));
  OAI21X1 g01298(.A0(n2684), .A1(n1842), .B0(n2826), .Y(n2827));
  XOR2X1  g01299(.A(n2827), .B(n2824), .Y(n2828));
  NOR3X1  g01300(.A(n2828), .B(n2819), .C(n2818), .Y(n2829));
  NOR2X1  g01301(.A(n2829), .B(n2821), .Y(n2830));
  AOI22X1 g01302(.A0(n2786), .A1(n2737), .B0(n2724), .B1(n2830), .Y(n2831));
  OAI21X1 g01303(.A0(n2725), .A1(n2751), .B0(n2830), .Y(n2832));
  AOI22X1 g01304(.A0(n2732), .A1(n2736), .B0(n2710), .B1(n2693), .Y(n2833));
  NAND4X1 g01305(.A(n2732), .B(n2710), .C(n2693), .D(n2736), .Y(n2834));
  AOI21X1 g01306(.A0(n2834), .A1(n2792), .B0(n2833), .Y(n2835));
  XOR2X1  g01307(.A(n2835), .B(n2828), .Y(n2836));
  OAI21X1 g01308(.A0(n2721), .A1(n2720), .B0(n2836), .Y(n2837));
  OAI21X1 g01309(.A0(n2715), .A1(n2714), .B0(n2836), .Y(n2838));
  NAND4X1 g01310(.A(n2837), .B(n2832), .C(n2831), .D(n2838), .Y(n2839));
  NAND4X1 g01311(.A(n2673), .B(n2656), .C(n2660), .D(n2830), .Y(n2840));
  NOR2X1  g01312(.A(n2757), .B(n2693), .Y(n2841));
  XOR2X1  g01313(.A(n2841), .B(n2814), .Y(n2842));
  AOI22X1 g01314(.A0(n2730), .A1(P1_REG0_REG_3__SCAN_IN), .B0(P1_REG2_REG_3__SCAN_IN), .B1(n2731), .Y(n2843));
  INVX1   g01315(.A(n2843), .Y(n2844));
  INVX1   g01316(.A(P1_REG1_REG_3__SCAN_IN), .Y(n2845));
  OAI22X1 g01317(.A0(n2707), .A1(n2845), .B0(P1_REG3_REG_3__SCAN_IN), .B1(n2708), .Y(n2846));
  NOR2X1  g01318(.A(n2846), .B(n2844), .Y(n2847));
  OAI22X1 g01319(.A0(n2814), .A1(n2744), .B0(n2791), .B1(n2847), .Y(n2848));
  AOI21X1 g01320(.A0(n2842), .A1(n2740), .B0(n2848), .Y(n2849));
  NAND2X1 g01321(.A(n2849), .B(n2840), .Y(n2850));
  NOR2X1  g01322(.A(n2850), .B(n2839), .Y(n2851));
  NAND2X1 g01323(.A(n2679), .B(P1_REG0_REG_2__SCAN_IN), .Y(n2852));
  OAI21X1 g01324(.A0(n2851), .A1(n2679), .B0(n2852), .Y(P1_U3465));
  INVX1   g01325(.A(n2786), .Y(n2854));
  AOI21X1 g01326(.A0(n2816), .A1(n2818), .B0(n2815), .Y(n2855));
  NAND2X1 g01327(.A(n2819), .B(n2816), .Y(n2856));
  NAND2X1 g01328(.A(n2856), .B(n2855), .Y(n2857));
  INVX1   g01329(.A(n2846), .Y(n2858));
  NAND2X1 g01330(.A(n2858), .B(n2843), .Y(n2859));
  INVX1   g01331(.A(n1849), .Y(n2860));
  XOR2X1  g01332(.A(n1862), .B(n1859), .Y(n2861));
  OAI21X1 g01333(.A0(n2861), .A1(n1837), .B0(n2860), .Y(n2862));
  NOR2X1  g01334(.A(P1_IR_REG_31__SCAN_IN), .B(n1866), .Y(n2863));
  AOI21X1 g01335(.A0(n1868), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2863), .Y(n2864));
  NOR4X1  g01336(.A(n2683), .B(n2682), .C(n2681), .D(n2864), .Y(n2865));
  AOI21X1 g01337(.A0(n2810), .A1(n2862), .B0(n2865), .Y(n2866));
  XOR2X1  g01338(.A(n2866), .B(n2859), .Y(n2867));
  NOR2X1  g01339(.A(n2867), .B(n2857), .Y(n2868));
  INVX1   g01340(.A(n2865), .Y(n2869));
  OAI21X1 g01341(.A0(n2684), .A1(n1865), .B0(n2869), .Y(n2870));
  XOR2X1  g01342(.A(n2870), .B(n2859), .Y(n2871));
  AOI21X1 g01343(.A0(n2856), .A1(n2855), .B0(n2871), .Y(n2872));
  NOR2X1  g01344(.A(n2872), .B(n2868), .Y(n2873));
  OAI22X1 g01345(.A0(n2799), .A1(n2854), .B0(n2723), .B1(n2873), .Y(n2874));
  INVX1   g01346(.A(n2725), .Y(n2875));
  AOI21X1 g01347(.A0(n2875), .A1(n2717), .B0(n2873), .Y(n2876));
  NOR2X1  g01348(.A(n2814), .B(n2824), .Y(n2877));
  NOR2X1  g01349(.A(n2827), .B(n2799), .Y(n2878));
  NAND2X1 g01350(.A(n2834), .B(n2792), .Y(n2879));
  OAI21X1 g01351(.A0(n2781), .A1(n2773), .B0(n2879), .Y(n2880));
  NOR2X1  g01352(.A(n2880), .B(n2878), .Y(n2881));
  NOR3X1  g01353(.A(n2881), .B(n2867), .C(n2877), .Y(n2882));
  NAND2X1 g01354(.A(n2827), .B(n2799), .Y(n2883));
  NAND2X1 g01355(.A(n2814), .B(n2824), .Y(n2884));
  NAND2X1 g01356(.A(n2867), .B(n2884), .Y(n2885));
  AOI21X1 g01357(.A0(n2880), .A1(n2883), .B0(n2885), .Y(n2886));
  OAI22X1 g01358(.A0(n2882), .A1(n2886), .B0(n2721), .B1(n2720), .Y(n2887));
  OAI22X1 g01359(.A0(n2882), .A1(n2886), .B0(n2715), .B1(n2714), .Y(n2888));
  NAND2X1 g01360(.A(n2888), .B(n2887), .Y(n2889));
  NAND3X1 g01361(.A(n2814), .B(n2792), .C(n2739), .Y(n2890));
  XOR2X1  g01362(.A(n2870), .B(n2890), .Y(n2891));
  AOI22X1 g01363(.A0(n2730), .A1(P1_REG0_REG_4__SCAN_IN), .B0(P1_REG2_REG_4__SCAN_IN), .B1(n2731), .Y(n2892));
  INVX1   g01364(.A(n2892), .Y(n2893));
  INVX1   g01365(.A(P1_REG1_REG_4__SCAN_IN), .Y(n2894));
  INVX1   g01366(.A(P1_REG3_REG_4__SCAN_IN), .Y(n2895));
  XOR2X1  g01367(.A(P1_REG3_REG_3__SCAN_IN), .B(n2895), .Y(n2896));
  OAI22X1 g01368(.A0(n2708), .A1(n2896), .B0(n2707), .B1(n2894), .Y(n2897));
  NOR2X1  g01369(.A(n2897), .B(n2893), .Y(n2898));
  OAI22X1 g01370(.A0(n2866), .A1(n2744), .B0(n2791), .B1(n2898), .Y(n2899));
  AOI21X1 g01371(.A0(n2891), .A1(n2740), .B0(n2899), .Y(n2900));
  OAI21X1 g01372(.A0(n2873), .A1(n2728), .B0(n2900), .Y(n2901));
  NOR4X1  g01373(.A(n2889), .B(n2876), .C(n2874), .D(n2901), .Y(n2902));
  NAND2X1 g01374(.A(n2679), .B(P1_REG0_REG_3__SCAN_IN), .Y(n2903));
  OAI21X1 g01375(.A0(n2902), .A1(n2679), .B0(n2903), .Y(P1_U3468));
  OAI21X1 g01376(.A0(n2870), .A1(n2859), .B0(n2816), .Y(n2905));
  INVX1   g01377(.A(n2905), .Y(n2906));
  NOR2X1  g01378(.A(n2866), .B(n2847), .Y(n2907));
  INVX1   g01379(.A(n2907), .Y(n2908));
  NAND2X1 g01380(.A(n2866), .B(n2847), .Y(n2909));
  INVX1   g01381(.A(n2909), .Y(n2910));
  OAI21X1 g01382(.A0(n2910), .A1(n2855), .B0(n2908), .Y(n2911));
  AOI21X1 g01383(.A0(n2906), .A1(n2819), .B0(n2911), .Y(n2912));
  NOR2X1  g01384(.A(P1_IR_REG_31__SCAN_IN), .B(n1891), .Y(n2914));
  INVX1   g01385(.A(n2914), .Y(n2915));
  OAI21X1 g01386(.A0(n1894), .A1(n1827), .B0(n2915), .Y(n2916));
  INVX1   g01387(.A(n2916), .Y(n2917));
  NOR4X1  g01388(.A(n2683), .B(n2682), .C(n2681), .D(n2917), .Y(n2918));
  INVX1   g01389(.A(n2918), .Y(n2919));
  OAI21X1 g01390(.A0(n2684), .A1(n1890), .B0(n2919), .Y(n2920));
  XOR2X1  g01391(.A(n2920), .B(n2898), .Y(n2921));
  NOR2X1  g01392(.A(n3011), .B(n2921), .Y(n2922));
  AOI21X1 g01393(.A0(n2921), .A1(n3011), .B0(n2922), .Y(n2924));
  AOI21X1 g01394(.A0(n2875), .A1(n2717), .B0(n2924), .Y(n2925));
  AOI21X1 g01395(.A0(n2870), .A1(n2847), .B0(n2877), .Y(n2926));
  NAND2X1 g01396(.A(n2926), .B(n2880), .Y(n2927));
  AOI21X1 g01397(.A0(n2847), .A1(n2884), .B0(n2870), .Y(n2928));
  AOI21X1 g01398(.A0(n2859), .A1(n2878), .B0(n2928), .Y(n2929));
  NAND2X1 g01399(.A(n2929), .B(n2927), .Y(n2930));
  XOR2X1  g01400(.A(n2930), .B(n2921), .Y(n2931));
  NAND2X1 g01401(.A(n2931), .B(n2715), .Y(n2932));
  OAI21X1 g01402(.A0(n2924), .A1(n2723), .B0(n2932), .Y(n2933));
  AOI22X1 g01403(.A0(n2859), .A1(n2786), .B0(n2721), .B1(n2931), .Y(n2934));
  OAI21X1 g01404(.A0(n2720), .A1(n2714), .B0(n2931), .Y(n2935));
  NAND2X1 g01405(.A(n2935), .B(n2934), .Y(n2936));
  NOR2X1  g01406(.A(n2870), .B(n2890), .Y(n2937));
  INVX1   g01407(.A(n2920), .Y(n2938));
  XOR2X1  g01408(.A(n2938), .B(n2937), .Y(n2939));
  AOI22X1 g01409(.A0(n2730), .A1(P1_REG0_REG_5__SCAN_IN), .B0(P1_REG2_REG_5__SCAN_IN), .B1(n2731), .Y(n2940));
  INVX1   g01410(.A(n2940), .Y(n2941));
  INVX1   g01411(.A(P1_REG1_REG_5__SCAN_IN), .Y(n2942));
  NAND2X1 g01412(.A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), .Y(n2943));
  XOR2X1  g01413(.A(n2943), .B(P1_REG3_REG_5__SCAN_IN), .Y(n2944));
  OAI22X1 g01414(.A0(n2708), .A1(n2944), .B0(n2707), .B1(n2942), .Y(n2945));
  NOR2X1  g01415(.A(n2945), .B(n2941), .Y(n2946));
  OAI22X1 g01416(.A0(n2938), .A1(n2744), .B0(n2791), .B1(n2946), .Y(n2947));
  AOI21X1 g01417(.A0(n2939), .A1(n2740), .B0(n2947), .Y(n2948));
  OAI21X1 g01418(.A0(n2924), .A1(n2728), .B0(n2948), .Y(n2949));
  NOR4X1  g01419(.A(n2936), .B(n2933), .C(n2925), .D(n2949), .Y(n2950));
  NAND2X1 g01420(.A(n2679), .B(P1_REG0_REG_4__SCAN_IN), .Y(n2951));
  OAI21X1 g01421(.A0(n2950), .A1(n2679), .B0(n2951), .Y(P1_U3471));
  INVX1   g01422(.A(n2897), .Y(n2953));
  NAND2X1 g01423(.A(n2953), .B(n2892), .Y(n2954));
  XOR2X1  g01424(.A(n1888), .B(n1929), .Y(n2955));
  NOR2X1  g01425(.A(n2955), .B(n1837), .Y(n2956));
  OAI21X1 g01426(.A0(n2956), .A1(n1872), .B0(n2810), .Y(n2957));
  AOI21X1 g01427(.A0(n2957), .A1(n2919), .B0(n2898), .Y(n2958));
  INVX1   g01428(.A(n2945), .Y(n2959));
  NAND2X1 g01429(.A(n2959), .B(n2940), .Y(n2960));
  NOR2X1  g01430(.A(P1_IR_REG_31__SCAN_IN), .B(n1942), .Y(n2961));
  AOI21X1 g01431(.A0(n1924), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2961), .Y(n2962));
  NOR4X1  g01432(.A(n2683), .B(n2682), .C(n2681), .D(n2962), .Y(n2963));
  INVX1   g01433(.A(n2963), .Y(n2964));
  OAI21X1 g01434(.A0(n1922), .A1(n1899), .B0(n2810), .Y(n2965));
  NAND2X1 g01435(.A(n2965), .B(n2964), .Y(n2966));
  NOR2X1  g01436(.A(n1922), .B(n1899), .Y(n2967));
  NOR2X1  g01437(.A(n2684), .B(n2967), .Y(n2968));
  NOR2X1  g01438(.A(n2968), .B(n2963), .Y(n2969));
  AOI22X1 g01439(.A0(n2946), .A1(n2969), .B0(n2938), .B1(n2898), .Y(n2970));
  INVX1   g01440(.A(n2970), .Y(n2971));
  AOI21X1 g01441(.A0(n2966), .A1(n2960), .B0(n2971), .Y(n2972));
  OAI21X1 g01442(.A0(n2958), .A1(n3011), .B0(n2972), .Y(n2973));
  AOI21X1 g01443(.A0(n2938), .A1(n2898), .B0(n2912), .Y(n2974));
  XOR2X1  g01444(.A(n2966), .B(n2946), .Y(n2975));
  OAI21X1 g01445(.A0(n2938), .A1(n2898), .B0(n2975), .Y(n2976));
  OAI21X1 g01446(.A0(n2976), .A1(n2974), .B0(n2973), .Y(n2977));
  INVX1   g01447(.A(n2977), .Y(n2978));
  AOI22X1 g01448(.A0(n2954), .A1(n2786), .B0(n2724), .B1(n2978), .Y(n2979));
  OAI21X1 g01449(.A0(n2725), .A1(n2751), .B0(n2978), .Y(n2980));
  AOI22X1 g01450(.A0(n2927), .A1(n2929), .B0(n2920), .B1(n2898), .Y(n2981));
  AOI21X1 g01451(.A0(n2938), .A1(n2954), .B0(n2981), .Y(n2982));
  XOR2X1  g01452(.A(n2982), .B(n2975), .Y(n2983));
  INVX1   g01453(.A(n2983), .Y(n2984));
  OAI21X1 g01454(.A0(n2721), .A1(n2720), .B0(n2984), .Y(n2985));
  OAI21X1 g01455(.A0(n2715), .A1(n2714), .B0(n2984), .Y(n2986));
  NAND4X1 g01456(.A(n2985), .B(n2980), .C(n2979), .D(n2986), .Y(n2987));
  NOR2X1  g01457(.A(n2977), .B(n2728), .Y(n2988));
  NAND2X1 g01458(.A(n2938), .B(n2937), .Y(n2989));
  XOR2X1  g01459(.A(n2969), .B(n2989), .Y(n2990));
  NOR2X1  g01460(.A(n2990), .B(n2741), .Y(n2991));
  AOI22X1 g01461(.A0(n2730), .A1(P1_REG0_REG_6__SCAN_IN), .B0(P1_REG2_REG_6__SCAN_IN), .B1(n2731), .Y(n2992));
  INVX1   g01462(.A(n2992), .Y(n2993));
  INVX1   g01463(.A(P1_REG1_REG_6__SCAN_IN), .Y(n2994));
  NAND3X1 g01464(.A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_5__SCAN_IN), .C(P1_REG3_REG_4__SCAN_IN), .Y(n2995));
  XOR2X1  g01465(.A(n2995), .B(P1_REG3_REG_6__SCAN_IN), .Y(n2996));
  OAI22X1 g01466(.A0(n2708), .A1(n2996), .B0(n2707), .B1(n2994), .Y(n2997));
  NOR2X1  g01467(.A(n2997), .B(n2993), .Y(n2998));
  OAI22X1 g01468(.A0(n2969), .A1(n2744), .B0(n2791), .B1(n2998), .Y(n2999));
  NOR4X1  g01469(.A(n2991), .B(n2988), .C(n2987), .D(n2999), .Y(n3000));
  NAND2X1 g01470(.A(n2679), .B(P1_REG0_REG_5__SCAN_IN), .Y(n3001));
  OAI21X1 g01471(.A0(n3000), .A1(n2679), .B0(n3001), .Y(P1_U3474));
  NOR2X1  g01472(.A(P1_IR_REG_31__SCAN_IN), .B(n1944), .Y(n3003));
  AOI21X1 g01473(.A0(n1947), .A1(P1_IR_REG_31__SCAN_IN), .B0(n3003), .Y(n3004));
  NOR4X1  g01474(.A(n2683), .B(n2682), .C(n2681), .D(n3004), .Y(n3005));
  INVX1   g01475(.A(n3005), .Y(n3006));
  OAI21X1 g01476(.A0(n2684), .A1(n1941), .B0(n3006), .Y(n3007));
  XOR2X1  g01477(.A(n3007), .B(n2998), .Y(n3008));
  AOI21X1 g01478(.A0(n2909), .A1(n2815), .B0(n2907), .Y(n3010));
  OAI21X1 g01479(.A0(n2905), .A1(n2820), .B0(n3010), .Y(n3011));
  NAND2X1 g01480(.A(n2966), .B(n2958), .Y(n3012));
  OAI21X1 g01481(.A0(n2966), .A1(n2958), .B0(n2960), .Y(n3013));
  NAND2X1 g01482(.A(n3013), .B(n3012), .Y(n3014));
  AOI21X1 g01483(.A0(n3011), .A1(n2970), .B0(n3014), .Y(n3015));
  INVX1   g01484(.A(n2997), .Y(n3016));
  NAND2X1 g01485(.A(n3016), .B(n2992), .Y(n3017));
  XOR2X1  g01486(.A(n3007), .B(n3017), .Y(n3018));
  NOR2X1  g01487(.A(n3018), .B(n3015), .Y(n3019));
  AOI21X1 g01488(.A0(n3015), .A1(n3018), .B0(n3019), .Y(n3020));
  OAI22X1 g01489(.A0(n2946), .A1(n2854), .B0(n2723), .B1(n3020), .Y(n3021));
  AOI21X1 g01490(.A0(n2875), .A1(n2717), .B0(n3020), .Y(n3022));
  NOR2X1  g01491(.A(n2966), .B(n2946), .Y(n3023));
  INVX1   g01492(.A(n2982), .Y(n3024));
  AOI21X1 g01493(.A0(n2965), .A1(n2964), .B0(n2960), .Y(n3025));
  NOR2X1  g01494(.A(n3008), .B(n3025), .Y(n3026));
  OAI21X1 g01495(.A0(n3024), .A1(n3023), .B0(n3026), .Y(n3027));
  INVX1   g01496(.A(n1939), .Y(n3028));
  XOR2X1  g01497(.A(n3028), .B(n1934), .Y(n3029));
  NOR2X1  g01498(.A(n3029), .B(n1837), .Y(n3030));
  OAI21X1 g01499(.A0(n3030), .A1(n1928), .B0(n2810), .Y(n3031));
  AOI21X1 g01500(.A0(n3031), .A1(n3006), .B0(n3017), .Y(n3032));
  OAI22X1 g01501(.A0(n2998), .A1(n3007), .B0(n2966), .B1(n2946), .Y(n3033));
  NOR2X1  g01502(.A(n3033), .B(n3032), .Y(n3034));
  OAI21X1 g01503(.A0(n2982), .A1(n3025), .B0(n3034), .Y(n3035));
  NAND2X1 g01504(.A(n3035), .B(n3027), .Y(n3036));
  OAI21X1 g01505(.A0(n2721), .A1(n2720), .B0(n3036), .Y(n3037));
  OAI21X1 g01506(.A0(n2715), .A1(n2714), .B0(n3036), .Y(n3038));
  NAND2X1 g01507(.A(n3038), .B(n3037), .Y(n3039));
  NOR4X1  g01508(.A(n2920), .B(n2870), .C(n2890), .D(n2966), .Y(n3040));
  NOR2X1  g01509(.A(n2684), .B(n1941), .Y(n3041));
  NOR2X1  g01510(.A(n3041), .B(n3005), .Y(n3042));
  XOR2X1  g01511(.A(n3042), .B(n3040), .Y(n3043));
  AOI22X1 g01512(.A0(n2730), .A1(P1_REG0_REG_7__SCAN_IN), .B0(P1_REG2_REG_7__SCAN_IN), .B1(n2731), .Y(n3044));
  NAND4X1 g01513(.A(P1_REG3_REG_5__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), .C(P1_REG3_REG_6__SCAN_IN), .D(P1_REG3_REG_3__SCAN_IN), .Y(n3045));
  XOR2X1  g01514(.A(n3045), .B(P1_REG3_REG_7__SCAN_IN), .Y(n3046));
  INVX1   g01515(.A(n3046), .Y(n3047));
  AOI22X1 g01516(.A0(n2735), .A1(n3047), .B0(n2734), .B1(P1_REG1_REG_7__SCAN_IN), .Y(n3048));
  NAND2X1 g01517(.A(n3048), .B(n3044), .Y(n3049));
  INVX1   g01518(.A(n3049), .Y(n3050));
  OAI22X1 g01519(.A0(n3042), .A1(n2744), .B0(n2791), .B1(n3050), .Y(n3051));
  AOI21X1 g01520(.A0(n3043), .A1(n2740), .B0(n3051), .Y(n3052));
  OAI21X1 g01521(.A0(n3020), .A1(n2728), .B0(n3052), .Y(n3053));
  NOR4X1  g01522(.A(n3039), .B(n3022), .C(n3021), .D(n3053), .Y(n3054));
  NAND2X1 g01523(.A(n2679), .B(P1_REG0_REG_6__SCAN_IN), .Y(n3055));
  OAI21X1 g01524(.A0(n3054), .A1(n2679), .B0(n3055), .Y(P1_U3477));
  INVX1   g01525(.A(n3015), .Y(n3057));
  AOI21X1 g01526(.A0(n3031), .A1(n3006), .B0(n2998), .Y(n3058));
  NOR2X1  g01527(.A(n3058), .B(n3057), .Y(n3059));
  NOR2X1  g01528(.A(P1_IR_REG_31__SCAN_IN), .B(n1970), .Y(n3060));
  AOI21X1 g01529(.A0(n1971), .A1(P1_IR_REG_31__SCAN_IN), .B0(n3060), .Y(n3061));
  INVX1   g01530(.A(n3061), .Y(n3062));
  NOR2X1  g01531(.A(n2684), .B(n1969), .Y(n3063));
  AOI21X1 g01532(.A0(n3062), .A1(n2684), .B0(n3063), .Y(n3064));
  NOR2X1  g01533(.A(n3064), .B(n3050), .Y(n3065));
  NAND3X1 g01534(.A(n3062), .B(n2687), .C(n2686), .Y(n3066));
  OAI21X1 g01535(.A0(n2684), .A1(n1969), .B0(n3066), .Y(n3067));
  OAI22X1 g01536(.A0(n3049), .A1(n3067), .B0(n3007), .B1(n3017), .Y(n3068));
  NOR3X1  g01537(.A(n3068), .B(n3065), .C(n3059), .Y(n3069));
  OAI21X1 g01538(.A0(n3007), .A1(n3017), .B0(n3057), .Y(n3070));
  XOR2X1  g01539(.A(n3067), .B(n3050), .Y(n3071));
  INVX1   g01540(.A(n3071), .Y(n3072));
  NOR2X1  g01541(.A(n3072), .B(n3058), .Y(n3073));
  AOI21X1 g01542(.A0(n3073), .A1(n3070), .B0(n3069), .Y(n3074));
  INVX1   g01543(.A(n3074), .Y(n3075));
  OAI22X1 g01544(.A0(n2998), .A1(n2854), .B0(n2723), .B1(n3075), .Y(n3076));
  AOI21X1 g01545(.A0(n2875), .A1(n2717), .B0(n3075), .Y(n3077));
  AOI22X1 g01546(.A0(n3017), .A1(n3042), .B0(n2969), .B1(n2960), .Y(n3078));
  AOI21X1 g01547(.A0(n3007), .A1(n2998), .B0(n3025), .Y(n3079));
  NAND3X1 g01548(.A(n3079), .B(n2938), .C(n2954), .Y(n3080));
  AOI21X1 g01549(.A0(n3080), .A1(n3078), .B0(n3032), .Y(n3081));
  OAI21X1 g01550(.A0(n2866), .A1(n2859), .B0(n2883), .Y(n3082));
  NOR2X1  g01551(.A(n3082), .B(n2835), .Y(n3083));
  OAI21X1 g01552(.A0(n2859), .A1(n2878), .B0(n2866), .Y(n3084));
  OAI21X1 g01553(.A0(n2847), .A1(n2884), .B0(n3084), .Y(n3085));
  OAI22X1 g01554(.A0(n3083), .A1(n3085), .B0(n2938), .B1(n2954), .Y(n3086));
  NOR3X1  g01555(.A(n3032), .B(n3086), .C(n3025), .Y(n3087));
  NOR2X1  g01556(.A(n3087), .B(n3081), .Y(n3088));
  XOR2X1  g01557(.A(n3088), .B(n3071), .Y(n3089));
  INVX1   g01558(.A(n3089), .Y(n3090));
  OAI21X1 g01559(.A0(n2721), .A1(n2720), .B0(n3090), .Y(n3091));
  OAI21X1 g01560(.A0(n2715), .A1(n2714), .B0(n3090), .Y(n3092));
  NAND2X1 g01561(.A(n3092), .B(n3091), .Y(n3093));
  NAND2X1 g01562(.A(n3042), .B(n3040), .Y(n3094));
  XOR2X1  g01563(.A(n3067), .B(n3094), .Y(n3095));
  AOI22X1 g01564(.A0(n2730), .A1(P1_REG0_REG_8__SCAN_IN), .B0(P1_REG2_REG_8__SCAN_IN), .B1(n2731), .Y(n3096));
  INVX1   g01565(.A(P1_REG3_REG_8__SCAN_IN), .Y(n3097));
  INVX1   g01566(.A(P1_REG3_REG_7__SCAN_IN), .Y(n3098));
  NOR2X1  g01567(.A(n3045), .B(n3098), .Y(n3099));
  XOR2X1  g01568(.A(n3099), .B(n3097), .Y(n3100));
  INVX1   g01569(.A(n3100), .Y(n3101));
  AOI22X1 g01570(.A0(n2735), .A1(n3101), .B0(n2734), .B1(P1_REG1_REG_8__SCAN_IN), .Y(n3102));
  NAND2X1 g01571(.A(n3102), .B(n3096), .Y(n3103));
  INVX1   g01572(.A(n3103), .Y(n3104));
  OAI22X1 g01573(.A0(n3064), .A1(n2744), .B0(n2791), .B1(n3104), .Y(n3105));
  AOI21X1 g01574(.A0(n3095), .A1(n2740), .B0(n3105), .Y(n3106));
  OAI21X1 g01575(.A0(n3075), .A1(n2728), .B0(n3106), .Y(n3107));
  NOR4X1  g01576(.A(n3093), .B(n3077), .C(n3076), .D(n3107), .Y(n3108));
  NAND2X1 g01577(.A(n2679), .B(P1_REG0_REG_7__SCAN_IN), .Y(n3109));
  OAI21X1 g01578(.A0(n3108), .A1(n2679), .B0(n3109), .Y(P1_U3480));
  NOR3X1  g01579(.A(n3064), .B(n3042), .C(n2998), .Y(n3111));
  OAI21X1 g01580(.A0(n3042), .A1(n2998), .B0(n3064), .Y(n3112));
  AOI21X1 g01581(.A0(n3112), .A1(n3049), .B0(n3111), .Y(n3113));
  OAI21X1 g01582(.A0(n3068), .A1(n3015), .B0(n3113), .Y(n3114));
  INVX1   g01583(.A(n3114), .Y(n3115));
  NOR2X1  g01584(.A(P1_IR_REG_31__SCAN_IN), .B(n1991), .Y(n3116));
  AOI21X1 g01585(.A0(n1996), .A1(P1_IR_REG_31__SCAN_IN), .B0(n3116), .Y(n3117));
  NOR4X1  g01586(.A(n2683), .B(n2682), .C(n2681), .D(n3117), .Y(n3118));
  INVX1   g01587(.A(n3118), .Y(n3119));
  OAI21X1 g01588(.A0(n2684), .A1(n1990), .B0(n3119), .Y(n3120));
  XOR2X1  g01589(.A(n3120), .B(n3104), .Y(n3121));
  XOR2X1  g01590(.A(n3120), .B(n3103), .Y(n3123));
  NOR2X1  g01591(.A(n3123), .B(n3115), .Y(n3124));
  AOI21X1 g01592(.A0(n3123), .A1(n3115), .B0(n3124), .Y(n3125));
  OAI22X1 g01593(.A0(n3050), .A1(n2854), .B0(n2723), .B1(n3125), .Y(n3126));
  AOI21X1 g01594(.A0(n2875), .A1(n2717), .B0(n3125), .Y(n3127));
  NAND2X1 g01595(.A(n3064), .B(n3049), .Y(n3128));
  AOI21X1 g01596(.A0(n3067), .A1(n3050), .B0(n3121), .Y(n3129));
  INVX1   g01597(.A(n3129), .Y(n3130));
  AOI21X1 g01598(.A0(n3088), .A1(n3128), .B0(n3130), .Y(n3131));
  NOR2X1  g01599(.A(n3067), .B(n3050), .Y(n3132));
  NOR4X1  g01600(.A(n3025), .B(n2920), .C(n2898), .D(n3032), .Y(n3133));
  OAI22X1 g01601(.A0(n3033), .A1(n3133), .B0(n3042), .B1(n3017), .Y(n3134));
  NAND2X1 g01602(.A(n3079), .B(n2981), .Y(n3135));
  AOI22X1 g01603(.A0(n3134), .A1(n3135), .B0(n3067), .B1(n3050), .Y(n3136));
  NOR3X1  g01604(.A(n3136), .B(n3123), .C(n3132), .Y(n3137));
  OAI22X1 g01605(.A0(n3131), .A1(n3137), .B0(n2721), .B1(n2720), .Y(n3138));
  OAI22X1 g01606(.A0(n3131), .A1(n3137), .B0(n2715), .B1(n2714), .Y(n3139));
  NAND2X1 g01607(.A(n3139), .B(n3138), .Y(n3140));
  NOR4X1  g01608(.A(n3007), .B(n2966), .C(n2989), .D(n3067), .Y(n3141));
  NOR2X1  g01609(.A(n2684), .B(n1990), .Y(n3142));
  NOR2X1  g01610(.A(n3142), .B(n3118), .Y(n3143));
  XOR2X1  g01611(.A(n3143), .B(n3141), .Y(n3144));
  INVX1   g01612(.A(P1_REG3_REG_9__SCAN_IN), .Y(n3145));
  NOR3X1  g01613(.A(n3045), .B(n3098), .C(n3097), .Y(n3146));
  XOR2X1  g01614(.A(n3146), .B(n3145), .Y(n3147));
  INVX1   g01615(.A(n3147), .Y(n3148));
  AOI22X1 g01616(.A0(n2735), .A1(n3148), .B0(n2730), .B1(P1_REG0_REG_9__SCAN_IN), .Y(n3149));
  INVX1   g01617(.A(n3149), .Y(n3150));
  AOI22X1 g01618(.A0(n2731), .A1(P1_REG2_REG_9__SCAN_IN), .B0(P1_REG1_REG_9__SCAN_IN), .B1(n2734), .Y(n3151));
  INVX1   g01619(.A(n3151), .Y(n3152));
  NOR2X1  g01620(.A(n3152), .B(n3150), .Y(n3153));
  OAI22X1 g01621(.A0(n3143), .A1(n2744), .B0(n2791), .B1(n3153), .Y(n3154));
  AOI21X1 g01622(.A0(n3144), .A1(n2740), .B0(n3154), .Y(n3155));
  OAI21X1 g01623(.A0(n3125), .A1(n2728), .B0(n3155), .Y(n3156));
  NOR4X1  g01624(.A(n3140), .B(n3127), .C(n3126), .D(n3156), .Y(n3157));
  NAND2X1 g01625(.A(n2679), .B(P1_REG0_REG_8__SCAN_IN), .Y(n3158));
  OAI21X1 g01626(.A0(n3157), .A1(n2679), .B0(n3158), .Y(P1_U3483));
  NOR2X1  g01627(.A(n3120), .B(n3103), .Y(n3160));
  NAND2X1 g01628(.A(n3120), .B(n3103), .Y(n3161));
  OAI21X1 g01629(.A0(n3160), .A1(n3115), .B0(n3161), .Y(n3162));
  NOR2X1  g01630(.A(P1_IR_REG_31__SCAN_IN), .B(n2034), .Y(n3163));
  AOI21X1 g01631(.A0(n2015), .A1(P1_IR_REG_31__SCAN_IN), .B0(n3163), .Y(n3164));
  INVX1   g01632(.A(n3164), .Y(n3165));
  NAND3X1 g01633(.A(n3165), .B(n2687), .C(n2686), .Y(n3166));
  OAI21X1 g01634(.A0(n2684), .A1(n2014), .B0(n3166), .Y(n3167));
  XOR2X1  g01635(.A(n3167), .B(n3153), .Y(n3168));
  NOR2X1  g01636(.A(n3162), .B(n3168), .Y(n3169));
  INVX1   g01637(.A(n3153), .Y(n3170));
  XOR2X1  g01638(.A(n3167), .B(n3170), .Y(n3171));
  AOI21X1 g01639(.A0(n3168), .A1(n3162), .B0(n3169), .Y(n3173));
  INVX1   g01640(.A(n3173), .Y(n3174));
  OAI21X1 g01641(.A0(n2725), .A1(n2751), .B0(n3174), .Y(n3175));
  OAI22X1 g01642(.A0(n3103), .A1(n3143), .B0(n3064), .B1(n3049), .Y(n3176));
  AOI21X1 g01643(.A0(n3135), .A1(n3134), .B0(n3176), .Y(n3177));
  OAI21X1 g01644(.A0(n3103), .A1(n3132), .B0(n3143), .Y(n3178));
  OAI21X1 g01645(.A0(n3104), .A1(n3128), .B0(n3178), .Y(n3179));
  NOR2X1  g01646(.A(n3179), .B(n3177), .Y(n3180));
  XOR2X1  g01647(.A(n3180), .B(n3168), .Y(n3181));
  INVX1   g01648(.A(n3181), .Y(n3182));
  AOI22X1 g01649(.A0(n3174), .A1(n2724), .B0(n2715), .B1(n3182), .Y(n3183));
  AOI22X1 g01650(.A0(n3103), .A1(n2786), .B0(n2721), .B1(n3182), .Y(n3184));
  OAI21X1 g01651(.A0(n2720), .A1(n2714), .B0(n3182), .Y(n3185));
  NAND4X1 g01652(.A(n3184), .B(n3183), .C(n3175), .D(n3185), .Y(n3186));
  NAND2X1 g01653(.A(n3143), .B(n3141), .Y(n3187));
  XOR2X1  g01654(.A(n3167), .B(n3187), .Y(n3188));
  NOR2X1  g01655(.A(n2684), .B(n2014), .Y(n3189));
  AOI21X1 g01656(.A0(n3165), .A1(n2684), .B0(n3189), .Y(n3190));
  INVX1   g01657(.A(P1_REG3_REG_10__SCAN_IN), .Y(n3191));
  NOR4X1  g01658(.A(n3098), .B(n3097), .C(n3145), .D(n3045), .Y(n3192));
  XOR2X1  g01659(.A(n3192), .B(n3191), .Y(n3193));
  INVX1   g01660(.A(n3193), .Y(n3194));
  AOI22X1 g01661(.A0(n2735), .A1(n3194), .B0(n2730), .B1(P1_REG0_REG_10__SCAN_IN), .Y(n3195));
  INVX1   g01662(.A(n3195), .Y(n3196));
  AOI22X1 g01663(.A0(n2731), .A1(P1_REG2_REG_10__SCAN_IN), .B0(P1_REG1_REG_10__SCAN_IN), .B1(n2734), .Y(n3197));
  INVX1   g01664(.A(n3197), .Y(n3198));
  NOR2X1  g01665(.A(n3198), .B(n3196), .Y(n3199));
  OAI22X1 g01666(.A0(n3190), .A1(n2744), .B0(n2791), .B1(n3199), .Y(n3200));
  AOI21X1 g01667(.A0(n3188), .A1(n2740), .B0(n3200), .Y(n3201));
  OAI21X1 g01668(.A0(n3173), .A1(n2728), .B0(n3201), .Y(n3202));
  NOR2X1  g01669(.A(n3202), .B(n3186), .Y(n3203));
  NAND2X1 g01670(.A(n2679), .B(P1_REG0_REG_9__SCAN_IN), .Y(n3204));
  OAI21X1 g01671(.A0(n3203), .A1(n2679), .B0(n3204), .Y(P1_U3486));
  AOI21X1 g01672(.A0(n3167), .A1(n3170), .B0(n3162), .Y(n3206));
  NOR2X1  g01673(.A(P1_IR_REG_31__SCAN_IN), .B(n2035), .Y(n3207));
  AOI21X1 g01674(.A0(n2040), .A1(P1_IR_REG_31__SCAN_IN), .B0(n3207), .Y(n3208));
  INVX1   g01675(.A(n3208), .Y(n3209));
  NOR2X1  g01676(.A(n2684), .B(n2033), .Y(n3210));
  AOI21X1 g01677(.A0(n3209), .A1(n2684), .B0(n3210), .Y(n3211));
  NOR2X1  g01678(.A(n3211), .B(n3199), .Y(n3212));
  INVX1   g01679(.A(n3199), .Y(n3213));
  NAND2X1 g01680(.A(n3209), .B(n2684), .Y(n3214));
  OAI21X1 g01681(.A0(n2684), .A1(n2033), .B0(n3214), .Y(n3215));
  OAI22X1 g01682(.A0(n3213), .A1(n3215), .B0(n3167), .B1(n3170), .Y(n3216));
  NOR3X1  g01683(.A(n3216), .B(n3212), .C(n3206), .Y(n3217));
  OAI21X1 g01684(.A0(n3167), .A1(n3170), .B0(n3162), .Y(n3218));
  AOI21X1 g01685(.A0(n3167), .A1(n3170), .B0(n5495), .Y(n3221));
  AOI21X1 g01686(.A0(n3221), .A1(n3218), .B0(n3217), .Y(n3222));
  INVX1   g01687(.A(n3222), .Y(n3223));
  OAI22X1 g01688(.A0(n3153), .A1(n2854), .B0(n2723), .B1(n3223), .Y(n3224));
  AOI21X1 g01689(.A0(n2875), .A1(n2717), .B0(n3223), .Y(n3225));
  NOR2X1  g01690(.A(n3190), .B(n3170), .Y(n3226));
  NAND2X1 g01691(.A(n3190), .B(n3170), .Y(n3227));
  OAI21X1 g01692(.A0(n3180), .A1(n3226), .B0(n3227), .Y(n3228));
  XOR2X1  g01693(.A(n3228), .B(n5495), .Y(n3229));
  INVX1   g01694(.A(n3229), .Y(n3230));
  OAI21X1 g01695(.A0(n2721), .A1(n2720), .B0(n3230), .Y(n3231));
  OAI21X1 g01696(.A0(n2715), .A1(n2714), .B0(n3230), .Y(n3232));
  NAND2X1 g01697(.A(n3232), .B(n3231), .Y(n3233));
  NOR4X1  g01698(.A(n3120), .B(n3067), .C(n3094), .D(n3167), .Y(n3234));
  NOR2X1  g01699(.A(n3211), .B(n3234), .Y(n3235));
  NOR3X1  g01700(.A(n3215), .B(n3167), .C(n3187), .Y(n3236));
  NOR2X1  g01701(.A(n3236), .B(n3235), .Y(n3237));
  NAND2X1 g01702(.A(n3192), .B(P1_REG3_REG_10__SCAN_IN), .Y(n3238));
  XOR2X1  g01703(.A(n3238), .B(P1_REG3_REG_11__SCAN_IN), .Y(n3239));
  INVX1   g01704(.A(n3239), .Y(n3240));
  AOI22X1 g01705(.A0(n2735), .A1(n3240), .B0(n2730), .B1(P1_REG0_REG_11__SCAN_IN), .Y(n3241));
  INVX1   g01706(.A(n3241), .Y(n3242));
  AOI22X1 g01707(.A0(n2731), .A1(P1_REG2_REG_11__SCAN_IN), .B0(P1_REG1_REG_11__SCAN_IN), .B1(n2734), .Y(n3243));
  INVX1   g01708(.A(n3243), .Y(n3244));
  NOR2X1  g01709(.A(n3244), .B(n3242), .Y(n3245));
  OAI22X1 g01710(.A0(n3211), .A1(n2744), .B0(n2791), .B1(n3245), .Y(n3246));
  AOI21X1 g01711(.A0(n3237), .A1(n2740), .B0(n3246), .Y(n3247));
  OAI21X1 g01712(.A0(n3223), .A1(n2728), .B0(n3247), .Y(n3248));
  NOR4X1  g01713(.A(n3233), .B(n3225), .C(n3224), .D(n3248), .Y(n3249));
  NAND2X1 g01714(.A(n2679), .B(P1_REG0_REG_10__SCAN_IN), .Y(n3250));
  OAI21X1 g01715(.A0(n3249), .A1(n2679), .B0(n3250), .Y(P1_U3489));
  INVX1   g01716(.A(n2721), .Y(n3252));
  NOR2X1  g01717(.A(n3211), .B(n3213), .Y(n3253));
  AOI21X1 g01718(.A0(n3211), .A1(n3213), .B0(n3228), .Y(n3254));
  NOR2X1  g01719(.A(P1_IR_REG_31__SCAN_IN), .B(n2061), .Y(n3255));
  AOI21X1 g01720(.A0(n2062), .A1(P1_IR_REG_31__SCAN_IN), .B0(n3255), .Y(n3256));
  INVX1   g01721(.A(n3256), .Y(n3257));
  NAND3X1 g01722(.A(n3257), .B(n2687), .C(n2686), .Y(n3258));
  OAI21X1 g01723(.A0(n2684), .A1(n2060), .B0(n3258), .Y(n3259));
  XOR2X1  g01724(.A(n3259), .B(n3245), .Y(n3260));
  NOR3X1  g01725(.A(n3260), .B(n3254), .C(n3253), .Y(n3261));
  NAND2X1 g01726(.A(n3215), .B(n3199), .Y(n3262));
  NAND2X1 g01727(.A(n3228), .B(n3262), .Y(n3263));
  NAND2X1 g01728(.A(n3259), .B(n3245), .Y(n3264));
  INVX1   g01729(.A(n3264), .Y(n3265));
  INVX1   g01730(.A(n3245), .Y(n3266));
  NOR2X1  g01731(.A(n2684), .B(n2060), .Y(n3267));
  AOI21X1 g01732(.A0(n3257), .A1(n2684), .B0(n3267), .Y(n3268));
  AOI22X1 g01733(.A0(n3266), .A1(n3268), .B0(n3211), .B1(n3213), .Y(n3269));
  INVX1   g01734(.A(n3269), .Y(n3270));
  NOR2X1  g01735(.A(n3270), .B(n3265), .Y(n3271));
  AOI21X1 g01736(.A0(n3271), .A1(n3263), .B0(n3261), .Y(n3272));
  NAND2X1 g01737(.A(n3211), .B(n3199), .Y(n3274));
  AOI22X1 g01738(.A0(n3213), .A1(n3215), .B0(n3167), .B1(n3170), .Y(n3275));
  OAI21X1 g01739(.A0(n3216), .A1(n3161), .B0(n3275), .Y(n3276));
  NOR2X1  g01740(.A(n3216), .B(n3160), .Y(n3277));
  AOI22X1 g01741(.A0(n3276), .A1(n3274), .B0(n3114), .B1(n3277), .Y(n3278));
  XOR2X1  g01742(.A(n3259), .B(n3266), .Y(n3279));
  NOR2X1  g01743(.A(n3279), .B(n3278), .Y(n3280));
  AOI21X1 g01744(.A0(n3278), .A1(n3279), .B0(n3280), .Y(n3281));
  OAI22X1 g01745(.A0(n3199), .A1(n2854), .B0(n2723), .B1(n3281), .Y(n3282));
  NOR2X1  g01746(.A(n3281), .B(n2875), .Y(n3283));
  NOR2X1  g01747(.A(n3281), .B(n2717), .Y(n3284));
  NOR3X1  g01748(.A(n3284), .B(n3283), .C(n3282), .Y(n3285));
  OAI21X1 g01749(.A0(n3272), .A1(n3252), .B0(n3285), .Y(n3286));
  NOR2X1  g01750(.A(n3272), .B(n2716), .Y(n3287));
  INVX1   g01751(.A(n2714), .Y(n3288));
  NAND3X1 g01752(.A(n2673), .B(n2666), .C(n2654), .Y(n3289));
  AOI21X1 g01753(.A0(n3289), .A1(n3288), .B0(n3272), .Y(n3290));
  XOR2X1  g01754(.A(n3268), .B(n3236), .Y(n3291));
  NAND3X1 g01755(.A(n3192), .B(P1_REG3_REG_10__SCAN_IN), .C(P1_REG3_REG_11__SCAN_IN), .Y(n3292));
  XOR2X1  g01756(.A(n3292), .B(P1_REG3_REG_12__SCAN_IN), .Y(n3293));
  INVX1   g01757(.A(n3293), .Y(n3294));
  AOI22X1 g01758(.A0(n2735), .A1(n3294), .B0(n2730), .B1(P1_REG0_REG_12__SCAN_IN), .Y(n3295));
  INVX1   g01759(.A(n3295), .Y(n3296));
  AOI22X1 g01760(.A0(n2731), .A1(P1_REG2_REG_12__SCAN_IN), .B0(P1_REG1_REG_12__SCAN_IN), .B1(n2734), .Y(n3297));
  INVX1   g01761(.A(n3297), .Y(n3298));
  NOR2X1  g01762(.A(n3298), .B(n3296), .Y(n3299));
  OAI22X1 g01763(.A0(n3268), .A1(n2744), .B0(n2791), .B1(n3299), .Y(n3300));
  AOI21X1 g01764(.A0(n3291), .A1(n2740), .B0(n3300), .Y(n3301));
  OAI21X1 g01765(.A0(n3281), .A1(n2728), .B0(n3301), .Y(n3302));
  NOR4X1  g01766(.A(n3290), .B(n3287), .C(n3286), .D(n3302), .Y(n3303));
  NAND2X1 g01767(.A(n2679), .B(P1_REG0_REG_11__SCAN_IN), .Y(n3304));
  OAI21X1 g01768(.A0(n3303), .A1(n2679), .B0(n3304), .Y(P1_U3492));
  AOI21X1 g01769(.A0(n3268), .A1(n3245), .B0(n3278), .Y(n3306));
  AOI21X1 g01770(.A0(n3259), .A1(n3266), .B0(n3306), .Y(n3307));
  INVX1   g01771(.A(n3307), .Y(n3308));
  NOR2X1  g01772(.A(P1_IR_REG_31__SCAN_IN), .B(n2082), .Y(n3309));
  AOI21X1 g01773(.A0(n2085), .A1(P1_IR_REG_31__SCAN_IN), .B0(n3309), .Y(n3310));
  INVX1   g01774(.A(n3310), .Y(n3311));
  NAND2X1 g01775(.A(n3311), .B(n2684), .Y(n3312));
  OAI21X1 g01776(.A0(n2684), .A1(n2081), .B0(n3312), .Y(n3313));
  XOR2X1  g01777(.A(n3313), .B(n3299), .Y(n3314));
  NOR2X1  g01778(.A(n3308), .B(n3314), .Y(n3315));
  AOI21X1 g01779(.A0(n3314), .A1(n3308), .B0(n3315), .Y(n3317));
  INVX1   g01780(.A(n3317), .Y(n3318));
  OAI21X1 g01781(.A0(n2725), .A1(n2751), .B0(n3318), .Y(n3319));
  NAND4X1 g01782(.A(n3262), .B(n3190), .C(n3170), .D(n3264), .Y(n3320));
  AOI21X1 g01783(.A0(n3320), .A1(n3269), .B0(n3265), .Y(n3321));
  AOI22X1 g01784(.A0(n3104), .A1(n3120), .B0(n3067), .B1(n3050), .Y(n3322));
  OAI21X1 g01785(.A0(n3087), .A1(n3081), .B0(n3322), .Y(n3323));
  AOI21X1 g01786(.A0(n3104), .A1(n3128), .B0(n3120), .Y(n3324));
  AOI21X1 g01787(.A0(n3103), .A1(n3132), .B0(n3324), .Y(n3325));
  NAND2X1 g01788(.A(n3167), .B(n3153), .Y(n3326));
  NAND3X1 g01789(.A(n3264), .B(n3262), .C(n3326), .Y(n3327));
  AOI21X1 g01790(.A0(n3325), .A1(n3323), .B0(n3327), .Y(n3328));
  NOR2X1  g01791(.A(n3328), .B(n3321), .Y(n3329));
  XOR2X1  g01792(.A(n3329), .B(n3314), .Y(n3330));
  INVX1   g01793(.A(n3330), .Y(n3331));
  AOI22X1 g01794(.A0(n3318), .A1(n2724), .B0(n2715), .B1(n3331), .Y(n3332));
  AOI22X1 g01795(.A0(n3266), .A1(n2786), .B0(n2721), .B1(n3331), .Y(n3333));
  OAI21X1 g01796(.A0(n2720), .A1(n2714), .B0(n3331), .Y(n3334));
  NAND4X1 g01797(.A(n3333), .B(n3332), .C(n3319), .D(n3334), .Y(n3335));
  NOR4X1  g01798(.A(n3215), .B(n3167), .C(n3187), .D(n3259), .Y(n3336));
  NOR2X1  g01799(.A(n2684), .B(n2081), .Y(n3337));
  AOI21X1 g01800(.A0(n3311), .A1(n2684), .B0(n3337), .Y(n3338));
  XOR2X1  g01801(.A(n3338), .B(n3336), .Y(n3339));
  NAND4X1 g01802(.A(P1_REG3_REG_10__SCAN_IN), .B(P1_REG3_REG_12__SCAN_IN), .C(P1_REG3_REG_11__SCAN_IN), .D(n3192), .Y(n3340));
  XOR2X1  g01803(.A(n3340), .B(P1_REG3_REG_13__SCAN_IN), .Y(n3341));
  INVX1   g01804(.A(n3341), .Y(n3342));
  AOI22X1 g01805(.A0(n2735), .A1(n3342), .B0(n2730), .B1(P1_REG0_REG_13__SCAN_IN), .Y(n3343));
  AOI22X1 g01806(.A0(n2731), .A1(P1_REG2_REG_13__SCAN_IN), .B0(P1_REG1_REG_13__SCAN_IN), .B1(n2734), .Y(n3344));
  NAND2X1 g01807(.A(n3344), .B(n3343), .Y(n3345));
  INVX1   g01808(.A(n3345), .Y(n3346));
  OAI22X1 g01809(.A0(n3338), .A1(n2744), .B0(n2791), .B1(n3346), .Y(n3347));
  AOI21X1 g01810(.A0(n3339), .A1(n2740), .B0(n3347), .Y(n3348));
  OAI21X1 g01811(.A0(n3317), .A1(n2728), .B0(n3348), .Y(n3349));
  NOR2X1  g01812(.A(n3349), .B(n3335), .Y(n3350));
  NAND2X1 g01813(.A(n2679), .B(P1_REG0_REG_12__SCAN_IN), .Y(n3351));
  OAI21X1 g01814(.A0(n3350), .A1(n2679), .B0(n3351), .Y(P1_U3495));
  NOR2X1  g01815(.A(n3338), .B(n3299), .Y(n3353));
  NOR2X1  g01816(.A(P1_IR_REG_31__SCAN_IN), .B(n2105), .Y(n3354));
  AOI21X1 g01817(.A0(n2106), .A1(P1_IR_REG_31__SCAN_IN), .B0(n3354), .Y(n3355));
  INVX1   g01818(.A(n3355), .Y(n3356));
  NAND3X1 g01819(.A(n3356), .B(n2687), .C(n2686), .Y(n3357));
  OAI21X1 g01820(.A0(n2684), .A1(n2104), .B0(n3357), .Y(n3358));
  NOR2X1  g01821(.A(n2684), .B(n2104), .Y(n3359));
  AOI21X1 g01822(.A0(n3356), .A1(n2684), .B0(n3359), .Y(n3360));
  AOI22X1 g01823(.A0(n3346), .A1(n3360), .B0(n3338), .B1(n3299), .Y(n3361));
  INVX1   g01824(.A(n3361), .Y(n3362));
  AOI21X1 g01825(.A0(n3358), .A1(n3345), .B0(n3362), .Y(n3363));
  OAI21X1 g01826(.A0(n3353), .A1(n3308), .B0(n3363), .Y(n3364));
  INVX1   g01827(.A(n3299), .Y(n3365));
  NOR2X1  g01828(.A(n3313), .B(n3365), .Y(n3366));
  NOR2X1  g01829(.A(n3360), .B(n3345), .Y(n3367));
  NOR2X1  g01830(.A(n3358), .B(n3346), .Y(n3368));
  NOR3X1  g01831(.A(n3368), .B(n3367), .C(n3353), .Y(n3369));
  OAI21X1 g01832(.A0(n3366), .A1(n3307), .B0(n3369), .Y(n3370));
  NAND2X1 g01833(.A(n3370), .B(n3364), .Y(n3371));
  OAI22X1 g01834(.A0(n3299), .A1(n2854), .B0(n2723), .B1(n3371), .Y(n3372));
  AOI21X1 g01835(.A0(n2875), .A1(n2717), .B0(n3371), .Y(n3373));
  XOR2X1  g01836(.A(n3358), .B(n3346), .Y(n3374));
  NOR2X1  g01837(.A(n3313), .B(n3299), .Y(n3375));
  NAND2X1 g01838(.A(n3320), .B(n3269), .Y(n3376));
  NAND2X1 g01839(.A(n3376), .B(n3264), .Y(n3377));
  NOR3X1  g01840(.A(n3265), .B(n3253), .C(n3226), .Y(n3378));
  OAI21X1 g01841(.A0(n3179), .A1(n3177), .B0(n3378), .Y(n3379));
  AOI22X1 g01842(.A0(n3377), .A1(n3379), .B0(n3313), .B1(n3299), .Y(n3380));
  NOR2X1  g01843(.A(n3380), .B(n3375), .Y(n3381));
  XOR2X1  g01844(.A(n3381), .B(n3374), .Y(n3382));
  INVX1   g01845(.A(n3382), .Y(n3383));
  OAI21X1 g01846(.A0(n2721), .A1(n2720), .B0(n3383), .Y(n3384));
  OAI21X1 g01847(.A0(n2715), .A1(n2714), .B0(n3383), .Y(n3385));
  NAND2X1 g01848(.A(n3385), .B(n3384), .Y(n3386));
  INVX1   g01849(.A(n3336), .Y(n3387));
  NOR2X1  g01850(.A(n3313), .B(n3387), .Y(n3388));
  XOR2X1  g01851(.A(n3360), .B(n3388), .Y(n3389));
  INVX1   g01852(.A(P1_REG3_REG_14__SCAN_IN), .Y(n3390));
  INVX1   g01853(.A(P1_REG3_REG_13__SCAN_IN), .Y(n3391));
  NOR2X1  g01854(.A(n3340), .B(n3391), .Y(n3392));
  XOR2X1  g01855(.A(n3392), .B(n3390), .Y(n3393));
  INVX1   g01856(.A(n3393), .Y(n3394));
  INVX1   g01857(.A(P1_REG1_REG_14__SCAN_IN), .Y(n3395));
  AOI22X1 g01858(.A0(n2730), .A1(P1_REG0_REG_14__SCAN_IN), .B0(P1_REG2_REG_14__SCAN_IN), .B1(n2731), .Y(n3396));
  OAI21X1 g01859(.A0(n2707), .A1(n3395), .B0(n3396), .Y(n3397));
  AOI21X1 g01860(.A0(n3394), .A1(n2735), .B0(n3397), .Y(n3398));
  OAI22X1 g01861(.A0(n3360), .A1(n2744), .B0(n2791), .B1(n3398), .Y(n3399));
  AOI21X1 g01862(.A0(n3389), .A1(n2740), .B0(n3399), .Y(n3400));
  OAI21X1 g01863(.A0(n3371), .A1(n2728), .B0(n3400), .Y(n3401));
  NOR4X1  g01864(.A(n3386), .B(n3373), .C(n3372), .D(n3401), .Y(n3402));
  NAND2X1 g01865(.A(n2679), .B(P1_REG0_REG_13__SCAN_IN), .Y(n3403));
  OAI21X1 g01866(.A0(n3402), .A1(n2679), .B0(n3403), .Y(P1_U3498));
  INVX1   g01867(.A(n3398), .Y(n3405));
  NOR2X1  g01868(.A(P1_IR_REG_31__SCAN_IN), .B(n2121), .Y(n3406));
  AOI21X1 g01869(.A0(n2125), .A1(P1_IR_REG_31__SCAN_IN), .B0(n3406), .Y(n3407));
  INVX1   g01870(.A(n3407), .Y(n3408));
  NOR2X1  g01871(.A(n2684), .B(n2120), .Y(n3409));
  AOI21X1 g01872(.A0(n3408), .A1(n2684), .B0(n3409), .Y(n3410));
  XOR2X1  g01873(.A(n3410), .B(n3405), .Y(n3411));
  INVX1   g01874(.A(n3375), .Y(n3412));
  OAI22X1 g01875(.A0(n3321), .A1(n3328), .B0(n3338), .B1(n3365), .Y(n3413));
  AOI21X1 g01876(.A0(n3413), .A1(n3412), .B0(n3367), .Y(n3414));
  NOR2X1  g01877(.A(n3414), .B(n3368), .Y(n3415));
  XOR2X1  g01878(.A(n3415), .B(n3411), .Y(n3416));
  NOR2X1  g01879(.A(n3416), .B(n3252), .Y(n3417));
  NAND3X1 g01880(.A(n3361), .B(n3259), .C(n3266), .Y(n3418));
  AOI22X1 g01881(.A0(n3345), .A1(n3358), .B0(n3313), .B1(n3365), .Y(n3419));
  AOI22X1 g01882(.A0(n3418), .A1(n3419), .B0(n3360), .B1(n3346), .Y(n3420));
  AOI21X1 g01883(.A0(n3361), .A1(n3306), .B0(n3420), .Y(n3421));
  XOR2X1  g01884(.A(n3421), .B(n3411), .Y(n3422));
  AOI22X1 g01885(.A0(n3345), .A1(n2786), .B0(n2724), .B1(n3422), .Y(n3423));
  OAI21X1 g01886(.A0(n2725), .A1(n2751), .B0(n3422), .Y(n3424));
  NAND2X1 g01887(.A(n3424), .B(n3423), .Y(n3425));
  NOR2X1  g01888(.A(n3416), .B(n2716), .Y(n3426));
  AOI21X1 g01889(.A0(n3289), .A1(n3288), .B0(n3416), .Y(n3427));
  NOR4X1  g01890(.A(n3426), .B(n3425), .C(n3417), .D(n3427), .Y(n3428));
  INVX1   g01891(.A(n3428), .Y(n3429));
  INVX1   g01892(.A(n3422), .Y(n3430));
  NOR2X1  g01893(.A(n3430), .B(n2728), .Y(n3431));
  NOR3X1  g01894(.A(n3358), .B(n3313), .C(n3387), .Y(n3432));
  NAND4X1 g01895(.A(n3360), .B(n3338), .C(n3336), .D(n3410), .Y(n3433));
  OAI21X1 g01896(.A0(n3410), .A1(n3432), .B0(n3433), .Y(n3434));
  NOR2X1  g01897(.A(n3434), .B(n2741), .Y(n3435));
  INVX1   g01898(.A(P1_REG3_REG_15__SCAN_IN), .Y(n3436));
  NOR3X1  g01899(.A(n3340), .B(n3390), .C(n3391), .Y(n3437));
  XOR2X1  g01900(.A(n3437), .B(n3436), .Y(n3438));
  INVX1   g01901(.A(n3438), .Y(n3439));
  INVX1   g01902(.A(P1_REG1_REG_15__SCAN_IN), .Y(n3440));
  AOI22X1 g01903(.A0(n2730), .A1(P1_REG0_REG_15__SCAN_IN), .B0(P1_REG2_REG_15__SCAN_IN), .B1(n2731), .Y(n3441));
  OAI21X1 g01904(.A0(n2707), .A1(n3440), .B0(n3441), .Y(n3442));
  AOI21X1 g01905(.A0(n3439), .A1(n2735), .B0(n3442), .Y(n3443));
  OAI22X1 g01906(.A0(n3410), .A1(n2744), .B0(n2791), .B1(n3443), .Y(n3444));
  NOR4X1  g01907(.A(n3435), .B(n3431), .C(n3429), .D(n3444), .Y(n3445));
  NAND2X1 g01908(.A(n2679), .B(P1_REG0_REG_14__SCAN_IN), .Y(n3446));
  OAI21X1 g01909(.A0(n3445), .A1(n2679), .B0(n3446), .Y(P1_U3501));
  NOR2X1  g01910(.A(P1_IR_REG_31__SCAN_IN), .B(n2144), .Y(n3448));
  AOI21X1 g01911(.A0(n2145), .A1(P1_IR_REG_31__SCAN_IN), .B0(n3448), .Y(n3449));
  INVX1   g01912(.A(n3449), .Y(n3450));
  NAND2X1 g01913(.A(n3450), .B(n2684), .Y(n3451));
  OAI21X1 g01914(.A0(n2684), .A1(n2143), .B0(n3451), .Y(n3452));
  XOR2X1  g01915(.A(n3452), .B(n3443), .Y(n3453));
  INVX1   g01916(.A(n3453), .Y(n3454));
  NOR2X1  g01917(.A(n3410), .B(n3405), .Y(n3455));
  NAND2X1 g01918(.A(n3410), .B(n3405), .Y(n3456));
  OAI21X1 g01919(.A0(n3415), .A1(n3455), .B0(n3456), .Y(n3457));
  XOR2X1  g01920(.A(n3457), .B(n3454), .Y(n3458));
  NOR2X1  g01921(.A(n3458), .B(n3252), .Y(n3459));
  INVX1   g01922(.A(n3410), .Y(n3460));
  NAND2X1 g01923(.A(n3460), .B(n3405), .Y(n3461));
  NOR2X1  g01924(.A(n3460), .B(n3405), .Y(n3462));
  OAI21X1 g01925(.A0(n3462), .A1(n3421), .B0(n3461), .Y(n3463));
  XOR2X1  g01926(.A(n3463), .B(n3453), .Y(n3464));
  INVX1   g01927(.A(n3464), .Y(n3465));
  AOI22X1 g01928(.A0(n3405), .A1(n2786), .B0(n2724), .B1(n3465), .Y(n3466));
  OAI21X1 g01929(.A0(n2725), .A1(n2751), .B0(n3465), .Y(n3467));
  NAND2X1 g01930(.A(n3467), .B(n3466), .Y(n3468));
  NOR2X1  g01931(.A(n3458), .B(n2716), .Y(n3469));
  AOI21X1 g01932(.A0(n3289), .A1(n3288), .B0(n3458), .Y(n3470));
  NOR4X1  g01933(.A(n3469), .B(n3468), .C(n3459), .D(n3470), .Y(n3471));
  INVX1   g01934(.A(n3471), .Y(n3472));
  XOR2X1  g01935(.A(n3452), .B(n3433), .Y(n3473));
  INVX1   g01936(.A(n3452), .Y(n3474));
  INVX1   g01937(.A(P1_REG3_REG_16__SCAN_IN), .Y(n3475));
  NOR4X1  g01938(.A(n3390), .B(n3391), .C(n3436), .D(n3340), .Y(n3476));
  XOR2X1  g01939(.A(n3476), .B(n3475), .Y(n3477));
  INVX1   g01940(.A(n3477), .Y(n3478));
  INVX1   g01941(.A(P1_REG1_REG_16__SCAN_IN), .Y(n3479));
  AOI22X1 g01942(.A0(n2730), .A1(P1_REG0_REG_16__SCAN_IN), .B0(P1_REG2_REG_16__SCAN_IN), .B1(n2731), .Y(n3480));
  OAI21X1 g01943(.A0(n2707), .A1(n3479), .B0(n3480), .Y(n3481));
  AOI21X1 g01944(.A0(n3478), .A1(n2735), .B0(n3481), .Y(n3482));
  OAI22X1 g01945(.A0(n3474), .A1(n2744), .B0(n2791), .B1(n3482), .Y(n3483));
  AOI21X1 g01946(.A0(n3473), .A1(n2740), .B0(n3483), .Y(n3484));
  OAI21X1 g01947(.A0(n3464), .A1(n2728), .B0(n3484), .Y(n3485));
  NOR2X1  g01948(.A(n3485), .B(n3472), .Y(n3486));
  NAND2X1 g01949(.A(n2679), .B(P1_REG0_REG_15__SCAN_IN), .Y(n3487));
  OAI21X1 g01950(.A0(n3486), .A1(n2679), .B0(n3487), .Y(P1_U3504));
  INVX1   g01951(.A(n3443), .Y(n3489));
  NOR2X1  g01952(.A(n3474), .B(n3489), .Y(n3490));
  AOI21X1 g01953(.A0(n3474), .A1(n3489), .B0(n3457), .Y(n3491));
  NOR2X1  g01954(.A(P1_IR_REG_31__SCAN_IN), .B(n2166), .Y(n3492));
  AOI21X1 g01955(.A0(n2178), .A1(P1_IR_REG_31__SCAN_IN), .B0(n3492), .Y(n3493));
  INVX1   g01956(.A(n3493), .Y(n3494));
  NAND2X1 g01957(.A(n3494), .B(n2684), .Y(n3495));
  OAI21X1 g01958(.A0(n2684), .A1(n2165), .B0(n3495), .Y(n3496));
  XOR2X1  g01959(.A(n3496), .B(n3482), .Y(n3497));
  NOR3X1  g01960(.A(n3497), .B(n3491), .C(n3490), .Y(n3498));
  NAND2X1 g01961(.A(n3452), .B(n3443), .Y(n3499));
  NAND2X1 g01962(.A(n3457), .B(n3499), .Y(n3500));
  NAND2X1 g01963(.A(n3496), .B(n3482), .Y(n3501));
  INVX1   g01964(.A(n3501), .Y(n3502));
  INVX1   g01965(.A(n3482), .Y(n3503));
  INVX1   g01966(.A(n3496), .Y(n3504));
  AOI22X1 g01967(.A0(n3503), .A1(n3504), .B0(n3474), .B1(n3489), .Y(n3505));
  INVX1   g01968(.A(n3505), .Y(n3506));
  NOR2X1  g01969(.A(n3506), .B(n3502), .Y(n3507));
  AOI21X1 g01970(.A0(n3507), .A1(n3500), .B0(n3498), .Y(n3508));
  NOR2X1  g01971(.A(n3508), .B(n3252), .Y(n3509));
  INVX1   g01972(.A(n3509), .Y(n3510));
  NOR2X1  g01973(.A(n3474), .B(n3443), .Y(n3511));
  NAND2X1 g01974(.A(n3474), .B(n3443), .Y(n3512));
  AOI21X1 g01975(.A0(n3512), .A1(n3463), .B0(n3511), .Y(n3513));
  INVX1   g01976(.A(n3513), .Y(n3514));
  NOR2X1  g01977(.A(n3514), .B(n3497), .Y(n3515));
  AOI21X1 g01978(.A0(n3497), .A1(n3514), .B0(n3515), .Y(n3517));
  INVX1   g01979(.A(n3517), .Y(n3518));
  AOI22X1 g01980(.A0(n3489), .A1(n2786), .B0(n2724), .B1(n3518), .Y(n3519));
  OAI21X1 g01981(.A0(n2725), .A1(n2751), .B0(n3518), .Y(n3520));
  NAND3X1 g01982(.A(n3520), .B(n3519), .C(n3510), .Y(n3521));
  NOR2X1  g01983(.A(n3508), .B(n2716), .Y(n3522));
  AOI21X1 g01984(.A0(n3289), .A1(n3288), .B0(n3508), .Y(n3523));
  NOR2X1  g01985(.A(n3452), .B(n3433), .Y(n3524));
  XOR2X1  g01986(.A(n3504), .B(n3524), .Y(n3525));
  NAND2X1 g01987(.A(n3476), .B(P1_REG3_REG_16__SCAN_IN), .Y(n3526));
  XOR2X1  g01988(.A(n3526), .B(P1_REG3_REG_17__SCAN_IN), .Y(n3527));
  INVX1   g01989(.A(n3527), .Y(n3528));
  INVX1   g01990(.A(P1_REG1_REG_17__SCAN_IN), .Y(n3529));
  AOI22X1 g01991(.A0(n2730), .A1(P1_REG0_REG_17__SCAN_IN), .B0(P1_REG2_REG_17__SCAN_IN), .B1(n2731), .Y(n3530));
  OAI21X1 g01992(.A0(n2707), .A1(n3529), .B0(n3530), .Y(n3531));
  AOI21X1 g01993(.A0(n3528), .A1(n2735), .B0(n3531), .Y(n3532));
  OAI22X1 g01994(.A0(n3504), .A1(n2744), .B0(n2791), .B1(n3532), .Y(n3533));
  AOI21X1 g01995(.A0(n3525), .A1(n2740), .B0(n3533), .Y(n3534));
  OAI21X1 g01996(.A0(n3517), .A1(n2728), .B0(n3534), .Y(n3535));
  NOR4X1  g01997(.A(n3523), .B(n3522), .C(n3521), .D(n3535), .Y(n3536));
  NAND2X1 g01998(.A(n2679), .B(P1_REG0_REG_16__SCAN_IN), .Y(n3537));
  OAI21X1 g01999(.A0(n3536), .A1(n2679), .B0(n3537), .Y(P1_U3507));
  NAND2X1 g02000(.A(n3496), .B(n3503), .Y(n3539));
  INVX1   g02001(.A(n3539), .Y(n3540));
  INVX1   g02002(.A(n3532), .Y(n3541));
  NOR2X1  g02003(.A(P1_IR_REG_31__SCAN_IN), .B(n2195), .Y(n3542));
  AOI21X1 g02004(.A0(n2196), .A1(P1_IR_REG_31__SCAN_IN), .B0(n3542), .Y(n3543));
  INVX1   g02005(.A(n3543), .Y(n3544));
  NOR2X1  g02006(.A(n2684), .B(n2194), .Y(n3545));
  AOI21X1 g02007(.A0(n3544), .A1(n2684), .B0(n3545), .Y(n3546));
  INVX1   g02008(.A(n3546), .Y(n3547));
  OAI22X1 g02009(.A0(n3541), .A1(n3547), .B0(n3496), .B1(n3503), .Y(n3548));
  AOI21X1 g02010(.A0(n3547), .A1(n3541), .B0(n3548), .Y(n3549));
  OAI21X1 g02011(.A0(n3540), .A1(n3514), .B0(n3549), .Y(n3550));
  NOR2X1  g02012(.A(n3496), .B(n3503), .Y(n3551));
  NOR2X1  g02013(.A(n5484), .B(n3540), .Y(n3554));
  OAI21X1 g02014(.A0(n3551), .A1(n3513), .B0(n3554), .Y(n3555));
  NAND2X1 g02015(.A(n3555), .B(n3550), .Y(n3556));
  AOI21X1 g02016(.A0(n2875), .A1(n2717), .B0(n3556), .Y(n3557));
  NAND3X1 g02017(.A(n3499), .B(n3410), .C(n3405), .Y(n3558));
  AOI21X1 g02018(.A0(n3558), .A1(n3505), .B0(n3502), .Y(n3559));
  INVX1   g02019(.A(n3559), .Y(n3560));
  NOR3X1  g02020(.A(n3502), .B(n3490), .C(n3455), .Y(n3561));
  OAI21X1 g02021(.A0(n3414), .A1(n3368), .B0(n3561), .Y(n3562));
  NAND2X1 g02022(.A(n3562), .B(n3560), .Y(n3563));
  XOR2X1  g02023(.A(n3563), .B(n5484), .Y(n3564));
  OAI22X1 g02024(.A0(n3556), .A1(n2723), .B0(n2716), .B1(n3564), .Y(n3565));
  INVX1   g02025(.A(n3564), .Y(n3566));
  AOI22X1 g02026(.A0(n3503), .A1(n2786), .B0(n2721), .B1(n3566), .Y(n3567));
  OAI21X1 g02027(.A0(n2720), .A1(n2714), .B0(n3566), .Y(n3568));
  NAND2X1 g02028(.A(n3568), .B(n3567), .Y(n3569));
  NOR3X1  g02029(.A(n3496), .B(n3452), .C(n3433), .Y(n3570));
  XOR2X1  g02030(.A(n3546), .B(n3570), .Y(n3571));
  NAND3X1 g02031(.A(n3476), .B(P1_REG3_REG_16__SCAN_IN), .C(P1_REG3_REG_17__SCAN_IN), .Y(n3572));
  XOR2X1  g02032(.A(n3572), .B(P1_REG3_REG_18__SCAN_IN), .Y(n3573));
  INVX1   g02033(.A(n3573), .Y(n3574));
  INVX1   g02034(.A(P1_REG1_REG_18__SCAN_IN), .Y(n3575));
  AOI22X1 g02035(.A0(n2730), .A1(P1_REG0_REG_18__SCAN_IN), .B0(P1_REG2_REG_18__SCAN_IN), .B1(n2731), .Y(n3576));
  OAI21X1 g02036(.A0(n2707), .A1(n3575), .B0(n3576), .Y(n3577));
  AOI21X1 g02037(.A0(n3574), .A1(n2735), .B0(n3577), .Y(n3578));
  OAI22X1 g02038(.A0(n3546), .A1(n2744), .B0(n2791), .B1(n3578), .Y(n3579));
  AOI21X1 g02039(.A0(n3571), .A1(n2740), .B0(n3579), .Y(n3580));
  OAI21X1 g02040(.A0(n3556), .A1(n2728), .B0(n3580), .Y(n3581));
  NOR4X1  g02041(.A(n3569), .B(n3565), .C(n3557), .D(n3581), .Y(n3582));
  NAND2X1 g02042(.A(n2679), .B(P1_REG0_REG_17__SCAN_IN), .Y(n3583));
  OAI21X1 g02043(.A0(n3582), .A1(n2679), .B0(n3583), .Y(P1_U3510));
  AOI21X1 g02044(.A0(n3546), .A1(n3539), .B0(n3532), .Y(n3585));
  AOI21X1 g02045(.A0(n3547), .A1(n3540), .B0(n3585), .Y(n3586));
  OAI21X1 g02046(.A0(n3548), .A1(n3513), .B0(n3586), .Y(n3587));
  INVX1   g02047(.A(n3578), .Y(n3588));
  NOR2X1  g02048(.A(P1_IR_REG_31__SCAN_IN), .B(n2334), .Y(n3589));
  AOI21X1 g02049(.A0(n2224), .A1(P1_IR_REG_31__SCAN_IN), .B0(n3589), .Y(n3590));
  INVX1   g02050(.A(n3590), .Y(n3591));
  NOR2X1  g02051(.A(n2684), .B(n2212), .Y(n3592));
  AOI21X1 g02052(.A0(n3591), .A1(n2684), .B0(n3592), .Y(n3593));
  XOR2X1  g02053(.A(n3593), .B(n3588), .Y(n3594));
  NOR2X1  g02054(.A(n3594), .B(n3587), .Y(n3595));
  XOR2X1  g02055(.A(n3593), .B(n3578), .Y(n3596));
  AOI21X1 g02056(.A0(n3594), .A1(n3587), .B0(n3595), .Y(n3598));
  INVX1   g02057(.A(n3598), .Y(n3599));
  AOI22X1 g02058(.A0(n3541), .A1(n2786), .B0(n2724), .B1(n3599), .Y(n3600));
  OAI21X1 g02059(.A0(n2725), .A1(n2751), .B0(n3599), .Y(n3601));
  NOR2X1  g02060(.A(n3547), .B(n3532), .Y(n3602));
  AOI22X1 g02061(.A0(n3560), .A1(n3562), .B0(n3547), .B1(n3532), .Y(n3603));
  NOR2X1  g02062(.A(n3603), .B(n3602), .Y(n3604));
  XOR2X1  g02063(.A(n3604), .B(n3594), .Y(n3605));
  INVX1   g02064(.A(n3605), .Y(n3606));
  OAI21X1 g02065(.A0(n2721), .A1(n2720), .B0(n3606), .Y(n3607));
  OAI21X1 g02066(.A0(n2715), .A1(n2714), .B0(n3606), .Y(n3608));
  NAND4X1 g02067(.A(n3607), .B(n3601), .C(n3600), .D(n3608), .Y(n3609));
  NOR2X1  g02068(.A(n3598), .B(n2728), .Y(n3610));
  NOR4X1  g02069(.A(n3496), .B(n3452), .C(n3433), .D(n3547), .Y(n3611));
  NAND3X1 g02070(.A(n3593), .B(n3546), .C(n3570), .Y(n3612));
  OAI21X1 g02071(.A0(n3593), .A1(n3611), .B0(n3612), .Y(n3613));
  NOR2X1  g02072(.A(n3613), .B(n2741), .Y(n3614));
  NAND4X1 g02073(.A(P1_REG3_REG_16__SCAN_IN), .B(P1_REG3_REG_17__SCAN_IN), .C(P1_REG3_REG_18__SCAN_IN), .D(n3476), .Y(n3615));
  XOR2X1  g02074(.A(n3615), .B(P1_REG3_REG_19__SCAN_IN), .Y(n3616));
  INVX1   g02075(.A(n3616), .Y(n3617));
  NAND3X1 g02076(.A(n2765), .B(n2703), .C(P1_REG1_REG_19__SCAN_IN), .Y(n3618));
  AOI22X1 g02077(.A0(n2730), .A1(P1_REG0_REG_19__SCAN_IN), .B0(P1_REG2_REG_19__SCAN_IN), .B1(n2731), .Y(n3619));
  NAND2X1 g02078(.A(n3619), .B(n3618), .Y(n3620));
  AOI21X1 g02079(.A0(n3617), .A1(n2735), .B0(n3620), .Y(n3621));
  OAI22X1 g02080(.A0(n3593), .A1(n2744), .B0(n2791), .B1(n3621), .Y(n3622));
  NOR4X1  g02081(.A(n3614), .B(n3610), .C(n3609), .D(n3622), .Y(n3623));
  NAND2X1 g02082(.A(n2679), .B(P1_REG0_REG_18__SCAN_IN), .Y(n3624));
  OAI21X1 g02083(.A0(n3623), .A1(n2679), .B0(n3624), .Y(P1_U3513));
  NAND3X1 g02084(.A(n2687), .B(n2686), .C(n2673), .Y(n3626));
  OAI21X1 g02085(.A0(n2684), .A1(n2240), .B0(n3626), .Y(n3627));
  XOR2X1  g02086(.A(n3627), .B(n3621), .Y(n3628));
  INVX1   g02087(.A(n3602), .Y(n3629));
  INVX1   g02088(.A(n3368), .Y(n3630));
  OAI22X1 g02089(.A0(n3360), .A1(n3345), .B0(n3375), .B1(n3380), .Y(n3631));
  INVX1   g02090(.A(n3561), .Y(n3632));
  AOI21X1 g02091(.A0(n3631), .A1(n3630), .B0(n3632), .Y(n3633));
  OAI22X1 g02092(.A0(n3559), .A1(n3633), .B0(n3546), .B1(n3541), .Y(n3634));
  AOI21X1 g02093(.A0(n3634), .A1(n3629), .B0(n3578), .Y(n3635));
  NAND3X1 g02094(.A(n3634), .B(n3578), .C(n3629), .Y(n3636));
  AOI21X1 g02095(.A0(n3636), .A1(n3593), .B0(n3635), .Y(n3637));
  XOR2X1  g02096(.A(n3637), .B(n3628), .Y(n3638));
  NOR2X1  g02097(.A(n3638), .B(n3252), .Y(n3639));
  INVX1   g02098(.A(n3593), .Y(n3640));
  NOR2X1  g02099(.A(n3640), .B(n3588), .Y(n3641));
  INVX1   g02100(.A(n3641), .Y(n3642));
  NOR2X1  g02101(.A(n3593), .B(n3578), .Y(n3643));
  AOI21X1 g02102(.A0(n3642), .A1(n3587), .B0(n3643), .Y(n3644));
  INVX1   g02103(.A(n3644), .Y(n3645));
  NOR2X1  g02104(.A(n3645), .B(n3628), .Y(n3646));
  AOI21X1 g02105(.A0(n3628), .A1(n3645), .B0(n3646), .Y(n3648));
  OAI22X1 g02106(.A0(n3578), .A1(n2854), .B0(n2723), .B1(n3648), .Y(n3649));
  AOI21X1 g02107(.A0(n2875), .A1(n2717), .B0(n3648), .Y(n3650));
  NOR3X1  g02108(.A(n3650), .B(n3649), .C(n3639), .Y(n3651));
  NOR2X1  g02109(.A(n3638), .B(n2716), .Y(n3652));
  AOI21X1 g02110(.A0(n3289), .A1(n3288), .B0(n3638), .Y(n3653));
  NOR2X1  g02111(.A(n3653), .B(n3652), .Y(n3654));
  NAND2X1 g02112(.A(n3654), .B(n3651), .Y(n3655));
  XOR2X1  g02113(.A(n3627), .B(n3612), .Y(n3656));
  INVX1   g02114(.A(n3627), .Y(n3657));
  INVX1   g02115(.A(P1_REG3_REG_20__SCAN_IN), .Y(n3658));
  INVX1   g02116(.A(P1_REG3_REG_19__SCAN_IN), .Y(n3659));
  NOR2X1  g02117(.A(n3615), .B(n3659), .Y(n3660));
  XOR2X1  g02118(.A(n3660), .B(n3658), .Y(n3661));
  AOI22X1 g02119(.A0(n2730), .A1(P1_REG0_REG_20__SCAN_IN), .B0(P1_REG2_REG_20__SCAN_IN), .B1(n2731), .Y(n3662));
  INVX1   g02120(.A(n3662), .Y(n3663));
  AOI21X1 g02121(.A0(n2734), .A1(P1_REG1_REG_20__SCAN_IN), .B0(n3663), .Y(n3664));
  OAI21X1 g02122(.A0(n3661), .A1(n2708), .B0(n3664), .Y(n3665));
  INVX1   g02123(.A(n3665), .Y(n3666));
  OAI22X1 g02124(.A0(n3657), .A1(n2744), .B0(n2791), .B1(n3666), .Y(n3667));
  AOI21X1 g02125(.A0(n3656), .A1(n2740), .B0(n3667), .Y(n3668));
  OAI21X1 g02126(.A0(n3648), .A1(n2728), .B0(n3668), .Y(n3669));
  NOR2X1  g02127(.A(n3669), .B(n3655), .Y(n3670));
  NAND2X1 g02128(.A(n2679), .B(P1_REG0_REG_19__SCAN_IN), .Y(n3671));
  OAI21X1 g02129(.A0(n3670), .A1(n2679), .B0(n3671), .Y(P1_U3515));
  OAI21X1 g02130(.A0(n2262), .A1(n2251), .B0(n2810), .Y(n3673));
  XOR2X1  g02131(.A(n3673), .B(n3665), .Y(n3674));
  NAND2X1 g02132(.A(n3627), .B(n3621), .Y(n3675));
  NOR2X1  g02133(.A(n3627), .B(n3621), .Y(n3676));
  OAI21X1 g02134(.A0(n3603), .A1(n3602), .B0(n3588), .Y(n3677));
  NOR3X1  g02135(.A(n3603), .B(n3588), .C(n3602), .Y(n3678));
  OAI21X1 g02136(.A0(n3678), .A1(n3640), .B0(n3677), .Y(n3679));
  AOI21X1 g02137(.A0(n3679), .A1(n3675), .B0(n3676), .Y(n3680));
  XOR2X1  g02138(.A(n3680), .B(n3674), .Y(n3681));
  NOR2X1  g02139(.A(n3681), .B(n3252), .Y(n3682));
  INVX1   g02140(.A(n3682), .Y(n3683));
  INVX1   g02141(.A(n3621), .Y(n3684));
  AOI21X1 g02142(.A0(n3627), .A1(n3684), .B0(n3645), .Y(n3685));
  AOI22X1 g02143(.A0(n3666), .A1(n3673), .B0(n3657), .B1(n3621), .Y(n3686));
  OAI21X1 g02144(.A0(n3673), .A1(n3666), .B0(n3686), .Y(n3687));
  AOI21X1 g02145(.A0(n3657), .A1(n3621), .B0(n3644), .Y(n3688));
  NAND2X1 g02146(.A(n3627), .B(n3684), .Y(n3689));
  NAND2X1 g02147(.A(n3674), .B(n3689), .Y(n3690));
  OAI22X1 g02148(.A0(n3688), .A1(n3690), .B0(n3687), .B1(n3685), .Y(n3691));
  INVX1   g02149(.A(n3691), .Y(n3692));
  AOI22X1 g02150(.A0(n3684), .A1(n2786), .B0(n2724), .B1(n3692), .Y(n3693));
  OAI21X1 g02151(.A0(n2725), .A1(n2751), .B0(n3692), .Y(n3694));
  NOR2X1  g02152(.A(n3681), .B(n2716), .Y(n3695));
  AOI21X1 g02153(.A0(n3289), .A1(n3288), .B0(n3681), .Y(n3696));
  NOR2X1  g02154(.A(n3696), .B(n3695), .Y(n3697));
  NAND4X1 g02155(.A(n3694), .B(n3693), .C(n3683), .D(n3697), .Y(n3698));
  NOR2X1  g02156(.A(n3691), .B(n2728), .Y(n3699));
  NAND4X1 g02157(.A(n3593), .B(n3546), .C(n3570), .D(n3657), .Y(n3700));
  XOR2X1  g02158(.A(n3673), .B(n3700), .Y(n3701));
  NOR2X1  g02159(.A(n3701), .B(n2741), .Y(n3702));
  INVX1   g02160(.A(P1_REG3_REG_21__SCAN_IN), .Y(n3703));
  NOR3X1  g02161(.A(n3615), .B(n3659), .C(n3658), .Y(n3704));
  XOR2X1  g02162(.A(n3704), .B(n3703), .Y(n3705));
  AOI22X1 g02163(.A0(n2730), .A1(P1_REG0_REG_21__SCAN_IN), .B0(P1_REG2_REG_21__SCAN_IN), .B1(n2731), .Y(n3706));
  INVX1   g02164(.A(n3706), .Y(n3707));
  AOI21X1 g02165(.A0(n2734), .A1(P1_REG1_REG_21__SCAN_IN), .B0(n3707), .Y(n3708));
  OAI21X1 g02166(.A0(n3705), .A1(n2708), .B0(n3708), .Y(n3709));
  INVX1   g02167(.A(n3709), .Y(n3710));
  OAI22X1 g02168(.A0(n3673), .A1(n2744), .B0(n2791), .B1(n3710), .Y(n3711));
  NOR4X1  g02169(.A(n3702), .B(n3699), .C(n3698), .D(n3711), .Y(n3712));
  NAND2X1 g02170(.A(n2679), .B(P1_REG0_REG_20__SCAN_IN), .Y(n3713));
  OAI21X1 g02171(.A0(n3712), .A1(n2679), .B0(n3713), .Y(P1_U3516));
  NOR2X1  g02172(.A(n2684), .B(n2284), .Y(n3715));
  XOR2X1  g02173(.A(n3715), .B(n3710), .Y(n3716));
  NOR2X1  g02174(.A(n3673), .B(n3665), .Y(n3717));
  INVX1   g02175(.A(n3717), .Y(n3718));
  INVX1   g02176(.A(n3673), .Y(n3719));
  NOR2X1  g02177(.A(n3719), .B(n3666), .Y(n3720));
  INVX1   g02178(.A(n3675), .Y(n3721));
  INVX1   g02179(.A(n3676), .Y(n3722));
  OAI21X1 g02180(.A0(n3637), .A1(n3721), .B0(n3722), .Y(n3723));
  AOI21X1 g02181(.A0(n3723), .A1(n3718), .B0(n3720), .Y(n3724));
  XOR2X1  g02182(.A(n3724), .B(n3716), .Y(n3725));
  NOR2X1  g02183(.A(n3725), .B(n3252), .Y(n3726));
  INVX1   g02184(.A(n3716), .Y(n3727));
  INVX1   g02185(.A(n3686), .Y(n3728));
  NAND2X1 g02186(.A(n3673), .B(n3689), .Y(n3729));
  OAI21X1 g02187(.A0(n3673), .A1(n3689), .B0(n3666), .Y(n3730));
  NAND2X1 g02188(.A(n3730), .B(n3729), .Y(n3731));
  OAI21X1 g02189(.A0(n3728), .A1(n3644), .B0(n3731), .Y(n3732));
  NAND2X1 g02190(.A(n3732), .B(n3727), .Y(n3733));
  AOI21X1 g02191(.A0(n3730), .A1(n3729), .B0(n3727), .Y(n3734));
  OAI21X1 g02192(.A0(n3728), .A1(n3644), .B0(n3734), .Y(n3735));
  NAND2X1 g02193(.A(n3735), .B(n3733), .Y(n3736));
  OAI22X1 g02194(.A0(n3666), .A1(n2854), .B0(n2723), .B1(n3736), .Y(n3737));
  AOI21X1 g02195(.A0(n2875), .A1(n2717), .B0(n3736), .Y(n3738));
  NOR3X1  g02196(.A(n3738), .B(n3737), .C(n3726), .Y(n3739));
  INVX1   g02197(.A(n3725), .Y(n3740));
  AOI21X1 g02198(.A0(n3289), .A1(n3288), .B0(n3725), .Y(n3741));
  AOI21X1 g02199(.A0(n3740), .A1(n2715), .B0(n3741), .Y(n3742));
  NAND2X1 g02200(.A(n3742), .B(n3739), .Y(n3743));
  NOR2X1  g02201(.A(n3719), .B(n3700), .Y(n3744));
  INVX1   g02202(.A(n3715), .Y(n3745));
  XOR2X1  g02203(.A(n3745), .B(n3744), .Y(n3746));
  NOR4X1  g02204(.A(n3659), .B(n3703), .C(n3658), .D(n3615), .Y(n3747));
  XOR2X1  g02205(.A(n3747), .B(P1_REG3_REG_22__SCAN_IN), .Y(n3748));
  INVX1   g02206(.A(n3748), .Y(n3749));
  AOI22X1 g02207(.A0(n2730), .A1(P1_REG0_REG_22__SCAN_IN), .B0(P1_REG2_REG_22__SCAN_IN), .B1(n2731), .Y(n3750));
  INVX1   g02208(.A(n3750), .Y(n3751));
  AOI21X1 g02209(.A0(n2734), .A1(P1_REG1_REG_22__SCAN_IN), .B0(n3751), .Y(n3752));
  OAI21X1 g02210(.A0(n3749), .A1(n2708), .B0(n3752), .Y(n3753));
  INVX1   g02211(.A(n3753), .Y(n3754));
  OAI22X1 g02212(.A0(n3745), .A1(n2744), .B0(n2791), .B1(n3754), .Y(n3755));
  AOI21X1 g02213(.A0(n3746), .A1(n2740), .B0(n3755), .Y(n3756));
  OAI21X1 g02214(.A0(n3736), .A1(n2728), .B0(n3756), .Y(n3757));
  NOR2X1  g02215(.A(n3757), .B(n3743), .Y(n3758));
  NAND2X1 g02216(.A(n2679), .B(P1_REG0_REG_21__SCAN_IN), .Y(n3759));
  OAI21X1 g02217(.A0(n3758), .A1(n2679), .B0(n3759), .Y(P1_U3517));
  NOR2X1  g02218(.A(n2684), .B(n2306), .Y(n3761));
  NOR3X1  g02219(.A(n3709), .B(n2684), .C(n2284), .Y(n3764));
  OAI21X1 g02220(.A0(n2684), .A1(n2284), .B0(n3709), .Y(n3765));
  OAI21X1 g02221(.A0(n3724), .A1(n3764), .B0(n3765), .Y(n3766));
  XOR2X1  g02222(.A(n3766), .B(n5481), .Y(n3767));
  INVX1   g02223(.A(n3767), .Y(n3768));
  NAND2X1 g02224(.A(n3768), .B(n2721), .Y(n3769));
  NOR2X1  g02225(.A(n3715), .B(n3709), .Y(n3770));
  NOR3X1  g02226(.A(n3770), .B(n3728), .C(n3641), .Y(n3771));
  AOI22X1 g02227(.A0(n3729), .A1(n3730), .B0(n3686), .B1(n3643), .Y(n3772));
  NAND2X1 g02228(.A(n3715), .B(n3709), .Y(n3773));
  OAI21X1 g02229(.A0(n3772), .A1(n3770), .B0(n3773), .Y(n3774));
  AOI21X1 g02230(.A0(n3771), .A1(n3587), .B0(n3774), .Y(n3775));
  XOR2X1  g02231(.A(n3775), .B(n5481), .Y(n3776));
  INVX1   g02232(.A(n3776), .Y(n3777));
  AOI22X1 g02233(.A0(n3709), .A1(n2786), .B0(n2724), .B1(n3777), .Y(n3778));
  OAI21X1 g02234(.A0(n2725), .A1(n2751), .B0(n3777), .Y(n3779));
  NAND3X1 g02235(.A(n3779), .B(n3778), .C(n3769), .Y(n3780));
  NOR2X1  g02236(.A(n3767), .B(n2716), .Y(n3781));
  AOI21X1 g02237(.A0(n3289), .A1(n3288), .B0(n3767), .Y(n3782));
  NAND2X1 g02238(.A(n3745), .B(n3744), .Y(n3783));
  XOR2X1  g02239(.A(n3761), .B(n3783), .Y(n3784));
  NAND2X1 g02240(.A(n2325), .B(n2323), .Y(n3785));
  XOR2X1  g02241(.A(n2304), .B(n3785), .Y(n3786));
  NOR2X1  g02242(.A(n3786), .B(n1837), .Y(n3787));
  OAI21X1 g02243(.A0(n3787), .A1(n2290), .B0(n2810), .Y(n3788));
  NAND2X1 g02244(.A(n3747), .B(P1_REG3_REG_22__SCAN_IN), .Y(n3789));
  XOR2X1  g02245(.A(n3789), .B(P1_REG3_REG_23__SCAN_IN), .Y(n3790));
  AOI22X1 g02246(.A0(n2730), .A1(P1_REG0_REG_23__SCAN_IN), .B0(P1_REG2_REG_23__SCAN_IN), .B1(n2731), .Y(n3791));
  INVX1   g02247(.A(n3791), .Y(n3792));
  AOI21X1 g02248(.A0(n2734), .A1(P1_REG1_REG_23__SCAN_IN), .B0(n3792), .Y(n3793));
  OAI21X1 g02249(.A0(n3790), .A1(n2708), .B0(n3793), .Y(n3794));
  INVX1   g02250(.A(n3794), .Y(n3795));
  OAI22X1 g02251(.A0(n3788), .A1(n2744), .B0(n2791), .B1(n3795), .Y(n3796));
  AOI21X1 g02252(.A0(n3784), .A1(n2740), .B0(n3796), .Y(n3797));
  OAI21X1 g02253(.A0(n3776), .A1(n2728), .B0(n3797), .Y(n3798));
  NOR4X1  g02254(.A(n3782), .B(n3781), .C(n3780), .D(n3798), .Y(n3799));
  NAND2X1 g02255(.A(n2679), .B(P1_REG0_REG_22__SCAN_IN), .Y(n3800));
  OAI21X1 g02256(.A0(n3799), .A1(n2679), .B0(n3800), .Y(P1_U3518));
  NOR2X1  g02257(.A(n3761), .B(n3754), .Y(n3802));
  NOR3X1  g02258(.A(n3753), .B(n2684), .C(n2306), .Y(n3803));
  NOR2X1  g02259(.A(n2684), .B(n2332), .Y(n3804));
  XOR2X1  g02260(.A(n3804), .B(n3795), .Y(n3805));
  NOR2X1  g02261(.A(n3805), .B(n3803), .Y(n3806));
  OAI21X1 g02262(.A0(n3766), .A1(n3802), .B0(n3806), .Y(n3807));
  NOR3X1  g02263(.A(n3794), .B(n2684), .C(n2332), .Y(n3808));
  INVX1   g02264(.A(n3808), .Y(n3809));
  INVX1   g02265(.A(n3803), .Y(n3810));
  NAND2X1 g02266(.A(n3766), .B(n3810), .Y(n3811));
  NAND2X1 g02267(.A(n2351), .B(n2349), .Y(n3812));
  XOR2X1  g02268(.A(n2330), .B(n3812), .Y(n3813));
  NOR2X1  g02269(.A(n3813), .B(n1837), .Y(n3814));
  OAI21X1 g02270(.A0(n3814), .A1(n2320), .B0(n2810), .Y(n3815));
  AOI21X1 g02271(.A0(n3815), .A1(n3794), .B0(n3802), .Y(n3816));
  NAND3X1 g02272(.A(n3816), .B(n3811), .C(n3809), .Y(n3817));
  AOI21X1 g02273(.A0(n3817), .A1(n3807), .B0(n3252), .Y(n3818));
  NAND2X1 g02274(.A(n3761), .B(n3753), .Y(n3819));
  NOR2X1  g02275(.A(n3761), .B(n3753), .Y(n3820));
  OAI21X1 g02276(.A0(n3820), .A1(n3775), .B0(n3819), .Y(n3821));
  XOR2X1  g02277(.A(n3821), .B(n3805), .Y(n3822));
  OAI22X1 g02278(.A0(n3754), .A1(n2854), .B0(n2723), .B1(n3822), .Y(n3823));
  AOI21X1 g02279(.A0(n2875), .A1(n2717), .B0(n3822), .Y(n3824));
  NOR3X1  g02280(.A(n3824), .B(n3823), .C(n3818), .Y(n3825));
  AOI21X1 g02281(.A0(n3817), .A1(n3807), .B0(n2716), .Y(n3826));
  AOI22X1 g02282(.A0(n3807), .A1(n3817), .B0(n3289), .B1(n3288), .Y(n3827));
  NOR2X1  g02283(.A(n3827), .B(n3826), .Y(n3828));
  NAND2X1 g02284(.A(n3828), .B(n3825), .Y(n3829));
  NOR4X1  g02285(.A(n3715), .B(n3719), .C(n3700), .D(n3761), .Y(n3830));
  XOR2X1  g02286(.A(n3815), .B(n3830), .Y(n3831));
  NAND3X1 g02287(.A(n3747), .B(P1_REG3_REG_23__SCAN_IN), .C(P1_REG3_REG_22__SCAN_IN), .Y(n3832));
  XOR2X1  g02288(.A(n3832), .B(P1_REG3_REG_24__SCAN_IN), .Y(n3833));
  AOI22X1 g02289(.A0(n2730), .A1(P1_REG0_REG_24__SCAN_IN), .B0(P1_REG2_REG_24__SCAN_IN), .B1(n2731), .Y(n3834));
  INVX1   g02290(.A(n3834), .Y(n3835));
  AOI21X1 g02291(.A0(n2734), .A1(P1_REG1_REG_24__SCAN_IN), .B0(n3835), .Y(n3836));
  OAI21X1 g02292(.A0(n3833), .A1(n2708), .B0(n3836), .Y(n3837));
  INVX1   g02293(.A(n3837), .Y(n3838));
  OAI22X1 g02294(.A0(n3815), .A1(n2744), .B0(n2791), .B1(n3838), .Y(n3839));
  AOI21X1 g02295(.A0(n3831), .A1(n2740), .B0(n3839), .Y(n3840));
  OAI21X1 g02296(.A0(n3822), .A1(n2728), .B0(n3840), .Y(n3841));
  NOR2X1  g02297(.A(n3841), .B(n3829), .Y(n3842));
  NAND2X1 g02298(.A(n2679), .B(P1_REG0_REG_23__SCAN_IN), .Y(n3843));
  OAI21X1 g02299(.A0(n3842), .A1(n2679), .B0(n3843), .Y(P1_U3519));
  NOR2X1  g02300(.A(n2684), .B(n2358), .Y(n3845));
  OAI21X1 g02301(.A0(n3803), .A1(n3765), .B0(n3816), .Y(n3848));
  NAND2X1 g02302(.A(n3848), .B(n3809), .Y(n3849));
  NOR3X1  g02303(.A(n3808), .B(n3803), .C(n3764), .Y(n3850));
  INVX1   g02304(.A(n3850), .Y(n3851));
  OAI21X1 g02305(.A0(n3851), .A1(n3724), .B0(n3849), .Y(n3852));
  XOR2X1  g02306(.A(n3852), .B(n3864), .Y(n3853));
  INVX1   g02307(.A(n3853), .Y(n3854));
  NAND2X1 g02308(.A(n3854), .B(n2721), .Y(n3855));
  NOR3X1  g02309(.A(n3795), .B(n2684), .C(n2332), .Y(n3856));
  OAI21X1 g02310(.A0(n2684), .A1(n2332), .B0(n3795), .Y(n3857));
  AOI21X1 g02311(.A0(n3857), .A1(n3821), .B0(n3856), .Y(n3858));
  NAND2X1 g02312(.A(n3858), .B(n3864), .Y(n3859));
  NAND2X1 g02313(.A(n2377), .B(n2375), .Y(n3860));
  XOR2X1  g02314(.A(n2356), .B(n3860), .Y(n3861));
  NOR2X1  g02315(.A(n3861), .B(n1837), .Y(n3862));
  OAI21X1 g02316(.A0(n3862), .A1(n2346), .B0(n2810), .Y(n3863));
  XOR2X1  g02317(.A(n3863), .B(n3838), .Y(n3864));
  OAI21X1 g02318(.A0(n3864), .A1(n3858), .B0(n3859), .Y(n3865));
  AOI22X1 g02319(.A0(n3794), .A1(n2786), .B0(n2724), .B1(n3865), .Y(n3866));
  OAI21X1 g02320(.A0(n2725), .A1(n2751), .B0(n3865), .Y(n3867));
  NAND3X1 g02321(.A(n3867), .B(n3866), .C(n3855), .Y(n3868));
  NOR2X1  g02322(.A(n3853), .B(n2716), .Y(n3869));
  AOI21X1 g02323(.A0(n3289), .A1(n3288), .B0(n3853), .Y(n3870));
  NAND4X1 g02324(.A(n2673), .B(n2656), .C(n2660), .D(n3865), .Y(n3871));
  NOR3X1  g02325(.A(n3804), .B(n3761), .C(n3783), .Y(n3872));
  XOR2X1  g02326(.A(n3863), .B(n3872), .Y(n3873));
  NAND4X1 g02327(.A(P1_REG3_REG_23__SCAN_IN), .B(P1_REG3_REG_24__SCAN_IN), .C(P1_REG3_REG_22__SCAN_IN), .D(n3747), .Y(n3874));
  XOR2X1  g02328(.A(n3874), .B(P1_REG3_REG_25__SCAN_IN), .Y(n3875));
  AOI22X1 g02329(.A0(n2730), .A1(P1_REG0_REG_25__SCAN_IN), .B0(P1_REG2_REG_25__SCAN_IN), .B1(n2731), .Y(n3876));
  INVX1   g02330(.A(n3876), .Y(n3877));
  AOI21X1 g02331(.A0(n2734), .A1(P1_REG1_REG_25__SCAN_IN), .B0(n3877), .Y(n3878));
  OAI21X1 g02332(.A0(n3875), .A1(n2708), .B0(n3878), .Y(n3879));
  INVX1   g02333(.A(n3879), .Y(n3880));
  OAI22X1 g02334(.A0(n3863), .A1(n2744), .B0(n2791), .B1(n3880), .Y(n3881));
  AOI21X1 g02335(.A0(n3873), .A1(n2740), .B0(n3881), .Y(n3882));
  NAND2X1 g02336(.A(n3882), .B(n3871), .Y(n3883));
  NOR4X1  g02337(.A(n3870), .B(n3869), .C(n3868), .D(n3883), .Y(n3884));
  NAND2X1 g02338(.A(n2679), .B(P1_REG0_REG_24__SCAN_IN), .Y(n3885));
  OAI21X1 g02339(.A0(n3884), .A1(n2679), .B0(n3885), .Y(P1_U3520));
  NOR2X1  g02340(.A(n2684), .B(n2384), .Y(n3887));
  XOR2X1  g02341(.A(n3887), .B(n3880), .Y(n3888));
  NOR3X1  g02342(.A(n3837), .B(n2684), .C(n2358), .Y(n3889));
  INVX1   g02343(.A(n3889), .Y(n3890));
  NOR2X1  g02344(.A(n3845), .B(n3838), .Y(n3891));
  AOI21X1 g02345(.A0(n3852), .A1(n3890), .B0(n3891), .Y(n3892));
  XOR2X1  g02346(.A(n3892), .B(n3888), .Y(n3893));
  INVX1   g02347(.A(n3893), .Y(n3894));
  NAND2X1 g02348(.A(n3894), .B(n2721), .Y(n3895));
  NOR2X1  g02349(.A(n3845), .B(n3837), .Y(n3896));
  NOR3X1  g02350(.A(n3838), .B(n2684), .C(n2358), .Y(n3897));
  INVX1   g02351(.A(n3897), .Y(n3898));
  OAI21X1 g02352(.A0(n3896), .A1(n3858), .B0(n3898), .Y(n3899));
  NAND2X1 g02353(.A(n3888), .B(n3899), .Y(n3901));
  OAI21X1 g02354(.A0(n3899), .A1(n3888), .B0(n3901), .Y(n3902));
  AOI22X1 g02355(.A0(n3837), .A1(n2786), .B0(n2724), .B1(n3902), .Y(n3903));
  OAI21X1 g02356(.A0(n2725), .A1(n2751), .B0(n3902), .Y(n3904));
  NAND3X1 g02357(.A(n3904), .B(n3903), .C(n3895), .Y(n3905));
  NOR2X1  g02358(.A(n3893), .B(n2716), .Y(n3906));
  AOI21X1 g02359(.A0(n3289), .A1(n3288), .B0(n3893), .Y(n3907));
  NAND4X1 g02360(.A(n2673), .B(n2656), .C(n2660), .D(n3902), .Y(n3908));
  NAND2X1 g02361(.A(n3863), .B(n3872), .Y(n3909));
  XOR2X1  g02362(.A(n3887), .B(n3909), .Y(n3910));
  INVX1   g02363(.A(n2372), .Y(n3911));
  NAND2X1 g02364(.A(n2403), .B(n2401), .Y(n3912));
  XOR2X1  g02365(.A(n2382), .B(n3912), .Y(n3913));
  OAI21X1 g02366(.A0(n3913), .A1(n1837), .B0(n3911), .Y(n3914));
  NAND2X1 g02367(.A(n2810), .B(n3914), .Y(n3915));
  INVX1   g02368(.A(P1_REG3_REG_26__SCAN_IN), .Y(n3916));
  INVX1   g02369(.A(P1_REG3_REG_25__SCAN_IN), .Y(n3917));
  NOR2X1  g02370(.A(n3874), .B(n3917), .Y(n3918));
  XOR2X1  g02371(.A(n3918), .B(n3916), .Y(n3919));
  AOI22X1 g02372(.A0(n2730), .A1(P1_REG0_REG_26__SCAN_IN), .B0(P1_REG2_REG_26__SCAN_IN), .B1(n2731), .Y(n3920));
  INVX1   g02373(.A(n3920), .Y(n3921));
  AOI21X1 g02374(.A0(n2734), .A1(P1_REG1_REG_26__SCAN_IN), .B0(n3921), .Y(n3922));
  OAI21X1 g02375(.A0(n3919), .A1(n2708), .B0(n3922), .Y(n3923));
  INVX1   g02376(.A(n3923), .Y(n3924));
  OAI22X1 g02377(.A0(n3915), .A1(n2744), .B0(n2791), .B1(n3924), .Y(n3925));
  AOI21X1 g02378(.A0(n3910), .A1(n2740), .B0(n3925), .Y(n3926));
  NAND2X1 g02379(.A(n3926), .B(n3908), .Y(n3927));
  NOR4X1  g02380(.A(n3907), .B(n3906), .C(n3905), .D(n3927), .Y(n3928));
  NAND2X1 g02381(.A(n2679), .B(P1_REG0_REG_25__SCAN_IN), .Y(n3929));
  OAI21X1 g02382(.A0(n3928), .A1(n2679), .B0(n3929), .Y(P1_U3521));
  INVX1   g02383(.A(n2390), .Y(n3931));
  NOR3X1  g02384(.A(n2398), .B(n2404), .C(n2392), .Y(n3932));
  AOI21X1 g02385(.A0(n2395), .A1(n2393), .B0(n2399), .Y(n3933));
  OAI21X1 g02386(.A0(n3933), .A1(n3932), .B0(n1790), .Y(n3934));
  AOI21X1 g02387(.A0(n3934), .A1(n3931), .B0(n2684), .Y(n3935));
  XOR2X1  g02388(.A(n3935), .B(n3924), .Y(n3936));
  NOR3X1  g02389(.A(n3879), .B(n2684), .C(n2384), .Y(n3937));
  INVX1   g02390(.A(n3937), .Y(n3938));
  AOI21X1 g02391(.A0(n2810), .A1(n3914), .B0(n3880), .Y(n3939));
  INVX1   g02392(.A(n3891), .Y(n3940));
  INVX1   g02393(.A(n3720), .Y(n3941));
  OAI21X1 g02394(.A0(n3680), .A1(n3717), .B0(n3941), .Y(n3942));
  AOI22X1 g02395(.A0(n3848), .A1(n3809), .B0(n3942), .B1(n3850), .Y(n3943));
  OAI21X1 g02396(.A0(n3943), .A1(n3889), .B0(n3940), .Y(n3944));
  AOI21X1 g02397(.A0(n3944), .A1(n3938), .B0(n3939), .Y(n3945));
  XOR2X1  g02398(.A(n3945), .B(n3936), .Y(n3946));
  NOR3X1  g02399(.A(n3880), .B(n2684), .C(n2384), .Y(n3947));
  NOR2X1  g02400(.A(n3947), .B(n3899), .Y(n3948));
  AOI21X1 g02401(.A0(n2810), .A1(n3914), .B0(n3879), .Y(n3949));
  OAI21X1 g02402(.A0(n2406), .A1(n2390), .B0(n2810), .Y(n3950));
  AOI21X1 g02403(.A0(n3950), .A1(n3924), .B0(n3949), .Y(n3951));
  NAND2X1 g02404(.A(n3935), .B(n3923), .Y(n3952));
  NAND2X1 g02405(.A(n3952), .B(n3951), .Y(n3953));
  INVX1   g02406(.A(n3899), .Y(n3954));
  NOR2X1  g02407(.A(n3949), .B(n3954), .Y(n3955));
  OAI21X1 g02408(.A0(n3915), .A1(n3880), .B0(n3936), .Y(n3956));
  OAI22X1 g02409(.A0(n3955), .A1(n3956), .B0(n3953), .B1(n3948), .Y(n3957));
  OAI22X1 g02410(.A0(n3880), .A1(n2854), .B0(n2723), .B1(n3957), .Y(n3958));
  AOI21X1 g02411(.A0(n2875), .A1(n2717), .B0(n3957), .Y(n3959));
  NOR2X1  g02412(.A(n3959), .B(n3958), .Y(n3960));
  OAI21X1 g02413(.A0(n3946), .A1(n3252), .B0(n3960), .Y(n3961));
  NOR2X1  g02414(.A(n3946), .B(n2716), .Y(n3962));
  AOI21X1 g02415(.A0(n3289), .A1(n3288), .B0(n3946), .Y(n3963));
  NOR2X1  g02416(.A(n3887), .B(n3909), .Y(n3964));
  XOR2X1  g02417(.A(n3950), .B(n3964), .Y(n3965));
  INVX1   g02418(.A(P1_REG3_REG_27__SCAN_IN), .Y(n3966));
  NOR3X1  g02419(.A(n3874), .B(n3917), .C(n3916), .Y(n3967));
  XOR2X1  g02420(.A(n3967), .B(n3966), .Y(n3968));
  AOI22X1 g02421(.A0(n2730), .A1(P1_REG0_REG_27__SCAN_IN), .B0(P1_REG2_REG_27__SCAN_IN), .B1(n2731), .Y(n3969));
  INVX1   g02422(.A(n3969), .Y(n3970));
  AOI21X1 g02423(.A0(n2734), .A1(P1_REG1_REG_27__SCAN_IN), .B0(n3970), .Y(n3971));
  OAI21X1 g02424(.A0(n3968), .A1(n2708), .B0(n3971), .Y(n3972));
  INVX1   g02425(.A(n3972), .Y(n3973));
  OAI22X1 g02426(.A0(n3950), .A1(n2744), .B0(n2791), .B1(n3973), .Y(n3974));
  AOI21X1 g02427(.A0(n3965), .A1(n2740), .B0(n3974), .Y(n3975));
  OAI21X1 g02428(.A0(n3957), .A1(n2728), .B0(n3975), .Y(n3976));
  NOR4X1  g02429(.A(n3963), .B(n3962), .C(n3961), .D(n3976), .Y(n3977));
  NAND2X1 g02430(.A(n2679), .B(P1_REG0_REG_26__SCAN_IN), .Y(n3978));
  OAI21X1 g02431(.A0(n3977), .A1(n2679), .B0(n3978), .Y(P1_U3522));
  NOR2X1  g02432(.A(n3935), .B(n3924), .Y(n3980));
  INVX1   g02433(.A(n3980), .Y(n3981));
  NOR2X1  g02434(.A(n3950), .B(n3923), .Y(n3982));
  INVX1   g02435(.A(n3982), .Y(n3983));
  INVX1   g02436(.A(n2422), .Y(n3984));
  NOR3X1  g02437(.A(n2430), .B(n2433), .C(n2424), .Y(n3985));
  AOI21X1 g02438(.A0(n2427), .A1(n2425), .B0(n2431), .Y(n3986));
  OAI21X1 g02439(.A0(n3986), .A1(n3985), .B0(n1790), .Y(n3987));
  AOI21X1 g02440(.A0(n3987), .A1(n3984), .B0(n2684), .Y(n3988));
  XOR2X1  g02441(.A(n3988), .B(n3973), .Y(n3989));
  NAND2X1 g02442(.A(n5478), .B(n3983), .Y(n3991));
  AOI21X1 g02443(.A0(n3945), .A1(n3981), .B0(n3991), .Y(n3992));
  INVX1   g02444(.A(n3939), .Y(n3993));
  OAI21X1 g02445(.A0(n3892), .A1(n3937), .B0(n3993), .Y(n3994));
  NAND2X1 g02446(.A(n3989), .B(n3981), .Y(n3995));
  AOI21X1 g02447(.A0(n3994), .A1(n3983), .B0(n3995), .Y(n3996));
  OAI21X1 g02448(.A0(n3996), .A1(n3992), .B0(n2721), .Y(n3997));
  OAI21X1 g02449(.A0(n3947), .A1(n3897), .B0(n3951), .Y(n3998));
  NOR2X1  g02450(.A(n3896), .B(n3858), .Y(n3999));
  AOI22X1 g02451(.A0(n3935), .A1(n3923), .B0(n3999), .B1(n3951), .Y(n4000));
  NAND2X1 g02452(.A(n4000), .B(n3998), .Y(n4001));
  XOR2X1  g02453(.A(n4001), .B(n3989), .Y(n4002));
  INVX1   g02454(.A(n4002), .Y(n4003));
  AOI22X1 g02455(.A0(n3923), .A1(n2786), .B0(n2724), .B1(n4003), .Y(n4004));
  OAI21X1 g02456(.A0(n2725), .A1(n2751), .B0(n4003), .Y(n4005));
  NAND3X1 g02457(.A(n4005), .B(n4004), .C(n3997), .Y(n4006));
  NOR2X1  g02458(.A(n3996), .B(n3992), .Y(n4007));
  NOR2X1  g02459(.A(n4007), .B(n2716), .Y(n4008));
  AOI21X1 g02460(.A0(n3289), .A1(n3288), .B0(n4007), .Y(n4009));
  NOR3X1  g02461(.A(n3935), .B(n3887), .C(n3909), .Y(n4010));
  OAI21X1 g02462(.A0(n2435), .A1(n2422), .B0(n2810), .Y(n4011));
  XOR2X1  g02463(.A(n4011), .B(n4010), .Y(n4012));
  INVX1   g02464(.A(P1_REG3_REG_28__SCAN_IN), .Y(n4013));
  NOR4X1  g02465(.A(n3966), .B(n3917), .C(n3916), .D(n3874), .Y(n4014));
  XOR2X1  g02466(.A(n4014), .B(n4013), .Y(n4015));
  AOI22X1 g02467(.A0(n2730), .A1(P1_REG0_REG_28__SCAN_IN), .B0(P1_REG2_REG_28__SCAN_IN), .B1(n2731), .Y(n4016));
  INVX1   g02468(.A(n4016), .Y(n4017));
  AOI21X1 g02469(.A0(n2734), .A1(P1_REG1_REG_28__SCAN_IN), .B0(n4017), .Y(n4018));
  OAI21X1 g02470(.A0(n4015), .A1(n2708), .B0(n4018), .Y(n4019));
  INVX1   g02471(.A(n4019), .Y(n4020));
  OAI22X1 g02472(.A0(n4011), .A1(n2744), .B0(n2791), .B1(n4020), .Y(n4021));
  AOI21X1 g02473(.A0(n4012), .A1(n2740), .B0(n4021), .Y(n4022));
  OAI21X1 g02474(.A0(n4002), .A1(n2728), .B0(n4022), .Y(n4023));
  NOR4X1  g02475(.A(n4009), .B(n4008), .C(n4006), .D(n4023), .Y(n4024));
  NAND2X1 g02476(.A(n2679), .B(P1_REG0_REG_27__SCAN_IN), .Y(n4025));
  OAI21X1 g02477(.A0(n4024), .A1(n2679), .B0(n4025), .Y(P1_U3523));
  INVX1   g02478(.A(n2442), .Y(n4027));
  NOR3X1  g02479(.A(n2449), .B(n2445), .C(n2444), .Y(n4028));
  INVX1   g02480(.A(n2449), .Y(n4029));
  AOI21X1 g02481(.A0(n2480), .A1(n2478), .B0(n4029), .Y(n4030));
  OAI21X1 g02482(.A0(n4030), .A1(n4028), .B0(n1790), .Y(n4031));
  AOI21X1 g02483(.A0(n4031), .A1(n4027), .B0(n2684), .Y(n4032));
  XOR2X1  g02484(.A(n4032), .B(n4020), .Y(n4033));
  OAI21X1 g02485(.A0(n3972), .A1(n3980), .B0(n4011), .Y(n4034));
  OAI21X1 g02486(.A0(n3973), .A1(n3981), .B0(n4034), .Y(n4035));
  NOR2X1  g02487(.A(n4011), .B(n3972), .Y(n4036));
  NOR3X1  g02488(.A(n4036), .B(n3945), .C(n3982), .Y(n4037));
  NOR2X1  g02489(.A(n4037), .B(n4035), .Y(n4038));
  XOR2X1  g02490(.A(n4038), .B(n4033), .Y(n4039));
  NOR2X1  g02491(.A(n4039), .B(n3252), .Y(n4040));
  NOR2X1  g02492(.A(n3988), .B(n3972), .Y(n4042));
  NAND2X1 g02493(.A(n3988), .B(n3972), .Y(n4043));
  OAI21X1 g02494(.A0(n4042), .A1(n3998), .B0(n4043), .Y(n4044));
  AOI21X1 g02495(.A0(n4011), .A1(n3973), .B0(n3952), .Y(n4045));
  OAI22X1 g02496(.A0(n3923), .A1(n3935), .B0(n3887), .B1(n3879), .Y(n4046));
  NOR4X1  g02497(.A(n4046), .B(n3896), .C(n3858), .D(n4042), .Y(n4047));
  NOR3X1  g02498(.A(n4047), .B(n4045), .C(n4044), .Y(n4048));
  XOR2X1  g02499(.A(n4048), .B(n5477), .Y(n4049));
  INVX1   g02500(.A(n4049), .Y(n4050));
  AOI22X1 g02501(.A0(n3972), .A1(n2786), .B0(n2724), .B1(n4050), .Y(n4051));
  OAI21X1 g02502(.A0(n2725), .A1(n2751), .B0(n4050), .Y(n4052));
  NAND2X1 g02503(.A(n4052), .B(n4051), .Y(n4053));
  XOR2X1  g02504(.A(n4038), .B(n5477), .Y(n4054));
  OAI21X1 g02505(.A0(n2720), .A1(n2714), .B0(n4054), .Y(n4055));
  OAI21X1 g02506(.A0(n4039), .A1(n2716), .B0(n4055), .Y(n4056));
  NAND2X1 g02507(.A(n4011), .B(n4010), .Y(n4057));
  XOR2X1  g02508(.A(n4032), .B(n4057), .Y(n4058));
  INVX1   g02509(.A(n4032), .Y(n4059));
  NAND4X1 g02510(.A(n2735), .B(P1_REG3_REG_27__SCAN_IN), .C(P1_REG3_REG_28__SCAN_IN), .D(n3967), .Y(n4060));
  NAND2X1 g02511(.A(n2730), .B(P1_REG0_REG_29__SCAN_IN), .Y(n4061));
  AOI22X1 g02512(.A0(n2731), .A1(P1_REG2_REG_29__SCAN_IN), .B0(P1_REG1_REG_29__SCAN_IN), .B1(n2734), .Y(n4062));
  NAND3X1 g02513(.A(n4062), .B(n4061), .C(n4060), .Y(n4063));
  INVX1   g02514(.A(n4063), .Y(n4064));
  OAI22X1 g02515(.A0(n4059), .A1(n2744), .B0(n2791), .B1(n4064), .Y(n4065));
  AOI21X1 g02516(.A0(n4058), .A1(n2740), .B0(n4065), .Y(n4066));
  OAI21X1 g02517(.A0(n4049), .A1(n2728), .B0(n4066), .Y(n4067));
  NOR4X1  g02518(.A(n4056), .B(n4053), .C(n4040), .D(n4067), .Y(n4068));
  NAND2X1 g02519(.A(n2679), .B(P1_REG0_REG_28__SCAN_IN), .Y(n4069));
  OAI21X1 g02520(.A0(n4068), .A1(n2679), .B0(n4069), .Y(P1_U3524));
  NOR3X1  g02521(.A(n4019), .B(n2684), .C(n2451), .Y(n4071));
  OAI21X1 g02522(.A0(n2483), .A1(n2467), .B0(n2810), .Y(n4072));
  XOR2X1  g02523(.A(n4072), .B(n4063), .Y(n4073));
  NOR2X1  g02524(.A(n4073), .B(n4071), .Y(n4074));
  OAI21X1 g02525(.A0(n4037), .A1(n4035), .B0(n4074), .Y(n4075));
  NAND2X1 g02526(.A(n3994), .B(n3983), .Y(n4076));
  NOR2X1  g02527(.A(n4032), .B(n4020), .Y(n4077));
  XOR2X1  g02528(.A(n4072), .B(n4064), .Y(n4078));
  NOR3X1  g02529(.A(n4078), .B(n4035), .C(n4077), .Y(n4079));
  OAI21X1 g02530(.A0(n4076), .A1(n4036), .B0(n4079), .Y(n4080));
  NOR3X1  g02531(.A(n4078), .B(n4059), .C(n4019), .Y(n4081));
  AOI21X1 g02532(.A0(n4078), .A1(n4077), .B0(n4081), .Y(n4082));
  NAND3X1 g02533(.A(n4082), .B(n4080), .C(n4075), .Y(n4083));
  NAND2X1 g02534(.A(n4083), .B(n2721), .Y(n4084));
  NOR2X1  g02535(.A(n4048), .B(n4059), .Y(n4085));
  AOI21X1 g02536(.A0(n4048), .A1(n4059), .B0(n4020), .Y(n4086));
  NOR2X1  g02537(.A(n4086), .B(n4085), .Y(n4087));
  XOR2X1  g02538(.A(n4087), .B(n4078), .Y(n4088));
  NOR2X1  g02539(.A(n4088), .B(n2723), .Y(n4089));
  NOR2X1  g02540(.A(n2658), .B(n2660), .Y(n4090));
  NOR3X1  g02541(.A(n2683), .B(n2682), .C(P1_B_REG_SCAN_IN), .Y(n4091));
  OAI21X1 g02542(.A0(n4091), .A1(n2684), .B0(n4090), .Y(n4092));
  INVX1   g02543(.A(P1_REG1_REG_30__SCAN_IN), .Y(n4093));
  NOR2X1  g02544(.A(n2707), .B(n4093), .Y(n4094));
  INVX1   g02545(.A(P1_REG2_REG_30__SCAN_IN), .Y(n4095));
  NOR4X1  g02546(.A(n2699), .B(n2703), .C(n4095), .D(n2700), .Y(n4096));
  INVX1   g02547(.A(P1_REG0_REG_30__SCAN_IN), .Y(n4097));
  NOR4X1  g02548(.A(n2699), .B(n2698), .C(n4097), .D(n2700), .Y(n4098));
  NOR3X1  g02549(.A(n4098), .B(n4096), .C(n4094), .Y(n4099));
  OAI22X1 g02550(.A0(n4092), .A1(n4099), .B0(n4020), .B1(n2854), .Y(n4100));
  AOI21X1 g02551(.A0(n2875), .A1(n2717), .B0(n4088), .Y(n4101));
  NOR3X1  g02552(.A(n4101), .B(n4100), .C(n4089), .Y(n4102));
  NAND2X1 g02553(.A(n4102), .B(n4084), .Y(n4103));
  NAND2X1 g02554(.A(n4083), .B(n2715), .Y(n4104));
  OAI21X1 g02555(.A0(n2720), .A1(n2714), .B0(n4083), .Y(n4105));
  NAND2X1 g02556(.A(n4105), .B(n4104), .Y(n4106));
  NOR2X1  g02557(.A(n4088), .B(n2728), .Y(n4107));
  NOR2X1  g02558(.A(n4032), .B(n4057), .Y(n4108));
  INVX1   g02559(.A(n2467), .Y(n4109));
  NOR3X1  g02560(.A(n2475), .B(n2481), .C(n2469), .Y(n4110));
  AOI21X1 g02561(.A0(n2472), .A1(n2470), .B0(n2476), .Y(n4111));
  OAI21X1 g02562(.A0(n4111), .A1(n4110), .B0(n1790), .Y(n4112));
  AOI21X1 g02563(.A0(n4112), .A1(n4109), .B0(n2684), .Y(n4113));
  XOR2X1  g02564(.A(n4113), .B(n4108), .Y(n4114));
  OAI22X1 g02565(.A0(n4072), .A1(n2744), .B0(n2741), .B1(n4114), .Y(n4115));
  NOR4X1  g02566(.A(n4107), .B(n4106), .C(n4103), .D(n4115), .Y(n4116));
  NAND2X1 g02567(.A(n2679), .B(P1_REG0_REG_29__SCAN_IN), .Y(n4117));
  OAI21X1 g02568(.A0(n4116), .A1(n2679), .B0(n4117), .Y(P1_U3525));
  NAND2X1 g02569(.A(n4072), .B(n4108), .Y(n4119));
  INVX1   g02570(.A(n2503), .Y(n4120));
  NAND3X1 g02571(.A(n4120), .B(n2499), .C(n2497), .Y(n4121));
  OAI21X1 g02572(.A0(n2520), .A1(n2496), .B0(n2503), .Y(n4122));
  AOI21X1 g02573(.A0(n4122), .A1(n4121), .B0(n1837), .Y(n4123));
  OAI21X1 g02574(.A0(n4123), .A1(n2493), .B0(n2810), .Y(n4124));
  INVX1   g02575(.A(n4124), .Y(n4125));
  XOR2X1  g02576(.A(n4125), .B(n4119), .Y(n4126));
  INVX1   g02577(.A(P1_REG1_REG_31__SCAN_IN), .Y(n4127));
  NOR2X1  g02578(.A(n2707), .B(n4127), .Y(n4128));
  INVX1   g02579(.A(P1_REG2_REG_31__SCAN_IN), .Y(n4129));
  NOR4X1  g02580(.A(n2699), .B(n2703), .C(n4129), .D(n2700), .Y(n4130));
  INVX1   g02581(.A(P1_REG0_REG_31__SCAN_IN), .Y(n4131));
  NOR4X1  g02582(.A(n2699), .B(n2698), .C(n4131), .D(n2700), .Y(n4132));
  NOR3X1  g02583(.A(n4132), .B(n4130), .C(n4128), .Y(n4133));
  NOR2X1  g02584(.A(n4133), .B(n4092), .Y(n4134));
  INVX1   g02585(.A(n4134), .Y(n4135));
  OAI21X1 g02586(.A0(n4124), .A1(n2744), .B0(n4135), .Y(n4136));
  AOI21X1 g02587(.A0(n4126), .A1(n2740), .B0(n4136), .Y(n4137));
  NAND2X1 g02588(.A(n2679), .B(P1_REG0_REG_30__SCAN_IN), .Y(n4138));
  OAI21X1 g02589(.A0(n4137), .A1(n2679), .B0(n4138), .Y(P1_U3526));
  AOI21X1 g02590(.A0(n2810), .A1(n2505), .B0(n4119), .Y(n4140));
  OAI21X1 g02591(.A0(n2528), .A1(n2512), .B0(n2810), .Y(n4141));
  XOR2X1  g02592(.A(n4141), .B(n4140), .Y(n4142));
  OAI21X1 g02593(.A0(n4141), .A1(n2744), .B0(n4135), .Y(n4143));
  AOI21X1 g02594(.A0(n4142), .A1(n2740), .B0(n4143), .Y(n4144));
  NAND2X1 g02595(.A(n2679), .B(P1_REG0_REG_31__SCAN_IN), .Y(n4145));
  OAI21X1 g02596(.A0(n4144), .A1(n2679), .B0(n4145), .Y(P1_U3527));
  NOR2X1  g02597(.A(n2678), .B(n2561), .Y(n4147));
  NAND2X1 g02598(.A(n4147), .B(n2676), .Y(n4148));
  NAND2X1 g02599(.A(n4148), .B(P1_REG1_REG_0__SCAN_IN), .Y(n4149));
  OAI21X1 g02600(.A0(n4148), .A1(n2748), .B0(n4149), .Y(P1_U3528));
  NAND2X1 g02601(.A(n4148), .B(P1_REG1_REG_1__SCAN_IN), .Y(n4151));
  OAI21X1 g02602(.A0(n4148), .A1(n2803), .B0(n4151), .Y(P1_U3529));
  NAND2X1 g02603(.A(n4148), .B(P1_REG1_REG_2__SCAN_IN), .Y(n4153));
  OAI21X1 g02604(.A0(n4148), .A1(n2851), .B0(n4153), .Y(P1_U3530));
  NAND2X1 g02605(.A(n4148), .B(P1_REG1_REG_3__SCAN_IN), .Y(n4155));
  OAI21X1 g02606(.A0(n4148), .A1(n2902), .B0(n4155), .Y(P1_U3531));
  NAND2X1 g02607(.A(n4148), .B(P1_REG1_REG_4__SCAN_IN), .Y(n4157));
  OAI21X1 g02608(.A0(n4148), .A1(n2950), .B0(n4157), .Y(P1_U3532));
  NAND2X1 g02609(.A(n4148), .B(P1_REG1_REG_5__SCAN_IN), .Y(n4159));
  OAI21X1 g02610(.A0(n4148), .A1(n3000), .B0(n4159), .Y(P1_U3533));
  NAND2X1 g02611(.A(n4148), .B(P1_REG1_REG_6__SCAN_IN), .Y(n4161));
  OAI21X1 g02612(.A0(n4148), .A1(n3054), .B0(n4161), .Y(P1_U3534));
  NAND2X1 g02613(.A(n4148), .B(P1_REG1_REG_7__SCAN_IN), .Y(n4163));
  OAI21X1 g02614(.A0(n4148), .A1(n3108), .B0(n4163), .Y(P1_U3535));
  NAND2X1 g02615(.A(n4148), .B(P1_REG1_REG_8__SCAN_IN), .Y(n4165));
  OAI21X1 g02616(.A0(n4148), .A1(n3157), .B0(n4165), .Y(P1_U3536));
  NAND2X1 g02617(.A(n4148), .B(P1_REG1_REG_9__SCAN_IN), .Y(n4167));
  OAI21X1 g02618(.A0(n4148), .A1(n3203), .B0(n4167), .Y(P1_U3537));
  NAND2X1 g02619(.A(n4148), .B(P1_REG1_REG_10__SCAN_IN), .Y(n4169));
  OAI21X1 g02620(.A0(n4148), .A1(n3249), .B0(n4169), .Y(P1_U3538));
  NAND2X1 g02621(.A(n4148), .B(P1_REG1_REG_11__SCAN_IN), .Y(n4171));
  OAI21X1 g02622(.A0(n4148), .A1(n3303), .B0(n4171), .Y(P1_U3539));
  NAND2X1 g02623(.A(n4148), .B(P1_REG1_REG_12__SCAN_IN), .Y(n4173));
  OAI21X1 g02624(.A0(n4148), .A1(n3350), .B0(n4173), .Y(P1_U3540));
  NAND2X1 g02625(.A(n4148), .B(P1_REG1_REG_13__SCAN_IN), .Y(n4175));
  OAI21X1 g02626(.A0(n4148), .A1(n3402), .B0(n4175), .Y(P1_U3541));
  NAND2X1 g02627(.A(n4148), .B(P1_REG1_REG_14__SCAN_IN), .Y(n4177));
  OAI21X1 g02628(.A0(n4148), .A1(n3445), .B0(n4177), .Y(P1_U3542));
  NAND2X1 g02629(.A(n4148), .B(P1_REG1_REG_15__SCAN_IN), .Y(n4179));
  OAI21X1 g02630(.A0(n4148), .A1(n3486), .B0(n4179), .Y(P1_U3543));
  NAND2X1 g02631(.A(n4148), .B(P1_REG1_REG_16__SCAN_IN), .Y(n4181));
  OAI21X1 g02632(.A0(n4148), .A1(n3536), .B0(n4181), .Y(P1_U3544));
  NAND2X1 g02633(.A(n4148), .B(P1_REG1_REG_17__SCAN_IN), .Y(n4183));
  OAI21X1 g02634(.A0(n4148), .A1(n3582), .B0(n4183), .Y(P1_U3545));
  NAND2X1 g02635(.A(n4148), .B(P1_REG1_REG_18__SCAN_IN), .Y(n4185));
  OAI21X1 g02636(.A0(n4148), .A1(n3623), .B0(n4185), .Y(P1_U3546));
  NAND2X1 g02637(.A(n4148), .B(P1_REG1_REG_19__SCAN_IN), .Y(n4187));
  OAI21X1 g02638(.A0(n4148), .A1(n3670), .B0(n4187), .Y(P1_U3547));
  NAND2X1 g02639(.A(n4148), .B(P1_REG1_REG_20__SCAN_IN), .Y(n4189));
  OAI21X1 g02640(.A0(n4148), .A1(n3712), .B0(n4189), .Y(P1_U3548));
  NAND2X1 g02641(.A(n4148), .B(P1_REG1_REG_21__SCAN_IN), .Y(n4191));
  OAI21X1 g02642(.A0(n4148), .A1(n3758), .B0(n4191), .Y(P1_U3549));
  NAND2X1 g02643(.A(n4148), .B(P1_REG1_REG_22__SCAN_IN), .Y(n4193));
  OAI21X1 g02644(.A0(n4148), .A1(n3799), .B0(n4193), .Y(P1_U3550));
  NAND2X1 g02645(.A(n4148), .B(P1_REG1_REG_23__SCAN_IN), .Y(n4195));
  OAI21X1 g02646(.A0(n4148), .A1(n3842), .B0(n4195), .Y(P1_U3551));
  NAND2X1 g02647(.A(n4148), .B(P1_REG1_REG_24__SCAN_IN), .Y(n4197));
  OAI21X1 g02648(.A0(n4148), .A1(n3884), .B0(n4197), .Y(P1_U3552));
  NAND2X1 g02649(.A(n4148), .B(P1_REG1_REG_25__SCAN_IN), .Y(n4199));
  OAI21X1 g02650(.A0(n4148), .A1(n3928), .B0(n4199), .Y(P1_U3553));
  NAND2X1 g02651(.A(n4148), .B(P1_REG1_REG_26__SCAN_IN), .Y(n4201));
  OAI21X1 g02652(.A0(n4148), .A1(n3977), .B0(n4201), .Y(P1_U3554));
  NAND2X1 g02653(.A(n4148), .B(P1_REG1_REG_27__SCAN_IN), .Y(n4203));
  OAI21X1 g02654(.A0(n4148), .A1(n4024), .B0(n4203), .Y(P1_U3555));
  NAND2X1 g02655(.A(n4148), .B(P1_REG1_REG_28__SCAN_IN), .Y(n4205));
  OAI21X1 g02656(.A0(n4148), .A1(n4068), .B0(n4205), .Y(P1_U3556));
  NAND2X1 g02657(.A(n4148), .B(P1_REG1_REG_29__SCAN_IN), .Y(n4207));
  OAI21X1 g02658(.A0(n4148), .A1(n4116), .B0(n4207), .Y(P1_U3557));
  NAND2X1 g02659(.A(n4148), .B(P1_REG1_REG_30__SCAN_IN), .Y(n4209));
  OAI21X1 g02660(.A0(n4148), .A1(n4137), .B0(n4209), .Y(P1_U3558));
  NAND2X1 g02661(.A(n4148), .B(P1_REG1_REG_31__SCAN_IN), .Y(n4211));
  OAI21X1 g02662(.A0(n4148), .A1(n4144), .B0(n4211), .Y(P1_U3559));
  NOR4X1  g02663(.A(n2668), .B(n2666), .C(n2654), .D(n2713), .Y(n4213));
  INVX1   g02664(.A(n4213), .Y(n4214));
  NOR2X1  g02665(.A(n2673), .B(n2666), .Y(n4215));
  NOR3X1  g02666(.A(n4215), .B(n2658), .C(n2660), .Y(n4216));
  NOR2X1  g02667(.A(n4216), .B(n2650), .Y(n4217));
  NAND3X1 g02668(.A(n4217), .B(n2678), .C(n2647), .Y(n4218));
  NAND2X1 g02669(.A(n4218), .B(n4214), .Y(n4219));
  NAND4X1 g02670(.A(n2737), .B(n2729), .C(n2560), .D(n4219), .Y(n4220));
  NAND2X1 g02671(.A(n4219), .B(n2560), .Y(n4221));
  INVX1   g02672(.A(n4221), .Y(n4222));
  AOI21X1 g02673(.A0(n4219), .A1(n2560), .B0(n2702), .Y(n4223));
  AOI21X1 g02674(.A0(n4222), .A1(n2727), .B0(n4223), .Y(n4224));
  NAND3X1 g02675(.A(n2658), .B(n2666), .C(n2660), .Y(n4225));
  NOR2X1  g02676(.A(n4225), .B(n4221), .Y(n4226));
  NAND3X1 g02677(.A(n2673), .B(n2668), .C(n2656), .Y(n4227));
  NOR2X1  g02678(.A(n4227), .B(n4221), .Y(n4228));
  AOI22X1 g02679(.A0(n4226), .A1(n2693), .B0(n5490), .B1(n4228), .Y(n4229));
  NAND3X1 g02680(.A(n2713), .B(n2658), .C(n2660), .Y(n4230));
  NOR3X1  g02681(.A(n4221), .B(n4230), .C(n2666), .Y(n4231));
  NOR2X1  g02682(.A(n4221), .B(n4214), .Y(n4232));
  AOI22X1 g02683(.A0(n4231), .A1(n2693), .B0(P1_REG3_REG_0__SCAN_IN), .B1(n4232), .Y(n4233));
  NAND4X1 g02684(.A(n4229), .B(n4224), .C(n4220), .D(n4233), .Y(P1_U3293));
  NAND4X1 g02685(.A(n2824), .B(n2729), .C(n2560), .D(n4219), .Y(n4235));
  AOI21X1 g02686(.A0(n4219), .A1(n2560), .B0(n2774), .Y(n4236));
  AOI21X1 g02687(.A0(n4222), .A1(n2789), .B0(n4236), .Y(n4237));
  AOI22X1 g02688(.A0(n4226), .A1(n2757), .B0(n2771), .B1(n4228), .Y(n4238));
  AOI22X1 g02689(.A0(n4231), .A1(n2790), .B0(P1_REG3_REG_1__SCAN_IN), .B1(n4232), .Y(n4239));
  NAND4X1 g02690(.A(n4238), .B(n4237), .C(n4235), .D(n4239), .Y(P1_U3292));
  AOI22X1 g02691(.A0(n4228), .A1(n2830), .B0(P1_REG3_REG_2__SCAN_IN), .B1(n4232), .Y(n4241));
  AOI22X1 g02692(.A0(n4226), .A1(n2827), .B0(n2842), .B1(n4231), .Y(n4242));
  NAND2X1 g02693(.A(n4222), .B(n2839), .Y(n4243));
  NOR2X1  g02694(.A(n4221), .B(n2791), .Y(n4244));
  AOI22X1 g02695(.A0(n4221), .A1(P1_REG2_REG_2__SCAN_IN), .B0(n2859), .B1(n4244), .Y(n4245));
  NAND4X1 g02696(.A(n4243), .B(n4242), .C(n4241), .D(n4245), .Y(P1_U3291));
  NOR3X1  g02697(.A(n2889), .B(n2876), .C(n2874), .Y(n4247));
  INVX1   g02698(.A(P1_REG2_REG_3__SCAN_IN), .Y(n4248));
  INVX1   g02699(.A(n4244), .Y(n4249));
  OAI22X1 g02700(.A0(n4222), .A1(n4248), .B0(n2898), .B1(n4249), .Y(n4250));
  INVX1   g02701(.A(n4228), .Y(n4251));
  INVX1   g02702(.A(n4232), .Y(n4252));
  OAI22X1 g02703(.A0(n4251), .A1(n2873), .B0(P1_REG3_REG_3__SCAN_IN), .B1(n4252), .Y(n4253));
  INVX1   g02704(.A(n4226), .Y(n4254));
  NOR4X1  g02705(.A(n2668), .B(n2666), .C(n2654), .D(n2673), .Y(n4255));
  NAND4X1 g02706(.A(n4219), .B(n2891), .C(n2560), .D(n4255), .Y(n4256));
  OAI21X1 g02707(.A0(n4254), .A1(n2866), .B0(n4256), .Y(n4257));
  NOR3X1  g02708(.A(n4257), .B(n4253), .C(n4250), .Y(n4258));
  OAI21X1 g02709(.A0(n4221), .A1(n4247), .B0(n4258), .Y(P1_U3290));
  NOR3X1  g02710(.A(n2936), .B(n2933), .C(n2925), .Y(n4260));
  INVX1   g02711(.A(P1_REG2_REG_4__SCAN_IN), .Y(n4261));
  OAI22X1 g02712(.A0(n4222), .A1(n4261), .B0(n2946), .B1(n4249), .Y(n4262));
  OAI22X1 g02713(.A0(n4251), .A1(n2924), .B0(n2896), .B1(n4252), .Y(n4263));
  NAND4X1 g02714(.A(n4219), .B(n2939), .C(n2560), .D(n4255), .Y(n4264));
  OAI21X1 g02715(.A0(n4254), .A1(n2938), .B0(n4264), .Y(n4265));
  NOR3X1  g02716(.A(n4265), .B(n4263), .C(n4262), .Y(n4266));
  OAI21X1 g02717(.A0(n4221), .A1(n4260), .B0(n4266), .Y(P1_U3289));
  NAND2X1 g02718(.A(n4222), .B(n2987), .Y(n4268));
  INVX1   g02719(.A(P1_REG2_REG_5__SCAN_IN), .Y(n4269));
  OAI22X1 g02720(.A0(n4222), .A1(n4269), .B0(n2998), .B1(n4249), .Y(n4270));
  OAI22X1 g02721(.A0(n4251), .A1(n2977), .B0(n2944), .B1(n4252), .Y(n4271));
  INVX1   g02722(.A(n4231), .Y(n4272));
  OAI22X1 g02723(.A0(n4254), .A1(n2969), .B0(n2990), .B1(n4272), .Y(n4273));
  NOR3X1  g02724(.A(n4273), .B(n4271), .C(n4270), .Y(n4274));
  NAND2X1 g02725(.A(n4274), .B(n4268), .Y(P1_U3288));
  NOR3X1  g02726(.A(n3039), .B(n3022), .C(n3021), .Y(n4276));
  INVX1   g02727(.A(n2996), .Y(n4277));
  AOI22X1 g02728(.A0(n4231), .A1(n3043), .B0(n4277), .B1(n4232), .Y(n4278));
  OAI21X1 g02729(.A0(n4254), .A1(n3042), .B0(n4278), .Y(n4279));
  AOI22X1 g02730(.A0(n4221), .A1(P1_REG2_REG_6__SCAN_IN), .B0(n3049), .B1(n4244), .Y(n4280));
  OAI21X1 g02731(.A0(n4251), .A1(n3020), .B0(n4280), .Y(n4281));
  NOR2X1  g02732(.A(n4281), .B(n4279), .Y(n4282));
  OAI21X1 g02733(.A0(n4221), .A1(n4276), .B0(n4282), .Y(P1_U3287));
  NOR3X1  g02734(.A(n3093), .B(n3077), .C(n3076), .Y(n4284));
  AOI22X1 g02735(.A0(n4221), .A1(P1_REG2_REG_7__SCAN_IN), .B0(n3103), .B1(n4244), .Y(n4285));
  INVX1   g02736(.A(n4225), .Y(n4286));
  NAND4X1 g02737(.A(n4219), .B(n3067), .C(n2560), .D(n4286), .Y(n4287));
  AOI22X1 g02738(.A0(n4231), .A1(n3095), .B0(n3047), .B1(n4232), .Y(n4288));
  NAND3X1 g02739(.A(n4288), .B(n4287), .C(n4285), .Y(n4289));
  AOI21X1 g02740(.A0(n4228), .A1(n3074), .B0(n4289), .Y(n4290));
  OAI21X1 g02741(.A0(n4221), .A1(n4284), .B0(n4290), .Y(P1_U3286));
  NOR3X1  g02742(.A(n3140), .B(n3127), .C(n3126), .Y(n4292));
  NOR2X1  g02743(.A(n4251), .B(n3125), .Y(n4293));
  AOI22X1 g02744(.A0(n4221), .A1(P1_REG2_REG_8__SCAN_IN), .B0(n3170), .B1(n4244), .Y(n4294));
  NAND4X1 g02745(.A(n4219), .B(n3120), .C(n2560), .D(n4286), .Y(n4295));
  AOI22X1 g02746(.A0(n4231), .A1(n3144), .B0(n3101), .B1(n4232), .Y(n4296));
  NAND3X1 g02747(.A(n4296), .B(n4295), .C(n4294), .Y(n4297));
  NOR2X1  g02748(.A(n4297), .B(n4293), .Y(n4298));
  OAI21X1 g02749(.A0(n4221), .A1(n4292), .B0(n4298), .Y(P1_U3285));
  NAND2X1 g02750(.A(n4222), .B(n3186), .Y(n4300));
  NAND2X1 g02751(.A(n4231), .B(n3188), .Y(n4301));
  AOI22X1 g02752(.A0(n4221), .A1(P1_REG2_REG_9__SCAN_IN), .B0(n3167), .B1(n4226), .Y(n4302));
  AOI22X1 g02753(.A0(n4244), .A1(n3213), .B0(n3148), .B1(n4232), .Y(n4303));
  NAND3X1 g02754(.A(n4303), .B(n4302), .C(n4301), .Y(n4304));
  AOI21X1 g02755(.A0(n4228), .A1(n3174), .B0(n4304), .Y(n4305));
  NAND2X1 g02756(.A(n4305), .B(n4300), .Y(P1_U3284));
  NOR3X1  g02757(.A(n3233), .B(n3225), .C(n3224), .Y(n4307));
  NAND2X1 g02758(.A(n4231), .B(n3237), .Y(n4308));
  AOI22X1 g02759(.A0(n4221), .A1(P1_REG2_REG_10__SCAN_IN), .B0(n3215), .B1(n4226), .Y(n4309));
  AOI22X1 g02760(.A0(n4244), .A1(n3266), .B0(n3194), .B1(n4232), .Y(n4310));
  NAND3X1 g02761(.A(n4310), .B(n4309), .C(n4308), .Y(n4311));
  AOI21X1 g02762(.A0(n4228), .A1(n3222), .B0(n4311), .Y(n4312));
  OAI21X1 g02763(.A0(n4221), .A1(n4307), .B0(n4312), .Y(P1_U3283));
  NOR2X1  g02764(.A(n3272), .B(n3252), .Y(n4314));
  INVX1   g02765(.A(n3285), .Y(n4315));
  NOR4X1  g02766(.A(n3287), .B(n4315), .C(n4314), .D(n3290), .Y(n4316));
  NOR2X1  g02767(.A(n4251), .B(n3281), .Y(n4317));
  NAND2X1 g02768(.A(n4231), .B(n3291), .Y(n4318));
  AOI22X1 g02769(.A0(n4221), .A1(P1_REG2_REG_11__SCAN_IN), .B0(n3365), .B1(n4244), .Y(n4319));
  AOI22X1 g02770(.A0(n4226), .A1(n3259), .B0(n3240), .B1(n4232), .Y(n4320));
  NAND3X1 g02771(.A(n4320), .B(n4319), .C(n4318), .Y(n4321));
  NOR2X1  g02772(.A(n4321), .B(n4317), .Y(n4322));
  OAI21X1 g02773(.A0(n4221), .A1(n4316), .B0(n4322), .Y(P1_U3282));
  NAND2X1 g02774(.A(n4222), .B(n3335), .Y(n4324));
  NAND2X1 g02775(.A(n4231), .B(n3339), .Y(n4325));
  AOI22X1 g02776(.A0(n4221), .A1(P1_REG2_REG_12__SCAN_IN), .B0(n3345), .B1(n4244), .Y(n4326));
  AOI22X1 g02777(.A0(n4226), .A1(n3313), .B0(n3294), .B1(n4232), .Y(n4327));
  NAND3X1 g02778(.A(n4327), .B(n4326), .C(n4325), .Y(n4328));
  AOI21X1 g02779(.A0(n4228), .A1(n3318), .B0(n4328), .Y(n4329));
  NAND2X1 g02780(.A(n4329), .B(n4324), .Y(P1_U3281));
  NOR3X1  g02781(.A(n3386), .B(n3373), .C(n3372), .Y(n4331));
  NOR2X1  g02782(.A(n4251), .B(n3371), .Y(n4332));
  NAND2X1 g02783(.A(n4231), .B(n3389), .Y(n4333));
  AOI22X1 g02784(.A0(n4221), .A1(P1_REG2_REG_13__SCAN_IN), .B0(n3405), .B1(n4244), .Y(n4334));
  AOI22X1 g02785(.A0(n4226), .A1(n3358), .B0(n3342), .B1(n4232), .Y(n4335));
  NAND3X1 g02786(.A(n4335), .B(n4334), .C(n4333), .Y(n4336));
  NOR2X1  g02787(.A(n4336), .B(n4332), .Y(n4337));
  OAI21X1 g02788(.A0(n4221), .A1(n4331), .B0(n4337), .Y(P1_U3280));
  INVX1   g02789(.A(P1_REG2_REG_14__SCAN_IN), .Y(n4339));
  OAI22X1 g02790(.A0(n4222), .A1(n4339), .B0(n3443), .B1(n4249), .Y(n4340));
  OAI22X1 g02791(.A0(n4254), .A1(n3410), .B0(n3393), .B1(n4252), .Y(n4341));
  NOR2X1  g02792(.A(n4341), .B(n4340), .Y(n4342));
  OAI21X1 g02793(.A0(n4272), .A1(n3434), .B0(n4342), .Y(n4343));
  AOI21X1 g02794(.A0(n4228), .A1(n3422), .B0(n4343), .Y(n4344));
  OAI21X1 g02795(.A0(n4221), .A1(n3428), .B0(n4344), .Y(P1_U3279));
  NAND2X1 g02796(.A(n4231), .B(n3473), .Y(n4346));
  AOI22X1 g02797(.A0(n4221), .A1(P1_REG2_REG_15__SCAN_IN), .B0(n3452), .B1(n4226), .Y(n4347));
  AOI22X1 g02798(.A0(n4244), .A1(n3503), .B0(n3439), .B1(n4232), .Y(n4348));
  NAND3X1 g02799(.A(n4348), .B(n4347), .C(n4346), .Y(n4349));
  AOI21X1 g02800(.A0(n4228), .A1(n3465), .B0(n4349), .Y(n4350));
  OAI21X1 g02801(.A0(n4221), .A1(n3471), .B0(n4350), .Y(P1_U3278));
  NOR3X1  g02802(.A(n3523), .B(n3522), .C(n3521), .Y(n4352));
  NAND2X1 g02803(.A(n4231), .B(n3525), .Y(n4353));
  AOI22X1 g02804(.A0(n4221), .A1(P1_REG2_REG_16__SCAN_IN), .B0(n3496), .B1(n4226), .Y(n4354));
  AOI22X1 g02805(.A0(n4244), .A1(n3541), .B0(n3478), .B1(n4232), .Y(n4355));
  NAND3X1 g02806(.A(n4355), .B(n4354), .C(n4353), .Y(n4356));
  AOI21X1 g02807(.A0(n4228), .A1(n3518), .B0(n4356), .Y(n4357));
  OAI21X1 g02808(.A0(n4221), .A1(n4352), .B0(n4357), .Y(P1_U3277));
  NOR3X1  g02809(.A(n3569), .B(n3565), .C(n3557), .Y(n4359));
  NOR2X1  g02810(.A(n4251), .B(n3556), .Y(n4360));
  NAND2X1 g02811(.A(n4231), .B(n3571), .Y(n4361));
  AOI22X1 g02812(.A0(n4221), .A1(P1_REG2_REG_17__SCAN_IN), .B0(n3588), .B1(n4244), .Y(n4362));
  OAI21X1 g02813(.A0(n4252), .A1(n3527), .B0(n4362), .Y(n4363));
  AOI21X1 g02814(.A0(n4226), .A1(n3547), .B0(n4363), .Y(n4364));
  NAND2X1 g02815(.A(n4364), .B(n4361), .Y(n4365));
  NOR2X1  g02816(.A(n4365), .B(n4360), .Y(n4366));
  OAI21X1 g02817(.A0(n4221), .A1(n4359), .B0(n4366), .Y(P1_U3276));
  NAND2X1 g02818(.A(n4222), .B(n3609), .Y(n4368));
  AOI22X1 g02819(.A0(n4221), .A1(P1_REG2_REG_18__SCAN_IN), .B0(n3684), .B1(n4244), .Y(n4369));
  OAI21X1 g02820(.A0(n4252), .A1(n3573), .B0(n4369), .Y(n4370));
  AOI21X1 g02821(.A0(n4226), .A1(n3640), .B0(n4370), .Y(n4371));
  OAI21X1 g02822(.A0(n4272), .A1(n3613), .B0(n4371), .Y(n4372));
  AOI21X1 g02823(.A0(n4228), .A1(n3599), .B0(n4372), .Y(n4373));
  NAND2X1 g02824(.A(n4373), .B(n4368), .Y(P1_U3275));
  NAND2X1 g02825(.A(n4222), .B(n3655), .Y(n4375));
  INVX1   g02826(.A(n3648), .Y(n4376));
  NAND2X1 g02827(.A(n4228), .B(n4376), .Y(n4377));
  NAND2X1 g02828(.A(n4231), .B(n3656), .Y(n4378));
  AOI22X1 g02829(.A0(n4221), .A1(P1_REG2_REG_19__SCAN_IN), .B0(n3617), .B1(n4232), .Y(n4379));
  OAI21X1 g02830(.A0(n4249), .A1(n3666), .B0(n4379), .Y(n4380));
  AOI21X1 g02831(.A0(n4226), .A1(n3627), .B0(n4380), .Y(n4381));
  NAND4X1 g02832(.A(n4378), .B(n4377), .C(n4375), .D(n4381), .Y(P1_U3274));
  NAND2X1 g02833(.A(n4222), .B(n3698), .Y(n4383));
  INVX1   g02834(.A(n3661), .Y(n4384));
  AOI22X1 g02835(.A0(n4221), .A1(P1_REG2_REG_20__SCAN_IN), .B0(n4384), .B1(n4232), .Y(n4385));
  OAI21X1 g02836(.A0(n4249), .A1(n3710), .B0(n4385), .Y(n4386));
  AOI21X1 g02837(.A0(n4226), .A1(n3719), .B0(n4386), .Y(n4387));
  OAI21X1 g02838(.A0(n4272), .A1(n3701), .B0(n4387), .Y(n4388));
  AOI21X1 g02839(.A0(n4228), .A1(n3692), .B0(n4388), .Y(n4389));
  NAND2X1 g02840(.A(n4389), .B(n4383), .Y(P1_U3273));
  NAND2X1 g02841(.A(n4222), .B(n3743), .Y(n4391));
  NAND3X1 g02842(.A(n4228), .B(n3735), .C(n3733), .Y(n4392));
  NAND2X1 g02843(.A(n4231), .B(n3746), .Y(n4393));
  INVX1   g02844(.A(n3705), .Y(n4394));
  AOI22X1 g02845(.A0(n4221), .A1(P1_REG2_REG_21__SCAN_IN), .B0(n4394), .B1(n4232), .Y(n4395));
  OAI21X1 g02846(.A0(n4249), .A1(n3754), .B0(n4395), .Y(n4396));
  AOI21X1 g02847(.A0(n4226), .A1(n3715), .B0(n4396), .Y(n4397));
  NAND4X1 g02848(.A(n4393), .B(n4392), .C(n4391), .D(n4397), .Y(P1_U3272));
  NOR3X1  g02849(.A(n3782), .B(n3781), .C(n3780), .Y(n4399));
  NAND2X1 g02850(.A(n4231), .B(n3784), .Y(n4400));
  AOI22X1 g02851(.A0(n4221), .A1(P1_REG2_REG_22__SCAN_IN), .B0(n3748), .B1(n4232), .Y(n4401));
  OAI21X1 g02852(.A0(n4249), .A1(n3795), .B0(n4401), .Y(n4402));
  AOI21X1 g02853(.A0(n4226), .A1(n3761), .B0(n4402), .Y(n4403));
  NAND2X1 g02854(.A(n4403), .B(n4400), .Y(n4404));
  AOI21X1 g02855(.A0(n4228), .A1(n3777), .B0(n4404), .Y(n4405));
  OAI21X1 g02856(.A0(n4221), .A1(n4399), .B0(n4405), .Y(P1_U3271));
  NAND2X1 g02857(.A(n4222), .B(n3829), .Y(n4407));
  INVX1   g02858(.A(n3822), .Y(n4408));
  NAND2X1 g02859(.A(n4228), .B(n4408), .Y(n4409));
  NAND2X1 g02860(.A(n4231), .B(n3831), .Y(n4410));
  INVX1   g02861(.A(n3790), .Y(n4411));
  AOI22X1 g02862(.A0(n4221), .A1(P1_REG2_REG_23__SCAN_IN), .B0(n4411), .B1(n4232), .Y(n4412));
  OAI21X1 g02863(.A0(n4249), .A1(n3838), .B0(n4412), .Y(n4413));
  AOI21X1 g02864(.A0(n4226), .A1(n3804), .B0(n4413), .Y(n4414));
  NAND4X1 g02865(.A(n4410), .B(n4409), .C(n4407), .D(n4414), .Y(P1_U3270));
  NOR3X1  g02866(.A(n3870), .B(n3869), .C(n3868), .Y(n4416));
  NAND2X1 g02867(.A(n4231), .B(n3873), .Y(n4417));
  INVX1   g02868(.A(n3833), .Y(n4418));
  AOI22X1 g02869(.A0(n4221), .A1(P1_REG2_REG_24__SCAN_IN), .B0(n4418), .B1(n4232), .Y(n4419));
  OAI21X1 g02870(.A0(n4249), .A1(n3880), .B0(n4419), .Y(n4420));
  AOI21X1 g02871(.A0(n4226), .A1(n3845), .B0(n4420), .Y(n4421));
  NAND2X1 g02872(.A(n4421), .B(n4417), .Y(n4422));
  AOI21X1 g02873(.A0(n4228), .A1(n3865), .B0(n4422), .Y(n4423));
  OAI21X1 g02874(.A0(n4221), .A1(n4416), .B0(n4423), .Y(P1_U3269));
  NOR3X1  g02875(.A(n3907), .B(n3906), .C(n3905), .Y(n4425));
  NAND2X1 g02876(.A(n4231), .B(n3910), .Y(n4426));
  INVX1   g02877(.A(n3875), .Y(n4427));
  AOI22X1 g02878(.A0(n4221), .A1(P1_REG2_REG_25__SCAN_IN), .B0(n4427), .B1(n4232), .Y(n4428));
  OAI21X1 g02879(.A0(n4249), .A1(n3924), .B0(n4428), .Y(n4429));
  AOI21X1 g02880(.A0(n4226), .A1(n3887), .B0(n4429), .Y(n4430));
  NAND2X1 g02881(.A(n4430), .B(n4426), .Y(n4431));
  AOI21X1 g02882(.A0(n4228), .A1(n3902), .B0(n4431), .Y(n4432));
  OAI21X1 g02883(.A0(n4221), .A1(n4425), .B0(n4432), .Y(P1_U3268));
  NOR3X1  g02884(.A(n3963), .B(n3962), .C(n3961), .Y(n4434));
  NOR2X1  g02885(.A(n4251), .B(n3957), .Y(n4435));
  NAND2X1 g02886(.A(n4231), .B(n3965), .Y(n4436));
  INVX1   g02887(.A(n3919), .Y(n4437));
  AOI22X1 g02888(.A0(n4221), .A1(P1_REG2_REG_26__SCAN_IN), .B0(n4437), .B1(n4232), .Y(n4438));
  OAI21X1 g02889(.A0(n4249), .A1(n3973), .B0(n4438), .Y(n4439));
  AOI21X1 g02890(.A0(n4226), .A1(n3935), .B0(n4439), .Y(n4440));
  NAND2X1 g02891(.A(n4440), .B(n4436), .Y(n4441));
  NOR2X1  g02892(.A(n4441), .B(n4435), .Y(n4442));
  OAI21X1 g02893(.A0(n4221), .A1(n4434), .B0(n4442), .Y(P1_U3267));
  NOR3X1  g02894(.A(n4009), .B(n4008), .C(n4006), .Y(n4444));
  NAND2X1 g02895(.A(n4231), .B(n4012), .Y(n4445));
  INVX1   g02896(.A(n3968), .Y(n4446));
  AOI22X1 g02897(.A0(n4221), .A1(P1_REG2_REG_27__SCAN_IN), .B0(n4446), .B1(n4232), .Y(n4447));
  OAI21X1 g02898(.A0(n4249), .A1(n4020), .B0(n4447), .Y(n4448));
  AOI21X1 g02899(.A0(n4226), .A1(n3988), .B0(n4448), .Y(n4449));
  NAND2X1 g02900(.A(n4449), .B(n4445), .Y(n4450));
  AOI21X1 g02901(.A0(n4228), .A1(n4003), .B0(n4450), .Y(n4451));
  OAI21X1 g02902(.A0(n4221), .A1(n4444), .B0(n4451), .Y(P1_U3266));
  NOR3X1  g02903(.A(n4056), .B(n4053), .C(n4040), .Y(n4453));
  NAND2X1 g02904(.A(n4231), .B(n4058), .Y(n4454));
  INVX1   g02905(.A(n4015), .Y(n4455));
  AOI22X1 g02906(.A0(n4221), .A1(P1_REG2_REG_28__SCAN_IN), .B0(n4455), .B1(n4232), .Y(n4456));
  OAI21X1 g02907(.A0(n4249), .A1(n4064), .B0(n4456), .Y(n4457));
  AOI21X1 g02908(.A0(n4226), .A1(n4032), .B0(n4457), .Y(n4458));
  NAND2X1 g02909(.A(n4458), .B(n4454), .Y(n4459));
  AOI21X1 g02910(.A0(n4228), .A1(n4050), .B0(n4459), .Y(n4460));
  OAI21X1 g02911(.A0(n4221), .A1(n4453), .B0(n4460), .Y(P1_U3265));
  OAI21X1 g02912(.A0(n4106), .A1(n4103), .B0(n4222), .Y(n4462));
  NOR2X1  g02913(.A(n4251), .B(n4088), .Y(n4463));
  NAND2X1 g02914(.A(n4221), .B(P1_REG2_REG_29__SCAN_IN), .Y(n4464));
  NAND4X1 g02915(.A(n3967), .B(P1_REG3_REG_27__SCAN_IN), .C(P1_REG3_REG_28__SCAN_IN), .D(n4232), .Y(n4465));
  NAND2X1 g02916(.A(n4465), .B(n4464), .Y(n4466));
  AOI21X1 g02917(.A0(n4226), .A1(n4113), .B0(n4466), .Y(n4467));
  OAI21X1 g02918(.A0(n4272), .A1(n4114), .B0(n4467), .Y(n4468));
  NOR2X1  g02919(.A(n4468), .B(n4463), .Y(n4469));
  NAND2X1 g02920(.A(n4469), .B(n4462), .Y(P1_U3356));
  NAND2X1 g02921(.A(n4231), .B(n4126), .Y(n4471));
  NAND3X1 g02922(.A(n4219), .B(n4134), .C(n2560), .Y(n4472));
  OAI21X1 g02923(.A0(n4222), .A1(n4095), .B0(n4472), .Y(n4473));
  AOI21X1 g02924(.A0(n4226), .A1(n4125), .B0(n4473), .Y(n4474));
  NAND2X1 g02925(.A(n4474), .B(n4471), .Y(P1_U3264));
  NAND2X1 g02926(.A(n4231), .B(n4142), .Y(n4476));
  INVX1   g02927(.A(n2512), .Y(n4477));
  OAI21X1 g02928(.A0(n2520), .A1(n2496), .B0(n2517), .Y(n4478));
  NOR3X1  g02929(.A(n2522), .B(n2521), .C(n2496), .Y(n4479));
  NAND2X1 g02930(.A(n4479), .B(n2499), .Y(n4480));
  NAND4X1 g02931(.A(n4480), .B(n4478), .C(n1790), .D(n2526), .Y(n4481));
  AOI21X1 g02932(.A0(n4481), .A1(n4477), .B0(n2684), .Y(n4482));
  OAI21X1 g02933(.A0(n4222), .A1(n4129), .B0(n4472), .Y(n4483));
  AOI21X1 g02934(.A0(n4226), .A1(n4482), .B0(n4483), .Y(n4484));
  NAND2X1 g02935(.A(n4484), .B(n4476), .Y(P1_U3263));
  NOR2X1  g02936(.A(P1_IR_REG_31__SCAN_IN), .B(n2339), .Y(n4486));
  AOI21X1 g02937(.A0(n2342), .A1(P1_IR_REG_31__SCAN_IN), .B0(n4486), .Y(n4487));
  NOR2X1  g02938(.A(n4090), .B(n2538), .Y(n4488));
  NOR2X1  g02939(.A(n4488), .B(n2540), .Y(n4489));
  OAI21X1 g02940(.A0(n4489), .A1(n2684), .B0(P1_STATE_REG_SCAN_IN), .Y(P1_U3085));
  AOI21X1 g02941(.A0(n4487), .A1(n2538), .B0(P1_U3085), .Y(n4491));
  NOR2X1  g02942(.A(n4491), .B(n2561), .Y(n4492));
  INVX1   g02943(.A(P1_REG2_REG_18__SCAN_IN), .Y(n4493));
  INVX1   g02944(.A(P1_REG2_REG_16__SCAN_IN), .Y(n4494));
  INVX1   g02945(.A(P1_REG2_REG_17__SCAN_IN), .Y(n4495));
  AOI22X1 g02946(.A0(n3493), .A1(n4494), .B0(n4495), .B1(n3543), .Y(n4496));
  NOR2X1  g02947(.A(n3450), .B(P1_REG2_REG_15__SCAN_IN), .Y(n4497));
  NOR2X1  g02948(.A(n3407), .B(n4339), .Y(n4498));
  NAND2X1 g02949(.A(n3407), .B(n4339), .Y(n4499));
  INVX1   g02950(.A(P1_REG2_REG_11__SCAN_IN), .Y(n4500));
  NOR2X1  g02951(.A(n3256), .B(n4500), .Y(n4501));
  INVX1   g02952(.A(n4501), .Y(n4502));
  INVX1   g02953(.A(P1_REG2_REG_12__SCAN_IN), .Y(n4503));
  INVX1   g02954(.A(P1_REG2_REG_13__SCAN_IN), .Y(n4504));
  AOI22X1 g02955(.A0(n3310), .A1(n4503), .B0(n4504), .B1(n3355), .Y(n4505));
  INVX1   g02956(.A(n4505), .Y(n4506));
  NOR2X1  g02957(.A(n3310), .B(n4503), .Y(n4507));
  AOI21X1 g02958(.A0(n3356), .A1(P1_REG2_REG_13__SCAN_IN), .B0(n4507), .Y(n4508));
  OAI21X1 g02959(.A0(n4506), .A1(n4502), .B0(n4508), .Y(n4509));
  OAI21X1 g02960(.A0(n3356), .A1(P1_REG2_REG_13__SCAN_IN), .B0(n4509), .Y(n4510));
  INVX1   g02961(.A(P1_REG2_REG_10__SCAN_IN), .Y(n4511));
  INVX1   g02962(.A(P1_REG2_REG_8__SCAN_IN), .Y(n4512));
  NOR2X1  g02963(.A(n3117), .B(n4512), .Y(n4513));
  INVX1   g02964(.A(P1_REG2_REG_9__SCAN_IN), .Y(n4514));
  AOI22X1 g02965(.A0(n3164), .A1(n4514), .B0(n4511), .B1(n3208), .Y(n4515));
  NAND2X1 g02966(.A(n3165), .B(P1_REG2_REG_9__SCAN_IN), .Y(n4516));
  OAI21X1 g02967(.A0(n3208), .A1(n4511), .B0(n4516), .Y(n4517));
  AOI21X1 g02968(.A0(n4515), .A1(n4513), .B0(n4517), .Y(n4518));
  AOI21X1 g02969(.A0(n3208), .A1(n4511), .B0(n4518), .Y(n4519));
  INVX1   g02970(.A(P1_REG2_REG_6__SCAN_IN), .Y(n4520));
  INVX1   g02971(.A(P1_REG2_REG_7__SCAN_IN), .Y(n4521));
  AOI22X1 g02972(.A0(n3004), .A1(n4520), .B0(n4521), .B1(n3061), .Y(n4522));
  AOI22X1 g02973(.A0(n2917), .A1(n4261), .B0(n4269), .B1(n2962), .Y(n4523));
  INVX1   g02974(.A(n2864), .Y(n4524));
  OAI22X1 g02975(.A0(n2825), .A1(P1_REG2_REG_2__SCAN_IN), .B0(P1_REG2_REG_3__SCAN_IN), .B1(n4524), .Y(n4525));
  NOR2X1  g02976(.A(n2219), .B(n2702), .Y(n4526));
  INVX1   g02977(.A(n4526), .Y(n4527));
  AOI21X1 g02978(.A0(n2754), .A1(n2774), .B0(n4527), .Y(n4528));
  NOR2X1  g02979(.A(n2754), .B(n2774), .Y(n4529));
  NOR2X1  g02980(.A(n4529), .B(n4528), .Y(n4530));
  NOR2X1  g02981(.A(n2864), .B(n4248), .Y(n4531));
  NOR2X1  g02982(.A(n4524), .B(P1_REG2_REG_3__SCAN_IN), .Y(n4532));
  NOR3X1  g02983(.A(n4532), .B(n2812), .C(n2793), .Y(n4533));
  NOR2X1  g02984(.A(n4533), .B(n4531), .Y(n4534));
  OAI21X1 g02985(.A0(n4530), .A1(n4525), .B0(n4534), .Y(n4535));
  NAND2X1 g02986(.A(n4535), .B(n4523), .Y(n4536));
  NOR2X1  g02987(.A(n2917), .B(n4261), .Y(n4537));
  AOI21X1 g02988(.A0(n2916), .A1(P1_REG2_REG_4__SCAN_IN), .B0(P1_REG2_REG_5__SCAN_IN), .Y(n4538));
  NOR2X1  g02989(.A(n4538), .B(n2962), .Y(n4539));
  AOI21X1 g02990(.A0(n4537), .A1(P1_REG2_REG_5__SCAN_IN), .B0(n4539), .Y(n4540));
  NAND2X1 g02991(.A(n4540), .B(n4536), .Y(n4541));
  NAND2X1 g02992(.A(n4541), .B(n4522), .Y(n4542));
  NOR3X1  g02993(.A(n3004), .B(n4521), .C(n4520), .Y(n4543));
  OAI21X1 g02994(.A0(n3004), .A1(n4520), .B0(n4521), .Y(n4544));
  AOI21X1 g02995(.A0(n4544), .A1(n3062), .B0(n4543), .Y(n4545));
  NAND2X1 g02996(.A(n4545), .B(n4542), .Y(n4546));
  INVX1   g02997(.A(n4515), .Y(n4547));
  INVX1   g02998(.A(n3117), .Y(n4548));
  NOR2X1  g02999(.A(n4548), .B(P1_REG2_REG_8__SCAN_IN), .Y(n4549));
  NOR2X1  g03000(.A(n4549), .B(n4547), .Y(n4550));
  AOI21X1 g03001(.A0(n4550), .A1(n4546), .B0(n4519), .Y(n4551));
  OAI21X1 g03002(.A0(n3257), .A1(P1_REG2_REG_11__SCAN_IN), .B0(n4505), .Y(n4552));
  OAI21X1 g03003(.A0(n4552), .A1(n4551), .B0(n4510), .Y(n4553));
  AOI21X1 g03004(.A0(n4553), .A1(n4499), .B0(n4498), .Y(n4554));
  NOR2X1  g03005(.A(n4554), .B(n4497), .Y(n4555));
  AOI21X1 g03006(.A0(n3450), .A1(P1_REG2_REG_15__SCAN_IN), .B0(n4555), .Y(n4556));
  INVX1   g03007(.A(n4556), .Y(n4557));
  NOR2X1  g03008(.A(n3493), .B(n4494), .Y(n4558));
  INVX1   g03009(.A(n4558), .Y(n4559));
  AOI21X1 g03010(.A0(n4559), .A1(n4495), .B0(n3543), .Y(n4560));
  AOI21X1 g03011(.A0(n4558), .A1(P1_REG2_REG_17__SCAN_IN), .B0(n4560), .Y(n4561));
  INVX1   g03012(.A(n4561), .Y(n4562));
  AOI21X1 g03013(.A0(n4557), .A1(n4496), .B0(n4562), .Y(n4563));
  OAI21X1 g03014(.A0(n3590), .A1(n4493), .B0(n4563), .Y(n4564));
  XOR2X1  g03015(.A(n2713), .B(P1_REG2_REG_19__SCAN_IN), .Y(n4565));
  AOI21X1 g03016(.A0(n3590), .A1(n4493), .B0(n4565), .Y(n4566));
  NAND2X1 g03017(.A(n4566), .B(n4564), .Y(n4567));
  AOI21X1 g03018(.A0(n3590), .A1(n4493), .B0(n4563), .Y(n4568));
  OAI21X1 g03019(.A0(n3590), .A1(n4493), .B0(n4565), .Y(n4569));
  OAI21X1 g03020(.A0(n4569), .A1(n4568), .B0(n4567), .Y(n4570));
  AOI21X1 g03021(.A0(n2666), .A1(n2654), .B0(n2668), .Y(n4571));
  OAI21X1 g03022(.A0(n2658), .A1(n2654), .B0(n2656), .Y(n4572));
  NAND3X1 g03023(.A(n4572), .B(n4571), .C(n4225), .Y(n4573));
  INVX1   g03024(.A(n4573), .Y(n4574));
  NOR2X1  g03025(.A(n2687), .B(n2686), .Y(n4575));
  INVX1   g03026(.A(n4575), .Y(n4576));
  NOR2X1  g03027(.A(n4576), .B(n4570), .Y(n4579));
  AOI22X1 g03028(.A0(n3493), .A1(n3479), .B0(n3529), .B1(n3543), .Y(n4580));
  INVX1   g03029(.A(P1_REG1_REG_13__SCAN_IN), .Y(n4581));
  NAND2X1 g03030(.A(n3355), .B(n4581), .Y(n4582));
  INVX1   g03031(.A(P1_REG1_REG_11__SCAN_IN), .Y(n4583));
  NOR2X1  g03032(.A(n3256), .B(n4583), .Y(n4584));
  INVX1   g03033(.A(n4584), .Y(n4585));
  INVX1   g03034(.A(P1_REG1_REG_12__SCAN_IN), .Y(n4586));
  AOI22X1 g03035(.A0(n3310), .A1(n4586), .B0(n4581), .B1(n3355), .Y(n4587));
  INVX1   g03036(.A(n4587), .Y(n4588));
  AOI22X1 g03037(.A0(n3311), .A1(P1_REG1_REG_12__SCAN_IN), .B0(P1_REG1_REG_13__SCAN_IN), .B1(n3356), .Y(n4589));
  OAI21X1 g03038(.A0(n4588), .A1(n4585), .B0(n4589), .Y(n4590));
  INVX1   g03039(.A(P1_REG1_REG_10__SCAN_IN), .Y(n4591));
  INVX1   g03040(.A(P1_REG1_REG_8__SCAN_IN), .Y(n4592));
  NOR2X1  g03041(.A(n3117), .B(n4592), .Y(n4593));
  INVX1   g03042(.A(P1_REG1_REG_9__SCAN_IN), .Y(n4594));
  AOI22X1 g03043(.A0(n3164), .A1(n4594), .B0(n4591), .B1(n3208), .Y(n4595));
  NAND2X1 g03044(.A(n3165), .B(P1_REG1_REG_9__SCAN_IN), .Y(n4596));
  OAI21X1 g03045(.A0(n3208), .A1(n4591), .B0(n4596), .Y(n4597));
  AOI21X1 g03046(.A0(n4595), .A1(n4593), .B0(n4597), .Y(n4598));
  AOI21X1 g03047(.A0(n3208), .A1(n4591), .B0(n4598), .Y(n4599));
  INVX1   g03048(.A(P1_REG1_REG_7__SCAN_IN), .Y(n4600));
  AOI22X1 g03049(.A0(n3004), .A1(n2994), .B0(n4600), .B1(n3061), .Y(n4601));
  AOI22X1 g03050(.A0(n2917), .A1(n2894), .B0(n2942), .B1(n2962), .Y(n4602));
  OAI22X1 g03051(.A0(n2825), .A1(P1_REG1_REG_2__SCAN_IN), .B0(P1_REG1_REG_3__SCAN_IN), .B1(n4524), .Y(n4603));
  NOR2X1  g03052(.A(n2219), .B(n2705), .Y(n4604));
  INVX1   g03053(.A(n4604), .Y(n4605));
  AOI21X1 g03054(.A0(n2754), .A1(n2778), .B0(n4605), .Y(n4606));
  NOR2X1  g03055(.A(n2754), .B(n2778), .Y(n4607));
  NOR2X1  g03056(.A(n4607), .B(n4606), .Y(n4608));
  NOR2X1  g03057(.A(n2864), .B(n2845), .Y(n4609));
  NOR2X1  g03058(.A(n4524), .B(P1_REG1_REG_3__SCAN_IN), .Y(n4610));
  NOR3X1  g03059(.A(n4610), .B(n2812), .C(n2796), .Y(n4611));
  NOR2X1  g03060(.A(n4611), .B(n4609), .Y(n4612));
  OAI21X1 g03061(.A0(n4608), .A1(n4603), .B0(n4612), .Y(n4613));
  NAND2X1 g03062(.A(n4613), .B(n4602), .Y(n4614));
  NOR2X1  g03063(.A(n2917), .B(n2894), .Y(n4615));
  AOI21X1 g03064(.A0(n2916), .A1(P1_REG1_REG_4__SCAN_IN), .B0(P1_REG1_REG_5__SCAN_IN), .Y(n4616));
  NOR2X1  g03065(.A(n4616), .B(n2962), .Y(n4617));
  AOI21X1 g03066(.A0(n4615), .A1(P1_REG1_REG_5__SCAN_IN), .B0(n4617), .Y(n4618));
  NAND2X1 g03067(.A(n4618), .B(n4614), .Y(n4619));
  NAND2X1 g03068(.A(n4619), .B(n4601), .Y(n4620));
  NOR3X1  g03069(.A(n3004), .B(n4600), .C(n2994), .Y(n4621));
  OAI21X1 g03070(.A0(n3004), .A1(n2994), .B0(n4600), .Y(n4622));
  AOI21X1 g03071(.A0(n4622), .A1(n3062), .B0(n4621), .Y(n4623));
  NAND2X1 g03072(.A(n4623), .B(n4620), .Y(n4624));
  NOR2X1  g03073(.A(n4548), .B(P1_REG1_REG_8__SCAN_IN), .Y(n4625));
  INVX1   g03074(.A(n4625), .Y(n4626));
  NAND3X1 g03075(.A(n4626), .B(n4624), .C(n4595), .Y(n4627));
  INVX1   g03076(.A(n4627), .Y(n4628));
  NOR2X1  g03077(.A(n4628), .B(n4599), .Y(n4629));
  NOR2X1  g03078(.A(n3257), .B(P1_REG1_REG_11__SCAN_IN), .Y(n4630));
  NOR3X1  g03079(.A(n4630), .B(n4629), .C(n4588), .Y(n4631));
  AOI21X1 g03080(.A0(n4590), .A1(n4582), .B0(n4631), .Y(n4632));
  AOI21X1 g03081(.A0(n3407), .A1(n3395), .B0(n4632), .Y(n4633));
  AOI21X1 g03082(.A0(n3408), .A1(P1_REG1_REG_14__SCAN_IN), .B0(n4633), .Y(n4634));
  AOI21X1 g03083(.A0(n3449), .A1(n3440), .B0(n4634), .Y(n4635));
  AOI21X1 g03084(.A0(n3450), .A1(P1_REG1_REG_15__SCAN_IN), .B0(n4635), .Y(n4636));
  INVX1   g03085(.A(n4636), .Y(n4637));
  NOR2X1  g03086(.A(n3493), .B(n3479), .Y(n4638));
  INVX1   g03087(.A(n4638), .Y(n4639));
  AOI21X1 g03088(.A0(n4639), .A1(n3529), .B0(n3543), .Y(n4640));
  AOI21X1 g03089(.A0(n4638), .A1(P1_REG1_REG_17__SCAN_IN), .B0(n4640), .Y(n4641));
  INVX1   g03090(.A(n4641), .Y(n4642));
  AOI21X1 g03091(.A0(n4637), .A1(n4580), .B0(n4642), .Y(n4643));
  INVX1   g03092(.A(n4643), .Y(n4644));
  AOI21X1 g03093(.A0(n3591), .A1(P1_REG1_REG_18__SCAN_IN), .B0(n4644), .Y(n4645));
  XOR2X1  g03094(.A(n2713), .B(P1_REG1_REG_19__SCAN_IN), .Y(n4646));
  AOI21X1 g03095(.A0(n3590), .A1(n3575), .B0(n4646), .Y(n4647));
  INVX1   g03096(.A(n4647), .Y(n4648));
  AOI21X1 g03097(.A0(n3590), .A1(n3575), .B0(n4643), .Y(n4649));
  OAI21X1 g03098(.A0(n3590), .A1(n3575), .B0(n4646), .Y(n4650));
  OAI22X1 g03099(.A0(n4649), .A1(n4650), .B0(n4648), .B1(n4645), .Y(n4651));
  INVX1   g03100(.A(n2687), .Y(n4654));
  OAI22X1 g03101(.A0(n2681), .A1(n4651), .B0(n2713), .B1(n4654), .Y(n4657));
  OAI21X1 g03102(.A0(n4657), .A1(n4579), .B0(n4492), .Y(n4658));
  NOR2X1  g03103(.A(n4487), .B(P1_U3086), .Y(n4659));
  NOR3X1  g03104(.A(n2343), .B(n4491), .C(n2681), .Y(n4661));
  INVX1   g03105(.A(n4661), .Y(n4662));
  NOR2X1  g03106(.A(n4662), .B(n4651), .Y(n4663));
  NOR3X1  g03107(.A(n2343), .B(n4576), .C(n4491), .Y(n4664));
  INVX1   g03108(.A(n4664), .Y(n4665));
  NOR3X1  g03109(.A(n2343), .B(n4491), .C(n4654), .Y(n4666));
  INVX1   g03110(.A(n4491), .Y(n4667));
  OAI22X1 g03111(.A0(P1_STATE_REG_SCAN_IN), .A1(n3659), .B0(n1718), .B1(n4667), .Y(n4668));
  AOI21X1 g03112(.A0(n4666), .A1(n2673), .B0(n4668), .Y(n4669));
  OAI21X1 g03113(.A0(n4665), .A1(n4570), .B0(n4669), .Y(n4670));
  NOR2X1  g03114(.A(n4670), .B(n4663), .Y(n4671));
  NAND2X1 g03115(.A(n4671), .B(n4658), .Y(P1_U3262));
  XOR2X1  g03116(.A(n3590), .B(P1_REG2_REG_18__SCAN_IN), .Y(n4673));
  INVX1   g03117(.A(n4673), .Y(n4674));
  XOR2X1  g03118(.A(n4674), .B(n4563), .Y(n4675));
  NOR2X1  g03119(.A(n4675), .B(n4576), .Y(n4676));
  XOR2X1  g03120(.A(n3590), .B(n3575), .Y(n4677));
  XOR2X1  g03121(.A(n4677), .B(n4643), .Y(n4678));
  OAI22X1 g03122(.A0(n4654), .A1(n3590), .B0(n2681), .B1(n4678), .Y(n4679));
  OAI21X1 g03123(.A0(n4679), .A1(n4676), .B0(n4492), .Y(n4680));
  NOR2X1  g03124(.A(n4678), .B(n4662), .Y(n4681));
  NOR2X1  g03125(.A(n4675), .B(n4665), .Y(n4682));
  INVX1   g03126(.A(n4666), .Y(n4683));
  AOI22X1 g03127(.A0(P1_U3086), .A1(P1_REG3_REG_18__SCAN_IN), .B0(P1_ADDR_REG_18__SCAN_IN), .B1(n4491), .Y(n4684));
  OAI21X1 g03128(.A0(n4683), .A1(n3590), .B0(n4684), .Y(n4685));
  NOR3X1  g03129(.A(n4685), .B(n4682), .C(n4681), .Y(n4686));
  NAND2X1 g03130(.A(n4686), .B(n4680), .Y(P1_U3261));
  INVX1   g03131(.A(n4492), .Y(n4688));
  OAI21X1 g03132(.A0(n3543), .A1(n4495), .B0(n4496), .Y(n4689));
  AOI21X1 g03133(.A0(n4559), .A1(n4556), .B0(n4689), .Y(n4690));
  NOR2X1  g03134(.A(n3494), .B(P1_REG2_REG_16__SCAN_IN), .Y(n4691));
  INVX1   g03135(.A(n4691), .Y(n4692));
  XOR2X1  g03136(.A(n3543), .B(P1_REG2_REG_17__SCAN_IN), .Y(n4693));
  OAI21X1 g03137(.A0(n3493), .A1(n4494), .B0(n4693), .Y(n4694));
  AOI21X1 g03138(.A0(n4557), .A1(n4692), .B0(n4694), .Y(n4695));
  NOR3X1  g03139(.A(n4695), .B(n4690), .C(n4576), .Y(n4696));
  OAI21X1 g03140(.A0(n3543), .A1(n3529), .B0(n4580), .Y(n4697));
  AOI21X1 g03141(.A0(n4639), .A1(n4636), .B0(n4697), .Y(n4698));
  AOI21X1 g03142(.A0(n3493), .A1(n3479), .B0(n4636), .Y(n4699));
  XOR2X1  g03143(.A(n3543), .B(n3529), .Y(n4700));
  NOR3X1  g03144(.A(n4700), .B(n4699), .C(n4638), .Y(n4701));
  NOR3X1  g03145(.A(n4701), .B(n4698), .C(n2681), .Y(n4702));
  NOR3X1  g03146(.A(n4574), .B(n3543), .C(n4654), .Y(n4703));
  NOR3X1  g03147(.A(n4703), .B(n4702), .C(n4696), .Y(n4704));
  NOR3X1  g03148(.A(n4701), .B(n4698), .C(n4662), .Y(n4705));
  NOR3X1  g03149(.A(n4695), .B(n4690), .C(n4665), .Y(n4706));
  AOI22X1 g03150(.A0(P1_U3086), .A1(P1_REG3_REG_17__SCAN_IN), .B0(P1_ADDR_REG_17__SCAN_IN), .B1(n4491), .Y(n4707));
  OAI21X1 g03151(.A0(n4683), .A1(n3543), .B0(n4707), .Y(n4708));
  NOR3X1  g03152(.A(n4708), .B(n4706), .C(n4705), .Y(n4709));
  OAI21X1 g03153(.A0(n4704), .A1(n4688), .B0(n4709), .Y(P1_U3260));
  XOR2X1  g03154(.A(n3493), .B(n4494), .Y(n4711));
  AOI21X1 g03155(.A0(n4559), .A1(n4692), .B0(n4556), .Y(n4712));
  AOI21X1 g03156(.A0(n4711), .A1(n4556), .B0(n4712), .Y(n4713));
  NOR2X1  g03157(.A(n4713), .B(n4576), .Y(n4714));
  XOR2X1  g03158(.A(n3493), .B(n3479), .Y(n4715));
  NOR2X1  g03159(.A(n4715), .B(n4636), .Y(n4717));
  AOI21X1 g03160(.A0(n4715), .A1(n4636), .B0(n4717), .Y(n4718));
  OAI22X1 g03161(.A0(n4654), .A1(n3493), .B0(n2681), .B1(n4718), .Y(n4719));
  OAI21X1 g03162(.A0(n4719), .A1(n4714), .B0(n4492), .Y(n4720));
  NOR2X1  g03163(.A(n4718), .B(n4662), .Y(n4721));
  OAI22X1 g03164(.A0(P1_STATE_REG_SCAN_IN), .A1(n3475), .B0(n1526), .B1(n4667), .Y(n4722));
  AOI21X1 g03165(.A0(n4666), .A1(n3494), .B0(n4722), .Y(n4723));
  OAI21X1 g03166(.A0(n4713), .A1(n4665), .B0(n4723), .Y(n4724));
  NOR2X1  g03167(.A(n4724), .B(n4721), .Y(n4725));
  NAND2X1 g03168(.A(n4725), .B(n4720), .Y(P1_U3259));
  XOR2X1  g03169(.A(n3449), .B(P1_REG2_REG_15__SCAN_IN), .Y(n4727));
  XOR2X1  g03170(.A(n4727), .B(n4554), .Y(n4728));
  XOR2X1  g03171(.A(n3449), .B(n3440), .Y(n4729));
  XOR2X1  g03172(.A(n4729), .B(n4634), .Y(n4730));
  OAI22X1 g03173(.A0(n4654), .A1(n3449), .B0(n2681), .B1(n4730), .Y(n4731));
  AOI21X1 g03174(.A0(n4728), .A1(n4575), .B0(n4731), .Y(n4732));
  NOR2X1  g03175(.A(n4730), .B(n4662), .Y(n4733));
  NAND2X1 g03176(.A(n4728), .B(n4664), .Y(n4734));
  OAI22X1 g03177(.A0(P1_STATE_REG_SCAN_IN), .A1(n3436), .B0(n1528), .B1(n4667), .Y(n4735));
  AOI21X1 g03178(.A0(n4666), .A1(n3450), .B0(n4735), .Y(n4736));
  NAND2X1 g03179(.A(n4736), .B(n4734), .Y(n4737));
  NOR2X1  g03180(.A(n4737), .B(n4733), .Y(n4738));
  OAI21X1 g03181(.A0(n4732), .A1(n4688), .B0(n4738), .Y(P1_U3258));
  XOR2X1  g03182(.A(n3407), .B(P1_REG2_REG_14__SCAN_IN), .Y(n4740));
  XOR2X1  g03183(.A(n4740), .B(n4553), .Y(n4741));
  NOR2X1  g03184(.A(n4741), .B(n4576), .Y(n4742));
  XOR2X1  g03185(.A(n3407), .B(n3395), .Y(n4743));
  XOR2X1  g03186(.A(n4743), .B(n4632), .Y(n4744));
  OAI22X1 g03187(.A0(n4654), .A1(n3407), .B0(n2681), .B1(n4744), .Y(n4745));
  OAI21X1 g03188(.A0(n4745), .A1(n4742), .B0(n4492), .Y(n4746));
  NOR2X1  g03189(.A(n4744), .B(n4662), .Y(n4747));
  OAI22X1 g03190(.A0(P1_STATE_REG_SCAN_IN), .A1(n3390), .B0(n1533), .B1(n4667), .Y(n4748));
  AOI21X1 g03191(.A0(n4666), .A1(n3408), .B0(n4748), .Y(n4749));
  OAI21X1 g03192(.A0(n4741), .A1(n4665), .B0(n4749), .Y(n4750));
  NOR2X1  g03193(.A(n4750), .B(n4747), .Y(n4751));
  NAND2X1 g03194(.A(n4751), .B(n4746), .Y(P1_U3257));
  INVX1   g03195(.A(n4507), .Y(n4753));
  NOR2X1  g03196(.A(n3257), .B(P1_REG2_REG_11__SCAN_IN), .Y(n4754));
  OAI21X1 g03197(.A0(n4754), .A1(n4551), .B0(n4502), .Y(n4755));
  INVX1   g03198(.A(n4755), .Y(n4756));
  OAI21X1 g03199(.A0(n3355), .A1(n4504), .B0(n4505), .Y(n4757));
  AOI21X1 g03200(.A0(n4756), .A1(n4753), .B0(n4757), .Y(n4758));
  NOR2X1  g03201(.A(n3311), .B(P1_REG2_REG_12__SCAN_IN), .Y(n4759));
  INVX1   g03202(.A(n4759), .Y(n4760));
  XOR2X1  g03203(.A(n3355), .B(P1_REG2_REG_13__SCAN_IN), .Y(n4761));
  OAI21X1 g03204(.A0(n3310), .A1(n4503), .B0(n4761), .Y(n4762));
  AOI21X1 g03205(.A0(n4755), .A1(n4760), .B0(n4762), .Y(n4763));
  NOR3X1  g03206(.A(n4763), .B(n4758), .C(n4576), .Y(n4764));
  NAND2X1 g03207(.A(n3311), .B(P1_REG1_REG_12__SCAN_IN), .Y(n4765));
  NOR2X1  g03208(.A(n4630), .B(n4629), .Y(n4766));
  NOR2X1  g03209(.A(n4766), .B(n4584), .Y(n4767));
  OAI21X1 g03210(.A0(n3355), .A1(n4581), .B0(n4587), .Y(n4768));
  AOI21X1 g03211(.A0(n4767), .A1(n4765), .B0(n4768), .Y(n4769));
  AOI21X1 g03212(.A0(n3310), .A1(n4586), .B0(n4767), .Y(n4770));
  XOR2X1  g03213(.A(n3355), .B(P1_REG1_REG_13__SCAN_IN), .Y(n4771));
  OAI21X1 g03214(.A0(n3310), .A1(n4586), .B0(n4771), .Y(n4772));
  NOR2X1  g03215(.A(n4772), .B(n4770), .Y(n4773));
  NOR3X1  g03216(.A(n4773), .B(n4769), .C(n2681), .Y(n4774));
  NOR3X1  g03217(.A(n4574), .B(n3355), .C(n4654), .Y(n4775));
  NOR3X1  g03218(.A(n4775), .B(n4774), .C(n4764), .Y(n4776));
  NOR3X1  g03219(.A(n4773), .B(n4769), .C(n4662), .Y(n4777));
  NOR3X1  g03220(.A(n4763), .B(n4758), .C(n4665), .Y(n4778));
  AOI22X1 g03221(.A0(P1_U3086), .A1(P1_REG3_REG_13__SCAN_IN), .B0(P1_ADDR_REG_13__SCAN_IN), .B1(n4491), .Y(n4779));
  OAI21X1 g03222(.A0(n4683), .A1(n3355), .B0(n4779), .Y(n4780));
  NOR3X1  g03223(.A(n4780), .B(n4778), .C(n4777), .Y(n4781));
  OAI21X1 g03224(.A0(n4776), .A1(n4688), .B0(n4781), .Y(P1_U3256));
  XOR2X1  g03225(.A(n3310), .B(n4503), .Y(n4783));
  AOI21X1 g03226(.A0(n4753), .A1(n4760), .B0(n4756), .Y(n4784));
  AOI21X1 g03227(.A0(n4783), .A1(n4756), .B0(n4784), .Y(n4785));
  NOR2X1  g03228(.A(n4785), .B(n4576), .Y(n4786));
  XOR2X1  g03229(.A(n3310), .B(n4586), .Y(n4787));
  NOR2X1  g03230(.A(n4787), .B(n4767), .Y(n4789));
  AOI21X1 g03231(.A0(n4787), .A1(n4767), .B0(n4789), .Y(n4790));
  OAI22X1 g03232(.A0(n4654), .A1(n3310), .B0(n2681), .B1(n4790), .Y(n4791));
  OAI21X1 g03233(.A0(n4791), .A1(n4786), .B0(n4492), .Y(n4792));
  NOR2X1  g03234(.A(n4790), .B(n4662), .Y(n4793));
  NOR2X1  g03235(.A(n4785), .B(n4665), .Y(n4794));
  AOI22X1 g03236(.A0(P1_U3086), .A1(P1_REG3_REG_12__SCAN_IN), .B0(P1_ADDR_REG_12__SCAN_IN), .B1(n4491), .Y(n4795));
  OAI21X1 g03237(.A0(n4683), .A1(n3310), .B0(n4795), .Y(n4796));
  NOR3X1  g03238(.A(n4796), .B(n4794), .C(n4793), .Y(n4797));
  NAND2X1 g03239(.A(n4797), .B(n4792), .Y(P1_U3255));
  XOR2X1  g03240(.A(n3256), .B(n4500), .Y(n4799));
  NOR2X1  g03241(.A(n4799), .B(n4551), .Y(n4801));
  AOI21X1 g03242(.A0(n4799), .A1(n4551), .B0(n4801), .Y(n4802));
  NOR2X1  g03243(.A(n4802), .B(n4576), .Y(n4803));
  XOR2X1  g03244(.A(n3256), .B(n4583), .Y(n4804));
  NOR2X1  g03245(.A(n4804), .B(n4629), .Y(n4806));
  AOI21X1 g03246(.A0(n4804), .A1(n4629), .B0(n4806), .Y(n4807));
  OAI22X1 g03247(.A0(n4654), .A1(n3256), .B0(n2681), .B1(n4807), .Y(n4808));
  OAI21X1 g03248(.A0(n4808), .A1(n4803), .B0(n4492), .Y(n4809));
  AOI22X1 g03249(.A0(P1_U3086), .A1(P1_REG3_REG_11__SCAN_IN), .B0(P1_ADDR_REG_11__SCAN_IN), .B1(n4491), .Y(n4810));
  OAI21X1 g03250(.A0(n4802), .A1(n4665), .B0(n4810), .Y(n4811));
  OAI22X1 g03251(.A0(n4683), .A1(n3256), .B0(n4662), .B1(n4807), .Y(n4812));
  NOR2X1  g03252(.A(n4812), .B(n4811), .Y(n4813));
  NAND2X1 g03253(.A(n4813), .B(n4809), .Y(P1_U3254));
  AOI21X1 g03254(.A0(n4545), .A1(n4542), .B0(n4549), .Y(n4815));
  NOR2X1  g03255(.A(n4815), .B(n4513), .Y(n4816));
  OAI21X1 g03256(.A0(n3208), .A1(n4511), .B0(n4515), .Y(n4817));
  AOI21X1 g03257(.A0(n4816), .A1(n4516), .B0(n4817), .Y(n4818));
  AOI21X1 g03258(.A0(n3164), .A1(n4514), .B0(n4816), .Y(n4819));
  AOI22X1 g03259(.A0(n3165), .A1(P1_REG2_REG_9__SCAN_IN), .B0(n4511), .B1(n3209), .Y(n4820));
  OAI21X1 g03260(.A0(n3209), .A1(n4511), .B0(n4820), .Y(n4821));
  NOR2X1  g03261(.A(n4821), .B(n4819), .Y(n4822));
  NOR3X1  g03262(.A(n4822), .B(n4818), .C(n4576), .Y(n4823));
  AOI21X1 g03263(.A0(n4626), .A1(n4624), .B0(n4593), .Y(n4824));
  OAI21X1 g03264(.A0(n3208), .A1(n4591), .B0(n4595), .Y(n4825));
  AOI21X1 g03265(.A0(n4824), .A1(n4596), .B0(n4825), .Y(n4826));
  AOI21X1 g03266(.A0(n3164), .A1(n4594), .B0(n4824), .Y(n4827));
  AOI22X1 g03267(.A0(n3165), .A1(P1_REG1_REG_9__SCAN_IN), .B0(n4591), .B1(n3209), .Y(n4828));
  OAI21X1 g03268(.A0(n3209), .A1(n4591), .B0(n4828), .Y(n4829));
  NOR2X1  g03269(.A(n4829), .B(n4827), .Y(n4830));
  NOR3X1  g03270(.A(n4830), .B(n4826), .C(n2681), .Y(n4831));
  NOR3X1  g03271(.A(n4574), .B(n3208), .C(n4654), .Y(n4832));
  NOR3X1  g03272(.A(n4832), .B(n4831), .C(n4823), .Y(n4833));
  NOR3X1  g03273(.A(n4822), .B(n4818), .C(n4665), .Y(n4834));
  OAI22X1 g03274(.A0(P1_STATE_REG_SCAN_IN), .A1(n3191), .B0(n1547), .B1(n4667), .Y(n4835));
  NOR3X1  g03275(.A(n4830), .B(n4826), .C(n4662), .Y(n4836));
  NOR4X1  g03276(.A(n4491), .B(n3208), .C(n4654), .D(n2343), .Y(n4837));
  NOR4X1  g03277(.A(n4836), .B(n4835), .C(n4834), .D(n4837), .Y(n4838));
  OAI21X1 g03278(.A0(n4833), .A1(n4688), .B0(n4838), .Y(P1_U3253));
  XOR2X1  g03279(.A(n3164), .B(n4514), .Y(n4840));
  NOR2X1  g03280(.A(n4840), .B(n4816), .Y(n4842));
  AOI21X1 g03281(.A0(n4840), .A1(n4816), .B0(n4842), .Y(n4843));
  NOR2X1  g03282(.A(n4843), .B(n4576), .Y(n4844));
  XOR2X1  g03283(.A(n3164), .B(n4594), .Y(n4845));
  NOR2X1  g03284(.A(n4845), .B(n4824), .Y(n4847));
  AOI21X1 g03285(.A0(n4845), .A1(n4824), .B0(n4847), .Y(n4848));
  OAI22X1 g03286(.A0(n4654), .A1(n3164), .B0(n2681), .B1(n4848), .Y(n4849));
  OAI21X1 g03287(.A0(n4849), .A1(n4844), .B0(n4492), .Y(n4850));
  AOI22X1 g03288(.A0(P1_U3086), .A1(P1_REG3_REG_9__SCAN_IN), .B0(P1_ADDR_REG_9__SCAN_IN), .B1(n4491), .Y(n4851));
  OAI21X1 g03289(.A0(n4843), .A1(n4665), .B0(n4851), .Y(n4852));
  OAI22X1 g03290(.A0(n4683), .A1(n3164), .B0(n4662), .B1(n4848), .Y(n4853));
  NOR2X1  g03291(.A(n4853), .B(n4852), .Y(n4854));
  NAND2X1 g03292(.A(n4854), .B(n4850), .Y(P1_U3252));
  NOR3X1  g03293(.A(n4574), .B(n3117), .C(n4654), .Y(n4856));
  XOR2X1  g03294(.A(n3117), .B(P1_REG1_REG_8__SCAN_IN), .Y(n4857));
  NOR2X1  g03295(.A(n4857), .B(n4624), .Y(n4858));
  AOI21X1 g03296(.A0(n4857), .A1(n4624), .B0(n4858), .Y(n4860));
  XOR2X1  g03297(.A(n3117), .B(P1_REG2_REG_8__SCAN_IN), .Y(n4861));
  NOR2X1  g03298(.A(n4861), .B(n4546), .Y(n4862));
  AOI21X1 g03299(.A0(n4861), .A1(n4546), .B0(n4862), .Y(n4864));
  OAI22X1 g03300(.A0(n4860), .A1(n2681), .B0(n4576), .B1(n4864), .Y(n4865));
  OAI21X1 g03301(.A0(n4865), .A1(n4856), .B0(n4492), .Y(n4866));
  AOI22X1 g03302(.A0(P1_U3086), .A1(P1_REG3_REG_8__SCAN_IN), .B0(P1_ADDR_REG_8__SCAN_IN), .B1(n4491), .Y(n4867));
  OAI21X1 g03303(.A0(n4864), .A1(n4665), .B0(n4867), .Y(n4868));
  OAI22X1 g03304(.A0(n4683), .A1(n3117), .B0(n4662), .B1(n4860), .Y(n4869));
  NOR2X1  g03305(.A(n4869), .B(n4868), .Y(n4870));
  NAND2X1 g03306(.A(n4870), .B(n4866), .Y(P1_U3251));
  NOR3X1  g03307(.A(n4574), .B(n3061), .C(n4654), .Y(n4872));
  NOR2X1  g03308(.A(n3004), .B(n2994), .Y(n4873));
  INVX1   g03309(.A(n4601), .Y(n4874));
  AOI21X1 g03310(.A0(n3062), .A1(P1_REG1_REG_7__SCAN_IN), .B0(n4874), .Y(n4875));
  OAI21X1 g03311(.A0(n4873), .A1(n4619), .B0(n4875), .Y(n4876));
  AOI22X1 g03312(.A0(n4614), .A1(n4618), .B0(n3004), .B1(n2994), .Y(n4877));
  AOI21X1 g03313(.A0(n3062), .A1(n4600), .B0(n4873), .Y(n4878));
  OAI21X1 g03314(.A0(n3062), .A1(n4600), .B0(n4878), .Y(n4879));
  OAI21X1 g03315(.A0(n4879), .A1(n4877), .B0(n4876), .Y(n4880));
  NOR2X1  g03316(.A(n3004), .B(n4520), .Y(n4881));
  INVX1   g03317(.A(n4522), .Y(n4882));
  AOI21X1 g03318(.A0(n3062), .A1(P1_REG2_REG_7__SCAN_IN), .B0(n4882), .Y(n4883));
  OAI21X1 g03319(.A0(n4881), .A1(n4541), .B0(n4883), .Y(n4884));
  AOI22X1 g03320(.A0(n4536), .A1(n4540), .B0(n3004), .B1(n4520), .Y(n4885));
  AOI21X1 g03321(.A0(n3062), .A1(n4521), .B0(n4881), .Y(n4886));
  OAI21X1 g03322(.A0(n3062), .A1(n4521), .B0(n4886), .Y(n4887));
  OAI21X1 g03323(.A0(n4887), .A1(n4885), .B0(n4884), .Y(n4888));
  OAI22X1 g03324(.A0(n4880), .A1(n2681), .B0(n4576), .B1(n4888), .Y(n4889));
  OAI21X1 g03325(.A0(n4889), .A1(n4872), .B0(n4492), .Y(n4890));
  AOI22X1 g03326(.A0(P1_U3086), .A1(P1_REG3_REG_7__SCAN_IN), .B0(P1_ADDR_REG_7__SCAN_IN), .B1(n4491), .Y(n4891));
  OAI21X1 g03327(.A0(n4888), .A1(n4665), .B0(n4891), .Y(n4892));
  OAI22X1 g03328(.A0(n4683), .A1(n3061), .B0(n4662), .B1(n4880), .Y(n4893));
  NOR2X1  g03329(.A(n4893), .B(n4892), .Y(n4894));
  NAND2X1 g03330(.A(n4894), .B(n4890), .Y(P1_U3250));
  NOR3X1  g03331(.A(n4574), .B(n3004), .C(n4654), .Y(n4896));
  XOR2X1  g03332(.A(n3004), .B(P1_REG1_REG_6__SCAN_IN), .Y(n4897));
  NOR2X1  g03333(.A(n4897), .B(n4619), .Y(n4898));
  XOR2X1  g03334(.A(n3004), .B(n2994), .Y(n4899));
  AOI21X1 g03335(.A0(n4618), .A1(n4614), .B0(n4899), .Y(n4900));
  NOR2X1  g03336(.A(n4900), .B(n4898), .Y(n4901));
  XOR2X1  g03337(.A(n3004), .B(P1_REG2_REG_6__SCAN_IN), .Y(n4902));
  NOR2X1  g03338(.A(n4902), .B(n4541), .Y(n4903));
  XOR2X1  g03339(.A(n3004), .B(n4520), .Y(n4904));
  AOI21X1 g03340(.A0(n4540), .A1(n4536), .B0(n4904), .Y(n4905));
  NOR2X1  g03341(.A(n4905), .B(n4903), .Y(n4906));
  OAI22X1 g03342(.A0(n4901), .A1(n2681), .B0(n4576), .B1(n4906), .Y(n4907));
  OAI21X1 g03343(.A0(n4907), .A1(n4896), .B0(n4492), .Y(n4908));
  AOI22X1 g03344(.A0(P1_U3086), .A1(P1_REG3_REG_6__SCAN_IN), .B0(P1_ADDR_REG_6__SCAN_IN), .B1(n4491), .Y(n4909));
  OAI21X1 g03345(.A0(n4906), .A1(n4665), .B0(n4909), .Y(n4910));
  OAI22X1 g03346(.A0(n4683), .A1(n3004), .B0(n4662), .B1(n4901), .Y(n4911));
  NOR2X1  g03347(.A(n4911), .B(n4910), .Y(n4912));
  NAND2X1 g03348(.A(n4912), .B(n4908), .Y(P1_U3249));
  NOR3X1  g03349(.A(n4574), .B(n2962), .C(n4654), .Y(n4914));
  INVX1   g03350(.A(n4606), .Y(n4915));
  NOR2X1  g03351(.A(n4915), .B(n4603), .Y(n4916));
  NOR2X1  g03352(.A(n2825), .B(P1_REG1_REG_2__SCAN_IN), .Y(n4917));
  NOR3X1  g03353(.A(n4917), .B(n2754), .C(n2778), .Y(n4918));
  AOI21X1 g03354(.A0(n2825), .A1(P1_REG1_REG_2__SCAN_IN), .B0(n4918), .Y(n4919));
  NOR2X1  g03355(.A(n4919), .B(n4610), .Y(n4920));
  NOR4X1  g03356(.A(n4916), .B(n4615), .C(n4609), .D(n4920), .Y(n4921));
  OAI21X1 g03357(.A0(n2962), .A1(n2942), .B0(n4602), .Y(n4922));
  NOR3X1  g03358(.A(n4920), .B(n4916), .C(n4609), .Y(n4923));
  AOI21X1 g03359(.A0(n2917), .A1(n2894), .B0(n4923), .Y(n4924));
  INVX1   g03360(.A(n2962), .Y(n4925));
  AOI22X1 g03361(.A0(n2916), .A1(P1_REG1_REG_4__SCAN_IN), .B0(n2942), .B1(n4925), .Y(n4926));
  OAI21X1 g03362(.A0(n4925), .A1(n2942), .B0(n4926), .Y(n4927));
  OAI22X1 g03363(.A0(n4924), .A1(n4927), .B0(n4922), .B1(n4921), .Y(n4928));
  INVX1   g03364(.A(n4528), .Y(n4929));
  NOR2X1  g03365(.A(n4929), .B(n4525), .Y(n4930));
  NOR2X1  g03366(.A(n2825), .B(P1_REG2_REG_2__SCAN_IN), .Y(n4931));
  NOR3X1  g03367(.A(n4931), .B(n2754), .C(n2774), .Y(n4932));
  AOI21X1 g03368(.A0(n2825), .A1(P1_REG2_REG_2__SCAN_IN), .B0(n4932), .Y(n4933));
  NOR2X1  g03369(.A(n4933), .B(n4532), .Y(n4934));
  NOR4X1  g03370(.A(n4930), .B(n4537), .C(n4531), .D(n4934), .Y(n4935));
  OAI21X1 g03371(.A0(n2962), .A1(n4269), .B0(n4523), .Y(n4936));
  NOR3X1  g03372(.A(n4934), .B(n4930), .C(n4531), .Y(n4937));
  AOI21X1 g03373(.A0(n2917), .A1(n4261), .B0(n4937), .Y(n4938));
  AOI22X1 g03374(.A0(n2916), .A1(P1_REG2_REG_4__SCAN_IN), .B0(n4269), .B1(n4925), .Y(n4939));
  OAI21X1 g03375(.A0(n4925), .A1(n4269), .B0(n4939), .Y(n4940));
  OAI22X1 g03376(.A0(n4938), .A1(n4940), .B0(n4936), .B1(n4935), .Y(n4941));
  OAI22X1 g03377(.A0(n4928), .A1(n2681), .B0(n4576), .B1(n4941), .Y(n4942));
  OAI21X1 g03378(.A0(n4942), .A1(n4914), .B0(n4492), .Y(n4943));
  INVX1   g03379(.A(n4928), .Y(n4944));
  NAND2X1 g03380(.A(n4944), .B(n4661), .Y(n4945));
  AOI22X1 g03381(.A0(P1_U3086), .A1(P1_REG3_REG_5__SCAN_IN), .B0(P1_ADDR_REG_5__SCAN_IN), .B1(n4491), .Y(n4946));
  NOR4X1  g03382(.A(n2343), .B(n4576), .C(n4491), .D(n4941), .Y(n4947));
  AOI21X1 g03383(.A0(n4666), .A1(n4925), .B0(n4947), .Y(n4948));
  NAND4X1 g03384(.A(n4946), .B(n4945), .C(n4943), .D(n4948), .Y(P1_U3248));
  NAND3X1 g03385(.A(n2549), .B(n2543), .C(n2554), .Y(n4950));
  NOR3X1  g03386(.A(n2540), .B(n4950), .C(P1_U3086), .Y(P1_U4016));
  INVX1   g03387(.A(P1_U4016), .Y(n4952));
  NAND2X1 g03388(.A(n2658), .B(n2660), .Y(n4953));
  NOR2X1  g03389(.A(n2713), .B(n2668), .Y(n4954));
  AOI21X1 g03390(.A0(n2668), .A1(n2666), .B0(n4954), .Y(n4955));
  AOI21X1 g03391(.A0(n4955), .A1(n4953), .B0(n2538), .Y(n4956));
  NOR3X1  g03392(.A(n2673), .B(n2666), .C(n2660), .Y(n4957));
  AOI21X1 g03393(.A0(n2673), .A1(n2658), .B0(n2656), .Y(n4958));
  OAI21X1 g03394(.A0(n4958), .A1(n4957), .B0(n4950), .Y(n4959));
  NAND2X1 g03395(.A(n4954), .B(n4950), .Y(n4960));
  AOI21X1 g03396(.A0(n4960), .A1(n4959), .B0(n2710), .Y(n4961));
  NAND3X1 g03397(.A(n2668), .B(n2656), .C(n4950), .Y(n4962));
  OAI22X1 g03398(.A0(n2739), .A1(n4962), .B0(n2219), .B1(n4950), .Y(n4963));
  NOR2X1  g03399(.A(n4963), .B(n4961), .Y(n4964));
  XOR2X1  g03400(.A(n4964), .B(n4956), .Y(n4965));
  NOR2X1  g03401(.A(n2668), .B(n2654), .Y(n4966));
  NAND2X1 g03402(.A(n2673), .B(n2658), .Y(n4967));
  OAI21X1 g03403(.A0(n2658), .A1(n2656), .B0(n4967), .Y(n4968));
  OAI21X1 g03404(.A0(n4968), .A1(n4966), .B0(n4950), .Y(n4969));
  NOR2X1  g03405(.A(n4953), .B(n2538), .Y(n4970));
  NAND3X1 g03406(.A(n2713), .B(n2656), .C(n2654), .Y(n4971));
  OAI21X1 g03407(.A0(n2713), .A1(n2668), .B0(n2666), .Y(n4972));
  AOI21X1 g03408(.A0(n4972), .A1(n4971), .B0(n2538), .Y(n4973));
  NOR2X1  g03409(.A(n4967), .B(n2538), .Y(n4974));
  NOR3X1  g03410(.A(n4974), .B(n4973), .C(n4970), .Y(n4975));
  NOR3X1  g03411(.A(n2658), .B(n2666), .C(n2538), .Y(n4976));
  AOI22X1 g03412(.A0(n2768), .A1(n4976), .B0(n2538), .B1(P1_REG1_REG_0__SCAN_IN), .Y(n4977));
  OAI21X1 g03413(.A0(n4975), .A1(n2739), .B0(n4977), .Y(n4978));
  XOR2X1  g03414(.A(n4978), .B(n4969), .Y(n4979));
  XOR2X1  g03415(.A(n4979), .B(n4965), .Y(n4980));
  NOR2X1  g03416(.A(n2687), .B(n2681), .Y(n4981));
  NAND3X1 g03417(.A(n4575), .B(n2219), .C(P1_REG2_REG_0__SCAN_IN), .Y(n4982));
  AOI21X1 g03418(.A0(n2681), .A1(n2702), .B0(n2687), .Y(n4983));
  OAI21X1 g03419(.A0(n4983), .A1(n2219), .B0(n4982), .Y(n4984));
  AOI21X1 g03420(.A0(n4981), .A1(n4980), .B0(n4984), .Y(n4985));
  XOR2X1  g03421(.A(n2916), .B(P1_REG1_REG_4__SCAN_IN), .Y(n4986));
  NOR2X1  g03422(.A(n4986), .B(n4923), .Y(n4988));
  AOI21X1 g03423(.A0(n4986), .A1(n4923), .B0(n4988), .Y(n4989));
  XOR2X1  g03424(.A(n2916), .B(P1_REG2_REG_4__SCAN_IN), .Y(n4990));
  NOR2X1  g03425(.A(n4990), .B(n4937), .Y(n4992));
  AOI21X1 g03426(.A0(n4990), .A1(n4937), .B0(n4992), .Y(n4993));
  OAI22X1 g03427(.A0(n4989), .A1(n2681), .B0(n4576), .B1(n4993), .Y(n4994));
  AOI21X1 g03428(.A0(n2687), .A1(n2916), .B0(n4994), .Y(n4995));
  NOR2X1  g03429(.A(n4995), .B(n4688), .Y(n4996));
  AOI22X1 g03430(.A0(P1_U3086), .A1(P1_REG3_REG_4__SCAN_IN), .B0(P1_ADDR_REG_4__SCAN_IN), .B1(n4491), .Y(n4997));
  OAI21X1 g03431(.A0(n4989), .A1(n4662), .B0(n4997), .Y(n4998));
  OAI22X1 g03432(.A0(n4683), .A1(n2917), .B0(n4665), .B1(n4993), .Y(n4999));
  NOR3X1  g03433(.A(n4999), .B(n4998), .C(n4996), .Y(n5000));
  OAI21X1 g03434(.A0(n4985), .A1(n4952), .B0(n5000), .Y(P1_U3247));
  OAI21X1 g03435(.A0(n4915), .A1(n4917), .B0(n4919), .Y(n5002));
  XOR2X1  g03436(.A(n2864), .B(P1_REG1_REG_3__SCAN_IN), .Y(n5003));
  OAI21X1 g03437(.A0(n4609), .A1(n4610), .B0(n5002), .Y(n5004));
  OAI21X1 g03438(.A0(n5003), .A1(n5002), .B0(n5004), .Y(n5005));
  OAI21X1 g03439(.A0(n4929), .A1(n4931), .B0(n4933), .Y(n5006));
  XOR2X1  g03440(.A(n2864), .B(P1_REG2_REG_3__SCAN_IN), .Y(n5007));
  OAI21X1 g03441(.A0(n4531), .A1(n4532), .B0(n5006), .Y(n5008));
  OAI21X1 g03442(.A0(n5007), .A1(n5006), .B0(n5008), .Y(n5009));
  AOI22X1 g03443(.A0(n5005), .A1(n2686), .B0(n4575), .B1(n5009), .Y(n5010));
  OAI21X1 g03444(.A0(n4654), .A1(n2864), .B0(n5010), .Y(n5011));
  NAND2X1 g03445(.A(n5011), .B(n4492), .Y(n5012));
  NAND2X1 g03446(.A(n5005), .B(n4661), .Y(n5013));
  AOI22X1 g03447(.A0(P1_U3086), .A1(P1_REG3_REG_3__SCAN_IN), .B0(P1_ADDR_REG_3__SCAN_IN), .B1(n4491), .Y(n5014));
  AOI22X1 g03448(.A0(n4666), .A1(n4524), .B0(n4664), .B1(n5009), .Y(n5015));
  NAND4X1 g03449(.A(n5014), .B(n5013), .C(n5012), .D(n5015), .Y(P1_U3246));
  XOR2X1  g03450(.A(n2812), .B(P1_REG1_REG_2__SCAN_IN), .Y(n5017));
  NOR2X1  g03451(.A(n5017), .B(n4608), .Y(n5018));
  AOI21X1 g03452(.A0(n5017), .A1(n4608), .B0(n5018), .Y(n5020));
  XOR2X1  g03453(.A(n2812), .B(P1_REG2_REG_2__SCAN_IN), .Y(n5021));
  NOR2X1  g03454(.A(n5021), .B(n4530), .Y(n5022));
  AOI21X1 g03455(.A0(n5021), .A1(n4530), .B0(n5022), .Y(n5024));
  AOI22X1 g03456(.A0(n5020), .A1(n2686), .B0(n4575), .B1(n5024), .Y(n5025));
  OAI21X1 g03457(.A0(n4654), .A1(n2812), .B0(n5025), .Y(n5026));
  NAND2X1 g03458(.A(n5024), .B(n4664), .Y(n5027));
  AOI22X1 g03459(.A0(P1_U3086), .A1(P1_REG3_REG_2__SCAN_IN), .B0(P1_ADDR_REG_2__SCAN_IN), .B1(n4491), .Y(n5028));
  AOI22X1 g03460(.A0(n4666), .A1(n2825), .B0(n4661), .B1(n5020), .Y(n5029));
  NAND3X1 g03461(.A(n5029), .B(n5028), .C(n5027), .Y(n5030));
  AOI21X1 g03462(.A0(n5026), .A1(n4492), .B0(n5030), .Y(n5031));
  OAI21X1 g03463(.A0(n4985), .A1(n4952), .B0(n5031), .Y(P1_U3245));
  XOR2X1  g03464(.A(n2754), .B(P1_REG1_REG_1__SCAN_IN), .Y(n5033));
  XOR2X1  g03465(.A(n5033), .B(n4604), .Y(n5034));
  XOR2X1  g03466(.A(n2754), .B(P1_REG2_REG_1__SCAN_IN), .Y(n5035));
  XOR2X1  g03467(.A(n5035), .B(n4526), .Y(n5036));
  OAI22X1 g03468(.A0(n5034), .A1(n2681), .B0(n4576), .B1(n5036), .Y(n5037));
  AOI21X1 g03469(.A0(n2687), .A1(n2755), .B0(n5037), .Y(n5038));
  AOI22X1 g03470(.A0(P1_U3086), .A1(P1_REG3_REG_1__SCAN_IN), .B0(P1_ADDR_REG_1__SCAN_IN), .B1(n4491), .Y(n5039));
  OAI21X1 g03471(.A0(n5034), .A1(n4662), .B0(n5039), .Y(n5040));
  OAI22X1 g03472(.A0(n4683), .A1(n2754), .B0(n4665), .B1(n5036), .Y(n5041));
  NOR2X1  g03473(.A(n5041), .B(n5040), .Y(n5042));
  OAI21X1 g03474(.A0(n5038), .A1(n4688), .B0(n5042), .Y(P1_U3244));
  XOR2X1  g03475(.A(n2219), .B(P1_REG1_REG_0__SCAN_IN), .Y(n5044));
  XOR2X1  g03476(.A(n2219), .B(P1_REG2_REG_0__SCAN_IN), .Y(n5045));
  OAI22X1 g03477(.A0(n5044), .A1(n2681), .B0(n4576), .B1(n5045), .Y(n5046));
  AOI21X1 g03478(.A0(n2687), .A1(n2691), .B0(n5046), .Y(n5047));
  AOI22X1 g03479(.A0(P1_U3086), .A1(P1_REG3_REG_0__SCAN_IN), .B0(P1_ADDR_REG_0__SCAN_IN), .B1(n4491), .Y(n5048));
  OAI21X1 g03480(.A0(n5044), .A1(n4662), .B0(n5048), .Y(n5049));
  OAI22X1 g03481(.A0(n4683), .A1(n2219), .B0(n4665), .B1(n5045), .Y(n5050));
  NOR2X1  g03482(.A(n5050), .B(n5049), .Y(n5051));
  OAI21X1 g03483(.A0(n5047), .A1(n4688), .B0(n5051), .Y(P1_U3243));
  NAND2X1 g03484(.A(P1_U4016), .B(n2768), .Y(n5053));
  OAI21X1 g03485(.A0(P1_U4016), .A1(n1796), .B0(n5053), .Y(P1_U3560));
  OAI21X1 g03486(.A0(n2780), .A1(n2777), .B0(P1_U4016), .Y(n5055));
  OAI21X1 g03487(.A0(P1_U4016), .A1(n1808), .B0(n5055), .Y(P1_U3561));
  OAI21X1 g03488(.A0(n2798), .A1(n2795), .B0(P1_U4016), .Y(n5057));
  OAI21X1 g03489(.A0(P1_U4016), .A1(n1854), .B0(n5057), .Y(P1_U3562));
  OAI21X1 g03490(.A0(n2846), .A1(n2844), .B0(P1_U4016), .Y(n5059));
  OAI21X1 g03491(.A0(P1_U4016), .A1(n1875), .B0(n5059), .Y(P1_U3563));
  OAI21X1 g03492(.A0(n2897), .A1(n2893), .B0(P1_U4016), .Y(n5061));
  OAI21X1 g03493(.A0(P1_U4016), .A1(n1884), .B0(n5061), .Y(P1_U3564));
  OAI21X1 g03494(.A0(n2945), .A1(n2941), .B0(P1_U4016), .Y(n5063));
  OAI21X1 g03495(.A0(P1_U4016), .A1(n1904), .B0(n5063), .Y(P1_U3565));
  OAI21X1 g03496(.A0(n2997), .A1(n2993), .B0(P1_U4016), .Y(n5065));
  OAI21X1 g03497(.A0(P1_U4016), .A1(n1935), .B0(n5065), .Y(P1_U3566));
  NAND2X1 g03498(.A(P1_U4016), .B(n3049), .Y(n5067));
  OAI21X1 g03499(.A0(P1_U4016), .A1(n1963), .B0(n5067), .Y(P1_U3567));
  INVX1   g03500(.A(P1_DATAO_REG_8__SCAN_IN), .Y(n5069));
  NAND2X1 g03501(.A(P1_U4016), .B(n3103), .Y(n5070));
  OAI21X1 g03502(.A0(P1_U4016), .A1(n5069), .B0(n5070), .Y(P1_U3568));
  OAI21X1 g03503(.A0(n3152), .A1(n3150), .B0(P1_U4016), .Y(n5072));
  OAI21X1 g03504(.A0(P1_U4016), .A1(n2020), .B0(n5072), .Y(P1_U3569));
  OAI21X1 g03505(.A0(n3198), .A1(n3196), .B0(P1_U4016), .Y(n5074));
  OAI21X1 g03506(.A0(P1_U4016), .A1(n2045), .B0(n5074), .Y(P1_U3570));
  INVX1   g03507(.A(P1_DATAO_REG_11__SCAN_IN), .Y(n5076));
  OAI21X1 g03508(.A0(n3244), .A1(n3242), .B0(P1_U4016), .Y(n5077));
  OAI21X1 g03509(.A0(P1_U4016), .A1(n5076), .B0(n5077), .Y(P1_U3571));
  INVX1   g03510(.A(P1_DATAO_REG_12__SCAN_IN), .Y(n5079));
  OAI21X1 g03511(.A0(n3298), .A1(n3296), .B0(P1_U4016), .Y(n5080));
  OAI21X1 g03512(.A0(P1_U4016), .A1(n5079), .B0(n5080), .Y(P1_U3572));
  NAND2X1 g03513(.A(n4952), .B(P1_DATAO_REG_13__SCAN_IN), .Y(n5082));
  OAI21X1 g03514(.A0(n4952), .A1(n3346), .B0(n5082), .Y(P1_U3573));
  NAND2X1 g03515(.A(n4952), .B(P1_DATAO_REG_14__SCAN_IN), .Y(n5084));
  OAI21X1 g03516(.A0(n4952), .A1(n3398), .B0(n5084), .Y(P1_U3574));
  NAND2X1 g03517(.A(n4952), .B(P1_DATAO_REG_15__SCAN_IN), .Y(n5086));
  OAI21X1 g03518(.A0(n4952), .A1(n3443), .B0(n5086), .Y(P1_U3575));
  NAND2X1 g03519(.A(n4952), .B(P1_DATAO_REG_16__SCAN_IN), .Y(n5088));
  OAI21X1 g03520(.A0(n4952), .A1(n3482), .B0(n5088), .Y(P1_U3576));
  NAND2X1 g03521(.A(n4952), .B(P1_DATAO_REG_17__SCAN_IN), .Y(n5090));
  OAI21X1 g03522(.A0(n4952), .A1(n3532), .B0(n5090), .Y(P1_U3577));
  NAND2X1 g03523(.A(n4952), .B(P1_DATAO_REG_18__SCAN_IN), .Y(n5092));
  OAI21X1 g03524(.A0(n4952), .A1(n3578), .B0(n5092), .Y(P1_U3578));
  NAND2X1 g03525(.A(n4952), .B(P1_DATAO_REG_19__SCAN_IN), .Y(n5094));
  OAI21X1 g03526(.A0(n4952), .A1(n3621), .B0(n5094), .Y(P1_U3579));
  NAND2X1 g03527(.A(n4952), .B(P1_DATAO_REG_20__SCAN_IN), .Y(n5096));
  OAI21X1 g03528(.A0(n4952), .A1(n3666), .B0(n5096), .Y(P1_U3580));
  NAND2X1 g03529(.A(n4952), .B(P1_DATAO_REG_21__SCAN_IN), .Y(n5098));
  OAI21X1 g03530(.A0(n4952), .A1(n3710), .B0(n5098), .Y(P1_U3581));
  NAND2X1 g03531(.A(n4952), .B(P1_DATAO_REG_22__SCAN_IN), .Y(n5100));
  OAI21X1 g03532(.A0(n4952), .A1(n3754), .B0(n5100), .Y(P1_U3582));
  NAND2X1 g03533(.A(n4952), .B(P1_DATAO_REG_23__SCAN_IN), .Y(n5102));
  OAI21X1 g03534(.A0(n4952), .A1(n3795), .B0(n5102), .Y(P1_U3583));
  NAND2X1 g03535(.A(n4952), .B(P1_DATAO_REG_24__SCAN_IN), .Y(n5104));
  OAI21X1 g03536(.A0(n4952), .A1(n3838), .B0(n5104), .Y(P1_U3584));
  NAND2X1 g03537(.A(n4952), .B(P1_DATAO_REG_25__SCAN_IN), .Y(n5106));
  OAI21X1 g03538(.A0(n4952), .A1(n3880), .B0(n5106), .Y(P1_U3585));
  NAND2X1 g03539(.A(n4952), .B(P1_DATAO_REG_26__SCAN_IN), .Y(n5108));
  OAI21X1 g03540(.A0(n4952), .A1(n3924), .B0(n5108), .Y(P1_U3586));
  NAND2X1 g03541(.A(n4952), .B(P1_DATAO_REG_27__SCAN_IN), .Y(n5110));
  OAI21X1 g03542(.A0(n4952), .A1(n3973), .B0(n5110), .Y(P1_U3587));
  NAND2X1 g03543(.A(n4952), .B(P1_DATAO_REG_28__SCAN_IN), .Y(n5112));
  OAI21X1 g03544(.A0(n4952), .A1(n4020), .B0(n5112), .Y(P1_U3588));
  NAND2X1 g03545(.A(n4952), .B(P1_DATAO_REG_29__SCAN_IN), .Y(n5114));
  OAI21X1 g03546(.A0(n4952), .A1(n4064), .B0(n5114), .Y(P1_U3589));
  INVX1   g03547(.A(P1_DATAO_REG_30__SCAN_IN), .Y(n5116));
  NOR2X1  g03548(.A(n4098), .B(n4096), .Y(n5117));
  OAI21X1 g03549(.A0(n2707), .A1(n4093), .B0(n5117), .Y(n5118));
  NAND2X1 g03550(.A(P1_U4016), .B(n5118), .Y(n5119));
  OAI21X1 g03551(.A0(P1_U4016), .A1(n5116), .B0(n5119), .Y(P1_U3590));
  INVX1   g03552(.A(P1_DATAO_REG_31__SCAN_IN), .Y(n5121));
  NOR2X1  g03553(.A(n4132), .B(n4130), .Y(n5122));
  OAI21X1 g03554(.A0(n2707), .A1(n4127), .B0(n5122), .Y(n5123));
  NAND2X1 g03555(.A(P1_U4016), .B(n5123), .Y(n5124));
  OAI21X1 g03556(.A0(P1_U4016), .A1(n5121), .B0(n5124), .Y(P1_U3591));
  NAND3X1 g03557(.A(n2673), .B(n2666), .C(n2660), .Y(n5126));
  NAND2X1 g03558(.A(n5126), .B(n2717), .Y(n5127));
  NAND4X1 g03559(.A(n2668), .B(n2656), .C(n2654), .D(n2713), .Y(n5128));
  NOR2X1  g03560(.A(n5128), .B(n4487), .Y(n5129));
  NAND3X1 g03561(.A(n2673), .B(n2658), .C(n2654), .Y(n5130));
  NAND4X1 g03562(.A(n4227), .B(n4230), .C(n2723), .D(n5130), .Y(n5131));
  NOR3X1  g03563(.A(n5131), .B(n5129), .C(n5127), .Y(n5132));
  NAND3X1 g03564(.A(n2713), .B(n2658), .C(n2654), .Y(n5133));
  NAND3X1 g03565(.A(n2673), .B(n2658), .C(n2660), .Y(n5134));
  NAND2X1 g03566(.A(n5134), .B(n5133), .Y(n5135));
  INVX1   g03567(.A(n5135), .Y(n5136));
  NAND3X1 g03568(.A(n2713), .B(n2666), .C(n2660), .Y(n5137));
  NAND2X1 g03569(.A(n5137), .B(n3289), .Y(n5138));
  OAI21X1 g03570(.A0(n5123), .A1(n4099), .B0(n5138), .Y(n5139));
  NAND2X1 g03571(.A(n5139), .B(n5136), .Y(n5140));
  NOR3X1  g03572(.A(n2673), .B(n2656), .C(n2654), .Y(n5141));
  NOR2X1  g03573(.A(n5141), .B(n2720), .Y(n5142));
  NOR3X1  g03574(.A(n5142), .B(n5123), .C(n4099), .Y(n5143));
  XOR2X1  g03575(.A(n5123), .B(n4099), .Y(n5144));
  AOI22X1 g03576(.A0(n5143), .A1(n5144), .B0(n5140), .B1(n5123), .Y(n5145));
  OAI21X1 g03577(.A0(n5132), .A1(n4141), .B0(n5145), .Y(n5146));
  NOR2X1  g03578(.A(n5138), .B(n5135), .Y(n5147));
  NOR2X1  g03579(.A(n5131), .B(n5129), .Y(n5148));
  OAI21X1 g03580(.A0(n5123), .A1(n4099), .B0(n5127), .Y(n5149));
  NAND2X1 g03581(.A(n5149), .B(n5148), .Y(n5150));
  NOR3X1  g03582(.A(n2713), .B(n2656), .C(n2654), .Y(n5151));
  NOR2X1  g03583(.A(n5151), .B(n2751), .Y(n5152));
  NOR3X1  g03584(.A(n5152), .B(n5123), .C(n4099), .Y(n5153));
  AOI22X1 g03585(.A0(n5150), .A1(n5123), .B0(n5144), .B1(n5153), .Y(n5154));
  OAI21X1 g03586(.A0(n5147), .A1(n4141), .B0(n5154), .Y(n5155));
  XOR2X1  g03587(.A(n5155), .B(n5146), .Y(n5156));
  NAND4X1 g03588(.A(n5134), .B(n5133), .C(n3289), .D(n5137), .Y(n5157));
  NAND3X1 g03589(.A(n5157), .B(n2810), .C(n2505), .Y(n5158));
  NAND3X1 g03590(.A(n5127), .B(n4133), .C(n5118), .Y(n5159));
  NOR2X1  g03591(.A(n5159), .B(n5118), .Y(n5160));
  AOI21X1 g03592(.A0(n5150), .A1(n5118), .B0(n5160), .Y(n5161));
  NAND3X1 g03593(.A(n5138), .B(n4133), .C(n5118), .Y(n5162));
  NOR2X1  g03594(.A(n5162), .B(n5118), .Y(n5163));
  AOI21X1 g03595(.A0(n5140), .A1(n5118), .B0(n5163), .Y(n5164));
  OAI21X1 g03596(.A0(n5132), .A1(n4124), .B0(n5164), .Y(n5165));
  AOI21X1 g03597(.A0(n5161), .A1(n5158), .B0(n5165), .Y(n5166));
  OAI22X1 g03598(.A0(n5147), .A1(n2739), .B0(n2710), .B1(n5159), .Y(n5167));
  AOI21X1 g03599(.A0(n5150), .A1(n2768), .B0(n5167), .Y(n5168));
  AOI21X1 g03600(.A0(n4133), .A1(n5118), .B0(n5142), .Y(n5169));
  OAI21X1 g03601(.A0(n5169), .A1(n5135), .B0(n2768), .Y(n5170));
  NAND4X1 g03602(.A(n4133), .B(n5118), .C(n2768), .D(n5138), .Y(n5171));
  NOR3X1  g03603(.A(n2673), .B(n2658), .C(n2666), .Y(n5172));
  NAND3X1 g03604(.A(n5172), .B(n2654), .C(n2540), .Y(n5173));
  NOR3X1  g03605(.A(n2713), .B(n2658), .C(n2666), .Y(n5174));
  NOR3X1  g03606(.A(n2713), .B(n2668), .C(n2660), .Y(n5175));
  NOR3X1  g03607(.A(n5175), .B(n5174), .C(n2743), .Y(n5176));
  NAND4X1 g03608(.A(n5173), .B(n5152), .C(n2723), .D(n5176), .Y(n5177));
  AOI21X1 g03609(.A0(n5177), .A1(n2693), .B0(n4487), .Y(n5178));
  NAND3X1 g03610(.A(n5178), .B(n5171), .C(n5170), .Y(n5179));
  AOI21X1 g03611(.A0(n2668), .A1(n2656), .B0(n4487), .Y(n5180));
  NAND4X1 g03612(.A(n5142), .B(n5134), .C(n5133), .D(n5180), .Y(n5181));
  AOI21X1 g03613(.A0(n5181), .A1(n5179), .B0(n5168), .Y(n5182));
  OAI21X1 g03614(.A0(n5169), .A1(n5135), .B0(n2737), .Y(n5183));
  NAND2X1 g03615(.A(n5143), .B(n2737), .Y(n5184));
  AOI21X1 g03616(.A0(n5177), .A1(n2757), .B0(n4487), .Y(n5185));
  NAND3X1 g03617(.A(n5185), .B(n5184), .C(n5183), .Y(n5186));
  AOI22X1 g03618(.A0(n2757), .A1(n5157), .B0(n2768), .B1(n4487), .Y(n5187));
  OAI21X1 g03619(.A0(n5159), .A1(n2781), .B0(n5187), .Y(n5188));
  AOI21X1 g03620(.A0(n5150), .A1(n2737), .B0(n5188), .Y(n5189));
  OAI22X1 g03621(.A0(n5186), .A1(n5189), .B0(n5181), .B1(n5179), .Y(n5190));
  AOI21X1 g03622(.A0(n5149), .A1(n5148), .B0(n2799), .Y(n5191));
  NOR2X1  g03623(.A(n5159), .B(n2799), .Y(n5192));
  OAI22X1 g03624(.A0(n2814), .A1(n5147), .B0(n2781), .B1(n2540), .Y(n5193));
  NOR3X1  g03625(.A(n5193), .B(n5192), .C(n5191), .Y(n5194));
  OAI21X1 g03626(.A0(n5169), .A1(n5135), .B0(n2824), .Y(n5195));
  NAND2X1 g03627(.A(n5143), .B(n2824), .Y(n5196));
  AOI21X1 g03628(.A0(n5177), .A1(n2827), .B0(n4487), .Y(n5197));
  NAND3X1 g03629(.A(n5197), .B(n5196), .C(n5195), .Y(n5198));
  AOI22X1 g03630(.A0(n5194), .A1(n5198), .B0(n5189), .B1(n5186), .Y(n5199));
  OAI21X1 g03631(.A0(n5190), .A1(n5182), .B0(n5199), .Y(n5200));
  NOR2X1  g03632(.A(n5198), .B(n5194), .Y(n5201));
  AOI21X1 g03633(.A0(n5139), .A1(n5136), .B0(n2847), .Y(n5202));
  NOR2X1  g03634(.A(n5162), .B(n2847), .Y(n5203));
  OAI21X1 g03635(.A0(n5132), .A1(n2866), .B0(n2540), .Y(n5204));
  NOR3X1  g03636(.A(n5204), .B(n5203), .C(n5202), .Y(n5205));
  NAND3X1 g03637(.A(n5176), .B(n5173), .C(n2723), .Y(n5206));
  AOI21X1 g03638(.A0(n4133), .A1(n5118), .B0(n5152), .Y(n5207));
  OAI21X1 g03639(.A0(n5207), .A1(n5206), .B0(n2859), .Y(n5208));
  NAND2X1 g03640(.A(n5153), .B(n2859), .Y(n5209));
  AOI22X1 g03641(.A0(n2870), .A1(n5157), .B0(n2824), .B1(n4487), .Y(n5210));
  NAND3X1 g03642(.A(n5210), .B(n5209), .C(n5208), .Y(n5211));
  AOI21X1 g03643(.A0(n5211), .A1(n5205), .B0(n5201), .Y(n5212));
  OAI21X1 g03644(.A0(n5207), .A1(n5206), .B0(n2954), .Y(n5213));
  NAND2X1 g03645(.A(n5153), .B(n2954), .Y(n5214));
  AOI21X1 g03646(.A0(n2858), .A1(n2843), .B0(n2540), .Y(n5215));
  AOI21X1 g03647(.A0(n5157), .A1(n2920), .B0(n5215), .Y(n5216));
  NAND3X1 g03648(.A(n5216), .B(n5214), .C(n5213), .Y(n5217));
  AOI21X1 g03649(.A0(n5139), .A1(n5136), .B0(n2898), .Y(n5218));
  NOR2X1  g03650(.A(n5162), .B(n2898), .Y(n5219));
  AOI21X1 g03651(.A0(n2957), .A1(n2919), .B0(n5132), .Y(n5220));
  NOR4X1  g03652(.A(n5219), .B(n5218), .C(n4487), .D(n5220), .Y(n5221));
  OAI22X1 g03653(.A0(n5217), .A1(n5221), .B0(n5211), .B1(n5205), .Y(n5222));
  AOI21X1 g03654(.A0(n5212), .A1(n5200), .B0(n5222), .Y(n5223));
  NAND2X1 g03655(.A(n5221), .B(n5217), .Y(n5224));
  OAI21X1 g03656(.A0(n5162), .A1(n2946), .B0(n2540), .Y(n5225));
  AOI21X1 g03657(.A0(n5140), .A1(n2960), .B0(n5225), .Y(n5226));
  OAI21X1 g03658(.A0(n5132), .A1(n2969), .B0(n5226), .Y(n5227));
  NOR2X1  g03659(.A(n5207), .B(n5206), .Y(n5228));
  AOI22X1 g03660(.A0(n2960), .A1(n5153), .B0(n2954), .B1(n4487), .Y(n5229));
  OAI21X1 g03661(.A0(n5228), .A1(n2946), .B0(n5229), .Y(n5230));
  AOI21X1 g03662(.A0(n5157), .A1(n2966), .B0(n5230), .Y(n5231));
  OAI21X1 g03663(.A0(n5231), .A1(n5227), .B0(n5224), .Y(n5232));
  AOI22X1 g03664(.A0(n3017), .A1(n5153), .B0(n2960), .B1(n4487), .Y(n5233));
  OAI21X1 g03665(.A0(n5228), .A1(n2998), .B0(n5233), .Y(n5234));
  AOI21X1 g03666(.A0(n5157), .A1(n3007), .B0(n5234), .Y(n5235));
  OAI21X1 g03667(.A0(n5162), .A1(n2998), .B0(n2540), .Y(n5236));
  AOI21X1 g03668(.A0(n5140), .A1(n3017), .B0(n5236), .Y(n5237));
  OAI21X1 g03669(.A0(n5132), .A1(n3042), .B0(n5237), .Y(n5238));
  AOI22X1 g03670(.A0(n5235), .A1(n5238), .B0(n5231), .B1(n5227), .Y(n5239));
  OAI21X1 g03671(.A0(n5232), .A1(n5223), .B0(n5239), .Y(n5240));
  NOR2X1  g03672(.A(n5238), .B(n5235), .Y(n5241));
  INVX1   g03673(.A(n5140), .Y(n5242));
  AOI21X1 g03674(.A0(n5143), .A1(n3049), .B0(n4487), .Y(n5243));
  OAI21X1 g03675(.A0(n5242), .A1(n3050), .B0(n5243), .Y(n5244));
  AOI21X1 g03676(.A0(n5177), .A1(n3067), .B0(n5244), .Y(n5245));
  OAI22X1 g03677(.A0(n3050), .A1(n5159), .B0(n2998), .B1(n2540), .Y(n5246));
  AOI21X1 g03678(.A0(n5150), .A1(n3049), .B0(n5246), .Y(n5247));
  OAI21X1 g03679(.A0(n5147), .A1(n3064), .B0(n5247), .Y(n5248));
  AOI21X1 g03680(.A0(n5248), .A1(n5245), .B0(n5241), .Y(n5249));
  AOI22X1 g03681(.A0(n3103), .A1(n5153), .B0(n3049), .B1(n4487), .Y(n5250));
  OAI21X1 g03682(.A0(n5228), .A1(n3104), .B0(n5250), .Y(n5251));
  INVX1   g03683(.A(n5251), .Y(n5252));
  OAI21X1 g03684(.A0(n5147), .A1(n3143), .B0(n5252), .Y(n5253));
  AOI21X1 g03685(.A0(n5143), .A1(n3103), .B0(n4487), .Y(n5254));
  OAI21X1 g03686(.A0(n5242), .A1(n3104), .B0(n5254), .Y(n5255));
  AOI21X1 g03687(.A0(n5177), .A1(n3120), .B0(n5255), .Y(n5256));
  OAI22X1 g03688(.A0(n5253), .A1(n5256), .B0(n5248), .B1(n5245), .Y(n5257));
  AOI21X1 g03689(.A0(n5249), .A1(n5240), .B0(n5257), .Y(n5258));
  NAND2X1 g03690(.A(n5256), .B(n5253), .Y(n5259));
  OAI21X1 g03691(.A0(n5162), .A1(n3153), .B0(n2540), .Y(n5260));
  AOI21X1 g03692(.A0(n5140), .A1(n3170), .B0(n5260), .Y(n5261));
  OAI21X1 g03693(.A0(n5132), .A1(n3190), .B0(n5261), .Y(n5262));
  AOI22X1 g03694(.A0(n3170), .A1(n5153), .B0(n3103), .B1(n4487), .Y(n5263));
  OAI21X1 g03695(.A0(n5228), .A1(n3153), .B0(n5263), .Y(n5264));
  AOI21X1 g03696(.A0(n5157), .A1(n3167), .B0(n5264), .Y(n5265));
  OAI21X1 g03697(.A0(n5265), .A1(n5262), .B0(n5259), .Y(n5266));
  AOI22X1 g03698(.A0(n3213), .A1(n5153), .B0(n3170), .B1(n4487), .Y(n5267));
  OAI21X1 g03699(.A0(n5228), .A1(n3199), .B0(n5267), .Y(n5268));
  AOI21X1 g03700(.A0(n5157), .A1(n3215), .B0(n5268), .Y(n5269));
  OAI21X1 g03701(.A0(n5162), .A1(n3199), .B0(n2540), .Y(n5270));
  AOI21X1 g03702(.A0(n5140), .A1(n3213), .B0(n5270), .Y(n5271));
  OAI21X1 g03703(.A0(n5132), .A1(n3211), .B0(n5271), .Y(n5272));
  AOI22X1 g03704(.A0(n5269), .A1(n5272), .B0(n5265), .B1(n5262), .Y(n5273));
  OAI21X1 g03705(.A0(n5266), .A1(n5258), .B0(n5273), .Y(n5274));
  NOR2X1  g03706(.A(n5272), .B(n5269), .Y(n5275));
  AOI21X1 g03707(.A0(n5143), .A1(n3266), .B0(n4487), .Y(n5276));
  OAI21X1 g03708(.A0(n5242), .A1(n3245), .B0(n5276), .Y(n5277));
  AOI21X1 g03709(.A0(n5177), .A1(n3259), .B0(n5277), .Y(n5278));
  OAI22X1 g03710(.A0(n3245), .A1(n5159), .B0(n3199), .B1(n2540), .Y(n5279));
  AOI21X1 g03711(.A0(n5150), .A1(n3266), .B0(n5279), .Y(n5280));
  OAI21X1 g03712(.A0(n5147), .A1(n3268), .B0(n5280), .Y(n5281));
  AOI21X1 g03713(.A0(n5281), .A1(n5278), .B0(n5275), .Y(n5282));
  AOI22X1 g03714(.A0(n3365), .A1(n5153), .B0(n3266), .B1(n4487), .Y(n5283));
  OAI21X1 g03715(.A0(n5228), .A1(n3299), .B0(n5283), .Y(n5284));
  AOI21X1 g03716(.A0(n5157), .A1(n3313), .B0(n5284), .Y(n5285));
  INVX1   g03717(.A(n5285), .Y(n5286));
  AOI21X1 g03718(.A0(n5143), .A1(n3365), .B0(n4487), .Y(n5287));
  OAI21X1 g03719(.A0(n5242), .A1(n3299), .B0(n5287), .Y(n5288));
  AOI21X1 g03720(.A0(n5177), .A1(n3313), .B0(n5288), .Y(n5289));
  OAI22X1 g03721(.A0(n5286), .A1(n5289), .B0(n5281), .B1(n5278), .Y(n5290));
  AOI21X1 g03722(.A0(n5282), .A1(n5274), .B0(n5290), .Y(n5291));
  INVX1   g03723(.A(n5289), .Y(n5292));
  AOI21X1 g03724(.A0(n5143), .A1(n3345), .B0(n4487), .Y(n5293));
  OAI21X1 g03725(.A0(n5242), .A1(n3346), .B0(n5293), .Y(n5294));
  INVX1   g03726(.A(n5294), .Y(n5295));
  OAI21X1 g03727(.A0(n5132), .A1(n3360), .B0(n5295), .Y(n5296));
  AOI22X1 g03728(.A0(n3345), .A1(n5153), .B0(n3365), .B1(n4487), .Y(n5297));
  OAI21X1 g03729(.A0(n5228), .A1(n3346), .B0(n5297), .Y(n5298));
  AOI21X1 g03730(.A0(n5157), .A1(n3358), .B0(n5298), .Y(n5299));
  OAI22X1 g03731(.A0(n5296), .A1(n5299), .B0(n5292), .B1(n5285), .Y(n5300));
  AOI22X1 g03732(.A0(n3405), .A1(n5153), .B0(n3345), .B1(n4487), .Y(n5301));
  OAI21X1 g03733(.A0(n5228), .A1(n3398), .B0(n5301), .Y(n5302));
  AOI21X1 g03734(.A0(n5157), .A1(n3460), .B0(n5302), .Y(n5303));
  OAI21X1 g03735(.A0(n5162), .A1(n3398), .B0(n2540), .Y(n5304));
  AOI21X1 g03736(.A0(n5140), .A1(n3405), .B0(n5304), .Y(n5305));
  OAI21X1 g03737(.A0(n5132), .A1(n3410), .B0(n5305), .Y(n5306));
  AOI22X1 g03738(.A0(n5303), .A1(n5306), .B0(n5299), .B1(n5296), .Y(n5307));
  OAI21X1 g03739(.A0(n5300), .A1(n5291), .B0(n5307), .Y(n5308));
  NOR2X1  g03740(.A(n5306), .B(n5303), .Y(n5309));
  AOI21X1 g03741(.A0(n5143), .A1(n3489), .B0(n4487), .Y(n5310));
  OAI21X1 g03742(.A0(n5242), .A1(n3443), .B0(n5310), .Y(n5311));
  AOI21X1 g03743(.A0(n5177), .A1(n3452), .B0(n5311), .Y(n5312));
  AOI22X1 g03744(.A0(n3489), .A1(n5153), .B0(n3405), .B1(n4487), .Y(n5313));
  OAI21X1 g03745(.A0(n5228), .A1(n3443), .B0(n5313), .Y(n5314));
  INVX1   g03746(.A(n5314), .Y(n5315));
  OAI21X1 g03747(.A0(n5147), .A1(n3474), .B0(n5315), .Y(n5316));
  AOI21X1 g03748(.A0(n5316), .A1(n5312), .B0(n5309), .Y(n5317));
  AOI22X1 g03749(.A0(n3503), .A1(n5153), .B0(n3489), .B1(n4487), .Y(n5318));
  OAI21X1 g03750(.A0(n5228), .A1(n3482), .B0(n5318), .Y(n5319));
  AOI21X1 g03751(.A0(n5157), .A1(n3496), .B0(n5319), .Y(n5320));
  INVX1   g03752(.A(n5320), .Y(n5321));
  AOI21X1 g03753(.A0(n5143), .A1(n3503), .B0(n4487), .Y(n5322));
  OAI21X1 g03754(.A0(n5242), .A1(n3482), .B0(n5322), .Y(n5323));
  AOI21X1 g03755(.A0(n5177), .A1(n3496), .B0(n5323), .Y(n5324));
  OAI22X1 g03756(.A0(n5321), .A1(n5324), .B0(n5316), .B1(n5312), .Y(n5325));
  AOI21X1 g03757(.A0(n5317), .A1(n5308), .B0(n5325), .Y(n5326));
  NAND2X1 g03758(.A(n5324), .B(n5321), .Y(n5327));
  AOI21X1 g03759(.A0(n5143), .A1(n3541), .B0(n4487), .Y(n5328));
  OAI21X1 g03760(.A0(n5242), .A1(n3532), .B0(n5328), .Y(n5329));
  INVX1   g03761(.A(n5329), .Y(n5330));
  OAI21X1 g03762(.A0(n5132), .A1(n3546), .B0(n5330), .Y(n5331));
  AOI22X1 g03763(.A0(n3541), .A1(n5153), .B0(n3503), .B1(n4487), .Y(n5332));
  OAI21X1 g03764(.A0(n5228), .A1(n3532), .B0(n5332), .Y(n5333));
  AOI21X1 g03765(.A0(n5157), .A1(n3547), .B0(n5333), .Y(n5334));
  OAI21X1 g03766(.A0(n5334), .A1(n5331), .B0(n5327), .Y(n5335));
  AOI22X1 g03767(.A0(n3588), .A1(n5153), .B0(n3541), .B1(n4487), .Y(n5336));
  OAI21X1 g03768(.A0(n5228), .A1(n3578), .B0(n5336), .Y(n5337));
  AOI21X1 g03769(.A0(n5157), .A1(n3640), .B0(n5337), .Y(n5338));
  AOI21X1 g03770(.A0(n5143), .A1(n3588), .B0(n4487), .Y(n5339));
  OAI21X1 g03771(.A0(n5242), .A1(n3578), .B0(n5339), .Y(n5340));
  INVX1   g03772(.A(n5340), .Y(n5341));
  OAI21X1 g03773(.A0(n5132), .A1(n3593), .B0(n5341), .Y(n5342));
  AOI22X1 g03774(.A0(n5338), .A1(n5342), .B0(n5334), .B1(n5331), .Y(n5343));
  OAI21X1 g03775(.A0(n5335), .A1(n5326), .B0(n5343), .Y(n5344));
  NOR2X1  g03776(.A(n5342), .B(n5338), .Y(n5345));
  AOI21X1 g03777(.A0(n5143), .A1(n3684), .B0(n4487), .Y(n5346));
  OAI21X1 g03778(.A0(n5242), .A1(n3621), .B0(n5346), .Y(n5347));
  AOI21X1 g03779(.A0(n5177), .A1(n3627), .B0(n5347), .Y(n5348));
  AOI22X1 g03780(.A0(n3684), .A1(n5153), .B0(n3588), .B1(n4487), .Y(n5349));
  OAI21X1 g03781(.A0(n5228), .A1(n3621), .B0(n5349), .Y(n5350));
  INVX1   g03782(.A(n5350), .Y(n5351));
  OAI21X1 g03783(.A0(n5147), .A1(n3657), .B0(n5351), .Y(n5352));
  AOI21X1 g03784(.A0(n5352), .A1(n5348), .B0(n5345), .Y(n5353));
  AOI22X1 g03785(.A0(n3665), .A1(n5153), .B0(n3684), .B1(n4487), .Y(n5354));
  OAI21X1 g03786(.A0(n5228), .A1(n3666), .B0(n5354), .Y(n5355));
  INVX1   g03787(.A(n5355), .Y(n5356));
  OAI21X1 g03788(.A0(n5147), .A1(n3673), .B0(n5356), .Y(n5357));
  AOI21X1 g03789(.A0(n5143), .A1(n3665), .B0(n4487), .Y(n5358));
  OAI21X1 g03790(.A0(n5242), .A1(n3666), .B0(n5358), .Y(n5359));
  AOI21X1 g03791(.A0(n5177), .A1(n3719), .B0(n5359), .Y(n5360));
  OAI22X1 g03792(.A0(n5357), .A1(n5360), .B0(n5352), .B1(n5348), .Y(n5361));
  AOI21X1 g03793(.A0(n5353), .A1(n5344), .B0(n5361), .Y(n5362));
  NAND2X1 g03794(.A(n5360), .B(n5357), .Y(n5363));
  AOI21X1 g03795(.A0(n5143), .A1(n3709), .B0(n4487), .Y(n5364));
  OAI21X1 g03796(.A0(n5242), .A1(n3710), .B0(n5364), .Y(n5365));
  INVX1   g03797(.A(n5365), .Y(n5366));
  OAI21X1 g03798(.A0(n5132), .A1(n3745), .B0(n5366), .Y(n5367));
  AOI22X1 g03799(.A0(n3709), .A1(n5153), .B0(n3665), .B1(n4487), .Y(n5368));
  OAI21X1 g03800(.A0(n5228), .A1(n3710), .B0(n5368), .Y(n5369));
  AOI21X1 g03801(.A0(n5157), .A1(n3715), .B0(n5369), .Y(n5370));
  OAI21X1 g03802(.A0(n5370), .A1(n5367), .B0(n5363), .Y(n5371));
  AOI22X1 g03803(.A0(n3753), .A1(n5153), .B0(n3709), .B1(n4487), .Y(n5372));
  OAI21X1 g03804(.A0(n5228), .A1(n3754), .B0(n5372), .Y(n5373));
  AOI21X1 g03805(.A0(n5157), .A1(n3761), .B0(n5373), .Y(n5374));
  AOI21X1 g03806(.A0(n5143), .A1(n3753), .B0(n4487), .Y(n5375));
  OAI21X1 g03807(.A0(n5242), .A1(n3754), .B0(n5375), .Y(n5376));
  INVX1   g03808(.A(n5376), .Y(n5377));
  OAI21X1 g03809(.A0(n5132), .A1(n3788), .B0(n5377), .Y(n5378));
  AOI22X1 g03810(.A0(n5374), .A1(n5378), .B0(n5370), .B1(n5367), .Y(n5379));
  OAI21X1 g03811(.A0(n5371), .A1(n5362), .B0(n5379), .Y(n5380));
  NOR2X1  g03812(.A(n5378), .B(n5374), .Y(n5381));
  AOI21X1 g03813(.A0(n5143), .A1(n3794), .B0(n4487), .Y(n5382));
  OAI21X1 g03814(.A0(n5242), .A1(n3795), .B0(n5382), .Y(n5383));
  AOI21X1 g03815(.A0(n5177), .A1(n3804), .B0(n5383), .Y(n5384));
  AOI22X1 g03816(.A0(n3794), .A1(n5153), .B0(n3753), .B1(n4487), .Y(n5385));
  OAI21X1 g03817(.A0(n5228), .A1(n3795), .B0(n5385), .Y(n5386));
  INVX1   g03818(.A(n5386), .Y(n5387));
  OAI21X1 g03819(.A0(n5147), .A1(n3815), .B0(n5387), .Y(n5388));
  AOI21X1 g03820(.A0(n5388), .A1(n5384), .B0(n5381), .Y(n5389));
  AOI22X1 g03821(.A0(n3837), .A1(n5153), .B0(n3794), .B1(n4487), .Y(n5390));
  OAI21X1 g03822(.A0(n5228), .A1(n3838), .B0(n5390), .Y(n5391));
  INVX1   g03823(.A(n5391), .Y(n5392));
  OAI21X1 g03824(.A0(n5147), .A1(n3863), .B0(n5392), .Y(n5393));
  AOI21X1 g03825(.A0(n5143), .A1(n3837), .B0(n4487), .Y(n5394));
  OAI21X1 g03826(.A0(n5242), .A1(n3838), .B0(n5394), .Y(n5395));
  AOI21X1 g03827(.A0(n5177), .A1(n3845), .B0(n5395), .Y(n5396));
  OAI22X1 g03828(.A0(n5393), .A1(n5396), .B0(n5388), .B1(n5384), .Y(n5397));
  AOI21X1 g03829(.A0(n5389), .A1(n5380), .B0(n5397), .Y(n5398));
  AOI21X1 g03830(.A0(n5157), .A1(n3845), .B0(n5391), .Y(n5399));
  NOR3X1  g03831(.A(n5132), .B(n2684), .C(n2358), .Y(n5400));
  NOR3X1  g03832(.A(n5395), .B(n5400), .C(n5399), .Y(n5401));
  AOI21X1 g03833(.A0(n5143), .A1(n3879), .B0(n4487), .Y(n5402));
  OAI21X1 g03834(.A0(n5242), .A1(n3880), .B0(n5402), .Y(n5403));
  INVX1   g03835(.A(n5403), .Y(n5404));
  OAI21X1 g03836(.A0(n5132), .A1(n3915), .B0(n5404), .Y(n5405));
  NAND3X1 g03837(.A(n5157), .B(n2810), .C(n3914), .Y(n5406));
  OAI22X1 g03838(.A0(n3880), .A1(n5159), .B0(n3838), .B1(n2540), .Y(n5407));
  AOI21X1 g03839(.A0(n5150), .A1(n3879), .B0(n5407), .Y(n5408));
  AOI21X1 g03840(.A0(n5408), .A1(n5406), .B0(n5405), .Y(n5409));
  NOR3X1  g03841(.A(n5409), .B(n5401), .C(n5398), .Y(n5410));
  NAND3X1 g03842(.A(n5408), .B(n5406), .C(n5405), .Y(n5411));
  AOI22X1 g03843(.A0(n3923), .A1(n5153), .B0(n3879), .B1(n4487), .Y(n5412));
  OAI21X1 g03844(.A0(n5228), .A1(n3924), .B0(n5412), .Y(n5413));
  AOI21X1 g03845(.A0(n5157), .A1(n3935), .B0(n5413), .Y(n5414));
  NOR2X1  g03846(.A(n5132), .B(n3950), .Y(n5415));
  AOI21X1 g03847(.A0(n5143), .A1(n3923), .B0(n4487), .Y(n5416));
  OAI21X1 g03848(.A0(n5242), .A1(n3924), .B0(n5416), .Y(n5417));
  OAI21X1 g03849(.A0(n5417), .A1(n5415), .B0(n5414), .Y(n5418));
  NAND2X1 g03850(.A(n5418), .B(n5411), .Y(n5419));
  NOR3X1  g03851(.A(n5417), .B(n5415), .C(n5414), .Y(n5420));
  AOI21X1 g03852(.A0(n5143), .A1(n3972), .B0(n4487), .Y(n5421));
  OAI21X1 g03853(.A0(n5242), .A1(n3973), .B0(n5421), .Y(n5422));
  AOI21X1 g03854(.A0(n5177), .A1(n3988), .B0(n5422), .Y(n5423));
  AOI22X1 g03855(.A0(n3972), .A1(n5153), .B0(n3923), .B1(n4487), .Y(n5424));
  OAI21X1 g03856(.A0(n5228), .A1(n3973), .B0(n5424), .Y(n5425));
  INVX1   g03857(.A(n5425), .Y(n5426));
  OAI21X1 g03858(.A0(n5147), .A1(n4011), .B0(n5426), .Y(n5427));
  AOI21X1 g03859(.A0(n5427), .A1(n5423), .B0(n5420), .Y(n5428));
  OAI21X1 g03860(.A0(n5419), .A1(n5410), .B0(n5428), .Y(n5429));
  NOR2X1  g03861(.A(n5427), .B(n5423), .Y(n5430));
  NOR3X1  g03862(.A(n5132), .B(n2684), .C(n2451), .Y(n5431));
  NOR2X1  g03863(.A(n5242), .B(n4020), .Y(n5432));
  OAI21X1 g03864(.A0(n5162), .A1(n4020), .B0(n2540), .Y(n5433));
  NOR4X1  g03865(.A(n5432), .B(n5431), .C(n5430), .D(n5433), .Y(n5434));
  AOI22X1 g03866(.A0(n4019), .A1(n5153), .B0(n3972), .B1(n4487), .Y(n5435));
  OAI21X1 g03867(.A0(n5228), .A1(n4020), .B0(n5435), .Y(n5436));
  AOI21X1 g03868(.A0(n5157), .A1(n4032), .B0(n5436), .Y(n5437));
  NOR4X1  g03869(.A(n5433), .B(n5432), .C(n5431), .D(n5437), .Y(n5438));
  AOI21X1 g03870(.A0(n5434), .A1(n5429), .B0(n5438), .Y(n5439));
  OAI21X1 g03871(.A0(n5153), .A1(n5150), .B0(n4063), .Y(n5440));
  OAI21X1 g03872(.A0(n4020), .A1(n2540), .B0(n5440), .Y(n5441));
  INVX1   g03873(.A(n5441), .Y(n5442));
  OAI21X1 g03874(.A0(n5147), .A1(n4072), .B0(n5442), .Y(n5443));
  AOI21X1 g03875(.A0(n5143), .A1(n4063), .B0(n4487), .Y(n5444));
  OAI21X1 g03876(.A0(n5242), .A1(n4064), .B0(n5444), .Y(n5445));
  AOI21X1 g03877(.A0(n5177), .A1(n4113), .B0(n5445), .Y(n5446));
  NOR2X1  g03878(.A(n5437), .B(n5430), .Y(n5447));
  AOI22X1 g03879(.A0(n5446), .A1(n5443), .B0(n5429), .B1(n5447), .Y(n5448));
  NAND2X1 g03880(.A(n5448), .B(n5439), .Y(n5449));
  NOR3X1  g03881(.A(n5449), .B(n5166), .C(n5156), .Y(n5450));
  NOR4X1  g03882(.A(n5443), .B(n5166), .C(n5156), .D(n5446), .Y(n5451));
  NAND3X1 g03883(.A(n5165), .B(n5161), .C(n5158), .Y(n5452));
  NOR2X1  g03884(.A(n5452), .B(n5156), .Y(n5453));
  NOR2X1  g03885(.A(n5128), .B(n2540), .Y(n5454));
  NAND2X1 g03886(.A(n5454), .B(n5146), .Y(n5455));
  INVX1   g03887(.A(n5145), .Y(n5456));
  AOI21X1 g03888(.A0(n5177), .A1(n4482), .B0(n5456), .Y(n5457));
  INVX1   g03889(.A(n5454), .Y(n5458));
  NAND3X1 g03890(.A(n5458), .B(n5155), .C(n5457), .Y(n5459));
  OAI21X1 g03891(.A0(n5455), .A1(n5155), .B0(n5459), .Y(n5460));
  NOR4X1  g03892(.A(n5453), .B(n5451), .C(n5450), .D(n5460), .Y(n5461));
  NAND3X1 g03893(.A(n5461), .B(n2668), .C(n2660), .Y(n5462));
  XOR2X1  g03894(.A(n5155), .B(n5457), .Y(n5463));
  OAI21X1 g03895(.A0(n5147), .A1(n4124), .B0(n5161), .Y(n5464));
  NAND3X1 g03896(.A(n5177), .B(n2810), .C(n2505), .Y(n5465));
  NAND3X1 g03897(.A(n5164), .B(n5465), .C(n5464), .Y(n5466));
  NOR2X1  g03898(.A(n5446), .B(n5443), .Y(n5467));
  NAND3X1 g03899(.A(n5467), .B(n5466), .C(n5463), .Y(n5468));
  NAND4X1 g03900(.A(n5161), .B(n5158), .C(n5463), .D(n5165), .Y(n5469));
  NAND2X1 g03901(.A(n5157), .B(n4482), .Y(n5470));
  NAND4X1 g03902(.A(n5154), .B(n5470), .C(n5146), .D(n5454), .Y(n5471));
  NAND4X1 g03903(.A(n5471), .B(n5469), .C(n5468), .D(n5459), .Y(n5472));
  OAI21X1 g03904(.A0(n5472), .A1(n5450), .B0(n4090), .Y(n5473));
  XOR2X1  g03905(.A(n4141), .B(n5123), .Y(n5474));
  XOR2X1  g03906(.A(n4124), .B(n5118), .Y(n5475));
  XOR2X1  g03907(.A(n4032), .B(n4019), .Y(n5477));
  XOR2X1  g03908(.A(n4011), .B(n3973), .Y(n5478));
  XOR2X1  g03909(.A(n3815), .B(n3795), .Y(n5480));
  XOR2X1  g03910(.A(n3788), .B(n3754), .Y(n5481));
  XOR2X1  g03911(.A(n3546), .B(n3532), .Y(n5484));
  NAND3X1 g03912(.A(n3453), .B(n3411), .C(n3497), .Y(n5487));
  XOR2X1  g03913(.A(n2768), .B(n2693), .Y(n5490));
  NOR4X1  g03914(.A(n2871), .B(n2828), .C(n2758), .D(n5490), .Y(n5491));
  NAND3X1 g03915(.A(n5491), .B(n3071), .C(n2921), .Y(n5492));
  XOR2X1  g03916(.A(n2966), .B(n2960), .Y(n5493));
  NOR4X1  g03917(.A(n5492), .B(n3171), .C(n3018), .D(n5493), .Y(n5494));
  XOR2X1  g03918(.A(n3215), .B(n3213), .Y(n5495));
  NOR3X1  g03919(.A(n5495), .B(n3279), .C(n3123), .Y(n5496));
  NAND4X1 g03920(.A(n5496), .B(n5494), .C(n3314), .D(n3374), .Y(n5498));
  NOR4X1  g03921(.A(n5487), .B(n5484), .C(n3596), .D(n5498), .Y(n5499));
  NAND4X1 g03922(.A(n3674), .B(n3716), .C(n3628), .D(n5499), .Y(n5500));
  NOR4X1  g03923(.A(n5481), .B(n5480), .C(n3864), .D(n5500), .Y(n5501));
  NAND3X1 g03924(.A(n5501), .B(n3936), .C(n3888), .Y(n5502));
  NOR3X1  g03925(.A(n5502), .B(n5478), .C(n5477), .Y(n5503));
  NAND4X1 g03926(.A(n4073), .B(n5475), .C(n5474), .D(n5503), .Y(n5504));
  NOR3X1  g03927(.A(n5504), .B(n2673), .C(n2668), .Y(n5505));
  AOI21X1 g03928(.A0(n5504), .A1(n4954), .B0(n5505), .Y(n5506));
  NAND3X1 g03929(.A(n5506), .B(n5473), .C(n5462), .Y(n5507));
  OAI22X1 g03930(.A0(n5450), .A1(n5472), .B0(n2740), .B1(n5172), .Y(n5508));
  OAI21X1 g03931(.A0(n2668), .A1(n2660), .B0(n4227), .Y(n5509));
  NAND3X1 g03932(.A(n5509), .B(n5461), .C(n2656), .Y(n5510));
  NAND2X1 g03933(.A(n5510), .B(n5508), .Y(n5511));
  AOI21X1 g03934(.A0(n5507), .A1(n2666), .B0(n5511), .Y(n5512));
  OAI21X1 g03935(.A0(n5128), .A1(n4576), .B0(n4487), .Y(n5513));
  OAI21X1 g03936(.A0(n2660), .A1(n4487), .B0(P1_STATE_REG_SCAN_IN), .Y(n5514));
  AOI21X1 g03937(.A0(n4487), .A1(n2538), .B0(n5514), .Y(n5515));
  AOI21X1 g03938(.A0(n5515), .A1(n5513), .B0(n2541), .Y(n5516));
  NOR3X1  g03939(.A(n5128), .B(n4576), .C(n2561), .Y(n5517));
  AOI21X1 g03940(.A0(n5517), .A1(n5461), .B0(n5516), .Y(n5518));
  OAI21X1 g03941(.A0(n5512), .A1(n2343), .B0(n5518), .Y(P1_U3242));
  NAND2X1 g03942(.A(n4960), .B(n4959), .Y(n5520));
  AOI22X1 g03943(.A0(n5520), .A1(n3405), .B0(n3460), .B1(n4976), .Y(n5521));
  NAND2X1 g03944(.A(n4966), .B(n4950), .Y(n5522));
  NAND3X1 g03945(.A(n4960), .B(n4959), .C(n5522), .Y(n5523));
  AOI22X1 g03946(.A0(n4976), .A1(n3405), .B0(n3460), .B1(n5523), .Y(n5524));
  XOR2X1  g03947(.A(n5524), .B(n4956), .Y(n5525));
  NOR2X1  g03948(.A(n5525), .B(n5521), .Y(n5526));
  INVX1   g03949(.A(n5521), .Y(n5527));
  INVX1   g03950(.A(n5525), .Y(n5528));
  NOR2X1  g03951(.A(n5528), .B(n5527), .Y(n5529));
  INVX1   g03952(.A(n5529), .Y(n5530));
  AOI22X1 g03953(.A0(n4976), .A1(n3345), .B0(n3358), .B1(n5523), .Y(n5531));
  XOR2X1  g03954(.A(n5531), .B(n4956), .Y(n5532));
  INVX1   g03955(.A(n5532), .Y(n5533));
  AOI22X1 g03956(.A0(n5520), .A1(n3345), .B0(n3358), .B1(n4976), .Y(n5534));
  INVX1   g03957(.A(n5534), .Y(n5535));
  NOR2X1  g03958(.A(n5535), .B(n5533), .Y(n5536));
  AOI22X1 g03959(.A0(n5520), .A1(n3266), .B0(n3259), .B1(n4976), .Y(n5537));
  AOI22X1 g03960(.A0(n4976), .A1(n3266), .B0(n3259), .B1(n5523), .Y(n5538));
  XOR2X1  g03961(.A(n5538), .B(n4956), .Y(n5539));
  NOR2X1  g03962(.A(n5539), .B(n5537), .Y(n5540));
  INVX1   g03963(.A(n5520), .Y(n5541));
  OAI22X1 g03964(.A0(n5541), .A1(n3299), .B0(n3338), .B1(n4962), .Y(n5542));
  AOI22X1 g03965(.A0(n4976), .A1(n3365), .B0(n3313), .B1(n5523), .Y(n5543));
  XOR2X1  g03966(.A(n5543), .B(n4969), .Y(n5544));
  NOR2X1  g03967(.A(n5544), .B(n5542), .Y(n5545));
  AOI21X1 g03968(.A0(n5534), .A1(n5532), .B0(n5545), .Y(n5546));
  NAND2X1 g03969(.A(n5544), .B(n5542), .Y(n5547));
  OAI21X1 g03970(.A0(n5534), .A1(n5532), .B0(n5547), .Y(n5548));
  AOI21X1 g03971(.A0(n5546), .A1(n5540), .B0(n5548), .Y(n5549));
  AOI22X1 g03972(.A0(n5520), .A1(n3213), .B0(n3215), .B1(n4976), .Y(n5550));
  AOI22X1 g03973(.A0(n4976), .A1(n3213), .B0(n3215), .B1(n5523), .Y(n5551));
  XOR2X1  g03974(.A(n5551), .B(n4956), .Y(n5552));
  NOR2X1  g03975(.A(n5552), .B(n5550), .Y(n5553));
  NAND2X1 g03976(.A(n5552), .B(n5550), .Y(n5554));
  AOI22X1 g03977(.A0(n5520), .A1(n3170), .B0(n3167), .B1(n4976), .Y(n5555));
  INVX1   g03978(.A(n5555), .Y(n5556));
  AOI22X1 g03979(.A0(n5520), .A1(n3103), .B0(n3120), .B1(n4976), .Y(n5557));
  AOI22X1 g03980(.A0(n4976), .A1(n3103), .B0(n3120), .B1(n5523), .Y(n5558));
  XOR2X1  g03981(.A(n5558), .B(n4956), .Y(n5559));
  NOR2X1  g03982(.A(n5559), .B(n5557), .Y(n5560));
  AOI22X1 g03983(.A0(n5520), .A1(n3017), .B0(n3007), .B1(n4976), .Y(n5561));
  AOI22X1 g03984(.A0(n4976), .A1(n3017), .B0(n3007), .B1(n5523), .Y(n5562));
  XOR2X1  g03985(.A(n5562), .B(n4956), .Y(n5563));
  AOI22X1 g03986(.A0(n5520), .A1(n3049), .B0(n3067), .B1(n4976), .Y(n5564));
  AOI22X1 g03987(.A0(n4976), .A1(n3049), .B0(n3067), .B1(n5523), .Y(n5565));
  XOR2X1  g03988(.A(n5565), .B(n4956), .Y(n5566));
  AOI22X1 g03989(.A0(n5564), .A1(n5566), .B0(n5563), .B1(n5561), .Y(n5567));
  AOI22X1 g03990(.A0(n5520), .A1(n2960), .B0(n2966), .B1(n4976), .Y(n5568));
  AOI22X1 g03991(.A0(n4976), .A1(n2960), .B0(n2966), .B1(n5523), .Y(n5569));
  XOR2X1  g03992(.A(n5569), .B(n4956), .Y(n5570));
  NOR2X1  g03993(.A(n5570), .B(n5568), .Y(n5571));
  OAI22X1 g03994(.A0(n5541), .A1(n2898), .B0(n2938), .B1(n4962), .Y(n5572));
  AOI22X1 g03995(.A0(n5520), .A1(n2824), .B0(n2827), .B1(n4976), .Y(n5573));
  AOI22X1 g03996(.A0(n4976), .A1(n2824), .B0(n2827), .B1(n5523), .Y(n5574));
  XOR2X1  g03997(.A(n5574), .B(n4956), .Y(n5575));
  NAND2X1 g03998(.A(n5575), .B(n5573), .Y(n5576));
  OAI22X1 g03999(.A0(n5541), .A1(n2847), .B0(n2866), .B1(n4962), .Y(n5577));
  AOI22X1 g04000(.A0(n4976), .A1(n2859), .B0(n2870), .B1(n5523), .Y(n5578));
  XOR2X1  g04001(.A(n5578), .B(n4969), .Y(n5579));
  OAI21X1 g04002(.A0(n5579), .A1(n5577), .B0(n5576), .Y(n5580));
  AOI22X1 g04003(.A0(n5520), .A1(n2737), .B0(n2757), .B1(n4976), .Y(n5581));
  AOI22X1 g04004(.A0(n4976), .A1(n2737), .B0(n2757), .B1(n5523), .Y(n5582));
  XOR2X1  g04005(.A(n5582), .B(n4956), .Y(n5583));
  NOR2X1  g04006(.A(n5583), .B(n5581), .Y(n5584));
  NAND2X1 g04007(.A(n5583), .B(n5581), .Y(n5585));
  OAI21X1 g04008(.A0(n4963), .A1(n4961), .B0(n4956), .Y(n5586));
  NOR3X1  g04009(.A(n4963), .B(n4961), .C(n4956), .Y(n5587));
  OAI21X1 g04010(.A0(n5587), .A1(n4979), .B0(n5586), .Y(n5588));
  AOI21X1 g04011(.A0(n5588), .A1(n5585), .B0(n5584), .Y(n5589));
  AOI22X1 g04012(.A0(n5520), .A1(n2859), .B0(n2870), .B1(n4976), .Y(n5590));
  NOR3X1  g04013(.A(n5590), .B(n5575), .C(n5573), .Y(n5591));
  OAI21X1 g04014(.A0(n5575), .A1(n5573), .B0(n5590), .Y(n5592));
  AOI21X1 g04015(.A0(n5592), .A1(n5579), .B0(n5591), .Y(n5593));
  OAI21X1 g04016(.A0(n5589), .A1(n5580), .B0(n5593), .Y(n5594));
  NAND2X1 g04017(.A(n5594), .B(n5572), .Y(n5595));
  AOI22X1 g04018(.A0(n4976), .A1(n2954), .B0(n2920), .B1(n5523), .Y(n5596));
  XOR2X1  g04019(.A(n5596), .B(n4969), .Y(n5597));
  OAI21X1 g04020(.A0(n5594), .A1(n5572), .B0(n5597), .Y(n5598));
  AOI22X1 g04021(.A0(n5595), .A1(n5598), .B0(n5570), .B1(n5568), .Y(n5599));
  OAI21X1 g04022(.A0(n5599), .A1(n5571), .B0(n5567), .Y(n5600));
  INVX1   g04023(.A(n5566), .Y(n5601));
  NOR3X1  g04024(.A(n5564), .B(n5563), .C(n5561), .Y(n5602));
  OAI21X1 g04025(.A0(n5563), .A1(n5561), .B0(n5564), .Y(n5603));
  AOI21X1 g04026(.A0(n5603), .A1(n5601), .B0(n5602), .Y(n5604));
  AOI22X1 g04027(.A0(n5600), .A1(n5604), .B0(n5559), .B1(n5557), .Y(n5605));
  OAI21X1 g04028(.A0(n5605), .A1(n5560), .B0(n5556), .Y(n5606));
  AOI22X1 g04029(.A0(n4976), .A1(n3170), .B0(n3167), .B1(n5523), .Y(n5607));
  XOR2X1  g04030(.A(n5607), .B(n4956), .Y(n5608));
  NOR3X1  g04031(.A(n5605), .B(n5560), .C(n5556), .Y(n5609));
  OAI21X1 g04032(.A0(n5609), .A1(n5608), .B0(n5606), .Y(n5610));
  AOI21X1 g04033(.A0(n5610), .A1(n5554), .B0(n5553), .Y(n5611));
  NAND2X1 g04034(.A(n5539), .B(n5537), .Y(n5612));
  NAND2X1 g04035(.A(n5612), .B(n5546), .Y(n5613));
  OAI22X1 g04036(.A0(n5611), .A1(n5613), .B0(n5549), .B1(n5536), .Y(n5614));
  AOI21X1 g04037(.A0(n5614), .A1(n5530), .B0(n5526), .Y(n5615));
  AOI22X1 g04038(.A0(n4976), .A1(n3489), .B0(n3452), .B1(n5523), .Y(n5616));
  XOR2X1  g04039(.A(n5616), .B(n4956), .Y(n5617));
  AOI22X1 g04040(.A0(n5520), .A1(n3489), .B0(n3452), .B1(n4976), .Y(n5618));
  XOR2X1  g04041(.A(n5618), .B(n5617), .Y(n5619));
  XOR2X1  g04042(.A(n5619), .B(n5615), .Y(n5620));
  NOR3X1  g04043(.A(n2678), .B(n2650), .C(n2648), .Y(n5621));
  AOI22X1 g04044(.A0(n2751), .A1(n2658), .B0(n2660), .B1(n5174), .Y(n5622));
  NOR3X1  g04045(.A(n2658), .B(n2656), .C(n2654), .Y(n5623));
  NOR4X1  g04046(.A(n5175), .B(n4255), .C(n2725), .D(n5623), .Y(n5624));
  NAND3X1 g04047(.A(n5624), .B(n5622), .C(n2723), .Y(n5625));
  NAND3X1 g04048(.A(n5625), .B(n5621), .C(n2560), .Y(n5626));
  INVX1   g04049(.A(n5621), .Y(n5627));
  AOI21X1 g04050(.A0(n5625), .A1(n5627), .B0(n4216), .Y(n5628));
  NOR2X1  g04051(.A(n5628), .B(n2561), .Y(n5629));
  NOR3X1  g04052(.A(n5629), .B(P1_U4016), .C(n4659), .Y(n5630));
  INVX1   g04053(.A(n5630), .Y(n5631));
  NOR4X1  g04054(.A(n2540), .B(n2538), .C(P1_U3086), .D(n4225), .Y(n5632));
  AOI21X1 g04055(.A0(n5632), .A1(n5627), .B0(n5631), .Y(n5633));
  INVX1   g04056(.A(n5633), .Y(n5634));
  NOR4X1  g04057(.A(n2540), .B(n2538), .C(P1_U3086), .D(n5128), .Y(n5635));
  INVX1   g04058(.A(n5635), .Y(n5636));
  NOR4X1  g04059(.A(n2678), .B(n2650), .C(n2648), .D(n2687), .Y(n5637));
  NOR4X1  g04060(.A(n2678), .B(n2650), .C(n2648), .D(n4654), .Y(n5638));
  INVX1   g04061(.A(n5638), .Y(n5639));
  OAI22X1 g04062(.A0(n5621), .A1(n3438), .B0(n3482), .B1(n5639), .Y(n5640));
  AOI21X1 g04063(.A0(n5637), .A1(n3405), .B0(n5640), .Y(n5641));
  AOI22X1 g04064(.A0(n5621), .A1(n5632), .B0(n4213), .B1(n2560), .Y(n5642));
  INVX1   g04065(.A(n5642), .Y(n5643));
  AOI22X1 g04066(.A0(n3452), .A1(n5643), .B0(P1_U3086), .B1(P1_REG3_REG_15__SCAN_IN), .Y(n5644));
  OAI21X1 g04067(.A0(n5641), .A1(n5636), .B0(n5644), .Y(n5645));
  AOI21X1 g04068(.A0(n5634), .A1(n3439), .B0(n5645), .Y(n5646));
  OAI21X1 g04069(.A0(n5626), .A1(n5620), .B0(n5646), .Y(P1_U3241));
  AOI22X1 g04070(.A0(n5520), .A1(n3837), .B0(n3845), .B1(n4976), .Y(n5648));
  INVX1   g04071(.A(n5648), .Y(n5649));
  OAI22X1 g04072(.A0(n4962), .A1(n3838), .B0(n3863), .B1(n4975), .Y(n5650));
  XOR2X1  g04073(.A(n5650), .B(n4956), .Y(n5651));
  NAND2X1 g04074(.A(n5651), .B(n5649), .Y(n5652));
  INVX1   g04075(.A(n5652), .Y(n5653));
  NOR2X1  g04076(.A(n5651), .B(n5649), .Y(n5654));
  INVX1   g04077(.A(n5654), .Y(n5655));
  AOI22X1 g04078(.A0(n5520), .A1(n3794), .B0(n3804), .B1(n4976), .Y(n5656));
  INVX1   g04079(.A(n5656), .Y(n5657));
  AOI22X1 g04080(.A0(n4976), .A1(n3794), .B0(n3804), .B1(n5523), .Y(n5658));
  XOR2X1  g04081(.A(n5658), .B(n4956), .Y(n5659));
  INVX1   g04082(.A(n5659), .Y(n5660));
  NAND2X1 g04083(.A(n5660), .B(n5657), .Y(n5661));
  NOR2X1  g04084(.A(n5660), .B(n5657), .Y(n5662));
  AOI22X1 g04085(.A0(n5520), .A1(n3753), .B0(n3761), .B1(n4976), .Y(n5663));
  AOI22X1 g04086(.A0(n4976), .A1(n3753), .B0(n3761), .B1(n5523), .Y(n5664));
  XOR2X1  g04087(.A(n5664), .B(n4956), .Y(n5665));
  NOR2X1  g04088(.A(n5665), .B(n5663), .Y(n5666));
  NAND2X1 g04089(.A(n5665), .B(n5663), .Y(n5667));
  AOI22X1 g04090(.A0(n4976), .A1(n3709), .B0(n3715), .B1(n5523), .Y(n5668));
  XOR2X1  g04091(.A(n5668), .B(n4969), .Y(n5669));
  AOI22X1 g04092(.A0(n5520), .A1(n3709), .B0(n3715), .B1(n4976), .Y(n5670));
  INVX1   g04093(.A(n5670), .Y(n5671));
  OAI22X1 g04094(.A0(n4962), .A1(n3666), .B0(n3673), .B1(n4975), .Y(n5672));
  XOR2X1  g04095(.A(n5672), .B(n4969), .Y(n5673));
  AOI22X1 g04096(.A0(n5520), .A1(n3665), .B0(n3719), .B1(n4976), .Y(n5674));
  NAND2X1 g04097(.A(n5674), .B(n5673), .Y(n5675));
  OAI21X1 g04098(.A0(n5671), .A1(n5669), .B0(n5675), .Y(n5676));
  AOI22X1 g04099(.A0(n4976), .A1(n3684), .B0(n3627), .B1(n5523), .Y(n5677));
  XOR2X1  g04100(.A(n5677), .B(n4956), .Y(n5678));
  AOI22X1 g04101(.A0(n5520), .A1(n3684), .B0(n3627), .B1(n4976), .Y(n5679));
  NAND2X1 g04102(.A(n5679), .B(n5678), .Y(n5680));
  AOI22X1 g04103(.A0(n5520), .A1(n3588), .B0(n3640), .B1(n4976), .Y(n5681));
  OAI22X1 g04104(.A0(n4962), .A1(n3578), .B0(n3593), .B1(n4975), .Y(n5682));
  XOR2X1  g04105(.A(n5682), .B(n4969), .Y(n5683));
  NOR2X1  g04106(.A(n5683), .B(n5681), .Y(n5684));
  INVX1   g04107(.A(n5684), .Y(n5685));
  NAND2X1 g04108(.A(n5683), .B(n5681), .Y(n5686));
  INVX1   g04109(.A(n5686), .Y(n5687));
  AOI22X1 g04110(.A0(n5520), .A1(n3503), .B0(n3496), .B1(n4976), .Y(n5688));
  INVX1   g04111(.A(n5688), .Y(n5689));
  AOI22X1 g04112(.A0(n4976), .A1(n3503), .B0(n3496), .B1(n5523), .Y(n5690));
  XOR2X1  g04113(.A(n5690), .B(n4956), .Y(n5691));
  INVX1   g04114(.A(n5691), .Y(n5692));
  NOR2X1  g04115(.A(n5692), .B(n5689), .Y(n5693));
  AOI22X1 g04116(.A0(n5520), .A1(n3541), .B0(n3547), .B1(n4976), .Y(n5694));
  OAI22X1 g04117(.A0(n4962), .A1(n3532), .B0(n3546), .B1(n4975), .Y(n5695));
  XOR2X1  g04118(.A(n5695), .B(n4969), .Y(n5696));
  AOI21X1 g04119(.A0(n5696), .A1(n5694), .B0(n5693), .Y(n5697));
  NOR2X1  g04120(.A(n5618), .B(n5617), .Y(n5698));
  INVX1   g04121(.A(n5698), .Y(n5699));
  NAND2X1 g04122(.A(n5618), .B(n5617), .Y(n5700));
  INVX1   g04123(.A(n5700), .Y(n5701));
  OAI21X1 g04124(.A0(n5701), .A1(n5615), .B0(n5699), .Y(n5702));
  INVX1   g04125(.A(n5694), .Y(n5703));
  NOR2X1  g04126(.A(n5691), .B(n5688), .Y(n5704));
  INVX1   g04127(.A(n5704), .Y(n5705));
  AOI21X1 g04128(.A0(n5705), .A1(n5694), .B0(n5696), .Y(n5706));
  AOI21X1 g04129(.A0(n5704), .A1(n5703), .B0(n5706), .Y(n5707));
  INVX1   g04130(.A(n5707), .Y(n5708));
  AOI21X1 g04131(.A0(n5702), .A1(n5697), .B0(n5708), .Y(n5709));
  OAI21X1 g04132(.A0(n5709), .A1(n5687), .B0(n5685), .Y(n5710));
  NAND2X1 g04133(.A(n5710), .B(n5680), .Y(n5711));
  NOR2X1  g04134(.A(n5671), .B(n5669), .Y(n5712));
  INVX1   g04135(.A(n5712), .Y(n5713));
  NOR2X1  g04136(.A(n5674), .B(n5673), .Y(n5714));
  INVX1   g04137(.A(n5714), .Y(n5715));
  NOR2X1  g04138(.A(n5679), .B(n5678), .Y(n5716));
  INVX1   g04139(.A(n5716), .Y(n5717));
  OAI21X1 g04140(.A0(n5717), .A1(n5676), .B0(n5715), .Y(n5718));
  INVX1   g04141(.A(n5669), .Y(n5719));
  NOR2X1  g04142(.A(n5670), .B(n5719), .Y(n5720));
  AOI21X1 g04143(.A0(n5718), .A1(n5713), .B0(n5720), .Y(n5721));
  OAI21X1 g04144(.A0(n5711), .A1(n5676), .B0(n5721), .Y(n5722));
  AOI21X1 g04145(.A0(n5722), .A1(n5667), .B0(n5666), .Y(n5723));
  OAI21X1 g04146(.A0(n5723), .A1(n5662), .B0(n5661), .Y(n5724));
  AOI21X1 g04147(.A0(n5724), .A1(n5655), .B0(n5653), .Y(n5725));
  AOI22X1 g04148(.A0(n5520), .A1(n3879), .B0(n3887), .B1(n4976), .Y(n5726));
  INVX1   g04149(.A(n5726), .Y(n5727));
  AOI22X1 g04150(.A0(n4976), .A1(n3879), .B0(n3887), .B1(n5523), .Y(n5728));
  XOR2X1  g04151(.A(n5728), .B(n4956), .Y(n5729));
  INVX1   g04152(.A(n5729), .Y(n5730));
  NAND2X1 g04153(.A(n5730), .B(n5727), .Y(n5731));
  OAI22X1 g04154(.A0(n5541), .A1(n3924), .B0(n3950), .B1(n4962), .Y(n5732));
  AOI22X1 g04155(.A0(n4976), .A1(n3923), .B0(n3935), .B1(n5523), .Y(n5733));
  XOR2X1  g04156(.A(n5733), .B(n4956), .Y(n5734));
  INVX1   g04157(.A(n5734), .Y(n5735));
  OAI22X1 g04158(.A0(n5732), .A1(n5735), .B0(n5730), .B1(n5727), .Y(n5736));
  INVX1   g04159(.A(n5736), .Y(n5737));
  INVX1   g04160(.A(n5732), .Y(n5738));
  NOR2X1  g04161(.A(n5734), .B(n5738), .Y(n5739));
  INVX1   g04162(.A(n5739), .Y(n5740));
  NAND2X1 g04163(.A(n5740), .B(n5737), .Y(n5741));
  AOI21X1 g04164(.A0(n5731), .A1(n5725), .B0(n5741), .Y(n5742));
  INVX1   g04165(.A(n5626), .Y(n5743));
  AOI21X1 g04166(.A0(n5729), .A1(n5726), .B0(n5725), .Y(n5744));
  AOI22X1 g04167(.A0(n5738), .A1(n5735), .B0(n5730), .B1(n5727), .Y(n5745));
  OAI21X1 g04168(.A0(n5735), .A1(n5738), .B0(n5745), .Y(n5746));
  OAI21X1 g04169(.A0(n5746), .A1(n5744), .B0(n5743), .Y(n5747));
  NOR2X1  g04170(.A(n5639), .B(n3973), .Y(n5750));
  INVX1   g04171(.A(n5637), .Y(n5751));
  OAI22X1 g04172(.A0(n5621), .A1(n3919), .B0(n3880), .B1(n5751), .Y(n5752));
  OAI21X1 g04173(.A0(n5752), .A1(n5750), .B0(n5635), .Y(n5753));
  AOI22X1 g04174(.A0(n4437), .A1(n5634), .B0(P1_U3086), .B1(P1_REG3_REG_26__SCAN_IN), .Y(n5754));
  NAND2X1 g04175(.A(n5754), .B(n5753), .Y(n5755));
  AOI21X1 g04176(.A0(n5643), .A1(n3935), .B0(n5755), .Y(n5756));
  OAI21X1 g04177(.A0(n5747), .A1(n5742), .B0(n5756), .Y(P1_U3240));
  NOR2X1  g04178(.A(n5599), .B(n5571), .Y(n5758));
  XOR2X1  g04179(.A(n5563), .B(n5561), .Y(n5759));
  NOR2X1  g04180(.A(n5759), .B(n5758), .Y(n5761));
  AOI21X1 g04181(.A0(n5759), .A1(n5758), .B0(n5761), .Y(n5762));
  OAI22X1 g04182(.A0(n5621), .A1(n2996), .B0(n2946), .B1(n5751), .Y(n5763));
  AOI21X1 g04183(.A0(n5638), .A1(n3049), .B0(n5763), .Y(n5764));
  AOI22X1 g04184(.A0(n3007), .A1(n5643), .B0(P1_U3086), .B1(P1_REG3_REG_6__SCAN_IN), .Y(n5765));
  OAI21X1 g04185(.A0(n5764), .A1(n5636), .B0(n5765), .Y(n5766));
  AOI21X1 g04186(.A0(n5634), .A1(n4277), .B0(n5766), .Y(n5767));
  OAI21X1 g04187(.A0(n5762), .A1(n5626), .B0(n5767), .Y(P1_U3239));
  XOR2X1  g04188(.A(n5683), .B(n5681), .Y(n5769));
  XOR2X1  g04189(.A(n5769), .B(n5709), .Y(n5770));
  AOI22X1 g04190(.A0(n5627), .A1(n3574), .B0(n3684), .B1(n5638), .Y(n5771));
  OAI21X1 g04191(.A0(n5751), .A1(n3532), .B0(n5771), .Y(n5772));
  AOI22X1 g04192(.A0(n5635), .A1(n5772), .B0(P1_U3086), .B1(P1_REG3_REG_18__SCAN_IN), .Y(n5773));
  OAI21X1 g04193(.A0(n5633), .A1(n3573), .B0(n5773), .Y(n5774));
  AOI21X1 g04194(.A0(n5643), .A1(n3640), .B0(n5774), .Y(n5775));
  OAI21X1 g04195(.A0(n5770), .A1(n5626), .B0(n5775), .Y(P1_U3238));
  XOR2X1  g04196(.A(n5575), .B(n5573), .Y(n5777));
  NAND2X1 g04197(.A(n5777), .B(n5589), .Y(n5778));
  OAI21X1 g04198(.A0(n5777), .A1(n5589), .B0(n5778), .Y(n5780));
  NAND2X1 g04199(.A(n5780), .B(n5743), .Y(n5781));
  OAI22X1 g04200(.A0(n5621), .A1(n2797), .B0(n2781), .B1(n5751), .Y(n5782));
  AOI21X1 g04201(.A0(n5638), .A1(n2859), .B0(n5782), .Y(n5783));
  AOI22X1 g04202(.A0(n2827), .A1(n5643), .B0(P1_U3086), .B1(P1_REG3_REG_2__SCAN_IN), .Y(n5784));
  OAI21X1 g04203(.A0(n5783), .A1(n5636), .B0(n5784), .Y(n5785));
  AOI21X1 g04204(.A0(n5634), .A1(P1_REG3_REG_2__SCAN_IN), .B0(n5785), .Y(n5786));
  NAND2X1 g04205(.A(n5786), .B(n5781), .Y(P1_U3237));
  XOR2X1  g04206(.A(n5539), .B(n5537), .Y(n5788));
  NAND2X1 g04207(.A(n5788), .B(n5611), .Y(n5789));
  OAI21X1 g04208(.A0(n5788), .A1(n5611), .B0(n5789), .Y(n5791));
  NAND2X1 g04209(.A(n5791), .B(n5743), .Y(n5792));
  OAI22X1 g04210(.A0(n5621), .A1(n3239), .B0(n3199), .B1(n5751), .Y(n5793));
  AOI21X1 g04211(.A0(n5638), .A1(n3365), .B0(n5793), .Y(n5794));
  AOI22X1 g04212(.A0(n3259), .A1(n5643), .B0(P1_U3086), .B1(P1_REG3_REG_11__SCAN_IN), .Y(n5795));
  OAI21X1 g04213(.A0(n5794), .A1(n5636), .B0(n5795), .Y(n5796));
  AOI21X1 g04214(.A0(n5634), .A1(n3240), .B0(n5796), .Y(n5797));
  NAND2X1 g04215(.A(n5797), .B(n5792), .Y(P1_U3236));
  INVX1   g04216(.A(n5663), .Y(n5799));
  XOR2X1  g04217(.A(n5665), .B(n5799), .Y(n5800));
  XOR2X1  g04218(.A(n5800), .B(n5722), .Y(n5801));
  AOI22X1 g04219(.A0(n5627), .A1(n3748), .B0(n3709), .B1(n5637), .Y(n5802));
  OAI21X1 g04220(.A0(n5639), .A1(n3795), .B0(n5802), .Y(n5803));
  AOI22X1 g04221(.A0(n5635), .A1(n5803), .B0(P1_U3086), .B1(P1_REG3_REG_22__SCAN_IN), .Y(n5804));
  OAI21X1 g04222(.A0(n5633), .A1(n3749), .B0(n5804), .Y(n5805));
  AOI21X1 g04223(.A0(n5643), .A1(n3761), .B0(n5805), .Y(n5806));
  OAI21X1 g04224(.A0(n5801), .A1(n5626), .B0(n5806), .Y(P1_U3235));
  AOI21X1 g04225(.A0(n5539), .A1(n5537), .B0(n5611), .Y(n5808));
  NOR2X1  g04226(.A(n5808), .B(n5540), .Y(n5809));
  OAI21X1 g04227(.A0(n5534), .A1(n5532), .B0(n5546), .Y(n5810));
  AOI21X1 g04228(.A0(n5809), .A1(n5547), .B0(n5810), .Y(n5811));
  OAI21X1 g04229(.A0(n5535), .A1(n5532), .B0(n5547), .Y(n5812));
  AOI21X1 g04230(.A0(n5535), .A1(n5532), .B0(n5812), .Y(n5813));
  OAI21X1 g04231(.A0(n5809), .A1(n5545), .B0(n5813), .Y(n5814));
  NAND2X1 g04232(.A(n5814), .B(n5743), .Y(n5815));
  OAI22X1 g04233(.A0(n5621), .A1(n3341), .B0(n3398), .B1(n5639), .Y(n5816));
  AOI21X1 g04234(.A0(n5637), .A1(n3365), .B0(n5816), .Y(n5817));
  AOI22X1 g04235(.A0(n3358), .A1(n5643), .B0(P1_U3086), .B1(P1_REG3_REG_13__SCAN_IN), .Y(n5818));
  OAI21X1 g04236(.A0(n5817), .A1(n5636), .B0(n5818), .Y(n5819));
  AOI21X1 g04237(.A0(n5634), .A1(n3342), .B0(n5819), .Y(n5820));
  OAI21X1 g04238(.A0(n5815), .A1(n5811), .B0(n5820), .Y(P1_U3234));
  INVX1   g04239(.A(n5674), .Y(n5822));
  XOR2X1  g04240(.A(n5822), .B(n5673), .Y(n5823));
  AOI21X1 g04241(.A0(n5710), .A1(n5680), .B0(n5716), .Y(n5824));
  INVX1   g04242(.A(n5824), .Y(n5825));
  NOR2X1  g04243(.A(n5825), .B(n5823), .Y(n5826));
  AOI21X1 g04244(.A0(n5715), .A1(n5675), .B0(n5824), .Y(n5827));
  OAI21X1 g04245(.A0(n5827), .A1(n5826), .B0(n5743), .Y(n5828));
  NAND2X1 g04246(.A(n5643), .B(n3719), .Y(n5829));
  OAI22X1 g04247(.A0(n5621), .A1(n3661), .B0(n3710), .B1(n5639), .Y(n5830));
  AOI21X1 g04248(.A0(n5637), .A1(n3684), .B0(n5830), .Y(n5831));
  OAI22X1 g04249(.A0(n5636), .A1(n5831), .B0(P1_STATE_REG_SCAN_IN), .B1(n3658), .Y(n5832));
  AOI21X1 g04250(.A0(n5634), .A1(n4384), .B0(n5832), .Y(n5833));
  NAND3X1 g04251(.A(n5833), .B(n5829), .C(n5828), .Y(P1_U3233));
  OAI21X1 g04252(.A0(n4225), .A1(n2561), .B0(n5636), .Y(n5835));
  AOI21X1 g04253(.A0(n5835), .A1(n5627), .B0(n5631), .Y(n5836));
  NOR2X1  g04254(.A(n5636), .B(n2781), .Y(n5837));
  AOI22X1 g04255(.A0(n5638), .A1(n5837), .B0(P1_U3086), .B1(P1_REG3_REG_0__SCAN_IN), .Y(n5838));
  OAI21X1 g04256(.A0(n5642), .A1(n2739), .B0(n5838), .Y(n5839));
  AOI21X1 g04257(.A0(n5743), .A1(n4980), .B0(n5839), .Y(n5840));
  OAI21X1 g04258(.A0(n5836), .A1(n2706), .B0(n5840), .Y(P1_U3232));
  NOR2X1  g04259(.A(n5605), .B(n5560), .Y(n5842));
  XOR2X1  g04260(.A(n5608), .B(n5555), .Y(n5843));
  XOR2X1  g04261(.A(n5843), .B(n5842), .Y(n5844));
  OAI22X1 g04262(.A0(n5621), .A1(n3147), .B0(n3104), .B1(n5751), .Y(n5845));
  AOI21X1 g04263(.A0(n5638), .A1(n3213), .B0(n5845), .Y(n5846));
  AOI22X1 g04264(.A0(n3167), .A1(n5643), .B0(P1_U3086), .B1(P1_REG3_REG_9__SCAN_IN), .Y(n5847));
  OAI21X1 g04265(.A0(n5846), .A1(n5636), .B0(n5847), .Y(n5848));
  AOI21X1 g04266(.A0(n5634), .A1(n3148), .B0(n5848), .Y(n5849));
  OAI21X1 g04267(.A0(n5844), .A1(n5626), .B0(n5849), .Y(P1_U3231));
  XOR2X1  g04268(.A(n5597), .B(n5572), .Y(n5851));
  XOR2X1  g04269(.A(n5851), .B(n5594), .Y(n5852));
  NAND2X1 g04270(.A(n5852), .B(n5743), .Y(n5853));
  NOR2X1  g04271(.A(n5633), .B(n2896), .Y(n5854));
  OAI22X1 g04272(.A0(n5621), .A1(n2896), .B0(n2847), .B1(n5751), .Y(n5855));
  AOI21X1 g04273(.A0(n5638), .A1(n2960), .B0(n5855), .Y(n5856));
  AOI22X1 g04274(.A0(n2920), .A1(n5643), .B0(P1_U3086), .B1(P1_REG3_REG_4__SCAN_IN), .Y(n5857));
  OAI21X1 g04275(.A0(n5856), .A1(n5636), .B0(n5857), .Y(n5858));
  NOR2X1  g04276(.A(n5858), .B(n5854), .Y(n5859));
  NAND2X1 g04277(.A(n5859), .B(n5853), .Y(P1_U3230));
  XOR2X1  g04278(.A(n5651), .B(n5648), .Y(n5861));
  OAI21X1 g04279(.A0(n5654), .A1(n5653), .B0(n5724), .Y(n5862));
  OAI21X1 g04280(.A0(n5861), .A1(n5724), .B0(n5862), .Y(n5863));
  NAND2X1 g04281(.A(n5863), .B(n5743), .Y(n5864));
  NAND2X1 g04282(.A(n5643), .B(n3845), .Y(n5865));
  NOR2X1  g04283(.A(n5639), .B(n3880), .Y(n5866));
  OAI22X1 g04284(.A0(n5621), .A1(n3833), .B0(n3795), .B1(n5751), .Y(n5867));
  OAI21X1 g04285(.A0(n5867), .A1(n5866), .B0(n5635), .Y(n5868));
  AOI22X1 g04286(.A0(n4418), .A1(n5634), .B0(P1_U3086), .B1(P1_REG3_REG_24__SCAN_IN), .Y(n5869));
  NAND4X1 g04287(.A(n5868), .B(n5865), .C(n5864), .D(n5869), .Y(P1_U3229));
  NOR2X1  g04288(.A(n5704), .B(n5702), .Y(n5871));
  OAI21X1 g04289(.A0(n5696), .A1(n5694), .B0(n5697), .Y(n5872));
  OAI21X1 g04290(.A0(n5692), .A1(n5689), .B0(n5702), .Y(n5873));
  OAI21X1 g04291(.A0(n5696), .A1(n5703), .B0(n5705), .Y(n5874));
  AOI21X1 g04292(.A0(n5696), .A1(n5703), .B0(n5874), .Y(n5875));
  AOI21X1 g04293(.A0(n5875), .A1(n5873), .B0(n5626), .Y(n5876));
  OAI21X1 g04294(.A0(n5872), .A1(n5871), .B0(n5876), .Y(n5877));
  NAND2X1 g04295(.A(n5634), .B(n3528), .Y(n5878));
  NAND2X1 g04296(.A(P1_U3086), .B(P1_REG3_REG_17__SCAN_IN), .Y(n5879));
  OAI22X1 g04297(.A0(n5621), .A1(n3527), .B0(n3578), .B1(n5639), .Y(n5880));
  AOI21X1 g04298(.A0(n5637), .A1(n3503), .B0(n5880), .Y(n5881));
  OAI21X1 g04299(.A0(n5881), .A1(n5636), .B0(n5879), .Y(n5882));
  AOI21X1 g04300(.A0(n5643), .A1(n3547), .B0(n5882), .Y(n5883));
  NAND3X1 g04301(.A(n5883), .B(n5878), .C(n5877), .Y(P1_U3228));
  NAND2X1 g04302(.A(n5598), .B(n5595), .Y(n5885));
  XOR2X1  g04303(.A(n5570), .B(n5568), .Y(n5886));
  XOR2X1  g04304(.A(n5886), .B(n5885), .Y(n5887));
  NAND2X1 g04305(.A(n5887), .B(n5743), .Y(n5888));
  NOR2X1  g04306(.A(n5633), .B(n2944), .Y(n5889));
  OAI22X1 g04307(.A0(n5621), .A1(n2944), .B0(n2898), .B1(n5751), .Y(n5890));
  AOI21X1 g04308(.A0(n5638), .A1(n3017), .B0(n5890), .Y(n5891));
  AOI22X1 g04309(.A0(n2966), .A1(n5643), .B0(P1_U3086), .B1(P1_REG3_REG_5__SCAN_IN), .Y(n5892));
  OAI21X1 g04310(.A0(n5891), .A1(n5636), .B0(n5892), .Y(n5893));
  NOR2X1  g04311(.A(n5893), .B(n5889), .Y(n5894));
  NAND2X1 g04312(.A(n5894), .B(n5888), .Y(P1_U3227));
  XOR2X1  g04313(.A(n5691), .B(n5689), .Y(n5896));
  NOR2X1  g04314(.A(n5896), .B(n5702), .Y(n5897));
  AOI21X1 g04315(.A0(n5896), .A1(n5702), .B0(n5897), .Y(n5899));
  OAI22X1 g04316(.A0(n5621), .A1(n3477), .B0(n3532), .B1(n5639), .Y(n5900));
  AOI21X1 g04317(.A0(n5637), .A1(n3489), .B0(n5900), .Y(n5901));
  AOI22X1 g04318(.A0(n3496), .A1(n5643), .B0(P1_U3086), .B1(P1_REG3_REG_16__SCAN_IN), .Y(n5902));
  OAI21X1 g04319(.A0(n5901), .A1(n5636), .B0(n5902), .Y(n5903));
  AOI21X1 g04320(.A0(n5634), .A1(n3478), .B0(n5903), .Y(n5904));
  OAI21X1 g04321(.A0(n5899), .A1(n5626), .B0(n5904), .Y(P1_U3226));
  XOR2X1  g04322(.A(n5729), .B(n5726), .Y(n5906));
  NOR2X1  g04323(.A(n5906), .B(n5725), .Y(n5908));
  AOI21X1 g04324(.A0(n5906), .A1(n5725), .B0(n5908), .Y(n5909));
  NOR2X1  g04325(.A(n5639), .B(n3924), .Y(n5910));
  OAI22X1 g04326(.A0(n5621), .A1(n3875), .B0(n3838), .B1(n5751), .Y(n5911));
  OAI21X1 g04327(.A0(n5911), .A1(n5910), .B0(n5635), .Y(n5912));
  AOI22X1 g04328(.A0(n4427), .A1(n5634), .B0(P1_U3086), .B1(P1_REG3_REG_25__SCAN_IN), .Y(n5913));
  NAND2X1 g04329(.A(n5913), .B(n5912), .Y(n5914));
  AOI21X1 g04330(.A0(n5643), .A1(n3887), .B0(n5914), .Y(n5915));
  OAI21X1 g04331(.A0(n5909), .A1(n5626), .B0(n5915), .Y(P1_U3225));
  XOR2X1  g04332(.A(n5544), .B(n5542), .Y(n5917));
  NOR2X1  g04333(.A(n5917), .B(n5809), .Y(n5919));
  AOI21X1 g04334(.A0(n5917), .A1(n5809), .B0(n5919), .Y(n5920));
  OAI22X1 g04335(.A0(n5621), .A1(n3293), .B0(n3346), .B1(n5639), .Y(n5921));
  AOI21X1 g04336(.A0(n5637), .A1(n3266), .B0(n5921), .Y(n5922));
  AOI22X1 g04337(.A0(n3313), .A1(n5643), .B0(P1_U3086), .B1(P1_REG3_REG_12__SCAN_IN), .Y(n5923));
  OAI21X1 g04338(.A0(n5922), .A1(n5636), .B0(n5923), .Y(n5924));
  AOI21X1 g04339(.A0(n5634), .A1(n3294), .B0(n5924), .Y(n5925));
  OAI21X1 g04340(.A0(n5920), .A1(n5626), .B0(n5925), .Y(P1_U3224));
  AOI21X1 g04341(.A0(n5671), .A1(n5669), .B0(n5676), .Y(n5927));
  OAI21X1 g04342(.A0(n5825), .A1(n5714), .B0(n5927), .Y(n5928));
  INVX1   g04343(.A(n5675), .Y(n5929));
  OAI21X1 g04344(.A0(n5671), .A1(n5719), .B0(n5715), .Y(n5930));
  AOI21X1 g04345(.A0(n5671), .A1(n5719), .B0(n5930), .Y(n5931));
  OAI21X1 g04346(.A0(n5824), .A1(n5929), .B0(n5931), .Y(n5932));
  NAND3X1 g04347(.A(n5932), .B(n5928), .C(n5743), .Y(n5933));
  NAND2X1 g04348(.A(n5643), .B(n3715), .Y(n5934));
  OAI22X1 g04349(.A0(n5621), .A1(n3705), .B0(n3666), .B1(n5751), .Y(n5935));
  AOI21X1 g04350(.A0(n5638), .A1(n3753), .B0(n5935), .Y(n5936));
  OAI22X1 g04351(.A0(n5636), .A1(n5936), .B0(P1_STATE_REG_SCAN_IN), .B1(n3703), .Y(n5937));
  AOI21X1 g04352(.A0(n5634), .A1(n4394), .B0(n5937), .Y(n5938));
  NAND3X1 g04353(.A(n5938), .B(n5934), .C(n5933), .Y(P1_U3223));
  XOR2X1  g04354(.A(n5583), .B(n5581), .Y(n5940));
  XOR2X1  g04355(.A(n5940), .B(n5588), .Y(n5941));
  NAND4X1 g04356(.A(n5625), .B(n5621), .C(n2560), .D(n5941), .Y(n5942));
  NAND2X1 g04357(.A(n5634), .B(P1_REG3_REG_1__SCAN_IN), .Y(n5943));
  AOI22X1 g04358(.A0(n5627), .A1(P1_REG3_REG_1__SCAN_IN), .B0(n2768), .B1(n5637), .Y(n5944));
  OAI21X1 g04359(.A0(n5639), .A1(n2799), .B0(n5944), .Y(n5945));
  OAI22X1 g04360(.A0(n2792), .A1(n5642), .B0(P1_STATE_REG_SCAN_IN), .B1(n2779), .Y(n5946));
  AOI21X1 g04361(.A0(n5945), .A1(n5635), .B0(n5946), .Y(n5947));
  NAND3X1 g04362(.A(n5947), .B(n5943), .C(n5942), .Y(P1_U3222));
  NAND2X1 g04363(.A(n5604), .B(n5600), .Y(n5949));
  XOR2X1  g04364(.A(n5559), .B(n5557), .Y(n5950));
  XOR2X1  g04365(.A(n5950), .B(n5949), .Y(n5951));
  NAND2X1 g04366(.A(n5951), .B(n5743), .Y(n5952));
  OAI22X1 g04367(.A0(n5621), .A1(n3100), .B0(n3050), .B1(n5751), .Y(n5953));
  AOI21X1 g04368(.A0(n5638), .A1(n3170), .B0(n5953), .Y(n5954));
  AOI22X1 g04369(.A0(n3120), .A1(n5643), .B0(P1_U3086), .B1(P1_REG3_REG_8__SCAN_IN), .Y(n5955));
  OAI21X1 g04370(.A0(n5954), .A1(n5636), .B0(n5955), .Y(n5956));
  AOI21X1 g04371(.A0(n5634), .A1(n3101), .B0(n5956), .Y(n5957));
  NAND2X1 g04372(.A(n5957), .B(n5952), .Y(P1_U3221));
  OAI22X1 g04373(.A0(n4962), .A1(n3973), .B0(n4011), .B1(n4975), .Y(n5959));
  XOR2X1  g04374(.A(n5959), .B(n4956), .Y(n5960));
  AOI22X1 g04375(.A0(n5520), .A1(n3972), .B0(n3988), .B1(n4976), .Y(n5961));
  INVX1   g04376(.A(n5961), .Y(n5962));
  NOR2X1  g04377(.A(n5962), .B(n5960), .Y(n5963));
  NOR3X1  g04378(.A(n5963), .B(n5736), .C(n5654), .Y(n5964));
  AOI22X1 g04379(.A0(n5520), .A1(n4019), .B0(n4032), .B1(n4976), .Y(n5965));
  XOR2X1  g04380(.A(n5965), .B(n4969), .Y(n5966));
  OAI22X1 g04381(.A0(n4962), .A1(n4020), .B0(n4059), .B1(n4975), .Y(n5967));
  XOR2X1  g04382(.A(n5967), .B(n5966), .Y(n5968));
  OAI21X1 g04383(.A0(n5962), .A1(n5960), .B0(n5739), .Y(n5969));
  AOI21X1 g04384(.A0(n5731), .A1(n5652), .B0(n5736), .Y(n5970));
  OAI21X1 g04385(.A0(n5962), .A1(n5960), .B0(n5970), .Y(n5971));
  NAND2X1 g04386(.A(n5962), .B(n5960), .Y(n5972));
  NAND4X1 g04387(.A(n5971), .B(n5969), .C(n5968), .D(n5972), .Y(n5973));
  AOI21X1 g04388(.A0(n5964), .A1(n5724), .B0(n5973), .Y(n5974));
  INVX1   g04389(.A(n5970), .Y(n5975));
  NAND3X1 g04390(.A(n5737), .B(n5724), .C(n5655), .Y(n5976));
  NAND4X1 g04391(.A(n5972), .B(n5975), .C(n5740), .D(n5976), .Y(n5977));
  NOR2X1  g04392(.A(n5968), .B(n5963), .Y(n5978));
  AOI21X1 g04393(.A0(n5978), .A1(n5977), .B0(n5974), .Y(n5979));
  NOR2X1  g04394(.A(n5751), .B(n3973), .Y(n5980));
  OAI22X1 g04395(.A0(n5621), .A1(n4015), .B0(n4064), .B1(n5639), .Y(n5981));
  OAI21X1 g04396(.A0(n5981), .A1(n5980), .B0(n5635), .Y(n5982));
  AOI22X1 g04397(.A0(n4455), .A1(n5634), .B0(P1_U3086), .B1(P1_REG3_REG_28__SCAN_IN), .Y(n5983));
  NAND2X1 g04398(.A(n5983), .B(n5982), .Y(n5984));
  AOI21X1 g04399(.A0(n5643), .A1(n4032), .B0(n5984), .Y(n5985));
  OAI21X1 g04400(.A0(n5979), .A1(n5626), .B0(n5985), .Y(P1_U3220));
  INVX1   g04401(.A(n5679), .Y(n5987));
  XOR2X1  g04402(.A(n5987), .B(n5678), .Y(n5988));
  NOR2X1  g04403(.A(n5988), .B(n5710), .Y(n5989));
  AOI21X1 g04404(.A0(n5988), .A1(n5710), .B0(n5989), .Y(n5991));
  AOI22X1 g04405(.A0(n5627), .A1(n3617), .B0(n3665), .B1(n5638), .Y(n5992));
  OAI21X1 g04406(.A0(n5751), .A1(n3578), .B0(n5992), .Y(n5993));
  AOI22X1 g04407(.A0(n5635), .A1(n5993), .B0(P1_U3086), .B1(P1_REG3_REG_19__SCAN_IN), .Y(n5994));
  OAI21X1 g04408(.A0(n5633), .A1(n3616), .B0(n5994), .Y(n5995));
  AOI21X1 g04409(.A0(n5643), .A1(n3627), .B0(n5995), .Y(n5996));
  OAI21X1 g04410(.A0(n5991), .A1(n5626), .B0(n5996), .Y(P1_U3219));
  INVX1   g04411(.A(n5589), .Y(n5998));
  NOR2X1  g04412(.A(n5575), .B(n5573), .Y(n5999));
  AOI21X1 g04413(.A0(n5579), .A1(n5577), .B0(n5580), .Y(n6000));
  OAI21X1 g04414(.A0(n5999), .A1(n5998), .B0(n6000), .Y(n6001));
  AOI21X1 g04415(.A0(n5579), .A1(n5590), .B0(n5999), .Y(n6002));
  OAI21X1 g04416(.A0(n5579), .A1(n5590), .B0(n6002), .Y(n6003));
  AOI21X1 g04417(.A0(n5998), .A1(n5576), .B0(n6003), .Y(n6004));
  NOR2X1  g04418(.A(n6004), .B(n5626), .Y(n6005));
  NAND2X1 g04419(.A(n6005), .B(n6001), .Y(n6006));
  NOR2X1  g04420(.A(n5633), .B(P1_REG3_REG_3__SCAN_IN), .Y(n6007));
  OAI22X1 g04421(.A0(n5621), .A1(P1_REG3_REG_3__SCAN_IN), .B0(n2799), .B1(n5751), .Y(n6008));
  AOI21X1 g04422(.A0(n5638), .A1(n2954), .B0(n6008), .Y(n6009));
  AOI22X1 g04423(.A0(n2870), .A1(n5643), .B0(P1_U3086), .B1(P1_REG3_REG_3__SCAN_IN), .Y(n6010));
  OAI21X1 g04424(.A0(n6009), .A1(n5636), .B0(n6010), .Y(n6011));
  NOR2X1  g04425(.A(n6011), .B(n6007), .Y(n6012));
  NAND2X1 g04426(.A(n6012), .B(n6006), .Y(P1_U3218));
  INVX1   g04427(.A(n5550), .Y(n6014));
  XOR2X1  g04428(.A(n5552), .B(n6014), .Y(n6015));
  XOR2X1  g04429(.A(n6015), .B(n5610), .Y(n6016));
  OAI22X1 g04430(.A0(n5621), .A1(n3193), .B0(n3153), .B1(n5751), .Y(n6017));
  AOI21X1 g04431(.A0(n5638), .A1(n3266), .B0(n6017), .Y(n6018));
  AOI22X1 g04432(.A0(n3215), .A1(n5643), .B0(P1_U3086), .B1(P1_REG3_REG_10__SCAN_IN), .Y(n6019));
  OAI21X1 g04433(.A0(n6018), .A1(n5636), .B0(n6019), .Y(n6020));
  AOI21X1 g04434(.A0(n5634), .A1(n3194), .B0(n6020), .Y(n6021));
  OAI21X1 g04435(.A0(n6016), .A1(n5626), .B0(n6021), .Y(P1_U3217));
  XOR2X1  g04436(.A(n5659), .B(n5656), .Y(n6023));
  XOR2X1  g04437(.A(n6023), .B(n5723), .Y(n6024));
  NOR2X1  g04438(.A(n5639), .B(n3838), .Y(n6025));
  OAI22X1 g04439(.A0(n5621), .A1(n3790), .B0(n3754), .B1(n5751), .Y(n6026));
  OAI21X1 g04440(.A0(n6026), .A1(n6025), .B0(n5635), .Y(n6027));
  AOI22X1 g04441(.A0(n4411), .A1(n5634), .B0(P1_U3086), .B1(P1_REG3_REG_23__SCAN_IN), .Y(n6028));
  NAND2X1 g04442(.A(n6028), .B(n6027), .Y(n6029));
  AOI21X1 g04443(.A0(n5643), .A1(n3804), .B0(n6029), .Y(n6030));
  OAI21X1 g04444(.A0(n6024), .A1(n5626), .B0(n6030), .Y(P1_U3216));
  XOR2X1  g04445(.A(n5525), .B(n5527), .Y(n6032));
  XOR2X1  g04446(.A(n6032), .B(n5614), .Y(n6033));
  OAI22X1 g04447(.A0(n5621), .A1(n3393), .B0(n3443), .B1(n5639), .Y(n6034));
  AOI21X1 g04448(.A0(n5637), .A1(n3345), .B0(n6034), .Y(n6035));
  AOI22X1 g04449(.A0(n3460), .A1(n5643), .B0(P1_U3086), .B1(P1_REG3_REG_14__SCAN_IN), .Y(n6036));
  OAI21X1 g04450(.A0(n6035), .A1(n5636), .B0(n6036), .Y(n6037));
  AOI21X1 g04451(.A0(n5634), .A1(n3394), .B0(n6037), .Y(n6038));
  OAI21X1 g04452(.A0(n6033), .A1(n5626), .B0(n6038), .Y(P1_U3215));
  NAND3X1 g04453(.A(n5976), .B(n5975), .C(n5740), .Y(n6040));
  XOR2X1  g04454(.A(n5961), .B(n5960), .Y(n6041));
  XOR2X1  g04455(.A(n6041), .B(n6040), .Y(n6042));
  NOR2X1  g04456(.A(n5639), .B(n4020), .Y(n6043));
  OAI22X1 g04457(.A0(n5621), .A1(n3968), .B0(n3924), .B1(n5751), .Y(n6044));
  OAI21X1 g04458(.A0(n6044), .A1(n6043), .B0(n5635), .Y(n6045));
  AOI22X1 g04459(.A0(n4446), .A1(n5634), .B0(P1_U3086), .B1(P1_REG3_REG_27__SCAN_IN), .Y(n6046));
  NAND2X1 g04460(.A(n6046), .B(n6045), .Y(n6047));
  AOI21X1 g04461(.A0(n5643), .A1(n3988), .B0(n6047), .Y(n6048));
  OAI21X1 g04462(.A0(n6042), .A1(n5626), .B0(n6048), .Y(P1_U3214));
  NOR2X1  g04463(.A(n5563), .B(n5561), .Y(n6050));
  NOR3X1  g04464(.A(n6050), .B(n5599), .C(n5571), .Y(n6051));
  OAI21X1 g04465(.A0(n5566), .A1(n5564), .B0(n5567), .Y(n6052));
  NOR2X1  g04466(.A(n6052), .B(n6051), .Y(n6053));
  AOI21X1 g04467(.A0(n5563), .A1(n5561), .B0(n5758), .Y(n6054));
  AOI21X1 g04468(.A0(n5601), .A1(n5564), .B0(n6050), .Y(n6055));
  OAI21X1 g04469(.A0(n5601), .A1(n5564), .B0(n6055), .Y(n6056));
  OAI21X1 g04470(.A0(n6056), .A1(n6054), .B0(n5743), .Y(n6057));
  OAI22X1 g04471(.A0(n5621), .A1(n3046), .B0(n2998), .B1(n5751), .Y(n6058));
  AOI21X1 g04472(.A0(n5638), .A1(n3103), .B0(n6058), .Y(n6059));
  AOI22X1 g04473(.A0(n3067), .A1(n5643), .B0(P1_U3086), .B1(P1_REG3_REG_7__SCAN_IN), .Y(n6060));
  OAI21X1 g04474(.A0(n6059), .A1(n5636), .B0(n6060), .Y(n6061));
  AOI21X1 g04475(.A0(n5634), .A1(n3047), .B0(n6061), .Y(n6062));
  OAI21X1 g04476(.A0(n6057), .A1(n6053), .B0(n6062), .Y(P1_U3213));
  AOI21X1 g04477(.A0(n1789), .A1(n1786), .B0(n1796), .Y(n6064));
  AOI21X1 g04478(.A0(n1800), .A1(n1837), .B0(n6064), .Y(n6065));
  INVX1   g04479(.A(P2_STATE_REG_SCAN_IN), .Y(P2_U3088));
  NOR2X1  g04480(.A(P2_U3088), .B(P2_IR_REG_31__SCAN_IN), .Y(n6067));
  OAI21X1 g04481(.A0(n6067), .A1(P2_STATE_REG_SCAN_IN), .B0(P2_IR_REG_0__SCAN_IN), .Y(n6068));
  OAI21X1 g04482(.A0(n6065), .A1(P2_STATE_REG_SCAN_IN), .B0(n6068), .Y(P2_U3327));
  AOI21X1 g04483(.A0(n1789), .A1(n1786), .B0(n1808), .Y(n6070));
  AOI21X1 g04484(.A0(n1825), .A1(n1837), .B0(n6070), .Y(n6071));
  INVX1   g04485(.A(P2_IR_REG_31__SCAN_IN), .Y(n6072));
  NOR2X1  g04486(.A(P2_U3088), .B(n6072), .Y(n6073));
  XOR2X1  g04487(.A(P2_IR_REG_1__SCAN_IN), .B(P2_IR_REG_0__SCAN_IN), .Y(n6074));
  AOI22X1 g04488(.A0(n6073), .A1(n6074), .B0(n6067), .B1(P2_IR_REG_1__SCAN_IN), .Y(n6075));
  OAI21X1 g04489(.A0(n6071), .A1(P2_STATE_REG_SCAN_IN), .B0(n6075), .Y(P2_U3326));
  AOI21X1 g04490(.A0(n1789), .A1(n1786), .B0(n1854), .Y(n6077));
  AOI21X1 g04491(.A0(n1841), .A1(n1837), .B0(n6077), .Y(n6078));
  INVX1   g04492(.A(P2_IR_REG_2__SCAN_IN), .Y(n6079));
  NOR2X1  g04493(.A(P2_IR_REG_1__SCAN_IN), .B(P2_IR_REG_0__SCAN_IN), .Y(n6080));
  XOR2X1  g04494(.A(n6080), .B(n6079), .Y(n6081));
  AOI22X1 g04495(.A0(n6073), .A1(n6081), .B0(n6067), .B1(P2_IR_REG_2__SCAN_IN), .Y(n6082));
  OAI21X1 g04496(.A0(n6078), .A1(P2_STATE_REG_SCAN_IN), .B0(n6082), .Y(P2_U3325));
  AOI21X1 g04497(.A0(n1789), .A1(n1786), .B0(n1875), .Y(n6084));
  AOI21X1 g04498(.A0(n1864), .A1(n1837), .B0(n6084), .Y(n6085));
  INVX1   g04499(.A(P2_IR_REG_3__SCAN_IN), .Y(n6086));
  NOR3X1  g04500(.A(P2_IR_REG_2__SCAN_IN), .B(P2_IR_REG_1__SCAN_IN), .C(P2_IR_REG_0__SCAN_IN), .Y(n6087));
  XOR2X1  g04501(.A(n6087), .B(n6086), .Y(n6088));
  AOI22X1 g04502(.A0(n6073), .A1(n6088), .B0(n6067), .B1(P2_IR_REG_3__SCAN_IN), .Y(n6089));
  OAI21X1 g04503(.A0(n6085), .A1(P2_STATE_REG_SCAN_IN), .B0(n6089), .Y(P2_U3324));
  AOI21X1 g04504(.A0(n1789), .A1(n1786), .B0(n1884), .Y(n6091));
  AOI21X1 g04505(.A0(n1889), .A1(n1837), .B0(n6091), .Y(n6092));
  INVX1   g04506(.A(P2_IR_REG_4__SCAN_IN), .Y(n6093));
  NOR4X1  g04507(.A(P2_IR_REG_2__SCAN_IN), .B(P2_IR_REG_1__SCAN_IN), .C(P2_IR_REG_0__SCAN_IN), .D(P2_IR_REG_3__SCAN_IN), .Y(n6094));
  INVX1   g04508(.A(n6087), .Y(n6095));
  NOR3X1  g04509(.A(n6095), .B(P2_IR_REG_4__SCAN_IN), .C(P2_IR_REG_3__SCAN_IN), .Y(n6096));
  INVX1   g04510(.A(n6096), .Y(n6097));
  OAI21X1 g04511(.A0(n6094), .A1(n6093), .B0(n6097), .Y(n6098));
  NOR3X1  g04512(.A(n6098), .B(P2_U3088), .C(n6072), .Y(n6099));
  AOI21X1 g04513(.A0(n6067), .A1(P2_IR_REG_4__SCAN_IN), .B0(n6099), .Y(n6100));
  OAI21X1 g04514(.A0(n6092), .A1(P2_STATE_REG_SCAN_IN), .B0(n6100), .Y(P2_U3323));
  AOI21X1 g04515(.A0(n1921), .A1(n1910), .B0(n1790), .Y(n6102));
  AOI21X1 g04516(.A0(n1789), .A1(n1786), .B0(n1904), .Y(n6103));
  NOR2X1  g04517(.A(n6103), .B(n6102), .Y(n6104));
  INVX1   g04518(.A(P2_IR_REG_5__SCAN_IN), .Y(n6105));
  XOR2X1  g04519(.A(n6096), .B(n6105), .Y(n6106));
  AOI22X1 g04520(.A0(n6073), .A1(n6106), .B0(n6067), .B1(P2_IR_REG_5__SCAN_IN), .Y(n6107));
  OAI21X1 g04521(.A0(n6104), .A1(P2_STATE_REG_SCAN_IN), .B0(n6107), .Y(P2_U3322));
  AOI21X1 g04522(.A0(n1789), .A1(n1786), .B0(n1935), .Y(n6109));
  AOI21X1 g04523(.A0(n1940), .A1(n1837), .B0(n6109), .Y(n6110));
  INVX1   g04524(.A(P2_IR_REG_6__SCAN_IN), .Y(n6111));
  AOI21X1 g04525(.A0(n6096), .A1(n6105), .B0(n6111), .Y(n6112));
  NOR3X1  g04526(.A(n6097), .B(P2_IR_REG_6__SCAN_IN), .C(P2_IR_REG_5__SCAN_IN), .Y(n6113));
  NOR2X1  g04527(.A(n6113), .B(n6112), .Y(n6114));
  AOI22X1 g04528(.A0(n6073), .A1(n6114), .B0(n6067), .B1(P2_IR_REG_6__SCAN_IN), .Y(n6115));
  OAI21X1 g04529(.A0(n6110), .A1(P2_STATE_REG_SCAN_IN), .B0(n6115), .Y(P2_U3321));
  AOI21X1 g04530(.A0(n1789), .A1(n1786), .B0(n1963), .Y(n6117));
  AOI21X1 g04531(.A0(n1968), .A1(n1837), .B0(n6117), .Y(n6118));
  INVX1   g04532(.A(P2_IR_REG_7__SCAN_IN), .Y(n6119));
  XOR2X1  g04533(.A(n6113), .B(n6119), .Y(n6120));
  AOI22X1 g04534(.A0(n6073), .A1(n6120), .B0(n6067), .B1(P2_IR_REG_7__SCAN_IN), .Y(n6121));
  OAI21X1 g04535(.A0(n6118), .A1(P2_STATE_REG_SCAN_IN), .B0(n6121), .Y(P2_U3320));
  AOI21X1 g04536(.A0(n1789), .A1(n1786), .B0(n5069), .Y(n6123));
  AOI21X1 g04537(.A0(n1989), .A1(n1837), .B0(n6123), .Y(n6124));
  NAND4X1 g04538(.A(n6119), .B(n6111), .C(n6105), .D(n6096), .Y(n6125));
  NOR4X1  g04539(.A(P2_IR_REG_5__SCAN_IN), .B(P2_IR_REG_4__SCAN_IN), .C(P2_IR_REG_3__SCAN_IN), .D(P2_IR_REG_6__SCAN_IN), .Y(n6126));
  INVX1   g04540(.A(n6126), .Y(n6127));
  NOR4X1  g04541(.A(n6095), .B(P2_IR_REG_8__SCAN_IN), .C(P2_IR_REG_7__SCAN_IN), .D(n6127), .Y(n6128));
  AOI21X1 g04542(.A0(n6125), .A1(P2_IR_REG_8__SCAN_IN), .B0(n6128), .Y(n6129));
  AOI22X1 g04543(.A0(n6073), .A1(n6129), .B0(n6067), .B1(P2_IR_REG_8__SCAN_IN), .Y(n6130));
  OAI21X1 g04544(.A0(n6124), .A1(P2_STATE_REG_SCAN_IN), .B0(n6130), .Y(P2_U3319));
  AOI21X1 g04545(.A0(n1789), .A1(n1786), .B0(n2020), .Y(n6132));
  AOI21X1 g04546(.A0(n2013), .A1(n1837), .B0(n6132), .Y(n6133));
  INVX1   g04547(.A(P2_IR_REG_9__SCAN_IN), .Y(n6134));
  XOR2X1  g04548(.A(n6128), .B(n6134), .Y(n6135));
  AOI22X1 g04549(.A0(n6073), .A1(n6135), .B0(n6067), .B1(P2_IR_REG_9__SCAN_IN), .Y(n6136));
  OAI21X1 g04550(.A0(n6133), .A1(P2_STATE_REG_SCAN_IN), .B0(n6136), .Y(P2_U3318));
  AOI21X1 g04551(.A0(n1789), .A1(n1786), .B0(n2045), .Y(n6138));
  AOI21X1 g04552(.A0(n2032), .A1(n1837), .B0(n6138), .Y(n6139));
  INVX1   g04553(.A(P2_IR_REG_10__SCAN_IN), .Y(n6140));
  AOI21X1 g04554(.A0(n6128), .A1(n6134), .B0(n6140), .Y(n6141));
  NOR2X1  g04555(.A(P2_IR_REG_10__SCAN_IN), .B(P2_IR_REG_9__SCAN_IN), .Y(n6142));
  AOI21X1 g04556(.A0(n6142), .A1(n6128), .B0(n6141), .Y(n6143));
  AOI22X1 g04557(.A0(n6073), .A1(n6143), .B0(n6067), .B1(P2_IR_REG_10__SCAN_IN), .Y(n6144));
  OAI21X1 g04558(.A0(n6139), .A1(P2_STATE_REG_SCAN_IN), .B0(n6144), .Y(P2_U3317));
  AOI21X1 g04559(.A0(n1789), .A1(n1786), .B0(n5076), .Y(n6146));
  AOI21X1 g04560(.A0(n2059), .A1(n1837), .B0(n6146), .Y(n6147));
  INVX1   g04561(.A(P2_IR_REG_11__SCAN_IN), .Y(n6148));
  INVX1   g04562(.A(n6128), .Y(n6149));
  INVX1   g04563(.A(n6142), .Y(n6150));
  NOR2X1  g04564(.A(n6150), .B(n6149), .Y(n6151));
  XOR2X1  g04565(.A(n6151), .B(n6148), .Y(n6152));
  AOI22X1 g04566(.A0(n6073), .A1(n6152), .B0(n6067), .B1(P2_IR_REG_11__SCAN_IN), .Y(n6153));
  OAI21X1 g04567(.A0(n6147), .A1(P2_STATE_REG_SCAN_IN), .B0(n6153), .Y(P2_U3316));
  AOI21X1 g04568(.A0(n1789), .A1(n1786), .B0(n5079), .Y(n6155));
  AOI21X1 g04569(.A0(n2080), .A1(n1837), .B0(n6155), .Y(n6156));
  NAND3X1 g04570(.A(n6142), .B(n6128), .C(n6148), .Y(n6157));
  NOR4X1  g04571(.A(n6149), .B(P2_IR_REG_12__SCAN_IN), .C(P2_IR_REG_11__SCAN_IN), .D(n6150), .Y(n6158));
  AOI21X1 g04572(.A0(n6157), .A1(P2_IR_REG_12__SCAN_IN), .B0(n6158), .Y(n6159));
  AOI22X1 g04573(.A0(n6073), .A1(n6159), .B0(n6067), .B1(P2_IR_REG_12__SCAN_IN), .Y(n6160));
  OAI21X1 g04574(.A0(n6156), .A1(P2_STATE_REG_SCAN_IN), .B0(n6160), .Y(P2_U3315));
  AOI21X1 g04575(.A0(n1789), .A1(n1786), .B0(n2099), .Y(n6162));
  AOI21X1 g04576(.A0(n2103), .A1(n1837), .B0(n6162), .Y(n6163));
  INVX1   g04577(.A(P2_IR_REG_13__SCAN_IN), .Y(n6164));
  XOR2X1  g04578(.A(n6158), .B(n6164), .Y(n6165));
  AOI22X1 g04579(.A0(n6073), .A1(n6165), .B0(n6067), .B1(P2_IR_REG_13__SCAN_IN), .Y(n6166));
  OAI21X1 g04580(.A0(n6163), .A1(P2_STATE_REG_SCAN_IN), .B0(n6166), .Y(P2_U3314));
  AOI21X1 g04581(.A0(n1789), .A1(n1786), .B0(n2131), .Y(n6168));
  AOI21X1 g04582(.A0(n2119), .A1(n1837), .B0(n6168), .Y(n6169));
  INVX1   g04583(.A(P2_IR_REG_14__SCAN_IN), .Y(n6170));
  AOI21X1 g04584(.A0(n6158), .A1(n6164), .B0(n6170), .Y(n6171));
  INVX1   g04585(.A(n6158), .Y(n6172));
  NOR3X1  g04586(.A(n6172), .B(P2_IR_REG_14__SCAN_IN), .C(P2_IR_REG_13__SCAN_IN), .Y(n6173));
  NOR2X1  g04587(.A(n6173), .B(n6171), .Y(n6174));
  AOI22X1 g04588(.A0(n6073), .A1(n6174), .B0(n6067), .B1(P2_IR_REG_14__SCAN_IN), .Y(n6175));
  OAI21X1 g04589(.A0(n6169), .A1(P2_STATE_REG_SCAN_IN), .B0(n6175), .Y(P2_U3313));
  INVX1   g04590(.A(P1_DATAO_REG_15__SCAN_IN), .Y(n6177));
  AOI21X1 g04591(.A0(n1789), .A1(n1786), .B0(n6177), .Y(n6178));
  AOI21X1 g04592(.A0(n2142), .A1(n1837), .B0(n6178), .Y(n6179));
  INVX1   g04593(.A(P2_IR_REG_15__SCAN_IN), .Y(n6180));
  XOR2X1  g04594(.A(n6173), .B(n6180), .Y(n6181));
  AOI22X1 g04595(.A0(n6073), .A1(n6181), .B0(n6067), .B1(P2_IR_REG_15__SCAN_IN), .Y(n6182));
  OAI21X1 g04596(.A0(n6179), .A1(P2_STATE_REG_SCAN_IN), .B0(n6182), .Y(P2_U3312));
  INVX1   g04597(.A(P1_DATAO_REG_16__SCAN_IN), .Y(n6184));
  AOI21X1 g04598(.A0(n1789), .A1(n1786), .B0(n6184), .Y(n6185));
  AOI21X1 g04599(.A0(n2164), .A1(n1837), .B0(n6185), .Y(n6186));
  INVX1   g04600(.A(P2_IR_REG_16__SCAN_IN), .Y(n6187));
  NOR4X1  g04601(.A(P2_IR_REG_15__SCAN_IN), .B(P2_IR_REG_14__SCAN_IN), .C(P2_IR_REG_13__SCAN_IN), .D(n6172), .Y(n6188));
  NOR4X1  g04602(.A(P2_IR_REG_4__SCAN_IN), .B(P2_IR_REG_3__SCAN_IN), .C(P2_IR_REG_2__SCAN_IN), .D(P2_IR_REG_14__SCAN_IN), .Y(n6189));
  NAND2X1 g04603(.A(n6189), .B(n6080), .Y(n6190));
  INVX1   g04604(.A(P2_IR_REG_12__SCAN_IN), .Y(n6191));
  NAND4X1 g04605(.A(n6191), .B(n6148), .C(n6140), .D(n6164), .Y(n6192));
  NOR4X1  g04606(.A(P2_IR_REG_7__SCAN_IN), .B(P2_IR_REG_6__SCAN_IN), .C(P2_IR_REG_5__SCAN_IN), .D(P2_IR_REG_8__SCAN_IN), .Y(n6193));
  NAND4X1 g04607(.A(n6187), .B(n6180), .C(n6134), .D(n6193), .Y(n6194));
  NOR3X1  g04608(.A(n6194), .B(n6192), .C(n6190), .Y(n6195));
  INVX1   g04609(.A(n6195), .Y(n6196));
  OAI21X1 g04610(.A0(n6188), .A1(n6187), .B0(n6196), .Y(n6197));
  INVX1   g04611(.A(n6197), .Y(n6198));
  AOI22X1 g04612(.A0(n6073), .A1(n6198), .B0(n6067), .B1(P2_IR_REG_16__SCAN_IN), .Y(n6199));
  OAI21X1 g04613(.A0(n6186), .A1(P2_STATE_REG_SCAN_IN), .B0(n6199), .Y(P2_U3311));
  INVX1   g04614(.A(P1_DATAO_REG_17__SCAN_IN), .Y(n6201));
  AOI21X1 g04615(.A0(n1789), .A1(n1786), .B0(n6201), .Y(n6202));
  AOI21X1 g04616(.A0(n2193), .A1(n1837), .B0(n6202), .Y(n6203));
  INVX1   g04617(.A(P2_IR_REG_17__SCAN_IN), .Y(n6204));
  XOR2X1  g04618(.A(n6195), .B(n6204), .Y(n6205));
  AOI22X1 g04619(.A0(n6073), .A1(n6205), .B0(n6067), .B1(P2_IR_REG_17__SCAN_IN), .Y(n6206));
  OAI21X1 g04620(.A0(n6203), .A1(P2_STATE_REG_SCAN_IN), .B0(n6206), .Y(P2_U3310));
  INVX1   g04621(.A(P1_DATAO_REG_18__SCAN_IN), .Y(n6208));
  AOI21X1 g04622(.A0(n1789), .A1(n1786), .B0(n6208), .Y(n6209));
  AOI21X1 g04623(.A0(n2211), .A1(n1837), .B0(n6209), .Y(n6210));
  INVX1   g04624(.A(P2_IR_REG_18__SCAN_IN), .Y(n6211));
  NOR4X1  g04625(.A(n6192), .B(n6190), .C(P2_IR_REG_17__SCAN_IN), .D(n6194), .Y(n6212));
  NOR2X1  g04626(.A(P2_IR_REG_18__SCAN_IN), .B(P2_IR_REG_17__SCAN_IN), .Y(n6213));
  NAND2X1 g04627(.A(n6213), .B(n6195), .Y(n6214));
  OAI21X1 g04628(.A0(n6212), .A1(n6211), .B0(n6214), .Y(n6215));
  INVX1   g04629(.A(n6215), .Y(n6216));
  AOI22X1 g04630(.A0(n6073), .A1(n6216), .B0(n6067), .B1(P2_IR_REG_18__SCAN_IN), .Y(n6217));
  OAI21X1 g04631(.A0(n6210), .A1(P2_STATE_REG_SCAN_IN), .B0(n6217), .Y(P2_U3309));
  INVX1   g04632(.A(P1_DATAO_REG_19__SCAN_IN), .Y(n6219));
  AOI21X1 g04633(.A0(n1789), .A1(n1786), .B0(n6219), .Y(n6220));
  AOI21X1 g04634(.A0(n2239), .A1(n1837), .B0(n6220), .Y(n6221));
  XOR2X1  g04635(.A(n6214), .B(P2_IR_REG_19__SCAN_IN), .Y(n6222));
  AOI22X1 g04636(.A0(n6073), .A1(n6222), .B0(n6067), .B1(P2_IR_REG_19__SCAN_IN), .Y(n6223));
  OAI21X1 g04637(.A0(n6221), .A1(P2_STATE_REG_SCAN_IN), .B0(n6223), .Y(P2_U3308));
  NOR2X1  g04638(.A(n2261), .B(n1790), .Y(n6225));
  INVX1   g04639(.A(P1_DATAO_REG_20__SCAN_IN), .Y(n6226));
  AOI21X1 g04640(.A0(n1789), .A1(n1786), .B0(n6226), .Y(n6227));
  NOR2X1  g04641(.A(n6227), .B(n6225), .Y(n6228));
  INVX1   g04642(.A(P2_IR_REG_19__SCAN_IN), .Y(n6229));
  NAND3X1 g04643(.A(n6213), .B(n6195), .C(n6229), .Y(n6230));
  XOR2X1  g04644(.A(n6230), .B(P2_IR_REG_20__SCAN_IN), .Y(n6231));
  AOI22X1 g04645(.A0(n6073), .A1(n6231), .B0(n6067), .B1(P2_IR_REG_20__SCAN_IN), .Y(n6232));
  OAI21X1 g04646(.A0(n6228), .A1(P2_STATE_REG_SCAN_IN), .B0(n6232), .Y(P2_U3307));
  INVX1   g04647(.A(P1_DATAO_REG_21__SCAN_IN), .Y(n6234));
  AOI21X1 g04648(.A0(n1789), .A1(n1786), .B0(n6234), .Y(n6235));
  AOI21X1 g04649(.A0(n2283), .A1(n1837), .B0(n6235), .Y(n6236));
  INVX1   g04650(.A(P2_IR_REG_20__SCAN_IN), .Y(n6237));
  NAND4X1 g04651(.A(n6195), .B(n6237), .C(n6229), .D(n6213), .Y(n6238));
  XOR2X1  g04652(.A(n6238), .B(P2_IR_REG_21__SCAN_IN), .Y(n6239));
  AOI22X1 g04653(.A0(n6073), .A1(n6239), .B0(n6067), .B1(P2_IR_REG_21__SCAN_IN), .Y(n6240));
  OAI21X1 g04654(.A0(n6236), .A1(P2_STATE_REG_SCAN_IN), .B0(n6240), .Y(P2_U3306));
  INVX1   g04655(.A(P1_DATAO_REG_22__SCAN_IN), .Y(n6242));
  AOI21X1 g04656(.A0(n1789), .A1(n1786), .B0(n6242), .Y(n6243));
  AOI21X1 g04657(.A0(n2305), .A1(n1837), .B0(n6243), .Y(n6244));
  INVX1   g04658(.A(P2_IR_REG_22__SCAN_IN), .Y(n6245));
  NOR2X1  g04659(.A(n6238), .B(P2_IR_REG_21__SCAN_IN), .Y(n6246));
  XOR2X1  g04660(.A(n6246), .B(n6245), .Y(n6247));
  AOI22X1 g04661(.A0(n6073), .A1(n6247), .B0(n6067), .B1(P2_IR_REG_22__SCAN_IN), .Y(n6248));
  OAI21X1 g04662(.A0(n6244), .A1(P2_STATE_REG_SCAN_IN), .B0(n6248), .Y(P2_U3305));
  INVX1   g04663(.A(P1_DATAO_REG_23__SCAN_IN), .Y(n6250));
  AOI21X1 g04664(.A0(n1789), .A1(n1786), .B0(n6250), .Y(n6251));
  AOI21X1 g04665(.A0(n2331), .A1(n1837), .B0(n6251), .Y(n6252));
  INVX1   g04666(.A(P2_IR_REG_23__SCAN_IN), .Y(n6253));
  AOI21X1 g04667(.A0(n6246), .A1(n6245), .B0(n6253), .Y(n6254));
  NOR4X1  g04668(.A(P2_IR_REG_23__SCAN_IN), .B(P2_IR_REG_22__SCAN_IN), .C(P2_IR_REG_21__SCAN_IN), .D(n6238), .Y(n6255));
  NOR4X1  g04669(.A(n6254), .B(P2_U3088), .C(n6072), .D(n6255), .Y(n6256));
  AOI21X1 g04670(.A0(n6067), .A1(P2_IR_REG_23__SCAN_IN), .B0(n6256), .Y(n6257));
  OAI21X1 g04671(.A0(n6252), .A1(P2_STATE_REG_SCAN_IN), .B0(n6257), .Y(P2_U3304));
  INVX1   g04672(.A(P1_DATAO_REG_24__SCAN_IN), .Y(n6259));
  AOI21X1 g04673(.A0(n1789), .A1(n1786), .B0(n6259), .Y(n6260));
  AOI21X1 g04674(.A0(n2357), .A1(n1837), .B0(n6260), .Y(n6261));
  INVX1   g04675(.A(P2_IR_REG_24__SCAN_IN), .Y(n6262));
  XOR2X1  g04676(.A(n6255), .B(n6262), .Y(n6263));
  AOI22X1 g04677(.A0(n6073), .A1(n6263), .B0(n6067), .B1(P2_IR_REG_24__SCAN_IN), .Y(n6264));
  OAI21X1 g04678(.A0(n6261), .A1(P2_STATE_REG_SCAN_IN), .B0(n6264), .Y(P2_U3303));
  INVX1   g04679(.A(P1_DATAO_REG_25__SCAN_IN), .Y(n6266));
  AOI21X1 g04680(.A0(n1789), .A1(n1786), .B0(n6266), .Y(n6267));
  AOI21X1 g04681(.A0(n2383), .A1(n1837), .B0(n6267), .Y(n6268));
  NAND2X1 g04682(.A(n6255), .B(n6262), .Y(n6269));
  XOR2X1  g04683(.A(n6269), .B(P2_IR_REG_25__SCAN_IN), .Y(n6270));
  AOI22X1 g04684(.A0(n6073), .A1(n6270), .B0(n6067), .B1(P2_IR_REG_25__SCAN_IN), .Y(n6271));
  OAI21X1 g04685(.A0(n6268), .A1(P2_STATE_REG_SCAN_IN), .B0(n6271), .Y(P2_U3302));
  AOI21X1 g04686(.A0(n2405), .A1(n2400), .B0(n1790), .Y(n6273));
  INVX1   g04687(.A(P1_DATAO_REG_26__SCAN_IN), .Y(n6274));
  AOI21X1 g04688(.A0(n1789), .A1(n1786), .B0(n6274), .Y(n6275));
  NOR2X1  g04689(.A(n6275), .B(n6273), .Y(n6276));
  INVX1   g04690(.A(P2_IR_REG_26__SCAN_IN), .Y(n6277));
  NOR2X1  g04691(.A(n6269), .B(P2_IR_REG_25__SCAN_IN), .Y(n6278));
  NOR2X1  g04692(.A(n6278), .B(n6277), .Y(n6279));
  NOR3X1  g04693(.A(P2_IR_REG_21__SCAN_IN), .B(P2_IR_REG_20__SCAN_IN), .C(P2_IR_REG_19__SCAN_IN), .Y(n6280));
  NAND3X1 g04694(.A(n6187), .B(n6180), .C(n6170), .Y(n6281));
  NOR2X1  g04695(.A(n6281), .B(n6192), .Y(n6282));
  NAND4X1 g04696(.A(n6280), .B(n6213), .C(n6080), .D(n6282), .Y(n6283));
  NOR4X1  g04697(.A(P2_IR_REG_6__SCAN_IN), .B(P2_IR_REG_5__SCAN_IN), .C(P2_IR_REG_4__SCAN_IN), .D(P2_IR_REG_26__SCAN_IN), .Y(n6284));
  NAND3X1 g04698(.A(n6284), .B(n6086), .C(n6079), .Y(n6285));
  INVX1   g04699(.A(P2_IR_REG_25__SCAN_IN), .Y(n6286));
  NAND4X1 g04700(.A(n6262), .B(n6253), .C(n6245), .D(n6286), .Y(n6287));
  INVX1   g04701(.A(P2_IR_REG_8__SCAN_IN), .Y(n6288));
  NAND3X1 g04702(.A(n6134), .B(n6288), .C(n6119), .Y(n6289));
  NOR4X1  g04703(.A(n6287), .B(n6285), .C(n6283), .D(n6289), .Y(n6290));
  NOR2X1  g04704(.A(n6290), .B(n6279), .Y(n6291));
  AOI22X1 g04705(.A0(n6073), .A1(n6291), .B0(n6067), .B1(P2_IR_REG_26__SCAN_IN), .Y(n6292));
  OAI21X1 g04706(.A0(n6276), .A1(P2_STATE_REG_SCAN_IN), .B0(n6292), .Y(P2_U3301));
  AOI21X1 g04707(.A0(n2434), .A1(n2432), .B0(n1790), .Y(n6294));
  INVX1   g04708(.A(P1_DATAO_REG_27__SCAN_IN), .Y(n6295));
  AOI21X1 g04709(.A0(n1789), .A1(n1786), .B0(n6295), .Y(n6296));
  NOR2X1  g04710(.A(n6296), .B(n6294), .Y(n6297));
  INVX1   g04711(.A(P2_IR_REG_27__SCAN_IN), .Y(n6298));
  XOR2X1  g04712(.A(n6290), .B(n6298), .Y(n6299));
  AOI22X1 g04713(.A0(n6073), .A1(n6299), .B0(n6067), .B1(P2_IR_REG_27__SCAN_IN), .Y(n6300));
  OAI21X1 g04714(.A0(n6297), .A1(P2_STATE_REG_SCAN_IN), .B0(n6300), .Y(P2_U3300));
  INVX1   g04715(.A(P1_DATAO_REG_28__SCAN_IN), .Y(n6302));
  AOI21X1 g04716(.A0(n1789), .A1(n1786), .B0(n6302), .Y(n6303));
  AOI21X1 g04717(.A0(n2450), .A1(n1837), .B0(n6303), .Y(n6304));
  INVX1   g04718(.A(P2_IR_REG_28__SCAN_IN), .Y(n6305));
  NAND4X1 g04719(.A(n6134), .B(n6288), .C(n6119), .D(n6126), .Y(n6306));
  NAND3X1 g04720(.A(n6298), .B(n6277), .C(n6079), .Y(n6307));
  NOR4X1  g04721(.A(n6306), .B(n6287), .C(n6283), .D(n6307), .Y(n6308));
  XOR2X1  g04722(.A(n6308), .B(n6305), .Y(n6309));
  AOI22X1 g04723(.A0(n6073), .A1(n6309), .B0(n6067), .B1(P2_IR_REG_28__SCAN_IN), .Y(n6310));
  OAI21X1 g04724(.A0(n6304), .A1(P2_STATE_REG_SCAN_IN), .B0(n6310), .Y(P2_U3299));
  INVX1   g04725(.A(P1_DATAO_REG_29__SCAN_IN), .Y(n6312));
  OAI21X1 g04726(.A0(n4111), .A1(n4110), .B0(n1837), .Y(n6313));
  OAI21X1 g04727(.A0(n1837), .A1(n6312), .B0(n6313), .Y(n6314));
  INVX1   g04728(.A(n6314), .Y(n6315));
  NOR4X1  g04729(.A(P2_IR_REG_19__SCAN_IN), .B(P2_IR_REG_18__SCAN_IN), .C(P2_IR_REG_17__SCAN_IN), .D(P2_IR_REG_21__SCAN_IN), .Y(n6316));
  NAND4X1 g04730(.A(n6080), .B(n6245), .C(n6237), .D(n6316), .Y(n6317));
  NOR3X1  g04731(.A(n6317), .B(n6281), .C(n6192), .Y(n6318));
  NAND4X1 g04732(.A(n6286), .B(n6262), .C(n6253), .D(n6277), .Y(n6319));
  NAND3X1 g04733(.A(n6305), .B(n6298), .C(n6079), .Y(n6320));
  NOR3X1  g04734(.A(n6320), .B(n6319), .C(n6306), .Y(n6321));
  NAND2X1 g04735(.A(n6321), .B(n6318), .Y(n6322));
  NOR4X1  g04736(.A(n6319), .B(n6306), .C(P2_IR_REG_29__SCAN_IN), .D(n6320), .Y(n6323));
  AOI22X1 g04737(.A0(n6322), .A1(P2_IR_REG_29__SCAN_IN), .B0(n6318), .B1(n6323), .Y(n6324));
  AOI22X1 g04738(.A0(n6073), .A1(n6324), .B0(n6067), .B1(P2_IR_REG_29__SCAN_IN), .Y(n6325));
  OAI21X1 g04739(.A0(n6315), .A1(P2_STATE_REG_SCAN_IN), .B0(n6325), .Y(P2_U3298));
  AOI21X1 g04740(.A0(n4122), .A1(n4121), .B0(n1790), .Y(n6327));
  AOI21X1 g04741(.A0(n1789), .A1(n1786), .B0(n5116), .Y(n6328));
  OAI21X1 g04742(.A0(n6328), .A1(n6327), .B0(P2_U3088), .Y(n6329));
  NAND2X1 g04743(.A(n6323), .B(n6318), .Y(n6330));
  XOR2X1  g04744(.A(n6330), .B(P2_IR_REG_30__SCAN_IN), .Y(n6331));
  AOI22X1 g04745(.A0(n6073), .A1(n6331), .B0(n6067), .B1(P2_IR_REG_30__SCAN_IN), .Y(n6332));
  NAND2X1 g04746(.A(n6332), .B(n6329), .Y(P2_U3297));
  NOR4X1  g04747(.A(n2523), .B(n2519), .C(n1790), .D(n2527), .Y(n6334));
  AOI21X1 g04748(.A0(n1789), .A1(n1786), .B0(n5121), .Y(n6335));
  OAI21X1 g04749(.A0(n6335), .A1(n6334), .B0(P2_U3088), .Y(n6336));
  NOR2X1  g04750(.A(n6330), .B(P2_IR_REG_30__SCAN_IN), .Y(n6337));
  NAND3X1 g04751(.A(n6337), .B(P2_STATE_REG_SCAN_IN), .C(P2_IR_REG_31__SCAN_IN), .Y(n6338));
  NAND2X1 g04752(.A(n6338), .B(n6336), .Y(P2_U3296));
  NOR3X1  g04753(.A(n6255), .B(n6254), .C(n6072), .Y(n6340));
  AOI21X1 g04754(.A0(n6072), .A1(P2_IR_REG_23__SCAN_IN), .B0(n6340), .Y(n6341));
  INVX1   g04755(.A(n6341), .Y(n6342));
  NOR2X1  g04756(.A(P2_IR_REG_31__SCAN_IN), .B(n6277), .Y(n6343));
  AOI21X1 g04757(.A0(n6291), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6343), .Y(n6344));
  NOR2X1  g04758(.A(P2_IR_REG_31__SCAN_IN), .B(n6286), .Y(n6345));
  AOI21X1 g04759(.A0(n6270), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6345), .Y(n6346));
  NOR2X1  g04760(.A(P2_IR_REG_31__SCAN_IN), .B(n6262), .Y(n6347));
  AOI21X1 g04761(.A0(n6263), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6347), .Y(n6348));
  NOR3X1  g04762(.A(n6348), .B(n6346), .C(n6344), .Y(n6349));
  NOR3X1  g04763(.A(n6349), .B(n6342), .C(P2_U3088), .Y(n6350));
  INVX1   g04764(.A(n6344), .Y(n6351));
  INVX1   g04765(.A(n6346), .Y(n6352));
  XOR2X1  g04766(.A(n6348), .B(P2_B_REG_SCAN_IN), .Y(n6353));
  OAI21X1 g04767(.A0(n6353), .A1(n6352), .B0(n6351), .Y(n6354));
  OAI21X1 g04768(.A0(n6352), .A1(n6344), .B0(n6348), .Y(n6355));
  NAND3X1 g04769(.A(n6355), .B(n6354), .C(n6350), .Y(n6356));
  INVX1   g04770(.A(n6350), .Y(n6357));
  INVX1   g04771(.A(n6354), .Y(n6358));
  OAI21X1 g04772(.A0(n6358), .A1(n6357), .B0(P2_D_REG_0__SCAN_IN), .Y(n6359));
  NAND2X1 g04773(.A(n6359), .B(n6356), .Y(P2_U3416));
  NAND2X1 g04774(.A(n6354), .B(n6350), .Y(n6361));
  NOR2X1  g04775(.A(n6352), .B(n6351), .Y(n6362));
  OAI21X1 g04776(.A0(n6358), .A1(n6357), .B0(P2_D_REG_1__SCAN_IN), .Y(n6363));
  OAI21X1 g04777(.A0(n6362), .A1(n6361), .B0(n6363), .Y(P2_U3417));
  INVX1   g04778(.A(P2_D_REG_2__SCAN_IN), .Y(n6365));
  AOI21X1 g04779(.A0(n6354), .A1(n6350), .B0(n6365), .Y(P2_U3295));
  INVX1   g04780(.A(P2_D_REG_3__SCAN_IN), .Y(n6367));
  AOI21X1 g04781(.A0(n6354), .A1(n6350), .B0(n6367), .Y(P2_U3294));
  INVX1   g04782(.A(P2_D_REG_4__SCAN_IN), .Y(n6369));
  AOI21X1 g04783(.A0(n6354), .A1(n6350), .B0(n6369), .Y(P2_U3293));
  INVX1   g04784(.A(P2_D_REG_5__SCAN_IN), .Y(n6371));
  AOI21X1 g04785(.A0(n6354), .A1(n6350), .B0(n6371), .Y(P2_U3292));
  INVX1   g04786(.A(P2_D_REG_6__SCAN_IN), .Y(n6373));
  AOI21X1 g04787(.A0(n6354), .A1(n6350), .B0(n6373), .Y(P2_U3291));
  INVX1   g04788(.A(P2_D_REG_7__SCAN_IN), .Y(n6375));
  AOI21X1 g04789(.A0(n6354), .A1(n6350), .B0(n6375), .Y(P2_U3290));
  INVX1   g04790(.A(P2_D_REG_8__SCAN_IN), .Y(n6377));
  AOI21X1 g04791(.A0(n6354), .A1(n6350), .B0(n6377), .Y(P2_U3289));
  INVX1   g04792(.A(P2_D_REG_9__SCAN_IN), .Y(n6379));
  AOI21X1 g04793(.A0(n6354), .A1(n6350), .B0(n6379), .Y(P2_U3288));
  INVX1   g04794(.A(P2_D_REG_10__SCAN_IN), .Y(n6381));
  AOI21X1 g04795(.A0(n6354), .A1(n6350), .B0(n6381), .Y(P2_U3287));
  INVX1   g04796(.A(P2_D_REG_11__SCAN_IN), .Y(n6383));
  AOI21X1 g04797(.A0(n6354), .A1(n6350), .B0(n6383), .Y(P2_U3286));
  INVX1   g04798(.A(P2_D_REG_12__SCAN_IN), .Y(n6385));
  AOI21X1 g04799(.A0(n6354), .A1(n6350), .B0(n6385), .Y(P2_U3285));
  INVX1   g04800(.A(P2_D_REG_13__SCAN_IN), .Y(n6387));
  AOI21X1 g04801(.A0(n6354), .A1(n6350), .B0(n6387), .Y(P2_U3284));
  INVX1   g04802(.A(P2_D_REG_14__SCAN_IN), .Y(n6389));
  AOI21X1 g04803(.A0(n6354), .A1(n6350), .B0(n6389), .Y(P2_U3283));
  INVX1   g04804(.A(P2_D_REG_15__SCAN_IN), .Y(n6391));
  AOI21X1 g04805(.A0(n6354), .A1(n6350), .B0(n6391), .Y(P2_U3282));
  INVX1   g04806(.A(P2_D_REG_16__SCAN_IN), .Y(n6393));
  AOI21X1 g04807(.A0(n6354), .A1(n6350), .B0(n6393), .Y(P2_U3281));
  INVX1   g04808(.A(P2_D_REG_17__SCAN_IN), .Y(n6395));
  AOI21X1 g04809(.A0(n6354), .A1(n6350), .B0(n6395), .Y(P2_U3280));
  INVX1   g04810(.A(P2_D_REG_18__SCAN_IN), .Y(n6397));
  AOI21X1 g04811(.A0(n6354), .A1(n6350), .B0(n6397), .Y(P2_U3279));
  INVX1   g04812(.A(P2_D_REG_19__SCAN_IN), .Y(n6399));
  AOI21X1 g04813(.A0(n6354), .A1(n6350), .B0(n6399), .Y(P2_U3278));
  INVX1   g04814(.A(P2_D_REG_20__SCAN_IN), .Y(n6401));
  AOI21X1 g04815(.A0(n6354), .A1(n6350), .B0(n6401), .Y(P2_U3277));
  INVX1   g04816(.A(P2_D_REG_21__SCAN_IN), .Y(n6403));
  AOI21X1 g04817(.A0(n6354), .A1(n6350), .B0(n6403), .Y(P2_U3276));
  INVX1   g04818(.A(P2_D_REG_22__SCAN_IN), .Y(n6405));
  AOI21X1 g04819(.A0(n6354), .A1(n6350), .B0(n6405), .Y(P2_U3275));
  INVX1   g04820(.A(P2_D_REG_23__SCAN_IN), .Y(n6407));
  AOI21X1 g04821(.A0(n6354), .A1(n6350), .B0(n6407), .Y(P2_U3274));
  INVX1   g04822(.A(P2_D_REG_24__SCAN_IN), .Y(n6409));
  AOI21X1 g04823(.A0(n6354), .A1(n6350), .B0(n6409), .Y(P2_U3273));
  INVX1   g04824(.A(P2_D_REG_25__SCAN_IN), .Y(n6411));
  AOI21X1 g04825(.A0(n6354), .A1(n6350), .B0(n6411), .Y(P2_U3272));
  INVX1   g04826(.A(P2_D_REG_26__SCAN_IN), .Y(n6413));
  AOI21X1 g04827(.A0(n6354), .A1(n6350), .B0(n6413), .Y(P2_U3271));
  INVX1   g04828(.A(P2_D_REG_27__SCAN_IN), .Y(n6415));
  AOI21X1 g04829(.A0(n6354), .A1(n6350), .B0(n6415), .Y(P2_U3270));
  INVX1   g04830(.A(P2_D_REG_28__SCAN_IN), .Y(n6417));
  AOI21X1 g04831(.A0(n6354), .A1(n6350), .B0(n6417), .Y(P2_U3269));
  INVX1   g04832(.A(P2_D_REG_29__SCAN_IN), .Y(n6419));
  AOI21X1 g04833(.A0(n6354), .A1(n6350), .B0(n6419), .Y(P2_U3268));
  INVX1   g04834(.A(P2_D_REG_30__SCAN_IN), .Y(n6421));
  AOI21X1 g04835(.A0(n6354), .A1(n6350), .B0(n6421), .Y(P2_U3267));
  INVX1   g04836(.A(P2_D_REG_31__SCAN_IN), .Y(n6423));
  AOI21X1 g04837(.A0(n6354), .A1(n6350), .B0(n6423), .Y(P2_U3266));
  OAI21X1 g04838(.A0(P2_D_REG_7__SCAN_IN), .A1(P2_D_REG_3__SCAN_IN), .B0(n6358), .Y(n6425));
  OAI21X1 g04839(.A0(P2_D_REG_9__SCAN_IN), .A1(P2_D_REG_8__SCAN_IN), .B0(n6358), .Y(n6426));
  OAI21X1 g04840(.A0(P2_D_REG_10__SCAN_IN), .A1(P2_D_REG_5__SCAN_IN), .B0(n6358), .Y(n6427));
  OAI21X1 g04841(.A0(P2_D_REG_6__SCAN_IN), .A1(P2_D_REG_4__SCAN_IN), .B0(n6358), .Y(n6428));
  NAND4X1 g04842(.A(n6427), .B(n6426), .C(n6425), .D(n6428), .Y(n6429));
  OAI21X1 g04843(.A0(P2_D_REG_28__SCAN_IN), .A1(P2_D_REG_27__SCAN_IN), .B0(n6358), .Y(n6430));
  OAI21X1 g04844(.A0(P2_D_REG_26__SCAN_IN), .A1(P2_D_REG_25__SCAN_IN), .B0(n6358), .Y(n6431));
  OAI21X1 g04845(.A0(P2_D_REG_31__SCAN_IN), .A1(P2_D_REG_30__SCAN_IN), .B0(n6358), .Y(n6432));
  OAI21X1 g04846(.A0(P2_D_REG_29__SCAN_IN), .A1(P2_D_REG_2__SCAN_IN), .B0(n6358), .Y(n6433));
  NAND4X1 g04847(.A(n6432), .B(n6431), .C(n6430), .D(n6433), .Y(n6434));
  OAI21X1 g04848(.A0(P2_D_REG_21__SCAN_IN), .A1(P2_D_REG_20__SCAN_IN), .B0(n6358), .Y(n6435));
  OAI21X1 g04849(.A0(P2_D_REG_19__SCAN_IN), .A1(P2_D_REG_18__SCAN_IN), .B0(n6358), .Y(n6436));
  OAI21X1 g04850(.A0(P2_D_REG_23__SCAN_IN), .A1(P2_D_REG_22__SCAN_IN), .B0(n6358), .Y(n6437));
  AOI21X1 g04851(.A0(n6389), .A1(n6385), .B0(n6354), .Y(n6438));
  AOI21X1 g04852(.A0(n6387), .A1(n6383), .B0(n6354), .Y(n6439));
  AOI21X1 g04853(.A0(n6409), .A1(n6393), .B0(n6354), .Y(n6440));
  AOI21X1 g04854(.A0(n6395), .A1(n6391), .B0(n6354), .Y(n6441));
  NOR4X1  g04855(.A(n6440), .B(n6439), .C(n6438), .D(n6441), .Y(n6442));
  NAND4X1 g04856(.A(n6437), .B(n6436), .C(n6435), .D(n6442), .Y(n6443));
  NOR3X1  g04857(.A(n6443), .B(n6434), .C(n6429), .Y(n6444));
  NOR2X1  g04858(.A(n6362), .B(n6358), .Y(n6445));
  AOI21X1 g04859(.A0(n6358), .A1(P2_D_REG_1__SCAN_IN), .B0(n6445), .Y(n6446));
  INVX1   g04860(.A(n6446), .Y(n6447));
  NOR2X1  g04861(.A(P2_IR_REG_31__SCAN_IN), .B(n6245), .Y(n6448));
  AOI21X1 g04862(.A0(n6247), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6448), .Y(n6449));
  NOR2X1  g04863(.A(P2_IR_REG_31__SCAN_IN), .B(n6237), .Y(n6450));
  AOI21X1 g04864(.A0(n6231), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6450), .Y(n6451));
  INVX1   g04865(.A(n6451), .Y(n6452));
  INVX1   g04866(.A(P2_IR_REG_21__SCAN_IN), .Y(n6453));
  NOR2X1  g04867(.A(P2_IR_REG_31__SCAN_IN), .B(n6453), .Y(n6454));
  AOI21X1 g04868(.A0(n6239), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6454), .Y(n6455));
  INVX1   g04869(.A(n6455), .Y(n6456));
  OAI21X1 g04870(.A0(n6456), .A1(n6452), .B0(n6449), .Y(n6457));
  INVX1   g04871(.A(n6449), .Y(n6458));
  NOR2X1  g04872(.A(P2_IR_REG_31__SCAN_IN), .B(n6229), .Y(n6459));
  AOI21X1 g04873(.A0(n6222), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6459), .Y(n6460));
  AOI22X1 g04874(.A0(n6455), .A1(n6458), .B0(n6451), .B1(n6460), .Y(n6461));
  AOI21X1 g04875(.A0(n6461), .A1(n6457), .B0(n6447), .Y(n6462));
  AOI21X1 g04876(.A0(n6348), .A1(n6344), .B0(n6358), .Y(n6463));
  AOI21X1 g04877(.A0(n6358), .A1(P2_D_REG_0__SCAN_IN), .B0(n6463), .Y(n6464));
  NAND4X1 g04878(.A(n6462), .B(n6444), .C(n6350), .D(n6464), .Y(n6465));
  XOR2X1  g04879(.A(n6290), .B(P2_IR_REG_27__SCAN_IN), .Y(n6466));
  NOR2X1  g04880(.A(P2_IR_REG_31__SCAN_IN), .B(n6298), .Y(n6467));
  INVX1   g04881(.A(n6467), .Y(n6468));
  OAI21X1 g04882(.A0(n6466), .A1(n6072), .B0(n6468), .Y(n6469));
  XOR2X1  g04883(.A(n6308), .B(P2_IR_REG_28__SCAN_IN), .Y(n6470));
  NOR2X1  g04884(.A(P2_IR_REG_31__SCAN_IN), .B(n6305), .Y(n6471));
  INVX1   g04885(.A(n6471), .Y(n6472));
  OAI21X1 g04886(.A0(n6470), .A1(n6072), .B0(n6472), .Y(n6473));
  NOR2X1  g04887(.A(n6473), .B(n6469), .Y(n6474));
  INVX1   g04888(.A(P2_IR_REG_0__SCAN_IN), .Y(n6475));
  INVX1   g04889(.A(n6475), .Y(n6479));
  AOI21X1 g04890(.A0(n6299), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6467), .Y(n6480));
  AOI21X1 g04891(.A0(n6309), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6471), .Y(n6481));
  NAND3X1 g04892(.A(n6481), .B(n6480), .C(n6479), .Y(n6482));
  OAI21X1 g04893(.A0(n6474), .A1(n6065), .B0(n6482), .Y(n6483));
  INVX1   g04894(.A(P2_REG2_REG_0__SCAN_IN), .Y(n6484));
  INVX1   g04895(.A(P2_IR_REG_30__SCAN_IN), .Y(n6485));
  NAND2X1 g04896(.A(n6331), .B(P2_IR_REG_31__SCAN_IN), .Y(n6486));
  OAI21X1 g04897(.A0(P2_IR_REG_31__SCAN_IN), .A1(n6485), .B0(n6486), .Y(n6487));
  NAND2X1 g04898(.A(n6324), .B(P2_IR_REG_31__SCAN_IN), .Y(n6488));
  NAND2X1 g04899(.A(n6072), .B(P2_IR_REG_29__SCAN_IN), .Y(n6489));
  NAND3X1 g04900(.A(n6489), .B(n6488), .C(n6487), .Y(n6490));
  NOR2X1  g04901(.A(P2_IR_REG_31__SCAN_IN), .B(n6485), .Y(n6491));
  AOI21X1 g04902(.A0(n6331), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6491), .Y(n6492));
  NAND4X1 g04903(.A(n6488), .B(n6492), .C(P2_REG0_REG_0__SCAN_IN), .D(n6489), .Y(n6493));
  OAI21X1 g04904(.A0(n6490), .A1(n6484), .B0(n6493), .Y(n6494));
  INVX1   g04905(.A(P2_REG1_REG_0__SCAN_IN), .Y(n6495));
  INVX1   g04906(.A(P2_REG3_REG_0__SCAN_IN), .Y(n6496));
  NAND2X1 g04907(.A(n6322), .B(P2_IR_REG_29__SCAN_IN), .Y(n6497));
  NAND2X1 g04908(.A(n6330), .B(n6497), .Y(n6498));
  NOR2X1  g04909(.A(n6498), .B(n6072), .Y(n6499));
  INVX1   g04910(.A(n6489), .Y(n6500));
  OAI21X1 g04911(.A0(n6500), .A1(n6499), .B0(n6492), .Y(n6501));
  AOI21X1 g04912(.A0(n6489), .A1(n6488), .B0(n6492), .Y(n6502));
  INVX1   g04913(.A(n6502), .Y(n6503));
  OAI22X1 g04914(.A0(n6501), .A1(n6495), .B0(n6496), .B1(n6503), .Y(n6504));
  NOR2X1  g04915(.A(n6504), .B(n6494), .Y(n6505));
  XOR2X1  g04916(.A(n6505), .B(n6483), .Y(n6506));
  NOR3X1  g04917(.A(n6460), .B(n6451), .C(n6449), .Y(n6507));
  INVX1   g04918(.A(n6507), .Y(n6508));
  NOR2X1  g04919(.A(n6508), .B(n6506), .Y(n6509));
  INVX1   g04920(.A(n6509), .Y(n6510));
  NOR3X1  g04921(.A(n6460), .B(n6455), .C(n6451), .Y(n6512));
  INVX1   g04922(.A(n6460), .Y(n6513));
  NOR3X1  g04923(.A(n6513), .B(n6451), .C(n6449), .Y(n6514));
  OAI21X1 g04924(.A0(n6514), .A1(n6512), .B0(n9403), .Y(n6515));
  NOR3X1  g04925(.A(n6460), .B(n6452), .C(n6449), .Y(n6516));
  NAND2X1 g04926(.A(n6460), .B(n6451), .Y(n6517));
  NOR3X1  g04927(.A(n6517), .B(n6455), .C(n6458), .Y(n6518));
  OAI21X1 g04928(.A0(n6518), .A1(n6516), .B0(n9403), .Y(n6519));
  NOR4X1  g04929(.A(n6456), .B(n6452), .C(n6449), .D(n6513), .Y(n6520));
  NOR3X1  g04930(.A(n6513), .B(n6455), .C(n6451), .Y(n6521));
  OAI21X1 g04931(.A0(n6521), .A1(n6520), .B0(n9403), .Y(n6522));
  NAND4X1 g04932(.A(n6519), .B(n6515), .C(n6510), .D(n6522), .Y(n6523));
  NOR3X1  g04933(.A(n6460), .B(n6452), .C(n6458), .Y(n6524));
  INVX1   g04934(.A(n6524), .Y(n6525));
  NOR3X1  g04935(.A(n6460), .B(n6456), .C(n6458), .Y(n6526));
  NOR4X1  g04936(.A(n6456), .B(n6451), .C(n6458), .D(n6513), .Y(n6527));
  NOR2X1  g04937(.A(n6527), .B(n6526), .Y(n6528));
  INVX1   g04938(.A(n6528), .Y(n6529));
  AOI21X1 g04939(.A0(n6481), .A1(n6480), .B0(n6065), .Y(n6530));
  AOI21X1 g04940(.A0(n6474), .A1(n6479), .B0(n6530), .Y(n6531));
  NOR3X1  g04941(.A(n6456), .B(n6452), .C(n6458), .Y(n6532));
  INVX1   g04942(.A(n6532), .Y(n6533));
  NOR3X1  g04943(.A(n6473), .B(n6455), .C(n6449), .Y(n6534));
  INVX1   g04944(.A(n6534), .Y(n6535));
  INVX1   g04945(.A(P2_REG2_REG_1__SCAN_IN), .Y(n6536));
  NAND4X1 g04946(.A(n6488), .B(n6492), .C(P2_REG0_REG_1__SCAN_IN), .D(n6489), .Y(n6537));
  OAI21X1 g04947(.A0(n6490), .A1(n6536), .B0(n6537), .Y(n6538));
  INVX1   g04948(.A(P2_REG1_REG_1__SCAN_IN), .Y(n6539));
  INVX1   g04949(.A(P2_REG3_REG_1__SCAN_IN), .Y(n6540));
  OAI22X1 g04950(.A0(n6501), .A1(n6539), .B0(n6540), .B1(n6503), .Y(n6541));
  NOR2X1  g04951(.A(n6541), .B(n6538), .Y(n6542));
  OAI22X1 g04952(.A0(n6535), .A1(n6542), .B0(n6533), .B1(n6531), .Y(n6543));
  AOI21X1 g04953(.A0(n6529), .A1(n6483), .B0(n6543), .Y(n6544));
  OAI21X1 g04954(.A0(n6525), .A1(n6506), .B0(n6544), .Y(n6545));
  NOR2X1  g04955(.A(n6545), .B(n6523), .Y(n6546));
  NAND2X1 g04956(.A(n6465), .B(P2_REG0_REG_0__SCAN_IN), .Y(n6547));
  OAI21X1 g04957(.A0(n6546), .A1(n6465), .B0(n6547), .Y(P2_U3430));
  INVX1   g04958(.A(P2_IR_REG_1__SCAN_IN), .Y(n6549));
  NOR2X1  g04959(.A(P2_IR_REG_31__SCAN_IN), .B(n6549), .Y(n6550));
  AOI21X1 g04960(.A0(n6074), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6550), .Y(n6551));
  INVX1   g04961(.A(n6551), .Y(n6552));
  AOI21X1 g04962(.A0(n6481), .A1(n6480), .B0(n6071), .Y(n6553));
  AOI21X1 g04963(.A0(n6552), .A1(n6474), .B0(n6553), .Y(n6554));
  XOR2X1  g04964(.A(n6554), .B(n6542), .Y(n6555));
  NOR3X1  g04965(.A(n6500), .B(n6499), .C(n6492), .Y(n6556));
  NOR3X1  g04966(.A(n6500), .B(n6499), .C(n6487), .Y(n6557));
  AOI22X1 g04967(.A0(n6556), .A1(P2_REG2_REG_0__SCAN_IN), .B0(P2_REG0_REG_0__SCAN_IN), .B1(n6557), .Y(n6558));
  AOI21X1 g04968(.A0(n6489), .A1(n6488), .B0(n6487), .Y(n6559));
  AOI22X1 g04969(.A0(n6559), .A1(P2_REG1_REG_0__SCAN_IN), .B0(P2_REG3_REG_0__SCAN_IN), .B1(n6502), .Y(n6560));
  AOI21X1 g04970(.A0(n6560), .A1(n6558), .B0(n6531), .Y(n6561));
  INVX1   g04971(.A(n6561), .Y(n6562));
  XOR2X1  g04972(.A(n6562), .B(n6555), .Y(n6563));
  INVX1   g04973(.A(n6563), .Y(n6564));
  OAI21X1 g04974(.A0(n6520), .A1(n6514), .B0(n6564), .Y(n6565));
  NAND3X1 g04975(.A(n6560), .B(n6558), .C(n6483), .Y(n6566));
  AOI22X1 g04976(.A0(n6556), .A1(P2_REG2_REG_1__SCAN_IN), .B0(P2_REG0_REG_1__SCAN_IN), .B1(n6557), .Y(n6567));
  AOI22X1 g04977(.A0(n6559), .A1(P2_REG1_REG_1__SCAN_IN), .B0(P2_REG3_REG_1__SCAN_IN), .B1(n6502), .Y(n6568));
  NAND2X1 g04978(.A(n6568), .B(n6567), .Y(n6569));
  XOR2X1  g04979(.A(n6554), .B(n6569), .Y(n6570));
  XOR2X1  g04980(.A(n6570), .B(n6566), .Y(n6571));
  AOI22X1 g04981(.A0(n6564), .A1(n6518), .B0(n6512), .B1(n6571), .Y(n6572));
  INVX1   g04982(.A(n6505), .Y(n6573));
  NOR3X1  g04983(.A(n6481), .B(n6455), .C(n6449), .Y(n6574));
  AOI22X1 g04984(.A0(n6571), .A1(n6521), .B0(n6573), .B1(n6574), .Y(n6575));
  OAI21X1 g04985(.A0(n6516), .A1(n6507), .B0(n6571), .Y(n6576));
  NAND4X1 g04986(.A(n6575), .B(n6572), .C(n6565), .D(n6576), .Y(n6577));
  NOR2X1  g04987(.A(n6563), .B(n6525), .Y(n6578));
  XOR2X1  g04988(.A(n6554), .B(n6483), .Y(n6579));
  INVX1   g04989(.A(n6554), .Y(n6580));
  AOI22X1 g04990(.A0(n6556), .A1(P2_REG2_REG_2__SCAN_IN), .B0(P2_REG0_REG_2__SCAN_IN), .B1(n6557), .Y(n6581));
  AOI22X1 g04991(.A0(n6559), .A1(P2_REG1_REG_2__SCAN_IN), .B0(P2_REG3_REG_2__SCAN_IN), .B1(n6502), .Y(n6582));
  NAND2X1 g04992(.A(n6582), .B(n6581), .Y(n6583));
  AOI22X1 g04993(.A0(n6580), .A1(n6529), .B0(n6534), .B1(n6583), .Y(n6584));
  OAI21X1 g04994(.A0(n6579), .A1(n6533), .B0(n6584), .Y(n6585));
  NOR3X1  g04995(.A(n6585), .B(n6578), .C(n6577), .Y(n6586));
  NAND2X1 g04996(.A(n6465), .B(P2_REG0_REG_1__SCAN_IN), .Y(n6587));
  OAI21X1 g04997(.A0(n6586), .A1(n6465), .B0(n6587), .Y(P2_U3433));
  INVX1   g04998(.A(P2_REG2_REG_2__SCAN_IN), .Y(n6589));
  NAND4X1 g04999(.A(n6488), .B(n6492), .C(P2_REG0_REG_2__SCAN_IN), .D(n6489), .Y(n6590));
  OAI21X1 g05000(.A0(n6490), .A1(n6589), .B0(n6590), .Y(n6591));
  INVX1   g05001(.A(P2_REG1_REG_2__SCAN_IN), .Y(n6592));
  INVX1   g05002(.A(P2_REG3_REG_2__SCAN_IN), .Y(n6593));
  OAI22X1 g05003(.A0(n6501), .A1(n6592), .B0(n6593), .B1(n6503), .Y(n6594));
  NOR2X1  g05004(.A(n6594), .B(n6591), .Y(n6595));
  NOR2X1  g05005(.A(P2_IR_REG_31__SCAN_IN), .B(n6079), .Y(n6596));
  AOI21X1 g05006(.A0(n6081), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6596), .Y(n6597));
  INVX1   g05007(.A(n6597), .Y(n6598));
  NAND3X1 g05008(.A(n6598), .B(n6481), .C(n6480), .Y(n6599));
  OAI21X1 g05009(.A0(n6474), .A1(n6078), .B0(n6599), .Y(n6600));
  INVX1   g05010(.A(n6600), .Y(n6601));
  XOR2X1  g05011(.A(n6601), .B(n6595), .Y(n6602));
  OAI21X1 g05012(.A0(n6580), .A1(n6569), .B0(n6561), .Y(n6603));
  OAI21X1 g05013(.A0(n6554), .A1(n6542), .B0(n6603), .Y(n6604));
  XOR2X1  g05014(.A(n6600), .B(n6595), .Y(n6605));
  NOR2X1  g05015(.A(n6602), .B(n6604), .Y(n6607));
  AOI21X1 g05016(.A0(n6604), .A1(n6602), .B0(n6607), .Y(n6608));
  AOI22X1 g05017(.A0(n6574), .A1(n6569), .B0(n6518), .B1(n6608), .Y(n6609));
  OAI21X1 g05018(.A0(n6520), .A1(n6514), .B0(n6608), .Y(n6610));
  NAND2X1 g05019(.A(n6569), .B(n6566), .Y(n6611));
  OAI21X1 g05020(.A0(n6569), .A1(n6566), .B0(n6554), .Y(n6612));
  NAND2X1 g05021(.A(n6612), .B(n6611), .Y(n6613));
  XOR2X1  g05022(.A(n6613), .B(n6605), .Y(n6614));
  OAI21X1 g05023(.A0(n6521), .A1(n6507), .B0(n6614), .Y(n6615));
  OAI21X1 g05024(.A0(n6516), .A1(n6512), .B0(n6614), .Y(n6616));
  NAND4X1 g05025(.A(n6615), .B(n6610), .C(n6609), .D(n6616), .Y(n6617));
  NAND2X1 g05026(.A(n6608), .B(n6524), .Y(n6618));
  NAND2X1 g05027(.A(n6554), .B(n6531), .Y(n6619));
  XOR2X1  g05028(.A(n6619), .B(n6600), .Y(n6620));
  INVX1   g05029(.A(P2_REG2_REG_3__SCAN_IN), .Y(n6621));
  NAND4X1 g05030(.A(n6488), .B(n6492), .C(P2_REG0_REG_3__SCAN_IN), .D(n6489), .Y(n6622));
  OAI21X1 g05031(.A0(n6490), .A1(n6621), .B0(n6622), .Y(n6623));
  INVX1   g05032(.A(P2_REG1_REG_3__SCAN_IN), .Y(n6624));
  OAI22X1 g05033(.A0(n6501), .A1(n6624), .B0(P2_REG3_REG_3__SCAN_IN), .B1(n6503), .Y(n6625));
  NOR2X1  g05034(.A(n6625), .B(n6623), .Y(n6626));
  OAI22X1 g05035(.A0(n6601), .A1(n6528), .B0(n6535), .B1(n6626), .Y(n6627));
  AOI21X1 g05036(.A0(n6620), .A1(n6532), .B0(n6627), .Y(n6628));
  NAND2X1 g05037(.A(n6628), .B(n6618), .Y(n6629));
  NOR2X1  g05038(.A(n6629), .B(n6617), .Y(n6630));
  NAND2X1 g05039(.A(n6465), .B(P2_REG0_REG_2__SCAN_IN), .Y(n6631));
  OAI21X1 g05040(.A0(n6630), .A1(n6465), .B0(n6631), .Y(P2_U3436));
  INVX1   g05041(.A(n6518), .Y(n6633));
  INVX1   g05042(.A(n6574), .Y(n6634));
  NAND2X1 g05043(.A(n6601), .B(n6595), .Y(n6635));
  INVX1   g05044(.A(n6603), .Y(n6636));
  AOI21X1 g05045(.A0(n6568), .A1(n6567), .B0(n6554), .Y(n6637));
  NOR2X1  g05046(.A(n6601), .B(n6595), .Y(n6638));
  AOI21X1 g05047(.A0(n6635), .A1(n6637), .B0(n6638), .Y(n6639));
  INVX1   g05048(.A(n6639), .Y(n6640));
  AOI21X1 g05049(.A0(n6636), .A1(n6635), .B0(n6640), .Y(n6641));
  NOR2X1  g05050(.A(P2_IR_REG_31__SCAN_IN), .B(n6086), .Y(n6642));
  AOI21X1 g05051(.A0(n6088), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6642), .Y(n6643));
  INVX1   g05052(.A(n6643), .Y(n6644));
  NAND3X1 g05053(.A(n6644), .B(n6481), .C(n6480), .Y(n6645));
  OAI21X1 g05054(.A0(n6474), .A1(n6085), .B0(n6645), .Y(n6646));
  XOR2X1  g05055(.A(n6646), .B(n6626), .Y(n6647));
  AOI22X1 g05056(.A0(n6556), .A1(P2_REG2_REG_3__SCAN_IN), .B0(P2_REG0_REG_3__SCAN_IN), .B1(n6557), .Y(n6649));
  INVX1   g05057(.A(P2_REG3_REG_3__SCAN_IN), .Y(n6650));
  AOI22X1 g05058(.A0(n6559), .A1(P2_REG1_REG_3__SCAN_IN), .B0(n6650), .B1(n6502), .Y(n6651));
  NAND2X1 g05059(.A(n6651), .B(n6649), .Y(n6652));
  XOR2X1  g05060(.A(n6646), .B(n6652), .Y(n6653));
  NOR2X1  g05061(.A(n6653), .B(n6641), .Y(n6654));
  AOI21X1 g05062(.A0(n6653), .A1(n6641), .B0(n6654), .Y(n6655));
  OAI22X1 g05063(.A0(n6595), .A1(n6634), .B0(n6633), .B1(n6655), .Y(n6656));
  INVX1   g05064(.A(n6514), .Y(n6657));
  INVX1   g05065(.A(n6520), .Y(n6658));
  AOI21X1 g05066(.A0(n6658), .A1(n6657), .B0(n6655), .Y(n6659));
  NOR2X1  g05067(.A(n6659), .B(n6656), .Y(n6660));
  INVX1   g05068(.A(n6521), .Y(n6661));
  AOI21X1 g05069(.A0(n6582), .A1(n6581), .B0(n6600), .Y(n6662));
  AOI21X1 g05070(.A0(n6600), .A1(n6595), .B0(n6647), .Y(n6663));
  OAI21X1 g05071(.A0(n6613), .A1(n6662), .B0(n6663), .Y(n6664));
  INVX1   g05072(.A(n6662), .Y(n6665));
  OAI21X1 g05073(.A0(n6601), .A1(n6583), .B0(n6613), .Y(n6666));
  NAND3X1 g05074(.A(n6666), .B(n6647), .C(n6665), .Y(n6667));
  AOI22X1 g05075(.A0(n6664), .A1(n6667), .B0(n6661), .B1(n6508), .Y(n6668));
  INVX1   g05076(.A(n6512), .Y(n6669));
  INVX1   g05077(.A(n6516), .Y(n6670));
  AOI22X1 g05078(.A0(n6664), .A1(n6667), .B0(n6670), .B1(n6669), .Y(n6671));
  NOR2X1  g05079(.A(n6671), .B(n6668), .Y(n6672));
  NAND2X1 g05080(.A(n6672), .B(n6660), .Y(n6673));
  NAND3X1 g05081(.A(n6601), .B(n6554), .C(n6531), .Y(n6674));
  XOR2X1  g05082(.A(n6646), .B(n6674), .Y(n6675));
  NOR2X1  g05083(.A(n6474), .B(n6085), .Y(n6676));
  AOI21X1 g05084(.A0(n6644), .A1(n6474), .B0(n6676), .Y(n6677));
  INVX1   g05085(.A(P2_REG2_REG_4__SCAN_IN), .Y(n6678));
  NAND4X1 g05086(.A(n6488), .B(n6492), .C(P2_REG0_REG_4__SCAN_IN), .D(n6489), .Y(n6679));
  OAI21X1 g05087(.A0(n6490), .A1(n6678), .B0(n6679), .Y(n6680));
  INVX1   g05088(.A(P2_REG1_REG_4__SCAN_IN), .Y(n6681));
  INVX1   g05089(.A(P2_REG3_REG_4__SCAN_IN), .Y(n6682));
  XOR2X1  g05090(.A(P2_REG3_REG_3__SCAN_IN), .B(n6682), .Y(n6683));
  OAI22X1 g05091(.A0(n6503), .A1(n6683), .B0(n6501), .B1(n6681), .Y(n6684));
  NOR2X1  g05092(.A(n6684), .B(n6680), .Y(n6685));
  OAI22X1 g05093(.A0(n6677), .A1(n6528), .B0(n6535), .B1(n6685), .Y(n6686));
  AOI21X1 g05094(.A0(n6675), .A1(n6532), .B0(n6686), .Y(n6687));
  OAI21X1 g05095(.A0(n6655), .A1(n6525), .B0(n6687), .Y(n6688));
  NOR2X1  g05096(.A(n6688), .B(n6673), .Y(n6689));
  NAND2X1 g05097(.A(n6465), .B(P2_REG0_REG_3__SCAN_IN), .Y(n6690));
  OAI21X1 g05098(.A0(n6689), .A1(n6465), .B0(n6690), .Y(P2_U3439));
  NOR2X1  g05099(.A(n6646), .B(n6652), .Y(n6692));
  NOR2X1  g05100(.A(P2_IR_REG_31__SCAN_IN), .B(n6093), .Y(n6699));
  INVX1   g05101(.A(n6699), .Y(n6700));
  OAI21X1 g05102(.A0(n6098), .A1(n6072), .B0(n6700), .Y(n6701));
  NAND3X1 g05103(.A(n6701), .B(n6481), .C(n6480), .Y(n6702));
  OAI21X1 g05104(.A0(n6474), .A1(n6092), .B0(n6702), .Y(n6703));
  XOR2X1  g05105(.A(n6703), .B(n6685), .Y(n6704));
  NOR2X1  g05106(.A(n6805), .B(n6704), .Y(n6705));
  INVX1   g05107(.A(n6685), .Y(n6706));
  AOI21X1 g05108(.A0(n6704), .A1(n6805), .B0(n6705), .Y(n6709));
  INVX1   g05109(.A(n6709), .Y(n6710));
  OAI21X1 g05110(.A0(n6520), .A1(n6514), .B0(n6710), .Y(n6711));
  AOI22X1 g05111(.A0(n6626), .A1(n6646), .B0(n6600), .B1(n6595), .Y(n6712));
  NAND2X1 g05112(.A(n6712), .B(n6613), .Y(n6713));
  OAI21X1 g05113(.A0(n6652), .A1(n6662), .B0(n6677), .Y(n6714));
  NAND2X1 g05114(.A(n6652), .B(n6662), .Y(n6715));
  NAND3X1 g05115(.A(n6715), .B(n6714), .C(n6713), .Y(n6716));
  XOR2X1  g05116(.A(n6716), .B(n6704), .Y(n6717));
  AOI22X1 g05117(.A0(n6710), .A1(n6518), .B0(n6512), .B1(n6717), .Y(n6718));
  AOI22X1 g05118(.A0(n6652), .A1(n6574), .B0(n6521), .B1(n6717), .Y(n6719));
  OAI21X1 g05119(.A0(n6516), .A1(n6507), .B0(n6717), .Y(n6720));
  NAND4X1 g05120(.A(n6719), .B(n6718), .C(n6711), .D(n6720), .Y(n6721));
  NOR3X1  g05121(.A(n6646), .B(n6619), .C(n6600), .Y(n6722));
  INVX1   g05122(.A(n6703), .Y(n6723));
  XOR2X1  g05123(.A(n6723), .B(n6722), .Y(n6724));
  INVX1   g05124(.A(P2_REG2_REG_5__SCAN_IN), .Y(n6725));
  NAND4X1 g05125(.A(n6488), .B(n6492), .C(P2_REG0_REG_5__SCAN_IN), .D(n6489), .Y(n6726));
  OAI21X1 g05126(.A0(n6490), .A1(n6725), .B0(n6726), .Y(n6727));
  INVX1   g05127(.A(P2_REG1_REG_5__SCAN_IN), .Y(n6728));
  NAND2X1 g05128(.A(P2_REG3_REG_3__SCAN_IN), .B(P2_REG3_REG_4__SCAN_IN), .Y(n6729));
  XOR2X1  g05129(.A(n6729), .B(P2_REG3_REG_5__SCAN_IN), .Y(n6730));
  OAI22X1 g05130(.A0(n6503), .A1(n6730), .B0(n6501), .B1(n6728), .Y(n6731));
  NOR2X1  g05131(.A(n6731), .B(n6727), .Y(n6732));
  OAI22X1 g05132(.A0(n6723), .A1(n6528), .B0(n6535), .B1(n6732), .Y(n6733));
  AOI21X1 g05133(.A0(n6724), .A1(n6532), .B0(n6733), .Y(n6734));
  OAI21X1 g05134(.A0(n6709), .A1(n6525), .B0(n6734), .Y(n6735));
  NOR2X1  g05135(.A(n6735), .B(n6721), .Y(n6736));
  NAND2X1 g05136(.A(n6465), .B(P2_REG0_REG_4__SCAN_IN), .Y(n6737));
  OAI21X1 g05137(.A0(n6736), .A1(n6465), .B0(n6737), .Y(P2_U3442));
  NOR2X1  g05138(.A(n6723), .B(n6685), .Y(n6739));
  NOR2X1  g05139(.A(n6739), .B(n6805), .Y(n6740));
  INVX1   g05140(.A(n6740), .Y(n6741));
  AOI22X1 g05141(.A0(n6556), .A1(P2_REG2_REG_5__SCAN_IN), .B0(P2_REG0_REG_5__SCAN_IN), .B1(n6557), .Y(n6742));
  INVX1   g05142(.A(n6730), .Y(n6743));
  AOI22X1 g05143(.A0(n6502), .A1(n6743), .B0(n6559), .B1(P2_REG1_REG_5__SCAN_IN), .Y(n6744));
  NAND2X1 g05144(.A(n6744), .B(n6742), .Y(n6745));
  NOR2X1  g05145(.A(P2_IR_REG_31__SCAN_IN), .B(n6105), .Y(n6746));
  AOI21X1 g05146(.A0(n6106), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6746), .Y(n6747));
  NOR3X1  g05147(.A(n6747), .B(n6473), .C(n6469), .Y(n6748));
  INVX1   g05148(.A(n6748), .Y(n6749));
  NAND2X1 g05149(.A(n6481), .B(n6480), .Y(n6750));
  OAI21X1 g05150(.A0(n6103), .A1(n6102), .B0(n6750), .Y(n6751));
  NAND2X1 g05151(.A(n6751), .B(n6749), .Y(n6752));
  INVX1   g05152(.A(n6752), .Y(n6753));
  AOI22X1 g05153(.A0(n6732), .A1(n6753), .B0(n6723), .B1(n6685), .Y(n6754));
  INVX1   g05154(.A(n6754), .Y(n6755));
  AOI21X1 g05155(.A0(n6752), .A1(n6745), .B0(n6755), .Y(n6756));
  OAI21X1 g05156(.A0(n6703), .A1(n6706), .B0(n6805), .Y(n6757));
  AOI21X1 g05157(.A0(n6751), .A1(n6749), .B0(n6745), .Y(n6758));
  NOR2X1  g05158(.A(n6752), .B(n6732), .Y(n6759));
  NOR3X1  g05159(.A(n6759), .B(n6758), .C(n6739), .Y(n6760));
  AOI22X1 g05160(.A0(n6757), .A1(n6760), .B0(n6756), .B1(n6741), .Y(n6761));
  AOI22X1 g05161(.A0(n6706), .A1(n6574), .B0(n6518), .B1(n6761), .Y(n6762));
  OAI21X1 g05162(.A0(n6520), .A1(n6514), .B0(n6761), .Y(n6763));
  XOR2X1  g05163(.A(n6752), .B(n6732), .Y(n6764));
  NOR2X1  g05164(.A(n6723), .B(n6706), .Y(n6765));
  INVX1   g05165(.A(n6765), .Y(n6766));
  NOR2X1  g05166(.A(n6703), .B(n6685), .Y(n6767));
  AOI21X1 g05167(.A0(n6716), .A1(n6766), .B0(n6767), .Y(n6768));
  XOR2X1  g05168(.A(n6768), .B(n6764), .Y(n6769));
  INVX1   g05169(.A(n6769), .Y(n6770));
  OAI21X1 g05170(.A0(n6521), .A1(n6507), .B0(n6770), .Y(n6771));
  OAI21X1 g05171(.A0(n6516), .A1(n6512), .B0(n6770), .Y(n6772));
  NAND4X1 g05172(.A(n6771), .B(n6763), .C(n6762), .D(n6772), .Y(n6773));
  NAND2X1 g05173(.A(n6761), .B(n6524), .Y(n6774));
  NAND2X1 g05174(.A(n6723), .B(n6722), .Y(n6775));
  XOR2X1  g05175(.A(n6752), .B(n6775), .Y(n6776));
  INVX1   g05176(.A(P2_REG2_REG_6__SCAN_IN), .Y(n6777));
  NAND4X1 g05177(.A(n6488), .B(n6492), .C(P2_REG0_REG_6__SCAN_IN), .D(n6489), .Y(n6778));
  OAI21X1 g05178(.A0(n6490), .A1(n6777), .B0(n6778), .Y(n6779));
  INVX1   g05179(.A(P2_REG1_REG_6__SCAN_IN), .Y(n6780));
  INVX1   g05180(.A(P2_REG3_REG_6__SCAN_IN), .Y(n6781));
  INVX1   g05181(.A(P2_REG3_REG_5__SCAN_IN), .Y(n6782));
  NOR2X1  g05182(.A(n6729), .B(n6782), .Y(n6783));
  XOR2X1  g05183(.A(n6783), .B(n6781), .Y(n6784));
  OAI22X1 g05184(.A0(n6503), .A1(n6784), .B0(n6501), .B1(n6780), .Y(n6785));
  NOR2X1  g05185(.A(n6785), .B(n6779), .Y(n6786));
  OAI22X1 g05186(.A0(n6753), .A1(n6528), .B0(n6535), .B1(n6786), .Y(n6787));
  AOI21X1 g05187(.A0(n6776), .A1(n6532), .B0(n6787), .Y(n6788));
  NAND2X1 g05188(.A(n6788), .B(n6774), .Y(n6789));
  NOR2X1  g05189(.A(n6789), .B(n6773), .Y(n6790));
  NAND2X1 g05190(.A(n6465), .B(P2_REG0_REG_5__SCAN_IN), .Y(n6791));
  OAI21X1 g05191(.A0(n6790), .A1(n6465), .B0(n6791), .Y(P2_U3445));
  NOR2X1  g05192(.A(P2_IR_REG_31__SCAN_IN), .B(n6111), .Y(n6793));
  AOI21X1 g05193(.A0(n6114), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6793), .Y(n6794));
  INVX1   g05194(.A(n6794), .Y(n6795));
  NAND2X1 g05195(.A(n6795), .B(n6474), .Y(n6796));
  OAI21X1 g05196(.A0(n6474), .A1(n6110), .B0(n6796), .Y(n6797));
  XOR2X1  g05197(.A(n6797), .B(n6786), .Y(n6798));
  NAND3X1 g05198(.A(n6752), .B(n6703), .C(n6706), .Y(n6800));
  OAI21X1 g05199(.A0(n6752), .A1(n6739), .B0(n6745), .Y(n6801));
  NAND2X1 g05200(.A(n6801), .B(n6800), .Y(n6802));
  NAND2X1 g05201(.A(n6604), .B(n6635), .Y(n6803));
  AOI22X1 g05202(.A0(n6652), .A1(n6646), .B0(n6600), .B1(n6583), .Y(n6804));
  AOI21X1 g05203(.A0(n6804), .A1(n6803), .B0(n6692), .Y(n6805));
  AOI21X1 g05204(.A0(n6805), .A1(n6754), .B0(n6802), .Y(n6806));
  INVX1   g05205(.A(n6786), .Y(n6807));
  XOR2X1  g05206(.A(n6797), .B(n6807), .Y(n6808));
  NOR2X1  g05207(.A(n6808), .B(n6806), .Y(n6809));
  AOI21X1 g05208(.A0(n6806), .A1(n6808), .B0(n6809), .Y(n6810));
  INVX1   g05209(.A(n6810), .Y(n6811));
  AOI22X1 g05210(.A0(n6745), .A1(n6574), .B0(n6518), .B1(n6811), .Y(n6812));
  OAI21X1 g05211(.A0(n6520), .A1(n6514), .B0(n6811), .Y(n6813));
  INVX1   g05212(.A(n6768), .Y(n6814));
  NOR2X1  g05213(.A(n6798), .B(n6758), .Y(n6815));
  OAI21X1 g05214(.A0(n6814), .A1(n6759), .B0(n6815), .Y(n6816));
  OAI22X1 g05215(.A0(n6786), .A1(n6797), .B0(n6752), .B1(n6732), .Y(n6817));
  AOI21X1 g05216(.A0(n6797), .A1(n6786), .B0(n6817), .Y(n6818));
  OAI21X1 g05217(.A0(n6768), .A1(n6758), .B0(n6818), .Y(n6819));
  NAND2X1 g05218(.A(n6819), .B(n6816), .Y(n6820));
  OAI21X1 g05219(.A0(n6521), .A1(n6507), .B0(n6820), .Y(n6821));
  OAI21X1 g05220(.A0(n6516), .A1(n6512), .B0(n6820), .Y(n6822));
  NAND4X1 g05221(.A(n6821), .B(n6813), .C(n6812), .D(n6822), .Y(n6823));
  NOR4X1  g05222(.A(n6703), .B(n6646), .C(n6674), .D(n6752), .Y(n6830));
  NOR2X1  g05223(.A(n6474), .B(n6110), .Y(n6831));
  AOI21X1 g05224(.A0(n6795), .A1(n6474), .B0(n6831), .Y(n6832));
  XOR2X1  g05225(.A(n6832), .B(n6830), .Y(n6833));
  AOI22X1 g05226(.A0(n6556), .A1(P2_REG2_REG_7__SCAN_IN), .B0(P2_REG0_REG_7__SCAN_IN), .B1(n6557), .Y(n6834));
  NAND4X1 g05227(.A(P2_REG3_REG_5__SCAN_IN), .B(P2_REG3_REG_4__SCAN_IN), .C(P2_REG3_REG_6__SCAN_IN), .D(P2_REG3_REG_3__SCAN_IN), .Y(n6835));
  XOR2X1  g05228(.A(n6835), .B(P2_REG3_REG_7__SCAN_IN), .Y(n6836));
  INVX1   g05229(.A(n6836), .Y(n6837));
  AOI22X1 g05230(.A0(n6502), .A1(n6837), .B0(n6559), .B1(P2_REG1_REG_7__SCAN_IN), .Y(n6838));
  NAND2X1 g05231(.A(n6838), .B(n6834), .Y(n6839));
  INVX1   g05232(.A(n6839), .Y(n6840));
  OAI22X1 g05233(.A0(n6832), .A1(n6528), .B0(n6535), .B1(n6840), .Y(n6841));
  AOI21X1 g05234(.A0(n6833), .A1(n6532), .B0(n6841), .Y(n6842));
  OAI21X1 g05235(.A0(n6810), .A1(n6525), .B0(n6842), .Y(n6843));
  NOR2X1  g05236(.A(n6843), .B(n6823), .Y(n6844));
  NAND2X1 g05237(.A(n6465), .B(P2_REG0_REG_6__SCAN_IN), .Y(n6845));
  OAI21X1 g05238(.A0(n6844), .A1(n6465), .B0(n6845), .Y(P2_U3448));
  NOR2X1  g05239(.A(P2_IR_REG_31__SCAN_IN), .B(n6119), .Y(n6847));
  AOI21X1 g05240(.A0(n6120), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6847), .Y(n6848));
  INVX1   g05241(.A(n6848), .Y(n6849));
  NAND2X1 g05242(.A(n6849), .B(n6474), .Y(n6850));
  OAI21X1 g05243(.A0(n6474), .A1(n6118), .B0(n6850), .Y(n6851));
  OAI22X1 g05244(.A0(n6839), .A1(n6851), .B0(n6797), .B1(n6807), .Y(n6852));
  AOI21X1 g05245(.A0(n6851), .A1(n6839), .B0(n6852), .Y(n6853));
  INVX1   g05246(.A(n6853), .Y(n6854));
  INVX1   g05247(.A(n6806), .Y(n6855));
  NAND2X1 g05248(.A(n6797), .B(n6807), .Y(n6856));
  INVX1   g05249(.A(n6856), .Y(n6857));
  NOR2X1  g05250(.A(n6857), .B(n6855), .Y(n6858));
  XOR2X1  g05251(.A(n6851), .B(n6840), .Y(n6859));
  INVX1   g05252(.A(n6859), .Y(n6860));
  NOR2X1  g05253(.A(n6860), .B(n6857), .Y(n6861));
  INVX1   g05254(.A(n6861), .Y(n6862));
  AOI21X1 g05255(.A0(n6832), .A1(n6786), .B0(n6806), .Y(n6863));
  OAI22X1 g05256(.A0(n6862), .A1(n6863), .B0(n6858), .B1(n6854), .Y(n6864));
  INVX1   g05257(.A(n6864), .Y(n6865));
  OAI21X1 g05258(.A0(n6520), .A1(n6514), .B0(n6865), .Y(n6866));
  INVX1   g05259(.A(n6866), .Y(n6867));
  NOR2X1  g05260(.A(n6832), .B(n6807), .Y(n6868));
  NOR3X1  g05261(.A(n6758), .B(n6703), .C(n6685), .Y(n6869));
  NOR2X1  g05262(.A(n6869), .B(n6817), .Y(n6870));
  NOR2X1  g05263(.A(n6870), .B(n6868), .Y(n6871));
  NOR3X1  g05264(.A(n6868), .B(n6758), .C(n6765), .Y(n6872));
  AOI21X1 g05265(.A0(n6872), .A1(n6716), .B0(n6871), .Y(n6873));
  XOR2X1  g05266(.A(n6873), .B(n6859), .Y(n6874));
  OAI22X1 g05267(.A0(n6864), .A1(n6633), .B0(n6669), .B1(n6874), .Y(n6875));
  OAI22X1 g05268(.A0(n6786), .A1(n6634), .B0(n6661), .B1(n6874), .Y(n6876));
  AOI21X1 g05269(.A0(n6670), .A1(n6508), .B0(n6874), .Y(n6877));
  NOR4X1  g05270(.A(n6876), .B(n6875), .C(n6867), .D(n6877), .Y(n6878));
  INVX1   g05271(.A(n6878), .Y(n6879));
  NAND2X1 g05272(.A(n6832), .B(n6830), .Y(n6884));
  XOR2X1  g05273(.A(n6851), .B(n6884), .Y(n6885));
  INVX1   g05274(.A(n6851), .Y(n6886));
  AOI22X1 g05275(.A0(n6556), .A1(P2_REG2_REG_8__SCAN_IN), .B0(P2_REG0_REG_8__SCAN_IN), .B1(n6557), .Y(n6887));
  INVX1   g05276(.A(P2_REG3_REG_8__SCAN_IN), .Y(n6888));
  INVX1   g05277(.A(P2_REG3_REG_7__SCAN_IN), .Y(n6889));
  NOR4X1  g05278(.A(n6889), .B(n6782), .C(n6781), .D(n6729), .Y(n6890));
  XOR2X1  g05279(.A(n6890), .B(n6888), .Y(n6891));
  INVX1   g05280(.A(n6891), .Y(n6892));
  AOI22X1 g05281(.A0(n6502), .A1(n6892), .B0(n6559), .B1(P2_REG1_REG_8__SCAN_IN), .Y(n6893));
  NAND2X1 g05282(.A(n6893), .B(n6887), .Y(n6894));
  INVX1   g05283(.A(n6894), .Y(n6895));
  OAI22X1 g05284(.A0(n6886), .A1(n6528), .B0(n6535), .B1(n6895), .Y(n6896));
  AOI21X1 g05285(.A0(n6885), .A1(n6532), .B0(n6896), .Y(n6897));
  OAI21X1 g05286(.A0(n6864), .A1(n6525), .B0(n6897), .Y(n6898));
  NOR2X1  g05287(.A(n6898), .B(n6879), .Y(n6899));
  NAND2X1 g05288(.A(n6465), .B(P2_REG0_REG_7__SCAN_IN), .Y(n6900));
  OAI21X1 g05289(.A0(n6899), .A1(n6465), .B0(n6900), .Y(P2_U3451));
  AOI21X1 g05290(.A0(n6886), .A1(n6856), .B0(n6840), .Y(n6902));
  AOI21X1 g05291(.A0(n6851), .A1(n6857), .B0(n6902), .Y(n6903));
  OAI21X1 g05292(.A0(n6852), .A1(n6806), .B0(n6903), .Y(n6904));
  NOR2X1  g05293(.A(P2_IR_REG_31__SCAN_IN), .B(n6288), .Y(n6905));
  AOI21X1 g05294(.A0(n6129), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6905), .Y(n6906));
  INVX1   g05295(.A(n6906), .Y(n6907));
  NAND3X1 g05296(.A(n6907), .B(n6481), .C(n6480), .Y(n6908));
  OAI21X1 g05297(.A0(n6474), .A1(n6124), .B0(n6908), .Y(n6909));
  XOR2X1  g05298(.A(n6909), .B(n6895), .Y(n6910));
  NOR2X1  g05299(.A(n6904), .B(n6910), .Y(n6911));
  AOI21X1 g05300(.A0(n6910), .A1(n6904), .B0(n6911), .Y(n6913));
  INVX1   g05301(.A(n6913), .Y(n6914));
  OAI21X1 g05302(.A0(n6520), .A1(n6514), .B0(n6914), .Y(n6915));
  NOR2X1  g05303(.A(n6851), .B(n6840), .Y(n6916));
  NAND2X1 g05304(.A(n6715), .B(n6714), .Y(n6917));
  AOI21X1 g05305(.A0(n6712), .A1(n6613), .B0(n6917), .Y(n6918));
  NOR4X1  g05306(.A(n6758), .B(n6918), .C(n6765), .D(n6868), .Y(n6919));
  NOR3X1  g05307(.A(n6919), .B(n6871), .C(n6916), .Y(n6920));
  AOI21X1 g05308(.A0(n6851), .A1(n6840), .B0(n6910), .Y(n6921));
  INVX1   g05309(.A(n6921), .Y(n6922));
  AOI21X1 g05310(.A0(n6851), .A1(n6840), .B0(n6873), .Y(n6923));
  INVX1   g05311(.A(n6916), .Y(n6924));
  NAND2X1 g05312(.A(n6910), .B(n6924), .Y(n6925));
  OAI22X1 g05313(.A0(n6923), .A1(n6925), .B0(n6922), .B1(n6920), .Y(n6926));
  AOI22X1 g05314(.A0(n6914), .A1(n6518), .B0(n6512), .B1(n6926), .Y(n6927));
  AOI22X1 g05315(.A0(n6839), .A1(n6574), .B0(n6521), .B1(n6926), .Y(n6928));
  OAI21X1 g05316(.A0(n6516), .A1(n6507), .B0(n6926), .Y(n6929));
  NAND4X1 g05317(.A(n6928), .B(n6927), .C(n6915), .D(n6929), .Y(n6930));
  NOR4X1  g05318(.A(n6797), .B(n6752), .C(n6775), .D(n6851), .Y(n6934));
  INVX1   g05319(.A(n6909), .Y(n6935));
  XOR2X1  g05320(.A(n6935), .B(n6934), .Y(n6936));
  AOI22X1 g05321(.A0(n6556), .A1(P2_REG2_REG_9__SCAN_IN), .B0(P2_REG0_REG_9__SCAN_IN), .B1(n6557), .Y(n6937));
  INVX1   g05322(.A(P2_REG3_REG_9__SCAN_IN), .Y(n6938));
  INVX1   g05323(.A(n6890), .Y(n6939));
  NOR2X1  g05324(.A(n6939), .B(n6888), .Y(n6940));
  XOR2X1  g05325(.A(n6940), .B(n6938), .Y(n6941));
  INVX1   g05326(.A(n6941), .Y(n6942));
  AOI22X1 g05327(.A0(n6502), .A1(n6942), .B0(n6559), .B1(P2_REG1_REG_9__SCAN_IN), .Y(n6943));
  NAND2X1 g05328(.A(n6943), .B(n6937), .Y(n6944));
  INVX1   g05329(.A(n6944), .Y(n6945));
  OAI22X1 g05330(.A0(n6935), .A1(n6528), .B0(n6535), .B1(n6945), .Y(n6946));
  AOI21X1 g05331(.A0(n6936), .A1(n6532), .B0(n6946), .Y(n6947));
  OAI21X1 g05332(.A0(n6913), .A1(n6525), .B0(n6947), .Y(n6948));
  NOR2X1  g05333(.A(n6948), .B(n6930), .Y(n6949));
  NAND2X1 g05334(.A(n6465), .B(P2_REG0_REG_8__SCAN_IN), .Y(n6950));
  OAI21X1 g05335(.A0(n6949), .A1(n6465), .B0(n6950), .Y(P2_U3454));
  NOR2X1  g05336(.A(P2_IR_REG_31__SCAN_IN), .B(n6134), .Y(n6952));
  AOI21X1 g05337(.A0(n6135), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6952), .Y(n6953));
  INVX1   g05338(.A(n6953), .Y(n6954));
  NAND3X1 g05339(.A(n6954), .B(n6481), .C(n6480), .Y(n6955));
  OAI21X1 g05340(.A0(n6474), .A1(n6133), .B0(n6955), .Y(n6956));
  XOR2X1  g05341(.A(n6956), .B(n6945), .Y(n6957));
  AOI22X1 g05342(.A0(n6895), .A1(n6909), .B0(n6851), .B1(n6840), .Y(n6958));
  INVX1   g05343(.A(n6958), .Y(n6959));
  NOR2X1  g05344(.A(n6959), .B(n6873), .Y(n6960));
  OAI21X1 g05345(.A0(n6894), .A1(n6916), .B0(n6935), .Y(n6961));
  OAI21X1 g05346(.A0(n6895), .A1(n6924), .B0(n6961), .Y(n6962));
  NOR2X1  g05347(.A(n6962), .B(n6960), .Y(n6963));
  XOR2X1  g05348(.A(n6963), .B(n6957), .Y(n6964));
  INVX1   g05349(.A(n6964), .Y(n6965));
  OAI21X1 g05350(.A0(n6516), .A1(n6507), .B0(n6965), .Y(n6966));
  OAI21X1 g05351(.A0(n6964), .A1(n6669), .B0(n6966), .Y(n6967));
  NAND2X1 g05352(.A(n6935), .B(n6895), .Y(n6969));
  NOR2X1  g05353(.A(n6935), .B(n6895), .Y(n6970));
  AOI21X1 g05354(.A0(n6969), .A1(n6904), .B0(n6970), .Y(n6971));
  XOR2X1  g05355(.A(n6956), .B(n6944), .Y(n6972));
  NOR2X1  g05356(.A(n6972), .B(n6971), .Y(n6973));
  AOI21X1 g05357(.A0(n6971), .A1(n6972), .B0(n6973), .Y(n6974));
  NOR2X1  g05358(.A(n6974), .B(n6657), .Y(n6975));
  OAI22X1 g05359(.A0(n6895), .A1(n6634), .B0(n6661), .B1(n6964), .Y(n6976));
  AOI21X1 g05360(.A0(n6658), .A1(n6633), .B0(n6974), .Y(n6977));
  NOR4X1  g05361(.A(n6976), .B(n6975), .C(n6967), .D(n6977), .Y(n6978));
  INVX1   g05362(.A(n6978), .Y(n6979));
  NOR3X1  g05363(.A(n6909), .B(n6851), .C(n6884), .Y(n6983));
  INVX1   g05364(.A(n6956), .Y(n6984));
  XOR2X1  g05365(.A(n6984), .B(n6983), .Y(n6985));
  AOI22X1 g05366(.A0(n6556), .A1(P2_REG2_REG_10__SCAN_IN), .B0(P2_REG0_REG_10__SCAN_IN), .B1(n6557), .Y(n6986));
  INVX1   g05367(.A(P2_REG3_REG_10__SCAN_IN), .Y(n6987));
  NOR3X1  g05368(.A(n6939), .B(n6888), .C(n6938), .Y(n6988));
  XOR2X1  g05369(.A(n6988), .B(n6987), .Y(n6989));
  INVX1   g05370(.A(n6989), .Y(n6990));
  AOI22X1 g05371(.A0(n6502), .A1(n6990), .B0(n6559), .B1(P2_REG1_REG_10__SCAN_IN), .Y(n6991));
  NAND2X1 g05372(.A(n6991), .B(n6986), .Y(n6992));
  INVX1   g05373(.A(n6992), .Y(n6993));
  OAI22X1 g05374(.A0(n6984), .A1(n6528), .B0(n6535), .B1(n6993), .Y(n6994));
  AOI21X1 g05375(.A0(n6985), .A1(n6532), .B0(n6994), .Y(n6995));
  OAI21X1 g05376(.A0(n6974), .A1(n6525), .B0(n6995), .Y(n6996));
  NOR2X1  g05377(.A(n6996), .B(n6979), .Y(n6997));
  NAND2X1 g05378(.A(n6465), .B(P2_REG0_REG_9__SCAN_IN), .Y(n6998));
  OAI21X1 g05379(.A0(n6997), .A1(n6465), .B0(n6998), .Y(P2_U3457));
  NOR2X1  g05380(.A(P2_IR_REG_31__SCAN_IN), .B(n6140), .Y(n7000));
  AOI21X1 g05381(.A0(n6143), .A1(P2_IR_REG_31__SCAN_IN), .B0(n7000), .Y(n7001));
  INVX1   g05382(.A(n7001), .Y(n7002));
  NAND3X1 g05383(.A(n7002), .B(n6481), .C(n6480), .Y(n7003));
  OAI21X1 g05384(.A0(n6474), .A1(n6139), .B0(n7003), .Y(n7004));
  NOR2X1  g05385(.A(n6956), .B(n6944), .Y(n7005));
  INVX1   g05386(.A(n7004), .Y(n7006));
  AOI21X1 g05387(.A0(n7006), .A1(n6993), .B0(n7005), .Y(n7007));
  INVX1   g05388(.A(n7007), .Y(n7008));
  AOI21X1 g05389(.A0(n7004), .A1(n6992), .B0(n7008), .Y(n7009));
  INVX1   g05390(.A(n7009), .Y(n7010));
  INVX1   g05391(.A(n6971), .Y(n7011));
  NOR2X1  g05392(.A(n6984), .B(n6945), .Y(n7012));
  NOR2X1  g05393(.A(n7012), .B(n7011), .Y(n7013));
  XOR2X1  g05394(.A(n7004), .B(n6993), .Y(n7014));
  NOR2X1  g05395(.A(n9408), .B(n7012), .Y(n7016));
  INVX1   g05396(.A(n7016), .Y(n7017));
  NOR2X1  g05397(.A(n7005), .B(n6971), .Y(n7018));
  OAI22X1 g05398(.A0(n7017), .A1(n7018), .B0(n7013), .B1(n7010), .Y(n7019));
  INVX1   g05399(.A(n7019), .Y(n7020));
  OAI21X1 g05400(.A0(n6520), .A1(n6514), .B0(n7020), .Y(n7021));
  INVX1   g05401(.A(n7021), .Y(n7022));
  NAND2X1 g05402(.A(n6956), .B(n6945), .Y(n7023));
  INVX1   g05403(.A(n7023), .Y(n7024));
  OAI21X1 g05404(.A0(n6919), .A1(n6871), .B0(n6958), .Y(n7025));
  AOI21X1 g05405(.A0(n6895), .A1(n6924), .B0(n6909), .Y(n7026));
  AOI21X1 g05406(.A0(n6894), .A1(n6916), .B0(n7026), .Y(n7027));
  AOI21X1 g05407(.A0(n7027), .A1(n7025), .B0(n7024), .Y(n7028));
  AOI21X1 g05408(.A0(n6984), .A1(n6944), .B0(n7028), .Y(n7029));
  XOR2X1  g05409(.A(n7029), .B(n7014), .Y(n7030));
  OAI22X1 g05410(.A0(n7019), .A1(n6633), .B0(n6669), .B1(n7030), .Y(n7031));
  OAI22X1 g05411(.A0(n6945), .A1(n6634), .B0(n6661), .B1(n7030), .Y(n7032));
  AOI21X1 g05412(.A0(n6670), .A1(n6508), .B0(n7030), .Y(n7033));
  NOR4X1  g05413(.A(n7032), .B(n7031), .C(n7022), .D(n7033), .Y(n7034));
  INVX1   g05414(.A(n7034), .Y(n7035));
  NAND3X1 g05415(.A(n6984), .B(n6935), .C(n6934), .Y(n7040));
  NOR2X1  g05416(.A(n7004), .B(n6956), .Y(n7041));
  AOI22X1 g05417(.A0(n7004), .A1(n7040), .B0(n6983), .B1(n7041), .Y(n7042));
  AOI22X1 g05418(.A0(n6556), .A1(P2_REG2_REG_11__SCAN_IN), .B0(P2_REG0_REG_11__SCAN_IN), .B1(n6557), .Y(n7043));
  INVX1   g05419(.A(n7043), .Y(n7044));
  INVX1   g05420(.A(P2_REG3_REG_11__SCAN_IN), .Y(n7045));
  NOR4X1  g05421(.A(n6987), .B(n6888), .C(n6938), .D(n6939), .Y(n7046));
  XOR2X1  g05422(.A(n7046), .B(n7045), .Y(n7047));
  INVX1   g05423(.A(n7047), .Y(n7048));
  AOI22X1 g05424(.A0(n6502), .A1(n7048), .B0(n6559), .B1(P2_REG1_REG_11__SCAN_IN), .Y(n7049));
  INVX1   g05425(.A(n7049), .Y(n7050));
  NOR2X1  g05426(.A(n7050), .B(n7044), .Y(n7051));
  OAI22X1 g05427(.A0(n7006), .A1(n6528), .B0(n6535), .B1(n7051), .Y(n7052));
  AOI21X1 g05428(.A0(n7042), .A1(n6532), .B0(n7052), .Y(n7053));
  OAI21X1 g05429(.A0(n7019), .A1(n6525), .B0(n7053), .Y(n7054));
  NOR2X1  g05430(.A(n7054), .B(n7035), .Y(n7055));
  NAND2X1 g05431(.A(n6465), .B(P2_REG0_REG_10__SCAN_IN), .Y(n7056));
  OAI21X1 g05432(.A0(n7055), .A1(n6465), .B0(n7056), .Y(P2_U3460));
  OAI21X1 g05433(.A0(n7004), .A1(n6993), .B0(n7029), .Y(n7058));
  NOR2X1  g05434(.A(P2_IR_REG_31__SCAN_IN), .B(n6148), .Y(n7059));
  AOI21X1 g05435(.A0(n6152), .A1(P2_IR_REG_31__SCAN_IN), .B0(n7059), .Y(n7060));
  INVX1   g05436(.A(n7060), .Y(n7061));
  NAND2X1 g05437(.A(n7061), .B(n6474), .Y(n7062));
  OAI21X1 g05438(.A0(n6474), .A1(n6147), .B0(n7062), .Y(n7063));
  XOR2X1  g05439(.A(n7063), .B(n7051), .Y(n7064));
  AOI21X1 g05440(.A0(n7004), .A1(n6993), .B0(n7064), .Y(n7065));
  NAND2X1 g05441(.A(n7004), .B(n6993), .Y(n7066));
  INVX1   g05442(.A(n7066), .Y(n7067));
  NOR2X1  g05443(.A(n7029), .B(n7067), .Y(n7068));
  INVX1   g05444(.A(n7068), .Y(n7069));
  NAND2X1 g05445(.A(n7063), .B(n7051), .Y(n7070));
  INVX1   g05446(.A(n7070), .Y(n7071));
  INVX1   g05447(.A(n7051), .Y(n7072));
  INVX1   g05448(.A(n7063), .Y(n7073));
  AOI22X1 g05449(.A0(n7072), .A1(n7073), .B0(n7006), .B1(n6992), .Y(n7074));
  INVX1   g05450(.A(n7074), .Y(n7075));
  NOR2X1  g05451(.A(n7075), .B(n7071), .Y(n7076));
  AOI22X1 g05452(.A0(n7069), .A1(n7076), .B0(n7065), .B1(n7058), .Y(n7077));
  NAND2X1 g05453(.A(n7007), .B(n6970), .Y(n7079));
  AOI22X1 g05454(.A0(n6992), .A1(n7004), .B0(n6956), .B1(n6944), .Y(n7080));
  AOI22X1 g05455(.A0(n7079), .A1(n7080), .B0(n7006), .B1(n6993), .Y(n7081));
  AOI21X1 g05456(.A0(n6935), .A1(n6895), .B0(n7008), .Y(n7082));
  AOI21X1 g05457(.A0(n7082), .A1(n6904), .B0(n7081), .Y(n7083));
  XOR2X1  g05458(.A(n7063), .B(n7072), .Y(n7084));
  NOR2X1  g05459(.A(n7084), .B(n7083), .Y(n7085));
  AOI21X1 g05460(.A0(n7083), .A1(n7084), .B0(n7085), .Y(n7086));
  OAI22X1 g05461(.A0(n6993), .A1(n6634), .B0(n6633), .B1(n7086), .Y(n7087));
  AOI21X1 g05462(.A0(n6658), .A1(n6657), .B0(n7086), .Y(n7088));
  NOR2X1  g05463(.A(n7088), .B(n7087), .Y(n7089));
  OAI21X1 g05464(.A0(n7077), .A1(n6661), .B0(n7089), .Y(n7090));
  NOR2X1  g05465(.A(n7077), .B(n6669), .Y(n7091));
  AOI21X1 g05466(.A0(n6670), .A1(n6508), .B0(n7077), .Y(n7092));
  NAND3X1 g05467(.A(n7041), .B(n6935), .C(n6934), .Y(n7096));
  XOR2X1  g05468(.A(n7063), .B(n7096), .Y(n7097));
  AOI22X1 g05469(.A0(n6556), .A1(P2_REG2_REG_12__SCAN_IN), .B0(P2_REG0_REG_12__SCAN_IN), .B1(n6557), .Y(n7098));
  NAND2X1 g05470(.A(P2_REG3_REG_10__SCAN_IN), .B(P2_REG3_REG_11__SCAN_IN), .Y(n7099));
  NOR4X1  g05471(.A(n6939), .B(n6888), .C(n6938), .D(n7099), .Y(n7100));
  XOR2X1  g05472(.A(n7100), .B(P2_REG3_REG_12__SCAN_IN), .Y(n7101));
  AOI22X1 g05473(.A0(n6502), .A1(n7101), .B0(n6559), .B1(P2_REG1_REG_12__SCAN_IN), .Y(n7102));
  NAND2X1 g05474(.A(n7102), .B(n7098), .Y(n7103));
  INVX1   g05475(.A(n7103), .Y(n7104));
  OAI22X1 g05476(.A0(n7073), .A1(n6528), .B0(n6535), .B1(n7104), .Y(n7105));
  AOI21X1 g05477(.A0(n7097), .A1(n6532), .B0(n7105), .Y(n7106));
  OAI21X1 g05478(.A0(n7086), .A1(n6525), .B0(n7106), .Y(n7107));
  NOR4X1  g05479(.A(n7092), .B(n7091), .C(n7090), .D(n7107), .Y(n7108));
  NAND2X1 g05480(.A(n6465), .B(P2_REG0_REG_11__SCAN_IN), .Y(n7109));
  OAI21X1 g05481(.A0(n7108), .A1(n6465), .B0(n7109), .Y(P2_U3463));
  NOR2X1  g05482(.A(P2_IR_REG_31__SCAN_IN), .B(n6191), .Y(n7111));
  AOI21X1 g05483(.A0(n6159), .A1(P2_IR_REG_31__SCAN_IN), .B0(n7111), .Y(n7112));
  INVX1   g05484(.A(n7112), .Y(n7113));
  NAND2X1 g05485(.A(n7113), .B(n6474), .Y(n7114));
  OAI21X1 g05486(.A0(n6474), .A1(n6156), .B0(n7114), .Y(n7115));
  XOR2X1  g05487(.A(n7115), .B(n7104), .Y(n7116));
  NAND3X1 g05488(.A(n7066), .B(n6984), .C(n6944), .Y(n7117));
  AOI21X1 g05489(.A0(n7117), .A1(n7074), .B0(n7071), .Y(n7118));
  NAND3X1 g05490(.A(n7070), .B(n7066), .C(n7023), .Y(n7119));
  AOI21X1 g05491(.A0(n7027), .A1(n7025), .B0(n7119), .Y(n7120));
  NOR2X1  g05492(.A(n7120), .B(n7118), .Y(n7121));
  XOR2X1  g05493(.A(n7121), .B(n7116), .Y(n7122));
  INVX1   g05494(.A(n7122), .Y(n7123));
  OAI21X1 g05495(.A0(n6516), .A1(n6507), .B0(n7123), .Y(n7124));
  OAI21X1 g05496(.A0(n7122), .A1(n6669), .B0(n7124), .Y(n7125));
  INVX1   g05497(.A(n7083), .Y(n7127));
  NOR2X1  g05498(.A(n7063), .B(n7072), .Y(n7128));
  INVX1   g05499(.A(n7128), .Y(n7129));
  NOR2X1  g05500(.A(n7073), .B(n7051), .Y(n7130));
  AOI21X1 g05501(.A0(n7129), .A1(n7127), .B0(n7130), .Y(n7131));
  XOR2X1  g05502(.A(n7115), .B(n7103), .Y(n7132));
  NOR2X1  g05503(.A(n7132), .B(n7131), .Y(n7133));
  AOI21X1 g05504(.A0(n7131), .A1(n7132), .B0(n7133), .Y(n7134));
  NOR2X1  g05505(.A(n7134), .B(n6657), .Y(n7135));
  OAI22X1 g05506(.A0(n7051), .A1(n6634), .B0(n6661), .B1(n7122), .Y(n7136));
  AOI21X1 g05507(.A0(n6658), .A1(n6633), .B0(n7134), .Y(n7137));
  NOR4X1  g05508(.A(n7136), .B(n7135), .C(n7125), .D(n7137), .Y(n7138));
  INVX1   g05509(.A(n7138), .Y(n7139));
  NOR2X1  g05510(.A(n7134), .B(n6525), .Y(n7144));
  NAND4X1 g05511(.A(n7041), .B(n6935), .C(n6934), .D(n7073), .Y(n7145));
  NOR2X1  g05512(.A(n6474), .B(n6156), .Y(n7146));
  AOI21X1 g05513(.A0(n7113), .A1(n6474), .B0(n7146), .Y(n7147));
  XOR2X1  g05514(.A(n7147), .B(n7145), .Y(n7148));
  AOI22X1 g05515(.A0(n6556), .A1(P2_REG2_REG_13__SCAN_IN), .B0(P2_REG0_REG_13__SCAN_IN), .B1(n6557), .Y(n7149));
  NAND2X1 g05516(.A(n7100), .B(P2_REG3_REG_12__SCAN_IN), .Y(n7150));
  XOR2X1  g05517(.A(n7150), .B(P2_REG3_REG_13__SCAN_IN), .Y(n7151));
  INVX1   g05518(.A(n7151), .Y(n7152));
  AOI22X1 g05519(.A0(n6502), .A1(n7152), .B0(n6559), .B1(P2_REG1_REG_13__SCAN_IN), .Y(n7153));
  NAND2X1 g05520(.A(n7153), .B(n7149), .Y(n7154));
  AOI22X1 g05521(.A0(n7115), .A1(n6529), .B0(n6534), .B1(n7154), .Y(n7155));
  OAI21X1 g05522(.A0(n7148), .A1(n6533), .B0(n7155), .Y(n7156));
  NOR3X1  g05523(.A(n7156), .B(n7144), .C(n7139), .Y(n7157));
  NAND2X1 g05524(.A(n6465), .B(P2_REG0_REG_12__SCAN_IN), .Y(n7158));
  OAI21X1 g05525(.A0(n7157), .A1(n6465), .B0(n7158), .Y(P2_U3466));
  NOR2X1  g05526(.A(P2_IR_REG_31__SCAN_IN), .B(n6164), .Y(n7160));
  AOI21X1 g05527(.A0(n6165), .A1(P2_IR_REG_31__SCAN_IN), .B0(n7160), .Y(n7161));
  INVX1   g05528(.A(n7161), .Y(n7162));
  NAND2X1 g05529(.A(n7162), .B(n6474), .Y(n7163));
  OAI21X1 g05530(.A0(n6474), .A1(n6163), .B0(n7163), .Y(n7164));
  INVX1   g05531(.A(n7154), .Y(n7165));
  NOR2X1  g05532(.A(n6474), .B(n6163), .Y(n7166));
  AOI21X1 g05533(.A0(n7162), .A1(n6474), .B0(n7166), .Y(n7167));
  AOI22X1 g05534(.A0(n7165), .A1(n7167), .B0(n7147), .B1(n7104), .Y(n7168));
  INVX1   g05535(.A(n7168), .Y(n7169));
  AOI21X1 g05536(.A0(n7164), .A1(n7154), .B0(n7169), .Y(n7170));
  INVX1   g05537(.A(n7170), .Y(n7171));
  NOR2X1  g05538(.A(n7128), .B(n7083), .Y(n7172));
  NOR2X1  g05539(.A(n7147), .B(n7104), .Y(n7173));
  NOR3X1  g05540(.A(n7173), .B(n7172), .C(n7130), .Y(n7174));
  NAND2X1 g05541(.A(n7147), .B(n7104), .Y(n7175));
  INVX1   g05542(.A(n7175), .Y(n7176));
  XOR2X1  g05543(.A(n7164), .B(n7165), .Y(n7177));
  INVX1   g05544(.A(n7177), .Y(n7178));
  NOR2X1  g05545(.A(n7178), .B(n7173), .Y(n7179));
  OAI21X1 g05546(.A0(n7176), .A1(n7131), .B0(n7179), .Y(n7180));
  OAI21X1 g05547(.A0(n7174), .A1(n7171), .B0(n7180), .Y(n7181));
  INVX1   g05548(.A(n7181), .Y(n7182));
  OAI21X1 g05549(.A0(n6520), .A1(n6514), .B0(n7182), .Y(n7183));
  NOR2X1  g05550(.A(n7115), .B(n7104), .Y(n7184));
  INVX1   g05551(.A(n7184), .Y(n7185));
  OAI22X1 g05552(.A0(n7118), .A1(n7120), .B0(n7147), .B1(n7103), .Y(n7186));
  NAND2X1 g05553(.A(n7186), .B(n7185), .Y(n7187));
  XOR2X1  g05554(.A(n7187), .B(n7178), .Y(n7188));
  NOR2X1  g05555(.A(n7188), .B(n6669), .Y(n7189));
  AOI21X1 g05556(.A0(n7182), .A1(n6518), .B0(n7189), .Y(n7190));
  OAI22X1 g05557(.A0(n7104), .A1(n6634), .B0(n6661), .B1(n7188), .Y(n7191));
  AOI21X1 g05558(.A0(n6670), .A1(n6508), .B0(n7188), .Y(n7192));
  NOR2X1  g05559(.A(n7192), .B(n7191), .Y(n7193));
  NAND3X1 g05560(.A(n7193), .B(n7190), .C(n7183), .Y(n7194));
  NAND4X1 g05561(.A(n7073), .B(n7041), .C(n6983), .D(n7147), .Y(n7199));
  XOR2X1  g05562(.A(n7164), .B(n7199), .Y(n7200));
  AOI22X1 g05563(.A0(n6556), .A1(P2_REG2_REG_14__SCAN_IN), .B0(P2_REG0_REG_14__SCAN_IN), .B1(n6557), .Y(n7201));
  NAND3X1 g05564(.A(n7100), .B(P2_REG3_REG_12__SCAN_IN), .C(P2_REG3_REG_13__SCAN_IN), .Y(n7202));
  XOR2X1  g05565(.A(n7202), .B(P2_REG3_REG_14__SCAN_IN), .Y(n7203));
  INVX1   g05566(.A(n7203), .Y(n7204));
  AOI22X1 g05567(.A0(n6502), .A1(n7204), .B0(n6559), .B1(P2_REG1_REG_14__SCAN_IN), .Y(n7205));
  NAND2X1 g05568(.A(n7205), .B(n7201), .Y(n7206));
  INVX1   g05569(.A(n7206), .Y(n7207));
  OAI22X1 g05570(.A0(n7167), .A1(n6528), .B0(n6535), .B1(n7207), .Y(n7208));
  AOI21X1 g05571(.A0(n7200), .A1(n6532), .B0(n7208), .Y(n7209));
  OAI21X1 g05572(.A0(n7181), .A1(n6525), .B0(n7209), .Y(n7210));
  NOR2X1  g05573(.A(n7210), .B(n7194), .Y(n7211));
  NAND2X1 g05574(.A(n6465), .B(P2_REG0_REG_13__SCAN_IN), .Y(n7212));
  OAI21X1 g05575(.A0(n7211), .A1(n6465), .B0(n7212), .Y(P2_U3469));
  NOR2X1  g05576(.A(P2_IR_REG_31__SCAN_IN), .B(n6170), .Y(n7214));
  AOI21X1 g05577(.A0(n6174), .A1(P2_IR_REG_31__SCAN_IN), .B0(n7214), .Y(n7215));
  INVX1   g05578(.A(n7215), .Y(n7216));
  NOR2X1  g05579(.A(n6474), .B(n6169), .Y(n7217));
  AOI21X1 g05580(.A0(n7216), .A1(n6474), .B0(n7217), .Y(n7218));
  XOR2X1  g05581(.A(n7218), .B(n7206), .Y(n7219));
  NOR2X1  g05582(.A(n7164), .B(n7165), .Y(n7220));
  AOI22X1 g05583(.A0(n7164), .A1(n7165), .B0(n7185), .B1(n7186), .Y(n7221));
  NOR2X1  g05584(.A(n7221), .B(n7220), .Y(n7222));
  XOR2X1  g05585(.A(n7222), .B(n7219), .Y(n7223));
  NOR2X1  g05586(.A(n7223), .B(n6661), .Y(n7224));
  NAND2X1 g05587(.A(n7168), .B(n7130), .Y(n7225));
  AOI22X1 g05588(.A0(n7154), .A1(n7164), .B0(n7115), .B1(n7103), .Y(n7226));
  NAND2X1 g05589(.A(n7226), .B(n7225), .Y(n7227));
  OAI21X1 g05590(.A0(n7164), .A1(n7154), .B0(n7227), .Y(n7228));
  NAND2X1 g05591(.A(n7168), .B(n7129), .Y(n7229));
  OAI21X1 g05592(.A0(n7229), .A1(n7083), .B0(n7228), .Y(n7230));
  XOR2X1  g05593(.A(n7230), .B(n7219), .Y(n7231));
  INVX1   g05594(.A(n7231), .Y(n7232));
  AOI22X1 g05595(.A0(n7154), .A1(n6574), .B0(n6518), .B1(n7232), .Y(n7233));
  OAI21X1 g05596(.A0(n6520), .A1(n6514), .B0(n7232), .Y(n7234));
  NAND2X1 g05597(.A(n7234), .B(n7233), .Y(n7235));
  NOR2X1  g05598(.A(n7223), .B(n6669), .Y(n7236));
  AOI21X1 g05599(.A0(n6670), .A1(n6508), .B0(n7223), .Y(n7237));
  NOR4X1  g05600(.A(n7236), .B(n7235), .C(n7224), .D(n7237), .Y(n7238));
  INVX1   g05601(.A(n7238), .Y(n7239));
  AOI22X1 g05602(.A0(n7225), .A1(n7226), .B0(n7167), .B1(n7165), .Y(n7240));
  NOR2X1  g05603(.A(n7229), .B(n7083), .Y(n7241));
  NOR2X1  g05604(.A(n7241), .B(n7240), .Y(n7242));
  NOR2X1  g05605(.A(n7231), .B(n6525), .Y(n7245));
  NOR3X1  g05606(.A(n7164), .B(n7115), .C(n7145), .Y(n7246));
  NAND2X1 g05607(.A(n7218), .B(n7167), .Y(n7247));
  OAI22X1 g05608(.A0(n7218), .A1(n7246), .B0(n7199), .B1(n7247), .Y(n7248));
  INVX1   g05609(.A(n7218), .Y(n7249));
  AOI22X1 g05610(.A0(n6556), .A1(P2_REG2_REG_15__SCAN_IN), .B0(P2_REG0_REG_15__SCAN_IN), .B1(n6557), .Y(n7250));
  NAND4X1 g05611(.A(P2_REG3_REG_14__SCAN_IN), .B(P2_REG3_REG_12__SCAN_IN), .C(P2_REG3_REG_13__SCAN_IN), .D(n7100), .Y(n7251));
  XOR2X1  g05612(.A(n7251), .B(P2_REG3_REG_15__SCAN_IN), .Y(n7252));
  INVX1   g05613(.A(n7252), .Y(n7253));
  AOI22X1 g05614(.A0(n6502), .A1(n7253), .B0(n6559), .B1(P2_REG1_REG_15__SCAN_IN), .Y(n7254));
  NAND2X1 g05615(.A(n7254), .B(n7250), .Y(n7255));
  AOI22X1 g05616(.A0(n7249), .A1(n6529), .B0(n6534), .B1(n7255), .Y(n7256));
  OAI21X1 g05617(.A0(n7248), .A1(n6533), .B0(n7256), .Y(n7257));
  NOR3X1  g05618(.A(n7257), .B(n7245), .C(n7239), .Y(n7258));
  NAND2X1 g05619(.A(n6465), .B(P2_REG0_REG_14__SCAN_IN), .Y(n7259));
  OAI21X1 g05620(.A0(n7258), .A1(n6465), .B0(n7259), .Y(P2_U3472));
  NOR2X1  g05621(.A(P2_IR_REG_31__SCAN_IN), .B(n6180), .Y(n7261));
  AOI21X1 g05622(.A0(n6181), .A1(P2_IR_REG_31__SCAN_IN), .B0(n7261), .Y(n7262));
  INVX1   g05623(.A(n7262), .Y(n7263));
  NOR2X1  g05624(.A(n6474), .B(n6179), .Y(n7264));
  AOI21X1 g05625(.A0(n7263), .A1(n6474), .B0(n7264), .Y(n7265));
  XOR2X1  g05626(.A(n7265), .B(n7255), .Y(n7266));
  INVX1   g05627(.A(n7220), .Y(n7267));
  NOR2X1  g05628(.A(n7218), .B(n7206), .Y(n7268));
  INVX1   g05629(.A(n7118), .Y(n7269));
  INVX1   g05630(.A(n7119), .Y(n7270));
  OAI21X1 g05631(.A0(n6962), .A1(n6960), .B0(n7270), .Y(n7271));
  AOI22X1 g05632(.A0(n7269), .A1(n7271), .B0(n7115), .B1(n7104), .Y(n7272));
  OAI22X1 g05633(.A0(n7167), .A1(n7154), .B0(n7184), .B1(n7272), .Y(n7273));
  AOI21X1 g05634(.A0(n7273), .A1(n7267), .B0(n7268), .Y(n7274));
  AOI21X1 g05635(.A0(n7218), .A1(n7206), .B0(n7274), .Y(n7275));
  XOR2X1  g05636(.A(n7275), .B(n7266), .Y(n7276));
  NOR2X1  g05637(.A(n7276), .B(n6661), .Y(n7277));
  INVX1   g05638(.A(n7266), .Y(n7278));
  NOR2X1  g05639(.A(n7218), .B(n7207), .Y(n7279));
  NOR2X1  g05640(.A(n7249), .B(n7206), .Y(n7280));
  INVX1   g05641(.A(n7280), .Y(n7281));
  AOI21X1 g05642(.A0(n7281), .A1(n7230), .B0(n7279), .Y(n7282));
  XOR2X1  g05643(.A(n7282), .B(n7278), .Y(n7283));
  INVX1   g05644(.A(n7283), .Y(n7284));
  AOI22X1 g05645(.A0(n7206), .A1(n6574), .B0(n6518), .B1(n7284), .Y(n7285));
  OAI21X1 g05646(.A0(n6520), .A1(n6514), .B0(n7284), .Y(n7286));
  NAND2X1 g05647(.A(n7286), .B(n7285), .Y(n7287));
  NOR2X1  g05648(.A(n7276), .B(n6669), .Y(n7288));
  AOI21X1 g05649(.A0(n6670), .A1(n6508), .B0(n7276), .Y(n7289));
  NOR4X1  g05650(.A(n7288), .B(n7287), .C(n7277), .D(n7289), .Y(n7290));
  INVX1   g05651(.A(n7290), .Y(n7291));
  INVX1   g05652(.A(n7279), .Y(n7292));
  OAI21X1 g05653(.A0(n7280), .A1(n7242), .B0(n7292), .Y(n7293));
  NOR3X1  g05654(.A(n7249), .B(n7164), .C(n7199), .Y(n7295));
  XOR2X1  g05655(.A(n7265), .B(n7295), .Y(n7296));
  AOI22X1 g05656(.A0(n6556), .A1(P2_REG2_REG_16__SCAN_IN), .B0(P2_REG0_REG_16__SCAN_IN), .B1(n6557), .Y(n7297));
  INVX1   g05657(.A(P2_REG3_REG_16__SCAN_IN), .Y(n7298));
  INVX1   g05658(.A(P2_REG3_REG_15__SCAN_IN), .Y(n7299));
  NOR2X1  g05659(.A(n7251), .B(n7299), .Y(n7300));
  XOR2X1  g05660(.A(n7300), .B(n7298), .Y(n7301));
  INVX1   g05661(.A(n7301), .Y(n7302));
  AOI22X1 g05662(.A0(n6502), .A1(n7302), .B0(n6559), .B1(P2_REG1_REG_16__SCAN_IN), .Y(n7303));
  NAND2X1 g05663(.A(n7303), .B(n7297), .Y(n7304));
  INVX1   g05664(.A(n7304), .Y(n7305));
  OAI22X1 g05665(.A0(n7265), .A1(n6528), .B0(n6535), .B1(n7305), .Y(n7306));
  AOI21X1 g05666(.A0(n7296), .A1(n6532), .B0(n7306), .Y(n7307));
  OAI21X1 g05667(.A0(n7283), .A1(n6525), .B0(n7307), .Y(n7308));
  NOR2X1  g05668(.A(n7308), .B(n7291), .Y(n7309));
  NAND2X1 g05669(.A(n6465), .B(P2_REG0_REG_15__SCAN_IN), .Y(n7310));
  OAI21X1 g05670(.A0(n7309), .A1(n6465), .B0(n7310), .Y(P2_U3475));
  INVX1   g05671(.A(n7255), .Y(n7312));
  INVX1   g05672(.A(n7265), .Y(n7313));
  OAI21X1 g05673(.A0(n7313), .A1(n7312), .B0(n7275), .Y(n7314));
  NOR2X1  g05674(.A(n7265), .B(n7255), .Y(n7315));
  NOR2X1  g05675(.A(P2_IR_REG_31__SCAN_IN), .B(n6187), .Y(n7316));
  AOI21X1 g05676(.A0(n6198), .A1(P2_IR_REG_31__SCAN_IN), .B0(n7316), .Y(n7317));
  INVX1   g05677(.A(n7317), .Y(n7318));
  NOR2X1  g05678(.A(n6474), .B(n6186), .Y(n7319));
  AOI21X1 g05679(.A0(n7318), .A1(n6474), .B0(n7319), .Y(n7320));
  XOR2X1  g05680(.A(n7320), .B(n7304), .Y(n7321));
  NOR2X1  g05681(.A(n7321), .B(n7315), .Y(n7322));
  NOR2X1  g05682(.A(n7275), .B(n7315), .Y(n7323));
  INVX1   g05683(.A(n7323), .Y(n7324));
  NOR2X1  g05684(.A(n7320), .B(n7304), .Y(n7325));
  INVX1   g05685(.A(n7320), .Y(n7326));
  OAI22X1 g05686(.A0(n7305), .A1(n7326), .B0(n7313), .B1(n7312), .Y(n7327));
  NOR2X1  g05687(.A(n7327), .B(n7325), .Y(n7328));
  AOI22X1 g05688(.A0(n7324), .A1(n7328), .B0(n7322), .B1(n7314), .Y(n7329));
  INVX1   g05689(.A(n7329), .Y(n7330));
  NAND2X1 g05690(.A(n7330), .B(n6521), .Y(n7331));
  NOR2X1  g05691(.A(n7265), .B(n7312), .Y(n7333));
  INVX1   g05692(.A(n7333), .Y(n7334));
  NOR2X1  g05693(.A(n7313), .B(n7255), .Y(n7335));
  OAI21X1 g05694(.A0(n7335), .A1(n7282), .B0(n7334), .Y(n7336));
  XOR2X1  g05695(.A(n7320), .B(n7305), .Y(n7338));
  OAI22X1 g05696(.A0(n7312), .A1(n6634), .B0(n6633), .B1(n7350), .Y(n7341));
  AOI21X1 g05697(.A0(n6658), .A1(n6657), .B0(n7350), .Y(n7342));
  NOR2X1  g05698(.A(n7342), .B(n7341), .Y(n7343));
  AOI21X1 g05699(.A0(n6670), .A1(n6508), .B0(n7329), .Y(n7344));
  AOI21X1 g05700(.A0(n7330), .A1(n6512), .B0(n7344), .Y(n7345));
  NAND3X1 g05701(.A(n7345), .B(n7343), .C(n7331), .Y(n7346));
  INVX1   g05702(.A(n7335), .Y(n7347));
  AOI21X1 g05703(.A0(n7347), .A1(n7293), .B0(n7333), .Y(n7348));
  NOR2X1  g05704(.A(n7348), .B(n7338), .Y(n7349));
  AOI21X1 g05705(.A0(n7348), .A1(n7338), .B0(n7349), .Y(n7350));
  NOR3X1  g05706(.A(n7313), .B(n7247), .C(n7199), .Y(n7351));
  XOR2X1  g05707(.A(n7320), .B(n7351), .Y(n7352));
  INVX1   g05708(.A(P2_REG3_REG_17__SCAN_IN), .Y(n7353));
  NOR3X1  g05709(.A(n7251), .B(n7298), .C(n7299), .Y(n7354));
  XOR2X1  g05710(.A(n7354), .B(n7353), .Y(n7355));
  INVX1   g05711(.A(n7355), .Y(n7356));
  INVX1   g05712(.A(P2_REG1_REG_17__SCAN_IN), .Y(n7357));
  AOI22X1 g05713(.A0(n6556), .A1(P2_REG2_REG_17__SCAN_IN), .B0(P2_REG0_REG_17__SCAN_IN), .B1(n6557), .Y(n7358));
  OAI21X1 g05714(.A0(n6501), .A1(n7357), .B0(n7358), .Y(n7359));
  AOI21X1 g05715(.A0(n7356), .A1(n6502), .B0(n7359), .Y(n7360));
  OAI22X1 g05716(.A0(n7320), .A1(n6528), .B0(n6535), .B1(n7360), .Y(n7361));
  AOI21X1 g05717(.A0(n7352), .A1(n6532), .B0(n7361), .Y(n7362));
  OAI21X1 g05718(.A0(n7350), .A1(n6525), .B0(n7362), .Y(n7363));
  NOR2X1  g05719(.A(n7363), .B(n7346), .Y(n7364));
  NAND2X1 g05720(.A(n6465), .B(P2_REG0_REG_16__SCAN_IN), .Y(n7365));
  OAI21X1 g05721(.A0(n7364), .A1(n6465), .B0(n7365), .Y(P2_U3478));
  NOR2X1  g05722(.A(n7320), .B(n7305), .Y(n7367));
  INVX1   g05723(.A(n7360), .Y(n7368));
  NOR2X1  g05724(.A(P2_IR_REG_31__SCAN_IN), .B(n6204), .Y(n7369));
  AOI21X1 g05725(.A0(n6205), .A1(P2_IR_REG_31__SCAN_IN), .B0(n7369), .Y(n7370));
  INVX1   g05726(.A(n7370), .Y(n7371));
  NAND3X1 g05727(.A(n7371), .B(n6481), .C(n6480), .Y(n7372));
  OAI21X1 g05728(.A0(n6474), .A1(n6203), .B0(n7372), .Y(n7373));
  INVX1   g05729(.A(n7373), .Y(n7374));
  AOI22X1 g05730(.A0(n7360), .A1(n7374), .B0(n7320), .B1(n7305), .Y(n7375));
  INVX1   g05731(.A(n7375), .Y(n7376));
  AOI21X1 g05732(.A0(n7373), .A1(n7368), .B0(n7376), .Y(n7377));
  OAI21X1 g05733(.A0(n7367), .A1(n7336), .B0(n7377), .Y(n7378));
  XOR2X1  g05734(.A(n7373), .B(n7360), .Y(n7379));
  INVX1   g05735(.A(n7379), .Y(n7380));
  NOR2X1  g05736(.A(n7380), .B(n7367), .Y(n7381));
  INVX1   g05737(.A(n7381), .Y(n7382));
  OAI21X1 g05738(.A0(n7403), .A1(n7382), .B0(n7378), .Y(n7384));
  INVX1   g05739(.A(n7384), .Y(n7385));
  OAI21X1 g05740(.A0(n6520), .A1(n6514), .B0(n7385), .Y(n7386));
  NOR4X1  g05741(.A(n7315), .B(n7249), .C(n7207), .D(n7325), .Y(n7387));
  NOR2X1  g05742(.A(n7387), .B(n7327), .Y(n7388));
  NOR2X1  g05743(.A(n7388), .B(n7325), .Y(n7389));
  INVX1   g05744(.A(n7389), .Y(n7390));
  NOR3X1  g05745(.A(n7325), .B(n7315), .C(n7268), .Y(n7391));
  OAI21X1 g05746(.A0(n7221), .A1(n7220), .B0(n7391), .Y(n7392));
  NAND2X1 g05747(.A(n7392), .B(n7390), .Y(n7393));
  XOR2X1  g05748(.A(n7393), .B(n7380), .Y(n7394));
  NOR2X1  g05749(.A(n7394), .B(n6669), .Y(n7395));
  AOI21X1 g05750(.A0(n7385), .A1(n6518), .B0(n7395), .Y(n7396));
  OAI22X1 g05751(.A0(n7305), .A1(n6634), .B0(n6661), .B1(n7394), .Y(n7397));
  AOI21X1 g05752(.A0(n6670), .A1(n6508), .B0(n7394), .Y(n7398));
  NOR2X1  g05753(.A(n7398), .B(n7397), .Y(n7399));
  NAND3X1 g05754(.A(n7399), .B(n7396), .C(n7386), .Y(n7400));
  AOI21X1 g05755(.A0(n7320), .A1(n7305), .B0(n7348), .Y(n7403));
  NAND3X1 g05756(.A(n7320), .B(n7265), .C(n7295), .Y(n7405));
  XOR2X1  g05757(.A(n7373), .B(n7405), .Y(n7406));
  INVX1   g05758(.A(P2_REG3_REG_18__SCAN_IN), .Y(n7407));
  NOR4X1  g05759(.A(n7298), .B(n7353), .C(n7299), .D(n7251), .Y(n7408));
  XOR2X1  g05760(.A(n7408), .B(n7407), .Y(n7409));
  INVX1   g05761(.A(n7409), .Y(n7410));
  NAND2X1 g05762(.A(n6559), .B(P2_REG1_REG_18__SCAN_IN), .Y(n7411));
  AOI22X1 g05763(.A0(n6556), .A1(P2_REG2_REG_18__SCAN_IN), .B0(P2_REG0_REG_18__SCAN_IN), .B1(n6557), .Y(n7412));
  NAND2X1 g05764(.A(n7412), .B(n7411), .Y(n7413));
  AOI21X1 g05765(.A0(n7410), .A1(n6502), .B0(n7413), .Y(n7414));
  OAI22X1 g05766(.A0(n7374), .A1(n6528), .B0(n6535), .B1(n7414), .Y(n7415));
  AOI21X1 g05767(.A0(n7406), .A1(n6532), .B0(n7415), .Y(n7416));
  OAI21X1 g05768(.A0(n7384), .A1(n6525), .B0(n7416), .Y(n7417));
  NOR2X1  g05769(.A(n7417), .B(n7400), .Y(n7418));
  NAND2X1 g05770(.A(n6465), .B(P2_REG0_REG_17__SCAN_IN), .Y(n7419));
  OAI21X1 g05771(.A0(n7418), .A1(n6465), .B0(n7419), .Y(P2_U3481));
  NOR2X1  g05772(.A(P2_IR_REG_31__SCAN_IN), .B(n6211), .Y(n7421));
  AOI21X1 g05773(.A0(n6216), .A1(P2_IR_REG_31__SCAN_IN), .B0(n7421), .Y(n7422));
  INVX1   g05774(.A(n7422), .Y(n7423));
  NAND2X1 g05775(.A(n7423), .B(n6474), .Y(n7424));
  OAI21X1 g05776(.A0(n6474), .A1(n6210), .B0(n7424), .Y(n7425));
  XOR2X1  g05777(.A(n7425), .B(n7414), .Y(n7426));
  NAND2X1 g05778(.A(n7373), .B(n7367), .Y(n7428));
  OAI21X1 g05779(.A0(n7373), .A1(n7367), .B0(n7368), .Y(n7429));
  NAND2X1 g05780(.A(n7429), .B(n7428), .Y(n7430));
  AOI21X1 g05781(.A0(n7375), .A1(n7336), .B0(n7430), .Y(n7431));
  INVX1   g05782(.A(n7414), .Y(n7432));
  XOR2X1  g05783(.A(n7425), .B(n7432), .Y(n7433));
  NOR2X1  g05784(.A(n7433), .B(n7431), .Y(n7434));
  AOI21X1 g05785(.A0(n7431), .A1(n7433), .B0(n7434), .Y(n7435));
  INVX1   g05786(.A(n7435), .Y(n7436));
  AOI22X1 g05787(.A0(n7368), .A1(n6574), .B0(n6518), .B1(n7436), .Y(n7437));
  OAI21X1 g05788(.A0(n6520), .A1(n6514), .B0(n7436), .Y(n7438));
  NOR2X1  g05789(.A(n7373), .B(n7360), .Y(n7439));
  AOI22X1 g05790(.A0(n7390), .A1(n7392), .B0(n7373), .B1(n7360), .Y(n7440));
  NOR2X1  g05791(.A(n7440), .B(n7439), .Y(n7441));
  XOR2X1  g05792(.A(n7441), .B(n7426), .Y(n7442));
  INVX1   g05793(.A(n7442), .Y(n7443));
  OAI21X1 g05794(.A0(n6521), .A1(n6507), .B0(n7443), .Y(n7444));
  OAI21X1 g05795(.A0(n6516), .A1(n6512), .B0(n7443), .Y(n7445));
  NAND4X1 g05796(.A(n7444), .B(n7438), .C(n7437), .D(n7445), .Y(n7446));
  INVX1   g05797(.A(n7430), .Y(n7448));
  OAI21X1 g05798(.A0(n7376), .A1(n7348), .B0(n7448), .Y(n7449));
  NOR2X1  g05799(.A(n7435), .B(n6525), .Y(n7452));
  NOR2X1  g05800(.A(n7373), .B(n7405), .Y(n7453));
  INVX1   g05801(.A(n7425), .Y(n7454));
  NOR2X1  g05802(.A(n7454), .B(n7453), .Y(n7455));
  NOR3X1  g05803(.A(n7425), .B(n7373), .C(n7405), .Y(n7456));
  NOR3X1  g05804(.A(n7456), .B(n7455), .C(n6533), .Y(n7457));
  NAND2X1 g05805(.A(n7408), .B(P2_REG3_REG_18__SCAN_IN), .Y(n7458));
  XOR2X1  g05806(.A(n7458), .B(P2_REG3_REG_19__SCAN_IN), .Y(n7459));
  INVX1   g05807(.A(n7459), .Y(n7460));
  NAND2X1 g05808(.A(n6559), .B(P2_REG1_REG_19__SCAN_IN), .Y(n7461));
  AOI22X1 g05809(.A0(n6556), .A1(P2_REG2_REG_19__SCAN_IN), .B0(P2_REG0_REG_19__SCAN_IN), .B1(n6557), .Y(n7462));
  NAND2X1 g05810(.A(n7462), .B(n7461), .Y(n7463));
  AOI21X1 g05811(.A0(n7460), .A1(n6502), .B0(n7463), .Y(n7464));
  OAI22X1 g05812(.A0(n7454), .A1(n6528), .B0(n6535), .B1(n7464), .Y(n7465));
  NOR4X1  g05813(.A(n7457), .B(n7452), .C(n7446), .D(n7465), .Y(n7466));
  NAND2X1 g05814(.A(n6465), .B(P2_REG0_REG_18__SCAN_IN), .Y(n7467));
  OAI21X1 g05815(.A0(n7466), .A1(n6465), .B0(n7467), .Y(P2_U3484));
  NAND3X1 g05816(.A(n6481), .B(n6480), .C(n6513), .Y(n7469));
  OAI21X1 g05817(.A0(n6474), .A1(n6221), .B0(n7469), .Y(n7470));
  XOR2X1  g05818(.A(n7470), .B(n7464), .Y(n7471));
  INVX1   g05819(.A(n7439), .Y(n7472));
  INVX1   g05820(.A(n7391), .Y(n7473));
  AOI21X1 g05821(.A0(n7273), .A1(n7267), .B0(n7473), .Y(n7474));
  OAI22X1 g05822(.A0(n7389), .A1(n7474), .B0(n7374), .B1(n7368), .Y(n7475));
  AOI21X1 g05823(.A0(n7475), .A1(n7472), .B0(n7414), .Y(n7476));
  NAND3X1 g05824(.A(n7475), .B(n7414), .C(n7472), .Y(n7477));
  AOI21X1 g05825(.A0(n7477), .A1(n7454), .B0(n7476), .Y(n7478));
  XOR2X1  g05826(.A(n7478), .B(n7471), .Y(n7479));
  INVX1   g05827(.A(n7479), .Y(n7480));
  NAND2X1 g05828(.A(n7480), .B(n6521), .Y(n7481));
  NOR2X1  g05829(.A(n7425), .B(n7432), .Y(n7482));
  NAND2X1 g05830(.A(n7425), .B(n7432), .Y(n7483));
  OAI21X1 g05831(.A0(n7482), .A1(n7431), .B0(n7483), .Y(n7484));
  NOR2X1  g05832(.A(n7484), .B(n7471), .Y(n7485));
  INVX1   g05833(.A(n7464), .Y(n7486));
  XOR2X1  g05834(.A(n7470), .B(n7486), .Y(n7487));
  AOI21X1 g05835(.A0(n7471), .A1(n7484), .B0(n7485), .Y(n7489));
  OAI22X1 g05836(.A0(n7414), .A1(n6634), .B0(n6633), .B1(n7489), .Y(n7490));
  AOI21X1 g05837(.A0(n6658), .A1(n6657), .B0(n7489), .Y(n7491));
  NOR2X1  g05838(.A(n7491), .B(n7490), .Y(n7492));
  AOI21X1 g05839(.A0(n6670), .A1(n6508), .B0(n7479), .Y(n7493));
  AOI21X1 g05840(.A0(n7480), .A1(n6512), .B0(n7493), .Y(n7494));
  NAND3X1 g05841(.A(n7494), .B(n7492), .C(n7481), .Y(n7495));
  INVX1   g05842(.A(n7482), .Y(n7497));
  INVX1   g05843(.A(n7483), .Y(n7498));
  AOI21X1 g05844(.A0(n7449), .A1(n7497), .B0(n7498), .Y(n7499));
  NOR2X1  g05845(.A(n7499), .B(n7487), .Y(n7500));
  INVX1   g05846(.A(n7470), .Y(n7502));
  XOR2X1  g05847(.A(n7502), .B(n7456), .Y(n7503));
  NAND3X1 g05848(.A(n7408), .B(P2_REG3_REG_19__SCAN_IN), .C(P2_REG3_REG_18__SCAN_IN), .Y(n7504));
  XOR2X1  g05849(.A(n7504), .B(P2_REG3_REG_20__SCAN_IN), .Y(n7505));
  AOI22X1 g05850(.A0(n6556), .A1(P2_REG2_REG_20__SCAN_IN), .B0(P2_REG0_REG_20__SCAN_IN), .B1(n6557), .Y(n7506));
  INVX1   g05851(.A(n7506), .Y(n7507));
  AOI21X1 g05852(.A0(n6559), .A1(P2_REG1_REG_20__SCAN_IN), .B0(n7507), .Y(n7508));
  OAI21X1 g05853(.A0(n7505), .A1(n6503), .B0(n7508), .Y(n7509));
  INVX1   g05854(.A(n7509), .Y(n7510));
  OAI22X1 g05855(.A0(n7502), .A1(n6528), .B0(n6535), .B1(n7510), .Y(n7511));
  AOI21X1 g05856(.A0(n7503), .A1(n6532), .B0(n7511), .Y(n7512));
  OAI21X1 g05857(.A0(n7489), .A1(n6525), .B0(n7512), .Y(n7513));
  NOR2X1  g05858(.A(n7513), .B(n7495), .Y(n7514));
  NAND2X1 g05859(.A(n6465), .B(P2_REG0_REG_19__SCAN_IN), .Y(n7515));
  OAI21X1 g05860(.A0(n7514), .A1(n6465), .B0(n7515), .Y(P2_U3486));
  OAI21X1 g05861(.A0(n6227), .A1(n6225), .B0(n6750), .Y(n7517));
  NOR2X1  g05862(.A(n7502), .B(n7486), .Y(n7520));
  NOR2X1  g05863(.A(n7470), .B(n7464), .Y(n7521));
  INVX1   g05864(.A(n7521), .Y(n7522));
  OAI21X1 g05865(.A0(n7478), .A1(n7520), .B0(n7522), .Y(n7523));
  XOR2X1  g05866(.A(n7523), .B(n9398), .Y(n7524));
  INVX1   g05867(.A(n7524), .Y(n7525));
  NAND2X1 g05868(.A(n7525), .B(n6521), .Y(n7526));
  INVX1   g05869(.A(n7517), .Y(n7527));
  AOI22X1 g05870(.A0(n7510), .A1(n7517), .B0(n7502), .B1(n7464), .Y(n7528));
  INVX1   g05871(.A(n7528), .Y(n7529));
  AOI21X1 g05872(.A0(n7527), .A1(n7509), .B0(n7529), .Y(n7530));
  INVX1   g05873(.A(n7530), .Y(n7531));
  NAND2X1 g05874(.A(n7470), .B(n7486), .Y(n7532));
  INVX1   g05875(.A(n7532), .Y(n7533));
  NOR2X1  g05876(.A(n7533), .B(n7484), .Y(n7534));
  NOR2X1  g05877(.A(n7534), .B(n7531), .Y(n7535));
  NAND2X1 g05878(.A(n7502), .B(n7464), .Y(n7536));
  NOR2X1  g05879(.A(n9398), .B(n7533), .Y(n7537));
  INVX1   g05880(.A(n7537), .Y(n7538));
  AOI21X1 g05881(.A0(n7536), .A1(n7484), .B0(n7538), .Y(n7539));
  NOR2X1  g05882(.A(n7539), .B(n7535), .Y(n7540));
  AOI22X1 g05883(.A0(n7486), .A1(n6574), .B0(n6518), .B1(n7540), .Y(n7541));
  OAI21X1 g05884(.A0(n6520), .A1(n6514), .B0(n7540), .Y(n7542));
  AOI21X1 g05885(.A0(n6670), .A1(n6508), .B0(n7524), .Y(n7543));
  AOI21X1 g05886(.A0(n7525), .A1(n6512), .B0(n7543), .Y(n7544));
  NAND4X1 g05887(.A(n7542), .B(n7541), .C(n7526), .D(n7544), .Y(n7545));
  AOI21X1 g05888(.A0(n7502), .A1(n7464), .B0(n7499), .Y(n7548));
  OAI22X1 g05889(.A0(n7534), .A1(n7531), .B0(n7538), .B1(n7548), .Y(n7549));
  NAND2X1 g05890(.A(n7502), .B(n7456), .Y(n7550));
  XOR2X1  g05891(.A(n7527), .B(n7550), .Y(n7551));
  NAND4X1 g05892(.A(P2_REG3_REG_19__SCAN_IN), .B(P2_REG3_REG_20__SCAN_IN), .C(P2_REG3_REG_18__SCAN_IN), .D(n7408), .Y(n7552));
  XOR2X1  g05893(.A(n7552), .B(P2_REG3_REG_21__SCAN_IN), .Y(n7553));
  AOI22X1 g05894(.A0(n6556), .A1(P2_REG2_REG_21__SCAN_IN), .B0(P2_REG0_REG_21__SCAN_IN), .B1(n6557), .Y(n7554));
  INVX1   g05895(.A(n7554), .Y(n7555));
  AOI21X1 g05896(.A0(n6559), .A1(P2_REG1_REG_21__SCAN_IN), .B0(n7555), .Y(n7556));
  OAI21X1 g05897(.A0(n7553), .A1(n6503), .B0(n7556), .Y(n7557));
  INVX1   g05898(.A(n7557), .Y(n7558));
  OAI22X1 g05899(.A0(n7517), .A1(n6528), .B0(n6535), .B1(n7558), .Y(n7559));
  AOI21X1 g05900(.A0(n7551), .A1(n6532), .B0(n7559), .Y(n7560));
  OAI21X1 g05901(.A0(n7549), .A1(n6525), .B0(n7560), .Y(n7561));
  NOR2X1  g05902(.A(n7561), .B(n7545), .Y(n7562));
  NAND2X1 g05903(.A(n6465), .B(P2_REG0_REG_20__SCAN_IN), .Y(n7563));
  OAI21X1 g05904(.A0(n7562), .A1(n6465), .B0(n7563), .Y(P2_U3487));
  NOR2X1  g05905(.A(n6474), .B(n6236), .Y(n7565));
  XOR2X1  g05906(.A(n7565), .B(n7558), .Y(n7566));
  NOR2X1  g05907(.A(n7517), .B(n7509), .Y(n7567));
  INVX1   g05908(.A(n7567), .Y(n7568));
  NOR2X1  g05909(.A(n7527), .B(n7510), .Y(n7569));
  AOI21X1 g05910(.A0(n7523), .A1(n7568), .B0(n7569), .Y(n7570));
  XOR2X1  g05911(.A(n7570), .B(n7566), .Y(n7571));
  INVX1   g05912(.A(n7571), .Y(n7572));
  NAND2X1 g05913(.A(n7572), .B(n6521), .Y(n7573));
  NAND2X1 g05914(.A(n7528), .B(n7484), .Y(n7574));
  OAI21X1 g05915(.A0(n7517), .A1(n7532), .B0(n7510), .Y(n7575));
  OAI21X1 g05916(.A0(n7527), .A1(n7533), .B0(n7575), .Y(n7576));
  AOI21X1 g05917(.A0(n7574), .A1(n7576), .B0(n7566), .Y(n7577));
  INVX1   g05918(.A(n7576), .Y(n7579));
  NOR2X1  g05919(.A(n7579), .B(n9397), .Y(n7580));
  AOI21X1 g05920(.A0(n7580), .A1(n7574), .B0(n7577), .Y(n7581));
  AOI22X1 g05921(.A0(n7509), .A1(n6574), .B0(n6518), .B1(n7581), .Y(n7582));
  OAI21X1 g05922(.A0(n6520), .A1(n6514), .B0(n7581), .Y(n7583));
  NAND3X1 g05923(.A(n7583), .B(n7582), .C(n7573), .Y(n7584));
  NOR2X1  g05924(.A(n7571), .B(n6669), .Y(n7585));
  AOI21X1 g05925(.A0(n6670), .A1(n6508), .B0(n7571), .Y(n7586));
  AOI21X1 g05926(.A0(n7528), .A1(n7484), .B0(n7579), .Y(n7587));
  OAI21X1 g05927(.A0(n7529), .A1(n7499), .B0(n7580), .Y(n7588));
  OAI21X1 g05928(.A0(n7587), .A1(n7566), .B0(n7588), .Y(n7589));
  NAND3X1 g05929(.A(n7517), .B(n7502), .C(n7456), .Y(n7590));
  XOR2X1  g05930(.A(n7565), .B(n7590), .Y(n7591));
  INVX1   g05931(.A(n7565), .Y(n7592));
  INVX1   g05932(.A(P2_REG3_REG_22__SCAN_IN), .Y(n7593));
  INVX1   g05933(.A(P2_REG3_REG_21__SCAN_IN), .Y(n7594));
  NOR2X1  g05934(.A(n7552), .B(n7594), .Y(n7595));
  XOR2X1  g05935(.A(n7595), .B(n7593), .Y(n7596));
  AOI22X1 g05936(.A0(n6556), .A1(P2_REG2_REG_22__SCAN_IN), .B0(P2_REG0_REG_22__SCAN_IN), .B1(n6557), .Y(n7597));
  INVX1   g05937(.A(n7597), .Y(n7598));
  AOI21X1 g05938(.A0(n6559), .A1(P2_REG1_REG_22__SCAN_IN), .B0(n7598), .Y(n7599));
  OAI21X1 g05939(.A0(n7596), .A1(n6503), .B0(n7599), .Y(n7600));
  INVX1   g05940(.A(n7600), .Y(n7601));
  OAI22X1 g05941(.A0(n7592), .A1(n6528), .B0(n6535), .B1(n7601), .Y(n7602));
  AOI21X1 g05942(.A0(n7591), .A1(n6532), .B0(n7602), .Y(n7603));
  OAI21X1 g05943(.A0(n7589), .A1(n6525), .B0(n7603), .Y(n7604));
  NOR4X1  g05944(.A(n7586), .B(n7585), .C(n7584), .D(n7604), .Y(n7605));
  NAND2X1 g05945(.A(n6465), .B(P2_REG0_REG_21__SCAN_IN), .Y(n7606));
  OAI21X1 g05946(.A0(n7605), .A1(n6465), .B0(n7606), .Y(P2_U3488));
  NOR2X1  g05947(.A(n6474), .B(n6244), .Y(n7608));
  XOR2X1  g05948(.A(n7608), .B(n7601), .Y(n7609));
  NOR3X1  g05949(.A(n7557), .B(n6474), .C(n6236), .Y(n7611));
  OAI21X1 g05950(.A0(n6474), .A1(n6236), .B0(n7557), .Y(n7612));
  OAI21X1 g05951(.A0(n7570), .A1(n7611), .B0(n7612), .Y(n7613));
  XOR2X1  g05952(.A(n7613), .B(n9396), .Y(n7614));
  NOR2X1  g05953(.A(n7565), .B(n7557), .Y(n7615));
  INVX1   g05954(.A(n7615), .Y(n7616));
  OAI21X1 g05955(.A0(n7529), .A1(n7483), .B0(n7576), .Y(n7617));
  NOR3X1  g05956(.A(n7558), .B(n6474), .C(n6236), .Y(n7618));
  AOI21X1 g05957(.A0(n7617), .A1(n7616), .B0(n7618), .Y(n7619));
  NOR3X1  g05958(.A(n7615), .B(n7529), .C(n7482), .Y(n7620));
  INVX1   g05959(.A(n7620), .Y(n7621));
  OAI21X1 g05960(.A0(n7621), .A1(n7431), .B0(n7619), .Y(n7622));
  XOR2X1  g05961(.A(n7622), .B(n7609), .Y(n7623));
  OAI22X1 g05962(.A0(n7558), .A1(n6634), .B0(n6633), .B1(n7623), .Y(n7624));
  AOI21X1 g05963(.A0(n6658), .A1(n6657), .B0(n7623), .Y(n7625));
  NOR2X1  g05964(.A(n7625), .B(n7624), .Y(n7626));
  OAI21X1 g05965(.A0(n7614), .A1(n6661), .B0(n7626), .Y(n7627));
  NOR2X1  g05966(.A(n7614), .B(n6669), .Y(n7628));
  AOI21X1 g05967(.A0(n6670), .A1(n6508), .B0(n7614), .Y(n7629));
  INVX1   g05968(.A(n7619), .Y(n7630));
  AOI21X1 g05969(.A0(n7620), .A1(n7449), .B0(n7630), .Y(n7631));
  NAND4X1 g05970(.A(n7517), .B(n7502), .C(n7456), .D(n7592), .Y(n7633));
  XOR2X1  g05971(.A(n7608), .B(n7633), .Y(n7634));
  INVX1   g05972(.A(n7608), .Y(n7635));
  INVX1   g05973(.A(P2_REG3_REG_23__SCAN_IN), .Y(n7636));
  NOR3X1  g05974(.A(n7552), .B(n7594), .C(n7593), .Y(n7637));
  XOR2X1  g05975(.A(n7637), .B(n7636), .Y(n7638));
  AOI22X1 g05976(.A0(n6556), .A1(P2_REG2_REG_23__SCAN_IN), .B0(P2_REG0_REG_23__SCAN_IN), .B1(n6557), .Y(n7639));
  INVX1   g05977(.A(n7639), .Y(n7640));
  AOI21X1 g05978(.A0(n6559), .A1(P2_REG1_REG_23__SCAN_IN), .B0(n7640), .Y(n7641));
  OAI21X1 g05979(.A0(n7638), .A1(n6503), .B0(n7641), .Y(n7642));
  INVX1   g05980(.A(n7642), .Y(n7643));
  OAI22X1 g05981(.A0(n7635), .A1(n6528), .B0(n6535), .B1(n7643), .Y(n7644));
  AOI21X1 g05982(.A0(n7634), .A1(n6532), .B0(n7644), .Y(n7645));
  OAI21X1 g05983(.A0(n7623), .A1(n6525), .B0(n7645), .Y(n7646));
  NOR4X1  g05984(.A(n7629), .B(n7628), .C(n7627), .D(n7646), .Y(n7647));
  NAND2X1 g05985(.A(n6465), .B(P2_REG0_REG_22__SCAN_IN), .Y(n7648));
  OAI21X1 g05986(.A0(n7647), .A1(n6465), .B0(n7648), .Y(P2_U3489));
  NOR2X1  g05987(.A(n7608), .B(n7601), .Y(n7650));
  NOR3X1  g05988(.A(n7600), .B(n6474), .C(n6244), .Y(n7651));
  NOR2X1  g05989(.A(n6474), .B(n6252), .Y(n7652));
  XOR2X1  g05990(.A(n7652), .B(n7643), .Y(n7653));
  NOR2X1  g05991(.A(n7653), .B(n7651), .Y(n7654));
  OAI21X1 g05992(.A0(n7613), .A1(n7650), .B0(n7654), .Y(n7655));
  OAI21X1 g05993(.A0(n7635), .A1(n7600), .B0(n7613), .Y(n7656));
  NOR3X1  g05994(.A(n7642), .B(n6474), .C(n6252), .Y(n7657));
  OAI22X1 g05995(.A0(n7643), .A1(n7652), .B0(n7608), .B1(n7601), .Y(n7658));
  NOR2X1  g05996(.A(n7658), .B(n7657), .Y(n7659));
  NAND2X1 g05997(.A(n7659), .B(n7656), .Y(n7660));
  AOI21X1 g05998(.A0(n7660), .A1(n7655), .B0(n6661), .Y(n7661));
  INVX1   g05999(.A(n7653), .Y(n7662));
  NOR3X1  g06000(.A(n7601), .B(n6474), .C(n6244), .Y(n7663));
  OAI21X1 g06001(.A0(n6474), .A1(n6244), .B0(n7601), .Y(n7664));
  AOI21X1 g06002(.A0(n7664), .A1(n7622), .B0(n7663), .Y(n7665));
  XOR2X1  g06003(.A(n7665), .B(n7662), .Y(n7666));
  OAI22X1 g06004(.A0(n7601), .A1(n6634), .B0(n6633), .B1(n7666), .Y(n7667));
  AOI21X1 g06005(.A0(n6658), .A1(n6657), .B0(n7666), .Y(n7668));
  NOR2X1  g06006(.A(n7668), .B(n7667), .Y(n7669));
  INVX1   g06007(.A(n7669), .Y(n7670));
  AOI21X1 g06008(.A0(n7660), .A1(n7655), .B0(n6669), .Y(n7671));
  AOI22X1 g06009(.A0(n7655), .A1(n7660), .B0(n6670), .B1(n6508), .Y(n7672));
  NOR4X1  g06010(.A(n7671), .B(n7670), .C(n7661), .D(n7672), .Y(n7673));
  INVX1   g06011(.A(n7673), .Y(n7674));
  INVX1   g06012(.A(n7663), .Y(n7675));
  INVX1   g06013(.A(n7664), .Y(n7676));
  OAI21X1 g06014(.A0(n7676), .A1(n7631), .B0(n7675), .Y(n7677));
  NOR2X1  g06015(.A(n7666), .B(n6525), .Y(n7679));
  NOR3X1  g06016(.A(n7608), .B(n7565), .C(n7590), .Y(n7680));
  XOR2X1  g06017(.A(n7652), .B(n7680), .Y(n7681));
  NOR4X1  g06018(.A(n7636), .B(n7594), .C(n7593), .D(n7552), .Y(n7682));
  XOR2X1  g06019(.A(n7682), .B(P2_REG3_REG_24__SCAN_IN), .Y(n7683));
  INVX1   g06020(.A(n7683), .Y(n7684));
  AOI22X1 g06021(.A0(n6556), .A1(P2_REG2_REG_24__SCAN_IN), .B0(P2_REG0_REG_24__SCAN_IN), .B1(n6557), .Y(n7685));
  INVX1   g06022(.A(n7685), .Y(n7686));
  AOI21X1 g06023(.A0(n6559), .A1(P2_REG1_REG_24__SCAN_IN), .B0(n7686), .Y(n7687));
  OAI21X1 g06024(.A0(n7684), .A1(n6503), .B0(n7687), .Y(n7688));
  AOI22X1 g06025(.A0(n7652), .A1(n6529), .B0(n6534), .B1(n7688), .Y(n7689));
  OAI21X1 g06026(.A0(n7681), .A1(n6533), .B0(n7689), .Y(n7690));
  NOR3X1  g06027(.A(n7690), .B(n7679), .C(n7674), .Y(n7691));
  NAND2X1 g06028(.A(n6465), .B(P2_REG0_REG_23__SCAN_IN), .Y(n7692));
  OAI21X1 g06029(.A0(n7691), .A1(n6465), .B0(n7692), .Y(P2_U3490));
  INVX1   g06030(.A(n7688), .Y(n7694));
  NOR2X1  g06031(.A(n6474), .B(n6261), .Y(n7695));
  XOR2X1  g06032(.A(n7695), .B(n7694), .Y(n7696));
  NOR3X1  g06033(.A(n7657), .B(n7651), .C(n7612), .Y(n7698));
  NOR2X1  g06034(.A(n7698), .B(n7658), .Y(n7699));
  NOR3X1  g06035(.A(n7657), .B(n7651), .C(n7611), .Y(n7700));
  INVX1   g06036(.A(n7700), .Y(n7701));
  OAI22X1 g06037(.A0(n7699), .A1(n7657), .B0(n7570), .B1(n7701), .Y(n7702));
  XOR2X1  g06038(.A(n7702), .B(n7724), .Y(n7703));
  INVX1   g06039(.A(n7703), .Y(n7704));
  NAND2X1 g06040(.A(n7704), .B(n6521), .Y(n7705));
  NOR3X1  g06041(.A(n7643), .B(n6474), .C(n6252), .Y(n7706));
  INVX1   g06042(.A(n7706), .Y(n7707));
  OAI21X1 g06043(.A0(n6474), .A1(n6252), .B0(n7643), .Y(n7708));
  INVX1   g06044(.A(n7708), .Y(n7709));
  OAI21X1 g06045(.A0(n7709), .A1(n7665), .B0(n7707), .Y(n7710));
  OAI21X1 g06046(.A0(n6474), .A1(n6261), .B0(n7694), .Y(n7711));
  INVX1   g06047(.A(n7711), .Y(n7712));
  NOR3X1  g06048(.A(n7694), .B(n6474), .C(n6261), .Y(n7713));
  OAI21X1 g06049(.A0(n7713), .A1(n7712), .B0(n7710), .Y(n7714));
  OAI21X1 g06050(.A0(n7710), .A1(n7696), .B0(n7714), .Y(n7715));
  AOI22X1 g06051(.A0(n7642), .A1(n6574), .B0(n6518), .B1(n7715), .Y(n7716));
  OAI21X1 g06052(.A0(n6520), .A1(n6514), .B0(n7715), .Y(n7717));
  NAND3X1 g06053(.A(n7717), .B(n7716), .C(n7705), .Y(n7718));
  NOR2X1  g06054(.A(n7703), .B(n6669), .Y(n7719));
  AOI21X1 g06055(.A0(n6670), .A1(n6508), .B0(n7703), .Y(n7720));
  AOI21X1 g06056(.A0(n7708), .A1(n7677), .B0(n7706), .Y(n7721));
  NOR2X1  g06057(.A(n3861), .B(n1790), .Y(n7722));
  OAI21X1 g06058(.A0(n6260), .A1(n7722), .B0(n6750), .Y(n7723));
  XOR2X1  g06059(.A(n7723), .B(n7694), .Y(n7724));
  NOR2X1  g06060(.A(n7721), .B(n7724), .Y(n7725));
  AOI21X1 g06061(.A0(n7721), .A1(n7724), .B0(n7725), .Y(n7726));
  NOR3X1  g06062(.A(n7652), .B(n7608), .C(n7633), .Y(n7727));
  XOR2X1  g06063(.A(n7723), .B(n7727), .Y(n7728));
  NAND2X1 g06064(.A(n7682), .B(P2_REG3_REG_24__SCAN_IN), .Y(n7729));
  XOR2X1  g06065(.A(n7729), .B(P2_REG3_REG_25__SCAN_IN), .Y(n7730));
  AOI22X1 g06066(.A0(n6556), .A1(P2_REG2_REG_25__SCAN_IN), .B0(P2_REG0_REG_25__SCAN_IN), .B1(n6557), .Y(n7731));
  INVX1   g06067(.A(n7731), .Y(n7732));
  AOI21X1 g06068(.A0(n6559), .A1(P2_REG1_REG_25__SCAN_IN), .B0(n7732), .Y(n7733));
  OAI21X1 g06069(.A0(n7730), .A1(n6503), .B0(n7733), .Y(n7734));
  INVX1   g06070(.A(n7734), .Y(n7735));
  OAI22X1 g06071(.A0(n7723), .A1(n6528), .B0(n6535), .B1(n7735), .Y(n7736));
  AOI21X1 g06072(.A0(n7728), .A1(n6532), .B0(n7736), .Y(n7737));
  OAI21X1 g06073(.A0(n7726), .A1(n6525), .B0(n7737), .Y(n7738));
  NOR4X1  g06074(.A(n7720), .B(n7719), .C(n7718), .D(n7738), .Y(n7739));
  NAND2X1 g06075(.A(n6465), .B(P2_REG0_REG_24__SCAN_IN), .Y(n7740));
  OAI21X1 g06076(.A0(n7739), .A1(n6465), .B0(n7740), .Y(P2_U3491));
  NOR2X1  g06077(.A(n6474), .B(n6268), .Y(n7742));
  XOR2X1  g06078(.A(n7742), .B(n7735), .Y(n7743));
  NOR3X1  g06079(.A(n7688), .B(n6474), .C(n6261), .Y(n7744));
  INVX1   g06080(.A(n7744), .Y(n7745));
  OAI21X1 g06081(.A0(n6474), .A1(n6261), .B0(n7688), .Y(n7746));
  INVX1   g06082(.A(n7746), .Y(n7747));
  AOI21X1 g06083(.A0(n7702), .A1(n7745), .B0(n7747), .Y(n7748));
  XOR2X1  g06084(.A(n7748), .B(n7743), .Y(n7749));
  NOR2X1  g06085(.A(n7749), .B(n6661), .Y(n7750));
  INVX1   g06086(.A(n7750), .Y(n7751));
  AOI21X1 g06087(.A0(n7711), .A1(n7710), .B0(n7713), .Y(n7752));
  NOR3X1  g06088(.A(n7734), .B(n6474), .C(n6268), .Y(n7753));
  OAI21X1 g06089(.A0(n6474), .A1(n6268), .B0(n7734), .Y(n7754));
  INVX1   g06090(.A(n7754), .Y(n7755));
  OAI21X1 g06091(.A0(n7755), .A1(n7753), .B0(n7752), .Y(n7756));
  NOR2X1  g06092(.A(n3913), .B(n1790), .Y(n7757));
  OAI21X1 g06093(.A0(n6267), .A1(n7757), .B0(n6750), .Y(n7758));
  XOR2X1  g06094(.A(n7758), .B(n7735), .Y(n7759));
  OAI21X1 g06095(.A0(n7759), .A1(n7752), .B0(n7756), .Y(n7760));
  AOI22X1 g06096(.A0(n7688), .A1(n6574), .B0(n6518), .B1(n7760), .Y(n7761));
  OAI21X1 g06097(.A0(n6520), .A1(n6514), .B0(n7760), .Y(n7762));
  NAND3X1 g06098(.A(n7762), .B(n7761), .C(n7751), .Y(n7763));
  INVX1   g06099(.A(n7749), .Y(n7764));
  OAI21X1 g06100(.A0(n6516), .A1(n6507), .B0(n7764), .Y(n7765));
  OAI21X1 g06101(.A0(n7749), .A1(n6669), .B0(n7765), .Y(n7766));
  INVX1   g06102(.A(n7713), .Y(n7768));
  OAI21X1 g06103(.A0(n7721), .A1(n7712), .B0(n7768), .Y(n7769));
  NOR2X1  g06104(.A(n7769), .B(n7743), .Y(n7770));
  AOI21X1 g06105(.A0(n7769), .A1(n7743), .B0(n7770), .Y(n7771));
  NOR4X1  g06106(.A(n7652), .B(n7608), .C(n7633), .D(n7695), .Y(n7772));
  XOR2X1  g06107(.A(n7758), .B(n7772), .Y(n7773));
  NAND3X1 g06108(.A(n7682), .B(P2_REG3_REG_25__SCAN_IN), .C(P2_REG3_REG_24__SCAN_IN), .Y(n7774));
  XOR2X1  g06109(.A(n7774), .B(P2_REG3_REG_26__SCAN_IN), .Y(n7775));
  AOI22X1 g06110(.A0(n6556), .A1(P2_REG2_REG_26__SCAN_IN), .B0(P2_REG0_REG_26__SCAN_IN), .B1(n6557), .Y(n7776));
  INVX1   g06111(.A(n7776), .Y(n7777));
  AOI21X1 g06112(.A0(n6559), .A1(P2_REG1_REG_26__SCAN_IN), .B0(n7777), .Y(n7778));
  OAI21X1 g06113(.A0(n7775), .A1(n6503), .B0(n7778), .Y(n7779));
  INVX1   g06114(.A(n7779), .Y(n7780));
  OAI22X1 g06115(.A0(n7758), .A1(n6528), .B0(n6535), .B1(n7780), .Y(n7781));
  AOI21X1 g06116(.A0(n7773), .A1(n6532), .B0(n7781), .Y(n7782));
  OAI21X1 g06117(.A0(n7771), .A1(n6525), .B0(n7782), .Y(n7783));
  NOR3X1  g06118(.A(n7783), .B(n7766), .C(n7763), .Y(n7784));
  NAND2X1 g06119(.A(n6465), .B(P2_REG0_REG_25__SCAN_IN), .Y(n7785));
  OAI21X1 g06120(.A0(n7784), .A1(n6465), .B0(n7785), .Y(P2_U3492));
  OAI21X1 g06121(.A0(n6275), .A1(n6273), .B0(n6750), .Y(n7787));
  XOR2X1  g06122(.A(n7787), .B(n7779), .Y(n7788));
  OAI21X1 g06123(.A0(n7748), .A1(n7753), .B0(n7754), .Y(n7789));
  XOR2X1  g06124(.A(n7789), .B(n7788), .Y(n7790));
  INVX1   g06125(.A(n7790), .Y(n7791));
  NOR3X1  g06126(.A(n7735), .B(n6474), .C(n6268), .Y(n7795));
  AOI22X1 g06127(.A0(n7780), .A1(n7787), .B0(n7758), .B1(n7735), .Y(n7796));
  OAI21X1 g06128(.A0(n7787), .A1(n7780), .B0(n7796), .Y(n7797));
  INVX1   g06129(.A(n7797), .Y(n7798));
  NOR2X1  g06130(.A(n7742), .B(n7734), .Y(n7800));
  INVX1   g06131(.A(n7795), .Y(n7801));
  NAND2X1 g06132(.A(n7788), .B(n7801), .Y(n7802));
  INVX1   g06133(.A(n7802), .Y(n7803));
  OAI21X1 g06134(.A0(n7800), .A1(n7752), .B0(n7803), .Y(n7804));
  NAND2X1 g06135(.A(n7804), .B(n7812), .Y(n7805));
  OAI22X1 g06136(.A0(n7735), .A1(n6634), .B0(n6633), .B1(n7805), .Y(n7806));
  AOI21X1 g06137(.A0(n6658), .A1(n6657), .B0(n7805), .Y(n7807));
  NOR2X1  g06138(.A(n7807), .B(n7806), .Y(n7808));
  OAI21X1 g06139(.A0(n7791), .A1(n6661), .B0(n7808), .Y(n7809));
  OAI21X1 g06140(.A0(n6516), .A1(n6507), .B0(n7790), .Y(n7810));
  OAI21X1 g06141(.A0(n7791), .A1(n6669), .B0(n7810), .Y(n7811));
  OAI21X1 g06142(.A0(n7769), .A1(n7795), .B0(n7798), .Y(n7812));
  NAND3X1 g06143(.A(n7804), .B(n7812), .C(n6524), .Y(n7815));
  NAND2X1 g06144(.A(n7758), .B(n7772), .Y(n7816));
  NOR2X1  g06145(.A(n6474), .B(n6276), .Y(n7817));
  XOR2X1  g06146(.A(n7817), .B(n7816), .Y(n7818));
  NAND4X1 g06147(.A(P2_REG3_REG_25__SCAN_IN), .B(P2_REG3_REG_24__SCAN_IN), .C(P2_REG3_REG_26__SCAN_IN), .D(n7682), .Y(n7819));
  XOR2X1  g06148(.A(n7819), .B(P2_REG3_REG_27__SCAN_IN), .Y(n7820));
  AOI22X1 g06149(.A0(n6556), .A1(P2_REG2_REG_27__SCAN_IN), .B0(P2_REG0_REG_27__SCAN_IN), .B1(n6557), .Y(n7821));
  INVX1   g06150(.A(n7821), .Y(n7822));
  AOI21X1 g06151(.A0(n6559), .A1(P2_REG1_REG_27__SCAN_IN), .B0(n7822), .Y(n7823));
  OAI21X1 g06152(.A0(n7820), .A1(n6503), .B0(n7823), .Y(n7824));
  INVX1   g06153(.A(n7824), .Y(n7825));
  OAI22X1 g06154(.A0(n7787), .A1(n6528), .B0(n6535), .B1(n7825), .Y(n7826));
  AOI21X1 g06155(.A0(n7818), .A1(n6532), .B0(n7826), .Y(n7827));
  NAND2X1 g06156(.A(n7827), .B(n7815), .Y(n7828));
  NOR3X1  g06157(.A(n7828), .B(n7811), .C(n7809), .Y(n7829));
  NAND2X1 g06158(.A(n6465), .B(P2_REG0_REG_26__SCAN_IN), .Y(n7830));
  OAI21X1 g06159(.A0(n7829), .A1(n6465), .B0(n7830), .Y(P2_U3493));
  NOR2X1  g06160(.A(n7817), .B(n7780), .Y(n7832));
  INVX1   g06161(.A(n7832), .Y(n7833));
  INVX1   g06162(.A(n7753), .Y(n7834));
  INVX1   g06163(.A(n7569), .Y(n7835));
  INVX1   g06164(.A(n7520), .Y(n7836));
  OAI21X1 g06165(.A0(n7440), .A1(n7439), .B0(n7432), .Y(n7837));
  NOR3X1  g06166(.A(n7440), .B(n7432), .C(n7439), .Y(n7838));
  OAI21X1 g06167(.A0(n7838), .A1(n7425), .B0(n7837), .Y(n7839));
  AOI21X1 g06168(.A0(n7839), .A1(n7836), .B0(n7521), .Y(n7840));
  OAI21X1 g06169(.A0(n7840), .A1(n7567), .B0(n7835), .Y(n7841));
  NOR2X1  g06170(.A(n7699), .B(n7657), .Y(n7842));
  AOI21X1 g06171(.A0(n7700), .A1(n7841), .B0(n7842), .Y(n7843));
  OAI21X1 g06172(.A0(n7843), .A1(n7744), .B0(n7746), .Y(n7844));
  AOI21X1 g06173(.A0(n7844), .A1(n7834), .B0(n7755), .Y(n7845));
  NOR2X1  g06174(.A(n7787), .B(n7779), .Y(n7846));
  INVX1   g06175(.A(n7846), .Y(n7847));
  OAI21X1 g06176(.A0(n6296), .A1(n6294), .B0(n6750), .Y(n7848));
  XOR2X1  g06177(.A(n7848), .B(n7824), .Y(n7849));
  INVX1   g06178(.A(n7849), .Y(n7850));
  NAND2X1 g06179(.A(n7850), .B(n7847), .Y(n7851));
  AOI21X1 g06180(.A0(n7845), .A1(n7833), .B0(n7851), .Y(n7852));
  OAI21X1 g06181(.A0(n7817), .A1(n7780), .B0(n7849), .Y(n7853));
  AOI21X1 g06182(.A0(n7789), .A1(n7847), .B0(n7853), .Y(n7854));
  OAI21X1 g06183(.A0(n7854), .A1(n7852), .B0(n6521), .Y(n7855));
  NAND2X1 g06184(.A(n7817), .B(n7779), .Y(n7856));
  OAI21X1 g06185(.A0(n7795), .A1(n7713), .B0(n7796), .Y(n7857));
  NAND3X1 g06186(.A(n7796), .B(n7711), .C(n7710), .Y(n7858));
  NAND3X1 g06187(.A(n7858), .B(n7857), .C(n7856), .Y(n7859));
  XOR2X1  g06188(.A(n7859), .B(n7850), .Y(n7860));
  NAND2X1 g06189(.A(n7860), .B(n6518), .Y(n7861));
  NOR2X1  g06190(.A(n7780), .B(n6634), .Y(n7862));
  INVX1   g06191(.A(n7862), .Y(n7863));
  OAI21X1 g06192(.A0(n6520), .A1(n6514), .B0(n7860), .Y(n7864));
  NAND4X1 g06193(.A(n7863), .B(n7861), .C(n7855), .D(n7864), .Y(n7865));
  OAI21X1 g06194(.A0(n7854), .A1(n7852), .B0(n6512), .Y(n7866));
  OAI22X1 g06195(.A0(n7852), .A1(n7854), .B0(n6516), .B1(n6507), .Y(n7867));
  NAND2X1 g06196(.A(n7867), .B(n7866), .Y(n7868));
  INVX1   g06197(.A(n7856), .Y(n7869));
  INVX1   g06198(.A(n7857), .Y(n7870));
  INVX1   g06199(.A(n7796), .Y(n7871));
  NOR3X1  g06200(.A(n7871), .B(n7721), .C(n7712), .Y(n7872));
  NOR3X1  g06201(.A(n7872), .B(n7870), .C(n7869), .Y(n7873));
  XOR2X1  g06202(.A(n7873), .B(n7850), .Y(n7874));
  NAND3X1 g06203(.A(n7787), .B(n7758), .C(n7772), .Y(n7875));
  NOR2X1  g06204(.A(n6474), .B(n6297), .Y(n7876));
  XOR2X1  g06205(.A(n7876), .B(n7875), .Y(n7877));
  INVX1   g06206(.A(P2_REG3_REG_28__SCAN_IN), .Y(n7878));
  INVX1   g06207(.A(P2_REG3_REG_27__SCAN_IN), .Y(n7879));
  NOR2X1  g06208(.A(n7819), .B(n7879), .Y(n7880));
  XOR2X1  g06209(.A(n7880), .B(n7878), .Y(n7881));
  AOI22X1 g06210(.A0(n6556), .A1(P2_REG2_REG_28__SCAN_IN), .B0(P2_REG0_REG_28__SCAN_IN), .B1(n6557), .Y(n7882));
  INVX1   g06211(.A(n7882), .Y(n7883));
  AOI21X1 g06212(.A0(n6559), .A1(P2_REG1_REG_28__SCAN_IN), .B0(n7883), .Y(n7884));
  OAI21X1 g06213(.A0(n7881), .A1(n6503), .B0(n7884), .Y(n7885));
  INVX1   g06214(.A(n7885), .Y(n7886));
  OAI22X1 g06215(.A0(n7848), .A1(n6528), .B0(n6535), .B1(n7886), .Y(n7887));
  AOI21X1 g06216(.A0(n7877), .A1(n6532), .B0(n7887), .Y(n7888));
  OAI21X1 g06217(.A0(n7874), .A1(n6525), .B0(n7888), .Y(n7889));
  NOR3X1  g06218(.A(n7889), .B(n7868), .C(n7865), .Y(n7890));
  NAND2X1 g06219(.A(n6465), .B(P2_REG0_REG_27__SCAN_IN), .Y(n7891));
  OAI21X1 g06220(.A0(n7890), .A1(n6465), .B0(n7891), .Y(P2_U3494));
  NOR2X1  g06221(.A(n6474), .B(n6304), .Y(n7893));
  XOR2X1  g06222(.A(n7893), .B(n7886), .Y(n7894));
  NOR2X1  g06223(.A(n7848), .B(n7824), .Y(n7895));
  NOR3X1  g06224(.A(n7895), .B(n7845), .C(n7846), .Y(n7896));
  OAI21X1 g06225(.A0(n7824), .A1(n7832), .B0(n7848), .Y(n7897));
  NAND3X1 g06226(.A(n7824), .B(n7787), .C(n7779), .Y(n7898));
  NAND2X1 g06227(.A(n7898), .B(n7897), .Y(n7899));
  NOR2X1  g06228(.A(n7899), .B(n7896), .Y(n7900));
  XOR2X1  g06229(.A(n7900), .B(n7894), .Y(n7901));
  AOI21X1 g06230(.A0(n7848), .A1(n7825), .B0(n7857), .Y(n7902));
  NOR2X1  g06231(.A(n7848), .B(n7825), .Y(n7903));
  AOI21X1 g06232(.A0(n7848), .A1(n7825), .B0(n7856), .Y(n7904));
  NOR3X1  g06233(.A(n7904), .B(n7903), .C(n7902), .Y(n7905));
  NAND2X1 g06234(.A(n7848), .B(n7825), .Y(n7906));
  NAND4X1 g06235(.A(n7796), .B(n7711), .C(n7710), .D(n7906), .Y(n7907));
  NAND2X1 g06236(.A(n7907), .B(n7905), .Y(n7908));
  XOR2X1  g06237(.A(n7908), .B(n7894), .Y(n7909));
  OAI22X1 g06238(.A0(n7825), .A1(n6634), .B0(n6633), .B1(n7909), .Y(n7910));
  AOI21X1 g06239(.A0(n6658), .A1(n6657), .B0(n7909), .Y(n7911));
  NOR2X1  g06240(.A(n7911), .B(n7910), .Y(n7912));
  OAI21X1 g06241(.A0(n7901), .A1(n6661), .B0(n7912), .Y(n7913));
  NOR2X1  g06242(.A(n7901), .B(n6669), .Y(n7914));
  AOI21X1 g06243(.A0(n6670), .A1(n6508), .B0(n7901), .Y(n7915));
  NAND2X1 g06244(.A(n7906), .B(n7711), .Y(n7916));
  NOR3X1  g06245(.A(n7916), .B(n7871), .C(n7721), .Y(n7917));
  NOR4X1  g06246(.A(n7904), .B(n7903), .C(n7902), .D(n7917), .Y(n7918));
  XOR2X1  g06247(.A(n7918), .B(n7894), .Y(n7919));
  NAND2X1 g06248(.A(n7919), .B(n6524), .Y(n7920));
  NOR2X1  g06249(.A(n7876), .B(n7875), .Y(n7921));
  OAI21X1 g06250(.A0(n4030), .A1(n4028), .B0(n1837), .Y(n7922));
  OAI21X1 g06251(.A0(n1837), .A1(n6302), .B0(n7922), .Y(n7923));
  NAND2X1 g06252(.A(n6750), .B(n7923), .Y(n7924));
  XOR2X1  g06253(.A(n7924), .B(n7921), .Y(n7925));
  NOR3X1  g06254(.A(n7819), .B(n7879), .C(n7878), .Y(n7926));
  INVX1   g06255(.A(n7926), .Y(n7927));
  AOI22X1 g06256(.A0(n6556), .A1(P2_REG2_REG_29__SCAN_IN), .B0(P2_REG1_REG_29__SCAN_IN), .B1(n6559), .Y(n7928));
  INVX1   g06257(.A(n7928), .Y(n7929));
  AOI21X1 g06258(.A0(n6557), .A1(P2_REG0_REG_29__SCAN_IN), .B0(n7929), .Y(n7930));
  OAI21X1 g06259(.A0(n7927), .A1(n6503), .B0(n7930), .Y(n7931));
  INVX1   g06260(.A(n7931), .Y(n7932));
  OAI22X1 g06261(.A0(n7924), .A1(n6528), .B0(n6535), .B1(n7932), .Y(n7933));
  AOI21X1 g06262(.A0(n7925), .A1(n6532), .B0(n7933), .Y(n7934));
  NAND2X1 g06263(.A(n7934), .B(n7920), .Y(n7935));
  NOR4X1  g06264(.A(n7915), .B(n7914), .C(n7913), .D(n7935), .Y(n7936));
  NAND2X1 g06265(.A(n6465), .B(P2_REG0_REG_28__SCAN_IN), .Y(n7937));
  OAI21X1 g06266(.A0(n7936), .A1(n6465), .B0(n7937), .Y(P2_U3495));
  AOI21X1 g06267(.A0(n2482), .A1(n2477), .B0(n1790), .Y(n7939));
  AOI21X1 g06268(.A0(n1789), .A1(n1786), .B0(n6312), .Y(n7940));
  OAI21X1 g06269(.A0(n7940), .A1(n7939), .B0(n6750), .Y(n7941));
  XOR2X1  g06270(.A(n7941), .B(n7931), .Y(n7942));
  INVX1   g06271(.A(n7942), .Y(n7943));
  AOI21X1 g06272(.A0(n7907), .A1(n7905), .B0(n7924), .Y(n7944));
  INVX1   g06273(.A(n7944), .Y(n7945));
  OAI21X1 g06274(.A0(n7908), .A1(n7893), .B0(n7885), .Y(n7946));
  NAND2X1 g06275(.A(n7946), .B(n7945), .Y(n7947));
  XOR2X1  g06276(.A(n7947), .B(n7943), .Y(n7948));
  NOR2X1  g06277(.A(n6455), .B(n6449), .Y(n7949));
  NOR2X1  g06278(.A(n6473), .B(P2_B_REG_SCAN_IN), .Y(n7950));
  OAI21X1 g06279(.A0(n7950), .A1(n6474), .B0(n7949), .Y(n7951));
  AOI22X1 g06280(.A0(n6556), .A1(P2_REG2_REG_30__SCAN_IN), .B0(P2_REG0_REG_30__SCAN_IN), .B1(n6557), .Y(n7952));
  INVX1   g06281(.A(n7952), .Y(n7953));
  AOI21X1 g06282(.A0(n6559), .A1(P2_REG1_REG_30__SCAN_IN), .B0(n7953), .Y(n7954));
  OAI22X1 g06283(.A0(n7951), .A1(n7954), .B0(n7886), .B1(n6634), .Y(n7955));
  AOI21X1 g06284(.A0(n7948), .A1(n6518), .B0(n7955), .Y(n7956));
  NOR2X1  g06285(.A(n7947), .B(n7942), .Y(n7957));
  AOI21X1 g06286(.A0(n7946), .A1(n7945), .B0(n7943), .Y(n7958));
  OAI22X1 g06287(.A0(n7957), .A1(n7958), .B0(n6520), .B1(n6514), .Y(n7959));
  NAND2X1 g06288(.A(n7959), .B(n7956), .Y(n7960));
  OAI21X1 g06289(.A0(n6474), .A1(n6304), .B0(n7885), .Y(n7961));
  INVX1   g06290(.A(n7895), .Y(n7962));
  NAND3X1 g06291(.A(n7962), .B(n7789), .C(n7847), .Y(n7963));
  NAND4X1 g06292(.A(n7897), .B(n7963), .C(n7961), .D(n7898), .Y(n7964));
  AOI21X1 g06293(.A0(n7893), .A1(n7886), .B0(n7942), .Y(n7965));
  OAI22X1 g06294(.A0(n7896), .A1(n7899), .B0(n7924), .B1(n7885), .Y(n7966));
  AOI21X1 g06295(.A0(n7924), .A1(n7885), .B0(n7943), .Y(n7967));
  AOI22X1 g06296(.A0(n7966), .A1(n7967), .B0(n7965), .B1(n7964), .Y(n7968));
  AOI21X1 g06297(.A0(n6661), .A1(n6508), .B0(n7968), .Y(n7969));
  AOI21X1 g06298(.A0(n6670), .A1(n6669), .B0(n7968), .Y(n7970));
  AOI21X1 g06299(.A0(n7918), .A1(n7924), .B0(n7886), .Y(n7972));
  NOR2X1  g06300(.A(n7972), .B(n7944), .Y(n7973));
  XOR2X1  g06301(.A(n7973), .B(n7943), .Y(n7974));
  INVX1   g06302(.A(n7941), .Y(n7975));
  NAND2X1 g06303(.A(n7924), .B(n7921), .Y(n7976));
  XOR2X1  g06304(.A(n7975), .B(n7976), .Y(n7977));
  AOI22X1 g06305(.A0(n7975), .A1(n6529), .B0(n6532), .B1(n7977), .Y(n7978));
  OAI21X1 g06306(.A0(n7974), .A1(n6525), .B0(n7978), .Y(n7979));
  NOR4X1  g06307(.A(n7970), .B(n7969), .C(n7960), .D(n7979), .Y(n7980));
  NAND2X1 g06308(.A(n6465), .B(P2_REG0_REG_29__SCAN_IN), .Y(n7981));
  OAI21X1 g06309(.A0(n7980), .A1(n6465), .B0(n7981), .Y(P2_U3496));
  NOR2X1  g06310(.A(n7975), .B(n7976), .Y(n7983));
  OAI21X1 g06311(.A0(n6328), .A1(n6327), .B0(n6750), .Y(n7984));
  XOR2X1  g06312(.A(n7984), .B(n7983), .Y(n7985));
  AOI22X1 g06313(.A0(n6556), .A1(P2_REG2_REG_31__SCAN_IN), .B0(P2_REG0_REG_31__SCAN_IN), .B1(n6557), .Y(n7986));
  INVX1   g06314(.A(n7986), .Y(n7987));
  AOI21X1 g06315(.A0(n6559), .A1(P2_REG1_REG_31__SCAN_IN), .B0(n7987), .Y(n7988));
  NOR2X1  g06316(.A(n7988), .B(n7951), .Y(n7989));
  INVX1   g06317(.A(n7989), .Y(n7990));
  OAI21X1 g06318(.A0(n7984), .A1(n6528), .B0(n7990), .Y(n7991));
  AOI21X1 g06319(.A0(n7985), .A1(n6532), .B0(n7991), .Y(n7992));
  NAND2X1 g06320(.A(n6465), .B(P2_REG0_REG_30__SCAN_IN), .Y(n7993));
  OAI21X1 g06321(.A0(n7992), .A1(n6465), .B0(n7993), .Y(P2_U3497));
  NAND4X1 g06322(.A(n7941), .B(n7924), .C(n7921), .D(n7984), .Y(n7995));
  NAND4X1 g06323(.A(n4480), .B(n4478), .C(n1837), .D(n2526), .Y(n7996));
  INVX1   g06324(.A(n6335), .Y(n7997));
  AOI21X1 g06325(.A0(n7997), .A1(n7996), .B0(n6474), .Y(n7998));
  XOR2X1  g06326(.A(n7998), .B(n7995), .Y(n7999));
  NAND2X1 g06327(.A(n7998), .B(n6529), .Y(n8000));
  NAND2X1 g06328(.A(n8000), .B(n7990), .Y(n8001));
  AOI21X1 g06329(.A0(n7999), .A1(n6532), .B0(n8001), .Y(n8002));
  NAND2X1 g06330(.A(n6465), .B(P2_REG0_REG_31__SCAN_IN), .Y(n8003));
  OAI21X1 g06331(.A0(n8002), .A1(n6465), .B0(n8003), .Y(P2_U3498));
  INVX1   g06332(.A(n6464), .Y(n8005));
  NAND4X1 g06333(.A(n6462), .B(n6444), .C(n6350), .D(n8005), .Y(n8006));
  NAND2X1 g06334(.A(n8006), .B(P2_REG1_REG_0__SCAN_IN), .Y(n8007));
  OAI21X1 g06335(.A0(n8006), .A1(n6546), .B0(n8007), .Y(P2_U3499));
  NAND2X1 g06336(.A(n8006), .B(P2_REG1_REG_1__SCAN_IN), .Y(n8009));
  OAI21X1 g06337(.A0(n8006), .A1(n6586), .B0(n8009), .Y(P2_U3500));
  NAND2X1 g06338(.A(n8006), .B(P2_REG1_REG_2__SCAN_IN), .Y(n8011));
  OAI21X1 g06339(.A0(n8006), .A1(n6630), .B0(n8011), .Y(P2_U3501));
  NAND2X1 g06340(.A(n8006), .B(P2_REG1_REG_3__SCAN_IN), .Y(n8013));
  OAI21X1 g06341(.A0(n8006), .A1(n6689), .B0(n8013), .Y(P2_U3502));
  NAND2X1 g06342(.A(n8006), .B(P2_REG1_REG_4__SCAN_IN), .Y(n8015));
  OAI21X1 g06343(.A0(n8006), .A1(n6736), .B0(n8015), .Y(P2_U3503));
  NAND2X1 g06344(.A(n8006), .B(P2_REG1_REG_5__SCAN_IN), .Y(n8017));
  OAI21X1 g06345(.A0(n8006), .A1(n6790), .B0(n8017), .Y(P2_U3504));
  NAND2X1 g06346(.A(n8006), .B(P2_REG1_REG_6__SCAN_IN), .Y(n8019));
  OAI21X1 g06347(.A0(n8006), .A1(n6844), .B0(n8019), .Y(P2_U3505));
  NAND2X1 g06348(.A(n8006), .B(P2_REG1_REG_7__SCAN_IN), .Y(n8021));
  OAI21X1 g06349(.A0(n8006), .A1(n6899), .B0(n8021), .Y(P2_U3506));
  NAND2X1 g06350(.A(n8006), .B(P2_REG1_REG_8__SCAN_IN), .Y(n8023));
  OAI21X1 g06351(.A0(n8006), .A1(n6949), .B0(n8023), .Y(P2_U3507));
  NAND2X1 g06352(.A(n8006), .B(P2_REG1_REG_9__SCAN_IN), .Y(n8025));
  OAI21X1 g06353(.A0(n8006), .A1(n6997), .B0(n8025), .Y(P2_U3508));
  NAND2X1 g06354(.A(n8006), .B(P2_REG1_REG_10__SCAN_IN), .Y(n8027));
  OAI21X1 g06355(.A0(n8006), .A1(n7055), .B0(n8027), .Y(P2_U3509));
  NAND2X1 g06356(.A(n8006), .B(P2_REG1_REG_11__SCAN_IN), .Y(n8029));
  OAI21X1 g06357(.A0(n8006), .A1(n7108), .B0(n8029), .Y(P2_U3510));
  NAND2X1 g06358(.A(n8006), .B(P2_REG1_REG_12__SCAN_IN), .Y(n8031));
  OAI21X1 g06359(.A0(n8006), .A1(n7157), .B0(n8031), .Y(P2_U3511));
  NAND2X1 g06360(.A(n8006), .B(P2_REG1_REG_13__SCAN_IN), .Y(n8033));
  OAI21X1 g06361(.A0(n8006), .A1(n7211), .B0(n8033), .Y(P2_U3512));
  NAND2X1 g06362(.A(n8006), .B(P2_REG1_REG_14__SCAN_IN), .Y(n8035));
  OAI21X1 g06363(.A0(n8006), .A1(n7258), .B0(n8035), .Y(P2_U3513));
  NAND2X1 g06364(.A(n8006), .B(P2_REG1_REG_15__SCAN_IN), .Y(n8037));
  OAI21X1 g06365(.A0(n8006), .A1(n7309), .B0(n8037), .Y(P2_U3514));
  NAND2X1 g06366(.A(n8006), .B(P2_REG1_REG_16__SCAN_IN), .Y(n8039));
  OAI21X1 g06367(.A0(n8006), .A1(n7364), .B0(n8039), .Y(P2_U3515));
  NAND2X1 g06368(.A(n8006), .B(P2_REG1_REG_17__SCAN_IN), .Y(n8041));
  OAI21X1 g06369(.A0(n8006), .A1(n7418), .B0(n8041), .Y(P2_U3516));
  NAND2X1 g06370(.A(n8006), .B(P2_REG1_REG_18__SCAN_IN), .Y(n8043));
  OAI21X1 g06371(.A0(n8006), .A1(n7466), .B0(n8043), .Y(P2_U3517));
  NAND2X1 g06372(.A(n8006), .B(P2_REG1_REG_19__SCAN_IN), .Y(n8045));
  OAI21X1 g06373(.A0(n8006), .A1(n7514), .B0(n8045), .Y(P2_U3518));
  NAND2X1 g06374(.A(n8006), .B(P2_REG1_REG_20__SCAN_IN), .Y(n8047));
  OAI21X1 g06375(.A0(n8006), .A1(n7562), .B0(n8047), .Y(P2_U3519));
  NAND2X1 g06376(.A(n8006), .B(P2_REG1_REG_21__SCAN_IN), .Y(n8049));
  OAI21X1 g06377(.A0(n8006), .A1(n7605), .B0(n8049), .Y(P2_U3520));
  NAND2X1 g06378(.A(n8006), .B(P2_REG1_REG_22__SCAN_IN), .Y(n8051));
  OAI21X1 g06379(.A0(n8006), .A1(n7647), .B0(n8051), .Y(P2_U3521));
  NAND2X1 g06380(.A(n8006), .B(P2_REG1_REG_23__SCAN_IN), .Y(n8053));
  OAI21X1 g06381(.A0(n8006), .A1(n7691), .B0(n8053), .Y(P2_U3522));
  NAND2X1 g06382(.A(n8006), .B(P2_REG1_REG_24__SCAN_IN), .Y(n8055));
  OAI21X1 g06383(.A0(n8006), .A1(n7739), .B0(n8055), .Y(P2_U3523));
  NAND2X1 g06384(.A(n8006), .B(P2_REG1_REG_25__SCAN_IN), .Y(n8057));
  OAI21X1 g06385(.A0(n8006), .A1(n7784), .B0(n8057), .Y(P2_U3524));
  NAND2X1 g06386(.A(n8006), .B(P2_REG1_REG_26__SCAN_IN), .Y(n8059));
  OAI21X1 g06387(.A0(n8006), .A1(n7829), .B0(n8059), .Y(P2_U3525));
  NAND2X1 g06388(.A(n8006), .B(P2_REG1_REG_27__SCAN_IN), .Y(n8061));
  OAI21X1 g06389(.A0(n8006), .A1(n7890), .B0(n8061), .Y(P2_U3526));
  NAND2X1 g06390(.A(n8006), .B(P2_REG1_REG_28__SCAN_IN), .Y(n8063));
  OAI21X1 g06391(.A0(n8006), .A1(n7936), .B0(n8063), .Y(P2_U3527));
  NAND2X1 g06392(.A(n8006), .B(P2_REG1_REG_29__SCAN_IN), .Y(n8065));
  OAI21X1 g06393(.A0(n8006), .A1(n7980), .B0(n8065), .Y(P2_U3528));
  NAND2X1 g06394(.A(n8006), .B(P2_REG1_REG_30__SCAN_IN), .Y(n8067));
  OAI21X1 g06395(.A0(n8006), .A1(n7992), .B0(n8067), .Y(P2_U3529));
  NAND2X1 g06396(.A(n8006), .B(P2_REG1_REG_31__SCAN_IN), .Y(n8069));
  OAI21X1 g06397(.A0(n8006), .A1(n8002), .B0(n8069), .Y(P2_U3530));
  NOR4X1  g06398(.A(n6456), .B(n6452), .C(n6458), .D(n6460), .Y(n8071));
  INVX1   g06399(.A(n6444), .Y(n8072));
  INVX1   g06400(.A(n7949), .Y(n8073));
  AOI21X1 g06401(.A0(n6460), .A1(n6451), .B0(n8073), .Y(n8074));
  NOR4X1  g06402(.A(n8005), .B(n6446), .C(n8072), .D(n8074), .Y(n8075));
  OAI21X1 g06403(.A0(n8075), .A1(n8071), .B0(n6350), .Y(n8076));
  NOR2X1  g06404(.A(n8076), .B(n6535), .Y(n8077));
  NAND2X1 g06405(.A(n8077), .B(n6569), .Y(n8078));
  INVX1   g06406(.A(n8076), .Y(n8079));
  NOR2X1  g06407(.A(n8079), .B(n6484), .Y(n8080));
  AOI21X1 g06408(.A0(n8079), .A1(n6523), .B0(n8080), .Y(n8081));
  NAND3X1 g06409(.A(n6455), .B(n6452), .C(n6449), .Y(n8082));
  NOR2X1  g06410(.A(n8082), .B(n8076), .Y(n8083));
  INVX1   g06411(.A(n8071), .Y(n8084));
  NOR4X1  g06412(.A(n6349), .B(n6342), .C(P2_U3088), .D(n8084), .Y(n8085));
  AOI22X1 g06413(.A0(n8083), .A1(n6483), .B0(P2_REG3_REG_0__SCAN_IN), .B1(n8085), .Y(n8086));
  NOR4X1  g06414(.A(n6456), .B(n6452), .C(n6458), .D(n6513), .Y(n8087));
  NOR2X1  g06415(.A(n9432), .B(n8076), .Y(n8089));
  NOR4X1  g06416(.A(n6460), .B(n6455), .C(n6452), .D(n8076), .Y(n8090));
  AOI22X1 g06417(.A0(n8089), .A1(n6483), .B0(n9403), .B1(n8090), .Y(n8091));
  NAND4X1 g06418(.A(n8086), .B(n8081), .C(n8078), .D(n8091), .Y(P2_U3265));
  NAND2X1 g06419(.A(n8077), .B(n6583), .Y(n8093));
  NOR2X1  g06420(.A(n8079), .B(n6536), .Y(n8094));
  AOI21X1 g06421(.A0(n8079), .A1(n6577), .B0(n8094), .Y(n8095));
  AOI22X1 g06422(.A0(n8083), .A1(n6580), .B0(P2_REG3_REG_1__SCAN_IN), .B1(n8085), .Y(n8096));
  NOR3X1  g06423(.A(n9432), .B(n8076), .C(n6579), .Y(n8097));
  AOI21X1 g06424(.A0(n8090), .A1(n6564), .B0(n8097), .Y(n8098));
  NAND4X1 g06425(.A(n8096), .B(n8095), .C(n8093), .D(n8098), .Y(P2_U3264));
  NAND2X1 g06426(.A(n8077), .B(n6652), .Y(n8100));
  NOR2X1  g06427(.A(n8079), .B(n6589), .Y(n8101));
  AOI21X1 g06428(.A0(n8079), .A1(n6617), .B0(n8101), .Y(n8102));
  AOI22X1 g06429(.A0(n8083), .A1(n6600), .B0(P2_REG3_REG_2__SCAN_IN), .B1(n8085), .Y(n8103));
  AOI22X1 g06430(.A0(n8089), .A1(n6620), .B0(n6608), .B1(n8090), .Y(n8104));
  NAND4X1 g06431(.A(n8103), .B(n8102), .C(n8100), .D(n8104), .Y(P2_U3263));
  NAND2X1 g06432(.A(n8077), .B(n6706), .Y(n8106));
  AOI21X1 g06433(.A0(n6672), .A1(n6660), .B0(n8076), .Y(n8107));
  AOI21X1 g06434(.A0(n8076), .A1(P2_REG2_REG_3__SCAN_IN), .B0(n8107), .Y(n8108));
  AOI22X1 g06435(.A0(n8083), .A1(n6646), .B0(n6650), .B1(n8085), .Y(n8109));
  INVX1   g06436(.A(n6655), .Y(n8110));
  AOI22X1 g06437(.A0(n8089), .A1(n6675), .B0(n8110), .B1(n8090), .Y(n8111));
  NAND4X1 g06438(.A(n8109), .B(n8108), .C(n8106), .D(n8111), .Y(P2_U3262));
  NAND2X1 g06439(.A(n8077), .B(n6745), .Y(n8113));
  AOI22X1 g06440(.A0(n8083), .A1(n6703), .B0(n6724), .B1(n8089), .Y(n8114));
  NOR2X1  g06441(.A(n8079), .B(n6678), .Y(n8115));
  AOI21X1 g06442(.A0(n8079), .A1(n6721), .B0(n8115), .Y(n8116));
  INVX1   g06443(.A(n6683), .Y(n8117));
  AOI22X1 g06444(.A0(n8085), .A1(n8117), .B0(n6710), .B1(n8090), .Y(n8118));
  NAND4X1 g06445(.A(n8116), .B(n8114), .C(n8113), .D(n8118), .Y(P2_U3261));
  NAND2X1 g06446(.A(n8079), .B(n6773), .Y(n8120));
  AOI22X1 g06447(.A0(n8076), .A1(P2_REG2_REG_5__SCAN_IN), .B0(n6807), .B1(n8077), .Y(n8121));
  AOI22X1 g06448(.A0(n8085), .A1(n6743), .B0(n6761), .B1(n8090), .Y(n8122));
  AOI22X1 g06449(.A0(n8083), .A1(n6752), .B0(n6776), .B1(n8089), .Y(n8123));
  NAND4X1 g06450(.A(n8122), .B(n8121), .C(n8120), .D(n8123), .Y(P2_U3260));
  NAND2X1 g06451(.A(n8079), .B(n6823), .Y(n8125));
  AOI22X1 g06452(.A0(n8076), .A1(P2_REG2_REG_6__SCAN_IN), .B0(n6839), .B1(n8077), .Y(n8126));
  INVX1   g06453(.A(n6784), .Y(n8127));
  INVX1   g06454(.A(n8090), .Y(n8128));
  NOR2X1  g06455(.A(n8128), .B(n6810), .Y(n8129));
  AOI21X1 g06456(.A0(n8085), .A1(n8127), .B0(n8129), .Y(n8130));
  AOI22X1 g06457(.A0(n8083), .A1(n6797), .B0(n6833), .B1(n8089), .Y(n8131));
  NAND4X1 g06458(.A(n8130), .B(n8126), .C(n8125), .D(n8131), .Y(P2_U3259));
  INVX1   g06459(.A(P2_REG2_REG_7__SCAN_IN), .Y(n8133));
  INVX1   g06460(.A(n8077), .Y(n8134));
  OAI22X1 g06461(.A0(n8079), .A1(n8133), .B0(n6895), .B1(n8134), .Y(n8135));
  INVX1   g06462(.A(n8085), .Y(n8136));
  OAI22X1 g06463(.A0(n8136), .A1(n6836), .B0(n6864), .B1(n8128), .Y(n8137));
  INVX1   g06464(.A(n8083), .Y(n8138));
  NAND2X1 g06465(.A(n8089), .B(n6885), .Y(n8139));
  OAI21X1 g06466(.A0(n8138), .A1(n6886), .B0(n8139), .Y(n8140));
  NOR3X1  g06467(.A(n8140), .B(n8137), .C(n8135), .Y(n8141));
  OAI21X1 g06468(.A0(n8076), .A1(n6878), .B0(n8141), .Y(P2_U3258));
  NAND2X1 g06469(.A(n8079), .B(n6930), .Y(n8143));
  AOI22X1 g06470(.A0(n8076), .A1(P2_REG2_REG_8__SCAN_IN), .B0(n6944), .B1(n8077), .Y(n8144));
  NOR2X1  g06471(.A(n8128), .B(n6913), .Y(n8145));
  AOI21X1 g06472(.A0(n8085), .A1(n6892), .B0(n8145), .Y(n8146));
  AOI22X1 g06473(.A0(n8083), .A1(n6909), .B0(n6936), .B1(n8089), .Y(n8147));
  NAND4X1 g06474(.A(n8146), .B(n8144), .C(n8143), .D(n8147), .Y(P2_U3257));
  NOR2X1  g06475(.A(n8128), .B(n6974), .Y(n8149));
  AOI22X1 g06476(.A0(n8076), .A1(P2_REG2_REG_9__SCAN_IN), .B0(n6992), .B1(n8077), .Y(n8150));
  NAND2X1 g06477(.A(n8083), .B(n6956), .Y(n8151));
  AOI22X1 g06478(.A0(n8085), .A1(n6942), .B0(n6985), .B1(n8089), .Y(n8152));
  NAND3X1 g06479(.A(n8152), .B(n8151), .C(n8150), .Y(n8153));
  NOR2X1  g06480(.A(n8153), .B(n8149), .Y(n8154));
  OAI21X1 g06481(.A0(n8076), .A1(n6978), .B0(n8154), .Y(P2_U3256));
  NOR2X1  g06482(.A(n8128), .B(n7019), .Y(n8156));
  AOI22X1 g06483(.A0(n8076), .A1(P2_REG2_REG_10__SCAN_IN), .B0(n7072), .B1(n8077), .Y(n8157));
  NAND2X1 g06484(.A(n8083), .B(n7004), .Y(n8158));
  AOI22X1 g06485(.A0(n8085), .A1(n6990), .B0(n7042), .B1(n8089), .Y(n8159));
  NAND3X1 g06486(.A(n8159), .B(n8158), .C(n8157), .Y(n8160));
  NOR2X1  g06487(.A(n8160), .B(n8156), .Y(n8161));
  OAI21X1 g06488(.A0(n8076), .A1(n7034), .B0(n8161), .Y(P2_U3255));
  NOR3X1  g06489(.A(n7092), .B(n7091), .C(n7090), .Y(n8163));
  NOR2X1  g06490(.A(n8128), .B(n7086), .Y(n8164));
  AOI22X1 g06491(.A0(n8076), .A1(P2_REG2_REG_11__SCAN_IN), .B0(n7103), .B1(n8077), .Y(n8165));
  NAND2X1 g06492(.A(n8083), .B(n7063), .Y(n8166));
  AOI22X1 g06493(.A0(n8085), .A1(n7048), .B0(n7097), .B1(n8089), .Y(n8167));
  NAND3X1 g06494(.A(n8167), .B(n8166), .C(n8165), .Y(n8168));
  NOR2X1  g06495(.A(n8168), .B(n8164), .Y(n8169));
  OAI21X1 g06496(.A0(n8076), .A1(n8163), .B0(n8169), .Y(P2_U3254));
  NOR2X1  g06497(.A(n8128), .B(n7134), .Y(n8171));
  INVX1   g06498(.A(P2_REG2_REG_12__SCAN_IN), .Y(n8172));
  OAI22X1 g06499(.A0(n8079), .A1(n8172), .B0(n7165), .B1(n8134), .Y(n8173));
  NOR3X1  g06500(.A(n8082), .B(n8076), .C(n7147), .Y(n8174));
  INVX1   g06501(.A(n7101), .Y(n8175));
  INVX1   g06502(.A(n8089), .Y(n8176));
  OAI22X1 g06503(.A0(n8136), .A1(n8175), .B0(n7148), .B1(n8176), .Y(n8177));
  NOR4X1  g06504(.A(n8174), .B(n8173), .C(n8171), .D(n8177), .Y(n8178));
  OAI21X1 g06505(.A0(n8076), .A1(n7138), .B0(n8178), .Y(P2_U3253));
  NAND2X1 g06506(.A(n8079), .B(n7194), .Y(n8180));
  NOR2X1  g06507(.A(n8128), .B(n7181), .Y(n8181));
  NAND2X1 g06508(.A(n8089), .B(n7200), .Y(n8182));
  AOI22X1 g06509(.A0(n8076), .A1(P2_REG2_REG_13__SCAN_IN), .B0(n7206), .B1(n8077), .Y(n8183));
  AOI22X1 g06510(.A0(n8083), .A1(n7164), .B0(n7152), .B1(n8085), .Y(n8184));
  NAND3X1 g06511(.A(n8184), .B(n8183), .C(n8182), .Y(n8185));
  NOR2X1  g06512(.A(n8185), .B(n8181), .Y(n8186));
  NAND2X1 g06513(.A(n8186), .B(n8180), .Y(P2_U3252));
  NOR2X1  g06514(.A(n8128), .B(n7231), .Y(n8188));
  NOR3X1  g06515(.A(n9432), .B(n8076), .C(n7248), .Y(n8189));
  INVX1   g06516(.A(P2_REG2_REG_14__SCAN_IN), .Y(n8190));
  OAI22X1 g06517(.A0(n8079), .A1(n8190), .B0(n7312), .B1(n8134), .Y(n8191));
  OAI22X1 g06518(.A0(n8138), .A1(n7218), .B0(n7203), .B1(n8136), .Y(n8192));
  NOR4X1  g06519(.A(n8191), .B(n8189), .C(n8188), .D(n8192), .Y(n8193));
  OAI21X1 g06520(.A0(n8076), .A1(n7238), .B0(n8193), .Y(P2_U3251));
  NOR2X1  g06521(.A(n8128), .B(n7283), .Y(n8195));
  NAND2X1 g06522(.A(n8089), .B(n7296), .Y(n8196));
  AOI22X1 g06523(.A0(n8076), .A1(P2_REG2_REG_15__SCAN_IN), .B0(n7304), .B1(n8077), .Y(n8197));
  AOI22X1 g06524(.A0(n8083), .A1(n7313), .B0(n7253), .B1(n8085), .Y(n8198));
  NAND3X1 g06525(.A(n8198), .B(n8197), .C(n8196), .Y(n8199));
  NOR2X1  g06526(.A(n8199), .B(n8195), .Y(n8200));
  OAI21X1 g06527(.A0(n8076), .A1(n7290), .B0(n8200), .Y(P2_U3250));
  NAND2X1 g06528(.A(n8079), .B(n7346), .Y(n8202));
  NOR2X1  g06529(.A(n8128), .B(n7350), .Y(n8203));
  NAND2X1 g06530(.A(n8089), .B(n7352), .Y(n8204));
  AOI22X1 g06531(.A0(n8076), .A1(P2_REG2_REG_16__SCAN_IN), .B0(n7326), .B1(n8083), .Y(n8205));
  AOI22X1 g06532(.A0(n8077), .A1(n7368), .B0(n7302), .B1(n8085), .Y(n8206));
  NAND3X1 g06533(.A(n8206), .B(n8205), .C(n8204), .Y(n8207));
  NOR2X1  g06534(.A(n8207), .B(n8203), .Y(n8208));
  NAND2X1 g06535(.A(n8208), .B(n8202), .Y(P2_U3249));
  NAND2X1 g06536(.A(n8079), .B(n7400), .Y(n8210));
  NOR2X1  g06537(.A(n8128), .B(n7384), .Y(n8211));
  NAND2X1 g06538(.A(n8089), .B(n7406), .Y(n8212));
  AOI22X1 g06539(.A0(n8076), .A1(P2_REG2_REG_17__SCAN_IN), .B0(n7373), .B1(n8083), .Y(n8213));
  AOI22X1 g06540(.A0(n8077), .A1(n7432), .B0(n7356), .B1(n8085), .Y(n8214));
  NAND3X1 g06541(.A(n8214), .B(n8213), .C(n8212), .Y(n8215));
  NOR2X1  g06542(.A(n8215), .B(n8211), .Y(n8216));
  NAND2X1 g06543(.A(n8216), .B(n8210), .Y(P2_U3248));
  NAND2X1 g06544(.A(n8079), .B(n7446), .Y(n8218));
  NOR2X1  g06545(.A(n8128), .B(n7435), .Y(n8219));
  NOR4X1  g06546(.A(n8076), .B(n7456), .C(n7455), .D(n9432), .Y(n8220));
  AOI22X1 g06547(.A0(n8076), .A1(P2_REG2_REG_18__SCAN_IN), .B0(n7425), .B1(n8083), .Y(n8221));
  AOI22X1 g06548(.A0(n8077), .A1(n7486), .B0(n7410), .B1(n8085), .Y(n8222));
  NAND2X1 g06549(.A(n8222), .B(n8221), .Y(n8223));
  NOR3X1  g06550(.A(n8223), .B(n8220), .C(n8219), .Y(n8224));
  NAND2X1 g06551(.A(n8224), .B(n8218), .Y(P2_U3247));
  NAND2X1 g06552(.A(n8079), .B(n7495), .Y(n8226));
  OAI21X1 g06553(.A0(n7500), .A1(n7485), .B0(n8090), .Y(n8228));
  NAND2X1 g06554(.A(n8089), .B(n7503), .Y(n8229));
  AOI22X1 g06555(.A0(n8076), .A1(P2_REG2_REG_19__SCAN_IN), .B0(n7460), .B1(n8085), .Y(n8230));
  OAI21X1 g06556(.A0(n8134), .A1(n7510), .B0(n8230), .Y(n8231));
  AOI21X1 g06557(.A0(n8083), .A1(n7470), .B0(n8231), .Y(n8232));
  NAND4X1 g06558(.A(n8229), .B(n8228), .C(n8226), .D(n8232), .Y(P2_U3246));
  NAND2X1 g06559(.A(n8079), .B(n7545), .Y(n8234));
  NAND2X1 g06560(.A(n8090), .B(n7540), .Y(n8236));
  NAND2X1 g06561(.A(n8089), .B(n7551), .Y(n8237));
  INVX1   g06562(.A(n7505), .Y(n8238));
  AOI22X1 g06563(.A0(n8076), .A1(P2_REG2_REG_20__SCAN_IN), .B0(n8238), .B1(n8085), .Y(n8239));
  OAI21X1 g06564(.A0(n8134), .A1(n7558), .B0(n8239), .Y(n8240));
  AOI21X1 g06565(.A0(n8083), .A1(n7527), .B0(n8240), .Y(n8241));
  NAND4X1 g06566(.A(n8237), .B(n8236), .C(n8234), .D(n8241), .Y(P2_U3245));
  NOR3X1  g06567(.A(n7586), .B(n7585), .C(n7584), .Y(n8243));
  NOR2X1  g06568(.A(n8128), .B(n7589), .Y(n8244));
  NAND2X1 g06569(.A(n8089), .B(n7591), .Y(n8245));
  NAND2X1 g06570(.A(n8083), .B(n7565), .Y(n8246));
  NAND2X1 g06571(.A(n8077), .B(n7600), .Y(n8247));
  INVX1   g06572(.A(n7553), .Y(n8248));
  AOI22X1 g06573(.A0(n8076), .A1(P2_REG2_REG_21__SCAN_IN), .B0(n8248), .B1(n8085), .Y(n8249));
  NAND4X1 g06574(.A(n8247), .B(n8246), .C(n8245), .D(n8249), .Y(n8250));
  NOR2X1  g06575(.A(n8250), .B(n8244), .Y(n8251));
  OAI21X1 g06576(.A0(n8076), .A1(n8243), .B0(n8251), .Y(P2_U3244));
  NOR3X1  g06577(.A(n7629), .B(n7628), .C(n7627), .Y(n8253));
  NOR2X1  g06578(.A(n8128), .B(n7623), .Y(n8254));
  NAND2X1 g06579(.A(n8089), .B(n7634), .Y(n8255));
  NAND2X1 g06580(.A(n8083), .B(n7608), .Y(n8256));
  NAND2X1 g06581(.A(n8077), .B(n7642), .Y(n8257));
  INVX1   g06582(.A(n7596), .Y(n8258));
  AOI22X1 g06583(.A0(n8076), .A1(P2_REG2_REG_22__SCAN_IN), .B0(n8258), .B1(n8085), .Y(n8259));
  NAND4X1 g06584(.A(n8257), .B(n8256), .C(n8255), .D(n8259), .Y(n8260));
  NOR2X1  g06585(.A(n8260), .B(n8254), .Y(n8261));
  OAI21X1 g06586(.A0(n8076), .A1(n8253), .B0(n8261), .Y(P2_U3243));
  NOR2X1  g06587(.A(n8128), .B(n7666), .Y(n8263));
  INVX1   g06588(.A(n7638), .Y(n8264));
  AOI22X1 g06589(.A0(n8076), .A1(P2_REG2_REG_23__SCAN_IN), .B0(n8264), .B1(n8085), .Y(n8265));
  OAI21X1 g06590(.A0(n8134), .A1(n7694), .B0(n8265), .Y(n8266));
  AOI21X1 g06591(.A0(n8083), .A1(n7652), .B0(n8266), .Y(n8267));
  OAI21X1 g06592(.A0(n8176), .A1(n7681), .B0(n8267), .Y(n8268));
  NOR2X1  g06593(.A(n8268), .B(n8263), .Y(n8269));
  OAI21X1 g06594(.A0(n8076), .A1(n7673), .B0(n8269), .Y(P2_U3242));
  NOR3X1  g06595(.A(n7720), .B(n7719), .C(n7718), .Y(n8271));
  NOR2X1  g06596(.A(n8128), .B(n7726), .Y(n8272));
  NOR2X1  g06597(.A(n7723), .B(n7727), .Y(n8273));
  NOR3X1  g06598(.A(n8176), .B(n7772), .C(n8273), .Y(n8274));
  NOR4X1  g06599(.A(n8076), .B(n6474), .C(n6261), .D(n8082), .Y(n8275));
  AOI22X1 g06600(.A0(n8076), .A1(P2_REG2_REG_24__SCAN_IN), .B0(n7683), .B1(n8085), .Y(n8276));
  OAI21X1 g06601(.A0(n8134), .A1(n7735), .B0(n8276), .Y(n8277));
  NOR4X1  g06602(.A(n8275), .B(n8274), .C(n8272), .D(n8277), .Y(n8278));
  OAI21X1 g06603(.A0(n8076), .A1(n8271), .B0(n8278), .Y(P2_U3241));
  OAI21X1 g06604(.A0(n7766), .A1(n7763), .B0(n8079), .Y(n8280));
  NOR2X1  g06605(.A(n8128), .B(n7771), .Y(n8281));
  INVX1   g06606(.A(n7773), .Y(n8282));
  NOR2X1  g06607(.A(n8176), .B(n8282), .Y(n8283));
  NOR3X1  g06608(.A(n8138), .B(n6474), .C(n6268), .Y(n8284));
  INVX1   g06609(.A(n7730), .Y(n8285));
  AOI22X1 g06610(.A0(n8076), .A1(P2_REG2_REG_25__SCAN_IN), .B0(n8285), .B1(n8085), .Y(n8286));
  OAI21X1 g06611(.A0(n8134), .A1(n7780), .B0(n8286), .Y(n8287));
  NOR4X1  g06612(.A(n8284), .B(n8283), .C(n8281), .D(n8287), .Y(n8288));
  NAND2X1 g06613(.A(n8288), .B(n8280), .Y(P2_U3240));
  OAI21X1 g06614(.A0(n7811), .A1(n7809), .B0(n8079), .Y(n8290));
  NAND3X1 g06615(.A(n8090), .B(n7804), .C(n7812), .Y(n8291));
  NAND2X1 g06616(.A(n8089), .B(n7818), .Y(n8292));
  INVX1   g06617(.A(n7775), .Y(n8293));
  AOI22X1 g06618(.A0(n8076), .A1(P2_REG2_REG_26__SCAN_IN), .B0(n8293), .B1(n8085), .Y(n8294));
  OAI21X1 g06619(.A0(n8134), .A1(n7825), .B0(n8294), .Y(n8295));
  AOI21X1 g06620(.A0(n8083), .A1(n7817), .B0(n8295), .Y(n8296));
  NAND4X1 g06621(.A(n8292), .B(n8291), .C(n8290), .D(n8296), .Y(P2_U3239));
  OAI21X1 g06622(.A0(n7868), .A1(n7865), .B0(n8079), .Y(n8298));
  NAND2X1 g06623(.A(n8090), .B(n7860), .Y(n8300));
  NAND2X1 g06624(.A(n8089), .B(n7877), .Y(n8301));
  INVX1   g06625(.A(n7820), .Y(n8302));
  AOI22X1 g06626(.A0(n8076), .A1(P2_REG2_REG_27__SCAN_IN), .B0(n8302), .B1(n8085), .Y(n8303));
  OAI21X1 g06627(.A0(n8134), .A1(n7886), .B0(n8303), .Y(n8304));
  AOI21X1 g06628(.A0(n8083), .A1(n7876), .B0(n8304), .Y(n8305));
  NAND4X1 g06629(.A(n8301), .B(n8300), .C(n8298), .D(n8305), .Y(P2_U3238));
  NOR3X1  g06630(.A(n7915), .B(n7914), .C(n7913), .Y(n8307));
  NAND2X1 g06631(.A(n8089), .B(n7925), .Y(n8308));
  INVX1   g06632(.A(n7881), .Y(n8309));
  AOI22X1 g06633(.A0(n8076), .A1(P2_REG2_REG_28__SCAN_IN), .B0(n8309), .B1(n8085), .Y(n8310));
  OAI21X1 g06634(.A0(n8134), .A1(n7932), .B0(n8310), .Y(n8311));
  AOI21X1 g06635(.A0(n8083), .A1(n7893), .B0(n8311), .Y(n8312));
  NAND2X1 g06636(.A(n8312), .B(n8308), .Y(n8313));
  AOI21X1 g06637(.A0(n8090), .A1(n7919), .B0(n8313), .Y(n8314));
  OAI21X1 g06638(.A0(n8076), .A1(n8307), .B0(n8314), .Y(P2_U3237));
  NOR3X1  g06639(.A(n7970), .B(n7969), .C(n7960), .Y(n8316));
  NOR2X1  g06640(.A(n8128), .B(n7974), .Y(n8317));
  NAND2X1 g06641(.A(n8089), .B(n7977), .Y(n8318));
  NAND3X1 g06642(.A(n8083), .B(n6750), .C(n6314), .Y(n8319));
  AOI22X1 g06643(.A0(n8076), .A1(P2_REG2_REG_29__SCAN_IN), .B0(n7926), .B1(n8085), .Y(n8320));
  NAND3X1 g06644(.A(n8320), .B(n8319), .C(n8318), .Y(n8321));
  NOR2X1  g06645(.A(n8321), .B(n8317), .Y(n8322));
  OAI21X1 g06646(.A0(n8076), .A1(n8316), .B0(n8322), .Y(P2_U3236));
  NAND2X1 g06647(.A(n8089), .B(n7985), .Y(n8324));
  INVX1   g06648(.A(n6328), .Y(n8325));
  OAI21X1 g06649(.A0(n2504), .A1(n1790), .B0(n8325), .Y(n8326));
  NAND3X1 g06650(.A(n8083), .B(n6750), .C(n8326), .Y(n8327));
  NAND2X1 g06651(.A(n8079), .B(n7989), .Y(n8328));
  NAND2X1 g06652(.A(n8076), .B(P2_REG2_REG_30__SCAN_IN), .Y(n8329));
  NAND4X1 g06653(.A(n8328), .B(n8327), .C(n8324), .D(n8329), .Y(P2_U3235));
  NAND2X1 g06654(.A(n8089), .B(n7999), .Y(n8331));
  NAND2X1 g06655(.A(n8083), .B(n7998), .Y(n8332));
  NAND2X1 g06656(.A(n8076), .B(P2_REG2_REG_31__SCAN_IN), .Y(n8333));
  NAND4X1 g06657(.A(n8332), .B(n8331), .C(n8328), .D(n8333), .Y(P2_U3234));
  OAI21X1 g06658(.A0(n8073), .A1(n6342), .B0(n6750), .Y(n8335));
  NOR4X1  g06659(.A(n6349), .B(n6342), .C(P2_U3088), .D(n8335), .Y(n8336));
  INVX1   g06660(.A(P2_REG2_REG_16__SCAN_IN), .Y(n8337));
  INVX1   g06661(.A(P2_REG2_REG_17__SCAN_IN), .Y(n8338));
  AOI22X1 g06662(.A0(n7317), .A1(n8337), .B0(n8338), .B1(n7370), .Y(n8339));
  INVX1   g06663(.A(n8339), .Y(n8340));
  NOR2X1  g06664(.A(n7263), .B(P2_REG2_REG_15__SCAN_IN), .Y(n8341));
  INVX1   g06665(.A(P2_REG2_REG_13__SCAN_IN), .Y(n8342));
  NAND2X1 g06666(.A(n7161), .B(n8342), .Y(n8343));
  INVX1   g06667(.A(P2_REG2_REG_11__SCAN_IN), .Y(n8344));
  NOR2X1  g06668(.A(n7060), .B(n8344), .Y(n8345));
  INVX1   g06669(.A(n8345), .Y(n8346));
  AOI22X1 g06670(.A0(n7112), .A1(n8172), .B0(n8342), .B1(n7161), .Y(n8347));
  INVX1   g06671(.A(n8347), .Y(n8348));
  NOR2X1  g06672(.A(n7112), .B(n8172), .Y(n8349));
  AOI21X1 g06673(.A0(n7162), .A1(P2_REG2_REG_13__SCAN_IN), .B0(n8349), .Y(n8350));
  OAI21X1 g06674(.A0(n8348), .A1(n8346), .B0(n8350), .Y(n8351));
  INVX1   g06675(.A(P2_REG2_REG_10__SCAN_IN), .Y(n8352));
  INVX1   g06676(.A(P2_REG2_REG_8__SCAN_IN), .Y(n8353));
  NOR2X1  g06677(.A(n6906), .B(n8353), .Y(n8354));
  INVX1   g06678(.A(P2_REG2_REG_9__SCAN_IN), .Y(n8355));
  AOI22X1 g06679(.A0(n6953), .A1(n8355), .B0(n8352), .B1(n7001), .Y(n8356));
  OAI22X1 g06680(.A0(n6953), .A1(n8355), .B0(n8352), .B1(n7001), .Y(n8357));
  AOI21X1 g06681(.A0(n8356), .A1(n8354), .B0(n8357), .Y(n8358));
  AOI21X1 g06682(.A0(n7001), .A1(n8352), .B0(n8358), .Y(n8359));
  AOI22X1 g06683(.A0(n6794), .A1(n6777), .B0(n8133), .B1(n6848), .Y(n8360));
  INVX1   g06684(.A(n6701), .Y(n8361));
  AOI22X1 g06685(.A0(n8361), .A1(n6678), .B0(n6725), .B1(n6747), .Y(n8362));
  OAI22X1 g06686(.A0(n6598), .A1(P2_REG2_REG_2__SCAN_IN), .B0(P2_REG2_REG_3__SCAN_IN), .B1(n6644), .Y(n8363));
  NOR2X1  g06687(.A(n6475), .B(n6484), .Y(n8364));
  INVX1   g06688(.A(n8364), .Y(n8365));
  AOI21X1 g06689(.A0(n6551), .A1(n6536), .B0(n8365), .Y(n8366));
  NOR2X1  g06690(.A(n6551), .B(n6536), .Y(n8367));
  NOR2X1  g06691(.A(n8367), .B(n8366), .Y(n8368));
  NOR2X1  g06692(.A(n6643), .B(n6621), .Y(n8369));
  NOR2X1  g06693(.A(n6644), .B(P2_REG2_REG_3__SCAN_IN), .Y(n8370));
  NOR3X1  g06694(.A(n8370), .B(n6597), .C(n6589), .Y(n8371));
  NOR2X1  g06695(.A(n8371), .B(n8369), .Y(n8372));
  OAI21X1 g06696(.A0(n8368), .A1(n8363), .B0(n8372), .Y(n8373));
  NAND2X1 g06697(.A(n8373), .B(n8362), .Y(n8374));
  NOR2X1  g06698(.A(n8361), .B(n6678), .Y(n8375));
  AOI21X1 g06699(.A0(n6701), .A1(P2_REG2_REG_4__SCAN_IN), .B0(P2_REG2_REG_5__SCAN_IN), .Y(n8376));
  NOR2X1  g06700(.A(n8376), .B(n6747), .Y(n8377));
  AOI21X1 g06701(.A0(n8375), .A1(P2_REG2_REG_5__SCAN_IN), .B0(n8377), .Y(n8378));
  NAND2X1 g06702(.A(n8378), .B(n8374), .Y(n8379));
  NAND2X1 g06703(.A(n8379), .B(n8360), .Y(n8380));
  NOR3X1  g06704(.A(n6794), .B(n8133), .C(n6777), .Y(n8381));
  OAI21X1 g06705(.A0(n6794), .A1(n6777), .B0(n8133), .Y(n8382));
  AOI21X1 g06706(.A0(n8382), .A1(n6849), .B0(n8381), .Y(n8383));
  NAND2X1 g06707(.A(n8383), .B(n8380), .Y(n8384));
  NOR2X1  g06708(.A(n6907), .B(P2_REG2_REG_8__SCAN_IN), .Y(n8385));
  INVX1   g06709(.A(n8385), .Y(n8386));
  NAND3X1 g06710(.A(n8386), .B(n8384), .C(n8356), .Y(n8387));
  INVX1   g06711(.A(n8387), .Y(n8388));
  NOR2X1  g06712(.A(n8388), .B(n8359), .Y(n8389));
  INVX1   g06713(.A(n8389), .Y(n8390));
  AOI21X1 g06714(.A0(n7060), .A1(n8344), .B0(n8348), .Y(n8391));
  AOI22X1 g06715(.A0(n8390), .A1(n8391), .B0(n8351), .B1(n8343), .Y(n8392));
  AOI21X1 g06716(.A0(n7215), .A1(n8190), .B0(n8392), .Y(n8393));
  AOI21X1 g06717(.A0(n7216), .A1(P2_REG2_REG_14__SCAN_IN), .B0(n8393), .Y(n8394));
  NOR2X1  g06718(.A(n8394), .B(n8341), .Y(n8395));
  AOI21X1 g06719(.A0(n7263), .A1(P2_REG2_REG_15__SCAN_IN), .B0(n8395), .Y(n8396));
  NOR3X1  g06720(.A(n7317), .B(n8338), .C(n8337), .Y(n8397));
  OAI21X1 g06721(.A0(n7317), .A1(n8337), .B0(n8338), .Y(n8398));
  AOI21X1 g06722(.A0(n8398), .A1(n7371), .B0(n8397), .Y(n8399));
  OAI21X1 g06723(.A0(n8396), .A1(n8340), .B0(n8399), .Y(n8400));
  AOI21X1 g06724(.A0(n7423), .A1(P2_REG2_REG_18__SCAN_IN), .B0(n8400), .Y(n8401));
  XOR2X1  g06725(.A(n6460), .B(P2_REG2_REG_19__SCAN_IN), .Y(n8402));
  INVX1   g06726(.A(n8402), .Y(n8403));
  OAI21X1 g06727(.A0(n7423), .A1(P2_REG2_REG_18__SCAN_IN), .B0(n8403), .Y(n8404));
  OAI21X1 g06728(.A0(n7423), .A1(P2_REG2_REG_18__SCAN_IN), .B0(n8400), .Y(n8405));
  AOI21X1 g06729(.A0(n7423), .A1(P2_REG2_REG_18__SCAN_IN), .B0(n8403), .Y(n8406));
  NAND2X1 g06730(.A(n8406), .B(n8405), .Y(n8407));
  OAI21X1 g06731(.A0(n8404), .A1(n8401), .B0(n8407), .Y(n8408));
  NOR2X1  g06732(.A(n6481), .B(n6480), .Y(n8409));
  NAND3X1 g06733(.A(n6460), .B(n6451), .C(n6458), .Y(n8410));
  OAI21X1 g06734(.A0(n6460), .A1(n6451), .B0(n6456), .Y(n8411));
  INVX1   g06735(.A(n8082), .Y(n8412));
  NAND3X1 g06736(.A(n9432), .B(n6657), .C(n6508), .Y(n8413));
  NOR4X1  g06737(.A(n8412), .B(n8071), .C(n6516), .D(n8413), .Y(n8414));
  NAND4X1 g06738(.A(n8411), .B(n8410), .C(n6669), .D(n8414), .Y(n8415));
  NOR2X1  g06739(.A(n8498), .B(n8408), .Y(n8417));
  INVX1   g06740(.A(P2_REG1_REG_16__SCAN_IN), .Y(n8418));
  AOI22X1 g06741(.A0(n7317), .A1(n8418), .B0(n7357), .B1(n7370), .Y(n8419));
  INVX1   g06742(.A(n8419), .Y(n8420));
  NOR2X1  g06743(.A(n7263), .B(P2_REG1_REG_15__SCAN_IN), .Y(n8421));
  INVX1   g06744(.A(P2_REG1_REG_14__SCAN_IN), .Y(n8422));
  NOR2X1  g06745(.A(n7215), .B(n8422), .Y(n8423));
  NAND2X1 g06746(.A(n7215), .B(n8422), .Y(n8424));
  NAND2X1 g06747(.A(n7061), .B(P2_REG1_REG_11__SCAN_IN), .Y(n8425));
  INVX1   g06748(.A(P2_REG1_REG_12__SCAN_IN), .Y(n8426));
  INVX1   g06749(.A(P2_REG1_REG_13__SCAN_IN), .Y(n8427));
  AOI22X1 g06750(.A0(n7112), .A1(n8426), .B0(n8427), .B1(n7161), .Y(n8428));
  INVX1   g06751(.A(n8428), .Y(n8429));
  NOR2X1  g06752(.A(n7112), .B(n8426), .Y(n8430));
  AOI21X1 g06753(.A0(n7162), .A1(P2_REG1_REG_13__SCAN_IN), .B0(n8430), .Y(n8431));
  OAI21X1 g06754(.A0(n8429), .A1(n8425), .B0(n8431), .Y(n8432));
  OAI21X1 g06755(.A0(n7162), .A1(P2_REG1_REG_13__SCAN_IN), .B0(n8432), .Y(n8433));
  INVX1   g06756(.A(P2_REG1_REG_10__SCAN_IN), .Y(n8434));
  INVX1   g06757(.A(P2_REG1_REG_9__SCAN_IN), .Y(n8435));
  AOI22X1 g06758(.A0(n6953), .A1(n8435), .B0(n8434), .B1(n7001), .Y(n8436));
  NAND3X1 g06759(.A(n8436), .B(n6907), .C(P2_REG1_REG_8__SCAN_IN), .Y(n8437));
  AOI22X1 g06760(.A0(n6954), .A1(P2_REG1_REG_9__SCAN_IN), .B0(P2_REG1_REG_10__SCAN_IN), .B1(n7002), .Y(n8438));
  AOI22X1 g06761(.A0(n8437), .A1(n8438), .B0(n7001), .B1(n8434), .Y(n8439));
  INVX1   g06762(.A(n8439), .Y(n8440));
  INVX1   g06763(.A(P2_REG1_REG_7__SCAN_IN), .Y(n8441));
  AOI22X1 g06764(.A0(n6794), .A1(n6780), .B0(n8441), .B1(n6848), .Y(n8442));
  INVX1   g06765(.A(n8442), .Y(n8443));
  AOI22X1 g06766(.A0(n8361), .A1(n6681), .B0(n6728), .B1(n6747), .Y(n8444));
  OAI22X1 g06767(.A0(n6598), .A1(P2_REG1_REG_2__SCAN_IN), .B0(P2_REG1_REG_3__SCAN_IN), .B1(n6644), .Y(n8445));
  NOR2X1  g06768(.A(n6475), .B(n6495), .Y(n8446));
  INVX1   g06769(.A(n8446), .Y(n8447));
  AOI21X1 g06770(.A0(n6551), .A1(n6539), .B0(n8447), .Y(n8448));
  NOR2X1  g06771(.A(n6551), .B(n6539), .Y(n8449));
  NOR2X1  g06772(.A(n8449), .B(n8448), .Y(n8450));
  NOR2X1  g06773(.A(n6643), .B(n6624), .Y(n8451));
  NOR2X1  g06774(.A(n6644), .B(P2_REG1_REG_3__SCAN_IN), .Y(n8452));
  NOR3X1  g06775(.A(n8452), .B(n6597), .C(n6592), .Y(n8453));
  NOR2X1  g06776(.A(n8453), .B(n8451), .Y(n8454));
  OAI21X1 g06777(.A0(n8450), .A1(n8445), .B0(n8454), .Y(n8455));
  NAND2X1 g06778(.A(n8455), .B(n8444), .Y(n8456));
  NOR2X1  g06779(.A(n8361), .B(n6681), .Y(n8457));
  AOI21X1 g06780(.A0(n6701), .A1(P2_REG1_REG_4__SCAN_IN), .B0(P2_REG1_REG_5__SCAN_IN), .Y(n8458));
  NOR2X1  g06781(.A(n8458), .B(n6747), .Y(n8459));
  AOI21X1 g06782(.A0(n8457), .A1(P2_REG1_REG_5__SCAN_IN), .B0(n8459), .Y(n8460));
  NAND2X1 g06783(.A(n8460), .B(n8456), .Y(n8461));
  INVX1   g06784(.A(n8461), .Y(n8462));
  NOR3X1  g06785(.A(n6794), .B(n8441), .C(n6780), .Y(n8463));
  OAI21X1 g06786(.A0(n6794), .A1(n6780), .B0(n8441), .Y(n8464));
  AOI21X1 g06787(.A0(n8464), .A1(n6849), .B0(n8463), .Y(n8465));
  OAI21X1 g06788(.A0(n8462), .A1(n8443), .B0(n8465), .Y(n8466));
  INVX1   g06789(.A(n8466), .Y(n8467));
  OAI21X1 g06790(.A0(n6907), .A1(P2_REG1_REG_8__SCAN_IN), .B0(n8436), .Y(n8468));
  OAI21X1 g06791(.A0(n8468), .A1(n8467), .B0(n8440), .Y(n8469));
  INVX1   g06792(.A(n8469), .Y(n8470));
  OAI21X1 g06793(.A0(n7061), .A1(P2_REG1_REG_11__SCAN_IN), .B0(n8428), .Y(n8471));
  OAI21X1 g06794(.A0(n8471), .A1(n8470), .B0(n8433), .Y(n8472));
  AOI21X1 g06795(.A0(n8472), .A1(n8424), .B0(n8423), .Y(n8473));
  NOR2X1  g06796(.A(n8473), .B(n8421), .Y(n8474));
  AOI21X1 g06797(.A0(n7263), .A1(P2_REG1_REG_15__SCAN_IN), .B0(n8474), .Y(n8475));
  NOR3X1  g06798(.A(n7317), .B(n7357), .C(n8418), .Y(n8476));
  OAI21X1 g06799(.A0(n7317), .A1(n8418), .B0(n7357), .Y(n8477));
  AOI21X1 g06800(.A0(n8477), .A1(n7371), .B0(n8476), .Y(n8478));
  OAI21X1 g06801(.A0(n8475), .A1(n8420), .B0(n8478), .Y(n8479));
  AOI21X1 g06802(.A0(n7423), .A1(P2_REG1_REG_18__SCAN_IN), .B0(n8479), .Y(n8480));
  XOR2X1  g06803(.A(n6460), .B(P2_REG1_REG_19__SCAN_IN), .Y(n8481));
  INVX1   g06804(.A(n8481), .Y(n8482));
  OAI21X1 g06805(.A0(n7423), .A1(P2_REG1_REG_18__SCAN_IN), .B0(n8482), .Y(n8483));
  OAI21X1 g06806(.A0(n7423), .A1(P2_REG1_REG_18__SCAN_IN), .B0(n8479), .Y(n8484));
  AOI21X1 g06807(.A0(n7423), .A1(P2_REG1_REG_18__SCAN_IN), .B0(n8482), .Y(n8485));
  NAND2X1 g06808(.A(n8485), .B(n8484), .Y(n8486));
  OAI21X1 g06809(.A0(n8483), .A1(n8480), .B0(n8486), .Y(n8487));
  OAI22X1 g06810(.A0(n6469), .A1(n8487), .B0(n6460), .B1(n6473), .Y(n8490));
  OAI21X1 g06811(.A0(n8490), .A1(n8417), .B0(n8336), .Y(n8491));
  NOR4X1  g06812(.A(n6346), .B(n6344), .C(n6342), .D(n6348), .Y(n8492));
  INVX1   g06813(.A(n8492), .Y(n8493));
  NOR2X1  g06814(.A(n8493), .B(P2_U3088), .Y(P2_U3947));
  NOR2X1  g06815(.A(n6481), .B(n6469), .Y(n8495));
  INVX1   g06816(.A(n8495), .Y(n8496));
  NOR2X1  g06817(.A(n8496), .B(n8487), .Y(n8497));
  INVX1   g06818(.A(n8409), .Y(n8498));
  OAI22X1 g06819(.A0(n8408), .A1(n8498), .B0(n6473), .B1(n6460), .Y(n8499));
  OAI21X1 g06820(.A0(n8499), .A1(n8497), .B0(P2_U3947), .Y(n8500));
  NAND3X1 g06821(.A(n8335), .B(n8493), .C(P2_STATE_REG_SCAN_IN), .Y(n8501));
  INVX1   g06822(.A(n8501), .Y(n8502));
  NOR4X1  g06823(.A(n6469), .B(n6341), .C(P2_U3088), .D(n8502), .Y(n8503));
  INVX1   g06824(.A(n8503), .Y(n8504));
  NOR2X1  g06825(.A(n8504), .B(n8487), .Y(n8505));
  NOR4X1  g06826(.A(n8502), .B(n6341), .C(P2_U3088), .D(n8498), .Y(n8506));
  INVX1   g06827(.A(n8506), .Y(n8507));
  NOR2X1  g06828(.A(n8507), .B(n8408), .Y(n8508));
  NOR4X1  g06829(.A(n6473), .B(n6341), .C(P2_U3088), .D(n8502), .Y(n8509));
  INVX1   g06830(.A(n8509), .Y(n8510));
  AOI22X1 g06831(.A0(P2_U3088), .A1(P2_REG3_REG_19__SCAN_IN), .B0(P2_ADDR_REG_19__SCAN_IN), .B1(n8502), .Y(n8511));
  OAI21X1 g06832(.A0(n8510), .A1(n6460), .B0(n8511), .Y(n8512));
  NOR3X1  g06833(.A(n8512), .B(n8508), .C(n8505), .Y(n8513));
  NAND3X1 g06834(.A(n8513), .B(n8500), .C(n8491), .Y(P2_U3233));
  XOR2X1  g06835(.A(n7422), .B(P2_REG2_REG_18__SCAN_IN), .Y(n8515));
  XOR2X1  g06836(.A(n8515), .B(n8400), .Y(n8516));
  NOR2X1  g06837(.A(n8516), .B(n8498), .Y(n8517));
  XOR2X1  g06838(.A(n7422), .B(P2_REG1_REG_18__SCAN_IN), .Y(n8518));
  XOR2X1  g06839(.A(n8518), .B(n8479), .Y(n8519));
  OAI22X1 g06840(.A0(n6473), .A1(n7422), .B0(n6469), .B1(n8519), .Y(n8520));
  OAI21X1 g06841(.A0(n8520), .A1(n8517), .B0(n8336), .Y(n8521));
  NOR2X1  g06842(.A(n8519), .B(n8496), .Y(n8522));
  OAI22X1 g06843(.A0(n8498), .A1(n8516), .B0(n7422), .B1(n6473), .Y(n8523));
  OAI21X1 g06844(.A0(n8523), .A1(n8522), .B0(P2_U3947), .Y(n8524));
  NOR2X1  g06845(.A(n8519), .B(n8504), .Y(n8525));
  OAI22X1 g06846(.A0(P2_STATE_REG_SCAN_IN), .A1(n7407), .B0(n1524), .B1(n8501), .Y(n8526));
  AOI21X1 g06847(.A0(n8509), .A1(n7423), .B0(n8526), .Y(n8527));
  OAI21X1 g06848(.A0(n8516), .A1(n8507), .B0(n8527), .Y(n8528));
  NOR2X1  g06849(.A(n8528), .B(n8525), .Y(n8529));
  NAND3X1 g06850(.A(n8529), .B(n8524), .C(n8521), .Y(P2_U3232));
  OAI21X1 g06851(.A0(n7317), .A1(n8337), .B0(n8396), .Y(n8531));
  AOI21X1 g06852(.A0(n7371), .A1(P2_REG2_REG_17__SCAN_IN), .B0(n8340), .Y(n8532));
  NAND2X1 g06853(.A(n8532), .B(n8531), .Y(n8533));
  AOI21X1 g06854(.A0(n7317), .A1(n8337), .B0(n8396), .Y(n8534));
  XOR2X1  g06855(.A(n7370), .B(P2_REG2_REG_17__SCAN_IN), .Y(n8535));
  OAI21X1 g06856(.A0(n7317), .A1(n8337), .B0(n8535), .Y(n8536));
  OAI21X1 g06857(.A0(n8536), .A1(n8534), .B0(n8533), .Y(n8537));
  NOR2X1  g06858(.A(n8537), .B(n8498), .Y(n8538));
  INVX1   g06859(.A(n8475), .Y(n8539));
  NOR2X1  g06860(.A(n7317), .B(n8418), .Y(n8540));
  AOI21X1 g06861(.A0(n7371), .A1(P2_REG1_REG_17__SCAN_IN), .B0(n8420), .Y(n8541));
  OAI21X1 g06862(.A0(n8540), .A1(n8539), .B0(n8541), .Y(n8542));
  NOR2X1  g06863(.A(n7318), .B(P2_REG1_REG_16__SCAN_IN), .Y(n8543));
  XOR2X1  g06864(.A(n7370), .B(n7357), .Y(n8544));
  NOR2X1  g06865(.A(n8544), .B(n8540), .Y(n8545));
  OAI21X1 g06866(.A0(n8475), .A1(n8543), .B0(n8545), .Y(n8546));
  NAND2X1 g06867(.A(n8546), .B(n8542), .Y(n8547));
  OAI22X1 g06868(.A0(n6473), .A1(n7370), .B0(n6469), .B1(n8547), .Y(n8548));
  OAI21X1 g06869(.A0(n8548), .A1(n8538), .B0(n8336), .Y(n8549));
  NOR2X1  g06870(.A(n8547), .B(n8496), .Y(n8550));
  OAI22X1 g06871(.A0(n8498), .A1(n8537), .B0(n7370), .B1(n6473), .Y(n8551));
  OAI21X1 g06872(.A0(n8551), .A1(n8550), .B0(P2_U3947), .Y(n8552));
  NOR2X1  g06873(.A(n8547), .B(n8504), .Y(n8553));
  OAI22X1 g06874(.A0(P2_STATE_REG_SCAN_IN), .A1(n7353), .B0(n1525), .B1(n8501), .Y(n8554));
  AOI21X1 g06875(.A0(n8509), .A1(n7371), .B0(n8554), .Y(n8555));
  OAI21X1 g06876(.A0(n8537), .A1(n8507), .B0(n8555), .Y(n8556));
  NOR2X1  g06877(.A(n8556), .B(n8553), .Y(n8557));
  NAND3X1 g06878(.A(n8557), .B(n8552), .C(n8549), .Y(P2_U3231));
  XOR2X1  g06879(.A(n7317), .B(n8337), .Y(n8559));
  NOR2X1  g06880(.A(n8559), .B(n8396), .Y(n8561));
  AOI21X1 g06881(.A0(n8559), .A1(n8396), .B0(n8561), .Y(n8562));
  NOR2X1  g06882(.A(n8562), .B(n8498), .Y(n8563));
  XOR2X1  g06883(.A(n7317), .B(n8418), .Y(n8564));
  NOR2X1  g06884(.A(n8564), .B(n8475), .Y(n8566));
  AOI21X1 g06885(.A0(n8564), .A1(n8475), .B0(n8566), .Y(n8567));
  OAI22X1 g06886(.A0(n6473), .A1(n7317), .B0(n6469), .B1(n8567), .Y(n8568));
  OAI21X1 g06887(.A0(n8568), .A1(n8563), .B0(n8336), .Y(n8569));
  NOR2X1  g06888(.A(n8567), .B(n8496), .Y(n8570));
  OAI22X1 g06889(.A0(n8498), .A1(n8562), .B0(n7317), .B1(n6473), .Y(n8571));
  OAI21X1 g06890(.A0(n8571), .A1(n8570), .B0(P2_U3947), .Y(n8572));
  NOR2X1  g06891(.A(n8567), .B(n8504), .Y(n8573));
  OAI22X1 g06892(.A0(P2_STATE_REG_SCAN_IN), .A1(n7298), .B0(n1610), .B1(n8501), .Y(n8574));
  AOI21X1 g06893(.A0(n8509), .A1(n7318), .B0(n8574), .Y(n8575));
  OAI21X1 g06894(.A0(n8562), .A1(n8507), .B0(n8575), .Y(n8576));
  NOR2X1  g06895(.A(n8576), .B(n8573), .Y(n8577));
  NAND3X1 g06896(.A(n8577), .B(n8572), .C(n8569), .Y(P2_U3230));
  XOR2X1  g06897(.A(n7262), .B(P2_REG2_REG_15__SCAN_IN), .Y(n8579));
  XOR2X1  g06898(.A(n8579), .B(n8394), .Y(n8580));
  INVX1   g06899(.A(n8580), .Y(n8581));
  NOR2X1  g06900(.A(n8581), .B(n8498), .Y(n8582));
  XOR2X1  g06901(.A(n7262), .B(P2_REG1_REG_15__SCAN_IN), .Y(n8583));
  XOR2X1  g06902(.A(n8583), .B(n8473), .Y(n8584));
  INVX1   g06903(.A(n8584), .Y(n8585));
  OAI22X1 g06904(.A0(n6473), .A1(n7262), .B0(n6469), .B1(n8585), .Y(n8586));
  OAI21X1 g06905(.A0(n8586), .A1(n8582), .B0(n8336), .Y(n8587));
  AOI22X1 g06906(.A0(n8409), .A1(n8580), .B0(n7263), .B1(n6481), .Y(n8588));
  OAI21X1 g06907(.A0(n8585), .A1(n8496), .B0(n8588), .Y(n8589));
  NAND2X1 g06908(.A(n8589), .B(P2_U3947), .Y(n8590));
  NAND2X1 g06909(.A(n8584), .B(n8503), .Y(n8591));
  AOI22X1 g06910(.A0(P2_U3088), .A1(P2_REG3_REG_15__SCAN_IN), .B0(P2_ADDR_REG_15__SCAN_IN), .B1(n8502), .Y(n8592));
  OAI21X1 g06911(.A0(n8510), .A1(n7262), .B0(n8592), .Y(n8593));
  AOI21X1 g06912(.A0(n8580), .A1(n8506), .B0(n8593), .Y(n8594));
  NAND4X1 g06913(.A(n8591), .B(n8590), .C(n8587), .D(n8594), .Y(P2_U3229));
  XOR2X1  g06914(.A(n7215), .B(P2_REG2_REG_14__SCAN_IN), .Y(n8596));
  XOR2X1  g06915(.A(n8596), .B(n8392), .Y(n8597));
  INVX1   g06916(.A(n8597), .Y(n8598));
  NOR2X1  g06917(.A(n8598), .B(n8498), .Y(n8599));
  XOR2X1  g06918(.A(n7215), .B(P2_REG1_REG_14__SCAN_IN), .Y(n8600));
  XOR2X1  g06919(.A(n8600), .B(n8472), .Y(n8601));
  OAI22X1 g06920(.A0(n6473), .A1(n7215), .B0(n6469), .B1(n8601), .Y(n8602));
  OAI21X1 g06921(.A0(n8602), .A1(n8599), .B0(n8336), .Y(n8603));
  AOI22X1 g06922(.A0(n8409), .A1(n8597), .B0(n7216), .B1(n6481), .Y(n8604));
  OAI21X1 g06923(.A0(n8601), .A1(n8496), .B0(n8604), .Y(n8605));
  AOI22X1 g06924(.A0(P2_U3088), .A1(P2_REG3_REG_14__SCAN_IN), .B0(P2_ADDR_REG_14__SCAN_IN), .B1(n8502), .Y(n8606));
  OAI21X1 g06925(.A0(n8510), .A1(n7215), .B0(n8606), .Y(n8607));
  AOI21X1 g06926(.A0(n8597), .A1(n8506), .B0(n8607), .Y(n8608));
  OAI21X1 g06927(.A0(n8601), .A1(n8504), .B0(n8608), .Y(n8609));
  AOI21X1 g06928(.A0(n8605), .A1(P2_U3947), .B0(n8609), .Y(n8610));
  NAND2X1 g06929(.A(n8610), .B(n8603), .Y(P2_U3228));
  NAND2X1 g06930(.A(n7060), .B(n8344), .Y(n8612));
  AOI21X1 g06931(.A0(n8612), .A1(n8390), .B0(n8345), .Y(n8613));
  INVX1   g06932(.A(n8613), .Y(n8614));
  AOI21X1 g06933(.A0(n7162), .A1(P2_REG2_REG_13__SCAN_IN), .B0(n8348), .Y(n8615));
  OAI21X1 g06934(.A0(n8614), .A1(n8349), .B0(n8615), .Y(n8616));
  NOR2X1  g06935(.A(n7113), .B(P2_REG2_REG_12__SCAN_IN), .Y(n8617));
  XOR2X1  g06936(.A(n7161), .B(n8342), .Y(n8618));
  NOR2X1  g06937(.A(n8618), .B(n8349), .Y(n8619));
  OAI21X1 g06938(.A0(n8613), .A1(n8617), .B0(n8619), .Y(n8620));
  NAND2X1 g06939(.A(n8620), .B(n8616), .Y(n8621));
  NOR2X1  g06940(.A(n8621), .B(n8498), .Y(n8622));
  NOR2X1  g06941(.A(n7061), .B(P2_REG1_REG_11__SCAN_IN), .Y(n8623));
  OAI21X1 g06942(.A0(n8623), .A1(n8470), .B0(n8425), .Y(n8624));
  AOI21X1 g06943(.A0(n7162), .A1(P2_REG1_REG_13__SCAN_IN), .B0(n8429), .Y(n8625));
  OAI21X1 g06944(.A0(n8624), .A1(n8430), .B0(n8625), .Y(n8626));
  OAI21X1 g06945(.A0(n7113), .A1(P2_REG1_REG_12__SCAN_IN), .B0(n8624), .Y(n8627));
  XOR2X1  g06946(.A(n7161), .B(n8427), .Y(n8628));
  NOR2X1  g06947(.A(n8628), .B(n8430), .Y(n8629));
  NAND2X1 g06948(.A(n8629), .B(n8627), .Y(n8630));
  NAND2X1 g06949(.A(n8630), .B(n8626), .Y(n8631));
  OAI22X1 g06950(.A0(n6473), .A1(n7161), .B0(n6469), .B1(n8631), .Y(n8632));
  OAI21X1 g06951(.A0(n8632), .A1(n8622), .B0(n8336), .Y(n8633));
  NOR2X1  g06952(.A(n8631), .B(n8496), .Y(n8634));
  OAI22X1 g06953(.A0(n8498), .A1(n8621), .B0(n7161), .B1(n6473), .Y(n8635));
  OAI21X1 g06954(.A0(n8635), .A1(n8634), .B0(P2_U3947), .Y(n8636));
  NOR2X1  g06955(.A(n8631), .B(n8504), .Y(n8637));
  NOR2X1  g06956(.A(n8621), .B(n8507), .Y(n8638));
  AOI22X1 g06957(.A0(P2_U3088), .A1(P2_REG3_REG_13__SCAN_IN), .B0(P2_ADDR_REG_13__SCAN_IN), .B1(n8502), .Y(n8639));
  OAI21X1 g06958(.A0(n8510), .A1(n7161), .B0(n8639), .Y(n8640));
  NOR3X1  g06959(.A(n8640), .B(n8638), .C(n8637), .Y(n8641));
  NAND3X1 g06960(.A(n8641), .B(n8636), .C(n8633), .Y(P2_U3227));
  XOR2X1  g06961(.A(n7112), .B(n8172), .Y(n8643));
  NOR2X1  g06962(.A(n8643), .B(n8613), .Y(n8645));
  AOI21X1 g06963(.A0(n8643), .A1(n8613), .B0(n8645), .Y(n8646));
  NOR2X1  g06964(.A(n8646), .B(n8498), .Y(n8647));
  XOR2X1  g06965(.A(n7112), .B(P2_REG1_REG_12__SCAN_IN), .Y(n8648));
  NOR2X1  g06966(.A(n8648), .B(n8624), .Y(n8649));
  AOI21X1 g06967(.A0(n8648), .A1(n8624), .B0(n8649), .Y(n8651));
  OAI22X1 g06968(.A0(n6473), .A1(n7112), .B0(n6469), .B1(n8651), .Y(n8652));
  OAI21X1 g06969(.A0(n8652), .A1(n8647), .B0(n8336), .Y(n8653));
  NOR2X1  g06970(.A(n8651), .B(n8496), .Y(n8654));
  OAI22X1 g06971(.A0(n8498), .A1(n8646), .B0(n7112), .B1(n6473), .Y(n8655));
  OAI21X1 g06972(.A0(n8655), .A1(n8654), .B0(P2_U3947), .Y(n8656));
  NOR2X1  g06973(.A(n8651), .B(n8504), .Y(n8657));
  NOR2X1  g06974(.A(n8646), .B(n8507), .Y(n8658));
  AOI22X1 g06975(.A0(P2_U3088), .A1(P2_REG3_REG_12__SCAN_IN), .B0(P2_ADDR_REG_12__SCAN_IN), .B1(n8502), .Y(n8659));
  OAI21X1 g06976(.A0(n8510), .A1(n7112), .B0(n8659), .Y(n8660));
  NOR3X1  g06977(.A(n8660), .B(n8658), .C(n8657), .Y(n8661));
  NAND3X1 g06978(.A(n8661), .B(n8656), .C(n8653), .Y(P2_U3226));
  NOR2X1  g06979(.A(n6473), .B(n7060), .Y(n8663));
  XOR2X1  g06980(.A(n7060), .B(P2_REG1_REG_11__SCAN_IN), .Y(n8664));
  NOR2X1  g06981(.A(n8664), .B(n8469), .Y(n8665));
  AOI21X1 g06982(.A0(n8664), .A1(n8469), .B0(n8665), .Y(n8667));
  XOR2X1  g06983(.A(n7060), .B(n8344), .Y(n8668));
  AOI21X1 g06984(.A0(n8612), .A1(n8346), .B0(n8389), .Y(n8669));
  AOI21X1 g06985(.A0(n8668), .A1(n8389), .B0(n8669), .Y(n8670));
  OAI22X1 g06986(.A0(n8667), .A1(n6469), .B0(n8498), .B1(n8670), .Y(n8671));
  OAI21X1 g06987(.A0(n8671), .A1(n8663), .B0(n8336), .Y(n8672));
  NOR2X1  g06988(.A(n8667), .B(n8496), .Y(n8673));
  OAI22X1 g06989(.A0(n8498), .A1(n8670), .B0(n7060), .B1(n6473), .Y(n8674));
  OAI21X1 g06990(.A0(n8674), .A1(n8673), .B0(P2_U3947), .Y(n8675));
  AOI22X1 g06991(.A0(P2_U3088), .A1(P2_REG3_REG_11__SCAN_IN), .B0(P2_ADDR_REG_11__SCAN_IN), .B1(n8502), .Y(n8676));
  OAI21X1 g06992(.A0(n8670), .A1(n8507), .B0(n8676), .Y(n8677));
  OAI22X1 g06993(.A0(n8510), .A1(n7060), .B0(n8504), .B1(n8667), .Y(n8678));
  NOR2X1  g06994(.A(n8678), .B(n8677), .Y(n8679));
  NAND3X1 g06995(.A(n8679), .B(n8675), .C(n8672), .Y(P2_U3225));
  NOR2X1  g06996(.A(n6473), .B(n7001), .Y(n8681));
  NAND2X1 g06997(.A(n7002), .B(P2_REG1_REG_10__SCAN_IN), .Y(n8682));
  NOR2X1  g06998(.A(n6907), .B(P2_REG1_REG_8__SCAN_IN), .Y(n8683));
  NOR2X1  g06999(.A(n8683), .B(n8467), .Y(n8684));
  AOI21X1 g07000(.A0(n6907), .A1(P2_REG1_REG_8__SCAN_IN), .B0(n8684), .Y(n8685));
  OAI21X1 g07001(.A0(n6953), .A1(n8435), .B0(n8685), .Y(n8686));
  NAND3X1 g07002(.A(n8686), .B(n8682), .C(n8436), .Y(n8687));
  AOI21X1 g07003(.A0(n6953), .A1(n8435), .B0(n8685), .Y(n8688));
  AOI22X1 g07004(.A0(n6954), .A1(P2_REG1_REG_9__SCAN_IN), .B0(n8434), .B1(n7002), .Y(n8689));
  OAI21X1 g07005(.A0(n7002), .A1(n8434), .B0(n8689), .Y(n8690));
  OAI21X1 g07006(.A0(n8690), .A1(n8688), .B0(n8687), .Y(n8691));
  NAND2X1 g07007(.A(n7002), .B(P2_REG2_REG_10__SCAN_IN), .Y(n8692));
  AOI21X1 g07008(.A0(n8386), .A1(n8384), .B0(n8354), .Y(n8693));
  OAI21X1 g07009(.A0(n6953), .A1(n8355), .B0(n8693), .Y(n8694));
  NAND3X1 g07010(.A(n8694), .B(n8692), .C(n8356), .Y(n8695));
  AOI21X1 g07011(.A0(n6953), .A1(n8355), .B0(n8693), .Y(n8696));
  AOI22X1 g07012(.A0(n6954), .A1(P2_REG2_REG_9__SCAN_IN), .B0(n8352), .B1(n7002), .Y(n8697));
  OAI21X1 g07013(.A0(n7002), .A1(n8352), .B0(n8697), .Y(n8698));
  OAI21X1 g07014(.A0(n8698), .A1(n8696), .B0(n8695), .Y(n8699));
  OAI22X1 g07015(.A0(n8691), .A1(n6469), .B0(n8498), .B1(n8699), .Y(n8700));
  OAI21X1 g07016(.A0(n8700), .A1(n8681), .B0(n8336), .Y(n8701));
  NOR2X1  g07017(.A(n8691), .B(n8496), .Y(n8702));
  OAI22X1 g07018(.A0(n8498), .A1(n8699), .B0(n7001), .B1(n6473), .Y(n8703));
  OAI21X1 g07019(.A0(n8703), .A1(n8702), .B0(P2_U3947), .Y(n8704));
  AOI22X1 g07020(.A0(P2_U3088), .A1(P2_REG3_REG_10__SCAN_IN), .B0(P2_ADDR_REG_10__SCAN_IN), .B1(n8502), .Y(n8705));
  OAI21X1 g07021(.A0(n8699), .A1(n8507), .B0(n8705), .Y(n8706));
  OAI22X1 g07022(.A0(n8510), .A1(n7001), .B0(n8504), .B1(n8691), .Y(n8707));
  NOR2X1  g07023(.A(n8707), .B(n8706), .Y(n8708));
  NAND3X1 g07024(.A(n8708), .B(n8704), .C(n8701), .Y(P2_U3224));
  NOR2X1  g07025(.A(n6473), .B(n6953), .Y(n8710));
  XOR2X1  g07026(.A(n6953), .B(n8435), .Y(n8711));
  NOR2X1  g07027(.A(n8711), .B(n8685), .Y(n8713));
  AOI21X1 g07028(.A0(n8711), .A1(n8685), .B0(n8713), .Y(n8714));
  XOR2X1  g07029(.A(n6953), .B(n8355), .Y(n8715));
  NOR2X1  g07030(.A(n8715), .B(n8693), .Y(n8717));
  AOI21X1 g07031(.A0(n8715), .A1(n8693), .B0(n8717), .Y(n8718));
  OAI22X1 g07032(.A0(n8714), .A1(n6469), .B0(n8498), .B1(n8718), .Y(n8719));
  OAI21X1 g07033(.A0(n8719), .A1(n8710), .B0(n8336), .Y(n8720));
  NOR2X1  g07034(.A(n8714), .B(n8496), .Y(n8721));
  OAI22X1 g07035(.A0(n8498), .A1(n8718), .B0(n6953), .B1(n6473), .Y(n8722));
  OAI21X1 g07036(.A0(n8722), .A1(n8721), .B0(P2_U3947), .Y(n8723));
  AOI22X1 g07037(.A0(P2_U3088), .A1(P2_REG3_REG_9__SCAN_IN), .B0(P2_ADDR_REG_9__SCAN_IN), .B1(n8502), .Y(n8724));
  OAI21X1 g07038(.A0(n8718), .A1(n8507), .B0(n8724), .Y(n8725));
  OAI22X1 g07039(.A0(n8510), .A1(n6953), .B0(n8504), .B1(n8714), .Y(n8726));
  NOR2X1  g07040(.A(n8726), .B(n8725), .Y(n8727));
  NAND3X1 g07041(.A(n8727), .B(n8723), .C(n8720), .Y(P2_U3223));
  NOR2X1  g07042(.A(n6473), .B(n6906), .Y(n8729));
  XOR2X1  g07043(.A(n6906), .B(P2_REG1_REG_8__SCAN_IN), .Y(n8730));
  NOR2X1  g07044(.A(n8730), .B(n8466), .Y(n8731));
  AOI21X1 g07045(.A0(n8730), .A1(n8466), .B0(n8731), .Y(n8733));
  XOR2X1  g07046(.A(n6906), .B(P2_REG2_REG_8__SCAN_IN), .Y(n8734));
  NOR2X1  g07047(.A(n8734), .B(n8384), .Y(n8735));
  AOI21X1 g07048(.A0(n8734), .A1(n8384), .B0(n8735), .Y(n8737));
  OAI22X1 g07049(.A0(n8733), .A1(n6469), .B0(n8498), .B1(n8737), .Y(n8738));
  OAI21X1 g07050(.A0(n8738), .A1(n8729), .B0(n8336), .Y(n8739));
  NOR2X1  g07051(.A(n8733), .B(n8496), .Y(n8740));
  OAI22X1 g07052(.A0(n8498), .A1(n8737), .B0(n6906), .B1(n6473), .Y(n8741));
  OAI21X1 g07053(.A0(n8741), .A1(n8740), .B0(P2_U3947), .Y(n8742));
  AOI22X1 g07054(.A0(P2_U3088), .A1(P2_REG3_REG_8__SCAN_IN), .B0(P2_ADDR_REG_8__SCAN_IN), .B1(n8502), .Y(n8743));
  OAI22X1 g07055(.A0(n8733), .A1(n8504), .B0(n8507), .B1(n8737), .Y(n8744));
  AOI21X1 g07056(.A0(n8509), .A1(n6907), .B0(n8744), .Y(n8745));
  NAND4X1 g07057(.A(n8743), .B(n8742), .C(n8739), .D(n8745), .Y(P2_U3222));
  NOR2X1  g07058(.A(n6473), .B(n6848), .Y(n8747));
  NOR2X1  g07059(.A(n6794), .B(n6780), .Y(n8748));
  AOI21X1 g07060(.A0(n6849), .A1(P2_REG1_REG_7__SCAN_IN), .B0(n8443), .Y(n8749));
  OAI21X1 g07061(.A0(n8748), .A1(n8461), .B0(n8749), .Y(n8750));
  AOI22X1 g07062(.A0(n8456), .A1(n8460), .B0(n6794), .B1(n6780), .Y(n8751));
  AOI21X1 g07063(.A0(n6849), .A1(n8441), .B0(n8748), .Y(n8752));
  OAI21X1 g07064(.A0(n6849), .A1(n8441), .B0(n8752), .Y(n8753));
  OAI21X1 g07065(.A0(n8753), .A1(n8751), .B0(n8750), .Y(n8754));
  NOR2X1  g07066(.A(n6794), .B(n6777), .Y(n8755));
  INVX1   g07067(.A(n8360), .Y(n8756));
  AOI21X1 g07068(.A0(n6849), .A1(P2_REG2_REG_7__SCAN_IN), .B0(n8756), .Y(n8757));
  OAI21X1 g07069(.A0(n8755), .A1(n8379), .B0(n8757), .Y(n8758));
  AOI22X1 g07070(.A0(n8374), .A1(n8378), .B0(n6794), .B1(n6777), .Y(n8759));
  AOI21X1 g07071(.A0(n6849), .A1(n8133), .B0(n8755), .Y(n8760));
  OAI21X1 g07072(.A0(n6849), .A1(n8133), .B0(n8760), .Y(n8761));
  OAI21X1 g07073(.A0(n8761), .A1(n8759), .B0(n8758), .Y(n8762));
  OAI22X1 g07074(.A0(n8754), .A1(n6469), .B0(n8498), .B1(n8762), .Y(n8763));
  OAI21X1 g07075(.A0(n8763), .A1(n8747), .B0(n8336), .Y(n8764));
  INVX1   g07076(.A(n8762), .Y(n8765));
  NAND2X1 g07077(.A(n8765), .B(n8506), .Y(n8766));
  AOI22X1 g07078(.A0(n8409), .A1(n8765), .B0(n6849), .B1(n6481), .Y(n8767));
  OAI21X1 g07079(.A0(n8754), .A1(n8496), .B0(n8767), .Y(n8768));
  OAI22X1 g07080(.A0(P2_STATE_REG_SCAN_IN), .A1(n6889), .B0(n1632), .B1(n8501), .Y(n8769));
  AOI21X1 g07081(.A0(n8768), .A1(P2_U3947), .B0(n8769), .Y(n8770));
  INVX1   g07082(.A(n8754), .Y(n8771));
  AOI22X1 g07083(.A0(n8509), .A1(n6849), .B0(n8503), .B1(n8771), .Y(n8772));
  NAND4X1 g07084(.A(n8770), .B(n8766), .C(n8764), .D(n8772), .Y(P2_U3221));
  NOR2X1  g07085(.A(n6473), .B(n6794), .Y(n8774));
  XOR2X1  g07086(.A(n6794), .B(P2_REG1_REG_6__SCAN_IN), .Y(n8775));
  NOR2X1  g07087(.A(n8775), .B(n8461), .Y(n8776));
  AOI21X1 g07088(.A0(n8775), .A1(n8461), .B0(n8776), .Y(n8779));
  XOR2X1  g07089(.A(n6794), .B(P2_REG2_REG_6__SCAN_IN), .Y(n8780));
  NOR2X1  g07090(.A(n8780), .B(n8379), .Y(n8781));
  XOR2X1  g07091(.A(n6794), .B(n6777), .Y(n8782));
  AOI21X1 g07092(.A0(n8378), .A1(n8374), .B0(n8782), .Y(n8783));
  NOR2X1  g07093(.A(n8783), .B(n8781), .Y(n8784));
  OAI22X1 g07094(.A0(n8779), .A1(n6469), .B0(n8498), .B1(n8784), .Y(n8785));
  OAI21X1 g07095(.A0(n8785), .A1(n8774), .B0(n8336), .Y(n8786));
  NOR2X1  g07096(.A(n8784), .B(n8507), .Y(n8787));
  INVX1   g07097(.A(P2_U3947), .Y(n8788));
  NOR2X1  g07098(.A(n8779), .B(n8496), .Y(n8789));
  OAI22X1 g07099(.A0(n8498), .A1(n8784), .B0(n6794), .B1(n6473), .Y(n8790));
  NOR2X1  g07100(.A(n8790), .B(n8789), .Y(n8791));
  AOI22X1 g07101(.A0(P2_U3088), .A1(P2_REG3_REG_6__SCAN_IN), .B0(P2_ADDR_REG_6__SCAN_IN), .B1(n8502), .Y(n8792));
  OAI21X1 g07102(.A0(n8791), .A1(n8788), .B0(n8792), .Y(n8793));
  OAI22X1 g07103(.A0(n8510), .A1(n6794), .B0(n8504), .B1(n8779), .Y(n8794));
  NOR3X1  g07104(.A(n8794), .B(n8793), .C(n8787), .Y(n8795));
  NAND2X1 g07105(.A(n8795), .B(n8786), .Y(P2_U3220));
  NOR2X1  g07106(.A(n6473), .B(n6747), .Y(n8797));
  INVX1   g07107(.A(n8448), .Y(n8798));
  NOR2X1  g07108(.A(n8798), .B(n8445), .Y(n8799));
  NOR2X1  g07109(.A(n6598), .B(P2_REG1_REG_2__SCAN_IN), .Y(n8800));
  NOR3X1  g07110(.A(n8800), .B(n6551), .C(n6539), .Y(n8801));
  AOI21X1 g07111(.A0(n6598), .A1(P2_REG1_REG_2__SCAN_IN), .B0(n8801), .Y(n8802));
  NOR2X1  g07112(.A(n8802), .B(n8452), .Y(n8803));
  NOR4X1  g07113(.A(n8799), .B(n8457), .C(n8451), .D(n8803), .Y(n8804));
  OAI21X1 g07114(.A0(n6747), .A1(n6728), .B0(n8444), .Y(n8805));
  NOR3X1  g07115(.A(n8803), .B(n8799), .C(n8451), .Y(n8806));
  AOI21X1 g07116(.A0(n8361), .A1(n6681), .B0(n8806), .Y(n8807));
  INVX1   g07117(.A(n6747), .Y(n8808));
  AOI22X1 g07118(.A0(n6701), .A1(P2_REG1_REG_4__SCAN_IN), .B0(n6728), .B1(n8808), .Y(n8809));
  OAI21X1 g07119(.A0(n8808), .A1(n6728), .B0(n8809), .Y(n8810));
  OAI22X1 g07120(.A0(n8807), .A1(n8810), .B0(n8805), .B1(n8804), .Y(n8811));
  INVX1   g07121(.A(n8366), .Y(n8812));
  NOR2X1  g07122(.A(n8812), .B(n8363), .Y(n8813));
  NOR2X1  g07123(.A(n6598), .B(P2_REG2_REG_2__SCAN_IN), .Y(n8814));
  NOR3X1  g07124(.A(n8814), .B(n6551), .C(n6536), .Y(n8815));
  AOI21X1 g07125(.A0(n6598), .A1(P2_REG2_REG_2__SCAN_IN), .B0(n8815), .Y(n8816));
  NOR2X1  g07126(.A(n8816), .B(n8370), .Y(n8817));
  NOR4X1  g07127(.A(n8813), .B(n8375), .C(n8369), .D(n8817), .Y(n8818));
  OAI21X1 g07128(.A0(n6747), .A1(n6725), .B0(n8362), .Y(n8819));
  NOR3X1  g07129(.A(n8817), .B(n8813), .C(n8369), .Y(n8820));
  AOI21X1 g07130(.A0(n8361), .A1(n6678), .B0(n8820), .Y(n8821));
  AOI22X1 g07131(.A0(n6701), .A1(P2_REG2_REG_4__SCAN_IN), .B0(n6725), .B1(n8808), .Y(n8822));
  OAI21X1 g07132(.A0(n8808), .A1(n6725), .B0(n8822), .Y(n8823));
  OAI22X1 g07133(.A0(n8821), .A1(n8823), .B0(n8819), .B1(n8818), .Y(n8824));
  OAI22X1 g07134(.A0(n8811), .A1(n6469), .B0(n8498), .B1(n8824), .Y(n8825));
  OAI21X1 g07135(.A0(n8825), .A1(n8797), .B0(n8336), .Y(n8826));
  INVX1   g07136(.A(n8824), .Y(n8827));
  NAND2X1 g07137(.A(n8827), .B(n8506), .Y(n8828));
  AOI22X1 g07138(.A0(n8409), .A1(n8827), .B0(n8808), .B1(n6481), .Y(n8829));
  OAI21X1 g07139(.A0(n8811), .A1(n8496), .B0(n8829), .Y(n8830));
  OAI22X1 g07140(.A0(P2_STATE_REG_SCAN_IN), .A1(n6782), .B0(n1641), .B1(n8501), .Y(n8831));
  AOI21X1 g07141(.A0(n8830), .A1(P2_U3947), .B0(n8831), .Y(n8832));
  INVX1   g07142(.A(n8811), .Y(n8833));
  AOI22X1 g07143(.A0(n8509), .A1(n8808), .B0(n8503), .B1(n8833), .Y(n8834));
  NAND4X1 g07144(.A(n8832), .B(n8828), .C(n8826), .D(n8834), .Y(P2_U3219));
  NOR2X1  g07145(.A(n6473), .B(n8361), .Y(n8836));
  XOR2X1  g07146(.A(n6701), .B(P2_REG1_REG_4__SCAN_IN), .Y(n8837));
  NOR2X1  g07147(.A(n8837), .B(n8806), .Y(n8839));
  AOI21X1 g07148(.A0(n8837), .A1(n8806), .B0(n8839), .Y(n8840));
  XOR2X1  g07149(.A(n6701), .B(P2_REG2_REG_4__SCAN_IN), .Y(n8841));
  NOR2X1  g07150(.A(n8841), .B(n8820), .Y(n8843));
  AOI21X1 g07151(.A0(n8841), .A1(n8820), .B0(n8843), .Y(n8844));
  OAI22X1 g07152(.A0(n8840), .A1(n6469), .B0(n8498), .B1(n8844), .Y(n8845));
  OAI21X1 g07153(.A0(n8845), .A1(n8836), .B0(n8336), .Y(n8846));
  INVX1   g07154(.A(n8844), .Y(n8847));
  NAND2X1 g07155(.A(n8847), .B(n8506), .Y(n8848));
  INVX1   g07156(.A(n8840), .Y(n8849));
  OAI22X1 g07157(.A0(n8498), .A1(n8844), .B0(n8361), .B1(n6473), .Y(n8850));
  AOI21X1 g07158(.A0(n8849), .A1(n8495), .B0(n8850), .Y(n8851));
  OAI22X1 g07159(.A0(n8788), .A1(n8851), .B0(P2_STATE_REG_SCAN_IN), .B1(n6682), .Y(n8852));
  AOI21X1 g07160(.A0(n8502), .A1(P2_ADDR_REG_4__SCAN_IN), .B0(n8852), .Y(n8853));
  AOI22X1 g07161(.A0(n8509), .A1(n6701), .B0(n8503), .B1(n8849), .Y(n8854));
  NAND4X1 g07162(.A(n8853), .B(n8848), .C(n8846), .D(n8854), .Y(P2_U3218));
  NOR2X1  g07163(.A(n6473), .B(n6643), .Y(n8856));
  OAI21X1 g07164(.A0(n8798), .A1(n8800), .B0(n8802), .Y(n8857));
  XOR2X1  g07165(.A(n6643), .B(P2_REG1_REG_3__SCAN_IN), .Y(n8858));
  OAI21X1 g07166(.A0(n8451), .A1(n8452), .B0(n8857), .Y(n8859));
  OAI21X1 g07167(.A0(n8858), .A1(n8857), .B0(n8859), .Y(n8860));
  INVX1   g07168(.A(n8860), .Y(n8861));
  OAI21X1 g07169(.A0(n8812), .A1(n8814), .B0(n8816), .Y(n8862));
  XOR2X1  g07170(.A(n6643), .B(P2_REG2_REG_3__SCAN_IN), .Y(n8863));
  OAI21X1 g07171(.A0(n8369), .A1(n8370), .B0(n8862), .Y(n8864));
  OAI21X1 g07172(.A0(n8863), .A1(n8862), .B0(n8864), .Y(n8865));
  NAND3X1 g07173(.A(n8865), .B(n8415), .C(n8409), .Y(n8866));
  OAI21X1 g07174(.A0(n8861), .A1(n6469), .B0(n8866), .Y(n8867));
  OAI21X1 g07175(.A0(n8867), .A1(n8856), .B0(n8336), .Y(n8868));
  AOI22X1 g07176(.A0(n8409), .A1(n8865), .B0(n6644), .B1(n6481), .Y(n8869));
  OAI21X1 g07177(.A0(n8861), .A1(n8496), .B0(n8869), .Y(n8870));
  AOI22X1 g07178(.A0(P2_U3947), .A1(n8870), .B0(P2_U3088), .B1(P2_REG3_REG_3__SCAN_IN), .Y(n8871));
  OAI21X1 g07179(.A0(n8501), .A1(n1646), .B0(n8871), .Y(n8872));
  AOI21X1 g07180(.A0(n8865), .A1(n8506), .B0(n8872), .Y(n8873));
  AOI22X1 g07181(.A0(n8509), .A1(n6644), .B0(n8503), .B1(n8860), .Y(n8874));
  NAND3X1 g07182(.A(n8874), .B(n8873), .C(n8868), .Y(P2_U3217));
  NAND3X1 g07183(.A(n8415), .B(n6598), .C(n6481), .Y(n8876));
  XOR2X1  g07184(.A(n6597), .B(P2_REG1_REG_2__SCAN_IN), .Y(n8877));
  NOR2X1  g07185(.A(n8877), .B(n8450), .Y(n8878));
  AOI21X1 g07186(.A0(n8877), .A1(n8450), .B0(n8878), .Y(n8880));
  NAND3X1 g07187(.A(n8880), .B(n8415), .C(n6480), .Y(n8881));
  XOR2X1  g07188(.A(n6597), .B(P2_REG2_REG_2__SCAN_IN), .Y(n8882));
  NOR2X1  g07189(.A(n8882), .B(n8368), .Y(n8883));
  AOI21X1 g07190(.A0(n8882), .A1(n8368), .B0(n8883), .Y(n8885));
  NAND3X1 g07191(.A(n8885), .B(n8415), .C(n8409), .Y(n8886));
  NAND3X1 g07192(.A(n8886), .B(n8881), .C(n8876), .Y(n8887));
  NAND2X1 g07193(.A(n8887), .B(n8336), .Y(n8888));
  NAND2X1 g07194(.A(n8885), .B(n8506), .Y(n8889));
  NOR2X1  g07195(.A(n8501), .B(n1647), .Y(n8890));
  NOR2X1  g07196(.A(P2_STATE_REG_SCAN_IN), .B(n6593), .Y(n8891));
  NAND2X1 g07197(.A(n8880), .B(n8495), .Y(n8892));
  AOI22X1 g07198(.A0(n8409), .A1(n8885), .B0(n6598), .B1(n6481), .Y(n8893));
  AOI21X1 g07199(.A0(n8893), .A1(n8892), .B0(n8788), .Y(n8894));
  NOR3X1  g07200(.A(n8894), .B(n8891), .C(n8890), .Y(n8895));
  AOI22X1 g07201(.A0(n8509), .A1(n6598), .B0(n8503), .B1(n8880), .Y(n8896));
  NAND4X1 g07202(.A(n8895), .B(n8889), .C(n8888), .D(n8896), .Y(P2_U3216));
  NOR2X1  g07203(.A(n6473), .B(n6551), .Y(n8898));
  XOR2X1  g07204(.A(n6551), .B(n6539), .Y(n8899));
  XOR2X1  g07205(.A(n8899), .B(n8447), .Y(n8900));
  XOR2X1  g07206(.A(n6551), .B(n6536), .Y(n8901));
  XOR2X1  g07207(.A(n8901), .B(n8365), .Y(n8902));
  OAI22X1 g07208(.A0(n8900), .A1(n6469), .B0(n8498), .B1(n8902), .Y(n8903));
  OAI21X1 g07209(.A0(n8903), .A1(n8898), .B0(n8336), .Y(n8904));
  INVX1   g07210(.A(n8902), .Y(n8905));
  AOI22X1 g07211(.A0(n8409), .A1(n8905), .B0(n6552), .B1(n6481), .Y(n8906));
  OAI21X1 g07212(.A0(n8900), .A1(n8496), .B0(n8906), .Y(n8907));
  AOI22X1 g07213(.A0(P2_U3947), .A1(n8907), .B0(P2_U3088), .B1(P2_REG3_REG_1__SCAN_IN), .Y(n8908));
  OAI21X1 g07214(.A0(n8501), .A1(n1656), .B0(n8908), .Y(n8909));
  AOI21X1 g07215(.A0(n8905), .A1(n8506), .B0(n8909), .Y(n8910));
  INVX1   g07216(.A(n8900), .Y(n8911));
  AOI22X1 g07217(.A0(n8509), .A1(n6552), .B0(n8503), .B1(n8911), .Y(n8912));
  NAND3X1 g07218(.A(n8912), .B(n8910), .C(n8904), .Y(P2_U3215));
  NOR2X1  g07219(.A(n6473), .B(n6475), .Y(n8914));
  XOR2X1  g07220(.A(n6475), .B(P2_REG1_REG_0__SCAN_IN), .Y(n8915));
  XOR2X1  g07221(.A(n6475), .B(P2_REG2_REG_0__SCAN_IN), .Y(n8916));
  OAI22X1 g07222(.A0(n8915), .A1(n6469), .B0(n8498), .B1(n8916), .Y(n8917));
  OAI21X1 g07223(.A0(n8917), .A1(n8914), .B0(n8336), .Y(n8918));
  INVX1   g07224(.A(n8916), .Y(n8919));
  NAND4X1 g07225(.A(n8493), .B(P2_STATE_REG_SCAN_IN), .C(P2_ADDR_REG_0__SCAN_IN), .D(n8335), .Y(n8920));
  NOR2X1  g07226(.A(P2_STATE_REG_SCAN_IN), .B(n6496), .Y(n8921));
  AOI22X1 g07227(.A0(n8409), .A1(n8919), .B0(n6481), .B1(n6479), .Y(n8922));
  OAI21X1 g07228(.A0(n8915), .A1(n8496), .B0(n8922), .Y(n8923));
  AOI21X1 g07229(.A0(n8923), .A1(P2_U3947), .B0(n8921), .Y(n8924));
  NAND2X1 g07230(.A(n8924), .B(n8920), .Y(n8925));
  AOI21X1 g07231(.A0(n8919), .A1(n8506), .B0(n8925), .Y(n8926));
  INVX1   g07232(.A(n8915), .Y(n8927));
  AOI22X1 g07233(.A0(n8509), .A1(n6479), .B0(n8503), .B1(n8927), .Y(n8928));
  NAND3X1 g07234(.A(n8928), .B(n8926), .C(n8918), .Y(P2_U3214));
  NAND3X1 g07235(.A(n8492), .B(n6573), .C(P2_STATE_REG_SCAN_IN), .Y(n8930));
  OAI21X1 g07236(.A0(P2_U3947), .A1(n1791), .B0(n8930), .Y(P2_U3531));
  NAND3X1 g07237(.A(n8492), .B(n6569), .C(P2_STATE_REG_SCAN_IN), .Y(n8932));
  OAI21X1 g07238(.A0(P2_U3947), .A1(n1806), .B0(n8932), .Y(P2_U3532));
  NAND3X1 g07239(.A(n8492), .B(n6583), .C(P2_STATE_REG_SCAN_IN), .Y(n8934));
  OAI21X1 g07240(.A0(P2_U3947), .A1(n1832), .B0(n8934), .Y(P2_U3533));
  NAND3X1 g07241(.A(n8492), .B(n6652), .C(P2_STATE_REG_SCAN_IN), .Y(n8936));
  OAI21X1 g07242(.A0(P2_U3947), .A1(n1848), .B0(n8936), .Y(P2_U3534));
  NAND3X1 g07243(.A(n8492), .B(n6706), .C(P2_STATE_REG_SCAN_IN), .Y(n8938));
  OAI21X1 g07244(.A0(P2_U3947), .A1(n1871), .B0(n8938), .Y(P2_U3535));
  NAND3X1 g07245(.A(n8492), .B(n6745), .C(P2_STATE_REG_SCAN_IN), .Y(n8940));
  OAI21X1 g07246(.A0(P2_U3947), .A1(n1898), .B0(n8940), .Y(P2_U3536));
  NAND3X1 g07247(.A(n8492), .B(n6807), .C(P2_STATE_REG_SCAN_IN), .Y(n8942));
  OAI21X1 g07248(.A0(P2_U3947), .A1(n1927), .B0(n8942), .Y(P2_U3537));
  NAND3X1 g07249(.A(n8492), .B(n6839), .C(P2_STATE_REG_SCAN_IN), .Y(n8944));
  OAI21X1 g07250(.A0(P2_U3947), .A1(n1950), .B0(n8944), .Y(P2_U3538));
  NAND3X1 g07251(.A(n8492), .B(n6894), .C(P2_STATE_REG_SCAN_IN), .Y(n8946));
  OAI21X1 g07252(.A0(P2_U3947), .A1(n1974), .B0(n8946), .Y(P2_U3539));
  NAND3X1 g07253(.A(n8492), .B(n6944), .C(P2_STATE_REG_SCAN_IN), .Y(n8948));
  OAI21X1 g07254(.A0(P2_U3947), .A1(n1999), .B0(n8948), .Y(P2_U3540));
  NAND3X1 g07255(.A(n8492), .B(n6992), .C(P2_STATE_REG_SCAN_IN), .Y(n8950));
  OAI21X1 g07256(.A0(P2_U3947), .A1(n2018), .B0(n8950), .Y(P2_U3541));
  NAND3X1 g07257(.A(n8492), .B(n7072), .C(P2_STATE_REG_SCAN_IN), .Y(n8952));
  OAI21X1 g07258(.A0(P2_U3947), .A1(n2043), .B0(n8952), .Y(P2_U3542));
  NAND3X1 g07259(.A(n8492), .B(n7103), .C(P2_STATE_REG_SCAN_IN), .Y(n8954));
  OAI21X1 g07260(.A0(P2_U3947), .A1(n2065), .B0(n8954), .Y(P2_U3543));
  NAND3X1 g07261(.A(n8492), .B(n7154), .C(P2_STATE_REG_SCAN_IN), .Y(n8956));
  OAI21X1 g07262(.A0(P2_U3947), .A1(n2088), .B0(n8956), .Y(P2_U3544));
  NAND3X1 g07263(.A(n8492), .B(n7206), .C(P2_STATE_REG_SCAN_IN), .Y(n8958));
  OAI21X1 g07264(.A0(P2_U3947), .A1(n2109), .B0(n8958), .Y(P2_U3545));
  NAND3X1 g07265(.A(n8492), .B(n7255), .C(P2_STATE_REG_SCAN_IN), .Y(n8960));
  OAI21X1 g07266(.A0(P2_U3947), .A1(n2128), .B0(n8960), .Y(P2_U3546));
  NAND3X1 g07267(.A(n8492), .B(n7304), .C(P2_STATE_REG_SCAN_IN), .Y(n8962));
  OAI21X1 g07268(.A0(P2_U3947), .A1(n2148), .B0(n8962), .Y(P2_U3547));
  NAND3X1 g07269(.A(n8492), .B(n7368), .C(P2_STATE_REG_SCAN_IN), .Y(n8964));
  OAI21X1 g07270(.A0(P2_U3947), .A1(n2181), .B0(n8964), .Y(P2_U3548));
  NAND3X1 g07271(.A(n8492), .B(n7432), .C(P2_STATE_REG_SCAN_IN), .Y(n8966));
  OAI21X1 g07272(.A0(P2_U3947), .A1(n2199), .B0(n8966), .Y(P2_U3549));
  NAND3X1 g07273(.A(n8492), .B(n7486), .C(P2_STATE_REG_SCAN_IN), .Y(n8968));
  OAI21X1 g07274(.A0(P2_U3947), .A1(n2227), .B0(n8968), .Y(P2_U3550));
  NAND3X1 g07275(.A(n8492), .B(n7509), .C(P2_STATE_REG_SCAN_IN), .Y(n8970));
  OAI21X1 g07276(.A0(P2_U3947), .A1(n2250), .B0(n8970), .Y(P2_U3551));
  NAND3X1 g07277(.A(n8492), .B(n7557), .C(P2_STATE_REG_SCAN_IN), .Y(n8972));
  OAI21X1 g07278(.A0(P2_U3947), .A1(n2274), .B0(n8972), .Y(P2_U3552));
  NAND3X1 g07279(.A(n8492), .B(n7600), .C(P2_STATE_REG_SCAN_IN), .Y(n8974));
  OAI21X1 g07280(.A0(P2_U3947), .A1(n2289), .B0(n8974), .Y(P2_U3553));
  NAND3X1 g07281(.A(n8492), .B(n7642), .C(P2_STATE_REG_SCAN_IN), .Y(n8976));
  OAI21X1 g07282(.A0(P2_U3947), .A1(n2319), .B0(n8976), .Y(P2_U3554));
  NAND3X1 g07283(.A(n8492), .B(n7688), .C(P2_STATE_REG_SCAN_IN), .Y(n8978));
  OAI21X1 g07284(.A0(P2_U3947), .A1(n2345), .B0(n8978), .Y(P2_U3555));
  NAND3X1 g07285(.A(n8492), .B(n7734), .C(P2_STATE_REG_SCAN_IN), .Y(n8980));
  OAI21X1 g07286(.A0(P2_U3947), .A1(n2371), .B0(n8980), .Y(P2_U3556));
  NAND3X1 g07287(.A(n8492), .B(n7779), .C(P2_STATE_REG_SCAN_IN), .Y(n8982));
  OAI21X1 g07288(.A0(P2_U3947), .A1(n2389), .B0(n8982), .Y(P2_U3557));
  NAND3X1 g07289(.A(n8492), .B(n7824), .C(P2_STATE_REG_SCAN_IN), .Y(n8984));
  OAI21X1 g07290(.A0(P2_U3947), .A1(n2421), .B0(n8984), .Y(P2_U3558));
  NAND3X1 g07291(.A(n8492), .B(n7885), .C(P2_STATE_REG_SCAN_IN), .Y(n8986));
  OAI21X1 g07292(.A0(P2_U3947), .A1(n2441), .B0(n8986), .Y(P2_U3559));
  NAND3X1 g07293(.A(n8492), .B(n7931), .C(P2_STATE_REG_SCAN_IN), .Y(n8988));
  OAI21X1 g07294(.A0(P2_U3947), .A1(n2466), .B0(n8988), .Y(P2_U3560));
  INVX1   g07295(.A(n7954), .Y(n8990));
  NAND3X1 g07296(.A(n8492), .B(n8990), .C(P2_STATE_REG_SCAN_IN), .Y(n8991));
  OAI21X1 g07297(.A0(P2_U3947), .A1(n2492), .B0(n8991), .Y(P2_U3561));
  INVX1   g07298(.A(n7988), .Y(n8993));
  NAND3X1 g07299(.A(n8492), .B(n8993), .C(P2_STATE_REG_SCAN_IN), .Y(n8994));
  OAI21X1 g07300(.A0(P2_U3947), .A1(n2511), .B0(n8994), .Y(P2_U3562));
  NOR3X1  g07301(.A(n6517), .B(n6455), .C(n6449), .Y(n8996));
  NAND2X1 g07302(.A(n8996), .B(n6342), .Y(n8997));
  OAI21X1 g07303(.A0(n6460), .A1(n6458), .B0(n6455), .Y(n8998));
  NOR2X1  g07304(.A(n6526), .B(n6516), .Y(n8999));
  NAND4X1 g07305(.A(n8998), .B(n8997), .C(n6633), .D(n8999), .Y(n9000));
  NAND2X1 g07306(.A(n6452), .B(n6449), .Y(n9001));
  AOI21X1 g07307(.A0(n7988), .A1(n8990), .B0(n6451), .Y(n9004));
  NOR2X1  g07308(.A(n9004), .B(n9000), .Y(n9005));
  NOR2X1  g07309(.A(n9005), .B(n7988), .Y(n9006));
  NOR3X1  g07310(.A(n6451), .B(n8993), .C(n7954), .Y(n9007));
  XOR2X1  g07311(.A(n7988), .B(n8990), .Y(n9008));
  NAND2X1 g07312(.A(n9008), .B(n9007), .Y(n9009));
  INVX1   g07313(.A(n9009), .Y(n9010));
  NOR2X1  g07314(.A(n9010), .B(n9006), .Y(n9011));
  NAND3X1 g07315(.A(n9011), .B(n7997), .C(n7996), .Y(n9012));
  NOR4X1  g07316(.A(n6455), .B(n6452), .C(n6458), .D(n6460), .Y(n9013));
  NOR3X1  g07317(.A(n9013), .B(n9010), .C(n9006), .Y(n9014));
  AOI21X1 g07318(.A0(n9011), .A1(n6474), .B0(n9014), .Y(n9015));
  NAND2X1 g07319(.A(n9015), .B(n9012), .Y(n9016));
  INVX1   g07320(.A(n9013), .Y(n9017));
  NOR2X1  g07321(.A(n9017), .B(n7988), .Y(n9018));
  NOR2X1  g07322(.A(n6452), .B(n9000), .Y(n9019));
  NOR2X1  g07323(.A(n9019), .B(n6474), .Y(n9020));
  INVX1   g07324(.A(n9020), .Y(n9021));
  AOI21X1 g07325(.A0(n7997), .A1(n7996), .B0(n9021), .Y(n9022));
  NOR2X1  g07326(.A(n9022), .B(n9018), .Y(n9023));
  XOR2X1  g07327(.A(n9023), .B(n9016), .Y(n9024));
  NOR2X1  g07328(.A(n9017), .B(n6474), .Y(n9025));
  OAI21X1 g07329(.A0(n6328), .A1(n6327), .B0(n9025), .Y(n9026));
  INVX1   g07330(.A(n9005), .Y(n9027));
  INVX1   g07331(.A(n9007), .Y(n9028));
  NOR2X1  g07332(.A(n9028), .B(n8990), .Y(n9029));
  AOI21X1 g07333(.A0(n9027), .A1(n8990), .B0(n9029), .Y(n9030));
  NAND2X1 g07334(.A(n9030), .B(n9026), .Y(n9031));
  NAND2X1 g07335(.A(n9013), .B(n8990), .Y(n9032));
  INVX1   g07336(.A(n9019), .Y(n9033));
  NAND3X1 g07337(.A(n9033), .B(n6750), .C(n8326), .Y(n9034));
  AOI21X1 g07338(.A0(n9034), .A1(n9032), .B0(n9031), .Y(n9035));
  NAND3X1 g07339(.A(n9033), .B(n6750), .C(n6314), .Y(n9036));
  AOI22X1 g07340(.A0(n7931), .A1(n9013), .B0(n7885), .B1(n6341), .Y(n9037));
  OAI21X1 g07341(.A0(n9005), .A1(n7932), .B0(n6342), .Y(n9038));
  AOI21X1 g07342(.A0(n9007), .A1(n7931), .B0(n9038), .Y(n9039));
  OAI21X1 g07343(.A0(n9017), .A1(n7941), .B0(n9039), .Y(n9040));
  AOI21X1 g07344(.A0(n9037), .A1(n9036), .B0(n9040), .Y(n9041));
  AOI22X1 g07345(.A0(n7885), .A1(n9013), .B0(n7824), .B1(n6341), .Y(n9042));
  OAI21X1 g07346(.A0(n9019), .A1(n7924), .B0(n9042), .Y(n9043));
  AOI21X1 g07347(.A0(n9027), .A1(n7885), .B0(n6341), .Y(n9044));
  OAI21X1 g07348(.A0(n9028), .A1(n7886), .B0(n9044), .Y(n9045));
  AOI21X1 g07349(.A0(n9013), .A1(n7893), .B0(n9045), .Y(n9046));
  NAND2X1 g07350(.A(n9046), .B(n9043), .Y(n9047));
  NOR2X1  g07351(.A(n9046), .B(n9043), .Y(n9048));
  AOI22X1 g07352(.A0(n7824), .A1(n9013), .B0(n7779), .B1(n6341), .Y(n9049));
  OAI21X1 g07353(.A0(n9019), .A1(n7848), .B0(n9049), .Y(n9050));
  AOI21X1 g07354(.A0(n9027), .A1(n7824), .B0(n6341), .Y(n9051));
  OAI21X1 g07355(.A0(n9028), .A1(n7825), .B0(n9051), .Y(n9052));
  INVX1   g07356(.A(n9052), .Y(n9053));
  OAI21X1 g07357(.A0(n9017), .A1(n7848), .B0(n9053), .Y(n9054));
  INVX1   g07358(.A(n9054), .Y(n9055));
  INVX1   g07359(.A(n9049), .Y(n9056));
  AOI21X1 g07360(.A0(n9033), .A1(n7876), .B0(n9056), .Y(n9057));
  AOI22X1 g07361(.A0(n7779), .A1(n9013), .B0(n7734), .B1(n6341), .Y(n9058));
  OAI21X1 g07362(.A0(n9019), .A1(n7787), .B0(n9058), .Y(n9059));
  NOR2X1  g07363(.A(n9017), .B(n7787), .Y(n9060));
  AOI21X1 g07364(.A0(n9027), .A1(n7779), .B0(n6341), .Y(n9061));
  OAI21X1 g07365(.A0(n9028), .A1(n7780), .B0(n9061), .Y(n9062));
  NOR2X1  g07366(.A(n9062), .B(n9060), .Y(n9063));
  NAND2X1 g07367(.A(n9063), .B(n9059), .Y(n9064));
  OAI21X1 g07368(.A0(n9054), .A1(n9057), .B0(n9064), .Y(n9065));
  AOI22X1 g07369(.A0(n7734), .A1(n9013), .B0(n7688), .B1(n6341), .Y(n9066));
  OAI21X1 g07370(.A0(n9019), .A1(n7758), .B0(n9066), .Y(n9067));
  INVX1   g07371(.A(n9067), .Y(n9068));
  AOI21X1 g07372(.A0(n9027), .A1(n7734), .B0(n6341), .Y(n9069));
  OAI21X1 g07373(.A0(n9028), .A1(n7735), .B0(n9069), .Y(n9070));
  AOI21X1 g07374(.A0(n9013), .A1(n7742), .B0(n9070), .Y(n9071));
  INVX1   g07375(.A(n9071), .Y(n9072));
  NAND2X1 g07376(.A(n9072), .B(n9068), .Y(n9073));
  OAI22X1 g07377(.A0(n9065), .A1(n9073), .B0(n9055), .B1(n9050), .Y(n9074));
  OAI21X1 g07378(.A0(n9074), .A1(n9048), .B0(n9047), .Y(n9075));
  NOR4X1  g07379(.A(n9041), .B(n9035), .C(n9024), .D(n9075), .Y(n9076));
  INVX1   g07380(.A(n9018), .Y(n9077));
  OAI21X1 g07381(.A0(n6335), .A1(n6334), .B0(n9020), .Y(n9078));
  NAND4X1 g07382(.A(n9077), .B(n9015), .C(n9012), .D(n9078), .Y(n9079));
  NOR4X1  g07383(.A(n9006), .B(n6335), .C(n6334), .D(n9010), .Y(n9080));
  INVX1   g07384(.A(n9015), .Y(n9081));
  OAI22X1 g07385(.A0(n9018), .A1(n9022), .B0(n9081), .B1(n9080), .Y(n9082));
  NAND2X1 g07386(.A(n9055), .B(n9050), .Y(n9083));
  INVX1   g07387(.A(n9059), .Y(n9084));
  NOR3X1  g07388(.A(n9062), .B(n9060), .C(n9084), .Y(n9085));
  NAND2X1 g07389(.A(n9071), .B(n9067), .Y(n9086));
  AOI22X1 g07390(.A0(n7688), .A1(n9013), .B0(n7642), .B1(n6341), .Y(n9087));
  INVX1   g07391(.A(n9087), .Y(n9088));
  AOI21X1 g07392(.A0(n9033), .A1(n7695), .B0(n9088), .Y(n9089));
  AOI21X1 g07393(.A0(n9027), .A1(n7688), .B0(n6341), .Y(n9090));
  OAI21X1 g07394(.A0(n9028), .A1(n7694), .B0(n9090), .Y(n9091));
  INVX1   g07395(.A(n9091), .Y(n9092));
  OAI21X1 g07396(.A0(n9017), .A1(n7723), .B0(n9092), .Y(n9093));
  AOI22X1 g07397(.A0(n7600), .A1(n9013), .B0(n7557), .B1(n6341), .Y(n9094));
  OAI21X1 g07398(.A0(n9019), .A1(n7635), .B0(n9094), .Y(n9095));
  AOI21X1 g07399(.A0(n9027), .A1(n7600), .B0(n6341), .Y(n9096));
  OAI21X1 g07400(.A0(n9028), .A1(n7601), .B0(n9096), .Y(n9097));
  AOI21X1 g07401(.A0(n9013), .A1(n7608), .B0(n9097), .Y(n9098));
  NAND2X1 g07402(.A(n9033), .B(n7652), .Y(n9099));
  AOI22X1 g07403(.A0(n7642), .A1(n9013), .B0(n7600), .B1(n6341), .Y(n9100));
  NAND2X1 g07404(.A(n9100), .B(n9099), .Y(n9101));
  AOI21X1 g07405(.A0(n9027), .A1(n7642), .B0(n6341), .Y(n9102));
  OAI21X1 g07406(.A0(n9028), .A1(n7643), .B0(n9102), .Y(n9103));
  AOI21X1 g07407(.A0(n9013), .A1(n7652), .B0(n9103), .Y(n9104));
  AOI22X1 g07408(.A0(n9101), .A1(n9104), .B0(n9098), .B1(n9095), .Y(n9105));
  OAI21X1 g07409(.A0(n9093), .A1(n9089), .B0(n9105), .Y(n9106));
  AOI22X1 g07410(.A0(n7557), .A1(n9013), .B0(n7509), .B1(n6341), .Y(n9107));
  OAI21X1 g07411(.A0(n9019), .A1(n7592), .B0(n9107), .Y(n9108));
  AOI21X1 g07412(.A0(n9027), .A1(n7557), .B0(n6341), .Y(n9109));
  OAI21X1 g07413(.A0(n9028), .A1(n7558), .B0(n9109), .Y(n9110));
  AOI21X1 g07414(.A0(n9013), .A1(n7565), .B0(n9110), .Y(n9111));
  NAND2X1 g07415(.A(n9111), .B(n9108), .Y(n9112));
  AOI22X1 g07416(.A0(n7509), .A1(n9013), .B0(n7486), .B1(n6341), .Y(n9113));
  OAI21X1 g07417(.A0(n9019), .A1(n7517), .B0(n9113), .Y(n9114));
  AOI21X1 g07418(.A0(n9007), .A1(n7509), .B0(n6341), .Y(n9115));
  OAI21X1 g07419(.A0(n9005), .A1(n7510), .B0(n9115), .Y(n9116));
  AOI21X1 g07420(.A0(n9013), .A1(n7527), .B0(n9116), .Y(n9117));
  NAND2X1 g07421(.A(n9117), .B(n9114), .Y(n9118));
  NAND2X1 g07422(.A(n9118), .B(n9112), .Y(n9119));
  NOR2X1  g07423(.A(n9119), .B(n9106), .Y(n9120));
  NAND2X1 g07424(.A(n9120), .B(n9086), .Y(n9121));
  AOI22X1 g07425(.A0(n7304), .A1(n9013), .B0(n7255), .B1(n6341), .Y(n9122));
  OAI21X1 g07426(.A0(n9019), .A1(n7320), .B0(n9122), .Y(n9123));
  INVX1   g07427(.A(n9123), .Y(n9124));
  NOR2X1  g07428(.A(n9017), .B(n7320), .Y(n9125));
  AOI21X1 g07429(.A0(n9007), .A1(n7304), .B0(n6341), .Y(n9126));
  OAI21X1 g07430(.A0(n9005), .A1(n7305), .B0(n9126), .Y(n9127));
  NOR3X1  g07431(.A(n9127), .B(n9125), .C(n9124), .Y(n9128));
  AOI22X1 g07432(.A0(n7486), .A1(n9013), .B0(n7432), .B1(n6341), .Y(n9129));
  OAI21X1 g07433(.A0(n9019), .A1(n7502), .B0(n9129), .Y(n9130));
  AOI21X1 g07434(.A0(n9007), .A1(n7486), .B0(n6341), .Y(n9131));
  OAI21X1 g07435(.A0(n9005), .A1(n7464), .B0(n9131), .Y(n9132));
  AOI21X1 g07436(.A0(n9013), .A1(n7470), .B0(n9132), .Y(n9133));
  NAND2X1 g07437(.A(n9133), .B(n9130), .Y(n9134));
  AOI22X1 g07438(.A0(n7368), .A1(n9013), .B0(n7304), .B1(n6341), .Y(n9135));
  OAI21X1 g07439(.A0(n9019), .A1(n7374), .B0(n9135), .Y(n9136));
  AOI21X1 g07440(.A0(n9007), .A1(n7368), .B0(n6341), .Y(n9137));
  OAI21X1 g07441(.A0(n9005), .A1(n7360), .B0(n9137), .Y(n9138));
  AOI21X1 g07442(.A0(n9013), .A1(n7373), .B0(n9138), .Y(n9139));
  AOI22X1 g07443(.A0(n7432), .A1(n9013), .B0(n7368), .B1(n6341), .Y(n9140));
  OAI21X1 g07444(.A0(n9019), .A1(n7454), .B0(n9140), .Y(n9141));
  AOI21X1 g07445(.A0(n9007), .A1(n7432), .B0(n6341), .Y(n9142));
  OAI21X1 g07446(.A0(n9005), .A1(n7414), .B0(n9142), .Y(n9143));
  AOI21X1 g07447(.A0(n9013), .A1(n7425), .B0(n9143), .Y(n9144));
  AOI22X1 g07448(.A0(n9141), .A1(n9144), .B0(n9139), .B1(n9136), .Y(n9145));
  NAND2X1 g07449(.A(n9145), .B(n9134), .Y(n9146));
  NOR4X1  g07450(.A(n9128), .B(n9121), .C(n9085), .D(n9146), .Y(n9147));
  NAND4X1 g07451(.A(n9083), .B(n9082), .C(n9079), .D(n9147), .Y(n9148));
  AOI22X1 g07452(.A0(n7255), .A1(n9013), .B0(n7206), .B1(n6341), .Y(n9149));
  OAI21X1 g07453(.A0(n9019), .A1(n7265), .B0(n9149), .Y(n9150));
  INVX1   g07454(.A(n9150), .Y(n9151));
  AOI21X1 g07455(.A0(n9007), .A1(n7255), .B0(n6341), .Y(n9152));
  OAI21X1 g07456(.A0(n9005), .A1(n7312), .B0(n9152), .Y(n9153));
  AOI21X1 g07457(.A0(n9013), .A1(n7313), .B0(n9153), .Y(n9154));
  INVX1   g07458(.A(n9154), .Y(n9155));
  NOR2X1  g07459(.A(n9155), .B(n9151), .Y(n9156));
  AOI22X1 g07460(.A0(n7206), .A1(n9013), .B0(n7154), .B1(n6341), .Y(n9157));
  OAI21X1 g07461(.A0(n9019), .A1(n7218), .B0(n9157), .Y(n9158));
  AOI21X1 g07462(.A0(n9007), .A1(n7206), .B0(n6341), .Y(n9159));
  OAI21X1 g07463(.A0(n9005), .A1(n7207), .B0(n9159), .Y(n9160));
  AOI21X1 g07464(.A0(n9013), .A1(n7249), .B0(n9160), .Y(n9161));
  AOI22X1 g07465(.A0(n7103), .A1(n9013), .B0(n7072), .B1(n6341), .Y(n9162));
  OAI21X1 g07466(.A0(n9019), .A1(n7147), .B0(n9162), .Y(n9163));
  AOI21X1 g07467(.A0(n9007), .A1(n7103), .B0(n6341), .Y(n9164));
  OAI21X1 g07468(.A0(n9005), .A1(n7104), .B0(n9164), .Y(n9165));
  AOI21X1 g07469(.A0(n9013), .A1(n7115), .B0(n9165), .Y(n9166));
  AOI22X1 g07470(.A0(n9163), .A1(n9166), .B0(n9161), .B1(n9158), .Y(n9167));
  AOI22X1 g07471(.A0(n7154), .A1(n9013), .B0(n7103), .B1(n6341), .Y(n9168));
  OAI21X1 g07472(.A0(n9019), .A1(n7167), .B0(n9168), .Y(n9169));
  AOI21X1 g07473(.A0(n9007), .A1(n7154), .B0(n6341), .Y(n9170));
  OAI21X1 g07474(.A0(n9005), .A1(n7165), .B0(n9170), .Y(n9171));
  AOI21X1 g07475(.A0(n9013), .A1(n7164), .B0(n9171), .Y(n9172));
  NAND2X1 g07476(.A(n9172), .B(n9169), .Y(n9173));
  AOI22X1 g07477(.A0(n6944), .A1(n9013), .B0(n6894), .B1(n6341), .Y(n9174));
  OAI21X1 g07478(.A0(n9019), .A1(n6984), .B0(n9174), .Y(n9175));
  AOI21X1 g07479(.A0(n9007), .A1(n6944), .B0(n6341), .Y(n9176));
  OAI21X1 g07480(.A0(n9005), .A1(n6945), .B0(n9176), .Y(n9177));
  AOI21X1 g07481(.A0(n9013), .A1(n6956), .B0(n9177), .Y(n9178));
  AOI22X1 g07482(.A0(n6992), .A1(n9013), .B0(n6944), .B1(n6341), .Y(n9179));
  OAI21X1 g07483(.A0(n9019), .A1(n7006), .B0(n9179), .Y(n9180));
  INVX1   g07484(.A(n9180), .Y(n9181));
  NOR2X1  g07485(.A(n9017), .B(n7006), .Y(n9182));
  AOI21X1 g07486(.A0(n9007), .A1(n6992), .B0(n6341), .Y(n9183));
  OAI21X1 g07487(.A0(n9005), .A1(n6993), .B0(n9183), .Y(n9184));
  NOR3X1  g07488(.A(n9184), .B(n9182), .C(n9181), .Y(n9185));
  AOI21X1 g07489(.A0(n9178), .A1(n9175), .B0(n9185), .Y(n9186));
  AOI22X1 g07490(.A0(n6894), .A1(n9013), .B0(n6839), .B1(n6341), .Y(n9187));
  OAI21X1 g07491(.A0(n9019), .A1(n6935), .B0(n9187), .Y(n9188));
  AOI21X1 g07492(.A0(n9007), .A1(n6894), .B0(n6341), .Y(n9189));
  OAI21X1 g07493(.A0(n9005), .A1(n6895), .B0(n9189), .Y(n9190));
  AOI21X1 g07494(.A0(n9013), .A1(n6909), .B0(n9190), .Y(n9191));
  AOI22X1 g07495(.A0(n7072), .A1(n9013), .B0(n6992), .B1(n6341), .Y(n9192));
  OAI21X1 g07496(.A0(n9019), .A1(n7073), .B0(n9192), .Y(n9193));
  AOI21X1 g07497(.A0(n9007), .A1(n7072), .B0(n6341), .Y(n9194));
  OAI21X1 g07498(.A0(n9005), .A1(n7051), .B0(n9194), .Y(n9195));
  AOI21X1 g07499(.A0(n9013), .A1(n7063), .B0(n9195), .Y(n9196));
  AOI22X1 g07500(.A0(n9193), .A1(n9196), .B0(n9191), .B1(n9188), .Y(n9197));
  NAND4X1 g07501(.A(n9186), .B(n9173), .C(n9167), .D(n9197), .Y(n9198));
  NOR2X1  g07502(.A(n9198), .B(n9156), .Y(n9199));
  AOI22X1 g07503(.A0(n6839), .A1(n9013), .B0(n6807), .B1(n6341), .Y(n9200));
  OAI21X1 g07504(.A0(n9019), .A1(n6886), .B0(n9200), .Y(n9201));
  AOI21X1 g07505(.A0(n9007), .A1(n6839), .B0(n6341), .Y(n9202));
  OAI21X1 g07506(.A0(n9005), .A1(n6840), .B0(n9202), .Y(n9203));
  AOI21X1 g07507(.A0(n9013), .A1(n6851), .B0(n9203), .Y(n9204));
  AOI22X1 g07508(.A0(n6807), .A1(n9013), .B0(n6745), .B1(n6341), .Y(n9205));
  OAI21X1 g07509(.A0(n9019), .A1(n6832), .B0(n9205), .Y(n9206));
  AOI21X1 g07510(.A0(n9007), .A1(n6807), .B0(n6341), .Y(n9207));
  OAI21X1 g07511(.A0(n9005), .A1(n6786), .B0(n9207), .Y(n9208));
  AOI21X1 g07512(.A0(n9013), .A1(n6797), .B0(n9208), .Y(n9209));
  AOI22X1 g07513(.A0(n9206), .A1(n9209), .B0(n9204), .B1(n9201), .Y(n9210));
  INVX1   g07514(.A(n9210), .Y(n9211));
  AOI22X1 g07515(.A0(n6745), .A1(n9013), .B0(n6706), .B1(n6341), .Y(n9212));
  OAI21X1 g07516(.A0(n9019), .A1(n6753), .B0(n9212), .Y(n9213));
  INVX1   g07517(.A(n9213), .Y(n9214));
  AOI21X1 g07518(.A0(n9007), .A1(n6745), .B0(n6341), .Y(n9215));
  OAI21X1 g07519(.A0(n9005), .A1(n6732), .B0(n9215), .Y(n9216));
  AOI21X1 g07520(.A0(n9013), .A1(n6752), .B0(n9216), .Y(n9217));
  INVX1   g07521(.A(n9217), .Y(n9218));
  AOI21X1 g07522(.A0(n9007), .A1(n6706), .B0(n6341), .Y(n9219));
  OAI21X1 g07523(.A0(n9017), .A1(n6723), .B0(n9219), .Y(n9220));
  AOI21X1 g07524(.A0(n9027), .A1(n6706), .B0(n9220), .Y(n9221));
  INVX1   g07525(.A(n9221), .Y(n9222));
  AOI22X1 g07526(.A0(n6706), .A1(n9013), .B0(n6652), .B1(n6341), .Y(n9223));
  OAI21X1 g07527(.A0(n9019), .A1(n6723), .B0(n9223), .Y(n9224));
  INVX1   g07528(.A(n9224), .Y(n9225));
  OAI22X1 g07529(.A0(n9222), .A1(n9225), .B0(n9218), .B1(n9214), .Y(n9226));
  NOR2X1  g07530(.A(n9226), .B(n9211), .Y(n9227));
  AOI22X1 g07531(.A0(n6652), .A1(n9013), .B0(n6583), .B1(n6341), .Y(n9228));
  OAI21X1 g07532(.A0(n9019), .A1(n6677), .B0(n9228), .Y(n9229));
  AOI21X1 g07533(.A0(n9007), .A1(n6652), .B0(n6341), .Y(n9230));
  OAI21X1 g07534(.A0(n9017), .A1(n6677), .B0(n9230), .Y(n9231));
  AOI21X1 g07535(.A0(n9027), .A1(n6652), .B0(n9231), .Y(n9232));
  AOI21X1 g07536(.A0(n9013), .A1(n6600), .B0(n6341), .Y(n9233));
  OAI21X1 g07537(.A0(n9028), .A1(n6595), .B0(n9233), .Y(n9234));
  AOI21X1 g07538(.A0(n9027), .A1(n6583), .B0(n9234), .Y(n9235));
  AOI22X1 g07539(.A0(n6583), .A1(n9013), .B0(n6569), .B1(n6341), .Y(n9236));
  OAI21X1 g07540(.A0(n9019), .A1(n6601), .B0(n9236), .Y(n9237));
  AOI22X1 g07541(.A0(n9235), .A1(n9237), .B0(n9232), .B1(n9229), .Y(n9238));
  INVX1   g07542(.A(n9238), .Y(n9239));
  AOI22X1 g07543(.A0(n6569), .A1(n9013), .B0(n6573), .B1(n6341), .Y(n9240));
  OAI21X1 g07544(.A0(n9019), .A1(n6554), .B0(n9240), .Y(n9241));
  AOI21X1 g07545(.A0(n9013), .A1(n6580), .B0(n6341), .Y(n9242));
  OAI21X1 g07546(.A0(n9028), .A1(n6542), .B0(n9242), .Y(n9243));
  AOI21X1 g07547(.A0(n9027), .A1(n6569), .B0(n9243), .Y(n9244));
  NOR3X1  g07548(.A(n9244), .B(n9241), .C(n9239), .Y(n9245));
  NAND4X1 g07549(.A(n9227), .B(n9199), .C(n9047), .D(n9245), .Y(n9246));
  NOR4X1  g07550(.A(n9148), .B(n9041), .C(n9035), .D(n9246), .Y(n9247));
  OAI21X1 g07551(.A0(n9019), .A1(n7941), .B0(n9037), .Y(n9248));
  NAND3X1 g07552(.A(n9013), .B(n6750), .C(n6314), .Y(n9249));
  NAND3X1 g07553(.A(n9039), .B(n9249), .C(n9248), .Y(n9250));
  INVX1   g07554(.A(n9158), .Y(n9251));
  NOR2X1  g07555(.A(n9017), .B(n7218), .Y(n9252));
  NOR3X1  g07556(.A(n9160), .B(n9252), .C(n9251), .Y(n9253));
  NOR3X1  g07557(.A(n9166), .B(n9163), .C(n9253), .Y(n9254));
  AOI22X1 g07558(.A0(n9169), .A1(n9172), .B0(n9154), .B1(n9150), .Y(n9255));
  NAND4X1 g07559(.A(n9254), .B(n9047), .C(n9250), .D(n9255), .Y(n9256));
  NOR3X1  g07560(.A(n9256), .B(n9148), .C(n9035), .Y(n9257));
  INVX1   g07561(.A(n9193), .Y(n9258));
  INVX1   g07562(.A(n9196), .Y(n9259));
  NAND2X1 g07563(.A(n9255), .B(n9167), .Y(n9260));
  INVX1   g07564(.A(n9260), .Y(n9261));
  NAND4X1 g07565(.A(n9259), .B(n9258), .C(n9047), .D(n9261), .Y(n9262));
  NOR4X1  g07566(.A(n9148), .B(n9041), .C(n9035), .D(n9262), .Y(n9263));
  NOR4X1  g07567(.A(n9257), .B(n9247), .C(n9076), .D(n9263), .Y(n9264));
  AOI21X1 g07568(.A0(n9039), .A1(n9249), .B0(n9248), .Y(n9265));
  NOR2X1  g07569(.A(n9063), .B(n9059), .Y(n9266));
  OAI21X1 g07570(.A0(n9054), .A1(n9057), .B0(n9266), .Y(n9267));
  AOI21X1 g07571(.A0(n9046), .A1(n9043), .B0(n9267), .Y(n9268));
  AOI21X1 g07572(.A0(n9268), .A1(n9250), .B0(n9265), .Y(n9269));
  NOR3X1  g07573(.A(n9269), .B(n9035), .C(n9024), .Y(n9270));
  NAND4X1 g07574(.A(n9151), .B(n9047), .C(n9250), .D(n9155), .Y(n9271));
  NOR3X1  g07575(.A(n9271), .B(n9148), .C(n9035), .Y(n9272));
  OAI22X1 g07576(.A0(n9017), .A1(n6505), .B0(n6531), .B1(n9019), .Y(n9273));
  AOI21X1 g07577(.A0(n9013), .A1(n6483), .B0(n6341), .Y(n9274));
  OAI21X1 g07578(.A0(n9028), .A1(n6505), .B0(n9274), .Y(n9275));
  AOI21X1 g07579(.A0(n9027), .A1(n6573), .B0(n9275), .Y(n9276));
  NOR2X1  g07580(.A(n6460), .B(n6458), .Y(n9277));
  NOR4X1  g07581(.A(n6455), .B(n6452), .C(n6341), .D(n9277), .Y(n9278));
  OAI21X1 g07582(.A0(n9278), .A1(n9276), .B0(n9273), .Y(n9279));
  AOI22X1 g07583(.A0(n9276), .A1(n9278), .B0(n9244), .B1(n9241), .Y(n9280));
  NAND4X1 g07584(.A(n9279), .B(n9238), .C(n9227), .D(n9280), .Y(n9281));
  NOR3X1  g07585(.A(n9281), .B(n9198), .C(n9156), .Y(n9282));
  NAND3X1 g07586(.A(n9282), .B(n9047), .C(n9250), .Y(n9283));
  NOR3X1  g07587(.A(n9283), .B(n9148), .C(n9035), .Y(n9284));
  NOR4X1  g07588(.A(n9229), .B(n9226), .C(n9211), .D(n9232), .Y(n9285));
  NAND4X1 g07589(.A(n9199), .B(n9047), .C(n9250), .D(n9285), .Y(n9286));
  NOR3X1  g07590(.A(n9286), .B(n9148), .C(n9035), .Y(n9287));
  NOR4X1  g07591(.A(n9284), .B(n9272), .C(n9270), .D(n9287), .Y(n9288));
  AOI21X1 g07592(.A0(n9055), .A1(n9050), .B0(n9085), .Y(n9289));
  INVX1   g07593(.A(n9086), .Y(n9290));
  NOR4X1  g07594(.A(n9108), .B(n9106), .C(n9290), .D(n9111), .Y(n9291));
  NAND4X1 g07595(.A(n9289), .B(n9047), .C(n9250), .D(n9291), .Y(n9292));
  NOR3X1  g07596(.A(n9292), .B(n9035), .C(n9024), .Y(n9293));
  NOR2X1  g07597(.A(n9093), .B(n9089), .Y(n9294));
  NOR4X1  g07598(.A(n9101), .B(n9294), .C(n9290), .D(n9104), .Y(n9295));
  NAND4X1 g07599(.A(n9289), .B(n9047), .C(n9250), .D(n9295), .Y(n9296));
  NOR3X1  g07600(.A(n9296), .B(n9035), .C(n9024), .Y(n9297));
  INVX1   g07601(.A(n9134), .Y(n9298));
  NAND2X1 g07602(.A(n9144), .B(n9141), .Y(n9299));
  NOR2X1  g07603(.A(n9139), .B(n9136), .Y(n9300));
  NAND2X1 g07604(.A(n9300), .B(n9299), .Y(n9301));
  NOR4X1  g07605(.A(n9298), .B(n9121), .C(n9065), .D(n9301), .Y(n9302));
  NAND3X1 g07606(.A(n9302), .B(n9047), .C(n9250), .Y(n9303));
  NOR3X1  g07607(.A(n9303), .B(n9035), .C(n9024), .Y(n9304));
  NOR4X1  g07608(.A(n9141), .B(n9298), .C(n9065), .D(n9144), .Y(n9305));
  NAND3X1 g07609(.A(n9305), .B(n9047), .C(n9250), .Y(n9306));
  NOR4X1  g07610(.A(n9121), .B(n9035), .C(n9024), .D(n9306), .Y(n9307));
  NOR4X1  g07611(.A(n9304), .B(n9297), .C(n9293), .D(n9307), .Y(n9308));
  NAND3X1 g07612(.A(n9308), .B(n9288), .C(n9264), .Y(n9309));
  NOR3X1  g07613(.A(n9161), .B(n9158), .C(n9156), .Y(n9310));
  NAND3X1 g07614(.A(n9310), .B(n9047), .C(n9250), .Y(n9311));
  NOR3X1  g07615(.A(n9311), .B(n9148), .C(n9035), .Y(n9312));
  NOR2X1  g07616(.A(n9259), .B(n9258), .Y(n9313));
  NOR3X1  g07617(.A(n9313), .B(n9191), .C(n9188), .Y(n9314));
  NAND4X1 g07618(.A(n9261), .B(n9186), .C(n9047), .D(n9314), .Y(n9315));
  NOR4X1  g07619(.A(n9148), .B(n9041), .C(n9035), .D(n9315), .Y(n9316));
  INVX1   g07620(.A(n9201), .Y(n9317));
  INVX1   g07621(.A(n9204), .Y(n9318));
  NOR2X1  g07622(.A(n9318), .B(n9317), .Y(n9319));
  NOR3X1  g07623(.A(n9209), .B(n9206), .C(n9319), .Y(n9320));
  NAND4X1 g07624(.A(n9199), .B(n9047), .C(n9250), .D(n9320), .Y(n9321));
  NOR3X1  g07625(.A(n9321), .B(n9148), .C(n9035), .Y(n9322));
  NAND2X1 g07626(.A(n9232), .B(n9229), .Y(n9323));
  INVX1   g07627(.A(n9323), .Y(n9324));
  NOR3X1  g07628(.A(n9237), .B(n9235), .C(n9324), .Y(n9325));
  NAND4X1 g07629(.A(n9227), .B(n9199), .C(n9047), .D(n9325), .Y(n9326));
  NOR4X1  g07630(.A(n9148), .B(n9041), .C(n9035), .D(n9326), .Y(n9327));
  NOR4X1  g07631(.A(n9322), .B(n9316), .C(n9312), .D(n9327), .Y(n9328));
  OAI21X1 g07632(.A0(n9184), .A1(n9182), .B0(n9181), .Y(n9329));
  NOR3X1  g07633(.A(n9329), .B(n9260), .C(n9313), .Y(n9330));
  NAND3X1 g07634(.A(n9330), .B(n9047), .C(n9250), .Y(n9331));
  NOR3X1  g07635(.A(n9331), .B(n9148), .C(n9035), .Y(n9332));
  NAND3X1 g07636(.A(n9034), .B(n9032), .C(n9031), .Y(n9333));
  INVX1   g07637(.A(n8996), .Y(n9334));
  NOR2X1  g07638(.A(n9334), .B(n6342), .Y(n9335));
  NOR3X1  g07639(.A(n9335), .B(n9022), .C(n9018), .Y(n9336));
  OAI21X1 g07640(.A0(n9081), .A1(n9080), .B0(n9335), .Y(n9337));
  OAI21X1 g07641(.A0(n9023), .A1(n9016), .B0(n9337), .Y(n9338));
  OAI22X1 g07642(.A0(n9336), .A1(n9338), .B0(n9333), .B1(n9024), .Y(n9339));
  NOR2X1  g07643(.A(n9224), .B(n9221), .Y(n9340));
  OAI21X1 g07644(.A0(n9218), .A1(n9214), .B0(n9340), .Y(n9341));
  NOR4X1  g07645(.A(n9211), .B(n9198), .C(n9156), .D(n9341), .Y(n9342));
  NAND3X1 g07646(.A(n9342), .B(n9047), .C(n9250), .Y(n9343));
  NOR3X1  g07647(.A(n9343), .B(n9148), .C(n9035), .Y(n9344));
  OAI21X1 g07648(.A0(n9127), .A1(n9125), .B0(n9124), .Y(n9345));
  NOR4X1  g07649(.A(n9146), .B(n9121), .C(n9065), .D(n9345), .Y(n9346));
  NAND3X1 g07650(.A(n9346), .B(n9047), .C(n9250), .Y(n9347));
  NOR3X1  g07651(.A(n9347), .B(n9035), .C(n9024), .Y(n9348));
  NOR4X1  g07652(.A(n9344), .B(n9339), .C(n9332), .D(n9348), .Y(n9349));
  NAND4X1 g07653(.A(n9317), .B(n9199), .C(n9047), .D(n9318), .Y(n9350));
  NOR4X1  g07654(.A(n9148), .B(n9041), .C(n9035), .D(n9350), .Y(n9351));
  NAND2X1 g07655(.A(n9104), .B(n9101), .Y(n9352));
  NOR2X1  g07656(.A(n9098), .B(n9095), .Y(n9353));
  NAND2X1 g07657(.A(n9353), .B(n9352), .Y(n9354));
  NOR4X1  g07658(.A(n9294), .B(n9290), .C(n9065), .D(n9354), .Y(n9355));
  NAND3X1 g07659(.A(n9355), .B(n9047), .C(n9250), .Y(n9356));
  NOR3X1  g07660(.A(n9356), .B(n9035), .C(n9024), .Y(n9357));
  INVX1   g07661(.A(n9089), .Y(n9358));
  INVX1   g07662(.A(n9093), .Y(n9359));
  NOR4X1  g07663(.A(n9358), .B(n9290), .C(n9065), .D(n9359), .Y(n9360));
  NAND3X1 g07664(.A(n9360), .B(n9047), .C(n9250), .Y(n9361));
  NOR3X1  g07665(.A(n9361), .B(n9035), .C(n9024), .Y(n9362));
  NOR4X1  g07666(.A(n9185), .B(n9178), .C(n9175), .D(n9313), .Y(n9363));
  NAND4X1 g07667(.A(n9261), .B(n9047), .C(n9250), .D(n9363), .Y(n9364));
  NOR3X1  g07668(.A(n9364), .B(n9148), .C(n9035), .Y(n9365));
  NOR4X1  g07669(.A(n9362), .B(n9357), .C(n9351), .D(n9365), .Y(n9366));
  NOR3X1  g07670(.A(n9133), .B(n9130), .C(n9065), .Y(n9367));
  NAND3X1 g07671(.A(n9367), .B(n9047), .C(n9250), .Y(n9368));
  NOR4X1  g07672(.A(n9121), .B(n9035), .C(n9024), .D(n9368), .Y(n9369));
  NAND2X1 g07673(.A(n9209), .B(n9206), .Y(n9370));
  NOR3X1  g07674(.A(n9217), .B(n9213), .C(n9319), .Y(n9371));
  NAND4X1 g07675(.A(n9370), .B(n9199), .C(n9047), .D(n9371), .Y(n9372));
  NOR4X1  g07676(.A(n9148), .B(n9041), .C(n9035), .D(n9372), .Y(n9373));
  INVX1   g07677(.A(n9112), .Y(n9374));
  NOR4X1  g07678(.A(n9114), .B(n9374), .C(n9106), .D(n9117), .Y(n9375));
  NAND4X1 g07679(.A(n9086), .B(n9289), .C(n9047), .D(n9375), .Y(n9376));
  NOR4X1  g07680(.A(n9041), .B(n9035), .C(n9024), .D(n9376), .Y(n9377));
  NOR4X1  g07681(.A(n9169), .B(n9253), .C(n9156), .D(n9172), .Y(n9378));
  NAND3X1 g07682(.A(n9378), .B(n9047), .C(n9250), .Y(n9379));
  NOR3X1  g07683(.A(n9379), .B(n9148), .C(n9035), .Y(n9380));
  NOR4X1  g07684(.A(n9377), .B(n9373), .C(n9369), .D(n9380), .Y(n9381));
  NAND4X1 g07685(.A(n9366), .B(n9349), .C(n9328), .D(n9381), .Y(n9382));
  NAND3X1 g07686(.A(n6513), .B(n6455), .C(n6451), .Y(n9383));
  NAND3X1 g07687(.A(n9383), .B(n6670), .C(n6669), .Y(n9384));
  OAI21X1 g07688(.A0(n9382), .A1(n9309), .B0(n9384), .Y(n9385));
  NOR2X1  g07689(.A(n9382), .B(n9309), .Y(n9386));
  AOI21X1 g07690(.A0(n6451), .A1(n6449), .B0(n6460), .Y(n9387));
  OAI21X1 g07691(.A0(n9387), .A1(n6455), .B0(n6517), .Y(n9388));
  NAND3X1 g07692(.A(n6513), .B(n6455), .C(n6452), .Y(n9389));
  XOR2X1  g07693(.A(n7984), .B(n7954), .Y(n9390));
  XOR2X1  g07694(.A(n7998), .B(n8993), .Y(n9391));
  XOR2X1  g07695(.A(n7787), .B(n7780), .Y(n9395));
  XOR2X1  g07696(.A(n7608), .B(n7600), .Y(n9396));
  XOR2X1  g07697(.A(n7565), .B(n7557), .Y(n9397));
  XOR2X1  g07698(.A(n7517), .B(n7510), .Y(n9398));
  OAI21X1 g07699(.A0(n7173), .A1(n7176), .B0(n7177), .Y(n9401));
  XOR2X1  g07700(.A(n6505), .B(n6531), .Y(n9403));
  NOR4X1  g07701(.A(n6653), .B(n6602), .C(n6555), .D(n9403), .Y(n9404));
  NAND3X1 g07702(.A(n9404), .B(n6859), .C(n6704), .Y(n9405));
  XOR2X1  g07703(.A(n6752), .B(n6745), .Y(n9406));
  NOR3X1  g07704(.A(n9406), .B(n9405), .C(n6808), .Y(n9407));
  XOR2X1  g07705(.A(n7004), .B(n6992), .Y(n9408));
  NOR3X1  g07706(.A(n9408), .B(n7084), .C(n6972), .Y(n9409));
  NAND3X1 g07707(.A(n9409), .B(n9407), .C(n6910), .Y(n9410));
  OAI22X1 g07708(.A0(n7333), .A1(n7335), .B0(n7280), .B1(n7279), .Y(n9411));
  NOR4X1  g07709(.A(n9410), .B(n9401), .C(n7338), .D(n9411), .Y(n9412));
  NAND4X1 g07710(.A(n7379), .B(n7471), .C(n7426), .D(n9412), .Y(n9413));
  NOR4X1  g07711(.A(n9398), .B(n9397), .C(n9396), .D(n9413), .Y(n9414));
  OAI21X1 g07712(.A0(n7709), .A1(n7706), .B0(n9414), .Y(n9415));
  NOR4X1  g07713(.A(n9395), .B(n7759), .C(n7724), .D(n9415), .Y(n9416));
  NAND4X1 g07714(.A(n7849), .B(n7894), .C(n7942), .D(n9416), .Y(n9417));
  NOR3X1  g07715(.A(n9417), .B(n9391), .C(n9390), .Y(n9418));
  INVX1   g07716(.A(P2_B_REG_SCAN_IN), .Y(n9419));
  AOI21X1 g07717(.A0(n8996), .A1(n8409), .B0(n6342), .Y(n9420));
  NOR2X1  g07718(.A(n6449), .B(n6341), .Y(n9421));
  NOR4X1  g07719(.A(n9420), .B(n8492), .C(P2_U3088), .D(n9421), .Y(n9422));
  NOR2X1  g07720(.A(n9422), .B(n9419), .Y(n9423));
  NOR3X1  g07721(.A(n6513), .B(n6456), .C(n6451), .Y(n9424));
  AOI21X1 g07722(.A0(n9424), .A1(n9418), .B0(n9423), .Y(n9425));
  OAI21X1 g07723(.A0(n9418), .A1(n9389), .B0(n9425), .Y(n9426));
  AOI21X1 g07724(.A0(n9388), .A1(n9386), .B0(n9426), .Y(n9427));
  NAND3X1 g07725(.A(n8996), .B(n8409), .C(n6350), .Y(n9428));
  NAND2X1 g07726(.A(n9428), .B(n6341), .Y(n9429));
  AOI21X1 g07727(.A0(n9429), .A1(P2_STATE_REG_SCAN_IN), .B0(n9423), .Y(n9430));
  AOI21X1 g07728(.A0(n9427), .A1(n9385), .B0(n9430), .Y(P2_U3328));
  NAND4X1 g07729(.A(n6455), .B(n6451), .C(n6449), .D(n6460), .Y(n9432));
  AOI21X1 g07730(.A0(n6943), .A1(n6937), .B0(n8087), .Y(n9434));
  INVX1   g07731(.A(n9434), .Y(n9435));
  NOR2X1  g07732(.A(n8087), .B(n6685), .Y(n9436));
  OAI21X1 g07733(.A0(n6513), .A1(n6449), .B0(n6455), .Y(n9437));
  OAI21X1 g07734(.A0(n6455), .A1(n6451), .B0(n9437), .Y(n9438));
  XOR2X1  g07735(.A(n9438), .B(n6600), .Y(n9439));
  AOI21X1 g07736(.A0(n9432), .A1(n6583), .B0(n9439), .Y(n9440));
  AOI21X1 g07737(.A0(n6651), .A1(n6649), .B0(n8087), .Y(n9441));
  INVX1   g07738(.A(n9441), .Y(n9442));
  INVX1   g07739(.A(n9438), .Y(n9443));
  XOR2X1  g07740(.A(n9443), .B(n6646), .Y(n9444));
  AOI21X1 g07741(.A0(n9444), .A1(n9442), .B0(n9440), .Y(n9445));
  XOR2X1  g07742(.A(n9438), .B(n6554), .Y(n9446));
  OAI21X1 g07743(.A0(n8087), .A1(n6542), .B0(n9446), .Y(n9447));
  NAND3X1 g07744(.A(n9447), .B(n9438), .C(n6531), .Y(n9448));
  OAI21X1 g07745(.A0(n6504), .A1(n6494), .B0(n9432), .Y(n9449));
  AOI21X1 g07746(.A0(n9443), .A1(n6531), .B0(n9449), .Y(n9450));
  NAND2X1 g07747(.A(n9450), .B(n9447), .Y(n9451));
  INVX1   g07748(.A(n9446), .Y(n9452));
  AOI21X1 g07749(.A0(n6568), .A1(n6567), .B0(n8087), .Y(n9453));
  NAND2X1 g07750(.A(n9453), .B(n9452), .Y(n9454));
  NAND3X1 g07751(.A(n9454), .B(n9451), .C(n9448), .Y(n9455));
  NAND2X1 g07752(.A(n9455), .B(n9445), .Y(n9456));
  NAND3X1 g07753(.A(n9439), .B(n9432), .C(n6583), .Y(n9457));
  INVX1   g07754(.A(n9457), .Y(n9458));
  AOI21X1 g07755(.A0(n9457), .A1(n9442), .B0(n9444), .Y(n9459));
  AOI21X1 g07756(.A0(n9458), .A1(n9441), .B0(n9459), .Y(n9460));
  NAND2X1 g07757(.A(n9460), .B(n9456), .Y(n9461));
  NAND2X1 g07758(.A(n9461), .B(n9436), .Y(n9462));
  XOR2X1  g07759(.A(n9443), .B(n6703), .Y(n9463));
  INVX1   g07760(.A(n9463), .Y(n9464));
  OAI21X1 g07761(.A0(n9461), .A1(n9436), .B0(n9464), .Y(n9465));
  NAND2X1 g07762(.A(n9465), .B(n9462), .Y(n9466));
  XOR2X1  g07763(.A(n9443), .B(n6909), .Y(n9467));
  INVX1   g07764(.A(n9467), .Y(n9468));
  AOI21X1 g07765(.A0(n6893), .A1(n6887), .B0(n8087), .Y(n9469));
  NOR2X1  g07766(.A(n9469), .B(n9468), .Y(n9470));
  NOR2X1  g07767(.A(n8087), .B(n6786), .Y(n9471));
  XOR2X1  g07768(.A(n9443), .B(n6797), .Y(n9472));
  INVX1   g07769(.A(n9472), .Y(n9473));
  AOI21X1 g07770(.A0(n6838), .A1(n6834), .B0(n8087), .Y(n9474));
  XOR2X1  g07771(.A(n9443), .B(n6851), .Y(n9475));
  INVX1   g07772(.A(n9475), .Y(n9476));
  OAI22X1 g07773(.A0(n9474), .A1(n9476), .B0(n9473), .B1(n9471), .Y(n9477));
  AOI21X1 g07774(.A0(n6744), .A1(n6742), .B0(n8087), .Y(n9478));
  XOR2X1  g07775(.A(n9438), .B(n6752), .Y(n9479));
  NOR2X1  g07776(.A(n9479), .B(n9478), .Y(n9480));
  NOR3X1  g07777(.A(n9480), .B(n9477), .C(n9470), .Y(n9481));
  NOR3X1  g07778(.A(n9472), .B(n8087), .C(n6786), .Y(n9482));
  NOR2X1  g07779(.A(n9482), .B(n9474), .Y(n9483));
  NOR2X1  g07780(.A(n9483), .B(n9475), .Y(n9484));
  NAND2X1 g07781(.A(n9479), .B(n9478), .Y(n9485));
  NAND2X1 g07782(.A(n9482), .B(n9474), .Y(n9486));
  OAI21X1 g07783(.A0(n9485), .A1(n9477), .B0(n9486), .Y(n9487));
  OAI22X1 g07784(.A0(n9484), .A1(n9487), .B0(n9469), .B1(n9468), .Y(n9488));
  NAND2X1 g07785(.A(n9469), .B(n9468), .Y(n9489));
  NAND2X1 g07786(.A(n9489), .B(n9488), .Y(n9490));
  AOI21X1 g07787(.A0(n9481), .A1(n9466), .B0(n9490), .Y(n9491));
  NOR2X1  g07788(.A(n9491), .B(n9435), .Y(n9492));
  XOR2X1  g07789(.A(n9443), .B(n6956), .Y(n9493));
  AOI21X1 g07790(.A0(n9491), .A1(n9435), .B0(n9493), .Y(n9494));
  XOR2X1  g07791(.A(n9438), .B(n7218), .Y(n9495));
  INVX1   g07792(.A(n9495), .Y(n9496));
  AOI21X1 g07793(.A0(n7205), .A1(n7201), .B0(n8087), .Y(n9497));
  NOR2X1  g07794(.A(n9497), .B(n9496), .Y(n9498));
  XOR2X1  g07795(.A(n9443), .B(n7115), .Y(n9499));
  OAI21X1 g07796(.A0(n8087), .A1(n7104), .B0(n9499), .Y(n9500));
  XOR2X1  g07797(.A(n9443), .B(n7164), .Y(n9501));
  OAI21X1 g07798(.A0(n8087), .A1(n7165), .B0(n9501), .Y(n9502));
  XOR2X1  g07799(.A(n9438), .B(n7063), .Y(n9503));
  AOI21X1 g07800(.A0(n7049), .A1(n7043), .B0(n8087), .Y(n9504));
  NOR2X1  g07801(.A(n9504), .B(n9503), .Y(n9505));
  INVX1   g07802(.A(n9505), .Y(n9506));
  AOI21X1 g07803(.A0(n6991), .A1(n6986), .B0(n8087), .Y(n9507));
  XOR2X1  g07804(.A(n9443), .B(n7004), .Y(n9508));
  INVX1   g07805(.A(n9508), .Y(n9509));
  NOR2X1  g07806(.A(n9509), .B(n9507), .Y(n9510));
  INVX1   g07807(.A(n9510), .Y(n9511));
  NAND4X1 g07808(.A(n9506), .B(n9502), .C(n9500), .D(n9511), .Y(n9512));
  NOR2X1  g07809(.A(n9512), .B(n9498), .Y(n9513));
  OAI21X1 g07810(.A0(n9494), .A1(n9492), .B0(n9513), .Y(n9514));
  NAND2X1 g07811(.A(n9502), .B(n9500), .Y(n9515));
  INVX1   g07812(.A(n9507), .Y(n9516));
  NOR2X1  g07813(.A(n9508), .B(n9516), .Y(n9517));
  INVX1   g07814(.A(n9517), .Y(n9518));
  NOR3X1  g07815(.A(n9518), .B(n9505), .C(n9515), .Y(n9519));
  NAND2X1 g07816(.A(n9504), .B(n9503), .Y(n9520));
  INVX1   g07817(.A(n9501), .Y(n9521));
  AOI21X1 g07818(.A0(n7153), .A1(n7149), .B0(n8087), .Y(n9522));
  NOR3X1  g07819(.A(n9499), .B(n8087), .C(n7104), .Y(n9523));
  AOI21X1 g07820(.A0(n9522), .A1(n9521), .B0(n9523), .Y(n9524));
  OAI21X1 g07821(.A0(n9520), .A1(n9515), .B0(n9524), .Y(n9525));
  AOI21X1 g07822(.A0(n9525), .A1(n9502), .B0(n9519), .Y(n9526));
  NOR2X1  g07823(.A(n9526), .B(n9498), .Y(n9527));
  AOI21X1 g07824(.A0(n9497), .A1(n9496), .B0(n9527), .Y(n9528));
  NAND2X1 g07825(.A(n9528), .B(n9514), .Y(n9529));
  XOR2X1  g07826(.A(n9438), .B(n7265), .Y(n9530));
  AOI21X1 g07827(.A0(n7254), .A1(n7250), .B0(n8087), .Y(n9531));
  XOR2X1  g07828(.A(n9531), .B(n9530), .Y(n9532));
  XOR2X1  g07829(.A(n9532), .B(n9529), .Y(n9533));
  NOR3X1  g07830(.A(n6464), .B(n6446), .C(n8072), .Y(n9534));
  INVX1   g07831(.A(n9534), .Y(n9535));
  NOR2X1  g07832(.A(n9001), .B(n6455), .Y(n9536));
  NAND2X1 g07833(.A(n6455), .B(n6458), .Y(n9537));
  NAND4X1 g07834(.A(n9537), .B(n9432), .C(n6633), .D(n9017), .Y(n9538));
  NOR2X1  g07835(.A(n9538), .B(n9536), .Y(n9539));
  NOR3X1  g07836(.A(n9539), .B(n9535), .C(n6357), .Y(n9540));
  INVX1   g07837(.A(n9540), .Y(n9541));
  NOR4X1  g07838(.A(n6349), .B(n6342), .C(P2_U3088), .D(n8082), .Y(n9542));
  NOR3X1  g07839(.A(n8074), .B(n6349), .C(n6342), .Y(n9543));
  OAI21X1 g07840(.A0(n9539), .A1(n9534), .B0(n9543), .Y(n9544));
  AOI22X1 g07841(.A0(n9542), .A1(n9535), .B0(P2_STATE_REG_SCAN_IN), .B1(n9544), .Y(n9545));
  INVX1   g07842(.A(n9545), .Y(n9546));
  NOR4X1  g07843(.A(n6349), .B(n6342), .C(P2_U3088), .D(n9334), .Y(n9547));
  INVX1   g07844(.A(n9547), .Y(n9548));
  NOR4X1  g07845(.A(n6464), .B(n6446), .C(n8072), .D(n6473), .Y(n9549));
  NOR4X1  g07846(.A(n6464), .B(n6446), .C(n8072), .D(n6481), .Y(n9550));
  INVX1   g07847(.A(n9550), .Y(n9551));
  OAI22X1 g07848(.A0(n9534), .A1(n7252), .B0(n7207), .B1(n9551), .Y(n9552));
  AOI21X1 g07849(.A0(n9549), .A1(n7304), .B0(n9552), .Y(n9553));
  AOI22X1 g07850(.A0(n9534), .A1(n9542), .B0(n8071), .B1(n6350), .Y(n9554));
  AOI22X1 g07851(.A0(n7313), .A1(n9636), .B0(P2_U3088), .B1(P2_REG3_REG_15__SCAN_IN), .Y(n9556));
  OAI21X1 g07852(.A0(n9553), .A1(n9548), .B0(n9556), .Y(n9557));
  AOI21X1 g07853(.A0(n9546), .A1(n7253), .B0(n9557), .Y(n9558));
  OAI21X1 g07854(.A0(n9541), .A1(n9533), .B0(n9558), .Y(P2_U3213));
  NAND2X1 g07855(.A(n9432), .B(n7688), .Y(n9560));
  XOR2X1  g07856(.A(n9443), .B(n7695), .Y(n9561));
  NOR2X1  g07857(.A(n9561), .B(n9560), .Y(n9562));
  NAND2X1 g07858(.A(n9561), .B(n9560), .Y(n9563));
  INVX1   g07859(.A(n9563), .Y(n9564));
  NAND2X1 g07860(.A(n9432), .B(n7642), .Y(n9565));
  XOR2X1  g07861(.A(n9443), .B(n7652), .Y(n9566));
  NOR2X1  g07862(.A(n9566), .B(n9565), .Y(n9567));
  NAND2X1 g07863(.A(n9566), .B(n9565), .Y(n9568));
  NAND2X1 g07864(.A(n9432), .B(n7600), .Y(n9569));
  XOR2X1  g07865(.A(n9443), .B(n7608), .Y(n9570));
  NOR2X1  g07866(.A(n8087), .B(n7601), .Y(n9571));
  INVX1   g07867(.A(n9570), .Y(n9572));
  XOR2X1  g07868(.A(n9443), .B(n7565), .Y(n9573));
  NOR2X1  g07869(.A(n8087), .B(n7558), .Y(n9574));
  INVX1   g07870(.A(n9574), .Y(n9575));
  NOR2X1  g07871(.A(n8087), .B(n7464), .Y(n9576));
  INVX1   g07872(.A(n9576), .Y(n9577));
  XOR2X1  g07873(.A(n9443), .B(n7470), .Y(n9578));
  NOR2X1  g07874(.A(n9578), .B(n9577), .Y(n9579));
  NAND2X1 g07875(.A(n9432), .B(n7509), .Y(n9580));
  XOR2X1  g07876(.A(n9438), .B(n7517), .Y(n9581));
  AOI22X1 g07877(.A0(n9580), .A1(n9581), .B0(n9575), .B1(n9573), .Y(n9582));
  NAND2X1 g07878(.A(n9582), .B(n9579), .Y(n9583));
  INVX1   g07879(.A(n9573), .Y(n9584));
  NOR2X1  g07880(.A(n9581), .B(n9580), .Y(n9585));
  AOI21X1 g07881(.A0(n9574), .A1(n9584), .B0(n9585), .Y(n9586));
  AOI22X1 g07882(.A0(n9583), .A1(n9586), .B0(n9575), .B1(n9573), .Y(n9587));
  INVX1   g07883(.A(n9587), .Y(n9588));
  XOR2X1  g07884(.A(n9443), .B(n7425), .Y(n9589));
  NOR3X1  g07885(.A(n9589), .B(n8087), .C(n7414), .Y(n9590));
  OAI21X1 g07886(.A0(n8087), .A1(n7414), .B0(n9589), .Y(n9591));
  AOI21X1 g07887(.A0(n7303), .A1(n7297), .B0(n8087), .Y(n9592));
  INVX1   g07888(.A(n9592), .Y(n9593));
  XOR2X1  g07889(.A(n9438), .B(n7320), .Y(n9594));
  NOR2X1  g07890(.A(n8087), .B(n7360), .Y(n9595));
  INVX1   g07891(.A(n9595), .Y(n9596));
  XOR2X1  g07892(.A(n9443), .B(n7373), .Y(n9597));
  AOI22X1 g07893(.A0(n9596), .A1(n9597), .B0(n9594), .B1(n9593), .Y(n9598));
  INVX1   g07894(.A(n9531), .Y(n9599));
  NOR2X1  g07895(.A(n9599), .B(n9530), .Y(n9600));
  AOI22X1 g07896(.A0(n9530), .A1(n9599), .B0(n9528), .B1(n9514), .Y(n9601));
  OAI21X1 g07897(.A0(n9601), .A1(n9600), .B0(n9598), .Y(n9602));
  NOR2X1  g07898(.A(n9594), .B(n9593), .Y(n9603));
  INVX1   g07899(.A(n9603), .Y(n9604));
  AOI21X1 g07900(.A0(n9604), .A1(n9596), .B0(n9597), .Y(n9605));
  AOI21X1 g07901(.A0(n9603), .A1(n9595), .B0(n9605), .Y(n9606));
  NAND2X1 g07902(.A(n9606), .B(n9602), .Y(n9607));
  AOI21X1 g07903(.A0(n9607), .A1(n9591), .B0(n9590), .Y(n9608));
  NAND2X1 g07904(.A(n9578), .B(n9577), .Y(n9609));
  NAND2X1 g07905(.A(n9609), .B(n9582), .Y(n9610));
  OAI21X1 g07906(.A0(n9610), .A1(n9608), .B0(n9588), .Y(n9611));
  OAI21X1 g07907(.A0(n9572), .A1(n9571), .B0(n9611), .Y(n9612));
  OAI21X1 g07908(.A0(n9570), .A1(n9569), .B0(n9612), .Y(n9613));
  AOI21X1 g07909(.A0(n9613), .A1(n9568), .B0(n9567), .Y(n9614));
  NOR2X1  g07910(.A(n9614), .B(n9564), .Y(n9615));
  NOR2X1  g07911(.A(n9615), .B(n9562), .Y(n9616));
  XOR2X1  g07912(.A(n9438), .B(n7742), .Y(n9617));
  NOR2X1  g07913(.A(n8087), .B(n7735), .Y(n9618));
  NAND2X1 g07914(.A(n9618), .B(n9617), .Y(n9619));
  NOR2X1  g07915(.A(n8087), .B(n7780), .Y(n9620));
  XOR2X1  g07916(.A(n9438), .B(n7787), .Y(n9621));
  XOR2X1  g07917(.A(n9621), .B(n9620), .Y(n9622));
  NAND3X1 g07918(.A(n9622), .B(n9619), .C(n9616), .Y(n9623));
  AOI21X1 g07919(.A0(n9618), .A1(n9617), .B0(n9562), .Y(n9624));
  INVX1   g07920(.A(n9624), .Y(n9625));
  INVX1   g07921(.A(n9620), .Y(n9626));
  NOR2X1  g07922(.A(n9621), .B(n9626), .Y(n9627));
  NOR2X1  g07923(.A(n9618), .B(n9617), .Y(n9628));
  AOI21X1 g07924(.A0(n9621), .A1(n9626), .B0(n9628), .Y(n9629));
  INVX1   g07925(.A(n9629), .Y(n9630));
  NOR2X1  g07926(.A(n9630), .B(n9627), .Y(n9631));
  OAI21X1 g07927(.A0(n9625), .A1(n9615), .B0(n9631), .Y(n9632));
  AOI21X1 g07928(.A0(n9628), .A1(n9622), .B0(n9541), .Y(n9633));
  NAND3X1 g07929(.A(n9633), .B(n9632), .C(n9623), .Y(n9634));
  NAND4X1 g07930(.A(n8005), .B(n6447), .C(n6444), .D(n8412), .Y(n9635));
  AOI21X1 g07931(.A0(n9635), .A1(n8084), .B0(n6357), .Y(n9636));
  NAND2X1 g07932(.A(n9636), .B(n7817), .Y(n9637));
  NOR2X1  g07933(.A(n9551), .B(n7735), .Y(n9638));
  INVX1   g07934(.A(n9549), .Y(n9639));
  OAI22X1 g07935(.A0(n9534), .A1(n7775), .B0(n7825), .B1(n9639), .Y(n9640));
  OAI21X1 g07936(.A0(n9640), .A1(n9638), .B0(n9547), .Y(n9641));
  AOI22X1 g07937(.A0(n8293), .A1(n9546), .B0(P2_U3088), .B1(P2_REG3_REG_26__SCAN_IN), .Y(n9644));
  NAND4X1 g07938(.A(n9641), .B(n9637), .C(n9634), .D(n9644), .Y(P2_U3212));
  XOR2X1  g07939(.A(n9472), .B(n9471), .Y(n9646));
  INVX1   g07940(.A(n9466), .Y(n9647));
  OAI21X1 g07941(.A0(n9480), .A1(n9647), .B0(n9485), .Y(n9648));
  NAND2X1 g07942(.A(n9646), .B(n9648), .Y(n9650));
  OAI21X1 g07943(.A0(n9648), .A1(n9646), .B0(n9650), .Y(n9651));
  NAND2X1 g07944(.A(n9651), .B(n9540), .Y(n9652));
  NOR2X1  g07945(.A(n9639), .B(n6840), .Y(n9653));
  OAI22X1 g07946(.A0(n9534), .A1(n6784), .B0(n6732), .B1(n9551), .Y(n9654));
  OAI21X1 g07947(.A0(n9654), .A1(n9653), .B0(n9547), .Y(n9655));
  OAI22X1 g07948(.A0(n6832), .A1(n9554), .B0(P2_STATE_REG_SCAN_IN), .B1(n6781), .Y(n9656));
  AOI21X1 g07949(.A0(n9546), .A1(n8127), .B0(n9656), .Y(n9657));
  NAND3X1 g07950(.A(n9657), .B(n9655), .C(n9652), .Y(P2_U3211));
  NOR2X1  g07951(.A(n8087), .B(n7414), .Y(n9659));
  XOR2X1  g07952(.A(n9589), .B(n9659), .Y(n9660));
  XOR2X1  g07953(.A(n9660), .B(n9607), .Y(n9661));
  OAI22X1 g07954(.A0(n9534), .A1(n7409), .B0(n7360), .B1(n9551), .Y(n9662));
  AOI21X1 g07955(.A0(n9549), .A1(n7486), .B0(n9662), .Y(n9663));
  AOI22X1 g07956(.A0(n7425), .A1(n9636), .B0(P2_U3088), .B1(P2_REG3_REG_18__SCAN_IN), .Y(n9664));
  OAI21X1 g07957(.A0(n9663), .A1(n9548), .B0(n9664), .Y(n9665));
  AOI21X1 g07958(.A0(n9546), .A1(n7410), .B0(n9665), .Y(n9666));
  OAI21X1 g07959(.A0(n9661), .A1(n9541), .B0(n9666), .Y(P2_U3210));
  NOR2X1  g07960(.A(n9639), .B(n6626), .Y(n9668));
  OAI22X1 g07961(.A0(n9534), .A1(n6593), .B0(n6542), .B1(n9551), .Y(n9669));
  OAI21X1 g07962(.A0(n9669), .A1(n9668), .B0(n9547), .Y(n9670));
  NOR2X1  g07963(.A(n9545), .B(n6593), .Y(n9671));
  NOR2X1  g07964(.A(n9554), .B(n6601), .Y(n9672));
  OAI21X1 g07965(.A0(n6594), .A1(n6591), .B0(n9432), .Y(n9673));
  INVX1   g07966(.A(n9439), .Y(n9674));
  XOR2X1  g07967(.A(n9674), .B(n9673), .Y(n9675));
  NAND4X1 g07968(.A(n9454), .B(n9451), .C(n9448), .D(n9675), .Y(n9676));
  OAI21X1 g07969(.A0(n9458), .A1(n9440), .B0(n9455), .Y(n9677));
  AOI21X1 g07970(.A0(n9677), .A1(n9676), .B0(n9541), .Y(n9678));
  NOR4X1  g07971(.A(n9672), .B(n9671), .C(n8891), .D(n9678), .Y(n9679));
  NAND2X1 g07972(.A(n9679), .B(n9670), .Y(P2_U3209));
  NOR2X1  g07973(.A(n9494), .B(n9492), .Y(n9681));
  OAI21X1 g07974(.A0(n9510), .A1(n9681), .B0(n9518), .Y(n9682));
  INVX1   g07975(.A(n9504), .Y(n9683));
  XOR2X1  g07976(.A(n9683), .B(n9503), .Y(n9684));
  INVX1   g07977(.A(n9520), .Y(n9685));
  OAI21X1 g07978(.A0(n9685), .A1(n9505), .B0(n9682), .Y(n9686));
  OAI21X1 g07979(.A0(n9684), .A1(n9682), .B0(n9686), .Y(n9687));
  NAND2X1 g07980(.A(n9687), .B(n9540), .Y(n9688));
  NAND2X1 g07981(.A(n9546), .B(n7048), .Y(n9689));
  AOI22X1 g07982(.A0(n9535), .A1(n7048), .B0(n6992), .B1(n9550), .Y(n9690));
  OAI21X1 g07983(.A0(n9639), .A1(n7104), .B0(n9690), .Y(n9691));
  OAI22X1 g07984(.A0(n7073), .A1(n9554), .B0(P2_STATE_REG_SCAN_IN), .B1(n7045), .Y(n9692));
  AOI21X1 g07985(.A0(n9691), .A1(n9547), .B0(n9692), .Y(n9693));
  NAND3X1 g07986(.A(n9693), .B(n9689), .C(n9688), .Y(P2_U3208));
  XOR2X1  g07987(.A(n9570), .B(n9571), .Y(n9695));
  XOR2X1  g07988(.A(n9695), .B(n9611), .Y(n9696));
  NOR2X1  g07989(.A(n9639), .B(n7643), .Y(n9697));
  OAI22X1 g07990(.A0(n9534), .A1(n7596), .B0(n7558), .B1(n9551), .Y(n9698));
  OAI21X1 g07991(.A0(n9698), .A1(n9697), .B0(n9547), .Y(n9699));
  AOI22X1 g07992(.A0(n8258), .A1(n9546), .B0(P2_U3088), .B1(P2_REG3_REG_22__SCAN_IN), .Y(n9700));
  NAND2X1 g07993(.A(n9700), .B(n9699), .Y(n9701));
  AOI21X1 g07994(.A0(n9636), .A1(n7608), .B0(n9701), .Y(n9702));
  OAI21X1 g07995(.A0(n9696), .A1(n9541), .B0(n9702), .Y(P2_U3207));
  AOI21X1 g07996(.A0(n9682), .A1(n9506), .B0(n9685), .Y(n9704));
  INVX1   g07997(.A(n9704), .Y(n9705));
  AOI21X1 g07998(.A0(n9522), .A1(n9521), .B0(n9515), .Y(n9706));
  OAI21X1 g07999(.A0(n9705), .A1(n9523), .B0(n9706), .Y(n9707));
  INVX1   g08000(.A(n9500), .Y(n9708));
  INVX1   g08001(.A(n9523), .Y(n9709));
  OAI21X1 g08002(.A0(n9522), .A1(n9501), .B0(n9709), .Y(n9710));
  AOI21X1 g08003(.A0(n9522), .A1(n9501), .B0(n9710), .Y(n9711));
  OAI21X1 g08004(.A0(n9704), .A1(n9708), .B0(n9711), .Y(n9712));
  NAND3X1 g08005(.A(n9712), .B(n9707), .C(n9540), .Y(n9713));
  NAND2X1 g08006(.A(n9546), .B(n7152), .Y(n9714));
  NOR2X1  g08007(.A(n9639), .B(n7207), .Y(n9715));
  OAI22X1 g08008(.A0(n9534), .A1(n7151), .B0(n7104), .B1(n9551), .Y(n9716));
  OAI21X1 g08009(.A0(n9716), .A1(n9715), .B0(n9547), .Y(n9717));
  AOI22X1 g08010(.A0(n7164), .A1(n9636), .B0(P2_U3088), .B1(P2_REG3_REG_13__SCAN_IN), .Y(n9718));
  NAND4X1 g08011(.A(n9717), .B(n9714), .C(n9713), .D(n9718), .Y(P2_U3206));
  XOR2X1  g08012(.A(n9581), .B(n9580), .Y(n9720));
  AOI21X1 g08013(.A0(n9578), .A1(n9577), .B0(n9608), .Y(n9721));
  NOR2X1  g08014(.A(n9721), .B(n9579), .Y(n9722));
  NOR2X1  g08015(.A(n9720), .B(n9722), .Y(n9724));
  AOI21X1 g08016(.A0(n9722), .A1(n9720), .B0(n9724), .Y(n9725));
  NAND2X1 g08017(.A(n9546), .B(n8238), .Y(n9726));
  AOI22X1 g08018(.A0(n9535), .A1(n8238), .B0(n7486), .B1(n9550), .Y(n9727));
  OAI21X1 g08019(.A0(n9639), .A1(n7558), .B0(n9727), .Y(n9728));
  AOI22X1 g08020(.A0(n9547), .A1(n9728), .B0(P2_U3088), .B1(P2_REG3_REG_20__SCAN_IN), .Y(n9729));
  NAND2X1 g08021(.A(n9729), .B(n9726), .Y(n9730));
  AOI21X1 g08022(.A0(n9636), .A1(n7527), .B0(n9730), .Y(n9731));
  OAI21X1 g08023(.A0(n9725), .A1(n9541), .B0(n9731), .Y(P2_U3205));
  OAI21X1 g08024(.A0(n8082), .A1(n6357), .B0(n9548), .Y(n9733));
  AOI22X1 g08025(.A0(n9544), .A1(P2_STATE_REG_SCAN_IN), .B0(n9535), .B1(n9733), .Y(n9734));
  NOR2X1  g08026(.A(n9554), .B(n6531), .Y(n9735));
  XOR2X1  g08027(.A(n6483), .B(n9449), .Y(n9737));
  NOR4X1  g08028(.A(n9539), .B(n9535), .C(n6357), .D(n9737), .Y(n9738));
  NOR3X1  g08029(.A(n9639), .B(n9548), .C(n6542), .Y(n9739));
  NOR4X1  g08030(.A(n9738), .B(n9735), .C(n8921), .D(n9739), .Y(n9740));
  OAI21X1 g08031(.A0(n9734), .A1(n6496), .B0(n9740), .Y(P2_U3204));
  XOR2X1  g08032(.A(n9493), .B(n9435), .Y(n9742));
  XOR2X1  g08033(.A(n9742), .B(n9491), .Y(n9743));
  OAI22X1 g08034(.A0(n9534), .A1(n6941), .B0(n6895), .B1(n9551), .Y(n9744));
  AOI21X1 g08035(.A0(n9549), .A1(n6992), .B0(n9744), .Y(n9745));
  AOI22X1 g08036(.A0(n6956), .A1(n9636), .B0(P2_U3088), .B1(P2_REG3_REG_9__SCAN_IN), .Y(n9746));
  OAI21X1 g08037(.A0(n9745), .A1(n9548), .B0(n9746), .Y(n9747));
  AOI21X1 g08038(.A0(n9546), .A1(n6942), .B0(n9747), .Y(n9748));
  OAI21X1 g08039(.A0(n9743), .A1(n9541), .B0(n9748), .Y(P2_U3203));
  NOR2X1  g08040(.A(n9639), .B(n6732), .Y(n9750));
  OAI22X1 g08041(.A0(n9534), .A1(n6683), .B0(n6626), .B1(n9551), .Y(n9751));
  OAI21X1 g08042(.A0(n9751), .A1(n9750), .B0(n9547), .Y(n9752));
  NAND2X1 g08043(.A(n9546), .B(n8117), .Y(n9753));
  XOR2X1  g08044(.A(n9464), .B(n9436), .Y(n9754));
  XOR2X1  g08045(.A(n9754), .B(n9461), .Y(n9755));
  OAI22X1 g08046(.A0(n6723), .A1(n9554), .B0(P2_STATE_REG_SCAN_IN), .B1(n6682), .Y(n9756));
  AOI21X1 g08047(.A0(n9755), .A1(n9540), .B0(n9756), .Y(n9757));
  NAND3X1 g08048(.A(n9757), .B(n9753), .C(n9752), .Y(P2_U3202));
  XOR2X1  g08049(.A(n9561), .B(n9560), .Y(n9759));
  NOR2X1  g08050(.A(n9759), .B(n9614), .Y(n9761));
  AOI21X1 g08051(.A0(n9759), .A1(n9614), .B0(n9761), .Y(n9762));
  NOR2X1  g08052(.A(n9639), .B(n7735), .Y(n9763));
  OAI22X1 g08053(.A0(n9534), .A1(n7684), .B0(n7643), .B1(n9551), .Y(n9764));
  OAI21X1 g08054(.A0(n9764), .A1(n9763), .B0(n9547), .Y(n9765));
  AOI22X1 g08055(.A0(n7683), .A1(n9546), .B0(P2_U3088), .B1(P2_REG3_REG_24__SCAN_IN), .Y(n9766));
  NAND2X1 g08056(.A(n9766), .B(n9765), .Y(n9767));
  AOI21X1 g08057(.A0(n9636), .A1(n7695), .B0(n9767), .Y(n9768));
  OAI21X1 g08058(.A0(n9762), .A1(n9541), .B0(n9768), .Y(P2_U3201));
  NOR2X1  g08059(.A(n9601), .B(n9600), .Y(n9770));
  OAI21X1 g08060(.A0(n9597), .A1(n9596), .B0(n9598), .Y(n9771));
  AOI21X1 g08061(.A0(n9604), .A1(n9770), .B0(n9771), .Y(n9772));
  AOI21X1 g08062(.A0(n9594), .A1(n9593), .B0(n9770), .Y(n9773));
  INVX1   g08063(.A(n9597), .Y(n9774));
  AOI21X1 g08064(.A0(n9774), .A1(n9596), .B0(n9603), .Y(n9775));
  OAI21X1 g08065(.A0(n9774), .A1(n9596), .B0(n9775), .Y(n9776));
  OAI21X1 g08066(.A0(n9776), .A1(n9773), .B0(n9540), .Y(n9777));
  OAI22X1 g08067(.A0(n9534), .A1(n7355), .B0(n7305), .B1(n9551), .Y(n9778));
  AOI21X1 g08068(.A0(n9549), .A1(n7432), .B0(n9778), .Y(n9779));
  AOI22X1 g08069(.A0(n7373), .A1(n9636), .B0(P2_U3088), .B1(P2_REG3_REG_17__SCAN_IN), .Y(n9780));
  OAI21X1 g08070(.A0(n9779), .A1(n9548), .B0(n9780), .Y(n9781));
  AOI21X1 g08071(.A0(n9546), .A1(n7356), .B0(n9781), .Y(n9782));
  OAI21X1 g08072(.A0(n9777), .A1(n9772), .B0(n9782), .Y(P2_U3200));
  XOR2X1  g08073(.A(n9479), .B(n9478), .Y(n9784));
  XOR2X1  g08074(.A(n9784), .B(n9647), .Y(n9785));
  NAND2X1 g08075(.A(n9549), .B(n6807), .Y(n9786));
  AOI22X1 g08076(.A0(n9535), .A1(n6743), .B0(n6706), .B1(n9550), .Y(n9787));
  AOI21X1 g08077(.A0(n9787), .A1(n9786), .B0(n9548), .Y(n9788));
  NOR2X1  g08078(.A(n9545), .B(n6730), .Y(n9789));
  OAI22X1 g08079(.A0(n6753), .A1(n9554), .B0(P2_STATE_REG_SCAN_IN), .B1(n6782), .Y(n9790));
  NOR3X1  g08080(.A(n9790), .B(n9789), .C(n9788), .Y(n9791));
  OAI21X1 g08081(.A0(n9785), .A1(n9541), .B0(n9791), .Y(P2_U3199));
  XOR2X1  g08082(.A(n9594), .B(n9593), .Y(n9793));
  NOR2X1  g08083(.A(n9793), .B(n9770), .Y(n9795));
  AOI21X1 g08084(.A0(n9793), .A1(n9770), .B0(n9795), .Y(n9796));
  OAI22X1 g08085(.A0(n9534), .A1(n7301), .B0(n7312), .B1(n9551), .Y(n9797));
  AOI21X1 g08086(.A0(n9549), .A1(n7368), .B0(n9797), .Y(n9798));
  AOI22X1 g08087(.A0(n7326), .A1(n9636), .B0(P2_U3088), .B1(P2_REG3_REG_16__SCAN_IN), .Y(n9799));
  OAI21X1 g08088(.A0(n9798), .A1(n9548), .B0(n9799), .Y(n9800));
  AOI21X1 g08089(.A0(n9546), .A1(n7302), .B0(n9800), .Y(n9801));
  OAI21X1 g08090(.A0(n9796), .A1(n9541), .B0(n9801), .Y(P2_U3198));
  XOR2X1  g08091(.A(n9618), .B(n9617), .Y(n9803));
  NOR2X1  g08092(.A(n9803), .B(n9616), .Y(n9805));
  AOI21X1 g08093(.A0(n9803), .A1(n9616), .B0(n9805), .Y(n9806));
  NOR2X1  g08094(.A(n9639), .B(n7780), .Y(n9807));
  OAI22X1 g08095(.A0(n9534), .A1(n7730), .B0(n7694), .B1(n9551), .Y(n9808));
  OAI21X1 g08096(.A0(n9808), .A1(n9807), .B0(n9547), .Y(n9809));
  AOI22X1 g08097(.A0(n8285), .A1(n9546), .B0(P2_U3088), .B1(P2_REG3_REG_25__SCAN_IN), .Y(n9810));
  NAND2X1 g08098(.A(n9810), .B(n9809), .Y(n9811));
  AOI21X1 g08099(.A0(n9636), .A1(n7742), .B0(n9811), .Y(n9812));
  OAI21X1 g08100(.A0(n9806), .A1(n9541), .B0(n9812), .Y(P2_U3197));
  AOI21X1 g08101(.A0(n7102), .A1(n7098), .B0(n8087), .Y(n9814));
  XOR2X1  g08102(.A(n9814), .B(n9499), .Y(n9815));
  NOR2X1  g08103(.A(n9815), .B(n9705), .Y(n9816));
  AOI21X1 g08104(.A0(n9709), .A1(n9500), .B0(n9704), .Y(n9817));
  OAI21X1 g08105(.A0(n9817), .A1(n9816), .B0(n9540), .Y(n9818));
  NAND2X1 g08106(.A(n9546), .B(n7101), .Y(n9819));
  NOR2X1  g08107(.A(n9639), .B(n7165), .Y(n9820));
  OAI22X1 g08108(.A0(n9534), .A1(n8175), .B0(n7051), .B1(n9551), .Y(n9821));
  OAI21X1 g08109(.A0(n9821), .A1(n9820), .B0(n9547), .Y(n9822));
  AOI22X1 g08110(.A0(n7115), .A1(n9636), .B0(P2_U3088), .B1(P2_REG3_REG_12__SCAN_IN), .Y(n9823));
  NAND4X1 g08111(.A(n9822), .B(n9819), .C(n9818), .D(n9823), .Y(P2_U3196));
  NOR3X1  g08112(.A(n9721), .B(n9585), .C(n9579), .Y(n9825));
  OAI21X1 g08113(.A0(n9575), .A1(n9573), .B0(n9582), .Y(n9826));
  NOR2X1  g08114(.A(n9826), .B(n9825), .Y(n9827));
  AOI21X1 g08115(.A0(n9581), .A1(n9580), .B0(n9722), .Y(n9828));
  AOI21X1 g08116(.A0(n9575), .A1(n9584), .B0(n9585), .Y(n9829));
  OAI21X1 g08117(.A0(n9575), .A1(n9584), .B0(n9829), .Y(n9830));
  OAI21X1 g08118(.A0(n9830), .A1(n9828), .B0(n9540), .Y(n9831));
  NAND2X1 g08119(.A(n9546), .B(n8248), .Y(n9832));
  AOI22X1 g08120(.A0(n9535), .A1(n8248), .B0(n7509), .B1(n9550), .Y(n9833));
  OAI21X1 g08121(.A0(n9639), .A1(n7601), .B0(n9833), .Y(n9834));
  AOI22X1 g08122(.A0(n9547), .A1(n9834), .B0(P2_U3088), .B1(P2_REG3_REG_21__SCAN_IN), .Y(n9835));
  NAND2X1 g08123(.A(n9835), .B(n9832), .Y(n9836));
  AOI21X1 g08124(.A0(n9636), .A1(n7565), .B0(n9836), .Y(n9837));
  OAI21X1 g08125(.A0(n9831), .A1(n9827), .B0(n9837), .Y(P2_U3195));
  NOR2X1  g08126(.A(n9639), .B(n6595), .Y(n9839));
  OAI22X1 g08127(.A0(n9534), .A1(n6540), .B0(n6505), .B1(n9551), .Y(n9840));
  OAI21X1 g08128(.A0(n9840), .A1(n9839), .B0(n9547), .Y(n9841));
  NAND2X1 g08129(.A(n9546), .B(P2_REG3_REG_1__SCAN_IN), .Y(n9842));
  AOI21X1 g08130(.A0(n9438), .A1(n6531), .B0(n9450), .Y(n9843));
  XOR2X1  g08131(.A(n9453), .B(n9452), .Y(n9844));
  XOR2X1  g08132(.A(n9844), .B(n9843), .Y(n9845));
  OAI22X1 g08133(.A0(n9541), .A1(n9845), .B0(P2_STATE_REG_SCAN_IN), .B1(n6540), .Y(n9846));
  AOI21X1 g08134(.A0(n9636), .A1(n6580), .B0(n9846), .Y(n9847));
  NAND3X1 g08135(.A(n9847), .B(n9842), .C(n9841), .Y(P2_U3194));
  INVX1   g08136(.A(n9477), .Y(n9849));
  INVX1   g08137(.A(n9480), .Y(n9850));
  NAND2X1 g08138(.A(n9850), .B(n9849), .Y(n9851));
  AOI21X1 g08139(.A0(n9465), .A1(n9462), .B0(n9851), .Y(n9852));
  NOR3X1  g08140(.A(n9852), .B(n9487), .C(n9484), .Y(n9853));
  XOR2X1  g08141(.A(n9469), .B(n9468), .Y(n9854));
  XOR2X1  g08142(.A(n9854), .B(n9853), .Y(n9855));
  NAND2X1 g08143(.A(n9549), .B(n6944), .Y(n9856));
  AOI22X1 g08144(.A0(n9535), .A1(n6892), .B0(n6839), .B1(n9550), .Y(n9857));
  AOI21X1 g08145(.A0(n9857), .A1(n9856), .B0(n9548), .Y(n9858));
  NOR2X1  g08146(.A(n9545), .B(n6891), .Y(n9859));
  OAI22X1 g08147(.A0(n6935), .A1(n9554), .B0(P2_STATE_REG_SCAN_IN), .B1(n6888), .Y(n9860));
  NOR3X1  g08148(.A(n9860), .B(n9859), .C(n9858), .Y(n9861));
  OAI21X1 g08149(.A0(n9855), .A1(n9541), .B0(n9861), .Y(P2_U3193));
  XOR2X1  g08150(.A(n9443), .B(n7893), .Y(n9863));
  NOR2X1  g08151(.A(n8087), .B(n7886), .Y(n9864));
  XOR2X1  g08152(.A(n9864), .B(n9863), .Y(n9865));
  XOR2X1  g08153(.A(n9438), .B(n7848), .Y(n9866));
  INVX1   g08154(.A(n9866), .Y(n9867));
  NOR2X1  g08155(.A(n8087), .B(n7825), .Y(n9868));
  NOR2X1  g08156(.A(n9868), .B(n9867), .Y(n9869));
  NOR4X1  g08157(.A(n9630), .B(n9614), .C(n9564), .D(n9869), .Y(n9870));
  NOR2X1  g08158(.A(n9629), .B(n9627), .Y(n9871));
  NOR2X1  g08159(.A(n9627), .B(n9625), .Y(n9872));
  NOR3X1  g08160(.A(n9872), .B(n9871), .C(n9869), .Y(n9873));
  NOR3X1  g08161(.A(n9866), .B(n8087), .C(n7825), .Y(n9874));
  NOR4X1  g08162(.A(n9873), .B(n9870), .C(n9865), .D(n9874), .Y(n9875));
  INVX1   g08163(.A(n9614), .Y(n9876));
  NAND3X1 g08164(.A(n9629), .B(n9876), .C(n9563), .Y(n9877));
  OAI21X1 g08165(.A0(n9618), .A1(n9617), .B0(n9625), .Y(n9878));
  AOI21X1 g08166(.A0(n9621), .A1(n9626), .B0(n9878), .Y(n9879));
  NOR3X1  g08167(.A(n9879), .B(n9874), .C(n9627), .Y(n9880));
  AOI21X1 g08168(.A0(n9880), .A1(n9877), .B0(n9869), .Y(n9881));
  AOI21X1 g08169(.A0(n9881), .A1(n9865), .B0(n9875), .Y(n9882));
  NOR2X1  g08170(.A(n9639), .B(n7932), .Y(n9883));
  OAI22X1 g08171(.A0(n9534), .A1(n7881), .B0(n7825), .B1(n9551), .Y(n9884));
  OAI21X1 g08172(.A0(n9884), .A1(n9883), .B0(n9547), .Y(n9885));
  AOI22X1 g08173(.A0(n8309), .A1(n9546), .B0(P2_U3088), .B1(P2_REG3_REG_28__SCAN_IN), .Y(n9886));
  NAND2X1 g08174(.A(n9886), .B(n9885), .Y(n9887));
  AOI21X1 g08175(.A0(n9636), .A1(n7893), .B0(n9887), .Y(n9888));
  OAI21X1 g08176(.A0(n9882), .A1(n9541), .B0(n9888), .Y(P2_U3192));
  XOR2X1  g08177(.A(n9578), .B(n9577), .Y(n9890));
  NOR2X1  g08178(.A(n9890), .B(n9608), .Y(n9892));
  AOI21X1 g08179(.A0(n9890), .A1(n9608), .B0(n9892), .Y(n9893));
  AOI22X1 g08180(.A0(n9535), .A1(n7460), .B0(n7432), .B1(n9550), .Y(n9894));
  OAI21X1 g08181(.A0(n9639), .A1(n7510), .B0(n9894), .Y(n9895));
  AOI22X1 g08182(.A0(n9547), .A1(n9895), .B0(P2_U3088), .B1(P2_REG3_REG_19__SCAN_IN), .Y(n9896));
  OAI21X1 g08183(.A0(n9545), .A1(n7459), .B0(n9896), .Y(n9897));
  AOI21X1 g08184(.A0(n9636), .A1(n7470), .B0(n9897), .Y(n9898));
  OAI21X1 g08185(.A0(n9893), .A1(n9541), .B0(n9898), .Y(P2_U3191));
  NOR2X1  g08186(.A(n9639), .B(n6685), .Y(n9900));
  OAI22X1 g08187(.A0(n9534), .A1(P2_REG3_REG_3__SCAN_IN), .B0(n6595), .B1(n9551), .Y(n9901));
  OAI21X1 g08188(.A0(n9901), .A1(n9900), .B0(n9547), .Y(n9902));
  NAND2X1 g08189(.A(n9546), .B(n6650), .Y(n9903));
  NAND2X1 g08190(.A(n9636), .B(n6646), .Y(n9904));
  NAND4X1 g08191(.A(n9454), .B(n9451), .C(n9448), .D(n9457), .Y(n9905));
  INVX1   g08192(.A(n9444), .Y(n9906));
  NAND2X1 g08193(.A(n9906), .B(n9441), .Y(n9907));
  NAND3X1 g08194(.A(n9907), .B(n9905), .C(n9445), .Y(n9908));
  INVX1   g08195(.A(n9440), .Y(n9909));
  AOI21X1 g08196(.A0(n9906), .A1(n9442), .B0(n9458), .Y(n9910));
  OAI21X1 g08197(.A0(n9906), .A1(n9442), .B0(n9910), .Y(n9911));
  AOI21X1 g08198(.A0(n9455), .A1(n9909), .B0(n9911), .Y(n9912));
  NOR4X1  g08199(.A(n9539), .B(n9535), .C(n6357), .D(n9912), .Y(n9913));
  AOI22X1 g08200(.A0(n9908), .A1(n9913), .B0(P2_U3088), .B1(P2_REG3_REG_3__SCAN_IN), .Y(n9914));
  NAND4X1 g08201(.A(n9904), .B(n9903), .C(n9902), .D(n9914), .Y(P2_U3190));
  XOR2X1  g08202(.A(n9508), .B(n9516), .Y(n9916));
  XOR2X1  g08203(.A(n9916), .B(n9681), .Y(n9917));
  OAI22X1 g08204(.A0(n9534), .A1(n6989), .B0(n6945), .B1(n9551), .Y(n9918));
  AOI21X1 g08205(.A0(n9549), .A1(n7072), .B0(n9918), .Y(n9919));
  AOI22X1 g08206(.A0(n7004), .A1(n9636), .B0(P2_U3088), .B1(P2_REG3_REG_10__SCAN_IN), .Y(n9920));
  OAI21X1 g08207(.A0(n9919), .A1(n9548), .B0(n9920), .Y(n9921));
  AOI21X1 g08208(.A0(n9546), .A1(n6990), .B0(n9921), .Y(n9922));
  OAI21X1 g08209(.A0(n9917), .A1(n9541), .B0(n9922), .Y(P2_U3189));
  XOR2X1  g08210(.A(n9566), .B(n9565), .Y(n9924));
  XOR2X1  g08211(.A(n9924), .B(n9613), .Y(n9925));
  NAND2X1 g08212(.A(n9925), .B(n9540), .Y(n9926));
  NAND2X1 g08213(.A(n9636), .B(n7652), .Y(n9927));
  NOR2X1  g08214(.A(n9639), .B(n7694), .Y(n9928));
  OAI22X1 g08215(.A0(n9534), .A1(n7638), .B0(n7601), .B1(n9551), .Y(n9929));
  OAI21X1 g08216(.A0(n9929), .A1(n9928), .B0(n9547), .Y(n9930));
  AOI22X1 g08217(.A0(n8264), .A1(n9546), .B0(P2_U3088), .B1(P2_REG3_REG_23__SCAN_IN), .Y(n9931));
  NAND4X1 g08218(.A(n9930), .B(n9927), .C(n9926), .D(n9931), .Y(P2_U3188));
  OAI21X1 g08219(.A0(n9512), .A1(n9681), .B0(n9526), .Y(n9933));
  XOR2X1  g08220(.A(n9497), .B(n9495), .Y(n9934));
  XOR2X1  g08221(.A(n9934), .B(n9933), .Y(n9935));
  OAI22X1 g08222(.A0(n9534), .A1(n7203), .B0(n7165), .B1(n9551), .Y(n9936));
  AOI21X1 g08223(.A0(n9549), .A1(n7255), .B0(n9936), .Y(n9937));
  AOI22X1 g08224(.A0(n7249), .A1(n9636), .B0(P2_U3088), .B1(P2_REG3_REG_14__SCAN_IN), .Y(n9938));
  OAI21X1 g08225(.A0(n9937), .A1(n9548), .B0(n9938), .Y(n9939));
  AOI21X1 g08226(.A0(n9546), .A1(n7204), .B0(n9939), .Y(n9940));
  OAI21X1 g08227(.A0(n9935), .A1(n9541), .B0(n9940), .Y(P2_U3187));
  OAI21X1 g08228(.A0(n9872), .A1(n9871), .B0(n9877), .Y(n9942));
  XOR2X1  g08229(.A(n9868), .B(n9866), .Y(n9943));
  XOR2X1  g08230(.A(n9943), .B(n9942), .Y(n9944));
  NOR2X1  g08231(.A(n9639), .B(n7886), .Y(n9945));
  OAI22X1 g08232(.A0(n9534), .A1(n7820), .B0(n7780), .B1(n9551), .Y(n9946));
  OAI21X1 g08233(.A0(n9946), .A1(n9945), .B0(n9547), .Y(n9947));
  AOI22X1 g08234(.A0(n8302), .A1(n9546), .B0(P2_U3088), .B1(P2_REG3_REG_27__SCAN_IN), .Y(n9948));
  NAND2X1 g08235(.A(n9948), .B(n9947), .Y(n9949));
  AOI21X1 g08236(.A0(n9636), .A1(n7876), .B0(n9949), .Y(n9950));
  OAI21X1 g08237(.A0(n9944), .A1(n9541), .B0(n9950), .Y(P2_U3186));
  AOI21X1 g08238(.A0(n9476), .A1(n9474), .B0(n9477), .Y(n9952));
  OAI21X1 g08239(.A0(n9648), .A1(n9482), .B0(n9952), .Y(n9953));
  OAI21X1 g08240(.A0(n9473), .A1(n9471), .B0(n9648), .Y(n9954));
  OAI21X1 g08241(.A0(n6785), .A1(n6779), .B0(n9432), .Y(n9955));
  OAI22X1 g08242(.A0(n9474), .A1(n9475), .B0(n9472), .B1(n9955), .Y(n9956));
  AOI21X1 g08243(.A0(n9475), .A1(n9474), .B0(n9956), .Y(n9957));
  NAND2X1 g08244(.A(n9957), .B(n9954), .Y(n9958));
  NAND3X1 g08245(.A(n9958), .B(n9953), .C(n9540), .Y(n9959));
  NOR2X1  g08246(.A(n9639), .B(n6895), .Y(n9960));
  OAI22X1 g08247(.A0(n9534), .A1(n6836), .B0(n6786), .B1(n9551), .Y(n9961));
  OAI21X1 g08248(.A0(n9961), .A1(n9960), .B0(n9547), .Y(n9962));
  OAI22X1 g08249(.A0(n6886), .A1(n9554), .B0(P2_STATE_REG_SCAN_IN), .B1(n6889), .Y(n9963));
  AOI21X1 g08250(.A0(n9546), .A1(n6837), .B0(n9963), .Y(n9964));
  NAND3X1 g08251(.A(n9964), .B(n9962), .C(n9959), .Y(P2_U3185));
  NOR2X1  g08252(.A(n6349), .B(n6342), .Y(n9966));
  NAND3X1 g08253(.A(n8073), .B(n6750), .C(n9966), .Y(n9967));
  AOI21X1 g08254(.A0(n6750), .A1(n6342), .B0(P2_U3088), .Y(n9968));
  NAND2X1 g08255(.A(n9968), .B(n9967), .Y(P2_U3087));
  XOR2X1  g08256(.A(P2_DATAO_REG_0__SCAN_IN), .B(n1796), .Y(n9970));
  AOI21X1 g08257(.A0(n1789), .A1(n1786), .B0(n9970), .Y(n9971));
  AOI21X1 g08258(.A0(n1837), .A1(SI_0_), .B0(n9971), .Y(n9972));
  NAND2X1 g08259(.A(P3_IR_REG_0__SCAN_IN), .B(P3_STATE_REG_SCAN_IN), .Y(n9973));
  OAI21X1 g08260(.A0(n9972), .A1(P3_STATE_REG_SCAN_IN), .B0(n9973), .Y(P3_U3295));
  NOR3X1  g08261(.A(n1793), .B(n1792), .C(n1822), .Y(n9975));
  NAND2X1 g08262(.A(P2_DATAO_REG_0__SCAN_IN), .B(n1796), .Y(n9976));
  XOR2X1  g08263(.A(P2_DATAO_REG_1__SCAN_IN), .B(n1808), .Y(n9977));
  XOR2X1  g08264(.A(n9977), .B(n9976), .Y(n9978));
  AOI21X1 g08265(.A0(n9978), .A1(n1790), .B0(n9975), .Y(n9979));
  INVX1   g08266(.A(P3_STATE_REG_SCAN_IN), .Y(P3_U3151));
  NOR2X1  g08267(.A(P3_IR_REG_31__SCAN_IN), .B(P3_U3151), .Y(n9981));
  INVX1   g08268(.A(P3_IR_REG_31__SCAN_IN), .Y(n9982));
  NOR2X1  g08269(.A(n9982), .B(P3_U3151), .Y(n9983));
  INVX1   g08270(.A(P3_IR_REG_0__SCAN_IN), .Y(n9984));
  XOR2X1  g08271(.A(P3_IR_REG_1__SCAN_IN), .B(n9984), .Y(n9985));
  INVX1   g08272(.A(n9985), .Y(n9986));
  AOI22X1 g08273(.A0(n9983), .A1(n9986), .B0(n9981), .B1(P3_IR_REG_1__SCAN_IN), .Y(n9987));
  OAI21X1 g08274(.A0(n9979), .A1(P3_STATE_REG_SCAN_IN), .B0(n9987), .Y(P3_U3294));
  NOR3X1  g08275(.A(n1793), .B(n1792), .C(n1850), .Y(n9989));
  XOR2X1  g08276(.A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), .Y(n9990));
  NOR2X1  g08277(.A(n1791), .B(P1_DATAO_REG_0__SCAN_IN), .Y(n9991));
  AOI21X1 g08278(.A0(n9991), .A1(n1808), .B0(P2_DATAO_REG_1__SCAN_IN), .Y(n9992));
  AOI21X1 g08279(.A0(n9976), .A1(P1_DATAO_REG_1__SCAN_IN), .B0(n9992), .Y(n9993));
  XOR2X1  g08280(.A(n9993), .B(n9990), .Y(n9994));
  AOI21X1 g08281(.A0(n9994), .A1(n1790), .B0(n9989), .Y(n9995));
  INVX1   g08282(.A(P3_IR_REG_1__SCAN_IN), .Y(n9996));
  NAND2X1 g08283(.A(n9996), .B(n9984), .Y(n9997));
  XOR2X1  g08284(.A(n9997), .B(P3_IR_REG_2__SCAN_IN), .Y(n9998));
  AOI22X1 g08285(.A0(n9983), .A1(n9998), .B0(n9981), .B1(P3_IR_REG_2__SCAN_IN), .Y(n9999));
  OAI21X1 g08286(.A0(n9995), .A1(P3_STATE_REG_SCAN_IN), .B0(n9999), .Y(P3_U3293));
  NOR3X1  g08287(.A(n1793), .B(n1792), .C(n1912), .Y(n10001));
  XOR2X1  g08288(.A(P2_DATAO_REG_3__SCAN_IN), .B(P1_DATAO_REG_3__SCAN_IN), .Y(n10002));
  AOI21X1 g08289(.A0(P2_DATAO_REG_2__SCAN_IN), .A1(n1854), .B0(n9993), .Y(n10003));
  AOI21X1 g08290(.A0(n1832), .A1(P1_DATAO_REG_2__SCAN_IN), .B0(n10003), .Y(n10004));
  XOR2X1  g08291(.A(n10004), .B(n10002), .Y(n10005));
  AOI21X1 g08292(.A0(n10005), .A1(n1790), .B0(n10001), .Y(n10006));
  INVX1   g08293(.A(P3_IR_REG_3__SCAN_IN), .Y(n10007));
  NOR3X1  g08294(.A(P3_IR_REG_2__SCAN_IN), .B(P3_IR_REG_1__SCAN_IN), .C(P3_IR_REG_0__SCAN_IN), .Y(n10008));
  XOR2X1  g08295(.A(n10008), .B(n10007), .Y(n10009));
  AOI22X1 g08296(.A0(n9983), .A1(n10009), .B0(n9981), .B1(P3_IR_REG_3__SCAN_IN), .Y(n10010));
  OAI21X1 g08297(.A0(n10006), .A1(P3_STATE_REG_SCAN_IN), .B0(n10010), .Y(P3_U3292));
  NOR3X1  g08298(.A(n1793), .B(n1792), .C(n1901), .Y(n10012));
  XOR2X1  g08299(.A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), .Y(n10013));
  OAI21X1 g08300(.A0(n9976), .A1(P1_DATAO_REG_1__SCAN_IN), .B0(n1806), .Y(n10014));
  OAI21X1 g08301(.A0(n9991), .A1(n1808), .B0(n10014), .Y(n10015));
  AOI22X1 g08302(.A0(n1832), .A1(P1_DATAO_REG_2__SCAN_IN), .B0(P1_DATAO_REG_3__SCAN_IN), .B1(n1848), .Y(n10016));
  AOI21X1 g08303(.A0(P2_DATAO_REG_3__SCAN_IN), .A1(n1875), .B0(n10016), .Y(n10017));
  AOI22X1 g08304(.A0(P2_DATAO_REG_2__SCAN_IN), .A1(n1854), .B0(n1875), .B1(P2_DATAO_REG_3__SCAN_IN), .Y(n10018));
  AOI21X1 g08305(.A0(n10018), .A1(n10015), .B0(n10017), .Y(n10019));
  XOR2X1  g08306(.A(n10019), .B(n10013), .Y(n10020));
  AOI21X1 g08307(.A0(n10020), .A1(n1790), .B0(n10012), .Y(n10021));
  INVX1   g08308(.A(P3_IR_REG_4__SCAN_IN), .Y(n10022));
  NOR4X1  g08309(.A(P3_IR_REG_2__SCAN_IN), .B(P3_IR_REG_1__SCAN_IN), .C(P3_IR_REG_0__SCAN_IN), .D(P3_IR_REG_3__SCAN_IN), .Y(n10023));
  NAND3X1 g08310(.A(n10008), .B(n10022), .C(n10007), .Y(n10024));
  OAI21X1 g08311(.A0(n10023), .A1(n10022), .B0(n10024), .Y(n10025));
  NOR3X1  g08312(.A(n10025), .B(n9982), .C(P3_U3151), .Y(n10026));
  AOI21X1 g08313(.A0(n9981), .A1(P3_IR_REG_4__SCAN_IN), .B0(n10026), .Y(n10027));
  OAI21X1 g08314(.A0(n10021), .A1(P3_STATE_REG_SCAN_IN), .B0(n10027), .Y(P3_U3291));
  XOR2X1  g08315(.A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), .Y(n10029));
  OAI21X1 g08316(.A0(n1871), .A1(P1_DATAO_REG_4__SCAN_IN), .B0(n10018), .Y(n10030));
  OAI22X1 g08317(.A0(n1848), .A1(P1_DATAO_REG_3__SCAN_IN), .B0(P1_DATAO_REG_4__SCAN_IN), .B1(n1871), .Y(n10031));
  NOR2X1  g08318(.A(n10031), .B(n10016), .Y(n10032));
  AOI21X1 g08319(.A0(n1871), .A1(P1_DATAO_REG_4__SCAN_IN), .B0(n10032), .Y(n10033));
  OAI21X1 g08320(.A0(n10030), .A1(n9993), .B0(n10033), .Y(n10034));
  XOR2X1  g08321(.A(n10034), .B(n10029), .Y(n10035));
  NOR2X1  g08322(.A(n10035), .B(n1837), .Y(n10036));
  AOI21X1 g08323(.A0(n1837), .A1(SI_5_), .B0(n10036), .Y(n10037));
  XOR2X1  g08324(.A(n10024), .B(P3_IR_REG_5__SCAN_IN), .Y(n10038));
  AOI22X1 g08325(.A0(n9983), .A1(n10038), .B0(n9981), .B1(P3_IR_REG_5__SCAN_IN), .Y(n10039));
  OAI21X1 g08326(.A0(n10037), .A1(P3_STATE_REG_SCAN_IN), .B0(n10039), .Y(P3_U3290));
  NOR3X1  g08327(.A(n1793), .B(n1792), .C(n1955), .Y(n10041));
  XOR2X1  g08328(.A(P2_DATAO_REG_6__SCAN_IN), .B(n1935), .Y(n10042));
  OAI21X1 g08329(.A0(n1898), .A1(P1_DATAO_REG_5__SCAN_IN), .B0(n10034), .Y(n10043));
  OAI21X1 g08330(.A0(P2_DATAO_REG_5__SCAN_IN), .A1(n1904), .B0(n10043), .Y(n10044));
  XOR2X1  g08331(.A(n10044), .B(n10042), .Y(n10045));
  AOI21X1 g08332(.A0(n10045), .A1(n1790), .B0(n10041), .Y(n10046));
  INVX1   g08333(.A(P3_IR_REG_5__SCAN_IN), .Y(n10047));
  NAND4X1 g08334(.A(n10047), .B(n10022), .C(n10007), .D(n10008), .Y(n10048));
  INVX1   g08335(.A(P3_IR_REG_6__SCAN_IN), .Y(n10049));
  NAND2X1 g08336(.A(n10049), .B(n10047), .Y(n10050));
  NOR2X1  g08337(.A(n10050), .B(n10024), .Y(n10051));
  AOI21X1 g08338(.A0(n10048), .A1(P3_IR_REG_6__SCAN_IN), .B0(n10051), .Y(n10052));
  AOI22X1 g08339(.A0(n9983), .A1(n10052), .B0(n9981), .B1(P3_IR_REG_6__SCAN_IN), .Y(n10053));
  OAI21X1 g08340(.A0(n10046), .A1(P3_STATE_REG_SCAN_IN), .B0(n10053), .Y(P3_U3289));
  XOR2X1  g08341(.A(P2_DATAO_REG_7__SCAN_IN), .B(n1963), .Y(n10055));
  OAI22X1 g08342(.A0(n1898), .A1(P1_DATAO_REG_5__SCAN_IN), .B0(P1_DATAO_REG_6__SCAN_IN), .B1(n1927), .Y(n10056));
  INVX1   g08343(.A(n10056), .Y(n10057));
  NAND2X1 g08344(.A(P2_DATAO_REG_6__SCAN_IN), .B(n1935), .Y(n10058));
  NAND3X1 g08345(.A(n10058), .B(n1898), .C(P1_DATAO_REG_5__SCAN_IN), .Y(n10059));
  OAI21X1 g08346(.A0(P2_DATAO_REG_6__SCAN_IN), .A1(n1935), .B0(n10059), .Y(n10060));
  AOI21X1 g08347(.A0(n10057), .A1(n10034), .B0(n10060), .Y(n10061));
  XOR2X1  g08348(.A(n10061), .B(n10055), .Y(n10062));
  NOR2X1  g08349(.A(n10062), .B(n1837), .Y(n10063));
  AOI21X1 g08350(.A0(n1837), .A1(SI_7_), .B0(n10063), .Y(n10064));
  INVX1   g08351(.A(P3_IR_REG_7__SCAN_IN), .Y(n10065));
  XOR2X1  g08352(.A(n10051), .B(n10065), .Y(n10066));
  AOI22X1 g08353(.A0(n9983), .A1(n10066), .B0(n9981), .B1(P3_IR_REG_7__SCAN_IN), .Y(n10067));
  OAI21X1 g08354(.A0(n10064), .A1(P3_STATE_REG_SCAN_IN), .B0(n10067), .Y(P3_U3288));
  XOR2X1  g08355(.A(P2_DATAO_REG_8__SCAN_IN), .B(n5069), .Y(n10069));
  AOI21X1 g08356(.A0(P2_DATAO_REG_7__SCAN_IN), .A1(n1963), .B0(n10056), .Y(n10070));
  AOI22X1 g08357(.A0(n1927), .A1(P1_DATAO_REG_6__SCAN_IN), .B0(P1_DATAO_REG_7__SCAN_IN), .B1(n1950), .Y(n10071));
  AOI22X1 g08358(.A0(n10059), .A1(n10071), .B0(P2_DATAO_REG_7__SCAN_IN), .B1(n1963), .Y(n10072));
  AOI21X1 g08359(.A0(n10070), .A1(n10034), .B0(n10072), .Y(n10073));
  XOR2X1  g08360(.A(n10073), .B(n10069), .Y(n10074));
  NOR2X1  g08361(.A(n10074), .B(n1837), .Y(n10075));
  AOI21X1 g08362(.A0(n1837), .A1(SI_8_), .B0(n10075), .Y(n10076));
  INVX1   g08363(.A(P3_IR_REG_8__SCAN_IN), .Y(n10077));
  AOI21X1 g08364(.A0(n10051), .A1(n10065), .B0(n10077), .Y(n10078));
  NOR4X1  g08365(.A(n10024), .B(P3_IR_REG_8__SCAN_IN), .C(P3_IR_REG_7__SCAN_IN), .D(n10050), .Y(n10079));
  NOR2X1  g08366(.A(n10079), .B(n10078), .Y(n10080));
  AOI22X1 g08367(.A0(n9983), .A1(n10080), .B0(n9981), .B1(P3_IR_REG_8__SCAN_IN), .Y(n10081));
  OAI21X1 g08368(.A0(n10076), .A1(P3_STATE_REG_SCAN_IN), .B0(n10081), .Y(P3_U3287));
  INVX1   g08369(.A(SI_9_), .Y(n10083));
  NOR3X1  g08370(.A(n1793), .B(n1792), .C(n10083), .Y(n10084));
  XOR2X1  g08371(.A(P2_DATAO_REG_9__SCAN_IN), .B(n2020), .Y(n10085));
  OAI22X1 g08372(.A0(n1832), .A1(P1_DATAO_REG_2__SCAN_IN), .B0(P1_DATAO_REG_3__SCAN_IN), .B1(n1848), .Y(n10086));
  AOI21X1 g08373(.A0(P2_DATAO_REG_4__SCAN_IN), .A1(n1884), .B0(n10086), .Y(n10087));
  OAI22X1 g08374(.A0(n10016), .A1(n10031), .B0(P2_DATAO_REG_4__SCAN_IN), .B1(n1884), .Y(n10088));
  AOI21X1 g08375(.A0(n10087), .A1(n10015), .B0(n10088), .Y(n10089));
  NAND2X1 g08376(.A(P2_DATAO_REG_8__SCAN_IN), .B(n5069), .Y(n10090));
  NAND2X1 g08377(.A(n10070), .B(n10090), .Y(n10091));
  NOR2X1  g08378(.A(P2_DATAO_REG_8__SCAN_IN), .B(n5069), .Y(n10092));
  AOI21X1 g08379(.A0(n10072), .A1(n10090), .B0(n10092), .Y(n10093));
  OAI21X1 g08380(.A0(n10091), .A1(n10089), .B0(n10093), .Y(n10094));
  XOR2X1  g08381(.A(n10094), .B(n10085), .Y(n10095));
  AOI21X1 g08382(.A0(n10095), .A1(n1790), .B0(n10084), .Y(n10096));
  INVX1   g08383(.A(P3_IR_REG_9__SCAN_IN), .Y(n10097));
  XOR2X1  g08384(.A(n10079), .B(n10097), .Y(n10098));
  AOI22X1 g08385(.A0(n9983), .A1(n10098), .B0(n9981), .B1(P3_IR_REG_9__SCAN_IN), .Y(n10099));
  OAI21X1 g08386(.A0(n10096), .A1(P3_STATE_REG_SCAN_IN), .B0(n10099), .Y(P3_U3286));
  XOR2X1  g08387(.A(P2_DATAO_REG_10__SCAN_IN), .B(n2045), .Y(n10101));
  NOR2X1  g08388(.A(P2_DATAO_REG_9__SCAN_IN), .B(n2020), .Y(n10102));
  NAND2X1 g08389(.A(P2_DATAO_REG_9__SCAN_IN), .B(n2020), .Y(n10103));
  AOI21X1 g08390(.A0(n10094), .A1(n10103), .B0(n10102), .Y(n10104));
  XOR2X1  g08391(.A(n10104), .B(n10101), .Y(n10105));
  NOR2X1  g08392(.A(n10105), .B(n1837), .Y(n10106));
  AOI21X1 g08393(.A0(n1837), .A1(SI_10_), .B0(n10106), .Y(n10107));
  INVX1   g08394(.A(P3_IR_REG_10__SCAN_IN), .Y(n10108));
  AOI21X1 g08395(.A0(n10079), .A1(n10097), .B0(n10108), .Y(n10109));
  NOR2X1  g08396(.A(P3_IR_REG_10__SCAN_IN), .B(P3_IR_REG_9__SCAN_IN), .Y(n10110));
  AOI21X1 g08397(.A0(n10110), .A1(n10079), .B0(n10109), .Y(n10111));
  AOI22X1 g08398(.A0(n9983), .A1(n10111), .B0(n9981), .B1(P3_IR_REG_10__SCAN_IN), .Y(n10112));
  OAI21X1 g08399(.A0(n10107), .A1(P3_STATE_REG_SCAN_IN), .B0(n10112), .Y(P3_U3285));
  XOR2X1  g08400(.A(P2_DATAO_REG_11__SCAN_IN), .B(n5076), .Y(n10114));
  OAI21X1 g08401(.A0(n2018), .A1(P1_DATAO_REG_10__SCAN_IN), .B0(n10102), .Y(n10115));
  OAI21X1 g08402(.A0(P2_DATAO_REG_10__SCAN_IN), .A1(n2045), .B0(n10115), .Y(n10116));
  AOI22X1 g08403(.A0(P2_DATAO_REG_9__SCAN_IN), .A1(n2020), .B0(n2045), .B1(P2_DATAO_REG_10__SCAN_IN), .Y(n10117));
  AOI21X1 g08404(.A0(n10117), .A1(n10094), .B0(n10116), .Y(n10118));
  XOR2X1  g08405(.A(n10118), .B(n10114), .Y(n10119));
  NOR2X1  g08406(.A(n10119), .B(n1837), .Y(n10120));
  AOI21X1 g08407(.A0(n1837), .A1(SI_11_), .B0(n10120), .Y(n10121));
  INVX1   g08408(.A(P3_IR_REG_11__SCAN_IN), .Y(n10122));
  INVX1   g08409(.A(n10079), .Y(n10123));
  INVX1   g08410(.A(n10110), .Y(n10124));
  NOR2X1  g08411(.A(n10124), .B(n10123), .Y(n10125));
  XOR2X1  g08412(.A(n10125), .B(n10122), .Y(n10126));
  AOI22X1 g08413(.A0(n9983), .A1(n10126), .B0(n9981), .B1(P3_IR_REG_11__SCAN_IN), .Y(n10127));
  OAI21X1 g08414(.A0(n10121), .A1(P3_STATE_REG_SCAN_IN), .B0(n10127), .Y(P3_U3284));
  NOR3X1  g08415(.A(n1793), .B(n1792), .C(n2075), .Y(n10129));
  XOR2X1  g08416(.A(P2_DATAO_REG_12__SCAN_IN), .B(n5079), .Y(n10130));
  NOR2X1  g08417(.A(P2_DATAO_REG_11__SCAN_IN), .B(n5076), .Y(n10131));
  NOR2X1  g08418(.A(n2043), .B(P1_DATAO_REG_11__SCAN_IN), .Y(n10132));
  INVX1   g08419(.A(n10132), .Y(n10133));
  AOI21X1 g08420(.A0(n10116), .A1(n10133), .B0(n10131), .Y(n10134));
  INVX1   g08421(.A(n10117), .Y(n10135));
  NOR2X1  g08422(.A(n10135), .B(n10132), .Y(n10136));
  NAND2X1 g08423(.A(n10136), .B(n10094), .Y(n10137));
  NAND2X1 g08424(.A(n10137), .B(n10134), .Y(n10138));
  XOR2X1  g08425(.A(n10138), .B(n10130), .Y(n10139));
  AOI21X1 g08426(.A0(n10139), .A1(n1790), .B0(n10129), .Y(n10140));
  NAND3X1 g08427(.A(n10110), .B(n10079), .C(n10122), .Y(n10141));
  NOR4X1  g08428(.A(n10123), .B(P3_IR_REG_12__SCAN_IN), .C(P3_IR_REG_11__SCAN_IN), .D(n10124), .Y(n10142));
  AOI21X1 g08429(.A0(n10141), .A1(P3_IR_REG_12__SCAN_IN), .B0(n10142), .Y(n10143));
  AOI22X1 g08430(.A0(n9983), .A1(n10143), .B0(n9981), .B1(P3_IR_REG_12__SCAN_IN), .Y(n10144));
  OAI21X1 g08431(.A0(n10140), .A1(P3_STATE_REG_SCAN_IN), .B0(n10144), .Y(P3_U3283));
  NAND3X1 g08432(.A(n1789), .B(n1786), .C(SI_13_), .Y(n10146));
  XOR2X1  g08433(.A(P2_DATAO_REG_13__SCAN_IN), .B(n2099), .Y(n10147));
  NOR2X1  g08434(.A(n2065), .B(P1_DATAO_REG_12__SCAN_IN), .Y(n10148));
  NOR3X1  g08435(.A(n10148), .B(n10135), .C(n10132), .Y(n10149));
  NAND2X1 g08436(.A(n2065), .B(P1_DATAO_REG_12__SCAN_IN), .Y(n10150));
  OAI21X1 g08437(.A0(n10134), .A1(n10148), .B0(n10150), .Y(n10151));
  AOI21X1 g08438(.A0(n10149), .A1(n10094), .B0(n10151), .Y(n10152));
  XOR2X1  g08439(.A(n10152), .B(n10147), .Y(n10153));
  OAI21X1 g08440(.A0(n10153), .A1(n1837), .B0(n10146), .Y(n10154));
  NAND2X1 g08441(.A(n10154), .B(P3_U3151), .Y(n10155));
  INVX1   g08442(.A(P3_IR_REG_13__SCAN_IN), .Y(n10156));
  XOR2X1  g08443(.A(n10142), .B(n10156), .Y(n10157));
  AOI22X1 g08444(.A0(n9983), .A1(n10157), .B0(n9981), .B1(P3_IR_REG_13__SCAN_IN), .Y(n10158));
  NAND2X1 g08445(.A(n10158), .B(n10155), .Y(P3_U3282));
  NOR3X1  g08446(.A(n1793), .B(n1792), .C(n2130), .Y(n10160));
  XOR2X1  g08447(.A(P2_DATAO_REG_14__SCAN_IN), .B(n2131), .Y(n10161));
  NOR2X1  g08448(.A(P2_DATAO_REG_13__SCAN_IN), .B(n2099), .Y(n10162));
  INVX1   g08449(.A(n10162), .Y(n10163));
  NOR2X1  g08450(.A(n2088), .B(P1_DATAO_REG_13__SCAN_IN), .Y(n10164));
  OAI21X1 g08451(.A0(n10152), .A1(n10164), .B0(n10163), .Y(n10165));
  XOR2X1  g08452(.A(n10165), .B(n10161), .Y(n10166));
  AOI21X1 g08453(.A0(n10166), .A1(n1790), .B0(n10160), .Y(n10167));
  INVX1   g08454(.A(P3_IR_REG_14__SCAN_IN), .Y(n10168));
  AOI21X1 g08455(.A0(n10142), .A1(n10156), .B0(n10168), .Y(n10169));
  INVX1   g08456(.A(n10142), .Y(n10170));
  NOR3X1  g08457(.A(n10170), .B(P3_IR_REG_14__SCAN_IN), .C(P3_IR_REG_13__SCAN_IN), .Y(n10171));
  NOR2X1  g08458(.A(n10171), .B(n10169), .Y(n10172));
  AOI22X1 g08459(.A0(n9983), .A1(n10172), .B0(n9981), .B1(P3_IR_REG_14__SCAN_IN), .Y(n10173));
  OAI21X1 g08460(.A0(n10167), .A1(P3_STATE_REG_SCAN_IN), .B0(n10173), .Y(P3_U3281));
  XOR2X1  g08461(.A(P2_DATAO_REG_15__SCAN_IN), .B(n6177), .Y(n10175));
  NOR2X1  g08462(.A(P2_DATAO_REG_14__SCAN_IN), .B(n2131), .Y(n10176));
  NOR2X1  g08463(.A(n2109), .B(P1_DATAO_REG_14__SCAN_IN), .Y(n10177));
  INVX1   g08464(.A(n10177), .Y(n10178));
  AOI21X1 g08465(.A0(n10165), .A1(n10178), .B0(n10176), .Y(n10179));
  XOR2X1  g08466(.A(n10179), .B(n10175), .Y(n10180));
  NOR2X1  g08467(.A(n10180), .B(n1837), .Y(n10181));
  AOI21X1 g08468(.A0(n1837), .A1(SI_15_), .B0(n10181), .Y(n10182));
  INVX1   g08469(.A(P3_IR_REG_15__SCAN_IN), .Y(n10183));
  XOR2X1  g08470(.A(n10171), .B(n10183), .Y(n10184));
  AOI22X1 g08471(.A0(n9983), .A1(n10184), .B0(n9981), .B1(P3_IR_REG_15__SCAN_IN), .Y(n10185));
  OAI21X1 g08472(.A0(n10182), .A1(P3_STATE_REG_SCAN_IN), .B0(n10185), .Y(P3_U3280));
  NOR3X1  g08473(.A(n1793), .B(n1792), .C(n2183), .Y(n10187));
  XOR2X1  g08474(.A(P2_DATAO_REG_16__SCAN_IN), .B(n6184), .Y(n10188));
  NOR2X1  g08475(.A(P2_DATAO_REG_15__SCAN_IN), .B(n6177), .Y(n10189));
  INVX1   g08476(.A(n10189), .Y(n10190));
  NOR2X1  g08477(.A(n2128), .B(P1_DATAO_REG_15__SCAN_IN), .Y(n10191));
  OAI21X1 g08478(.A0(n10179), .A1(n10191), .B0(n10190), .Y(n10192));
  XOR2X1  g08479(.A(n10192), .B(n10188), .Y(n10193));
  AOI21X1 g08480(.A0(n10193), .A1(n1790), .B0(n10187), .Y(n10194));
  INVX1   g08481(.A(P3_IR_REG_16__SCAN_IN), .Y(n10195));
  NOR4X1  g08482(.A(P3_IR_REG_15__SCAN_IN), .B(P3_IR_REG_14__SCAN_IN), .C(P3_IR_REG_13__SCAN_IN), .D(n10170), .Y(n10196));
  INVX1   g08483(.A(P3_IR_REG_2__SCAN_IN), .Y(n10197));
  NAND4X1 g08484(.A(n10022), .B(n10007), .C(n10197), .D(n10047), .Y(n10198));
  NOR3X1  g08485(.A(P3_IR_REG_12__SCAN_IN), .B(P3_IR_REG_11__SCAN_IN), .C(P3_IR_REG_10__SCAN_IN), .Y(n10199));
  NOR4X1  g08486(.A(P3_IR_REG_15__SCAN_IN), .B(P3_IR_REG_14__SCAN_IN), .C(P3_IR_REG_13__SCAN_IN), .D(P3_IR_REG_16__SCAN_IN), .Y(n10200));
  NOR4X1  g08487(.A(P3_IR_REG_8__SCAN_IN), .B(P3_IR_REG_7__SCAN_IN), .C(P3_IR_REG_6__SCAN_IN), .D(P3_IR_REG_9__SCAN_IN), .Y(n10201));
  NAND3X1 g08488(.A(n10201), .B(n10200), .C(n10199), .Y(n10202));
  NOR3X1  g08489(.A(n10202), .B(n10198), .C(n9997), .Y(n10203));
  INVX1   g08490(.A(n10203), .Y(n10204));
  OAI21X1 g08491(.A0(n10196), .A1(n10195), .B0(n10204), .Y(n10205));
  INVX1   g08492(.A(n10205), .Y(n10206));
  AOI22X1 g08493(.A0(n9983), .A1(n10206), .B0(n9981), .B1(P3_IR_REG_16__SCAN_IN), .Y(n10207));
  OAI21X1 g08494(.A0(n10194), .A1(P3_STATE_REG_SCAN_IN), .B0(n10207), .Y(P3_U3279));
  XOR2X1  g08495(.A(P2_DATAO_REG_17__SCAN_IN), .B(n6201), .Y(n10209));
  NOR2X1  g08496(.A(P2_DATAO_REG_16__SCAN_IN), .B(n6184), .Y(n10210));
  NOR2X1  g08497(.A(n2148), .B(P1_DATAO_REG_16__SCAN_IN), .Y(n10211));
  INVX1   g08498(.A(n10211), .Y(n10212));
  AOI21X1 g08499(.A0(n10192), .A1(n10212), .B0(n10210), .Y(n10213));
  XOR2X1  g08500(.A(n10213), .B(n10209), .Y(n10214));
  NOR2X1  g08501(.A(n10214), .B(n1837), .Y(n10215));
  AOI21X1 g08502(.A0(n1837), .A1(SI_17_), .B0(n10215), .Y(n10216));
  INVX1   g08503(.A(P3_IR_REG_17__SCAN_IN), .Y(n10217));
  XOR2X1  g08504(.A(n10203), .B(n10217), .Y(n10218));
  AOI22X1 g08505(.A0(n9983), .A1(n10218), .B0(n9981), .B1(P3_IR_REG_17__SCAN_IN), .Y(n10219));
  OAI21X1 g08506(.A0(n10216), .A1(P3_STATE_REG_SCAN_IN), .B0(n10219), .Y(P3_U3278));
  NOR3X1  g08507(.A(n1793), .B(n1792), .C(n2229), .Y(n10221));
  XOR2X1  g08508(.A(P2_DATAO_REG_18__SCAN_IN), .B(n6208), .Y(n10222));
  NOR2X1  g08509(.A(P2_DATAO_REG_17__SCAN_IN), .B(n6201), .Y(n10223));
  INVX1   g08510(.A(n10223), .Y(n10224));
  NOR2X1  g08511(.A(n2181), .B(P1_DATAO_REG_17__SCAN_IN), .Y(n10225));
  OAI21X1 g08512(.A0(n10213), .A1(n10225), .B0(n10224), .Y(n10226));
  XOR2X1  g08513(.A(n10226), .B(n10222), .Y(n10227));
  AOI21X1 g08514(.A0(n10227), .A1(n1790), .B0(n10221), .Y(n10228));
  INVX1   g08515(.A(P3_IR_REG_18__SCAN_IN), .Y(n10229));
  NOR4X1  g08516(.A(n10198), .B(n9997), .C(P3_IR_REG_17__SCAN_IN), .D(n10202), .Y(n10230));
  NAND3X1 g08517(.A(n10203), .B(n10229), .C(n10217), .Y(n10231));
  OAI21X1 g08518(.A0(n10230), .A1(n10229), .B0(n10231), .Y(n10232));
  INVX1   g08519(.A(n10232), .Y(n10233));
  AOI22X1 g08520(.A0(n9983), .A1(n10233), .B0(n9981), .B1(P3_IR_REG_18__SCAN_IN), .Y(n10234));
  OAI21X1 g08521(.A0(n10228), .A1(P3_STATE_REG_SCAN_IN), .B0(n10234), .Y(P3_U3277));
  NOR3X1  g08522(.A(n1793), .B(n1792), .C(n2252), .Y(n10236));
  XOR2X1  g08523(.A(P2_DATAO_REG_19__SCAN_IN), .B(n6219), .Y(n10237));
  NOR2X1  g08524(.A(P2_DATAO_REG_18__SCAN_IN), .B(n6208), .Y(n10238));
  NOR2X1  g08525(.A(n2199), .B(P1_DATAO_REG_18__SCAN_IN), .Y(n10239));
  INVX1   g08526(.A(n10239), .Y(n10240));
  AOI21X1 g08527(.A0(n10226), .A1(n10240), .B0(n10238), .Y(n10241));
  XOR2X1  g08528(.A(n10241), .B(n10237), .Y(n10242));
  NOR2X1  g08529(.A(n10242), .B(n1837), .Y(n10243));
  NOR2X1  g08530(.A(n10243), .B(n10236), .Y(n10244));
  XOR2X1  g08531(.A(n10231), .B(P3_IR_REG_19__SCAN_IN), .Y(n10245));
  AOI22X1 g08532(.A0(n9983), .A1(n10245), .B0(n9981), .B1(P3_IR_REG_19__SCAN_IN), .Y(n10246));
  OAI21X1 g08533(.A0(n10244), .A1(P3_STATE_REG_SCAN_IN), .B0(n10246), .Y(P3_U3276));
  NOR3X1  g08534(.A(n1793), .B(n1792), .C(n2276), .Y(n10248));
  XOR2X1  g08535(.A(P2_DATAO_REG_20__SCAN_IN), .B(n6226), .Y(n10249));
  NOR2X1  g08536(.A(P2_DATAO_REG_19__SCAN_IN), .B(n6219), .Y(n10250));
  INVX1   g08537(.A(n10250), .Y(n10251));
  NOR2X1  g08538(.A(n2227), .B(P1_DATAO_REG_19__SCAN_IN), .Y(n10252));
  OAI21X1 g08539(.A0(n10241), .A1(n10252), .B0(n10251), .Y(n10253));
  XOR2X1  g08540(.A(n10253), .B(n10249), .Y(n10254));
  AOI21X1 g08541(.A0(n10254), .A1(n1790), .B0(n10248), .Y(n10255));
  OAI21X1 g08542(.A0(n10231), .A1(P3_IR_REG_19__SCAN_IN), .B0(P3_IR_REG_20__SCAN_IN), .Y(n10256));
  NOR4X1  g08543(.A(P3_IR_REG_19__SCAN_IN), .B(P3_IR_REG_18__SCAN_IN), .C(P3_IR_REG_17__SCAN_IN), .D(P3_IR_REG_20__SCAN_IN), .Y(n10257));
  NAND2X1 g08544(.A(n10257), .B(n10203), .Y(n10258));
  NAND2X1 g08545(.A(n10258), .B(n10256), .Y(n10259));
  NOR3X1  g08546(.A(n10259), .B(n9982), .C(P3_U3151), .Y(n10260));
  AOI21X1 g08547(.A0(n9981), .A1(P3_IR_REG_20__SCAN_IN), .B0(n10260), .Y(n10261));
  OAI21X1 g08548(.A0(n10255), .A1(P3_STATE_REG_SCAN_IN), .B0(n10261), .Y(P3_U3275));
  NOR3X1  g08549(.A(n1793), .B(n1792), .C(n2291), .Y(n10263));
  XOR2X1  g08550(.A(P2_DATAO_REG_21__SCAN_IN), .B(n6234), .Y(n10264));
  NOR2X1  g08551(.A(P2_DATAO_REG_20__SCAN_IN), .B(n6226), .Y(n10265));
  NOR2X1  g08552(.A(n2250), .B(P1_DATAO_REG_20__SCAN_IN), .Y(n10266));
  INVX1   g08553(.A(n10266), .Y(n10267));
  AOI21X1 g08554(.A0(n10253), .A1(n10267), .B0(n10265), .Y(n10268));
  XOR2X1  g08555(.A(n10268), .B(n10264), .Y(n10269));
  NOR2X1  g08556(.A(n10269), .B(n1837), .Y(n10270));
  NOR2X1  g08557(.A(n10270), .B(n10263), .Y(n10271));
  XOR2X1  g08558(.A(n10258), .B(P3_IR_REG_21__SCAN_IN), .Y(n10272));
  AOI22X1 g08559(.A0(n9983), .A1(n10272), .B0(n9981), .B1(P3_IR_REG_21__SCAN_IN), .Y(n10273));
  OAI21X1 g08560(.A0(n10271), .A1(P3_STATE_REG_SCAN_IN), .B0(n10273), .Y(P3_U3274));
  NOR3X1  g08561(.A(n1793), .B(n1792), .C(n2321), .Y(n10275));
  XOR2X1  g08562(.A(P2_DATAO_REG_22__SCAN_IN), .B(n6242), .Y(n10276));
  NOR2X1  g08563(.A(P2_DATAO_REG_21__SCAN_IN), .B(n6234), .Y(n10277));
  INVX1   g08564(.A(n10277), .Y(n10278));
  NOR2X1  g08565(.A(n2274), .B(P1_DATAO_REG_21__SCAN_IN), .Y(n10279));
  OAI21X1 g08566(.A0(n10268), .A1(n10279), .B0(n10278), .Y(n10280));
  XOR2X1  g08567(.A(n10280), .B(n10276), .Y(n10281));
  AOI21X1 g08568(.A0(n10281), .A1(n1790), .B0(n10275), .Y(n10282));
  OAI21X1 g08569(.A0(n10258), .A1(P3_IR_REG_21__SCAN_IN), .B0(P3_IR_REG_22__SCAN_IN), .Y(n10283));
  NOR2X1  g08570(.A(P3_IR_REG_22__SCAN_IN), .B(P3_IR_REG_21__SCAN_IN), .Y(n10284));
  INVX1   g08571(.A(n10284), .Y(n10285));
  OAI21X1 g08572(.A0(n10285), .A1(n10258), .B0(n10283), .Y(n10286));
  NOR3X1  g08573(.A(n10286), .B(n9982), .C(P3_U3151), .Y(n10287));
  AOI21X1 g08574(.A0(n9981), .A1(P3_IR_REG_22__SCAN_IN), .B0(n10287), .Y(n10288));
  OAI21X1 g08575(.A0(n10282), .A1(P3_STATE_REG_SCAN_IN), .B0(n10288), .Y(P3_U3273));
  NOR3X1  g08576(.A(n1793), .B(n1792), .C(n2347), .Y(n10290));
  XOR2X1  g08577(.A(P2_DATAO_REG_23__SCAN_IN), .B(n6250), .Y(n10291));
  NOR2X1  g08578(.A(P2_DATAO_REG_22__SCAN_IN), .B(n6242), .Y(n10292));
  NOR2X1  g08579(.A(n2289), .B(P1_DATAO_REG_22__SCAN_IN), .Y(n10293));
  INVX1   g08580(.A(n10293), .Y(n10294));
  AOI21X1 g08581(.A0(n10280), .A1(n10294), .B0(n10292), .Y(n10295));
  XOR2X1  g08582(.A(n10295), .B(n10291), .Y(n10296));
  NOR2X1  g08583(.A(n10296), .B(n1837), .Y(n10297));
  NOR2X1  g08584(.A(n10297), .B(n10290), .Y(n10298));
  INVX1   g08585(.A(P3_IR_REG_23__SCAN_IN), .Y(n10299));
  NOR2X1  g08586(.A(n10285), .B(n10258), .Y(n10300));
  XOR2X1  g08587(.A(n10300), .B(n10299), .Y(n10301));
  AOI22X1 g08588(.A0(n9983), .A1(n10301), .B0(n9981), .B1(P3_IR_REG_23__SCAN_IN), .Y(n10302));
  OAI21X1 g08589(.A0(n10298), .A1(P3_STATE_REG_SCAN_IN), .B0(n10302), .Y(P3_U3272));
  NOR3X1  g08590(.A(n1793), .B(n1792), .C(n2373), .Y(n10304));
  XOR2X1  g08591(.A(P2_DATAO_REG_24__SCAN_IN), .B(n6259), .Y(n10305));
  NOR2X1  g08592(.A(P2_DATAO_REG_23__SCAN_IN), .B(n6250), .Y(n10306));
  INVX1   g08593(.A(n10306), .Y(n10307));
  NOR2X1  g08594(.A(n2319), .B(P1_DATAO_REG_23__SCAN_IN), .Y(n10308));
  OAI21X1 g08595(.A0(n10295), .A1(n10308), .B0(n10307), .Y(n10309));
  XOR2X1  g08596(.A(n10309), .B(n10305), .Y(n10310));
  AOI21X1 g08597(.A0(n10310), .A1(n1790), .B0(n10304), .Y(n10311));
  NAND4X1 g08598(.A(n10257), .B(n10203), .C(n10299), .D(n10284), .Y(n10312));
  NOR4X1  g08599(.A(P3_IR_REG_23__SCAN_IN), .B(P3_IR_REG_22__SCAN_IN), .C(P3_IR_REG_21__SCAN_IN), .D(P3_IR_REG_24__SCAN_IN), .Y(n10313));
  NAND2X1 g08600(.A(n10313), .B(n10257), .Y(n10314));
  NOR4X1  g08601(.A(n10202), .B(n10198), .C(n9997), .D(n10314), .Y(n10315));
  AOI21X1 g08602(.A0(n10312), .A1(P3_IR_REG_24__SCAN_IN), .B0(n10315), .Y(n10316));
  AOI22X1 g08603(.A0(n9983), .A1(n10316), .B0(n9981), .B1(P3_IR_REG_24__SCAN_IN), .Y(n10317));
  OAI21X1 g08604(.A0(n10311), .A1(P3_STATE_REG_SCAN_IN), .B0(n10317), .Y(P3_U3271));
  NOR3X1  g08605(.A(n1793), .B(n1792), .C(n2391), .Y(n10319));
  XOR2X1  g08606(.A(P2_DATAO_REG_25__SCAN_IN), .B(n6266), .Y(n10320));
  NOR2X1  g08607(.A(P2_DATAO_REG_24__SCAN_IN), .B(n6259), .Y(n10321));
  NOR2X1  g08608(.A(n2345), .B(P1_DATAO_REG_24__SCAN_IN), .Y(n10322));
  INVX1   g08609(.A(n10322), .Y(n10323));
  AOI21X1 g08610(.A0(n10309), .A1(n10323), .B0(n10321), .Y(n10324));
  XOR2X1  g08611(.A(n10324), .B(n10320), .Y(n10325));
  NOR2X1  g08612(.A(n10325), .B(n1837), .Y(n10326));
  NOR2X1  g08613(.A(n10326), .B(n10319), .Y(n10327));
  INVX1   g08614(.A(P3_IR_REG_25__SCAN_IN), .Y(n10328));
  XOR2X1  g08615(.A(n10315), .B(n10328), .Y(n10329));
  AOI22X1 g08616(.A0(n9983), .A1(n10329), .B0(n9981), .B1(P3_IR_REG_25__SCAN_IN), .Y(n10330));
  OAI21X1 g08617(.A0(n10327), .A1(P3_STATE_REG_SCAN_IN), .B0(n10330), .Y(P3_U3270));
  NOR3X1  g08618(.A(n1793), .B(n1792), .C(n2423), .Y(n10332));
  XOR2X1  g08619(.A(P2_DATAO_REG_26__SCAN_IN), .B(n6274), .Y(n10333));
  NOR2X1  g08620(.A(P2_DATAO_REG_25__SCAN_IN), .B(n6266), .Y(n10334));
  INVX1   g08621(.A(n10334), .Y(n10335));
  NOR2X1  g08622(.A(n2371), .B(P1_DATAO_REG_25__SCAN_IN), .Y(n10336));
  OAI21X1 g08623(.A0(n10324), .A1(n10336), .B0(n10335), .Y(n10337));
  XOR2X1  g08624(.A(n10337), .B(n10333), .Y(n10338));
  AOI21X1 g08625(.A0(n10338), .A1(n1790), .B0(n10332), .Y(n10339));
  INVX1   g08626(.A(P3_IR_REG_26__SCAN_IN), .Y(n10340));
  AOI21X1 g08627(.A0(n10315), .A1(n10328), .B0(n10340), .Y(n10341));
  NAND3X1 g08628(.A(n10313), .B(n10257), .C(n10203), .Y(n10342));
  NAND2X1 g08629(.A(n10340), .B(n10328), .Y(n10343));
  NOR2X1  g08630(.A(n10343), .B(n10342), .Y(n10344));
  NOR2X1  g08631(.A(n10344), .B(n10341), .Y(n10345));
  AOI22X1 g08632(.A0(n9983), .A1(n10345), .B0(n9981), .B1(P3_IR_REG_26__SCAN_IN), .Y(n10346));
  OAI21X1 g08633(.A0(n10339), .A1(P3_STATE_REG_SCAN_IN), .B0(n10346), .Y(P3_U3269));
  NOR3X1  g08634(.A(n1793), .B(n1792), .C(n2443), .Y(n10348));
  XOR2X1  g08635(.A(P2_DATAO_REG_27__SCAN_IN), .B(n6295), .Y(n10349));
  NOR2X1  g08636(.A(P2_DATAO_REG_26__SCAN_IN), .B(n6274), .Y(n10350));
  NOR2X1  g08637(.A(n2389), .B(P1_DATAO_REG_26__SCAN_IN), .Y(n10351));
  INVX1   g08638(.A(n10351), .Y(n10352));
  AOI21X1 g08639(.A0(n10337), .A1(n10352), .B0(n10350), .Y(n10353));
  XOR2X1  g08640(.A(n10353), .B(n10349), .Y(n10354));
  NOR2X1  g08641(.A(n10354), .B(n1837), .Y(n10355));
  NOR2X1  g08642(.A(n10355), .B(n10348), .Y(n10356));
  INVX1   g08643(.A(P3_IR_REG_27__SCAN_IN), .Y(n10357));
  XOR2X1  g08644(.A(n10344), .B(n10357), .Y(n10358));
  AOI22X1 g08645(.A0(n9983), .A1(n10358), .B0(n9981), .B1(P3_IR_REG_27__SCAN_IN), .Y(n10359));
  OAI21X1 g08646(.A0(n10356), .A1(P3_STATE_REG_SCAN_IN), .B0(n10359), .Y(P3_U3268));
  NOR3X1  g08647(.A(n1793), .B(n1792), .C(n2468), .Y(n10361));
  NOR2X1  g08648(.A(P2_DATAO_REG_27__SCAN_IN), .B(n6295), .Y(n10362));
  XOR2X1  g08649(.A(P2_DATAO_REG_28__SCAN_IN), .B(n6302), .Y(n10363));
  INVX1   g08650(.A(n10363), .Y(n10364));
  AOI21X1 g08651(.A0(P2_DATAO_REG_27__SCAN_IN), .A1(n6295), .B0(n10353), .Y(n10365));
  OAI21X1 g08652(.A0(n10365), .A1(n10362), .B0(n10364), .Y(n10366));
  INVX1   g08653(.A(n10362), .Y(n10367));
  NAND3X1 g08654(.A(n10070), .B(n10090), .C(n10034), .Y(n10368));
  INVX1   g08655(.A(n10149), .Y(n10369));
  AOI21X1 g08656(.A0(n10093), .A1(n10368), .B0(n10369), .Y(n10370));
  OAI22X1 g08657(.A0(n10370), .A1(n10151), .B0(n2088), .B1(P1_DATAO_REG_13__SCAN_IN), .Y(n10371));
  AOI21X1 g08658(.A0(n10371), .A1(n10163), .B0(n10177), .Y(n10372));
  OAI22X1 g08659(.A0(n10176), .A1(n10372), .B0(n2128), .B1(P1_DATAO_REG_15__SCAN_IN), .Y(n10373));
  AOI21X1 g08660(.A0(n10373), .A1(n10190), .B0(n10211), .Y(n10374));
  OAI22X1 g08661(.A0(n10210), .A1(n10374), .B0(n2181), .B1(P1_DATAO_REG_17__SCAN_IN), .Y(n10375));
  AOI21X1 g08662(.A0(n10375), .A1(n10224), .B0(n10239), .Y(n10376));
  OAI22X1 g08663(.A0(n10238), .A1(n10376), .B0(n2227), .B1(P1_DATAO_REG_19__SCAN_IN), .Y(n10377));
  AOI21X1 g08664(.A0(n10377), .A1(n10251), .B0(n10266), .Y(n10378));
  OAI22X1 g08665(.A0(n10265), .A1(n10378), .B0(n2274), .B1(P1_DATAO_REG_21__SCAN_IN), .Y(n10379));
  AOI21X1 g08666(.A0(n10379), .A1(n10278), .B0(n10293), .Y(n10380));
  OAI22X1 g08667(.A0(n10292), .A1(n10380), .B0(n2319), .B1(P1_DATAO_REG_23__SCAN_IN), .Y(n10381));
  AOI21X1 g08668(.A0(n10381), .A1(n10307), .B0(n10322), .Y(n10382));
  OAI22X1 g08669(.A0(n10321), .A1(n10382), .B0(n2371), .B1(P1_DATAO_REG_25__SCAN_IN), .Y(n10383));
  AOI21X1 g08670(.A0(n10383), .A1(n10335), .B0(n10351), .Y(n10384));
  OAI22X1 g08671(.A0(n10350), .A1(n10384), .B0(n2421), .B1(P1_DATAO_REG_27__SCAN_IN), .Y(n10385));
  NAND3X1 g08672(.A(n10385), .B(n10363), .C(n10367), .Y(n10386));
  AOI21X1 g08673(.A0(n10386), .A1(n10366), .B0(n1837), .Y(n10387));
  OAI21X1 g08674(.A0(n10387), .A1(n10361), .B0(P3_U3151), .Y(n10388));
  OAI21X1 g08675(.A0(n10343), .A1(n10342), .B0(P3_IR_REG_28__SCAN_IN), .Y(n10389));
  NOR4X1  g08676(.A(n10342), .B(P3_IR_REG_28__SCAN_IN), .C(P3_IR_REG_27__SCAN_IN), .D(n10343), .Y(n10390));
  AOI21X1 g08677(.A0(P3_IR_REG_28__SCAN_IN), .A1(P3_IR_REG_27__SCAN_IN), .B0(n10390), .Y(n10391));
  NAND2X1 g08678(.A(n10391), .B(n10389), .Y(n10392));
  NOR3X1  g08679(.A(n10392), .B(n9982), .C(P3_U3151), .Y(n10393));
  AOI21X1 g08680(.A0(n9981), .A1(P3_IR_REG_28__SCAN_IN), .B0(n10393), .Y(n10394));
  NAND2X1 g08681(.A(n10394), .B(n10388), .Y(P3_U3267));
  NOR3X1  g08682(.A(n1793), .B(n1792), .C(n2495), .Y(n10396));
  NOR2X1  g08683(.A(P2_DATAO_REG_28__SCAN_IN), .B(n6302), .Y(n10397));
  XOR2X1  g08684(.A(P2_DATAO_REG_29__SCAN_IN), .B(n6312), .Y(n10398));
  INVX1   g08685(.A(n10398), .Y(n10399));
  AOI22X1 g08686(.A0(n10367), .A1(n10385), .B0(P2_DATAO_REG_28__SCAN_IN), .B1(n6302), .Y(n10400));
  OAI21X1 g08687(.A0(n10400), .A1(n10397), .B0(n10399), .Y(n10401));
  INVX1   g08688(.A(n10397), .Y(n10402));
  OAI22X1 g08689(.A0(n10362), .A1(n10365), .B0(n2441), .B1(P1_DATAO_REG_28__SCAN_IN), .Y(n10403));
  NAND3X1 g08690(.A(n10403), .B(n10398), .C(n10402), .Y(n10404));
  AOI21X1 g08691(.A0(n10404), .A1(n10401), .B0(n1837), .Y(n10405));
  OAI21X1 g08692(.A0(n10405), .A1(n10396), .B0(P3_U3151), .Y(n10406));
  INVX1   g08693(.A(P3_IR_REG_29__SCAN_IN), .Y(n10407));
  XOR2X1  g08694(.A(n10390), .B(n10407), .Y(n10408));
  AOI22X1 g08695(.A0(n9983), .A1(n10408), .B0(n9981), .B1(P3_IR_REG_29__SCAN_IN), .Y(n10409));
  NAND2X1 g08696(.A(n10409), .B(n10406), .Y(P3_U3266));
  NOR3X1  g08697(.A(n1793), .B(n1792), .C(n2513), .Y(n10411));
  NOR2X1  g08698(.A(P2_DATAO_REG_29__SCAN_IN), .B(n6312), .Y(n10412));
  XOR2X1  g08699(.A(P2_DATAO_REG_30__SCAN_IN), .B(n5116), .Y(n10413));
  INVX1   g08700(.A(n10413), .Y(n10414));
  AOI22X1 g08701(.A0(n10402), .A1(n10403), .B0(P2_DATAO_REG_29__SCAN_IN), .B1(n6312), .Y(n10415));
  OAI21X1 g08702(.A0(n10415), .A1(n10412), .B0(n10414), .Y(n10416));
  INVX1   g08703(.A(n10412), .Y(n10417));
  OAI22X1 g08704(.A0(n10397), .A1(n10400), .B0(n2466), .B1(P1_DATAO_REG_29__SCAN_IN), .Y(n10418));
  NAND3X1 g08705(.A(n10418), .B(n10413), .C(n10417), .Y(n10419));
  AOI21X1 g08706(.A0(n10419), .A1(n10416), .B0(n1837), .Y(n10420));
  OAI21X1 g08707(.A0(n10420), .A1(n10411), .B0(P3_U3151), .Y(n10421));
  NAND2X1 g08708(.A(n10390), .B(n10407), .Y(n10422));
  XOR2X1  g08709(.A(n10422), .B(P3_IR_REG_30__SCAN_IN), .Y(n10423));
  AOI22X1 g08710(.A0(n9983), .A1(n10423), .B0(n9981), .B1(P3_IR_REG_30__SCAN_IN), .Y(n10424));
  NAND2X1 g08711(.A(n10424), .B(n10421), .Y(P3_U3265));
  NAND3X1 g08712(.A(n1789), .B(n1786), .C(SI_31_), .Y(n10426));
  INVX1   g08713(.A(n10426), .Y(n10427));
  XOR2X1  g08714(.A(P2_DATAO_REG_31__SCAN_IN), .B(n5121), .Y(n10428));
  AOI21X1 g08715(.A0(P2_DATAO_REG_30__SCAN_IN), .A1(n5116), .B0(n10428), .Y(n10429));
  OAI21X1 g08716(.A0(n10415), .A1(n10412), .B0(n10429), .Y(n10430));
  NOR2X1  g08717(.A(P2_DATAO_REG_30__SCAN_IN), .B(n5116), .Y(n10431));
  INVX1   g08718(.A(n10428), .Y(n10432));
  NOR3X1  g08719(.A(n10432), .B(n10431), .C(n10412), .Y(n10433));
  NOR3X1  g08720(.A(n10432), .B(n2492), .C(P1_DATAO_REG_30__SCAN_IN), .Y(n10434));
  AOI21X1 g08721(.A0(n10432), .A1(n10431), .B0(n10434), .Y(n10435));
  INVX1   g08722(.A(n10435), .Y(n10436));
  AOI21X1 g08723(.A0(n10433), .A1(n10418), .B0(n10436), .Y(n10437));
  AOI21X1 g08724(.A0(n10437), .A1(n10430), .B0(n1837), .Y(n10438));
  OAI21X1 g08725(.A0(n10438), .A1(n10427), .B0(P3_U3151), .Y(n10439));
  NOR2X1  g08726(.A(n10422), .B(P3_IR_REG_30__SCAN_IN), .Y(n10440));
  NAND3X1 g08727(.A(n10440), .B(P3_IR_REG_31__SCAN_IN), .C(P3_STATE_REG_SCAN_IN), .Y(n10441));
  NAND2X1 g08728(.A(n10441), .B(n10439), .Y(P3_U3264));
  INVX1   g08729(.A(P3_D_REG_0__SCAN_IN), .Y(n10443));
  NOR2X1  g08730(.A(P3_IR_REG_31__SCAN_IN), .B(n10299), .Y(n10444));
  AOI21X1 g08731(.A0(n10301), .A1(P3_IR_REG_31__SCAN_IN), .B0(n10444), .Y(n10445));
  INVX1   g08732(.A(n10445), .Y(n10446));
  NAND2X1 g08733(.A(n9982), .B(P3_IR_REG_24__SCAN_IN), .Y(n10447));
  INVX1   g08734(.A(n10447), .Y(n10448));
  AOI21X1 g08735(.A0(n10316), .A1(P3_IR_REG_31__SCAN_IN), .B0(n10448), .Y(n10449));
  NOR2X1  g08736(.A(P3_IR_REG_31__SCAN_IN), .B(n10328), .Y(n10450));
  AOI21X1 g08737(.A0(n10329), .A1(P3_IR_REG_31__SCAN_IN), .B0(n10450), .Y(n10451));
  NOR2X1  g08738(.A(P3_IR_REG_31__SCAN_IN), .B(n10340), .Y(n10452));
  AOI21X1 g08739(.A0(n10345), .A1(P3_IR_REG_31__SCAN_IN), .B0(n10452), .Y(n10453));
  NOR3X1  g08740(.A(n10453), .B(n10451), .C(n10449), .Y(n10454));
  INVX1   g08741(.A(P3_B_REG_SCAN_IN), .Y(n10455));
  XOR2X1  g08742(.A(n10449), .B(n10455), .Y(n10456));
  AOI21X1 g08743(.A0(n10456), .A1(n10451), .B0(n10453), .Y(n10457));
  NOR4X1  g08744(.A(n10454), .B(n10446), .C(P3_U3151), .D(n10457), .Y(n10458));
  INVX1   g08745(.A(n10451), .Y(n10459));
  OAI21X1 g08746(.A0(n10453), .A1(n10459), .B0(n10449), .Y(n10460));
  NAND2X1 g08747(.A(n10460), .B(n10458), .Y(n10461));
  OAI21X1 g08748(.A0(n10458), .A1(n10443), .B0(n10461), .Y(P3_U3376));
  INVX1   g08749(.A(P3_D_REG_1__SCAN_IN), .Y(n10463));
  INVX1   g08750(.A(n10453), .Y(n10464));
  OAI21X1 g08751(.A0(n10464), .A1(n10459), .B0(n10458), .Y(n10465));
  OAI21X1 g08752(.A0(n10458), .A1(n10463), .B0(n10465), .Y(P3_U3377));
  INVX1   g08753(.A(P3_D_REG_2__SCAN_IN), .Y(n10467));
  NOR2X1  g08754(.A(n10458), .B(n10467), .Y(P3_U3263));
  INVX1   g08755(.A(P3_D_REG_3__SCAN_IN), .Y(n10469));
  NOR2X1  g08756(.A(n10458), .B(n10469), .Y(P3_U3262));
  INVX1   g08757(.A(P3_D_REG_4__SCAN_IN), .Y(n10471));
  NOR2X1  g08758(.A(n10458), .B(n10471), .Y(P3_U3261));
  INVX1   g08759(.A(P3_D_REG_5__SCAN_IN), .Y(n10473));
  NOR2X1  g08760(.A(n10458), .B(n10473), .Y(P3_U3260));
  INVX1   g08761(.A(P3_D_REG_6__SCAN_IN), .Y(n10475));
  NOR2X1  g08762(.A(n10458), .B(n10475), .Y(P3_U3259));
  INVX1   g08763(.A(P3_D_REG_7__SCAN_IN), .Y(n10477));
  NOR2X1  g08764(.A(n10458), .B(n10477), .Y(P3_U3258));
  INVX1   g08765(.A(P3_D_REG_8__SCAN_IN), .Y(n10479));
  NOR2X1  g08766(.A(n10458), .B(n10479), .Y(P3_U3257));
  INVX1   g08767(.A(P3_D_REG_9__SCAN_IN), .Y(n10481));
  NOR2X1  g08768(.A(n10458), .B(n10481), .Y(P3_U3256));
  INVX1   g08769(.A(P3_D_REG_10__SCAN_IN), .Y(n10483));
  NOR2X1  g08770(.A(n10458), .B(n10483), .Y(P3_U3255));
  INVX1   g08771(.A(P3_D_REG_11__SCAN_IN), .Y(n10485));
  NOR2X1  g08772(.A(n10458), .B(n10485), .Y(P3_U3254));
  INVX1   g08773(.A(P3_D_REG_12__SCAN_IN), .Y(n10487));
  NOR2X1  g08774(.A(n10458), .B(n10487), .Y(P3_U3253));
  INVX1   g08775(.A(P3_D_REG_13__SCAN_IN), .Y(n10489));
  NOR2X1  g08776(.A(n10458), .B(n10489), .Y(P3_U3252));
  INVX1   g08777(.A(P3_D_REG_14__SCAN_IN), .Y(n10491));
  NOR2X1  g08778(.A(n10458), .B(n10491), .Y(P3_U3251));
  INVX1   g08779(.A(P3_D_REG_15__SCAN_IN), .Y(n10493));
  NOR2X1  g08780(.A(n10458), .B(n10493), .Y(P3_U3250));
  INVX1   g08781(.A(P3_D_REG_16__SCAN_IN), .Y(n10495));
  NOR2X1  g08782(.A(n10458), .B(n10495), .Y(P3_U3249));
  INVX1   g08783(.A(P3_D_REG_17__SCAN_IN), .Y(n10497));
  NOR2X1  g08784(.A(n10458), .B(n10497), .Y(P3_U3248));
  INVX1   g08785(.A(P3_D_REG_18__SCAN_IN), .Y(n10499));
  NOR2X1  g08786(.A(n10458), .B(n10499), .Y(P3_U3247));
  INVX1   g08787(.A(P3_D_REG_19__SCAN_IN), .Y(n10501));
  NOR2X1  g08788(.A(n10458), .B(n10501), .Y(P3_U3246));
  INVX1   g08789(.A(P3_D_REG_20__SCAN_IN), .Y(n10503));
  NOR2X1  g08790(.A(n10458), .B(n10503), .Y(P3_U3245));
  INVX1   g08791(.A(P3_D_REG_21__SCAN_IN), .Y(n10505));
  NOR2X1  g08792(.A(n10458), .B(n10505), .Y(P3_U3244));
  INVX1   g08793(.A(P3_D_REG_22__SCAN_IN), .Y(n10507));
  NOR2X1  g08794(.A(n10458), .B(n10507), .Y(P3_U3243));
  INVX1   g08795(.A(P3_D_REG_23__SCAN_IN), .Y(n10509));
  NOR2X1  g08796(.A(n10458), .B(n10509), .Y(P3_U3242));
  INVX1   g08797(.A(P3_D_REG_24__SCAN_IN), .Y(n10511));
  NOR2X1  g08798(.A(n10458), .B(n10511), .Y(P3_U3241));
  INVX1   g08799(.A(P3_D_REG_25__SCAN_IN), .Y(n10513));
  NOR2X1  g08800(.A(n10458), .B(n10513), .Y(P3_U3240));
  INVX1   g08801(.A(P3_D_REG_26__SCAN_IN), .Y(n10515));
  NOR2X1  g08802(.A(n10458), .B(n10515), .Y(P3_U3239));
  INVX1   g08803(.A(P3_D_REG_27__SCAN_IN), .Y(n10517));
  NOR2X1  g08804(.A(n10458), .B(n10517), .Y(P3_U3238));
  INVX1   g08805(.A(P3_D_REG_28__SCAN_IN), .Y(n10519));
  NOR2X1  g08806(.A(n10458), .B(n10519), .Y(P3_U3237));
  INVX1   g08807(.A(P3_D_REG_29__SCAN_IN), .Y(n10521));
  NOR2X1  g08808(.A(n10458), .B(n10521), .Y(P3_U3236));
  INVX1   g08809(.A(P3_D_REG_30__SCAN_IN), .Y(n10523));
  NOR2X1  g08810(.A(n10458), .B(n10523), .Y(P3_U3235));
  INVX1   g08811(.A(P3_D_REG_31__SCAN_IN), .Y(n10525));
  NOR2X1  g08812(.A(n10458), .B(n10525), .Y(P3_U3234));
  INVX1   g08813(.A(P3_REG0_REG_0__SCAN_IN), .Y(n10527));
  NOR3X1  g08814(.A(n10454), .B(n10446), .C(P3_U3151), .Y(n10528));
  INVX1   g08815(.A(n10528), .Y(n10529));
  OAI21X1 g08816(.A0(P3_D_REG_7__SCAN_IN), .A1(P3_D_REG_3__SCAN_IN), .B0(n10457), .Y(n10530));
  OAI21X1 g08817(.A0(P3_D_REG_9__SCAN_IN), .A1(P3_D_REG_8__SCAN_IN), .B0(n10457), .Y(n10531));
  OAI21X1 g08818(.A0(P3_D_REG_10__SCAN_IN), .A1(P3_D_REG_5__SCAN_IN), .B0(n10457), .Y(n10532));
  OAI21X1 g08819(.A0(P3_D_REG_6__SCAN_IN), .A1(P3_D_REG_4__SCAN_IN), .B0(n10457), .Y(n10533));
  NAND4X1 g08820(.A(n10532), .B(n10531), .C(n10530), .D(n10533), .Y(n10534));
  OAI21X1 g08821(.A0(P3_D_REG_28__SCAN_IN), .A1(P3_D_REG_27__SCAN_IN), .B0(n10457), .Y(n10535));
  OAI21X1 g08822(.A0(P3_D_REG_26__SCAN_IN), .A1(P3_D_REG_25__SCAN_IN), .B0(n10457), .Y(n10536));
  OAI21X1 g08823(.A0(P3_D_REG_31__SCAN_IN), .A1(P3_D_REG_30__SCAN_IN), .B0(n10457), .Y(n10537));
  OAI21X1 g08824(.A0(P3_D_REG_29__SCAN_IN), .A1(P3_D_REG_2__SCAN_IN), .B0(n10457), .Y(n10538));
  NAND4X1 g08825(.A(n10537), .B(n10536), .C(n10535), .D(n10538), .Y(n10539));
  OAI21X1 g08826(.A0(P3_D_REG_21__SCAN_IN), .A1(P3_D_REG_20__SCAN_IN), .B0(n10457), .Y(n10540));
  OAI21X1 g08827(.A0(P3_D_REG_19__SCAN_IN), .A1(P3_D_REG_18__SCAN_IN), .B0(n10457), .Y(n10541));
  OAI21X1 g08828(.A0(P3_D_REG_23__SCAN_IN), .A1(P3_D_REG_22__SCAN_IN), .B0(n10457), .Y(n10542));
  NAND3X1 g08829(.A(n10542), .B(n10541), .C(n10540), .Y(n10543));
  OAI21X1 g08830(.A0(P3_D_REG_14__SCAN_IN), .A1(P3_D_REG_12__SCAN_IN), .B0(n10457), .Y(n10544));
  OAI21X1 g08831(.A0(P3_D_REG_13__SCAN_IN), .A1(P3_D_REG_11__SCAN_IN), .B0(n10457), .Y(n10545));
  OAI21X1 g08832(.A0(P3_D_REG_24__SCAN_IN), .A1(P3_D_REG_16__SCAN_IN), .B0(n10457), .Y(n10546));
  OAI21X1 g08833(.A0(P3_D_REG_17__SCAN_IN), .A1(P3_D_REG_15__SCAN_IN), .B0(n10457), .Y(n10547));
  NAND4X1 g08834(.A(n10546), .B(n10545), .C(n10544), .D(n10547), .Y(n10548));
  NOR4X1  g08835(.A(n10543), .B(n10539), .C(n10534), .D(n10548), .Y(n10549));
  INVX1   g08836(.A(n10549), .Y(n10550));
  AOI21X1 g08837(.A0(n10453), .A1(n10451), .B0(n10457), .Y(n10551));
  AOI21X1 g08838(.A0(n10457), .A1(P3_D_REG_1__SCAN_IN), .B0(n10551), .Y(n10552));
  INVX1   g08839(.A(n10552), .Y(n10553));
  NAND2X1 g08840(.A(n10457), .B(P3_D_REG_0__SCAN_IN), .Y(n10554));
  INVX1   g08841(.A(n10449), .Y(n10555));
  NOR2X1  g08842(.A(n10464), .B(n10555), .Y(n10556));
  OAI21X1 g08843(.A0(n10556), .A1(n10457), .B0(n10554), .Y(n10557));
  INVX1   g08844(.A(P3_IR_REG_21__SCAN_IN), .Y(n10558));
  NOR2X1  g08845(.A(P3_IR_REG_31__SCAN_IN), .B(n10558), .Y(n10559));
  AOI21X1 g08846(.A0(n10272), .A1(P3_IR_REG_31__SCAN_IN), .B0(n10559), .Y(n10560));
  NAND2X1 g08847(.A(n9982), .B(P3_IR_REG_22__SCAN_IN), .Y(n10561));
  OAI21X1 g08848(.A0(n10286), .A1(n9982), .B0(n10561), .Y(n10562));
  INVX1   g08849(.A(n10562), .Y(n10563));
  INVX1   g08850(.A(n10560), .Y(n10564));
  NAND2X1 g08851(.A(n9982), .B(P3_IR_REG_20__SCAN_IN), .Y(n10565));
  OAI21X1 g08852(.A0(n10259), .A1(n9982), .B0(n10565), .Y(n10566));
  NOR2X1  g08853(.A(n10566), .B(n10564), .Y(n10567));
  XOR2X1  g08854(.A(n10567), .B(n10563), .Y(n10568));
  NAND2X1 g08855(.A(n9982), .B(P3_IR_REG_19__SCAN_IN), .Y(n10569));
  INVX1   g08856(.A(n10569), .Y(n10570));
  AOI21X1 g08857(.A0(n10245), .A1(P3_IR_REG_31__SCAN_IN), .B0(n10570), .Y(n10571));
  AOI21X1 g08858(.A0(n10571), .A1(n10560), .B0(n10568), .Y(n10572));
  NOR4X1  g08859(.A(n10557), .B(n10553), .C(n10550), .D(n10572), .Y(n10573));
  INVX1   g08860(.A(n10573), .Y(n10574));
  INVX1   g08861(.A(n10566), .Y(n10575));
  INVX1   g08862(.A(n10571), .Y(n10576));
  NAND2X1 g08863(.A(n10576), .B(n10562), .Y(n10577));
  NOR2X1  g08864(.A(n10577), .B(n10564), .Y(n10578));
  INVX1   g08865(.A(n10578), .Y(n10579));
  NAND2X1 g08866(.A(n10571), .B(n10562), .Y(n10580));
  NOR3X1  g08867(.A(n10580), .B(n10566), .C(n10560), .Y(n10581));
  INVX1   g08868(.A(n10581), .Y(n10582));
  OAI21X1 g08869(.A0(n10579), .A1(n10575), .B0(n10582), .Y(n10583));
  NAND4X1 g08870(.A(n10557), .B(n10553), .C(n10549), .D(n10583), .Y(n10584));
  AOI21X1 g08871(.A0(n10584), .A1(n10574), .B0(n10529), .Y(n10585));
  NAND2X1 g08872(.A(n10358), .B(P3_IR_REG_31__SCAN_IN), .Y(n10586));
  OAI21X1 g08873(.A0(P3_IR_REG_31__SCAN_IN), .A1(n10357), .B0(n10586), .Y(n10587));
  NAND2X1 g08874(.A(n9982), .B(P3_IR_REG_28__SCAN_IN), .Y(n10588));
  OAI21X1 g08875(.A0(n10392), .A1(n9982), .B0(n10588), .Y(n10589));
  NOR2X1  g08876(.A(n10589), .B(n10587), .Y(n10590));
  NAND2X1 g08877(.A(P3_IR_REG_31__SCAN_IN), .B(P3_IR_REG_0__SCAN_IN), .Y(n10591));
  NAND2X1 g08878(.A(n9982), .B(P3_IR_REG_0__SCAN_IN), .Y(n10592));
  NAND2X1 g08879(.A(n10592), .B(n10591), .Y(n10593));
  NAND2X1 g08880(.A(n10593), .B(n10590), .Y(n10594));
  OAI21X1 g08881(.A0(n10590), .A1(n9972), .B0(n10594), .Y(n10595));
  INVX1   g08882(.A(P3_REG2_REG_0__SCAN_IN), .Y(n10596));
  INVX1   g08883(.A(P3_IR_REG_30__SCAN_IN), .Y(n10597));
  NOR2X1  g08884(.A(P3_IR_REG_31__SCAN_IN), .B(n10597), .Y(n10598));
  AOI21X1 g08885(.A0(n10423), .A1(P3_IR_REG_31__SCAN_IN), .B0(n10598), .Y(n10599));
  NOR2X1  g08886(.A(P3_IR_REG_31__SCAN_IN), .B(n10407), .Y(n10600));
  AOI21X1 g08887(.A0(n10408), .A1(P3_IR_REG_31__SCAN_IN), .B0(n10600), .Y(n10601));
  NAND2X1 g08888(.A(n10601), .B(n10599), .Y(n10602));
  XOR2X1  g08889(.A(n10422), .B(n10597), .Y(n10603));
  INVX1   g08890(.A(n10598), .Y(n10604));
  OAI21X1 g08891(.A0(n10603), .A1(n9982), .B0(n10604), .Y(n10605));
  NAND2X1 g08892(.A(n10601), .B(n10605), .Y(n10606));
  OAI22X1 g08893(.A0(n10602), .A1(n10527), .B0(n10596), .B1(n10606), .Y(n10607));
  INVX1   g08894(.A(P3_REG3_REG_0__SCAN_IN), .Y(n10608));
  INVX1   g08895(.A(P3_REG1_REG_0__SCAN_IN), .Y(n10609));
  NAND2X1 g08896(.A(n10408), .B(P3_IR_REG_31__SCAN_IN), .Y(n10610));
  OAI21X1 g08897(.A0(P3_IR_REG_31__SCAN_IN), .A1(n10407), .B0(n10610), .Y(n10611));
  NAND2X1 g08898(.A(n10611), .B(n10599), .Y(n10612));
  NAND2X1 g08899(.A(n10611), .B(n10605), .Y(n10613));
  OAI22X1 g08900(.A0(n10612), .A1(n10609), .B0(n10608), .B1(n10613), .Y(n10614));
  NOR2X1  g08901(.A(n10614), .B(n10607), .Y(n10615));
  XOR2X1  g08902(.A(n10615), .B(n10595), .Y(n10616));
  NOR2X1  g08903(.A(n10577), .B(n10566), .Y(n10617));
  INVX1   g08904(.A(n10617), .Y(n10618));
  NOR2X1  g08905(.A(n10618), .B(n10616), .Y(n10619));
  INVX1   g08906(.A(n10619), .Y(n10620));
  NOR3X1  g08907(.A(n10571), .B(n10575), .C(n10560), .Y(n10622));
  NOR2X1  g08908(.A(n10580), .B(n10575), .Y(n10623));
  OAI21X1 g08909(.A0(n10623), .A1(n10622), .B0(n13412), .Y(n10624));
  NOR2X1  g08910(.A(n10577), .B(n10575), .Y(n10625));
  NOR3X1  g08911(.A(n10576), .B(n10575), .C(n10560), .Y(n10626));
  OAI21X1 g08912(.A0(n10626), .A1(n10625), .B0(n13412), .Y(n10627));
  NOR4X1  g08913(.A(n10566), .B(n10560), .C(n10562), .D(n10576), .Y(n10628));
  NOR3X1  g08914(.A(n10580), .B(n10566), .C(n10564), .Y(n10629));
  OAI21X1 g08915(.A0(n10629), .A1(n10628), .B0(n13412), .Y(n10630));
  NAND4X1 g08916(.A(n10627), .B(n10624), .C(n10620), .D(n10630), .Y(n10631));
  INVX1   g08917(.A(n10631), .Y(n10632));
  NOR3X1  g08918(.A(n10571), .B(n10566), .C(n10562), .Y(n10633));
  NOR2X1  g08919(.A(n10590), .B(n9972), .Y(n10634));
  AOI21X1 g08920(.A0(n10593), .A1(n10590), .B0(n10634), .Y(n10635));
  XOR2X1  g08921(.A(n10589), .B(n10587), .Y(n10636));
  NOR3X1  g08922(.A(n10636), .B(n10560), .C(n10563), .Y(n10637));
  INVX1   g08923(.A(n10637), .Y(n10638));
  INVX1   g08924(.A(P3_REG0_REG_1__SCAN_IN), .Y(n10639));
  INVX1   g08925(.A(P3_REG2_REG_1__SCAN_IN), .Y(n10640));
  OAI22X1 g08926(.A0(n10602), .A1(n10639), .B0(n10640), .B1(n10606), .Y(n10641));
  INVX1   g08927(.A(P3_REG3_REG_1__SCAN_IN), .Y(n10642));
  INVX1   g08928(.A(P3_REG1_REG_1__SCAN_IN), .Y(n10643));
  OAI22X1 g08929(.A0(n10612), .A1(n10643), .B0(n10642), .B1(n10613), .Y(n10644));
  NOR2X1  g08930(.A(n10644), .B(n10641), .Y(n10645));
  NAND2X1 g08931(.A(n10560), .B(n10563), .Y(n10646));
  OAI22X1 g08932(.A0(n10645), .A1(n10638), .B0(n10635), .B1(n10646), .Y(n10647));
  AOI21X1 g08933(.A0(n10633), .A1(n13412), .B0(n10647), .Y(n10648));
  NAND2X1 g08934(.A(n10648), .B(n10632), .Y(n10649));
  NAND2X1 g08935(.A(n10649), .B(n10585), .Y(n10650));
  OAI21X1 g08936(.A0(n10585), .A1(n10527), .B0(n10650), .Y(P3_U3390));
  NOR2X1  g08937(.A(n10611), .B(n10605), .Y(n10652));
  NOR2X1  g08938(.A(n10611), .B(n10599), .Y(n10653));
  AOI22X1 g08939(.A0(n10652), .A1(P3_REG0_REG_0__SCAN_IN), .B0(P3_REG2_REG_0__SCAN_IN), .B1(n10653), .Y(n10654));
  NOR2X1  g08940(.A(n10601), .B(n10605), .Y(n10655));
  NOR2X1  g08941(.A(n10601), .B(n10599), .Y(n10656));
  AOI22X1 g08942(.A0(n10655), .A1(P3_REG1_REG_0__SCAN_IN), .B0(P3_REG3_REG_0__SCAN_IN), .B1(n10656), .Y(n10657));
  NAND2X1 g08943(.A(n10657), .B(n10654), .Y(n10658));
  NOR2X1  g08944(.A(n10658), .B(n10635), .Y(n10659));
  AOI22X1 g08945(.A0(n10652), .A1(P3_REG0_REG_1__SCAN_IN), .B0(P3_REG2_REG_1__SCAN_IN), .B1(n10653), .Y(n10660));
  AOI22X1 g08946(.A0(n10655), .A1(P3_REG1_REG_1__SCAN_IN), .B0(P3_REG3_REG_1__SCAN_IN), .B1(n10656), .Y(n10661));
  NAND2X1 g08947(.A(n10661), .B(n10660), .Y(n10662));
  NOR2X1  g08948(.A(P3_IR_REG_31__SCAN_IN), .B(n9996), .Y(n10663));
  AOI21X1 g08949(.A0(n9986), .A1(P3_IR_REG_31__SCAN_IN), .B0(n10663), .Y(n10664));
  INVX1   g08950(.A(n10664), .Y(n10665));
  NOR2X1  g08951(.A(n10590), .B(n9979), .Y(n10666));
  AOI21X1 g08952(.A0(n10665), .A1(n10590), .B0(n10666), .Y(n10667));
  XOR2X1  g08953(.A(n10667), .B(n10662), .Y(n10668));
  XOR2X1  g08954(.A(n10668), .B(n10659), .Y(n10669));
  INVX1   g08955(.A(n10669), .Y(n10670));
  OAI21X1 g08956(.A0(n10629), .A1(n10623), .B0(n10670), .Y(n10671));
  XOR2X1  g08957(.A(n10667), .B(n10645), .Y(n10672));
  NOR2X1  g08958(.A(n10615), .B(n10635), .Y(n10673));
  INVX1   g08959(.A(n10673), .Y(n10674));
  XOR2X1  g08960(.A(n10674), .B(n10672), .Y(n10675));
  INVX1   g08961(.A(n10675), .Y(n10676));
  AOI22X1 g08962(.A0(n10670), .A1(n10628), .B0(n10622), .B1(n10676), .Y(n10677));
  INVX1   g08963(.A(n10587), .Y(n10678));
  XOR2X1  g08964(.A(n10589), .B(n10678), .Y(n10679));
  NOR3X1  g08965(.A(n10679), .B(n10560), .C(n10563), .Y(n10680));
  AOI22X1 g08966(.A0(n10676), .A1(n10626), .B0(n10658), .B1(n10680), .Y(n10681));
  OAI21X1 g08967(.A0(n10625), .A1(n10617), .B0(n10676), .Y(n10682));
  NAND4X1 g08968(.A(n10681), .B(n10677), .C(n10671), .D(n10682), .Y(n10683));
  INVX1   g08969(.A(n10683), .Y(n10684));
  INVX1   g08970(.A(P3_REG2_REG_2__SCAN_IN), .Y(n10685));
  NAND3X1 g08971(.A(n10601), .B(n10599), .C(P3_REG0_REG_2__SCAN_IN), .Y(n10686));
  OAI21X1 g08972(.A0(n10606), .A1(n10685), .B0(n10686), .Y(n10687));
  INVX1   g08973(.A(P3_REG3_REG_2__SCAN_IN), .Y(n10688));
  INVX1   g08974(.A(P3_REG1_REG_2__SCAN_IN), .Y(n10689));
  OAI22X1 g08975(.A0(n10612), .A1(n10689), .B0(n10688), .B1(n10613), .Y(n10690));
  NOR2X1  g08976(.A(n10690), .B(n10687), .Y(n10691));
  OAI22X1 g08977(.A0(n10667), .A1(n10646), .B0(n10638), .B1(n10691), .Y(n10692));
  AOI21X1 g08978(.A0(n10670), .A1(n10633), .B0(n10692), .Y(n10693));
  NAND2X1 g08979(.A(n10693), .B(n10684), .Y(n10694));
  NAND2X1 g08980(.A(n10694), .B(n10585), .Y(n10695));
  OAI21X1 g08981(.A0(n10585), .A1(n10639), .B0(n10695), .Y(P3_U3393));
  INVX1   g08982(.A(n10585), .Y(n10697));
  NOR2X1  g08983(.A(n10667), .B(n10645), .Y(n10698));
  NAND2X1 g08984(.A(n10667), .B(n10645), .Y(n10699));
  AOI21X1 g08985(.A0(n10673), .A1(n10699), .B0(n10698), .Y(n10700));
  NOR2X1  g08986(.A(P3_IR_REG_31__SCAN_IN), .B(n10197), .Y(n10701));
  AOI21X1 g08987(.A0(n9998), .A1(P3_IR_REG_31__SCAN_IN), .B0(n10701), .Y(n10702));
  INVX1   g08988(.A(n10702), .Y(n10703));
  NOR2X1  g08989(.A(n10590), .B(n9995), .Y(n10704));
  AOI21X1 g08990(.A0(n10703), .A1(n10590), .B0(n10704), .Y(n10705));
  NOR2X1  g08991(.A(n10705), .B(n10691), .Y(n10706));
  AOI22X1 g08992(.A0(n10652), .A1(P3_REG0_REG_2__SCAN_IN), .B0(P3_REG2_REG_2__SCAN_IN), .B1(n10653), .Y(n10707));
  AOI22X1 g08993(.A0(n10655), .A1(P3_REG1_REG_2__SCAN_IN), .B0(P3_REG3_REG_2__SCAN_IN), .B1(n10656), .Y(n10708));
  NAND2X1 g08994(.A(n10708), .B(n10707), .Y(n10709));
  NAND2X1 g08995(.A(n10703), .B(n10590), .Y(n10710));
  OAI21X1 g08996(.A0(n10590), .A1(n9995), .B0(n10710), .Y(n10711));
  NOR2X1  g08997(.A(n10711), .B(n10709), .Y(n10712));
  NOR3X1  g08998(.A(n10700), .B(n10712), .C(n10706), .Y(n10713));
  XOR2X1  g08999(.A(n10705), .B(n10709), .Y(n10714));
  AOI21X1 g09000(.A0(n10714), .A1(n10700), .B0(n10713), .Y(n10715));
  NAND2X1 g09001(.A(n10715), .B(n10622), .Y(n10716));
  OAI21X1 g09002(.A0(n10625), .A1(n10617), .B0(n10715), .Y(n10717));
  INVX1   g09003(.A(n10623), .Y(n10718));
  NAND2X1 g09004(.A(n10665), .B(n10590), .Y(n10719));
  OAI21X1 g09005(.A0(n10590), .A1(n9979), .B0(n10719), .Y(n10720));
  NOR2X1  g09006(.A(n10720), .B(n10645), .Y(n10721));
  AOI21X1 g09007(.A0(n10615), .A1(n10595), .B0(n10645), .Y(n10722));
  AOI21X1 g09008(.A0(n10615), .A1(n10595), .B0(n10720), .Y(n10723));
  NOR3X1  g09009(.A(n10723), .B(n10722), .C(n10721), .Y(n10724));
  XOR2X1  g09010(.A(n10724), .B(n10714), .Y(n10725));
  AOI22X1 g09011(.A0(n10680), .A1(n10662), .B0(n10626), .B1(n10715), .Y(n10726));
  OAI21X1 g09012(.A0(n10725), .A1(n10718), .B0(n10726), .Y(n10727));
  INVX1   g09013(.A(n10628), .Y(n10728));
  INVX1   g09014(.A(n10629), .Y(n10729));
  AOI21X1 g09015(.A0(n10729), .A1(n10728), .B0(n10725), .Y(n10730));
  NOR2X1  g09016(.A(n10730), .B(n10727), .Y(n10731));
  NAND3X1 g09017(.A(n10731), .B(n10717), .C(n10716), .Y(n10732));
  INVX1   g09018(.A(n10633), .Y(n10733));
  INVX1   g09019(.A(n10646), .Y(n10734));
  AOI22X1 g09020(.A0(n10652), .A1(P3_REG0_REG_3__SCAN_IN), .B0(P3_REG2_REG_3__SCAN_IN), .B1(n10653), .Y(n10735));
  INVX1   g09021(.A(P3_REG3_REG_3__SCAN_IN), .Y(n10736));
  AOI22X1 g09022(.A0(n10655), .A1(P3_REG1_REG_3__SCAN_IN), .B0(n10736), .B1(n10656), .Y(n10737));
  NAND2X1 g09023(.A(n10737), .B(n10735), .Y(n10738));
  AOI22X1 g09024(.A0(n10711), .A1(n10734), .B0(n10637), .B1(n10738), .Y(n10739));
  OAI21X1 g09025(.A0(n10725), .A1(n10733), .B0(n10739), .Y(n10740));
  NOR2X1  g09026(.A(n10740), .B(n10732), .Y(n10741));
  NAND2X1 g09027(.A(n10697), .B(P3_REG0_REG_2__SCAN_IN), .Y(n10742));
  OAI21X1 g09028(.A0(n10741), .A1(n10697), .B0(n10742), .Y(P3_U3396));
  INVX1   g09029(.A(n10622), .Y(n10744));
  OAI21X1 g09030(.A0(n10720), .A1(n10662), .B0(n10673), .Y(n10745));
  NOR3X1  g09031(.A(n10712), .B(n10667), .C(n10645), .Y(n10746));
  NOR2X1  g09032(.A(n10746), .B(n10706), .Y(n10747));
  OAI21X1 g09033(.A0(n10745), .A1(n10712), .B0(n10747), .Y(n10748));
  NOR2X1  g09034(.A(P3_IR_REG_31__SCAN_IN), .B(n10007), .Y(n10749));
  AOI21X1 g09035(.A0(n10009), .A1(P3_IR_REG_31__SCAN_IN), .B0(n10749), .Y(n10750));
  INVX1   g09036(.A(n10750), .Y(n10751));
  NOR2X1  g09037(.A(n10590), .B(n10006), .Y(n10752));
  AOI21X1 g09038(.A0(n10751), .A1(n10590), .B0(n10752), .Y(n10753));
  XOR2X1  g09039(.A(n10753), .B(n10738), .Y(n10754));
  NOR2X1  g09040(.A(n10748), .B(n10754), .Y(n10755));
  INVX1   g09041(.A(P3_REG2_REG_3__SCAN_IN), .Y(n10756));
  NAND3X1 g09042(.A(n10601), .B(n10599), .C(P3_REG0_REG_3__SCAN_IN), .Y(n10757));
  OAI21X1 g09043(.A0(n10606), .A1(n10756), .B0(n10757), .Y(n10758));
  INVX1   g09044(.A(P3_REG1_REG_3__SCAN_IN), .Y(n10759));
  OAI22X1 g09045(.A0(n10612), .A1(n10759), .B0(P3_REG3_REG_3__SCAN_IN), .B1(n10613), .Y(n10760));
  NOR2X1  g09046(.A(n10760), .B(n10758), .Y(n10761));
  XOR2X1  g09047(.A(n10753), .B(n10761), .Y(n10762));
  AOI21X1 g09048(.A0(n10754), .A1(n10748), .B0(n10755), .Y(n10764));
  NOR2X1  g09049(.A(n10764), .B(n10744), .Y(n10765));
  INVX1   g09050(.A(n10625), .Y(n10766));
  AOI21X1 g09051(.A0(n10766), .A1(n10618), .B0(n10764), .Y(n10767));
  NOR2X1  g09052(.A(n10767), .B(n10765), .Y(n10768));
  NOR2X1  g09053(.A(n10711), .B(n10691), .Y(n10769));
  NAND2X1 g09054(.A(n10667), .B(n10662), .Y(n10770));
  OAI21X1 g09055(.A0(n10658), .A1(n10635), .B0(n10662), .Y(n10771));
  OAI21X1 g09056(.A0(n10658), .A1(n10635), .B0(n10667), .Y(n10772));
  NAND3X1 g09057(.A(n10772), .B(n10771), .C(n10770), .Y(n10773));
  NOR2X1  g09058(.A(n10705), .B(n10709), .Y(n10774));
  NOR2X1  g09059(.A(n10754), .B(n10774), .Y(n10775));
  OAI21X1 g09060(.A0(n10773), .A1(n10769), .B0(n10775), .Y(n10776));
  NOR2X1  g09061(.A(n10724), .B(n10774), .Y(n10777));
  OAI21X1 g09062(.A0(n10711), .A1(n10691), .B0(n10754), .Y(n10778));
  OAI21X1 g09063(.A0(n10778), .A1(n10777), .B0(n10776), .Y(n10779));
  INVX1   g09064(.A(n10626), .Y(n10780));
  INVX1   g09065(.A(n10680), .Y(n10781));
  OAI22X1 g09066(.A0(n10691), .A1(n10781), .B0(n10780), .B1(n10764), .Y(n10782));
  AOI21X1 g09067(.A0(n10779), .A1(n10623), .B0(n10782), .Y(n10783));
  OAI21X1 g09068(.A0(n10629), .A1(n10628), .B0(n10779), .Y(n10784));
  NAND3X1 g09069(.A(n10784), .B(n10783), .C(n10768), .Y(n10785));
  NAND2X1 g09070(.A(n10779), .B(n10633), .Y(n10786));
  NAND2X1 g09071(.A(n10751), .B(n10590), .Y(n10787));
  OAI21X1 g09072(.A0(n10590), .A1(n10006), .B0(n10787), .Y(n10788));
  AOI22X1 g09073(.A0(n10652), .A1(P3_REG0_REG_4__SCAN_IN), .B0(P3_REG2_REG_4__SCAN_IN), .B1(n10653), .Y(n10789));
  XOR2X1  g09074(.A(P3_REG3_REG_4__SCAN_IN), .B(P3_REG3_REG_3__SCAN_IN), .Y(n10790));
  INVX1   g09075(.A(n10790), .Y(n10791));
  AOI22X1 g09076(.A0(n10656), .A1(n10791), .B0(n10655), .B1(P3_REG1_REG_4__SCAN_IN), .Y(n10792));
  NAND2X1 g09077(.A(n10792), .B(n10789), .Y(n10793));
  AOI22X1 g09078(.A0(n10788), .A1(n10734), .B0(n10637), .B1(n10793), .Y(n10794));
  NAND2X1 g09079(.A(n10794), .B(n10786), .Y(n10795));
  NOR2X1  g09080(.A(n10795), .B(n10785), .Y(n10796));
  NAND2X1 g09081(.A(n10697), .B(P3_REG0_REG_3__SCAN_IN), .Y(n10797));
  OAI21X1 g09082(.A0(n10796), .A1(n10697), .B0(n10797), .Y(P3_U3399));
  NOR2X1  g09083(.A(P3_IR_REG_31__SCAN_IN), .B(n10022), .Y(n10799));
  INVX1   g09084(.A(n10799), .Y(n10800));
  OAI21X1 g09085(.A0(n10025), .A1(n9982), .B0(n10800), .Y(n10801));
  NOR2X1  g09086(.A(n10590), .B(n10021), .Y(n10802));
  AOI21X1 g09087(.A0(n10801), .A1(n10590), .B0(n10802), .Y(n10803));
  XOR2X1  g09088(.A(n10803), .B(n10793), .Y(n10804));
  NOR2X1  g09089(.A(n10753), .B(n10761), .Y(n10806));
  NOR2X1  g09090(.A(n10788), .B(n10738), .Y(n10807));
  NOR2X1  g09091(.A(n10807), .B(n10747), .Y(n10808));
  NOR3X1  g09092(.A(n10807), .B(n10745), .C(n10712), .Y(n10809));
  NOR3X1  g09093(.A(n10809), .B(n10808), .C(n10806), .Y(n10810));
  INVX1   g09094(.A(P3_REG2_REG_4__SCAN_IN), .Y(n10811));
  NAND3X1 g09095(.A(n10601), .B(n10599), .C(P3_REG0_REG_4__SCAN_IN), .Y(n10812));
  OAI21X1 g09096(.A0(n10606), .A1(n10811), .B0(n10812), .Y(n10813));
  INVX1   g09097(.A(P3_REG1_REG_4__SCAN_IN), .Y(n10814));
  OAI22X1 g09098(.A0(n10613), .A1(n10790), .B0(n10612), .B1(n10814), .Y(n10815));
  NOR2X1  g09099(.A(n10815), .B(n10813), .Y(n10816));
  XOR2X1  g09100(.A(n10803), .B(n10816), .Y(n10817));
  NOR2X1  g09101(.A(n10817), .B(n10810), .Y(n10818));
  AOI21X1 g09102(.A0(n10810), .A1(n10817), .B0(n10818), .Y(n10819));
  NOR2X1  g09103(.A(n10819), .B(n10744), .Y(n10820));
  AOI21X1 g09104(.A0(n10766), .A1(n10618), .B0(n10819), .Y(n10821));
  NOR2X1  g09105(.A(n10821), .B(n10820), .Y(n10822));
  AOI22X1 g09106(.A0(n10761), .A1(n10788), .B0(n10711), .B1(n10691), .Y(n10823));
  AOI21X1 g09107(.A0(n10705), .A1(n10709), .B0(n10738), .Y(n10824));
  NAND3X1 g09108(.A(n10738), .B(n10705), .C(n10709), .Y(n10825));
  OAI21X1 g09109(.A0(n10824), .A1(n10788), .B0(n10825), .Y(n10826));
  AOI21X1 g09110(.A0(n10823), .A1(n10773), .B0(n10826), .Y(n10827));
  XOR2X1  g09111(.A(n10827), .B(n10804), .Y(n10828));
  INVX1   g09112(.A(n10828), .Y(n10829));
  OAI22X1 g09113(.A0(n10761), .A1(n10781), .B0(n10780), .B1(n10819), .Y(n10830));
  AOI21X1 g09114(.A0(n10829), .A1(n10623), .B0(n10830), .Y(n10831));
  OAI21X1 g09115(.A0(n10629), .A1(n10628), .B0(n10829), .Y(n10832));
  NAND3X1 g09116(.A(n10832), .B(n10831), .C(n10822), .Y(n10833));
  NAND2X1 g09117(.A(n10801), .B(n10590), .Y(n10834));
  OAI21X1 g09118(.A0(n10590), .A1(n10021), .B0(n10834), .Y(n10835));
  NAND3X1 g09119(.A(n10601), .B(n10599), .C(P3_REG0_REG_5__SCAN_IN), .Y(n10836));
  NAND3X1 g09120(.A(n10601), .B(n10605), .C(P3_REG2_REG_5__SCAN_IN), .Y(n10837));
  NAND3X1 g09121(.A(n10611), .B(n10599), .C(P3_REG1_REG_5__SCAN_IN), .Y(n10838));
  INVX1   g09122(.A(P3_REG3_REG_5__SCAN_IN), .Y(n10839));
  NOR2X1  g09123(.A(P3_REG3_REG_4__SCAN_IN), .B(P3_REG3_REG_3__SCAN_IN), .Y(n10840));
  XOR2X1  g09124(.A(n10840), .B(n10839), .Y(n10841));
  INVX1   g09125(.A(n10841), .Y(n10842));
  NAND3X1 g09126(.A(n10842), .B(n10611), .C(n10605), .Y(n10843));
  NAND4X1 g09127(.A(n10838), .B(n10837), .C(n10836), .D(n10843), .Y(n10844));
  AOI22X1 g09128(.A0(n10835), .A1(n10734), .B0(n10637), .B1(n10844), .Y(n10845));
  OAI21X1 g09129(.A0(n10828), .A1(n10733), .B0(n10845), .Y(n10846));
  NOR2X1  g09130(.A(n10846), .B(n10833), .Y(n10847));
  NAND2X1 g09131(.A(n10697), .B(P3_REG0_REG_4__SCAN_IN), .Y(n10848));
  OAI21X1 g09132(.A0(n10847), .A1(n10697), .B0(n10848), .Y(P3_U3402));
  NAND2X1 g09133(.A(n10835), .B(n10793), .Y(n10850));
  NOR2X1  g09134(.A(P3_IR_REG_31__SCAN_IN), .B(n10047), .Y(n10851));
  AOI21X1 g09135(.A0(n10038), .A1(P3_IR_REG_31__SCAN_IN), .B0(n10851), .Y(n10852));
  INVX1   g09136(.A(n10852), .Y(n10853));
  NAND2X1 g09137(.A(n10853), .B(n10590), .Y(n10854));
  OAI21X1 g09138(.A0(n10590), .A1(n10037), .B0(n10854), .Y(n10855));
  INVX1   g09139(.A(P3_REG2_REG_5__SCAN_IN), .Y(n10856));
  OAI21X1 g09140(.A0(n10606), .A1(n10856), .B0(n10836), .Y(n10857));
  OAI21X1 g09141(.A0(n10841), .A1(n10613), .B0(n10838), .Y(n10858));
  NOR2X1  g09142(.A(n10858), .B(n10857), .Y(n10859));
  NOR2X1  g09143(.A(n10590), .B(n10037), .Y(n10860));
  AOI21X1 g09144(.A0(n10853), .A1(n10590), .B0(n10860), .Y(n10861));
  AOI22X1 g09145(.A0(n10859), .A1(n10861), .B0(n10803), .B1(n10816), .Y(n10862));
  INVX1   g09146(.A(n10862), .Y(n10863));
  AOI21X1 g09147(.A0(n10855), .A1(n10844), .B0(n10863), .Y(n10864));
  INVX1   g09148(.A(n10864), .Y(n10865));
  AOI21X1 g09149(.A0(n10850), .A1(n10810), .B0(n10865), .Y(n10866));
  INVX1   g09150(.A(n10850), .Y(n10867));
  AOI21X1 g09151(.A0(n10803), .A1(n10816), .B0(n10810), .Y(n10868));
  NOR2X1  g09152(.A(n10855), .B(n10859), .Y(n10869));
  NOR2X1  g09153(.A(n10861), .B(n10844), .Y(n10870));
  NOR4X1  g09154(.A(n10869), .B(n10868), .C(n10867), .D(n10870), .Y(n10871));
  NOR2X1  g09155(.A(n10871), .B(n10866), .Y(n10872));
  INVX1   g09156(.A(n10872), .Y(n10873));
  OAI22X1 g09157(.A0(n10816), .A1(n10781), .B0(n10780), .B1(n10873), .Y(n10874));
  OAI21X1 g09158(.A0(n10625), .A1(n10617), .B0(n10872), .Y(n10875));
  OAI21X1 g09159(.A0(n10873), .A1(n10744), .B0(n10875), .Y(n10876));
  XOR2X1  g09160(.A(n10861), .B(n10844), .Y(n10877));
  NOR2X1  g09161(.A(n10835), .B(n10816), .Y(n10878));
  NAND2X1 g09162(.A(n10835), .B(n10816), .Y(n10879));
  OAI22X1 g09163(.A0(n10738), .A1(n10753), .B0(n10705), .B1(n10709), .Y(n10880));
  OAI21X1 g09164(.A0(n10711), .A1(n10691), .B0(n10761), .Y(n10881));
  NOR3X1  g09165(.A(n10761), .B(n10711), .C(n10691), .Y(n10882));
  AOI21X1 g09166(.A0(n10881), .A1(n10753), .B0(n10882), .Y(n10883));
  OAI21X1 g09167(.A0(n10880), .A1(n10724), .B0(n10883), .Y(n10884));
  AOI21X1 g09168(.A0(n10884), .A1(n10879), .B0(n10878), .Y(n10885));
  XOR2X1  g09169(.A(n10885), .B(n10877), .Y(n10886));
  INVX1   g09170(.A(n10886), .Y(n10887));
  OAI21X1 g09171(.A0(n10628), .A1(n10623), .B0(n10887), .Y(n10888));
  OAI21X1 g09172(.A0(n10886), .A1(n10729), .B0(n10888), .Y(n10889));
  AOI22X1 g09173(.A0(n10652), .A1(P3_REG0_REG_6__SCAN_IN), .B0(P3_REG2_REG_6__SCAN_IN), .B1(n10653), .Y(n10890));
  NOR4X1  g09174(.A(P3_REG3_REG_4__SCAN_IN), .B(P3_REG3_REG_5__SCAN_IN), .C(P3_REG3_REG_3__SCAN_IN), .D(P3_REG3_REG_6__SCAN_IN), .Y(n10891));
  INVX1   g09175(.A(P3_REG3_REG_6__SCAN_IN), .Y(n10892));
  AOI21X1 g09176(.A0(n10840), .A1(n10839), .B0(n10892), .Y(n10893));
  NOR2X1  g09177(.A(n10893), .B(n10891), .Y(n10894));
  INVX1   g09178(.A(n10894), .Y(n10895));
  AOI22X1 g09179(.A0(n10656), .A1(n10895), .B0(n10655), .B1(P3_REG1_REG_6__SCAN_IN), .Y(n10896));
  NAND2X1 g09180(.A(n10896), .B(n10890), .Y(n10897));
  AOI22X1 g09181(.A0(n10855), .A1(n10734), .B0(n10637), .B1(n10897), .Y(n10898));
  OAI21X1 g09182(.A0(n10886), .A1(n10733), .B0(n10898), .Y(n10899));
  NOR4X1  g09183(.A(n10889), .B(n10876), .C(n10874), .D(n10899), .Y(n10900));
  NAND2X1 g09184(.A(n10697), .B(P3_REG0_REG_5__SCAN_IN), .Y(n10901));
  OAI21X1 g09185(.A0(n10900), .A1(n10697), .B0(n10901), .Y(P3_U3405));
  NOR2X1  g09186(.A(n10700), .B(n10712), .Y(n10903));
  NOR3X1  g09187(.A(n10903), .B(n10806), .C(n10706), .Y(n10904));
  OAI21X1 g09188(.A0(n10788), .A1(n10738), .B0(n10862), .Y(n10905));
  AOI21X1 g09189(.A0(n10861), .A1(n10850), .B0(n10859), .Y(n10906));
  AOI21X1 g09190(.A0(n10855), .A1(n10867), .B0(n10906), .Y(n10907));
  OAI21X1 g09191(.A0(n10905), .A1(n10904), .B0(n10907), .Y(n10908));
  INVX1   g09192(.A(P3_REG2_REG_6__SCAN_IN), .Y(n10909));
  NAND3X1 g09193(.A(n10601), .B(n10599), .C(P3_REG0_REG_6__SCAN_IN), .Y(n10910));
  OAI21X1 g09194(.A0(n10606), .A1(n10909), .B0(n10910), .Y(n10911));
  INVX1   g09195(.A(P3_REG1_REG_6__SCAN_IN), .Y(n10912));
  OAI22X1 g09196(.A0(n10613), .A1(n10894), .B0(n10612), .B1(n10912), .Y(n10913));
  NOR2X1  g09197(.A(n10913), .B(n10911), .Y(n10914));
  NOR2X1  g09198(.A(P3_IR_REG_31__SCAN_IN), .B(n10049), .Y(n10915));
  AOI21X1 g09199(.A0(n10052), .A1(P3_IR_REG_31__SCAN_IN), .B0(n10915), .Y(n10916));
  INVX1   g09200(.A(n10916), .Y(n10917));
  NAND2X1 g09201(.A(n10917), .B(n10590), .Y(n10918));
  OAI21X1 g09202(.A0(n10590), .A1(n10046), .B0(n10918), .Y(n10919));
  XOR2X1  g09203(.A(n10919), .B(n10914), .Y(n10920));
  NOR2X1  g09204(.A(n10908), .B(n10920), .Y(n10921));
  AOI21X1 g09205(.A0(n10920), .A1(n10908), .B0(n10921), .Y(n10923));
  OAI22X1 g09206(.A0(n10859), .A1(n10781), .B0(n10780), .B1(n10923), .Y(n10924));
  INVX1   g09207(.A(n10923), .Y(n10925));
  OAI21X1 g09208(.A0(n10625), .A1(n10617), .B0(n10925), .Y(n10926));
  OAI21X1 g09209(.A0(n10923), .A1(n10744), .B0(n10926), .Y(n10927));
  OAI21X1 g09210(.A0(n10855), .A1(n10859), .B0(n10885), .Y(n10928));
  NOR2X1  g09211(.A(n10920), .B(n10870), .Y(n10929));
  NAND2X1 g09212(.A(n10929), .B(n10928), .Y(n10930));
  NOR2X1  g09213(.A(n10590), .B(n10046), .Y(n10931));
  AOI21X1 g09214(.A0(n10917), .A1(n10590), .B0(n10931), .Y(n10932));
  NOR2X1  g09215(.A(n10932), .B(n10897), .Y(n10933));
  OAI22X1 g09216(.A0(n10914), .A1(n10919), .B0(n10855), .B1(n10859), .Y(n10934));
  NOR2X1  g09217(.A(n10934), .B(n10933), .Y(n10935));
  OAI21X1 g09218(.A0(n10885), .A1(n10870), .B0(n10935), .Y(n10936));
  NAND2X1 g09219(.A(n10936), .B(n10930), .Y(n10937));
  INVX1   g09220(.A(n10937), .Y(n10938));
  OAI21X1 g09221(.A0(n10628), .A1(n10623), .B0(n10937), .Y(n10939));
  OAI21X1 g09222(.A0(n10938), .A1(n10729), .B0(n10939), .Y(n10940));
  AOI22X1 g09223(.A0(n10652), .A1(P3_REG0_REG_7__SCAN_IN), .B0(P3_REG2_REG_7__SCAN_IN), .B1(n10653), .Y(n10941));
  INVX1   g09224(.A(P3_REG3_REG_7__SCAN_IN), .Y(n10942));
  XOR2X1  g09225(.A(n10891), .B(n10942), .Y(n10943));
  INVX1   g09226(.A(n10943), .Y(n10944));
  AOI22X1 g09227(.A0(n10656), .A1(n10944), .B0(n10655), .B1(P3_REG1_REG_7__SCAN_IN), .Y(n10945));
  NAND2X1 g09228(.A(n10945), .B(n10941), .Y(n10946));
  AOI22X1 g09229(.A0(n10919), .A1(n10734), .B0(n10637), .B1(n10946), .Y(n10947));
  OAI21X1 g09230(.A0(n10938), .A1(n10733), .B0(n10947), .Y(n10948));
  NOR4X1  g09231(.A(n10940), .B(n10927), .C(n10924), .D(n10948), .Y(n10949));
  NAND2X1 g09232(.A(n10697), .B(P3_REG0_REG_6__SCAN_IN), .Y(n10950));
  OAI21X1 g09233(.A0(n10949), .A1(n10697), .B0(n10950), .Y(P3_U3408));
  INVX1   g09234(.A(P3_REG2_REG_7__SCAN_IN), .Y(n10952));
  NAND3X1 g09235(.A(n10601), .B(n10599), .C(P3_REG0_REG_7__SCAN_IN), .Y(n10953));
  OAI21X1 g09236(.A0(n10606), .A1(n10952), .B0(n10953), .Y(n10954));
  INVX1   g09237(.A(P3_REG1_REG_7__SCAN_IN), .Y(n10955));
  OAI22X1 g09238(.A0(n10613), .A1(n10943), .B0(n10612), .B1(n10955), .Y(n10956));
  NOR2X1  g09239(.A(n10956), .B(n10954), .Y(n10957));
  NOR2X1  g09240(.A(P3_IR_REG_31__SCAN_IN), .B(n10065), .Y(n10958));
  AOI21X1 g09241(.A0(n10066), .A1(P3_IR_REG_31__SCAN_IN), .B0(n10958), .Y(n10959));
  INVX1   g09242(.A(n10959), .Y(n10960));
  NAND2X1 g09243(.A(n10960), .B(n10590), .Y(n10961));
  OAI21X1 g09244(.A0(n10590), .A1(n10064), .B0(n10961), .Y(n10962));
  XOR2X1  g09245(.A(n10962), .B(n10957), .Y(n10963));
  NAND2X1 g09246(.A(n10855), .B(n10859), .Y(n10964));
  AOI21X1 g09247(.A0(n10964), .A1(n10878), .B0(n10934), .Y(n10965));
  NOR2X1  g09248(.A(n10965), .B(n10933), .Y(n10966));
  OAI22X1 g09249(.A0(n10897), .A1(n10932), .B0(n10803), .B1(n10793), .Y(n10967));
  NOR2X1  g09250(.A(n10967), .B(n10870), .Y(n10968));
  AOI21X1 g09251(.A0(n10968), .A1(n10884), .B0(n10966), .Y(n10969));
  XOR2X1  g09252(.A(n10969), .B(n10963), .Y(n10970));
  INVX1   g09253(.A(n10970), .Y(n10971));
  OAI21X1 g09254(.A0(n10629), .A1(n10623), .B0(n10971), .Y(n10972));
  INVX1   g09255(.A(n10908), .Y(n10973));
  NOR2X1  g09256(.A(n10932), .B(n10914), .Y(n10974));
  INVX1   g09257(.A(n10974), .Y(n10975));
  NOR2X1  g09258(.A(n10590), .B(n10064), .Y(n10976));
  AOI21X1 g09259(.A0(n10960), .A1(n10590), .B0(n10976), .Y(n10977));
  AOI22X1 g09260(.A0(n10957), .A1(n10977), .B0(n10932), .B1(n10914), .Y(n10978));
  OAI21X1 g09261(.A0(n10977), .A1(n10957), .B0(n10978), .Y(n10979));
  AOI21X1 g09262(.A0(n10975), .A1(n10973), .B0(n10979), .Y(n10980));
  OAI21X1 g09263(.A0(n10919), .A1(n10897), .B0(n10908), .Y(n10981));
  NAND2X1 g09264(.A(n10977), .B(n10946), .Y(n10982));
  INVX1   g09265(.A(n10982), .Y(n10983));
  NOR2X1  g09266(.A(n10977), .B(n10946), .Y(n10984));
  NOR3X1  g09267(.A(n10984), .B(n10983), .C(n10974), .Y(n10985));
  AOI21X1 g09268(.A0(n10985), .A1(n10981), .B0(n10980), .Y(n10986));
  AOI22X1 g09269(.A0(n10971), .A1(n10628), .B0(n10622), .B1(n10986), .Y(n10987));
  AOI22X1 g09270(.A0(n10897), .A1(n10680), .B0(n10626), .B1(n10986), .Y(n10988));
  OAI21X1 g09271(.A0(n10625), .A1(n10617), .B0(n10986), .Y(n10989));
  NAND4X1 g09272(.A(n10988), .B(n10987), .C(n10972), .D(n10989), .Y(n10990));
  AOI22X1 g09273(.A0(n10652), .A1(P3_REG0_REG_8__SCAN_IN), .B0(P3_REG2_REG_8__SCAN_IN), .B1(n10653), .Y(n10991));
  NAND2X1 g09274(.A(n10891), .B(n10942), .Y(n10992));
  XOR2X1  g09275(.A(n10992), .B(P3_REG3_REG_8__SCAN_IN), .Y(n10993));
  INVX1   g09276(.A(n10993), .Y(n10994));
  AOI22X1 g09277(.A0(n10656), .A1(n10994), .B0(n10655), .B1(P3_REG1_REG_8__SCAN_IN), .Y(n10995));
  NAND2X1 g09278(.A(n10995), .B(n10991), .Y(n10996));
  AOI22X1 g09279(.A0(n10962), .A1(n10734), .B0(n10637), .B1(n10996), .Y(n10997));
  OAI21X1 g09280(.A0(n10970), .A1(n10733), .B0(n10997), .Y(n10998));
  NOR2X1  g09281(.A(n10998), .B(n10990), .Y(n10999));
  NAND2X1 g09282(.A(n10697), .B(P3_REG0_REG_7__SCAN_IN), .Y(n11000));
  OAI21X1 g09283(.A0(n10999), .A1(n10697), .B0(n11000), .Y(P3_U3411));
  NOR2X1  g09284(.A(P3_IR_REG_31__SCAN_IN), .B(n10077), .Y(n11002));
  AOI21X1 g09285(.A0(n10080), .A1(P3_IR_REG_31__SCAN_IN), .B0(n11002), .Y(n11003));
  INVX1   g09286(.A(n11003), .Y(n11004));
  NAND2X1 g09287(.A(n11004), .B(n10590), .Y(n11005));
  OAI21X1 g09288(.A0(n10590), .A1(n10076), .B0(n11005), .Y(n11006));
  XOR2X1  g09289(.A(n11006), .B(n10996), .Y(n11007));
  OAI21X1 g09290(.A0(n10977), .A1(n10946), .B0(n11007), .Y(n11008));
  AOI21X1 g09291(.A0(n10969), .A1(n10982), .B0(n11008), .Y(n11009));
  NOR2X1  g09292(.A(n10969), .B(n10984), .Y(n11010));
  NOR3X1  g09293(.A(n11010), .B(n11007), .C(n10983), .Y(n11011));
  NOR2X1  g09294(.A(n11011), .B(n11009), .Y(n11012));
  AOI21X1 g09295(.A0(n10729), .A1(n10718), .B0(n11012), .Y(n11013));
  OAI21X1 g09296(.A0(n10962), .A1(n10974), .B0(n10946), .Y(n11014));
  OAI21X1 g09297(.A0(n10977), .A1(n10975), .B0(n11014), .Y(n11015));
  AOI21X1 g09298(.A0(n10978), .A1(n10908), .B0(n11015), .Y(n11016));
  NOR2X1  g09299(.A(n11007), .B(n11016), .Y(n11018));
  AOI21X1 g09300(.A0(n11016), .A1(n11007), .B0(n11018), .Y(n11019));
  OAI22X1 g09301(.A0(n11012), .A1(n10728), .B0(n10744), .B1(n11019), .Y(n11020));
  NOR2X1  g09302(.A(n11020), .B(n11013), .Y(n11021));
  INVX1   g09303(.A(n11019), .Y(n11022));
  AOI22X1 g09304(.A0(n10946), .A1(n10680), .B0(n10626), .B1(n11022), .Y(n11023));
  OAI21X1 g09305(.A0(n10625), .A1(n10617), .B0(n11022), .Y(n11024));
  NAND3X1 g09306(.A(n11024), .B(n11023), .C(n11021), .Y(n11025));
  AOI22X1 g09307(.A0(n10652), .A1(P3_REG0_REG_9__SCAN_IN), .B0(P3_REG2_REG_9__SCAN_IN), .B1(n10653), .Y(n11026));
  INVX1   g09308(.A(P3_REG1_REG_9__SCAN_IN), .Y(n11027));
  NOR3X1  g09309(.A(n10601), .B(n10605), .C(n11027), .Y(n11028));
  NOR3X1  g09310(.A(n10992), .B(P3_REG3_REG_9__SCAN_IN), .C(P3_REG3_REG_8__SCAN_IN), .Y(n11029));
  INVX1   g09311(.A(n11029), .Y(n11030));
  OAI21X1 g09312(.A0(n10992), .A1(P3_REG3_REG_8__SCAN_IN), .B0(P3_REG3_REG_9__SCAN_IN), .Y(n11031));
  NAND2X1 g09313(.A(n11031), .B(n11030), .Y(n11032));
  INVX1   g09314(.A(n11032), .Y(n11033));
  NOR3X1  g09315(.A(n11033), .B(n10601), .C(n10599), .Y(n11034));
  NOR2X1  g09316(.A(n11034), .B(n11028), .Y(n11035));
  NAND2X1 g09317(.A(n11035), .B(n11026), .Y(n11036));
  AOI22X1 g09318(.A0(n11006), .A1(n10734), .B0(n10637), .B1(n11036), .Y(n11037));
  OAI21X1 g09319(.A0(n11012), .A1(n10733), .B0(n11037), .Y(n11038));
  NOR2X1  g09320(.A(n11038), .B(n11025), .Y(n11039));
  NAND2X1 g09321(.A(n10697), .B(P3_REG0_REG_8__SCAN_IN), .Y(n11040));
  OAI21X1 g09322(.A0(n11039), .A1(n10697), .B0(n11040), .Y(P3_U3414));
  NOR2X1  g09323(.A(n11006), .B(n10996), .Y(n11042));
  NAND2X1 g09324(.A(n11006), .B(n10996), .Y(n11043));
  OAI21X1 g09325(.A0(n11042), .A1(n11016), .B0(n11043), .Y(n11044));
  INVX1   g09326(.A(n11036), .Y(n11045));
  NOR2X1  g09327(.A(P3_IR_REG_31__SCAN_IN), .B(n10097), .Y(n11046));
  AOI21X1 g09328(.A0(n10098), .A1(P3_IR_REG_31__SCAN_IN), .B0(n11046), .Y(n11047));
  INVX1   g09329(.A(n11047), .Y(n11048));
  NAND2X1 g09330(.A(n11048), .B(n10590), .Y(n11049));
  OAI21X1 g09331(.A0(n10590), .A1(n10096), .B0(n11049), .Y(n11050));
  XOR2X1  g09332(.A(n11050), .B(n11045), .Y(n11051));
  NOR2X1  g09333(.A(n11044), .B(n11051), .Y(n11052));
  AOI21X1 g09334(.A0(n11051), .A1(n11044), .B0(n11052), .Y(n11054));
  NOR2X1  g09335(.A(n11054), .B(n10780), .Y(n11055));
  INVX1   g09336(.A(P3_REG2_REG_8__SCAN_IN), .Y(n11056));
  NAND3X1 g09337(.A(n10601), .B(n10599), .C(P3_REG0_REG_8__SCAN_IN), .Y(n11057));
  OAI21X1 g09338(.A0(n10606), .A1(n11056), .B0(n11057), .Y(n11058));
  INVX1   g09339(.A(P3_REG1_REG_8__SCAN_IN), .Y(n11059));
  OAI22X1 g09340(.A0(n10613), .A1(n10993), .B0(n10612), .B1(n11059), .Y(n11060));
  NOR2X1  g09341(.A(n11060), .B(n11058), .Y(n11061));
  AOI22X1 g09342(.A0(n11061), .A1(n11006), .B0(n10962), .B1(n10957), .Y(n11062));
  INVX1   g09343(.A(n11062), .Y(n11063));
  NOR4X1  g09344(.A(n10967), .B(n10870), .C(n10827), .D(n11063), .Y(n11064));
  NOR3X1  g09345(.A(n10870), .B(n10835), .C(n10816), .Y(n11065));
  OAI22X1 g09346(.A0(n10934), .A1(n11065), .B0(n10932), .B1(n10897), .Y(n11066));
  OAI21X1 g09347(.A0(n11061), .A1(n10982), .B0(n11006), .Y(n11067));
  OAI21X1 g09348(.A0(n10962), .A1(n10957), .B0(n11061), .Y(n11068));
  NAND2X1 g09349(.A(n11068), .B(n11067), .Y(n11069));
  OAI21X1 g09350(.A0(n11063), .A1(n11066), .B0(n11069), .Y(n11070));
  NOR2X1  g09351(.A(n11070), .B(n11064), .Y(n11071));
  XOR2X1  g09352(.A(n11071), .B(n11051), .Y(n11072));
  INVX1   g09353(.A(n11072), .Y(n11073));
  AOI22X1 g09354(.A0(n10996), .A1(n10680), .B0(n10628), .B1(n11073), .Y(n11074));
  OAI21X1 g09355(.A0(n10629), .A1(n10623), .B0(n11073), .Y(n11075));
  NAND2X1 g09356(.A(n11075), .B(n11074), .Y(n11076));
  NOR2X1  g09357(.A(n11054), .B(n10744), .Y(n11077));
  AOI21X1 g09358(.A0(n10766), .A1(n10618), .B0(n11054), .Y(n11078));
  NOR4X1  g09359(.A(n11077), .B(n11076), .C(n11055), .D(n11078), .Y(n11079));
  INVX1   g09360(.A(n11079), .Y(n11080));
  AOI22X1 g09361(.A0(n10652), .A1(P3_REG0_REG_10__SCAN_IN), .B0(P3_REG2_REG_10__SCAN_IN), .B1(n10653), .Y(n11081));
  INVX1   g09362(.A(P3_REG3_REG_10__SCAN_IN), .Y(n11082));
  XOR2X1  g09363(.A(n11029), .B(n11082), .Y(n11083));
  INVX1   g09364(.A(n11083), .Y(n11084));
  AOI22X1 g09365(.A0(n10656), .A1(n11084), .B0(n10655), .B1(P3_REG1_REG_10__SCAN_IN), .Y(n11085));
  NAND2X1 g09366(.A(n11085), .B(n11081), .Y(n11086));
  AOI22X1 g09367(.A0(n11050), .A1(n10734), .B0(n10637), .B1(n11086), .Y(n11087));
  OAI21X1 g09368(.A0(n11072), .A1(n10733), .B0(n11087), .Y(n11088));
  NOR2X1  g09369(.A(n11088), .B(n11080), .Y(n11089));
  NAND2X1 g09370(.A(n10697), .B(P3_REG0_REG_9__SCAN_IN), .Y(n11090));
  OAI21X1 g09371(.A0(n11089), .A1(n10697), .B0(n11090), .Y(P3_U3417));
  INVX1   g09372(.A(n11050), .Y(n11092));
  NOR2X1  g09373(.A(n11092), .B(n11045), .Y(n11093));
  NOR2X1  g09374(.A(n11093), .B(n11044), .Y(n11094));
  INVX1   g09375(.A(n11086), .Y(n11095));
  NOR2X1  g09376(.A(P3_IR_REG_31__SCAN_IN), .B(n10108), .Y(n11096));
  AOI21X1 g09377(.A0(n10111), .A1(P3_IR_REG_31__SCAN_IN), .B0(n11096), .Y(n11097));
  INVX1   g09378(.A(n11097), .Y(n11098));
  NOR2X1  g09379(.A(n10590), .B(n10107), .Y(n11099));
  AOI21X1 g09380(.A0(n11098), .A1(n10590), .B0(n11099), .Y(n11100));
  NAND2X1 g09381(.A(n11098), .B(n10590), .Y(n11101));
  OAI21X1 g09382(.A0(n10590), .A1(n10107), .B0(n11101), .Y(n11102));
  OAI22X1 g09383(.A0(n11086), .A1(n11102), .B0(n11050), .B1(n11036), .Y(n11103));
  INVX1   g09384(.A(n11103), .Y(n11104));
  OAI21X1 g09385(.A0(n11100), .A1(n11095), .B0(n11104), .Y(n11105));
  INVX1   g09386(.A(n11044), .Y(n11106));
  AOI21X1 g09387(.A0(n11092), .A1(n11045), .B0(n11106), .Y(n11107));
  XOR2X1  g09388(.A(n11102), .B(n11095), .Y(n11108));
  OAI21X1 g09389(.A0(n11092), .A1(n11045), .B0(n11108), .Y(n11109));
  OAI22X1 g09390(.A0(n11107), .A1(n11109), .B0(n11105), .B1(n11094), .Y(n11110));
  AOI21X1 g09391(.A0(n11035), .A1(n11026), .B0(n11050), .Y(n11111));
  NAND3X1 g09392(.A(n11050), .B(n11035), .C(n11026), .Y(n11112));
  INVX1   g09393(.A(n11071), .Y(n11113));
  AOI21X1 g09394(.A0(n11113), .A1(n11112), .B0(n11111), .Y(n11114));
  XOR2X1  g09395(.A(n11114), .B(n11108), .Y(n11115));
  OAI22X1 g09396(.A0(n11045), .A1(n10781), .B0(n10728), .B1(n11115), .Y(n11116));
  AOI21X1 g09397(.A0(n10729), .A1(n10718), .B0(n11115), .Y(n11117));
  NOR2X1  g09398(.A(n11117), .B(n11116), .Y(n11118));
  OAI21X1 g09399(.A0(n11110), .A1(n10780), .B0(n11118), .Y(n11119));
  NOR2X1  g09400(.A(n11110), .B(n10744), .Y(n11120));
  AOI21X1 g09401(.A0(n10766), .A1(n10618), .B0(n11110), .Y(n11121));
  AOI22X1 g09402(.A0(n10652), .A1(P3_REG0_REG_11__SCAN_IN), .B0(P3_REG2_REG_11__SCAN_IN), .B1(n10653), .Y(n11122));
  INVX1   g09403(.A(P3_REG1_REG_11__SCAN_IN), .Y(n11123));
  NOR3X1  g09404(.A(n10601), .B(n10605), .C(n11123), .Y(n11124));
  NOR3X1  g09405(.A(n11030), .B(P3_REG3_REG_11__SCAN_IN), .C(P3_REG3_REG_10__SCAN_IN), .Y(n11125));
  INVX1   g09406(.A(P3_REG3_REG_11__SCAN_IN), .Y(n11126));
  AOI21X1 g09407(.A0(n11029), .A1(n11082), .B0(n11126), .Y(n11127));
  NOR2X1  g09408(.A(n11127), .B(n11125), .Y(n11128));
  NOR3X1  g09409(.A(n11128), .B(n10601), .C(n10599), .Y(n11129));
  NOR2X1  g09410(.A(n11129), .B(n11124), .Y(n11130));
  NAND2X1 g09411(.A(n11130), .B(n11122), .Y(n11131));
  AOI22X1 g09412(.A0(n11102), .A1(n10734), .B0(n10637), .B1(n11131), .Y(n11132));
  OAI21X1 g09413(.A0(n11115), .A1(n10733), .B0(n11132), .Y(n11133));
  NOR4X1  g09414(.A(n11121), .B(n11120), .C(n11119), .D(n11133), .Y(n11134));
  NAND2X1 g09415(.A(n10697), .B(P3_REG0_REG_10__SCAN_IN), .Y(n11135));
  OAI21X1 g09416(.A0(n11134), .A1(n10697), .B0(n11135), .Y(P3_U3420));
  AOI21X1 g09417(.A0(n11085), .A1(n11081), .B0(n11102), .Y(n11137));
  INVX1   g09418(.A(n11114), .Y(n11138));
  NOR2X1  g09419(.A(n11100), .B(n11086), .Y(n11139));
  INVX1   g09420(.A(n11131), .Y(n11140));
  NOR2X1  g09421(.A(P3_IR_REG_31__SCAN_IN), .B(n10122), .Y(n11141));
  AOI21X1 g09422(.A0(n10126), .A1(P3_IR_REG_31__SCAN_IN), .B0(n11141), .Y(n11142));
  INVX1   g09423(.A(n11142), .Y(n11143));
  NAND2X1 g09424(.A(n11143), .B(n10590), .Y(n11144));
  OAI21X1 g09425(.A0(n10590), .A1(n10121), .B0(n11144), .Y(n11145));
  XOR2X1  g09426(.A(n11145), .B(n11140), .Y(n11146));
  NOR2X1  g09427(.A(n11146), .B(n11139), .Y(n11147));
  OAI21X1 g09428(.A0(n11138), .A1(n11137), .B0(n11147), .Y(n11148));
  NOR2X1  g09429(.A(n10590), .B(n10121), .Y(n11149));
  AOI21X1 g09430(.A0(n11143), .A1(n10590), .B0(n11149), .Y(n11150));
  NOR2X1  g09431(.A(n11150), .B(n11131), .Y(n11151));
  OAI22X1 g09432(.A0(n11140), .A1(n11145), .B0(n11102), .B1(n11095), .Y(n11152));
  NOR2X1  g09433(.A(n11152), .B(n11151), .Y(n11153));
  OAI21X1 g09434(.A0(n11114), .A1(n11139), .B0(n11153), .Y(n11154));
  NAND2X1 g09435(.A(n11154), .B(n11148), .Y(n11155));
  OAI21X1 g09436(.A0(n10629), .A1(n10623), .B0(n11155), .Y(n11156));
  NOR2X1  g09437(.A(n11103), .B(n11042), .Y(n11157));
  INVX1   g09438(.A(n11157), .Y(n11158));
  NOR2X1  g09439(.A(n11100), .B(n11095), .Y(n11159));
  NAND2X1 g09440(.A(n11100), .B(n11095), .Y(n11160));
  OAI22X1 g09441(.A0(n11092), .A1(n11045), .B0(n11043), .B1(n11103), .Y(n11161));
  AOI21X1 g09442(.A0(n11161), .A1(n11160), .B0(n11159), .Y(n11162));
  OAI21X1 g09443(.A0(n11158), .A1(n11016), .B0(n11162), .Y(n11163));
  NOR2X1  g09444(.A(n11163), .B(n11146), .Y(n11164));
  INVX1   g09445(.A(n11163), .Y(n11165));
  XOR2X1  g09446(.A(n11145), .B(n11131), .Y(n11166));
  NOR2X1  g09447(.A(n11166), .B(n11165), .Y(n11167));
  OAI21X1 g09448(.A0(n11167), .A1(n11164), .B0(n10622), .Y(n11168));
  NAND2X1 g09449(.A(n11155), .B(n10628), .Y(n11169));
  NAND3X1 g09450(.A(n11169), .B(n11168), .C(n11156), .Y(n11170));
  OAI21X1 g09451(.A0(n11167), .A1(n11164), .B0(n10626), .Y(n11171));
  OAI21X1 g09452(.A0(n11095), .A1(n10781), .B0(n11171), .Y(n11172));
  NAND2X1 g09453(.A(n11165), .B(n11166), .Y(n11180));
  NOR2X1  g09454(.A(n11145), .B(n11131), .Y(n11181));
  NOR2X1  g09455(.A(n11150), .B(n11140), .Y(n11182));
  OAI21X1 g09456(.A0(n11182), .A1(n11181), .B0(n11163), .Y(n11183));
  AOI22X1 g09457(.A0(n11180), .A1(n11183), .B0(n10766), .B1(n10618), .Y(n11184));
  NAND2X1 g09458(.A(n11155), .B(n10633), .Y(n11185));
  AOI22X1 g09459(.A0(n10652), .A1(P3_REG0_REG_12__SCAN_IN), .B0(P3_REG2_REG_12__SCAN_IN), .B1(n10653), .Y(n11186));
  INVX1   g09460(.A(P3_REG3_REG_12__SCAN_IN), .Y(n11187));
  XOR2X1  g09461(.A(n11125), .B(n11187), .Y(n11188));
  INVX1   g09462(.A(n11188), .Y(n11189));
  AOI22X1 g09463(.A0(n10656), .A1(n11189), .B0(n10655), .B1(P3_REG1_REG_12__SCAN_IN), .Y(n11190));
  NAND2X1 g09464(.A(n11190), .B(n11186), .Y(n11191));
  AOI22X1 g09465(.A0(n11145), .A1(n10734), .B0(n10637), .B1(n11191), .Y(n11192));
  NAND2X1 g09466(.A(n11192), .B(n11185), .Y(n11193));
  NOR4X1  g09467(.A(n11184), .B(n11172), .C(n11170), .D(n11193), .Y(n11194));
  NAND2X1 g09468(.A(n10697), .B(P3_REG0_REG_11__SCAN_IN), .Y(n11195));
  OAI21X1 g09469(.A0(n11194), .A1(n10697), .B0(n11195), .Y(P3_U3423));
  INVX1   g09470(.A(P3_IR_REG_12__SCAN_IN), .Y(n11197));
  NOR2X1  g09471(.A(P3_IR_REG_31__SCAN_IN), .B(n11197), .Y(n11198));
  AOI21X1 g09472(.A0(n10143), .A1(P3_IR_REG_31__SCAN_IN), .B0(n11198), .Y(n11199));
  INVX1   g09473(.A(n11199), .Y(n11200));
  NOR2X1  g09474(.A(n10590), .B(n10140), .Y(n11201));
  AOI21X1 g09475(.A0(n11200), .A1(n10590), .B0(n11201), .Y(n11202));
  XOR2X1  g09476(.A(n11202), .B(n11191), .Y(n11203));
  INVX1   g09477(.A(n11181), .Y(n11205));
  AOI21X1 g09478(.A0(n11205), .A1(n11163), .B0(n11182), .Y(n11206));
  INVX1   g09479(.A(n11191), .Y(n11207));
  XOR2X1  g09480(.A(n11202), .B(n11207), .Y(n11208));
  NOR2X1  g09481(.A(n11208), .B(n11206), .Y(n11209));
  AOI21X1 g09482(.A0(n11206), .A1(n11208), .B0(n11209), .Y(n11210));
  NOR2X1  g09483(.A(n11210), .B(n10780), .Y(n11211));
  AOI22X1 g09484(.A0(n11140), .A1(n11145), .B0(n11102), .B1(n11095), .Y(n11212));
  AOI21X1 g09485(.A0(n11212), .A1(n11111), .B0(n11152), .Y(n11213));
  NOR2X1  g09486(.A(n11213), .B(n11151), .Y(n11214));
  NAND3X1 g09487(.A(n11062), .B(n10968), .C(n10884), .Y(n11215));
  AOI22X1 g09488(.A0(n11067), .A1(n11068), .B0(n11062), .B1(n10966), .Y(n11216));
  NAND2X1 g09489(.A(n11212), .B(n11112), .Y(n11217));
  AOI21X1 g09490(.A0(n11216), .A1(n11215), .B0(n11217), .Y(n11218));
  NOR2X1  g09491(.A(n11218), .B(n11214), .Y(n11219));
  XOR2X1  g09492(.A(n11219), .B(n11203), .Y(n11220));
  INVX1   g09493(.A(n11220), .Y(n11221));
  AOI22X1 g09494(.A0(n11131), .A1(n10680), .B0(n10628), .B1(n11221), .Y(n11222));
  OAI21X1 g09495(.A0(n10629), .A1(n10623), .B0(n11221), .Y(n11223));
  NAND2X1 g09496(.A(n11223), .B(n11222), .Y(n11224));
  NOR2X1  g09497(.A(n11210), .B(n10744), .Y(n11225));
  AOI21X1 g09498(.A0(n10766), .A1(n10618), .B0(n11210), .Y(n11229));
  NOR4X1  g09499(.A(n11225), .B(n11224), .C(n11211), .D(n11229), .Y(n11230));
  INVX1   g09500(.A(n11230), .Y(n11231));
  INVX1   g09501(.A(n11202), .Y(n11232));
  AOI22X1 g09502(.A0(n10652), .A1(P3_REG0_REG_13__SCAN_IN), .B0(P3_REG2_REG_13__SCAN_IN), .B1(n10653), .Y(n11233));
  INVX1   g09503(.A(P3_REG3_REG_13__SCAN_IN), .Y(n11234));
  NOR4X1  g09504(.A(P3_REG3_REG_11__SCAN_IN), .B(P3_REG3_REG_12__SCAN_IN), .C(P3_REG3_REG_10__SCAN_IN), .D(n11030), .Y(n11235));
  NAND3X1 g09505(.A(n11125), .B(n11234), .C(n11187), .Y(n11236));
  OAI21X1 g09506(.A0(n11235), .A1(n11234), .B0(n11236), .Y(n11237));
  AOI22X1 g09507(.A0(n10656), .A1(n11237), .B0(n10655), .B1(P3_REG1_REG_13__SCAN_IN), .Y(n11238));
  NAND2X1 g09508(.A(n11238), .B(n11233), .Y(n11239));
  AOI22X1 g09509(.A0(n11232), .A1(n10734), .B0(n10637), .B1(n11239), .Y(n11240));
  OAI21X1 g09510(.A0(n11220), .A1(n10733), .B0(n11240), .Y(n11241));
  NOR2X1  g09511(.A(n11241), .B(n11231), .Y(n11242));
  NAND2X1 g09512(.A(n10697), .B(P3_REG0_REG_12__SCAN_IN), .Y(n11243));
  OAI21X1 g09513(.A0(n11242), .A1(n10697), .B0(n11243), .Y(P3_U3426));
  NOR2X1  g09514(.A(n11202), .B(n11207), .Y(n11245));
  INVX1   g09515(.A(n11245), .Y(n11246));
  INVX1   g09516(.A(n10590), .Y(n11247));
  NOR2X1  g09517(.A(P3_IR_REG_31__SCAN_IN), .B(n10156), .Y(n11248));
  AOI21X1 g09518(.A0(n10157), .A1(P3_IR_REG_31__SCAN_IN), .B0(n11248), .Y(n11249));
  OAI21X1 g09519(.A0(n10589), .A1(n10587), .B0(n10154), .Y(n11250));
  OAI21X1 g09520(.A0(n11249), .A1(n11247), .B0(n11250), .Y(n11251));
  NOR2X1  g09521(.A(n11251), .B(n11239), .Y(n11252));
  AOI21X1 g09522(.A0(n11202), .A1(n11207), .B0(n11252), .Y(n11253));
  INVX1   g09523(.A(n11253), .Y(n11254));
  AOI21X1 g09524(.A0(n11251), .A1(n11239), .B0(n11254), .Y(n11255));
  INVX1   g09525(.A(n11255), .Y(n11256));
  AOI21X1 g09526(.A0(n11246), .A1(n11206), .B0(n11256), .Y(n11257));
  INVX1   g09527(.A(n11257), .Y(n11258));
  NOR2X1  g09528(.A(n11232), .B(n11191), .Y(n11259));
  AOI21X1 g09529(.A0(n11238), .A1(n11233), .B0(n11251), .Y(n11260));
  INVX1   g09530(.A(n11251), .Y(n11261));
  NOR2X1  g09531(.A(n11261), .B(n11239), .Y(n11262));
  NOR3X1  g09532(.A(n11262), .B(n11260), .C(n11245), .Y(n11263));
  OAI21X1 g09533(.A0(n11259), .A1(n11206), .B0(n11263), .Y(n11264));
  NAND3X1 g09534(.A(n11264), .B(n11258), .C(n10626), .Y(n11265));
  INVX1   g09535(.A(n11239), .Y(n11266));
  XOR2X1  g09536(.A(n11251), .B(n11266), .Y(n11267));
  NOR2X1  g09537(.A(n11232), .B(n11207), .Y(n11268));
  NOR4X1  g09538(.A(n11139), .B(n11050), .C(n11045), .D(n11151), .Y(n11269));
  OAI22X1 g09539(.A0(n11152), .A1(n11269), .B0(n11150), .B1(n11131), .Y(n11270));
  INVX1   g09540(.A(n11112), .Y(n11271));
  NOR3X1  g09541(.A(n11151), .B(n11139), .C(n11271), .Y(n11272));
  OAI21X1 g09542(.A0(n11070), .A1(n11064), .B0(n11272), .Y(n11273));
  AOI22X1 g09543(.A0(n11270), .A1(n11273), .B0(n11232), .B1(n11207), .Y(n11274));
  NOR2X1  g09544(.A(n11274), .B(n11268), .Y(n11275));
  XOR2X1  g09545(.A(n11275), .B(n11267), .Y(n11276));
  INVX1   g09546(.A(n11276), .Y(n11277));
  AOI22X1 g09547(.A0(n11191), .A1(n10680), .B0(n10628), .B1(n11277), .Y(n11278));
  OAI21X1 g09548(.A0(n10629), .A1(n10623), .B0(n11277), .Y(n11279));
  NAND3X1 g09549(.A(n11279), .B(n11278), .C(n11265), .Y(n11280));
  INVX1   g09550(.A(n11264), .Y(n11281));
  NOR3X1  g09551(.A(n11281), .B(n11257), .C(n10744), .Y(n11282));
  NAND2X1 g09552(.A(n11264), .B(n11258), .Y(n11286));
  AOI21X1 g09553(.A0(n10766), .A1(n10618), .B0(n11286), .Y(n11287));
  AOI22X1 g09554(.A0(n10652), .A1(P3_REG0_REG_14__SCAN_IN), .B0(P3_REG2_REG_14__SCAN_IN), .B1(n10653), .Y(n11288));
  XOR2X1  g09555(.A(n11236), .B(P3_REG3_REG_14__SCAN_IN), .Y(n11289));
  INVX1   g09556(.A(n11289), .Y(n11290));
  AOI22X1 g09557(.A0(n10656), .A1(n11290), .B0(n10655), .B1(P3_REG1_REG_14__SCAN_IN), .Y(n11291));
  NAND2X1 g09558(.A(n11291), .B(n11288), .Y(n11292));
  AOI22X1 g09559(.A0(n11251), .A1(n10734), .B0(n10637), .B1(n11292), .Y(n11293));
  OAI21X1 g09560(.A0(n11276), .A1(n10733), .B0(n11293), .Y(n11294));
  NOR4X1  g09561(.A(n11287), .B(n11282), .C(n11280), .D(n11294), .Y(n11295));
  NAND2X1 g09562(.A(n10697), .B(P3_REG0_REG_13__SCAN_IN), .Y(n11296));
  OAI21X1 g09563(.A0(n11295), .A1(n10697), .B0(n11296), .Y(P3_U3429));
  NOR2X1  g09564(.A(P3_IR_REG_31__SCAN_IN), .B(n10168), .Y(n11298));
  AOI21X1 g09565(.A0(n10172), .A1(P3_IR_REG_31__SCAN_IN), .B0(n11298), .Y(n11299));
  INVX1   g09566(.A(n11299), .Y(n11300));
  NOR2X1  g09567(.A(n10590), .B(n10167), .Y(n11301));
  AOI21X1 g09568(.A0(n11300), .A1(n10590), .B0(n11301), .Y(n11302));
  XOR2X1  g09569(.A(n11302), .B(n11292), .Y(n11303));
  NAND2X1 g09570(.A(n11253), .B(n11182), .Y(n11305));
  AOI21X1 g09571(.A0(n11251), .A1(n11239), .B0(n11245), .Y(n11306));
  AOI21X1 g09572(.A0(n11306), .A1(n11305), .B0(n11252), .Y(n11307));
  NOR2X1  g09573(.A(n11254), .B(n11181), .Y(n11308));
  AOI21X1 g09574(.A0(n11308), .A1(n11163), .B0(n11307), .Y(n11309));
  XOR2X1  g09575(.A(n11309), .B(n13411), .Y(n11310));
  XOR2X1  g09576(.A(n11309), .B(n11303), .Y(n11312));
  OAI21X1 g09577(.A0(n10625), .A1(n10617), .B0(n11312), .Y(n11313));
  OAI21X1 g09578(.A0(n11310), .A1(n10744), .B0(n11313), .Y(n11314));
  INVX1   g09579(.A(n11260), .Y(n11315));
  OAI22X1 g09580(.A0(n11261), .A1(n11239), .B0(n11268), .B1(n11274), .Y(n11316));
  NAND2X1 g09581(.A(n11316), .B(n11315), .Y(n11317));
  XOR2X1  g09582(.A(n11317), .B(n13411), .Y(n11318));
  NOR2X1  g09583(.A(n11310), .B(n10780), .Y(n11319));
  AOI21X1 g09584(.A0(n11239), .A1(n10680), .B0(n11319), .Y(n11320));
  OAI21X1 g09585(.A0(n11318), .A1(n10718), .B0(n11320), .Y(n11321));
  AOI21X1 g09586(.A0(n10729), .A1(n10728), .B0(n11318), .Y(n11322));
  INVX1   g09587(.A(n11302), .Y(n11323));
  AOI22X1 g09588(.A0(n10652), .A1(P3_REG0_REG_15__SCAN_IN), .B0(P3_REG2_REG_15__SCAN_IN), .B1(n10653), .Y(n11324));
  INVX1   g09589(.A(P3_REG3_REG_15__SCAN_IN), .Y(n11325));
  NOR2X1  g09590(.A(n11236), .B(P3_REG3_REG_14__SCAN_IN), .Y(n11326));
  NOR3X1  g09591(.A(n11236), .B(P3_REG3_REG_15__SCAN_IN), .C(P3_REG3_REG_14__SCAN_IN), .Y(n11327));
  INVX1   g09592(.A(n11327), .Y(n11328));
  OAI21X1 g09593(.A0(n11326), .A1(n11325), .B0(n11328), .Y(n11329));
  AOI22X1 g09594(.A0(n10656), .A1(n11329), .B0(n10655), .B1(P3_REG1_REG_15__SCAN_IN), .Y(n11330));
  NAND2X1 g09595(.A(n11330), .B(n11324), .Y(n11331));
  AOI22X1 g09596(.A0(n11323), .A1(n10734), .B0(n10637), .B1(n11331), .Y(n11332));
  OAI21X1 g09597(.A0(n11318), .A1(n10733), .B0(n11332), .Y(n11333));
  NOR4X1  g09598(.A(n11322), .B(n11321), .C(n11314), .D(n11333), .Y(n11334));
  NAND2X1 g09599(.A(n10697), .B(P3_REG0_REG_14__SCAN_IN), .Y(n11335));
  OAI21X1 g09600(.A0(n11334), .A1(n10697), .B0(n11335), .Y(P3_U3432));
  INVX1   g09601(.A(n11331), .Y(n11337));
  NOR2X1  g09602(.A(P3_IR_REG_31__SCAN_IN), .B(n10183), .Y(n11338));
  AOI21X1 g09603(.A0(n10184), .A1(P3_IR_REG_31__SCAN_IN), .B0(n11338), .Y(n11339));
  INVX1   g09604(.A(n11339), .Y(n11340));
  NAND2X1 g09605(.A(n11340), .B(n10590), .Y(n11341));
  OAI21X1 g09606(.A0(n10590), .A1(n10182), .B0(n11341), .Y(n11342));
  XOR2X1  g09607(.A(n11342), .B(n11337), .Y(n11343));
  INVX1   g09608(.A(n11292), .Y(n11344));
  NOR2X1  g09609(.A(n11302), .B(n11344), .Y(n11345));
  INVX1   g09610(.A(n11345), .Y(n11346));
  NOR2X1  g09611(.A(n11323), .B(n11292), .Y(n11347));
  OAI21X1 g09612(.A0(n11347), .A1(n11309), .B0(n11346), .Y(n11348));
  XOR2X1  g09613(.A(n11348), .B(n11343), .Y(n11349));
  INVX1   g09614(.A(n11348), .Y(n11351));
  XOR2X1  g09615(.A(n11351), .B(n11343), .Y(n11352));
  OAI21X1 g09616(.A0(n10625), .A1(n10617), .B0(n11352), .Y(n11353));
  OAI21X1 g09617(.A0(n11349), .A1(n10744), .B0(n11353), .Y(n11354));
  NOR2X1  g09618(.A(n11323), .B(n11344), .Y(n11355));
  NOR2X1  g09619(.A(n11302), .B(n11292), .Y(n11356));
  INVX1   g09620(.A(n11356), .Y(n11357));
  AOI21X1 g09621(.A0(n11317), .A1(n11357), .B0(n11355), .Y(n11358));
  XOR2X1  g09622(.A(n11358), .B(n11343), .Y(n11359));
  NOR2X1  g09623(.A(n11349), .B(n10780), .Y(n11360));
  AOI21X1 g09624(.A0(n11292), .A1(n10680), .B0(n11360), .Y(n11361));
  OAI21X1 g09625(.A0(n11359), .A1(n10718), .B0(n11361), .Y(n11362));
  AOI21X1 g09626(.A0(n10729), .A1(n10728), .B0(n11359), .Y(n11363));
  AOI22X1 g09627(.A0(n10652), .A1(P3_REG0_REG_16__SCAN_IN), .B0(P3_REG2_REG_16__SCAN_IN), .B1(n10653), .Y(n11364));
  INVX1   g09628(.A(P3_REG3_REG_16__SCAN_IN), .Y(n11365));
  XOR2X1  g09629(.A(n11327), .B(n11365), .Y(n11366));
  INVX1   g09630(.A(n11366), .Y(n11367));
  AOI22X1 g09631(.A0(n10656), .A1(n11367), .B0(n10655), .B1(P3_REG1_REG_16__SCAN_IN), .Y(n11368));
  NAND2X1 g09632(.A(n11368), .B(n11364), .Y(n11369));
  AOI22X1 g09633(.A0(n11342), .A1(n10734), .B0(n10637), .B1(n11369), .Y(n11370));
  OAI21X1 g09634(.A0(n11359), .A1(n10733), .B0(n11370), .Y(n11371));
  NOR4X1  g09635(.A(n11363), .B(n11362), .C(n11354), .D(n11371), .Y(n11372));
  NAND2X1 g09636(.A(n10697), .B(P3_REG0_REG_15__SCAN_IN), .Y(n11373));
  OAI21X1 g09637(.A0(n11372), .A1(n10697), .B0(n11373), .Y(P3_U3435));
  NOR2X1  g09638(.A(n11342), .B(n11337), .Y(n11375));
  INVX1   g09639(.A(n11358), .Y(n11376));
  INVX1   g09640(.A(n11369), .Y(n11377));
  NOR2X1  g09641(.A(P3_IR_REG_31__SCAN_IN), .B(n10195), .Y(n11378));
  AOI21X1 g09642(.A0(n10206), .A1(P3_IR_REG_31__SCAN_IN), .B0(n11378), .Y(n11379));
  INVX1   g09643(.A(n11379), .Y(n11380));
  NAND2X1 g09644(.A(n11380), .B(n10590), .Y(n11381));
  OAI21X1 g09645(.A0(n10590), .A1(n10194), .B0(n11381), .Y(n11382));
  XOR2X1  g09646(.A(n11382), .B(n11377), .Y(n11383));
  AOI21X1 g09647(.A0(n11342), .A1(n11337), .B0(n11383), .Y(n11384));
  OAI21X1 g09648(.A0(n11376), .A1(n11375), .B0(n11384), .Y(n11385));
  NAND2X1 g09649(.A(n11342), .B(n11337), .Y(n11386));
  INVX1   g09650(.A(n11386), .Y(n11387));
  NAND2X1 g09651(.A(n11382), .B(n11377), .Y(n11388));
  INVX1   g09652(.A(n11388), .Y(n11389));
  INVX1   g09653(.A(n11342), .Y(n11390));
  INVX1   g09654(.A(n11382), .Y(n11391));
  AOI22X1 g09655(.A0(n11369), .A1(n11391), .B0(n11390), .B1(n11331), .Y(n11392));
  INVX1   g09656(.A(n11392), .Y(n11393));
  NOR2X1  g09657(.A(n11393), .B(n11389), .Y(n11394));
  OAI21X1 g09658(.A0(n11358), .A1(n11387), .B0(n11394), .Y(n11395));
  NAND2X1 g09659(.A(n11395), .B(n11385), .Y(n11396));
  OAI21X1 g09660(.A0(n10629), .A1(n10623), .B0(n11396), .Y(n11397));
  NOR2X1  g09661(.A(n11390), .B(n11337), .Y(n11398));
  NOR2X1  g09662(.A(n11342), .B(n11331), .Y(n11399));
  INVX1   g09663(.A(n11399), .Y(n11400));
  AOI21X1 g09664(.A0(n11400), .A1(n11348), .B0(n11398), .Y(n11401));
  INVX1   g09665(.A(n11401), .Y(n11402));
  NOR2X1  g09666(.A(n11402), .B(n11383), .Y(n11403));
  XOR2X1  g09667(.A(n11382), .B(n11369), .Y(n11404));
  NOR2X1  g09668(.A(n11404), .B(n11401), .Y(n11405));
  OAI21X1 g09669(.A0(n11405), .A1(n11403), .B0(n10622), .Y(n11406));
  NAND2X1 g09670(.A(n11396), .B(n10628), .Y(n11407));
  NAND3X1 g09671(.A(n11407), .B(n11406), .C(n11397), .Y(n11408));
  OAI21X1 g09672(.A0(n11405), .A1(n11403), .B0(n10626), .Y(n11409));
  OAI21X1 g09673(.A0(n11337), .A1(n10781), .B0(n11409), .Y(n11410));
  AOI21X1 g09674(.A0(n11401), .A1(n11404), .B0(n11405), .Y(n11414));
  AOI21X1 g09675(.A0(n10766), .A1(n10618), .B0(n11414), .Y(n11415));
  NAND2X1 g09676(.A(n11396), .B(n10633), .Y(n11416));
  AOI22X1 g09677(.A0(n10652), .A1(P3_REG0_REG_17__SCAN_IN), .B0(P3_REG2_REG_17__SCAN_IN), .B1(n10653), .Y(n11417));
  INVX1   g09678(.A(P3_REG3_REG_17__SCAN_IN), .Y(n11418));
  NOR4X1  g09679(.A(P3_REG3_REG_15__SCAN_IN), .B(P3_REG3_REG_16__SCAN_IN), .C(P3_REG3_REG_14__SCAN_IN), .D(n11236), .Y(n11419));
  NOR3X1  g09680(.A(n11328), .B(P3_REG3_REG_17__SCAN_IN), .C(P3_REG3_REG_16__SCAN_IN), .Y(n11420));
  INVX1   g09681(.A(n11420), .Y(n11421));
  OAI21X1 g09682(.A0(n11419), .A1(n11418), .B0(n11421), .Y(n11422));
  AOI22X1 g09683(.A0(n10656), .A1(n11422), .B0(n10655), .B1(P3_REG1_REG_17__SCAN_IN), .Y(n11423));
  NAND2X1 g09684(.A(n11423), .B(n11417), .Y(n11424));
  AOI22X1 g09685(.A0(n11382), .A1(n10734), .B0(n10637), .B1(n11424), .Y(n11425));
  NAND2X1 g09686(.A(n11425), .B(n11416), .Y(n11426));
  NOR4X1  g09687(.A(n11415), .B(n11410), .C(n11408), .D(n11426), .Y(n11427));
  NAND2X1 g09688(.A(n10697), .B(P3_REG0_REG_16__SCAN_IN), .Y(n11428));
  OAI21X1 g09689(.A0(n11427), .A1(n10697), .B0(n11428), .Y(P3_U3438));
  NAND2X1 g09690(.A(n11382), .B(n11369), .Y(n11430));
  NOR2X1  g09691(.A(P3_IR_REG_31__SCAN_IN), .B(n10217), .Y(n11431));
  AOI21X1 g09692(.A0(n10218), .A1(P3_IR_REG_31__SCAN_IN), .B0(n11431), .Y(n11432));
  INVX1   g09693(.A(n11432), .Y(n11433));
  NOR2X1  g09694(.A(n10590), .B(n10216), .Y(n11434));
  AOI21X1 g09695(.A0(n11433), .A1(n10590), .B0(n11434), .Y(n11435));
  INVX1   g09696(.A(n11435), .Y(n11436));
  NOR2X1  g09697(.A(n11382), .B(n11369), .Y(n11437));
  INVX1   g09698(.A(n11437), .Y(n11438));
  OAI21X1 g09699(.A0(n11436), .A1(n11424), .B0(n11438), .Y(n11439));
  AOI21X1 g09700(.A0(n11436), .A1(n11424), .B0(n11439), .Y(n11440));
  INVX1   g09701(.A(n11440), .Y(n11441));
  AOI21X1 g09702(.A0(n11430), .A1(n11401), .B0(n11441), .Y(n11442));
  INVX1   g09703(.A(n11430), .Y(n11443));
  XOR2X1  g09704(.A(n11435), .B(n11424), .Y(n11444));
  NOR2X1  g09705(.A(n13405), .B(n11443), .Y(n11446));
  INVX1   g09706(.A(n11446), .Y(n11447));
  AOI21X1 g09707(.A0(n11438), .A1(n11402), .B0(n11447), .Y(n11448));
  NOR2X1  g09708(.A(n11448), .B(n11442), .Y(n11449));
  NAND2X1 g09709(.A(n11449), .B(n10626), .Y(n11450));
  NAND3X1 g09710(.A(n11388), .B(n11386), .C(n11355), .Y(n11451));
  AOI21X1 g09711(.A0(n11451), .A1(n11392), .B0(n11389), .Y(n11452));
  NOR3X1  g09712(.A(n11389), .B(n11387), .C(n11356), .Y(n11453));
  INVX1   g09713(.A(n11453), .Y(n11454));
  AOI21X1 g09714(.A0(n11316), .A1(n11315), .B0(n11454), .Y(n11455));
  NOR2X1  g09715(.A(n11455), .B(n11452), .Y(n11456));
  XOR2X1  g09716(.A(n11456), .B(n11444), .Y(n11457));
  INVX1   g09717(.A(n11457), .Y(n11458));
  AOI22X1 g09718(.A0(n11369), .A1(n10680), .B0(n10628), .B1(n11458), .Y(n11459));
  OAI21X1 g09719(.A0(n10629), .A1(n10623), .B0(n11458), .Y(n11460));
  NAND3X1 g09720(.A(n11460), .B(n11459), .C(n11450), .Y(n11461));
  NOR3X1  g09721(.A(n11448), .B(n11442), .C(n10744), .Y(n11462));
  NAND2X1 g09722(.A(n11401), .B(n11430), .Y(n11463));
  NAND2X1 g09723(.A(n11463), .B(n11440), .Y(n11464));
  OAI21X1 g09724(.A0(n11401), .A1(n11437), .B0(n11446), .Y(n11465));
  NAND2X1 g09725(.A(n11465), .B(n11464), .Y(n11466));
  AOI21X1 g09726(.A0(n10766), .A1(n10618), .B0(n11466), .Y(n11467));
  AOI22X1 g09727(.A0(n10652), .A1(P3_REG0_REG_18__SCAN_IN), .B0(P3_REG2_REG_18__SCAN_IN), .B1(n10653), .Y(n11468));
  INVX1   g09728(.A(P3_REG3_REG_18__SCAN_IN), .Y(n11469));
  XOR2X1  g09729(.A(n11420), .B(n11469), .Y(n11470));
  INVX1   g09730(.A(n11470), .Y(n11471));
  AOI22X1 g09731(.A0(n10656), .A1(n11471), .B0(n10655), .B1(P3_REG1_REG_18__SCAN_IN), .Y(n11472));
  NAND2X1 g09732(.A(n11472), .B(n11468), .Y(n11473));
  AOI22X1 g09733(.A0(n11436), .A1(n10734), .B0(n10637), .B1(n11473), .Y(n11474));
  OAI21X1 g09734(.A0(n11457), .A1(n10733), .B0(n11474), .Y(n11475));
  NOR4X1  g09735(.A(n11467), .B(n11462), .C(n11461), .D(n11475), .Y(n11476));
  NAND2X1 g09736(.A(n10697), .B(P3_REG0_REG_17__SCAN_IN), .Y(n11477));
  OAI21X1 g09737(.A0(n11476), .A1(n10697), .B0(n11477), .Y(P3_U3441));
  NOR2X1  g09738(.A(P3_IR_REG_31__SCAN_IN), .B(n10229), .Y(n11479));
  AOI21X1 g09739(.A0(n10233), .A1(P3_IR_REG_31__SCAN_IN), .B0(n11479), .Y(n11480));
  INVX1   g09740(.A(n11480), .Y(n11481));
  NOR2X1  g09741(.A(n10590), .B(n10228), .Y(n11482));
  AOI21X1 g09742(.A0(n11481), .A1(n10590), .B0(n11482), .Y(n11483));
  XOR2X1  g09743(.A(n11483), .B(n11473), .Y(n11484));
  INVX1   g09744(.A(n11424), .Y(n11485));
  NOR2X1  g09745(.A(n11436), .B(n11485), .Y(n11486));
  INVX1   g09746(.A(n11486), .Y(n11487));
  OAI22X1 g09747(.A0(n11452), .A1(n11455), .B0(n11435), .B1(n11424), .Y(n11488));
  NAND2X1 g09748(.A(n11488), .B(n11487), .Y(n11489));
  XOR2X1  g09749(.A(n11489), .B(n11484), .Y(n11490));
  AOI22X1 g09750(.A0(n11424), .A1(n10680), .B0(n10628), .B1(n11490), .Y(n11491));
  OAI21X1 g09751(.A0(n10629), .A1(n10623), .B0(n11490), .Y(n11492));
  NAND2X1 g09752(.A(n11492), .B(n11491), .Y(n11493));
  AOI21X1 g09753(.A0(n11435), .A1(n11430), .B0(n11485), .Y(n11494));
  AOI21X1 g09754(.A0(n11436), .A1(n11443), .B0(n11494), .Y(n11495));
  OAI21X1 g09755(.A0(n11439), .A1(n11401), .B0(n11495), .Y(n11496));
  NOR2X1  g09756(.A(n11496), .B(n11484), .Y(n11497));
  INVX1   g09757(.A(n11473), .Y(n11498));
  XOR2X1  g09758(.A(n11483), .B(n11498), .Y(n11499));
  AOI21X1 g09759(.A0(n11484), .A1(n11496), .B0(n11497), .Y(n11501));
  OAI22X1 g09760(.A0(n11501), .A1(n10780), .B0(n10766), .B1(n11501), .Y(n11505));
  OAI22X1 g09761(.A0(n11501), .A1(n10744), .B0(n10618), .B1(n11501), .Y(n11506));
  NAND2X1 g09762(.A(n11490), .B(n10633), .Y(n11507));
  INVX1   g09763(.A(n11483), .Y(n11508));
  AOI22X1 g09764(.A0(n10652), .A1(P3_REG0_REG_19__SCAN_IN), .B0(P3_REG2_REG_19__SCAN_IN), .B1(n10653), .Y(n11509));
  INVX1   g09765(.A(P3_REG3_REG_19__SCAN_IN), .Y(n11510));
  NOR4X1  g09766(.A(P3_REG3_REG_18__SCAN_IN), .B(P3_REG3_REG_17__SCAN_IN), .C(P3_REG3_REG_16__SCAN_IN), .D(n11328), .Y(n11511));
  NAND3X1 g09767(.A(n11420), .B(n11469), .C(n11510), .Y(n11512));
  OAI21X1 g09768(.A0(n11511), .A1(n11510), .B0(n11512), .Y(n11513));
  AOI22X1 g09769(.A0(n10656), .A1(n11513), .B0(n10655), .B1(P3_REG1_REG_19__SCAN_IN), .Y(n11514));
  NAND2X1 g09770(.A(n11514), .B(n11509), .Y(n11515));
  AOI22X1 g09771(.A0(n11508), .A1(n10734), .B0(n10637), .B1(n11515), .Y(n11516));
  NAND2X1 g09772(.A(n11516), .B(n11507), .Y(n11517));
  NOR4X1  g09773(.A(n11506), .B(n11505), .C(n11493), .D(n11517), .Y(n11518));
  NAND2X1 g09774(.A(n10697), .B(P3_REG0_REG_18__SCAN_IN), .Y(n11519));
  OAI21X1 g09775(.A0(n11518), .A1(n10697), .B0(n11519), .Y(P3_U3444));
  INVX1   g09776(.A(n11515), .Y(n11521));
  OAI21X1 g09777(.A0(n10243), .A1(n10236), .B0(n11247), .Y(n11522));
  OAI21X1 g09778(.A0(n11247), .A1(n10571), .B0(n11522), .Y(n11523));
  XOR2X1  g09779(.A(n11523), .B(n11521), .Y(n11524));
  NOR2X1  g09780(.A(n11508), .B(n11498), .Y(n11525));
  AOI21X1 g09781(.A0(n11488), .A1(n11487), .B0(n11498), .Y(n11526));
  AOI21X1 g09782(.A0(n11488), .A1(n11487), .B0(n11508), .Y(n11527));
  NOR3X1  g09783(.A(n11527), .B(n11526), .C(n11525), .Y(n11528));
  XOR2X1  g09784(.A(n11528), .B(n11524), .Y(n11529));
  INVX1   g09785(.A(n11529), .Y(n11530));
  OAI21X1 g09786(.A0(n10629), .A1(n10623), .B0(n11530), .Y(n11531));
  INVX1   g09787(.A(n11531), .Y(n11532));
  INVX1   g09788(.A(n11524), .Y(n11533));
  NOR2X1  g09789(.A(n11508), .B(n11473), .Y(n11534));
  INVX1   g09790(.A(n11534), .Y(n11535));
  NOR2X1  g09791(.A(n11483), .B(n11498), .Y(n11536));
  AOI21X1 g09792(.A0(n11535), .A1(n11496), .B0(n11536), .Y(n11537));
  NOR2X1  g09793(.A(n11533), .B(n11537), .Y(n11540));
  AOI21X1 g09794(.A0(n11537), .A1(n11533), .B0(n11540), .Y(n11541));
  OAI22X1 g09795(.A0(n11529), .A1(n10728), .B0(n10744), .B1(n11541), .Y(n11542));
  OAI22X1 g09796(.A0(n11498), .A1(n10781), .B0(n10780), .B1(n11541), .Y(n11543));
  AOI21X1 g09797(.A0(n10766), .A1(n10618), .B0(n11541), .Y(n11547));
  NOR4X1  g09798(.A(n11543), .B(n11542), .C(n11532), .D(n11547), .Y(n11548));
  INVX1   g09799(.A(n11548), .Y(n11549));
  AOI22X1 g09800(.A0(n10652), .A1(P3_REG0_REG_20__SCAN_IN), .B0(P3_REG2_REG_20__SCAN_IN), .B1(n10653), .Y(n11550));
  XOR2X1  g09801(.A(n11512), .B(P3_REG3_REG_20__SCAN_IN), .Y(n11551));
  INVX1   g09802(.A(n11551), .Y(n11552));
  AOI22X1 g09803(.A0(n10656), .A1(n11552), .B0(n10655), .B1(P3_REG1_REG_20__SCAN_IN), .Y(n11553));
  NAND2X1 g09804(.A(n11553), .B(n11550), .Y(n11554));
  AOI22X1 g09805(.A0(n11523), .A1(n10734), .B0(n10637), .B1(n11554), .Y(n11555));
  OAI21X1 g09806(.A0(n11529), .A1(n10733), .B0(n11555), .Y(n11556));
  NOR2X1  g09807(.A(n11556), .B(n11549), .Y(n11557));
  NAND2X1 g09808(.A(n10697), .B(P3_REG0_REG_19__SCAN_IN), .Y(n11558));
  OAI21X1 g09809(.A0(n11557), .A1(n10697), .B0(n11558), .Y(P3_U3446));
  NOR2X1  g09810(.A(n10590), .B(n10255), .Y(n11560));
  NOR2X1  g09811(.A(n11523), .B(n11515), .Y(n11561));
  INVX1   g09812(.A(n11554), .Y(n11562));
  INVX1   g09813(.A(n11560), .Y(n11563));
  AOI21X1 g09814(.A0(n11563), .A1(n11562), .B0(n11561), .Y(n11564));
  INVX1   g09815(.A(n11564), .Y(n11565));
  AOI21X1 g09816(.A0(n11560), .A1(n11554), .B0(n11565), .Y(n11566));
  NAND2X1 g09817(.A(n11523), .B(n11515), .Y(n11567));
  NAND2X1 g09818(.A(n11567), .B(n11537), .Y(n11568));
  INVX1   g09819(.A(n11567), .Y(n11569));
  XOR2X1  g09820(.A(n11560), .B(n11562), .Y(n11570));
  INVX1   g09821(.A(n11570), .Y(n11571));
  NOR2X1  g09822(.A(n11561), .B(n11537), .Y(n11572));
  NOR3X1  g09823(.A(n11572), .B(n11571), .C(n11569), .Y(n11573));
  AOI21X1 g09824(.A0(n11568), .A1(n11566), .B0(n11573), .Y(n11574));
  NAND2X1 g09825(.A(n11574), .B(n10622), .Y(n11575));
  INVX1   g09826(.A(n11537), .Y(n11576));
  OAI21X1 g09827(.A0(n11576), .A1(n11569), .B0(n11566), .Y(n11577));
  NOR2X1  g09828(.A(n11571), .B(n11569), .Y(n11578));
  OAI21X1 g09829(.A0(n11537), .A1(n11561), .B0(n11578), .Y(n11579));
  NAND3X1 g09830(.A(n11579), .B(n11577), .C(n10625), .Y(n11580));
  NAND3X1 g09831(.A(n11579), .B(n11577), .C(n10617), .Y(n11581));
  NAND3X1 g09832(.A(n11581), .B(n11580), .C(n11575), .Y(n11582));
  NOR2X1  g09833(.A(n11523), .B(n11521), .Y(n11583));
  INVX1   g09834(.A(n11583), .Y(n11584));
  INVX1   g09835(.A(n11523), .Y(n11585));
  NOR2X1  g09836(.A(n11585), .B(n11515), .Y(n11586));
  OAI21X1 g09837(.A0(n11528), .A1(n11586), .B0(n11584), .Y(n11587));
  XOR2X1  g09838(.A(n11587), .B(n11571), .Y(n11588));
  NOR2X1  g09839(.A(n11588), .B(n10718), .Y(n11589));
  INVX1   g09840(.A(n11589), .Y(n11590));
  AOI22X1 g09841(.A0(n11515), .A1(n10680), .B0(n10626), .B1(n11574), .Y(n11591));
  INVX1   g09842(.A(n11588), .Y(n11592));
  OAI21X1 g09843(.A0(n10629), .A1(n10628), .B0(n11592), .Y(n11593));
  NAND3X1 g09844(.A(n11593), .B(n11591), .C(n11590), .Y(n11594));
  AOI22X1 g09845(.A0(n10652), .A1(P3_REG0_REG_21__SCAN_IN), .B0(P3_REG2_REG_21__SCAN_IN), .B1(n10653), .Y(n11595));
  NOR3X1  g09846(.A(n11512), .B(P3_REG3_REG_20__SCAN_IN), .C(P3_REG3_REG_21__SCAN_IN), .Y(n11596));
  INVX1   g09847(.A(n11596), .Y(n11597));
  OAI21X1 g09848(.A0(n11512), .A1(P3_REG3_REG_20__SCAN_IN), .B0(P3_REG3_REG_21__SCAN_IN), .Y(n11598));
  NAND2X1 g09849(.A(n11598), .B(n11597), .Y(n11599));
  AOI22X1 g09850(.A0(n10656), .A1(n11599), .B0(n10655), .B1(P3_REG1_REG_21__SCAN_IN), .Y(n11600));
  NAND2X1 g09851(.A(n11600), .B(n11595), .Y(n11601));
  AOI22X1 g09852(.A0(n11560), .A1(n10734), .B0(n10637), .B1(n11601), .Y(n11602));
  OAI21X1 g09853(.A0(n11588), .A1(n10733), .B0(n11602), .Y(n11603));
  NOR3X1  g09854(.A(n11603), .B(n11594), .C(n11582), .Y(n11604));
  NAND2X1 g09855(.A(n10697), .B(P3_REG0_REG_20__SCAN_IN), .Y(n11605));
  OAI21X1 g09856(.A0(n11604), .A1(n10697), .B0(n11605), .Y(P3_U3447));
  INVX1   g09857(.A(n11601), .Y(n11607));
  NOR2X1  g09858(.A(n10590), .B(n10271), .Y(n11608));
  XOR2X1  g09859(.A(n11608), .B(n11607), .Y(n11609));
  INVX1   g09860(.A(n11609), .Y(n11610));
  NAND2X1 g09861(.A(n11563), .B(n11567), .Y(n11611));
  OAI21X1 g09862(.A0(n11563), .A1(n11567), .B0(n11562), .Y(n11612));
  NAND2X1 g09863(.A(n11612), .B(n11611), .Y(n11613));
  OAI21X1 g09864(.A0(n11565), .A1(n11537), .B0(n11613), .Y(n11614));
  NOR2X1  g09865(.A(n11565), .B(n11537), .Y(n11615));
  NAND2X1 g09866(.A(n11613), .B(n11609), .Y(n11616));
  NOR2X1  g09867(.A(n11616), .B(n11615), .Y(n11617));
  AOI21X1 g09868(.A0(n11614), .A1(n11610), .B0(n11617), .Y(n11618));
  AOI22X1 g09869(.A0(n11554), .A1(n10680), .B0(n10626), .B1(n11618), .Y(n11619));
  NAND2X1 g09870(.A(n11618), .B(n10622), .Y(n11620));
  OAI21X1 g09871(.A0(n10625), .A1(n10617), .B0(n11618), .Y(n11624));
  NOR2X1  g09872(.A(n11560), .B(n11562), .Y(n11625));
  NOR3X1  g09873(.A(n11554), .B(n10590), .C(n10255), .Y(n11626));
  INVX1   g09874(.A(n11626), .Y(n11627));
  AOI21X1 g09875(.A0(n11587), .A1(n11627), .B0(n11625), .Y(n11628));
  XOR2X1  g09876(.A(n11628), .B(n11609), .Y(n11629));
  NOR2X1  g09877(.A(n11629), .B(n10729), .Y(n11630));
  AOI21X1 g09878(.A0(n10728), .A1(n10718), .B0(n11629), .Y(n11631));
  NOR2X1  g09879(.A(n11631), .B(n11630), .Y(n11632));
  NAND4X1 g09880(.A(n11624), .B(n11620), .C(n11619), .D(n11632), .Y(n11633));
  AOI22X1 g09881(.A0(n10652), .A1(P3_REG0_REG_22__SCAN_IN), .B0(P3_REG2_REG_22__SCAN_IN), .B1(n10653), .Y(n11634));
  INVX1   g09882(.A(P3_REG3_REG_22__SCAN_IN), .Y(n11635));
  XOR2X1  g09883(.A(n11596), .B(n11635), .Y(n11636));
  INVX1   g09884(.A(n11636), .Y(n11637));
  AOI22X1 g09885(.A0(n10656), .A1(n11637), .B0(n10655), .B1(P3_REG1_REG_22__SCAN_IN), .Y(n11638));
  NAND2X1 g09886(.A(n11638), .B(n11634), .Y(n11639));
  AOI22X1 g09887(.A0(n11608), .A1(n10734), .B0(n10637), .B1(n11639), .Y(n11640));
  OAI21X1 g09888(.A0(n11629), .A1(n10733), .B0(n11640), .Y(n11641));
  NOR2X1  g09889(.A(n11641), .B(n11633), .Y(n11642));
  NAND2X1 g09890(.A(n10697), .B(P3_REG0_REG_21__SCAN_IN), .Y(n11643));
  OAI21X1 g09891(.A0(n11642), .A1(n10697), .B0(n11643), .Y(P3_U3448));
  INVX1   g09892(.A(n11639), .Y(n11645));
  NOR2X1  g09893(.A(n10590), .B(n10282), .Y(n11646));
  XOR2X1  g09894(.A(n11646), .B(n11645), .Y(n11647));
  NOR2X1  g09895(.A(n11608), .B(n11607), .Y(n11648));
  NOR3X1  g09896(.A(n11601), .B(n10590), .C(n10271), .Y(n11649));
  INVX1   g09897(.A(n11649), .Y(n11650));
  INVX1   g09898(.A(n11625), .Y(n11651));
  INVX1   g09899(.A(n11586), .Y(n11652));
  INVX1   g09900(.A(n11525), .Y(n11653));
  INVX1   g09901(.A(n11452), .Y(n11654));
  INVX1   g09902(.A(n11268), .Y(n11655));
  OAI22X1 g09903(.A0(n11214), .A1(n11218), .B0(n11202), .B1(n11191), .Y(n11656));
  AOI21X1 g09904(.A0(n11656), .A1(n11655), .B0(n11262), .Y(n11657));
  OAI21X1 g09905(.A0(n11657), .A1(n11260), .B0(n11453), .Y(n11658));
  AOI22X1 g09906(.A0(n11654), .A1(n11658), .B0(n11436), .B1(n11485), .Y(n11659));
  OAI21X1 g09907(.A0(n11659), .A1(n11486), .B0(n11473), .Y(n11660));
  OAI21X1 g09908(.A0(n11659), .A1(n11486), .B0(n11483), .Y(n11661));
  NAND3X1 g09909(.A(n11661), .B(n11660), .C(n11653), .Y(n11662));
  AOI21X1 g09910(.A0(n11662), .A1(n11652), .B0(n11583), .Y(n11663));
  OAI21X1 g09911(.A0(n11663), .A1(n11626), .B0(n11651), .Y(n11664));
  AOI21X1 g09912(.A0(n11664), .A1(n11650), .B0(n11648), .Y(n11665));
  XOR2X1  g09913(.A(n11665), .B(n11647), .Y(n11666));
  INVX1   g09914(.A(n11666), .Y(n11667));
  NOR2X1  g09915(.A(n11608), .B(n11601), .Y(n11668));
  AOI22X1 g09916(.A0(n11611), .A1(n11612), .B0(n11564), .B1(n11536), .Y(n11669));
  NOR3X1  g09917(.A(n11607), .B(n10590), .C(n10271), .Y(n11670));
  INVX1   g09918(.A(n11670), .Y(n11671));
  OAI21X1 g09919(.A0(n11669), .A1(n11668), .B0(n11671), .Y(n11672));
  NOR3X1  g09920(.A(n11668), .B(n11565), .C(n11534), .Y(n11673));
  AOI21X1 g09921(.A0(n11673), .A1(n11496), .B0(n11672), .Y(n11674));
  XOR2X1  g09922(.A(n11674), .B(n11647), .Y(n11675));
  AOI22X1 g09923(.A0(n11601), .A1(n10680), .B0(n10626), .B1(n11675), .Y(n11676));
  NAND2X1 g09924(.A(n11675), .B(n10622), .Y(n11677));
  OAI21X1 g09925(.A0(n10625), .A1(n10617), .B0(n11675), .Y(n11680));
  NAND3X1 g09926(.A(n11680), .B(n11677), .C(n11676), .Y(n11681));
  AOI21X1 g09927(.A0(n11667), .A1(n10623), .B0(n11681), .Y(n11682));
  OAI21X1 g09928(.A0(n10629), .A1(n10628), .B0(n11667), .Y(n11683));
  NAND2X1 g09929(.A(n11683), .B(n11682), .Y(n11684));
  AOI22X1 g09930(.A0(n10652), .A1(P3_REG0_REG_23__SCAN_IN), .B0(P3_REG2_REG_23__SCAN_IN), .B1(n10653), .Y(n11685));
  NAND3X1 g09931(.A(n10611), .B(n10599), .C(P3_REG1_REG_23__SCAN_IN), .Y(n11686));
  NOR3X1  g09932(.A(n11597), .B(P3_REG3_REG_22__SCAN_IN), .C(P3_REG3_REG_23__SCAN_IN), .Y(n11687));
  INVX1   g09933(.A(P3_REG3_REG_23__SCAN_IN), .Y(n11688));
  AOI21X1 g09934(.A0(n11596), .A1(n11635), .B0(n11688), .Y(n11689));
  OAI21X1 g09935(.A0(n11689), .A1(n11687), .B0(n10656), .Y(n11690));
  NAND3X1 g09936(.A(n11690), .B(n11686), .C(n11685), .Y(n11691));
  AOI22X1 g09937(.A0(n11646), .A1(n10734), .B0(n10637), .B1(n11691), .Y(n11692));
  OAI21X1 g09938(.A0(n11666), .A1(n10733), .B0(n11692), .Y(n11693));
  NOR2X1  g09939(.A(n11693), .B(n11684), .Y(n11694));
  NAND2X1 g09940(.A(n10697), .B(P3_REG0_REG_22__SCAN_IN), .Y(n11695));
  OAI21X1 g09941(.A0(n11694), .A1(n10697), .B0(n11695), .Y(P3_U3449));
  OAI21X1 g09942(.A0(n11646), .A1(n11645), .B0(n11665), .Y(n11697));
  NOR3X1  g09943(.A(n11639), .B(n10590), .C(n10282), .Y(n11698));
  OAI21X1 g09944(.A0(n10297), .A1(n10290), .B0(n11247), .Y(n11699));
  XOR2X1  g09945(.A(n11699), .B(n11691), .Y(n11700));
  NOR2X1  g09946(.A(n11700), .B(n11698), .Y(n11701));
  NAND2X1 g09947(.A(n11701), .B(n11697), .Y(n11702));
  NOR2X1  g09948(.A(n11699), .B(n11691), .Y(n11703));
  INVX1   g09949(.A(n11646), .Y(n11704));
  AOI22X1 g09950(.A0(n11691), .A1(n11699), .B0(n11704), .B1(n11639), .Y(n11705));
  INVX1   g09951(.A(n11705), .Y(n11706));
  NOR2X1  g09952(.A(n11706), .B(n11703), .Y(n11707));
  OAI21X1 g09953(.A0(n11665), .A1(n11698), .B0(n11707), .Y(n11708));
  NAND2X1 g09954(.A(n11708), .B(n11702), .Y(n11709));
  NAND2X1 g09955(.A(n11709), .B(n10623), .Y(n11710));
  NOR3X1  g09956(.A(n11645), .B(n10590), .C(n10282), .Y(n11711));
  INVX1   g09957(.A(n11711), .Y(n11712));
  NOR2X1  g09958(.A(n11646), .B(n11639), .Y(n11713));
  OAI21X1 g09959(.A0(n11713), .A1(n11674), .B0(n11712), .Y(n11714));
  XOR2X1  g09960(.A(n11714), .B(n11700), .Y(n11715));
  INVX1   g09961(.A(n11715), .Y(n11716));
  AOI22X1 g09962(.A0(n11639), .A1(n10680), .B0(n10626), .B1(n11716), .Y(n11717));
  AOI21X1 g09963(.A0(n10766), .A1(n10618), .B0(n11715), .Y(n11720));
  AOI21X1 g09964(.A0(n11716), .A1(n10622), .B0(n11720), .Y(n11721));
  NAND3X1 g09965(.A(n11721), .B(n11717), .C(n11710), .Y(n11722));
  AOI22X1 g09966(.A0(n11702), .A1(n11708), .B0(n10729), .B1(n10728), .Y(n11723));
  AOI21X1 g09967(.A0(n11708), .A1(n11702), .B0(n10733), .Y(n11724));
  AOI22X1 g09968(.A0(n10652), .A1(P3_REG0_REG_24__SCAN_IN), .B0(P3_REG2_REG_24__SCAN_IN), .B1(n10653), .Y(n11725));
  INVX1   g09969(.A(P3_REG3_REG_24__SCAN_IN), .Y(n11726));
  XOR2X1  g09970(.A(n11687), .B(n11726), .Y(n11727));
  INVX1   g09971(.A(n11727), .Y(n11728));
  AOI22X1 g09972(.A0(n10656), .A1(n11728), .B0(n10655), .B1(P3_REG1_REG_24__SCAN_IN), .Y(n11729));
  NAND2X1 g09973(.A(n11729), .B(n11725), .Y(n11730));
  INVX1   g09974(.A(n11730), .Y(n11731));
  OAI22X1 g09975(.A0(n11699), .A1(n10646), .B0(n10638), .B1(n11731), .Y(n11732));
  NOR4X1  g09976(.A(n11724), .B(n11723), .C(n11722), .D(n11732), .Y(n11733));
  NAND2X1 g09977(.A(n10697), .B(P3_REG0_REG_23__SCAN_IN), .Y(n11734));
  OAI21X1 g09978(.A0(n11733), .A1(n10697), .B0(n11734), .Y(P3_U3450));
  INVX1   g09979(.A(n11691), .Y(n11736));
  NOR2X1  g09980(.A(n10590), .B(n10311), .Y(n11737));
  XOR2X1  g09981(.A(n11737), .B(n11731), .Y(n11738));
  INVX1   g09982(.A(n11738), .Y(n11739));
  NOR2X1  g09983(.A(n11699), .B(n11736), .Y(n11740));
  NAND2X1 g09984(.A(n11699), .B(n11736), .Y(n11741));
  AOI21X1 g09985(.A0(n11741), .A1(n11714), .B0(n11740), .Y(n11742));
  NOR2X1  g09986(.A(n11739), .B(n11742), .Y(n11745));
  AOI21X1 g09987(.A0(n11742), .A1(n11739), .B0(n11745), .Y(n11746));
  OAI22X1 g09988(.A0(n11736), .A1(n10781), .B0(n10780), .B1(n11746), .Y(n11747));
  NAND2X1 g09989(.A(n11742), .B(n11739), .Y(n11749));
  OAI21X1 g09990(.A0(n11742), .A1(n11739), .B0(n11749), .Y(n11750));
  OAI21X1 g09991(.A0(n10625), .A1(n10617), .B0(n11750), .Y(n11751));
  OAI21X1 g09992(.A0(n11746), .A1(n10744), .B0(n11751), .Y(n11752));
  INVX1   g09993(.A(n11703), .Y(n11753));
  INVX1   g09994(.A(n11648), .Y(n11754));
  INVX1   g09995(.A(n11698), .Y(n11755));
  OAI21X1 g09996(.A0(n11699), .A1(n11691), .B0(n11755), .Y(n11756));
  OAI21X1 g09997(.A0(n11756), .A1(n11754), .B0(n11705), .Y(n11757));
  NAND2X1 g09998(.A(n11757), .B(n11753), .Y(n11758));
  NOR2X1  g09999(.A(n11756), .B(n11649), .Y(n11759));
  INVX1   g10000(.A(n11759), .Y(n11760));
  OAI21X1 g10001(.A0(n11760), .A1(n11628), .B0(n11758), .Y(n11761));
  XOR2X1  g10002(.A(n11761), .B(n11738), .Y(n11762));
  INVX1   g10003(.A(n11762), .Y(n11763));
  OAI21X1 g10004(.A0(n10628), .A1(n10623), .B0(n11762), .Y(n11764));
  OAI21X1 g10005(.A0(n11763), .A1(n10729), .B0(n11764), .Y(n11765));
  NOR4X1  g10006(.A(P3_REG3_REG_22__SCAN_IN), .B(P3_REG3_REG_24__SCAN_IN), .C(P3_REG3_REG_23__SCAN_IN), .D(n11597), .Y(n11766));
  INVX1   g10007(.A(n11766), .Y(n11767));
  INVX1   g10008(.A(n11687), .Y(n11768));
  NOR3X1  g10009(.A(n11768), .B(P3_REG3_REG_24__SCAN_IN), .C(P3_REG3_REG_25__SCAN_IN), .Y(n11769));
  AOI21X1 g10010(.A0(n11767), .A1(P3_REG3_REG_25__SCAN_IN), .B0(n11769), .Y(n11770));
  NOR2X1  g10011(.A(n11770), .B(n10613), .Y(n11771));
  INVX1   g10012(.A(P3_REG1_REG_25__SCAN_IN), .Y(n11772));
  NOR3X1  g10013(.A(n10601), .B(n10605), .C(n11772), .Y(n11773));
  INVX1   g10014(.A(P3_REG2_REG_25__SCAN_IN), .Y(n11774));
  NAND3X1 g10015(.A(n10601), .B(n10599), .C(P3_REG0_REG_25__SCAN_IN), .Y(n11775));
  OAI21X1 g10016(.A0(n10606), .A1(n11774), .B0(n11775), .Y(n11776));
  NOR3X1  g10017(.A(n11776), .B(n11773), .C(n11771), .Y(n11777));
  INVX1   g10018(.A(n11777), .Y(n11778));
  AOI22X1 g10019(.A0(n11737), .A1(n10734), .B0(n10637), .B1(n11778), .Y(n11779));
  OAI21X1 g10020(.A0(n11763), .A1(n10733), .B0(n11779), .Y(n11780));
  NOR4X1  g10021(.A(n11765), .B(n11752), .C(n11747), .D(n11780), .Y(n11781));
  NAND2X1 g10022(.A(n10697), .B(P3_REG0_REG_24__SCAN_IN), .Y(n11782));
  OAI21X1 g10023(.A0(n11781), .A1(n10697), .B0(n11782), .Y(P3_U3451));
  OAI21X1 g10024(.A0(n10590), .A1(n10311), .B0(n11731), .Y(n11784));
  INVX1   g10025(.A(n11784), .Y(n11785));
  NOR3X1  g10026(.A(n11731), .B(n10590), .C(n10311), .Y(n11786));
  INVX1   g10027(.A(n11786), .Y(n11787));
  OAI21X1 g10028(.A0(n11785), .A1(n11742), .B0(n11787), .Y(n11788));
  OAI21X1 g10029(.A0(n10326), .A1(n10319), .B0(n11247), .Y(n11789));
  XOR2X1  g10030(.A(n11789), .B(n11778), .Y(n11790));
  NOR2X1  g10031(.A(n11788), .B(n11790), .Y(n11791));
  AOI21X1 g10032(.A0(n11790), .A1(n11788), .B0(n11791), .Y(n11793));
  OAI22X1 g10033(.A0(n11731), .A1(n10781), .B0(n10780), .B1(n11793), .Y(n11794));
  NAND2X1 g10034(.A(n11788), .B(n11790), .Y(n11796));
  OAI21X1 g10035(.A0(n11788), .A1(n11790), .B0(n11796), .Y(n11797));
  OAI21X1 g10036(.A0(n10625), .A1(n10617), .B0(n11797), .Y(n11798));
  OAI21X1 g10037(.A0(n11793), .A1(n10744), .B0(n11798), .Y(n11799));
  NOR2X1  g10038(.A(n11737), .B(n11731), .Y(n11800));
  NOR3X1  g10039(.A(n11730), .B(n10590), .C(n10311), .Y(n11801));
  INVX1   g10040(.A(n11801), .Y(n11802));
  AOI21X1 g10041(.A0(n11761), .A1(n11802), .B0(n11800), .Y(n11803));
  XOR2X1  g10042(.A(n11803), .B(n11790), .Y(n11804));
  INVX1   g10043(.A(n11804), .Y(n11805));
  OAI21X1 g10044(.A0(n10628), .A1(n10623), .B0(n11805), .Y(n11806));
  OAI21X1 g10045(.A0(n11804), .A1(n10729), .B0(n11806), .Y(n11807));
  NOR2X1  g10046(.A(n10590), .B(n10327), .Y(n11808));
  INVX1   g10047(.A(P3_REG3_REG_26__SCAN_IN), .Y(n11809));
  XOR2X1  g10048(.A(n11769), .B(n11809), .Y(n11810));
  AOI22X1 g10049(.A0(n10652), .A1(P3_REG0_REG_26__SCAN_IN), .B0(P3_REG2_REG_26__SCAN_IN), .B1(n10653), .Y(n11811));
  INVX1   g10050(.A(n11811), .Y(n11812));
  AOI21X1 g10051(.A0(n10655), .A1(P3_REG1_REG_26__SCAN_IN), .B0(n11812), .Y(n11813));
  OAI21X1 g10052(.A0(n11810), .A1(n10613), .B0(n11813), .Y(n11814));
  AOI22X1 g10053(.A0(n11808), .A1(n10734), .B0(n10637), .B1(n11814), .Y(n11815));
  OAI21X1 g10054(.A0(n11804), .A1(n10733), .B0(n11815), .Y(n11816));
  NOR4X1  g10055(.A(n11807), .B(n11799), .C(n11794), .D(n11816), .Y(n11817));
  NAND2X1 g10056(.A(n10697), .B(P3_REG0_REG_25__SCAN_IN), .Y(n11818));
  OAI21X1 g10057(.A0(n11817), .A1(n10697), .B0(n11818), .Y(P3_U3452));
  INVX1   g10058(.A(n11814), .Y(n11820));
  NOR2X1  g10059(.A(n10590), .B(n10339), .Y(n11821));
  XOR2X1  g10060(.A(n11821), .B(n11820), .Y(n11822));
  NOR2X1  g10061(.A(n11789), .B(n11778), .Y(n11824));
  INVX1   g10062(.A(n11824), .Y(n11825));
  XOR2X1  g10063(.A(n13383), .B(n11822), .Y(n11830));
  NOR2X1  g10064(.A(n11830), .B(n10718), .Y(n11831));
  INVX1   g10065(.A(n11831), .Y(n11832));
  NAND2X1 g10066(.A(n11808), .B(n11778), .Y(n11833));
  INVX1   g10067(.A(n11833), .Y(n11834));
  NOR2X1  g10068(.A(n11834), .B(n11788), .Y(n11835));
  INVX1   g10069(.A(n11821), .Y(n11836));
  NAND2X1 g10070(.A(n11789), .B(n11777), .Y(n11837));
  OAI21X1 g10071(.A0(n11821), .A1(n11814), .B0(n11837), .Y(n11838));
  INVX1   g10072(.A(n11838), .Y(n11839));
  OAI21X1 g10073(.A0(n11836), .A1(n11820), .B0(n11839), .Y(n11840));
  NOR2X1  g10074(.A(n11840), .B(n11835), .Y(n11841));
  NAND2X1 g10075(.A(n11822), .B(n11833), .Y(n11842));
  AOI21X1 g10076(.A0(n11837), .A1(n11788), .B0(n11842), .Y(n11843));
  NOR3X1  g10077(.A(n11843), .B(n11841), .C(n10780), .Y(n11844));
  AOI21X1 g10078(.A0(n11778), .A1(n10680), .B0(n11844), .Y(n11845));
  NOR3X1  g10079(.A(n11843), .B(n11841), .C(n10744), .Y(n11846));
  NOR3X1  g10080(.A(n11843), .B(n11841), .C(n10766), .Y(n11850));
  NOR3X1  g10081(.A(n11843), .B(n11841), .C(n10618), .Y(n11851));
  NOR3X1  g10082(.A(n11851), .B(n11850), .C(n11846), .Y(n11852));
  NAND3X1 g10083(.A(n11852), .B(n11845), .C(n11832), .Y(n11853));
  AOI21X1 g10084(.A0(n10729), .A1(n10728), .B0(n11830), .Y(n11854));
  INVX1   g10085(.A(P3_REG3_REG_27__SCAN_IN), .Y(n11855));
  NOR4X1  g10086(.A(P3_REG3_REG_26__SCAN_IN), .B(P3_REG3_REG_24__SCAN_IN), .C(P3_REG3_REG_25__SCAN_IN), .D(n11768), .Y(n11856));
  NAND3X1 g10087(.A(n11769), .B(n11809), .C(n11855), .Y(n11857));
  OAI21X1 g10088(.A0(n11856), .A1(n11855), .B0(n11857), .Y(n11858));
  INVX1   g10089(.A(n11858), .Y(n11859));
  AOI22X1 g10090(.A0(n10652), .A1(P3_REG0_REG_27__SCAN_IN), .B0(P3_REG2_REG_27__SCAN_IN), .B1(n10653), .Y(n11860));
  INVX1   g10091(.A(n11860), .Y(n11861));
  AOI21X1 g10092(.A0(n10655), .A1(P3_REG1_REG_27__SCAN_IN), .B0(n11861), .Y(n11862));
  OAI21X1 g10093(.A0(n11859), .A1(n10613), .B0(n11862), .Y(n11863));
  AOI22X1 g10094(.A0(n11821), .A1(n10734), .B0(n10637), .B1(n11863), .Y(n11864));
  OAI21X1 g10095(.A0(n11830), .A1(n10733), .B0(n11864), .Y(n11865));
  NOR3X1  g10096(.A(n11865), .B(n11854), .C(n11853), .Y(n11866));
  NAND2X1 g10097(.A(n10697), .B(P3_REG0_REG_26__SCAN_IN), .Y(n11867));
  OAI21X1 g10098(.A0(n11866), .A1(n10697), .B0(n11867), .Y(P3_U3453));
  OAI21X1 g10099(.A0(n10355), .A1(n10348), .B0(n11247), .Y(n11869));
  XOR2X1  g10100(.A(n11869), .B(n11863), .Y(n11870));
  INVX1   g10101(.A(n11870), .Y(n11871));
  NOR3X1  g10102(.A(n11820), .B(n10590), .C(n10339), .Y(n11872));
  AOI21X1 g10103(.A0(n11833), .A1(n11787), .B0(n11838), .Y(n11873));
  NOR3X1  g10104(.A(n11838), .B(n11785), .C(n11742), .Y(n11874));
  NOR3X1  g10105(.A(n11874), .B(n11873), .C(n11872), .Y(n11875));
  XOR2X1  g10106(.A(n11875), .B(n11871), .Y(n11876));
  OAI22X1 g10107(.A0(n11820), .A1(n10781), .B0(n10780), .B1(n11876), .Y(n11877));
  XOR2X1  g10108(.A(n11875), .B(n11870), .Y(n11880));
  OAI21X1 g10109(.A0(n10625), .A1(n10617), .B0(n11880), .Y(n11881));
  OAI21X1 g10110(.A0(n11876), .A1(n10744), .B0(n11881), .Y(n11882));
  NOR2X1  g10111(.A(n11882), .B(n11877), .Y(n11883));
  OAI21X1 g10112(.A0(n10590), .A1(n10339), .B0(n11814), .Y(n11884));
  INVX1   g10113(.A(n11884), .Y(n11885));
  OAI21X1 g10114(.A0(n11803), .A1(n11824), .B0(n13309), .Y(n11887));
  NOR3X1  g10115(.A(n11814), .B(n10590), .C(n10339), .Y(n11888));
  NOR2X1  g10116(.A(n11870), .B(n11888), .Y(n11889));
  OAI21X1 g10117(.A0(n11887), .A1(n11885), .B0(n11889), .Y(n11890));
  NOR2X1  g10118(.A(n11871), .B(n11885), .Y(n11891));
  OAI21X1 g10119(.A0(n13383), .A1(n11888), .B0(n11891), .Y(n11892));
  AOI21X1 g10120(.A0(n11892), .A1(n11890), .B0(n10729), .Y(n11893));
  AOI22X1 g10121(.A0(n11890), .A1(n11892), .B0(n10728), .B1(n10718), .Y(n11894));
  NOR2X1  g10122(.A(n11894), .B(n11893), .Y(n11895));
  NAND2X1 g10123(.A(n11895), .B(n11883), .Y(n11896));
  AOI21X1 g10124(.A0(n11892), .A1(n11890), .B0(n10733), .Y(n11897));
  XOR2X1  g10125(.A(n11857), .B(P3_REG3_REG_28__SCAN_IN), .Y(n11898));
  AOI22X1 g10126(.A0(n10652), .A1(P3_REG0_REG_28__SCAN_IN), .B0(P3_REG2_REG_28__SCAN_IN), .B1(n10653), .Y(n11899));
  INVX1   g10127(.A(n11899), .Y(n11900));
  AOI21X1 g10128(.A0(n10655), .A1(P3_REG1_REG_28__SCAN_IN), .B0(n11900), .Y(n11901));
  OAI21X1 g10129(.A0(n11898), .A1(n10613), .B0(n11901), .Y(n11902));
  INVX1   g10130(.A(n11902), .Y(n11903));
  OAI22X1 g10131(.A0(n11869), .A1(n10646), .B0(n10638), .B1(n11903), .Y(n11904));
  NOR3X1  g10132(.A(n11904), .B(n11897), .C(n11896), .Y(n11905));
  NAND2X1 g10133(.A(n10697), .B(P3_REG0_REG_27__SCAN_IN), .Y(n11906));
  OAI21X1 g10134(.A0(n11905), .A1(n10697), .B0(n11906), .Y(P3_U3454));
  OAI21X1 g10135(.A0(n10387), .A1(n10361), .B0(n11247), .Y(n11908));
  XOR2X1  g10136(.A(n11908), .B(n11902), .Y(n11909));
  INVX1   g10137(.A(n11863), .Y(n11910));
  NAND2X1 g10138(.A(n11869), .B(n11910), .Y(n11911));
  NAND2X1 g10139(.A(n11911), .B(n11784), .Y(n11912));
  NOR3X1  g10140(.A(n11912), .B(n11838), .C(n11742), .Y(n11913));
  NAND2X1 g10141(.A(n11911), .B(n11873), .Y(n11914));
  NOR2X1  g10142(.A(n10590), .B(n10356), .Y(n11915));
  NAND2X1 g10143(.A(n11915), .B(n11863), .Y(n11916));
  NAND2X1 g10144(.A(n11911), .B(n11872), .Y(n11917));
  NAND3X1 g10145(.A(n11917), .B(n11916), .C(n11914), .Y(n11918));
  NOR2X1  g10146(.A(n11918), .B(n11913), .Y(n11919));
  XOR2X1  g10147(.A(n11919), .B(n11909), .Y(n11920));
  NAND2X1 g10148(.A(n11920), .B(n10622), .Y(n11921));
  INVX1   g10149(.A(n11909), .Y(n11922));
  NOR2X1  g10150(.A(n11838), .B(n11742), .Y(n11923));
  NAND3X1 g10151(.A(n11923), .B(n11911), .C(n11784), .Y(n11924));
  NAND4X1 g10152(.A(n11917), .B(n11916), .C(n11914), .D(n11924), .Y(n11925));
  OAI21X1 g10153(.A0(n10625), .A1(n10617), .B0(n11920), .Y(n11927));
  NAND2X1 g10154(.A(n11927), .B(n11921), .Y(n11928));
  OAI22X1 g10155(.A0(n11863), .A1(n11869), .B0(n11836), .B1(n11814), .Y(n11929));
  AOI21X1 g10156(.A0(n11910), .A1(n11884), .B0(n11915), .Y(n11930));
  AOI21X1 g10157(.A0(n11863), .A1(n11885), .B0(n11930), .Y(n11931));
  OAI21X1 g10158(.A0(n11929), .A1(n13383), .B0(n11931), .Y(n11932));
  XOR2X1  g10159(.A(n11932), .B(n11922), .Y(n11933));
  AOI22X1 g10160(.A0(n11863), .A1(n10680), .B0(n10626), .B1(n11920), .Y(n11934));
  OAI21X1 g10161(.A0(n11933), .A1(n10718), .B0(n11934), .Y(n11935));
  AOI21X1 g10162(.A0(n10729), .A1(n10728), .B0(n11933), .Y(n11936));
  INVX1   g10163(.A(n10361), .Y(n11937));
  AOI21X1 g10164(.A0(n10385), .A1(n10367), .B0(n10363), .Y(n11938));
  NOR3X1  g10165(.A(n10365), .B(n10364), .C(n10362), .Y(n11939));
  OAI21X1 g10166(.A0(n11939), .A1(n11938), .B0(n1790), .Y(n11940));
  AOI21X1 g10167(.A0(n11940), .A1(n11937), .B0(n10590), .Y(n11941));
  INVX1   g10168(.A(P3_REG3_REG_28__SCAN_IN), .Y(n11942));
  NAND4X1 g10169(.A(n11809), .B(n11942), .C(n11855), .D(n11769), .Y(n11943));
  NOR2X1  g10170(.A(n11943), .B(n10613), .Y(n11944));
  NAND3X1 g10171(.A(n10601), .B(n10599), .C(P3_REG0_REG_29__SCAN_IN), .Y(n11945));
  INVX1   g10172(.A(n11945), .Y(n11946));
  AOI22X1 g10173(.A0(n10653), .A1(P3_REG2_REG_29__SCAN_IN), .B0(P3_REG1_REG_29__SCAN_IN), .B1(n10655), .Y(n11947));
  INVX1   g10174(.A(n11947), .Y(n11948));
  NOR3X1  g10175(.A(n11948), .B(n11946), .C(n11944), .Y(n11949));
  INVX1   g10176(.A(n11949), .Y(n11950));
  AOI22X1 g10177(.A0(n11941), .A1(n10734), .B0(n10637), .B1(n11950), .Y(n11951));
  OAI21X1 g10178(.A0(n11933), .A1(n10733), .B0(n11951), .Y(n11952));
  NOR4X1  g10179(.A(n11936), .B(n11935), .C(n11928), .D(n11952), .Y(n11953));
  NAND2X1 g10180(.A(n10697), .B(P3_REG0_REG_28__SCAN_IN), .Y(n11954));
  OAI21X1 g10181(.A0(n11953), .A1(n10697), .B0(n11954), .Y(P3_U3455));
  NAND2X1 g10182(.A(n11941), .B(n11903), .Y(n11956));
  OAI21X1 g10183(.A0(n10405), .A1(n10396), .B0(n11247), .Y(n11957));
  XOR2X1  g10184(.A(n11957), .B(n11949), .Y(n11958));
  NAND3X1 g10185(.A(n11958), .B(n11932), .C(n11956), .Y(n11959));
  NAND2X1 g10186(.A(n11908), .B(n11902), .Y(n11960));
  INVX1   g10187(.A(n11929), .Y(n11961));
  OAI21X1 g10188(.A0(n11863), .A1(n11885), .B0(n11869), .Y(n11962));
  OAI21X1 g10189(.A0(n11910), .A1(n11884), .B0(n11962), .Y(n11963));
  AOI21X1 g10190(.A0(n11961), .A1(n11887), .B0(n11963), .Y(n11964));
  XOR2X1  g10191(.A(n11957), .B(n11950), .Y(n11965));
  NAND3X1 g10192(.A(n11965), .B(n11964), .C(n11960), .Y(n11966));
  NOR2X1  g10193(.A(n11958), .B(n11956), .Y(n11967));
  NOR2X1  g10194(.A(n11965), .B(n11960), .Y(n11968));
  NOR2X1  g10195(.A(n11968), .B(n11967), .Y(n11969));
  NAND3X1 g10196(.A(n11969), .B(n11966), .C(n11959), .Y(n11970));
  OAI21X1 g10197(.A0(n10629), .A1(n10628), .B0(n11970), .Y(n11971));
  NOR2X1  g10198(.A(n11919), .B(n11908), .Y(n11972));
  AOI21X1 g10199(.A0(n11919), .A1(n11908), .B0(n11903), .Y(n11973));
  NOR3X1  g10200(.A(n11973), .B(n11972), .C(n11965), .Y(n11974));
  OAI21X1 g10201(.A0(n11918), .A1(n11913), .B0(n11941), .Y(n11975));
  OAI21X1 g10202(.A0(n11925), .A1(n11941), .B0(n11902), .Y(n11979));
  AOI21X1 g10203(.A0(n11979), .A1(n11975), .B0(n11958), .Y(n11980));
  OAI22X1 g10204(.A0(n11974), .A1(n11980), .B0(n10626), .B1(n10622), .Y(n11981));
  NAND2X1 g10205(.A(n11981), .B(n11971), .Y(n11982));
  NAND2X1 g10206(.A(n11979), .B(n11975), .Y(n11985));
  XOR2X1  g10207(.A(n11985), .B(n11965), .Y(n11986));
  INVX1   g10208(.A(n11944), .Y(n11987));
  NAND3X1 g10209(.A(n10611), .B(n10599), .C(P3_REG1_REG_30__SCAN_IN), .Y(n11988));
  AOI22X1 g10210(.A0(n10652), .A1(P3_REG0_REG_30__SCAN_IN), .B0(P3_REG2_REG_30__SCAN_IN), .B1(n10653), .Y(n11989));
  NAND3X1 g10211(.A(n11989), .B(n11988), .C(n11987), .Y(n11990));
  NOR2X1  g10212(.A(n10560), .B(n10563), .Y(n11991));
  INVX1   g10213(.A(n10589), .Y(n11992));
  NOR3X1  g10214(.A(n11992), .B(n10678), .C(P3_B_REG_SCAN_IN), .Y(n11993));
  OAI21X1 g10215(.A0(n11993), .A1(n10590), .B0(n11991), .Y(n11994));
  INVX1   g10216(.A(n11994), .Y(n11995));
  AOI22X1 g10217(.A0(n11990), .A1(n11995), .B0(n11902), .B1(n10680), .Y(n11996));
  OAI21X1 g10218(.A0(n11986), .A1(n10618), .B0(n11996), .Y(n11997));
  INVX1   g10219(.A(n11956), .Y(n11998));
  NOR3X1  g10220(.A(n11965), .B(n11964), .C(n11998), .Y(n11999));
  NAND2X1 g10221(.A(n11969), .B(n11966), .Y(n12000));
  NOR2X1  g10222(.A(n12000), .B(n11999), .Y(n12001));
  OAI22X1 g10223(.A0(n12001), .A1(n10718), .B0(n10766), .B1(n11986), .Y(n12002));
  OAI22X1 g10224(.A0(n11957), .A1(n10646), .B0(n10733), .B1(n12001), .Y(n12003));
  NOR4X1  g10225(.A(n12002), .B(n11997), .C(n11982), .D(n12003), .Y(n12004));
  NAND2X1 g10226(.A(n10697), .B(P3_REG0_REG_29__SCAN_IN), .Y(n12005));
  OAI21X1 g10227(.A0(n12004), .A1(n10697), .B0(n12005), .Y(P3_U3456));
  NAND3X1 g10228(.A(n10601), .B(n10599), .C(P3_REG0_REG_31__SCAN_IN), .Y(n12007));
  AOI22X1 g10229(.A0(n10653), .A1(P3_REG2_REG_31__SCAN_IN), .B0(P3_REG1_REG_31__SCAN_IN), .B1(n10655), .Y(n12008));
  NAND3X1 g10230(.A(n12008), .B(n12007), .C(n11987), .Y(n12009));
  INVX1   g10231(.A(n12009), .Y(n12010));
  NOR2X1  g10232(.A(n12010), .B(n11994), .Y(n12011));
  INVX1   g10233(.A(n10411), .Y(n12012));
  AOI21X1 g10234(.A0(n10418), .A1(n10417), .B0(n10413), .Y(n12013));
  NOR3X1  g10235(.A(n10415), .B(n10414), .C(n10412), .Y(n12014));
  OAI21X1 g10236(.A0(n12014), .A1(n12013), .B0(n1790), .Y(n12015));
  AOI21X1 g10237(.A0(n12015), .A1(n12012), .B0(n10590), .Y(n12016));
  AOI21X1 g10238(.A0(n12016), .A1(n10734), .B0(n12011), .Y(n12017));
  NAND2X1 g10239(.A(n10697), .B(P3_REG0_REG_30__SCAN_IN), .Y(n12018));
  OAI21X1 g10240(.A0(n12017), .A1(n10697), .B0(n12018), .Y(P3_U3457));
  INVX1   g10241(.A(n10429), .Y(n12020));
  AOI21X1 g10242(.A0(n10418), .A1(n10417), .B0(n12020), .Y(n12021));
  INVX1   g10243(.A(n10433), .Y(n12022));
  OAI21X1 g10244(.A0(n12022), .A1(n10415), .B0(n10435), .Y(n12023));
  OAI21X1 g10245(.A0(n12023), .A1(n12021), .B0(n1790), .Y(n12024));
  AOI21X1 g10246(.A0(n12024), .A1(n10426), .B0(n10590), .Y(n12025));
  AOI21X1 g10247(.A0(n12025), .A1(n10734), .B0(n12011), .Y(n12026));
  NAND2X1 g10248(.A(n10697), .B(P3_REG0_REG_31__SCAN_IN), .Y(n12027));
  OAI21X1 g10249(.A0(n12026), .A1(n10697), .B0(n12027), .Y(P3_U3458));
  INVX1   g10250(.A(n10567), .Y(n12029));
  AOI21X1 g10251(.A0(n12029), .A1(n10563), .B0(n10578), .Y(n12030));
  OAI21X1 g10252(.A0(n10576), .A1(n12029), .B0(n12030), .Y(n12031));
  NAND4X1 g10253(.A(n10557), .B(n10552), .C(n10549), .D(n12031), .Y(n12032));
  NOR3X1  g10254(.A(n10580), .B(n10575), .C(n10564), .Y(n12033));
  NOR2X1  g10255(.A(n12033), .B(n10581), .Y(n12034));
  NOR4X1  g10256(.A(n10557), .B(n10552), .C(n10550), .D(n12034), .Y(n12035));
  INVX1   g10257(.A(n12035), .Y(n12036));
  AOI21X1 g10258(.A0(n12036), .A1(n12032), .B0(n10529), .Y(n12037));
  NAND2X1 g10259(.A(n12037), .B(n10649), .Y(n12038));
  OAI21X1 g10260(.A0(n12037), .A1(n10609), .B0(n12038), .Y(P3_U3459));
  NAND2X1 g10261(.A(n12037), .B(n10694), .Y(n12040));
  OAI21X1 g10262(.A0(n12037), .A1(n10643), .B0(n12040), .Y(P3_U3460));
  INVX1   g10263(.A(n12037), .Y(n12042));
  NAND2X1 g10264(.A(n12042), .B(P3_REG1_REG_2__SCAN_IN), .Y(n12043));
  OAI21X1 g10265(.A0(n12042), .A1(n10741), .B0(n12043), .Y(P3_U3461));
  NAND2X1 g10266(.A(n12042), .B(P3_REG1_REG_3__SCAN_IN), .Y(n12045));
  OAI21X1 g10267(.A0(n12042), .A1(n10796), .B0(n12045), .Y(P3_U3462));
  NAND2X1 g10268(.A(n12042), .B(P3_REG1_REG_4__SCAN_IN), .Y(n12047));
  OAI21X1 g10269(.A0(n12042), .A1(n10847), .B0(n12047), .Y(P3_U3463));
  NAND2X1 g10270(.A(n12042), .B(P3_REG1_REG_5__SCAN_IN), .Y(n12049));
  OAI21X1 g10271(.A0(n12042), .A1(n10900), .B0(n12049), .Y(P3_U3464));
  NAND2X1 g10272(.A(n12042), .B(P3_REG1_REG_6__SCAN_IN), .Y(n12051));
  OAI21X1 g10273(.A0(n12042), .A1(n10949), .B0(n12051), .Y(P3_U3465));
  NAND2X1 g10274(.A(n12042), .B(P3_REG1_REG_7__SCAN_IN), .Y(n12053));
  OAI21X1 g10275(.A0(n12042), .A1(n10999), .B0(n12053), .Y(P3_U3466));
  NAND2X1 g10276(.A(n12042), .B(P3_REG1_REG_8__SCAN_IN), .Y(n12055));
  OAI21X1 g10277(.A0(n12042), .A1(n11039), .B0(n12055), .Y(P3_U3467));
  NAND2X1 g10278(.A(n12042), .B(P3_REG1_REG_9__SCAN_IN), .Y(n12057));
  OAI21X1 g10279(.A0(n12042), .A1(n11089), .B0(n12057), .Y(P3_U3468));
  NAND2X1 g10280(.A(n12042), .B(P3_REG1_REG_10__SCAN_IN), .Y(n12059));
  OAI21X1 g10281(.A0(n12042), .A1(n11134), .B0(n12059), .Y(P3_U3469));
  NAND2X1 g10282(.A(n12042), .B(P3_REG1_REG_11__SCAN_IN), .Y(n12061));
  OAI21X1 g10283(.A0(n12042), .A1(n11194), .B0(n12061), .Y(P3_U3470));
  NAND2X1 g10284(.A(n12042), .B(P3_REG1_REG_12__SCAN_IN), .Y(n12063));
  OAI21X1 g10285(.A0(n12042), .A1(n11242), .B0(n12063), .Y(P3_U3471));
  NAND2X1 g10286(.A(n12042), .B(P3_REG1_REG_13__SCAN_IN), .Y(n12065));
  OAI21X1 g10287(.A0(n12042), .A1(n11295), .B0(n12065), .Y(P3_U3472));
  NAND2X1 g10288(.A(n12042), .B(P3_REG1_REG_14__SCAN_IN), .Y(n12067));
  OAI21X1 g10289(.A0(n12042), .A1(n11334), .B0(n12067), .Y(P3_U3473));
  NAND2X1 g10290(.A(n12042), .B(P3_REG1_REG_15__SCAN_IN), .Y(n12069));
  OAI21X1 g10291(.A0(n12042), .A1(n11372), .B0(n12069), .Y(P3_U3474));
  NAND2X1 g10292(.A(n12042), .B(P3_REG1_REG_16__SCAN_IN), .Y(n12071));
  OAI21X1 g10293(.A0(n12042), .A1(n11427), .B0(n12071), .Y(P3_U3475));
  NAND2X1 g10294(.A(n12042), .B(P3_REG1_REG_17__SCAN_IN), .Y(n12073));
  OAI21X1 g10295(.A0(n12042), .A1(n11476), .B0(n12073), .Y(P3_U3476));
  NAND2X1 g10296(.A(n12042), .B(P3_REG1_REG_18__SCAN_IN), .Y(n12075));
  OAI21X1 g10297(.A0(n12042), .A1(n11518), .B0(n12075), .Y(P3_U3477));
  NAND2X1 g10298(.A(n12042), .B(P3_REG1_REG_19__SCAN_IN), .Y(n12077));
  OAI21X1 g10299(.A0(n12042), .A1(n11557), .B0(n12077), .Y(P3_U3478));
  NAND2X1 g10300(.A(n12042), .B(P3_REG1_REG_20__SCAN_IN), .Y(n12079));
  OAI21X1 g10301(.A0(n12042), .A1(n11604), .B0(n12079), .Y(P3_U3479));
  NAND2X1 g10302(.A(n12042), .B(P3_REG1_REG_21__SCAN_IN), .Y(n12081));
  OAI21X1 g10303(.A0(n12042), .A1(n11642), .B0(n12081), .Y(P3_U3480));
  NAND2X1 g10304(.A(n12042), .B(P3_REG1_REG_22__SCAN_IN), .Y(n12083));
  OAI21X1 g10305(.A0(n12042), .A1(n11694), .B0(n12083), .Y(P3_U3481));
  NAND2X1 g10306(.A(n12042), .B(P3_REG1_REG_23__SCAN_IN), .Y(n12085));
  OAI21X1 g10307(.A0(n12042), .A1(n11733), .B0(n12085), .Y(P3_U3482));
  NAND2X1 g10308(.A(n12042), .B(P3_REG1_REG_24__SCAN_IN), .Y(n12087));
  OAI21X1 g10309(.A0(n12042), .A1(n11781), .B0(n12087), .Y(P3_U3483));
  NAND2X1 g10310(.A(n12042), .B(P3_REG1_REG_25__SCAN_IN), .Y(n12089));
  OAI21X1 g10311(.A0(n12042), .A1(n11817), .B0(n12089), .Y(P3_U3484));
  NAND2X1 g10312(.A(n12042), .B(P3_REG1_REG_26__SCAN_IN), .Y(n12091));
  OAI21X1 g10313(.A0(n12042), .A1(n11866), .B0(n12091), .Y(P3_U3485));
  NAND2X1 g10314(.A(n12042), .B(P3_REG1_REG_27__SCAN_IN), .Y(n12093));
  OAI21X1 g10315(.A0(n12042), .A1(n11905), .B0(n12093), .Y(P3_U3486));
  NAND2X1 g10316(.A(n12042), .B(P3_REG1_REG_28__SCAN_IN), .Y(n12095));
  OAI21X1 g10317(.A0(n12042), .A1(n11953), .B0(n12095), .Y(P3_U3487));
  NAND2X1 g10318(.A(n12042), .B(P3_REG1_REG_29__SCAN_IN), .Y(n12097));
  OAI21X1 g10319(.A0(n12042), .A1(n12004), .B0(n12097), .Y(P3_U3488));
  NAND2X1 g10320(.A(n12042), .B(P3_REG1_REG_30__SCAN_IN), .Y(n12099));
  OAI21X1 g10321(.A0(n12042), .A1(n12017), .B0(n12099), .Y(P3_U3489));
  NAND2X1 g10322(.A(n12042), .B(P3_REG1_REG_31__SCAN_IN), .Y(n12101));
  OAI21X1 g10323(.A0(n12042), .A1(n12026), .B0(n12101), .Y(P3_U3490));
  NOR4X1  g10324(.A(n10566), .B(n10564), .C(n10562), .D(n10571), .Y(n12103));
  AOI21X1 g10325(.A0(n10453), .A1(n10449), .B0(n10457), .Y(n12104));
  AOI21X1 g10326(.A0(n10457), .A1(P3_D_REG_0__SCAN_IN), .B0(n12104), .Y(n12105));
  AOI21X1 g10327(.A0(n10576), .A1(n10560), .B0(n10563), .Y(n12106));
  NAND2X1 g10328(.A(n12106), .B(n12029), .Y(n12107));
  NAND4X1 g10329(.A(n12105), .B(n10553), .C(n10549), .D(n12107), .Y(n12108));
  INVX1   g10330(.A(n12108), .Y(n12109));
  NOR4X1  g10331(.A(n12105), .B(n10553), .C(n10550), .D(n12034), .Y(n12110));
  NAND3X1 g10332(.A(n12103), .B(n10528), .C(P3_REG3_REG_0__SCAN_IN), .Y(n12111));
  NOR3X1  g10333(.A(n12110), .B(n12109), .C(n12103), .Y(n12112));
  NOR2X1  g10334(.A(n12112), .B(n10529), .Y(n12113));
  NOR2X1  g10335(.A(n12113), .B(n10596), .Y(n12114));
  AOI21X1 g10336(.A0(n12113), .A1(n10631), .B0(n12114), .Y(n12115));
  NOR3X1  g10337(.A(n12112), .B(n10638), .C(n10529), .Y(n12116));
  NAND2X1 g10338(.A(n12116), .B(n10662), .Y(n12117));
  NOR3X1  g10339(.A(n10576), .B(n10564), .C(n10562), .Y(n12118));
  NOR3X1  g10340(.A(n10571), .B(n10564), .C(n10562), .Y(n12119));
  AOI21X1 g10341(.A0(n12119), .A1(n10566), .B0(n12118), .Y(n12120));
  NOR3X1  g10342(.A(n12120), .B(n12112), .C(n10529), .Y(n12121));
  NOR2X1  g10343(.A(n10566), .B(n10560), .Y(n12122));
  INVX1   g10344(.A(n12122), .Y(n12123));
  NOR4X1  g10345(.A(n12112), .B(n10571), .C(n10529), .D(n12123), .Y(n12124));
  AOI22X1 g10346(.A0(n12121), .A1(n10595), .B0(n13412), .B1(n12124), .Y(n12125));
  NAND4X1 g10347(.A(n12117), .B(n12115), .C(n12111), .D(n12125), .Y(P3_U3233));
  NAND3X1 g10348(.A(n12103), .B(n10528), .C(P3_REG3_REG_1__SCAN_IN), .Y(n12127));
  NOR2X1  g10349(.A(n12113), .B(n10640), .Y(n12128));
  AOI21X1 g10350(.A0(n12113), .A1(n10683), .B0(n12128), .Y(n12129));
  INVX1   g10351(.A(n12121), .Y(n12130));
  INVX1   g10352(.A(n12124), .Y(n12131));
  OAI22X1 g10353(.A0(n12130), .A1(n10667), .B0(n10669), .B1(n12131), .Y(n12132));
  AOI21X1 g10354(.A0(n12116), .A1(n10709), .B0(n12132), .Y(n12133));
  NAND3X1 g10355(.A(n12133), .B(n12129), .C(n12127), .Y(P3_U3232));
  NAND3X1 g10356(.A(n12103), .B(n10528), .C(P3_REG3_REG_2__SCAN_IN), .Y(n12135));
  NOR2X1  g10357(.A(n12113), .B(n10685), .Y(n12136));
  AOI21X1 g10358(.A0(n12113), .A1(n10732), .B0(n12136), .Y(n12137));
  OAI22X1 g10359(.A0(n12130), .A1(n10705), .B0(n10725), .B1(n12131), .Y(n12138));
  AOI21X1 g10360(.A0(n12116), .A1(n10738), .B0(n12138), .Y(n12139));
  NAND3X1 g10361(.A(n12139), .B(n12137), .C(n12135), .Y(P3_U3231));
  NAND3X1 g10362(.A(n12103), .B(n10528), .C(n10736), .Y(n12141));
  NOR2X1  g10363(.A(n12113), .B(n10756), .Y(n12142));
  AOI21X1 g10364(.A0(n12113), .A1(n10785), .B0(n12142), .Y(n12143));
  NAND2X1 g10365(.A(n12116), .B(n10793), .Y(n12144));
  AOI22X1 g10366(.A0(n12121), .A1(n10788), .B0(n10779), .B1(n12124), .Y(n12145));
  NAND4X1 g10367(.A(n12144), .B(n12143), .C(n12141), .D(n12145), .Y(P3_U3230));
  INVX1   g10368(.A(n12113), .Y(n12147));
  INVX1   g10369(.A(n12103), .Y(n12148));
  NOR2X1  g10370(.A(n12148), .B(n10529), .Y(n12149));
  AOI22X1 g10371(.A0(n12147), .A1(P3_REG2_REG_4__SCAN_IN), .B0(n10791), .B1(n12149), .Y(n12150));
  AOI22X1 g10372(.A0(n12121), .A1(n10835), .B0(n10829), .B1(n12124), .Y(n12151));
  AOI22X1 g10373(.A0(n12113), .A1(n10833), .B0(n10844), .B1(n12116), .Y(n12152));
  NAND3X1 g10374(.A(n12152), .B(n12151), .C(n12150), .Y(P3_U3229));
  NOR3X1  g10375(.A(n10889), .B(n10876), .C(n10874), .Y(n12154));
  INVX1   g10376(.A(n12149), .Y(n12155));
  OAI22X1 g10377(.A0(n12113), .A1(n10856), .B0(n10841), .B1(n12155), .Y(n12156));
  NOR4X1  g10378(.A(n10914), .B(n10638), .C(n10529), .D(n12112), .Y(n12157));
  OAI22X1 g10379(.A0(n12130), .A1(n10861), .B0(n10886), .B1(n12131), .Y(n12158));
  NOR3X1  g10380(.A(n12158), .B(n12157), .C(n12156), .Y(n12159));
  OAI21X1 g10381(.A0(n12147), .A1(n12154), .B0(n12159), .Y(P3_U3228));
  NOR3X1  g10382(.A(n10940), .B(n10927), .C(n10924), .Y(n12161));
  OAI22X1 g10383(.A0(n12113), .A1(n10909), .B0(n10894), .B1(n12155), .Y(n12162));
  INVX1   g10384(.A(n12116), .Y(n12163));
  AOI22X1 g10385(.A0(n12121), .A1(n10919), .B0(n10937), .B1(n12124), .Y(n12164));
  OAI21X1 g10386(.A0(n12163), .A1(n10957), .B0(n12164), .Y(n12165));
  NOR2X1  g10387(.A(n12165), .B(n12162), .Y(n12166));
  OAI21X1 g10388(.A0(n12147), .A1(n12161), .B0(n12166), .Y(P3_U3227));
  NAND2X1 g10389(.A(n12113), .B(n10990), .Y(n12168));
  AOI22X1 g10390(.A0(n12147), .A1(P3_REG2_REG_7__SCAN_IN), .B0(n10944), .B1(n12149), .Y(n12169));
  OAI22X1 g10391(.A0(n12130), .A1(n10977), .B0(n10970), .B1(n12131), .Y(n12170));
  AOI21X1 g10392(.A0(n12116), .A1(n10996), .B0(n12170), .Y(n12171));
  NAND3X1 g10393(.A(n12171), .B(n12169), .C(n12168), .Y(P3_U3226));
  NAND2X1 g10394(.A(n12113), .B(n11025), .Y(n12173));
  OAI22X1 g10395(.A0(n12113), .A1(n11056), .B0(n10993), .B1(n12155), .Y(n12174));
  NOR4X1  g10396(.A(n11045), .B(n10638), .C(n10529), .D(n12112), .Y(n12175));
  INVX1   g10397(.A(n11006), .Y(n12176));
  OAI22X1 g10398(.A0(n12130), .A1(n12176), .B0(n11012), .B1(n12131), .Y(n12177));
  NOR3X1  g10399(.A(n12177), .B(n12175), .C(n12174), .Y(n12178));
  NAND2X1 g10400(.A(n12178), .B(n12173), .Y(P3_U3225));
  INVX1   g10401(.A(P3_REG2_REG_9__SCAN_IN), .Y(n12180));
  OAI22X1 g10402(.A0(n12113), .A1(n12180), .B0(n11033), .B1(n12155), .Y(n12181));
  NOR4X1  g10403(.A(n11095), .B(n10638), .C(n10529), .D(n12112), .Y(n12182));
  OAI22X1 g10404(.A0(n12130), .A1(n11092), .B0(n11072), .B1(n12131), .Y(n12183));
  NOR3X1  g10405(.A(n12183), .B(n12182), .C(n12181), .Y(n12184));
  OAI21X1 g10406(.A0(n12147), .A1(n11079), .B0(n12184), .Y(P3_U3224));
  NOR3X1  g10407(.A(n11121), .B(n11120), .C(n11119), .Y(n12186));
  INVX1   g10408(.A(P3_REG2_REG_10__SCAN_IN), .Y(n12187));
  OAI22X1 g10409(.A0(n12113), .A1(n12187), .B0(n11100), .B1(n12130), .Y(n12188));
  NOR4X1  g10410(.A(n11140), .B(n10638), .C(n10529), .D(n12112), .Y(n12189));
  OAI22X1 g10411(.A0(n12155), .A1(n11083), .B0(n11115), .B1(n12131), .Y(n12190));
  NOR3X1  g10412(.A(n12190), .B(n12189), .C(n12188), .Y(n12191));
  OAI21X1 g10413(.A0(n12147), .A1(n12186), .B0(n12191), .Y(P3_U3223));
  NOR3X1  g10414(.A(n11184), .B(n11172), .C(n11170), .Y(n12193));
  AOI22X1 g10415(.A0(n12147), .A1(P3_REG2_REG_11__SCAN_IN), .B0(n11191), .B1(n12116), .Y(n12194));
  INVX1   g10416(.A(n11128), .Y(n12195));
  AOI22X1 g10417(.A0(n12149), .A1(n12195), .B0(n11145), .B1(n12121), .Y(n12196));
  NAND2X1 g10418(.A(n12196), .B(n12194), .Y(n12197));
  AOI21X1 g10419(.A0(n12124), .A1(n11155), .B0(n12197), .Y(n12198));
  OAI21X1 g10420(.A0(n12147), .A1(n12193), .B0(n12198), .Y(P3_U3222));
  INVX1   g10421(.A(P3_REG2_REG_12__SCAN_IN), .Y(n12200));
  OAI22X1 g10422(.A0(n12113), .A1(n12200), .B0(n11202), .B1(n12130), .Y(n12201));
  NOR4X1  g10423(.A(n11266), .B(n10638), .C(n10529), .D(n12112), .Y(n12202));
  OAI22X1 g10424(.A0(n12155), .A1(n11188), .B0(n11220), .B1(n12131), .Y(n12203));
  NOR3X1  g10425(.A(n12203), .B(n12202), .C(n12201), .Y(n12204));
  OAI21X1 g10426(.A0(n12147), .A1(n11230), .B0(n12204), .Y(P3_U3221));
  NOR3X1  g10427(.A(n11287), .B(n11282), .C(n11280), .Y(n12206));
  AOI22X1 g10428(.A0(n12147), .A1(P3_REG2_REG_13__SCAN_IN), .B0(n11292), .B1(n12116), .Y(n12207));
  AOI22X1 g10429(.A0(n12149), .A1(n11237), .B0(n11251), .B1(n12121), .Y(n12208));
  NAND2X1 g10430(.A(n12208), .B(n12207), .Y(n12209));
  AOI21X1 g10431(.A0(n12124), .A1(n11277), .B0(n12209), .Y(n12210));
  OAI21X1 g10432(.A0(n12147), .A1(n12206), .B0(n12210), .Y(P3_U3220));
  NOR3X1  g10433(.A(n11322), .B(n11321), .C(n11314), .Y(n12212));
  NOR2X1  g10434(.A(n12131), .B(n11318), .Y(n12213));
  INVX1   g10435(.A(P3_REG2_REG_14__SCAN_IN), .Y(n12214));
  OAI22X1 g10436(.A0(n12113), .A1(n12214), .B0(n11337), .B1(n12163), .Y(n12215));
  OAI22X1 g10437(.A0(n12155), .A1(n11289), .B0(n11302), .B1(n12130), .Y(n12216));
  NOR3X1  g10438(.A(n12216), .B(n12215), .C(n12213), .Y(n12217));
  OAI21X1 g10439(.A0(n12147), .A1(n12212), .B0(n12217), .Y(P3_U3219));
  NOR3X1  g10440(.A(n11363), .B(n11362), .C(n11354), .Y(n12219));
  NOR2X1  g10441(.A(n12131), .B(n11359), .Y(n12220));
  INVX1   g10442(.A(P3_REG2_REG_15__SCAN_IN), .Y(n12221));
  OAI22X1 g10443(.A0(n12113), .A1(n12221), .B0(n11377), .B1(n12163), .Y(n12222));
  INVX1   g10444(.A(n11329), .Y(n12223));
  OAI22X1 g10445(.A0(n12155), .A1(n12223), .B0(n11390), .B1(n12130), .Y(n12224));
  NOR3X1  g10446(.A(n12224), .B(n12222), .C(n12220), .Y(n12225));
  OAI21X1 g10447(.A0(n12147), .A1(n12219), .B0(n12225), .Y(P3_U3218));
  NOR3X1  g10448(.A(n11415), .B(n11410), .C(n11408), .Y(n12227));
  AOI22X1 g10449(.A0(n12147), .A1(P3_REG2_REG_16__SCAN_IN), .B0(n11424), .B1(n12116), .Y(n12228));
  AOI22X1 g10450(.A0(n12149), .A1(n11367), .B0(n11382), .B1(n12121), .Y(n12229));
  NAND2X1 g10451(.A(n12229), .B(n12228), .Y(n12230));
  AOI21X1 g10452(.A0(n12124), .A1(n11396), .B0(n12230), .Y(n12231));
  OAI21X1 g10453(.A0(n12147), .A1(n12227), .B0(n12231), .Y(P3_U3217));
  NOR3X1  g10454(.A(n11467), .B(n11462), .C(n11461), .Y(n12233));
  AOI22X1 g10455(.A0(n12147), .A1(P3_REG2_REG_17__SCAN_IN), .B0(n11473), .B1(n12116), .Y(n12234));
  AOI22X1 g10456(.A0(n12149), .A1(n11422), .B0(n11436), .B1(n12121), .Y(n12235));
  NAND2X1 g10457(.A(n12235), .B(n12234), .Y(n12236));
  AOI21X1 g10458(.A0(n12124), .A1(n11458), .B0(n12236), .Y(n12237));
  OAI21X1 g10459(.A0(n12147), .A1(n12233), .B0(n12237), .Y(P3_U3216));
  NOR3X1  g10460(.A(n11506), .B(n11505), .C(n11493), .Y(n12239));
  AOI22X1 g10461(.A0(n12147), .A1(P3_REG2_REG_18__SCAN_IN), .B0(n11515), .B1(n12116), .Y(n12240));
  AOI22X1 g10462(.A0(n12149), .A1(n11471), .B0(n11508), .B1(n12121), .Y(n12241));
  NAND2X1 g10463(.A(n12241), .B(n12240), .Y(n12242));
  AOI21X1 g10464(.A0(n12124), .A1(n11490), .B0(n12242), .Y(n12243));
  OAI21X1 g10465(.A0(n12147), .A1(n12239), .B0(n12243), .Y(P3_U3215));
  AOI22X1 g10466(.A0(n12147), .A1(P3_REG2_REG_19__SCAN_IN), .B0(n11554), .B1(n12116), .Y(n12245));
  AOI22X1 g10467(.A0(n12149), .A1(n11513), .B0(n11523), .B1(n12121), .Y(n12246));
  NAND2X1 g10468(.A(n12246), .B(n12245), .Y(n12247));
  AOI21X1 g10469(.A0(n12124), .A1(n11530), .B0(n12247), .Y(n12248));
  OAI21X1 g10470(.A0(n12147), .A1(n11548), .B0(n12248), .Y(P3_U3214));
  OAI21X1 g10471(.A0(n11594), .A1(n11582), .B0(n12113), .Y(n12250));
  OAI21X1 g10472(.A0(n12112), .A1(n10529), .B0(P3_REG2_REG_20__SCAN_IN), .Y(n12251));
  OAI21X1 g10473(.A0(n12163), .A1(n11607), .B0(n12251), .Y(n12252));
  AOI21X1 g10474(.A0(n12149), .A1(n11552), .B0(n12252), .Y(n12253));
  OAI21X1 g10475(.A0(n12130), .A1(n11563), .B0(n12253), .Y(n12254));
  AOI21X1 g10476(.A0(n12124), .A1(n11592), .B0(n12254), .Y(n12255));
  NAND2X1 g10477(.A(n12255), .B(n12250), .Y(P3_U3213));
  NAND2X1 g10478(.A(n12113), .B(n11633), .Y(n12257));
  NOR2X1  g10479(.A(n12131), .B(n11629), .Y(n12258));
  NOR3X1  g10480(.A(n12130), .B(n10590), .C(n10271), .Y(n12259));
  INVX1   g10481(.A(n11599), .Y(n12260));
  AOI22X1 g10482(.A0(n12147), .A1(P3_REG2_REG_21__SCAN_IN), .B0(n11639), .B1(n12116), .Y(n12261));
  OAI21X1 g10483(.A0(n12155), .A1(n12260), .B0(n12261), .Y(n12262));
  NOR3X1  g10484(.A(n12262), .B(n12259), .C(n12258), .Y(n12263));
  NAND2X1 g10485(.A(n12263), .B(n12257), .Y(P3_U3212));
  NAND2X1 g10486(.A(n12113), .B(n11684), .Y(n12265));
  NAND2X1 g10487(.A(n12124), .B(n11667), .Y(n12266));
  AOI22X1 g10488(.A0(n12147), .A1(P3_REG2_REG_22__SCAN_IN), .B0(n11691), .B1(n12116), .Y(n12267));
  OAI21X1 g10489(.A0(n12155), .A1(n11636), .B0(n12267), .Y(n12268));
  AOI21X1 g10490(.A0(n12121), .A1(n11646), .B0(n12268), .Y(n12269));
  NAND3X1 g10491(.A(n12269), .B(n12266), .C(n12265), .Y(P3_U3211));
  OAI21X1 g10492(.A0(n11723), .A1(n11722), .B0(n12113), .Y(n12271));
  AOI21X1 g10493(.A0(n11708), .A1(n11702), .B0(n12131), .Y(n12272));
  NOR2X1  g10494(.A(n12130), .B(n11699), .Y(n12273));
  NOR2X1  g10495(.A(n11689), .B(n11687), .Y(n12274));
  AOI22X1 g10496(.A0(n12147), .A1(P3_REG2_REG_23__SCAN_IN), .B0(n11730), .B1(n12116), .Y(n12275));
  OAI21X1 g10497(.A0(n12155), .A1(n12274), .B0(n12275), .Y(n12276));
  NOR3X1  g10498(.A(n12276), .B(n12273), .C(n12272), .Y(n12277));
  NAND2X1 g10499(.A(n12277), .B(n12271), .Y(P3_U3210));
  NOR3X1  g10500(.A(n11765), .B(n11752), .C(n11747), .Y(n12279));
  INVX1   g10501(.A(n11737), .Y(n12280));
  OAI21X1 g10502(.A0(n12112), .A1(n10529), .B0(P3_REG2_REG_24__SCAN_IN), .Y(n12281));
  OAI21X1 g10503(.A0(n12163), .A1(n11777), .B0(n12281), .Y(n12282));
  AOI21X1 g10504(.A0(n12149), .A1(n11728), .B0(n12282), .Y(n12283));
  OAI21X1 g10505(.A0(n12130), .A1(n12280), .B0(n12283), .Y(n12284));
  AOI21X1 g10506(.A0(n12124), .A1(n11762), .B0(n12284), .Y(n12285));
  OAI21X1 g10507(.A0(n12147), .A1(n12279), .B0(n12285), .Y(P3_U3209));
  NOR3X1  g10508(.A(n11807), .B(n11799), .C(n11794), .Y(n12287));
  INVX1   g10509(.A(n11770), .Y(n12288));
  OAI22X1 g10510(.A0(n12113), .A1(n11774), .B0(n11820), .B1(n12163), .Y(n12289));
  AOI21X1 g10511(.A0(n12149), .A1(n12288), .B0(n12289), .Y(n12290));
  OAI21X1 g10512(.A0(n12130), .A1(n11789), .B0(n12290), .Y(n12291));
  AOI21X1 g10513(.A0(n12124), .A1(n11805), .B0(n12291), .Y(n12292));
  OAI21X1 g10514(.A0(n12147), .A1(n12287), .B0(n12292), .Y(P3_U3208));
  OAI21X1 g10515(.A0(n11854), .A1(n11853), .B0(n12113), .Y(n12294));
  NOR2X1  g10516(.A(n12131), .B(n11830), .Y(n12295));
  NOR3X1  g10517(.A(n12130), .B(n10590), .C(n10339), .Y(n12296));
  AOI22X1 g10518(.A0(n12147), .A1(P3_REG2_REG_26__SCAN_IN), .B0(n11863), .B1(n12116), .Y(n12297));
  OAI21X1 g10519(.A0(n12155), .A1(n11810), .B0(n12297), .Y(n12298));
  NOR3X1  g10520(.A(n12298), .B(n12296), .C(n12295), .Y(n12299));
  NAND2X1 g10521(.A(n12299), .B(n12294), .Y(P3_U3207));
  NOR4X1  g10522(.A(n11893), .B(n11882), .C(n11877), .D(n11894), .Y(n12301));
  AOI21X1 g10523(.A0(n11892), .A1(n11890), .B0(n12131), .Y(n12302));
  NOR2X1  g10524(.A(n12130), .B(n11869), .Y(n12303));
  AOI22X1 g10525(.A0(n12147), .A1(P3_REG2_REG_27__SCAN_IN), .B0(n11902), .B1(n12116), .Y(n12304));
  OAI21X1 g10526(.A0(n12155), .A1(n11859), .B0(n12304), .Y(n12305));
  NOR3X1  g10527(.A(n12305), .B(n12303), .C(n12302), .Y(n12306));
  OAI21X1 g10528(.A0(n12147), .A1(n12301), .B0(n12306), .Y(P3_U3206));
  NOR3X1  g10529(.A(n11936), .B(n11935), .C(n11928), .Y(n12308));
  NOR2X1  g10530(.A(n12131), .B(n11933), .Y(n12309));
  NOR2X1  g10531(.A(n12130), .B(n11908), .Y(n12310));
  AOI22X1 g10532(.A0(n12147), .A1(P3_REG2_REG_28__SCAN_IN), .B0(n11950), .B1(n12116), .Y(n12311));
  OAI21X1 g10533(.A0(n12155), .A1(n11898), .B0(n12311), .Y(n12312));
  NOR3X1  g10534(.A(n12312), .B(n12310), .C(n12309), .Y(n12313));
  OAI21X1 g10535(.A0(n12147), .A1(n12308), .B0(n12313), .Y(P3_U3205));
  NOR3X1  g10536(.A(n12002), .B(n11997), .C(n11982), .Y(n12315));
  NOR2X1  g10537(.A(n12155), .B(n11943), .Y(n12316));
  AOI21X1 g10538(.A0(n12147), .A1(P3_REG2_REG_29__SCAN_IN), .B0(n12316), .Y(n12317));
  OAI21X1 g10539(.A0(n12130), .A1(n11957), .B0(n12317), .Y(n12318));
  AOI21X1 g10540(.A0(n12124), .A1(n11970), .B0(n12318), .Y(n12319));
  OAI21X1 g10541(.A0(n12147), .A1(n12315), .B0(n12319), .Y(P3_U3204));
  OAI21X1 g10542(.A0(n10420), .A1(n10411), .B0(n11247), .Y(n12321));
  NAND3X1 g10543(.A(n12113), .B(n12009), .C(n11995), .Y(n12322));
  OAI21X1 g10544(.A0(n12155), .A1(n11943), .B0(n12322), .Y(n12323));
  AOI21X1 g10545(.A0(n12147), .A1(P3_REG2_REG_30__SCAN_IN), .B0(n12323), .Y(n12324));
  OAI21X1 g10546(.A0(n12130), .A1(n12321), .B0(n12324), .Y(P3_U3203));
  OAI21X1 g10547(.A0(n10438), .A1(n10427), .B0(n11247), .Y(n12326));
  AOI21X1 g10548(.A0(n12147), .A1(P3_REG2_REG_31__SCAN_IN), .B0(n12323), .Y(n12327));
  OAI21X1 g10549(.A0(n12130), .A1(n12326), .B0(n12327), .Y(P3_U3202));
  AOI21X1 g10550(.A0(n10454), .A1(n10445), .B0(P3_U3151), .Y(n12329));
  OAI21X1 g10551(.A0(n10589), .A1(n10587), .B0(n10446), .Y(n12330));
  OAI22X1 g10552(.A0(n10587), .A1(n10589), .B0(n10560), .B1(n10563), .Y(n12331));
  NAND3X1 g10553(.A(n12331), .B(n12330), .C(n12329), .Y(n12332));
  INVX1   g10554(.A(n12332), .Y(n12333));
  NOR2X1  g10555(.A(n12333), .B(n10529), .Y(n12334));
  INVX1   g10556(.A(P3_REG2_REG_17__SCAN_IN), .Y(n12335));
  NOR2X1  g10557(.A(n11379), .B(P3_REG2_REG_16__SCAN_IN), .Y(n12336));
  NAND2X1 g10558(.A(n11300), .B(n12214), .Y(n12337));
  NOR2X1  g10559(.A(n11300), .B(n12214), .Y(n12338));
  NOR2X1  g10560(.A(n11249), .B(P3_REG2_REG_13__SCAN_IN), .Y(n12339));
  NAND2X1 g10561(.A(n11249), .B(P3_REG2_REG_13__SCAN_IN), .Y(n12340));
  NAND2X1 g10562(.A(n11200), .B(n12200), .Y(n12341));
  NOR2X1  g10563(.A(n11200), .B(n12200), .Y(n12342));
  NOR2X1  g10564(.A(n11142), .B(P3_REG2_REG_11__SCAN_IN), .Y(n12343));
  NAND2X1 g10565(.A(n11142), .B(P3_REG2_REG_11__SCAN_IN), .Y(n12344));
  NAND2X1 g10566(.A(n11098), .B(n12187), .Y(n12345));
  NOR2X1  g10567(.A(n11098), .B(n12187), .Y(n12346));
  NOR2X1  g10568(.A(n11047), .B(P3_REG2_REG_9__SCAN_IN), .Y(n12347));
  NAND2X1 g10569(.A(n11047), .B(P3_REG2_REG_9__SCAN_IN), .Y(n12348));
  NAND2X1 g10570(.A(n11004), .B(n11056), .Y(n12349));
  NOR2X1  g10571(.A(n11004), .B(n11056), .Y(n12350));
  NOR2X1  g10572(.A(n10959), .B(P3_REG2_REG_7__SCAN_IN), .Y(n12351));
  NAND2X1 g10573(.A(n10959), .B(P3_REG2_REG_7__SCAN_IN), .Y(n12352));
  NAND2X1 g10574(.A(n10917), .B(n10909), .Y(n12353));
  NOR2X1  g10575(.A(n10917), .B(n10909), .Y(n12354));
  NOR2X1  g10576(.A(n10852), .B(P3_REG2_REG_5__SCAN_IN), .Y(n12355));
  NAND2X1 g10577(.A(n10852), .B(P3_REG2_REG_5__SCAN_IN), .Y(n12356));
  NAND2X1 g10578(.A(n10801), .B(n10811), .Y(n12357));
  NOR2X1  g10579(.A(n10801), .B(n10811), .Y(n12358));
  NOR2X1  g10580(.A(n10702), .B(P3_REG2_REG_2__SCAN_IN), .Y(n12359));
  INVX1   g10581(.A(n12359), .Y(n12360));
  NOR2X1  g10582(.A(n10593), .B(n10596), .Y(n12361));
  NOR2X1  g10583(.A(n12361), .B(P3_REG2_REG_1__SCAN_IN), .Y(n12362));
  AOI21X1 g10584(.A0(n12361), .A1(P3_REG2_REG_1__SCAN_IN), .B0(n10664), .Y(n12363));
  OAI22X1 g10585(.A0(n12362), .A1(n12363), .B0(n10703), .B1(n10685), .Y(n12364));
  AOI22X1 g10586(.A0(n12360), .A1(n12364), .B0(n10750), .B1(P3_REG2_REG_3__SCAN_IN), .Y(n12365));
  AOI21X1 g10587(.A0(n10751), .A1(n10756), .B0(n12365), .Y(n12366));
  OAI21X1 g10588(.A0(n12366), .A1(n12358), .B0(n12357), .Y(n12367));
  AOI21X1 g10589(.A0(n12367), .A1(n12356), .B0(n12355), .Y(n12368));
  OAI21X1 g10590(.A0(n12368), .A1(n12354), .B0(n12353), .Y(n12369));
  AOI21X1 g10591(.A0(n12369), .A1(n12352), .B0(n12351), .Y(n12370));
  OAI21X1 g10592(.A0(n12370), .A1(n12350), .B0(n12349), .Y(n12371));
  AOI21X1 g10593(.A0(n12371), .A1(n12348), .B0(n12347), .Y(n12372));
  OAI21X1 g10594(.A0(n12372), .A1(n12346), .B0(n12345), .Y(n12373));
  AOI21X1 g10595(.A0(n12373), .A1(n12344), .B0(n12343), .Y(n12374));
  OAI21X1 g10596(.A0(n12374), .A1(n12342), .B0(n12341), .Y(n12375));
  AOI21X1 g10597(.A0(n12375), .A1(n12340), .B0(n12339), .Y(n12376));
  OAI21X1 g10598(.A0(n12376), .A1(n12338), .B0(n12337), .Y(n12377));
  NAND2X1 g10599(.A(n12377), .B(n12221), .Y(n12378));
  OAI21X1 g10600(.A0(n12377), .A1(n12221), .B0(n11340), .Y(n12379));
  AOI22X1 g10601(.A0(n12378), .A1(n12379), .B0(n11379), .B1(P3_REG2_REG_16__SCAN_IN), .Y(n12380));
  OAI22X1 g10602(.A0(n12336), .A1(n12380), .B0(n11433), .B1(n12335), .Y(n12381));
  OAI21X1 g10603(.A0(n11432), .A1(P3_REG2_REG_17__SCAN_IN), .B0(n12381), .Y(n12382));
  NOR2X1  g10604(.A(n11480), .B(P3_REG2_REG_18__SCAN_IN), .Y(n12383));
  XOR2X1  g10605(.A(n10571), .B(P3_REG2_REG_19__SCAN_IN), .Y(n12384));
  AOI21X1 g10606(.A0(n11480), .A1(P3_REG2_REG_18__SCAN_IN), .B0(n12384), .Y(n12385));
  OAI21X1 g10607(.A0(n12383), .A1(n12382), .B0(n12385), .Y(n12386));
  INVX1   g10608(.A(n12383), .Y(n12387));
  INVX1   g10609(.A(P3_REG2_REG_18__SCAN_IN), .Y(n12388));
  OAI21X1 g10610(.A0(n11481), .A1(n12388), .B0(n12382), .Y(n12389));
  NAND3X1 g10611(.A(n12389), .B(n12384), .C(n12387), .Y(n12390));
  NOR2X1  g10612(.A(n11992), .B(n10678), .Y(n12391));
  INVX1   g10613(.A(n12391), .Y(n12392));
  INVX1   g10614(.A(n12120), .Y(n12393));
  AOI21X1 g10615(.A0(n12390), .A1(n12386), .B0(n12392), .Y(n12400));
  NOR2X1  g10616(.A(n11432), .B(P3_REG1_REG_17__SCAN_IN), .Y(n12401));
  INVX1   g10617(.A(P3_REG1_REG_17__SCAN_IN), .Y(n12402));
  NOR2X1  g10618(.A(n11433), .B(n12402), .Y(n12403));
  INVX1   g10619(.A(n12403), .Y(n12404));
  INVX1   g10620(.A(P3_REG1_REG_16__SCAN_IN), .Y(n12405));
  INVX1   g10621(.A(P3_REG1_REG_14__SCAN_IN), .Y(n12406));
  NOR2X1  g10622(.A(n11300), .B(n12406), .Y(n12407));
  NOR2X1  g10623(.A(n11249), .B(P3_REG1_REG_13__SCAN_IN), .Y(n12408));
  NAND2X1 g10624(.A(n11249), .B(P3_REG1_REG_13__SCAN_IN), .Y(n12409));
  INVX1   g10625(.A(P3_REG1_REG_12__SCAN_IN), .Y(n12410));
  NAND2X1 g10626(.A(n11200), .B(n12410), .Y(n12411));
  NOR2X1  g10627(.A(n11200), .B(n12410), .Y(n12412));
  NOR2X1  g10628(.A(n11142), .B(P3_REG1_REG_11__SCAN_IN), .Y(n12413));
  NAND2X1 g10629(.A(n11142), .B(P3_REG1_REG_11__SCAN_IN), .Y(n12414));
  INVX1   g10630(.A(P3_REG1_REG_10__SCAN_IN), .Y(n12415));
  NAND2X1 g10631(.A(n11098), .B(n12415), .Y(n12416));
  NOR2X1  g10632(.A(n11098), .B(n12415), .Y(n12417));
  NOR2X1  g10633(.A(n11047), .B(P3_REG1_REG_9__SCAN_IN), .Y(n12418));
  NAND2X1 g10634(.A(n11047), .B(P3_REG1_REG_9__SCAN_IN), .Y(n12419));
  NAND2X1 g10635(.A(n11004), .B(n11059), .Y(n12420));
  NOR2X1  g10636(.A(n11004), .B(n11059), .Y(n12421));
  NOR2X1  g10637(.A(n10959), .B(P3_REG1_REG_7__SCAN_IN), .Y(n12422));
  NAND2X1 g10638(.A(n10959), .B(P3_REG1_REG_7__SCAN_IN), .Y(n12423));
  NAND2X1 g10639(.A(n10917), .B(n10912), .Y(n12424));
  NOR2X1  g10640(.A(n10917), .B(n10912), .Y(n12425));
  NOR2X1  g10641(.A(n10852), .B(P3_REG1_REG_5__SCAN_IN), .Y(n12426));
  NAND2X1 g10642(.A(n10852), .B(P3_REG1_REG_5__SCAN_IN), .Y(n12427));
  NAND2X1 g10643(.A(n10801), .B(n10814), .Y(n12428));
  NOR2X1  g10644(.A(n10801), .B(n10814), .Y(n12429));
  NOR2X1  g10645(.A(n10702), .B(P3_REG1_REG_2__SCAN_IN), .Y(n12430));
  INVX1   g10646(.A(n12430), .Y(n12431));
  NOR2X1  g10647(.A(n10593), .B(n10609), .Y(n12432));
  NOR2X1  g10648(.A(n12432), .B(P3_REG1_REG_1__SCAN_IN), .Y(n12433));
  AOI21X1 g10649(.A0(n12432), .A1(P3_REG1_REG_1__SCAN_IN), .B0(n10664), .Y(n12434));
  OAI22X1 g10650(.A0(n12433), .A1(n12434), .B0(n10703), .B1(n10689), .Y(n12435));
  AOI22X1 g10651(.A0(n12431), .A1(n12435), .B0(n10750), .B1(P3_REG1_REG_3__SCAN_IN), .Y(n12436));
  AOI21X1 g10652(.A0(n10751), .A1(n10759), .B0(n12436), .Y(n12437));
  OAI21X1 g10653(.A0(n12437), .A1(n12429), .B0(n12428), .Y(n12438));
  AOI21X1 g10654(.A0(n12438), .A1(n12427), .B0(n12426), .Y(n12439));
  OAI21X1 g10655(.A0(n12439), .A1(n12425), .B0(n12424), .Y(n12440));
  AOI21X1 g10656(.A0(n12440), .A1(n12423), .B0(n12422), .Y(n12441));
  OAI21X1 g10657(.A0(n12441), .A1(n12421), .B0(n12420), .Y(n12442));
  AOI21X1 g10658(.A0(n12442), .A1(n12419), .B0(n12418), .Y(n12443));
  OAI21X1 g10659(.A0(n12443), .A1(n12417), .B0(n12416), .Y(n12444));
  AOI21X1 g10660(.A0(n12444), .A1(n12414), .B0(n12413), .Y(n12445));
  OAI21X1 g10661(.A0(n12445), .A1(n12412), .B0(n12411), .Y(n12446));
  AOI21X1 g10662(.A0(n12446), .A1(n12409), .B0(n12408), .Y(n12447));
  NOR2X1  g10663(.A(n12447), .B(n12407), .Y(n12448));
  AOI21X1 g10664(.A0(n11300), .A1(n12406), .B0(n12448), .Y(n12449));
  NOR2X1  g10665(.A(n12449), .B(P3_REG1_REG_15__SCAN_IN), .Y(n12450));
  AOI21X1 g10666(.A0(n12449), .A1(P3_REG1_REG_15__SCAN_IN), .B0(n11339), .Y(n12451));
  OAI22X1 g10667(.A0(n12450), .A1(n12451), .B0(n11380), .B1(n12405), .Y(n12452));
  OAI21X1 g10668(.A0(n11379), .A1(P3_REG1_REG_16__SCAN_IN), .B0(n12452), .Y(n12453));
  AOI21X1 g10669(.A0(n12453), .A1(n12404), .B0(n12401), .Y(n12454));
  OAI21X1 g10670(.A0(n11480), .A1(P3_REG1_REG_18__SCAN_IN), .B0(n12454), .Y(n12455));
  XOR2X1  g10671(.A(n10571), .B(P3_REG1_REG_19__SCAN_IN), .Y(n12456));
  AOI21X1 g10672(.A0(n11480), .A1(P3_REG1_REG_18__SCAN_IN), .B0(n12456), .Y(n12457));
  AOI21X1 g10673(.A0(n11480), .A1(P3_REG1_REG_18__SCAN_IN), .B0(n12454), .Y(n12458));
  OAI21X1 g10674(.A0(n11480), .A1(P3_REG1_REG_18__SCAN_IN), .B0(n12456), .Y(n12459));
  NOR2X1  g10675(.A(n12459), .B(n12458), .Y(n12460));
  AOI21X1 g10676(.A0(n12457), .A1(n12455), .B0(n12460), .Y(n12461));
  OAI22X1 g10677(.A0(n10587), .A1(n12461), .B0(n10571), .B1(n10589), .Y(n12466));
  OAI21X1 g10678(.A0(n12466), .A1(n12400), .B0(n12334), .Y(n12467));
  NOR4X1  g10679(.A(n10587), .B(n10445), .C(P3_U3151), .D(n12333), .Y(n12468));
  INVX1   g10680(.A(n12468), .Y(n12469));
  NOR2X1  g10681(.A(n12469), .B(n12461), .Y(n12470));
  NOR4X1  g10682(.A(n12392), .B(n10445), .C(P3_U3151), .D(n12333), .Y(n12471));
  INVX1   g10683(.A(n12471), .Y(n12472));
  AOI21X1 g10684(.A0(n12390), .A1(n12386), .B0(n12472), .Y(n12473));
  INVX1   g10685(.A(P3_REG1_REG_19__SCAN_IN), .Y(n12474));
  NOR2X1  g10686(.A(n10587), .B(n12474), .Y(n12475));
  AOI21X1 g10687(.A0(n10587), .A1(P3_REG2_REG_19__SCAN_IN), .B0(n12475), .Y(n12476));
  XOR2X1  g10688(.A(n12476), .B(n10571), .Y(n12477));
  NAND2X1 g10689(.A(n10678), .B(P3_REG1_REG_18__SCAN_IN), .Y(n12478));
  OAI21X1 g10690(.A0(n10678), .A1(n12388), .B0(n12478), .Y(n12479));
  NOR2X1  g10691(.A(n10678), .B(n12335), .Y(n12480));
  AOI21X1 g10692(.A0(n10678), .A1(P3_REG1_REG_17__SCAN_IN), .B0(n12480), .Y(n12481));
  INVX1   g10693(.A(n12481), .Y(n12482));
  NAND2X1 g10694(.A(n12482), .B(n11432), .Y(n12483));
  NOR2X1  g10695(.A(n12482), .B(n11432), .Y(n12484));
  NOR2X1  g10696(.A(n10587), .B(n12405), .Y(n12485));
  AOI21X1 g10697(.A0(n10587), .A1(P3_REG2_REG_16__SCAN_IN), .B0(n12485), .Y(n12486));
  INVX1   g10698(.A(n12486), .Y(n12487));
  NOR2X1  g10699(.A(n12487), .B(n11379), .Y(n12488));
  INVX1   g10700(.A(n12488), .Y(n12489));
  NOR2X1  g10701(.A(n10678), .B(n12221), .Y(n12490));
  AOI21X1 g10702(.A0(n10678), .A1(P3_REG1_REG_15__SCAN_IN), .B0(n12490), .Y(n12491));
  NOR2X1  g10703(.A(n12491), .B(n11340), .Y(n12492));
  AOI21X1 g10704(.A0(n12487), .A1(n11379), .B0(n12492), .Y(n12493));
  NOR2X1  g10705(.A(n10678), .B(n12214), .Y(n12494));
  AOI21X1 g10706(.A0(n10678), .A1(P3_REG1_REG_14__SCAN_IN), .B0(n12494), .Y(n12495));
  NOR2X1  g10707(.A(n12495), .B(n11300), .Y(n12496));
  INVX1   g10708(.A(n12496), .Y(n12497));
  INVX1   g10709(.A(n12491), .Y(n12498));
  OAI22X1 g10710(.A0(n12487), .A1(n11379), .B0(n11339), .B1(n12498), .Y(n12499));
  OAI21X1 g10711(.A0(n12499), .A1(n12497), .B0(n12493), .Y(n12500));
  INVX1   g10712(.A(n11249), .Y(n12501));
  INVX1   g10713(.A(P3_REG1_REG_13__SCAN_IN), .Y(n12502));
  NOR2X1  g10714(.A(n10587), .B(n12502), .Y(n12503));
  AOI21X1 g10715(.A0(n10587), .A1(P3_REG2_REG_13__SCAN_IN), .B0(n12503), .Y(n12504));
  NAND2X1 g10716(.A(n12504), .B(n12501), .Y(n12505));
  NOR2X1  g10717(.A(n10678), .B(n12200), .Y(n12506));
  AOI21X1 g10718(.A0(n10678), .A1(P3_REG1_REG_12__SCAN_IN), .B0(n12506), .Y(n12507));
  NOR2X1  g10719(.A(n12507), .B(n11200), .Y(n12508));
  INVX1   g10720(.A(P3_REG2_REG_11__SCAN_IN), .Y(n12509));
  NOR2X1  g10721(.A(n10678), .B(n12509), .Y(n12510));
  AOI21X1 g10722(.A0(n10678), .A1(P3_REG1_REG_11__SCAN_IN), .B0(n12510), .Y(n12511));
  INVX1   g10723(.A(n12511), .Y(n12512));
  NOR2X1  g10724(.A(n12512), .B(n11142), .Y(n12513));
  NOR2X1  g10725(.A(n10678), .B(n12187), .Y(n12514));
  AOI21X1 g10726(.A0(n10678), .A1(P3_REG1_REG_10__SCAN_IN), .B0(n12514), .Y(n12515));
  INVX1   g10727(.A(n12515), .Y(n12516));
  AOI22X1 g10728(.A0(n12512), .A1(n11142), .B0(n11097), .B1(n12516), .Y(n12517));
  NOR2X1  g10729(.A(n10587), .B(n11027), .Y(n12518));
  AOI21X1 g10730(.A0(n10587), .A1(P3_REG2_REG_9__SCAN_IN), .B0(n12518), .Y(n12519));
  NOR2X1  g10731(.A(n12519), .B(n11048), .Y(n12520));
  AOI22X1 g10732(.A0(n12511), .A1(n11143), .B0(n11098), .B1(n12515), .Y(n12521));
  NAND2X1 g10733(.A(n12521), .B(n12520), .Y(n12522));
  AOI21X1 g10734(.A0(n12522), .A1(n12517), .B0(n12513), .Y(n12523));
  NOR2X1  g10735(.A(n10678), .B(n10909), .Y(n12524));
  AOI21X1 g10736(.A0(n10678), .A1(P3_REG1_REG_6__SCAN_IN), .B0(n12524), .Y(n12525));
  INVX1   g10737(.A(n12525), .Y(n12526));
  NOR2X1  g10738(.A(n12526), .B(n10916), .Y(n12527));
  INVX1   g10739(.A(n12527), .Y(n12528));
  NOR2X1  g10740(.A(n10678), .B(n10856), .Y(n12529));
  AOI21X1 g10741(.A0(n10678), .A1(P3_REG1_REG_5__SCAN_IN), .B0(n12529), .Y(n12530));
  NOR2X1  g10742(.A(n12530), .B(n10853), .Y(n12531));
  AOI21X1 g10743(.A0(n12526), .A1(n10916), .B0(n12531), .Y(n12532));
  INVX1   g10744(.A(n12532), .Y(n12533));
  NOR2X1  g10745(.A(n10587), .B(n10814), .Y(n12534));
  AOI21X1 g10746(.A0(n10587), .A1(P3_REG2_REG_4__SCAN_IN), .B0(n12534), .Y(n12535));
  NAND2X1 g10747(.A(n12530), .B(n10853), .Y(n12536));
  INVX1   g10748(.A(n12536), .Y(n12537));
  NOR4X1  g10749(.A(n12535), .B(n12527), .C(n10801), .D(n12537), .Y(n12538));
  OAI21X1 g10750(.A0(n12538), .A1(n12533), .B0(n12528), .Y(n12539));
  NOR2X1  g10751(.A(n10587), .B(n10643), .Y(n12540));
  AOI21X1 g10752(.A0(n10587), .A1(P3_REG2_REG_1__SCAN_IN), .B0(n12540), .Y(n12541));
  NOR2X1  g10753(.A(n10587), .B(n10609), .Y(n12542));
  AOI21X1 g10754(.A0(n10587), .A1(P3_REG2_REG_0__SCAN_IN), .B0(n12542), .Y(n12543));
  AOI21X1 g10755(.A0(n12543), .A1(n10593), .B0(n12541), .Y(n12544));
  NAND2X1 g10756(.A(n12543), .B(n10593), .Y(n12545));
  INVX1   g10757(.A(n12545), .Y(n12546));
  AOI21X1 g10758(.A0(n12546), .A1(n12541), .B0(n10665), .Y(n12547));
  NOR2X1  g10759(.A(n12547), .B(n12544), .Y(n12548));
  NOR2X1  g10760(.A(n10678), .B(n10756), .Y(n12549));
  AOI21X1 g10761(.A0(n10678), .A1(P3_REG1_REG_3__SCAN_IN), .B0(n12549), .Y(n12550));
  INVX1   g10762(.A(n12550), .Y(n12551));
  NOR2X1  g10763(.A(n10678), .B(n10685), .Y(n12552));
  AOI21X1 g10764(.A0(n10678), .A1(P3_REG1_REG_2__SCAN_IN), .B0(n12552), .Y(n12553));
  INVX1   g10765(.A(n12553), .Y(n12554));
  OAI22X1 g10766(.A0(n12551), .A1(n10750), .B0(n10702), .B1(n12554), .Y(n12555));
  OAI21X1 g10767(.A0(n12553), .A1(n10703), .B0(n12550), .Y(n12556));
  NOR3X1  g10768(.A(n12553), .B(n12550), .C(n10703), .Y(n12557));
  AOI21X1 g10769(.A0(n12556), .A1(n10750), .B0(n12557), .Y(n12558));
  OAI21X1 g10770(.A0(n12555), .A1(n12548), .B0(n12558), .Y(n12559));
  INVX1   g10771(.A(n12559), .Y(n12560));
  NAND2X1 g10772(.A(n12535), .B(n10801), .Y(n12561));
  NAND3X1 g10773(.A(n12561), .B(n12536), .C(n12528), .Y(n12562));
  OAI21X1 g10774(.A0(n12562), .A1(n12560), .B0(n12539), .Y(n12563));
  INVX1   g10775(.A(n12563), .Y(n12564));
  NOR2X1  g10776(.A(n10678), .B(n11056), .Y(n12565));
  AOI21X1 g10777(.A0(n10678), .A1(P3_REG1_REG_8__SCAN_IN), .B0(n12565), .Y(n12566));
  INVX1   g10778(.A(n12566), .Y(n12567));
  NOR2X1  g10779(.A(n10678), .B(n10952), .Y(n12568));
  AOI21X1 g10780(.A0(n10678), .A1(P3_REG1_REG_7__SCAN_IN), .B0(n12568), .Y(n12569));
  INVX1   g10781(.A(n12569), .Y(n12570));
  OAI22X1 g10782(.A0(n12567), .A1(n11003), .B0(n10959), .B1(n12570), .Y(n12571));
  OAI21X1 g10783(.A0(n12569), .A1(n10960), .B0(n12566), .Y(n12572));
  NOR3X1  g10784(.A(n12569), .B(n12566), .C(n10960), .Y(n12573));
  AOI21X1 g10785(.A0(n12572), .A1(n11003), .B0(n12573), .Y(n12574));
  OAI21X1 g10786(.A0(n12571), .A1(n12564), .B0(n12574), .Y(n12575));
  NOR2X1  g10787(.A(n12516), .B(n11097), .Y(n12576));
  NAND2X1 g10788(.A(n12519), .B(n11048), .Y(n12577));
  INVX1   g10789(.A(n12577), .Y(n12578));
  NOR3X1  g10790(.A(n12578), .B(n12576), .C(n12513), .Y(n12579));
  AOI21X1 g10791(.A0(n12579), .A1(n12575), .B0(n12523), .Y(n12580));
  AOI21X1 g10792(.A0(n12507), .A1(n11200), .B0(n12580), .Y(n12581));
  OAI21X1 g10793(.A0(n12581), .A1(n12508), .B0(n12505), .Y(n12582));
  OAI21X1 g10794(.A0(n12504), .A1(n12501), .B0(n12582), .Y(n12583));
  NOR2X1  g10795(.A(n10587), .B(n12406), .Y(n12584));
  NOR3X1  g10796(.A(n12584), .B(n12494), .C(n11299), .Y(n12585));
  NOR2X1  g10797(.A(n12585), .B(n12499), .Y(n12586));
  AOI22X1 g10798(.A0(n12583), .A1(n12586), .B0(n12500), .B1(n12489), .Y(n12587));
  OAI21X1 g10799(.A0(n12587), .A1(n12484), .B0(n12483), .Y(n12588));
  NAND2X1 g10800(.A(n12588), .B(n12479), .Y(n12589));
  OAI21X1 g10801(.A0(n12588), .A1(n12479), .B0(n11480), .Y(n12590));
  NAND2X1 g10802(.A(n12590), .B(n12589), .Y(n12591));
  XOR2X1  g10803(.A(n12591), .B(n12477), .Y(n12592));
  NOR2X1  g10804(.A(n10589), .B(n10678), .Y(n12593));
  NAND3X1 g10805(.A(n10454), .B(n10445), .C(P3_STATE_REG_SCAN_IN), .Y(n12594));
  INVX1   g10806(.A(n12594), .Y(P3_U3897));
  OAI21X1 g10807(.A0(n12593), .A1(n10590), .B0(P3_U3897), .Y(n12596));
  NOR4X1  g10808(.A(n10589), .B(n10445), .C(P3_U3151), .D(n12333), .Y(n12597));
  AOI21X1 g10809(.A0(P3_U3897), .A1(n10589), .B0(n12597), .Y(n12598));
  INVX1   g10810(.A(n12598), .Y(n12599));
  OAI22X1 g10811(.A0(n1788), .A1(n12332), .B0(n11510), .B1(P3_STATE_REG_SCAN_IN), .Y(n12600));
  AOI21X1 g10812(.A0(n12599), .A1(n10576), .B0(n12600), .Y(n12601));
  OAI21X1 g10813(.A0(n12596), .A1(n12592), .B0(n12601), .Y(n12602));
  NOR3X1  g10814(.A(n12602), .B(n12473), .C(n12470), .Y(n12603));
  NAND2X1 g10815(.A(n12603), .B(n12467), .Y(P3_U3201));
  INVX1   g10816(.A(n12334), .Y(n12605));
  XOR2X1  g10817(.A(n11480), .B(P3_REG2_REG_18__SCAN_IN), .Y(n12606));
  XOR2X1  g10818(.A(n12606), .B(n12382), .Y(n12607));
  XOR2X1  g10819(.A(n11480), .B(P3_REG1_REG_18__SCAN_IN), .Y(n12608));
  XOR2X1  g10820(.A(n12608), .B(n12454), .Y(n12609));
  OAI22X1 g10821(.A0(n10589), .A1(n11480), .B0(n10587), .B1(n12609), .Y(n12610));
  AOI21X1 g10822(.A0(n12607), .A1(n12391), .B0(n12610), .Y(n12611));
  NOR2X1  g10823(.A(n12609), .B(n12469), .Y(n12612));
  INVX1   g10824(.A(n12607), .Y(n12613));
  NOR2X1  g10825(.A(n12613), .B(n12472), .Y(n12614));
  XOR2X1  g10826(.A(n12479), .B(n11481), .Y(n12615));
  XOR2X1  g10827(.A(n12615), .B(n12588), .Y(n12616));
  NOR2X1  g10828(.A(n12616), .B(n12596), .Y(n12617));
  AOI22X1 g10829(.A0(P3_ADDR_REG_18__SCAN_IN), .A1(n12333), .B0(P3_REG3_REG_18__SCAN_IN), .B1(P3_U3151), .Y(n12618));
  OAI21X1 g10830(.A0(n12598), .A1(n11480), .B0(n12618), .Y(n12619));
  NOR4X1  g10831(.A(n12617), .B(n12614), .C(n12612), .D(n12619), .Y(n12620));
  OAI21X1 g10832(.A0(n12611), .A1(n12605), .B0(n12620), .Y(P3_U3200));
  INVX1   g10833(.A(P3_REG2_REG_16__SCAN_IN), .Y(n12622));
  AOI21X1 g10834(.A0(n11380), .A1(n12622), .B0(n12380), .Y(n12623));
  XOR2X1  g10835(.A(n11432), .B(P3_REG2_REG_17__SCAN_IN), .Y(n12624));
  XOR2X1  g10836(.A(n12624), .B(n12623), .Y(n12625));
  XOR2X1  g10837(.A(n11432), .B(P3_REG1_REG_17__SCAN_IN), .Y(n12626));
  XOR2X1  g10838(.A(n12626), .B(n12453), .Y(n12627));
  AOI22X1 g10839(.A0(n11992), .A1(n11433), .B0(n10678), .B1(n12627), .Y(n12628));
  OAI21X1 g10840(.A0(n12625), .A1(n12392), .B0(n12628), .Y(n12629));
  NAND2X1 g10841(.A(n12629), .B(n12334), .Y(n12630));
  NAND2X1 g10842(.A(n12627), .B(n12468), .Y(n12631));
  NOR2X1  g10843(.A(n12625), .B(n12472), .Y(n12632));
  XOR2X1  g10844(.A(n12481), .B(n11433), .Y(n12633));
  XOR2X1  g10845(.A(n12633), .B(n12587), .Y(n12634));
  OAI22X1 g10846(.A0(n1710), .A1(n12332), .B0(n11418), .B1(P3_STATE_REG_SCAN_IN), .Y(n12635));
  AOI21X1 g10847(.A0(n12599), .A1(n11433), .B0(n12635), .Y(n12636));
  OAI21X1 g10848(.A0(n12634), .A1(n12596), .B0(n12636), .Y(n12637));
  NOR2X1  g10849(.A(n12637), .B(n12632), .Y(n12638));
  NAND3X1 g10850(.A(n12638), .B(n12631), .C(n12630), .Y(P3_U3199));
  NAND2X1 g10851(.A(n12379), .B(n12378), .Y(n12640));
  XOR2X1  g10852(.A(n11379), .B(P3_REG2_REG_16__SCAN_IN), .Y(n12641));
  XOR2X1  g10853(.A(n12641), .B(n12640), .Y(n12642));
  INVX1   g10854(.A(P3_REG1_REG_15__SCAN_IN), .Y(n12643));
  INVX1   g10855(.A(n12449), .Y(n12644));
  AOI21X1 g10856(.A0(n12644), .A1(n12643), .B0(n12451), .Y(n12645));
  XOR2X1  g10857(.A(n11379), .B(P3_REG1_REG_16__SCAN_IN), .Y(n12646));
  XOR2X1  g10858(.A(n12646), .B(n12645), .Y(n12647));
  OAI22X1 g10859(.A0(n10589), .A1(n11379), .B0(n10587), .B1(n12647), .Y(n12648));
  AOI21X1 g10860(.A0(n12642), .A1(n12391), .B0(n12648), .Y(n12649));
  NOR2X1  g10861(.A(n12647), .B(n12469), .Y(n12650));
  INVX1   g10862(.A(n12642), .Y(n12651));
  NOR2X1  g10863(.A(n12651), .B(n12472), .Y(n12652));
  INVX1   g10864(.A(n12583), .Y(n12653));
  OAI21X1 g10865(.A0(n12585), .A1(n12653), .B0(n12497), .Y(n12654));
  XOR2X1  g10866(.A(n12487), .B(n11379), .Y(n12655));
  AOI21X1 g10867(.A0(n12491), .A1(n11340), .B0(n12655), .Y(n12656));
  OAI21X1 g10868(.A0(n12654), .A1(n12492), .B0(n12656), .Y(n12657));
  OAI21X1 g10869(.A0(n12498), .A1(n11339), .B0(n12654), .Y(n12658));
  NAND3X1 g10870(.A(n12658), .B(n12493), .C(n12489), .Y(n12659));
  AOI21X1 g10871(.A0(n12659), .A1(n12657), .B0(n12596), .Y(n12660));
  AOI22X1 g10872(.A0(P3_ADDR_REG_16__SCAN_IN), .A1(n12333), .B0(P3_REG3_REG_16__SCAN_IN), .B1(P3_U3151), .Y(n12661));
  OAI21X1 g10873(.A0(n12598), .A1(n11379), .B0(n12661), .Y(n12662));
  NOR4X1  g10874(.A(n12660), .B(n12652), .C(n12650), .D(n12662), .Y(n12663));
  OAI21X1 g10875(.A0(n12649), .A1(n12605), .B0(n12663), .Y(P3_U3198));
  XOR2X1  g10876(.A(n11339), .B(P3_REG2_REG_15__SCAN_IN), .Y(n12665));
  XOR2X1  g10877(.A(n12665), .B(n12377), .Y(n12666));
  XOR2X1  g10878(.A(n11339), .B(P3_REG1_REG_15__SCAN_IN), .Y(n12667));
  XOR2X1  g10879(.A(n12667), .B(n12449), .Y(n12668));
  OAI22X1 g10880(.A0(n10589), .A1(n11339), .B0(n10587), .B1(n12668), .Y(n12669));
  AOI21X1 g10881(.A0(n12666), .A1(n12391), .B0(n12669), .Y(n12670));
  NOR2X1  g10882(.A(n12668), .B(n12469), .Y(n12671));
  INVX1   g10883(.A(n12666), .Y(n12672));
  NOR2X1  g10884(.A(n12672), .B(n12472), .Y(n12673));
  XOR2X1  g10885(.A(n12491), .B(n11339), .Y(n12674));
  XOR2X1  g10886(.A(n12674), .B(n12654), .Y(n12675));
  OAI22X1 g10887(.A0(n1530), .A1(n12332), .B0(n11325), .B1(P3_STATE_REG_SCAN_IN), .Y(n12676));
  AOI21X1 g10888(.A0(n12599), .A1(n11340), .B0(n12676), .Y(n12677));
  OAI21X1 g10889(.A0(n12675), .A1(n12596), .B0(n12677), .Y(n12678));
  NOR3X1  g10890(.A(n12678), .B(n12673), .C(n12671), .Y(n12679));
  OAI21X1 g10891(.A0(n12670), .A1(n12605), .B0(n12679), .Y(P3_U3197));
  XOR2X1  g10892(.A(n11299), .B(P3_REG2_REG_14__SCAN_IN), .Y(n12681));
  XOR2X1  g10893(.A(n12681), .B(n12376), .Y(n12682));
  NOR2X1  g10894(.A(n12682), .B(n12392), .Y(n12683));
  XOR2X1  g10895(.A(n11299), .B(P3_REG1_REG_14__SCAN_IN), .Y(n12684));
  XOR2X1  g10896(.A(n12684), .B(n12447), .Y(n12685));
  OAI22X1 g10897(.A0(n10589), .A1(n11299), .B0(n10587), .B1(n12685), .Y(n12686));
  OAI21X1 g10898(.A0(n12686), .A1(n12683), .B0(n12334), .Y(n12687));
  NOR2X1  g10899(.A(n12685), .B(n12469), .Y(n12688));
  NOR2X1  g10900(.A(n12682), .B(n12472), .Y(n12689));
  XOR2X1  g10901(.A(n12495), .B(n11299), .Y(n12690));
  XOR2X1  g10902(.A(n12690), .B(n12583), .Y(n12691));
  NOR2X1  g10903(.A(n12691), .B(n12596), .Y(n12692));
  AOI22X1 g10904(.A0(P3_ADDR_REG_14__SCAN_IN), .A1(n12333), .B0(P3_REG3_REG_14__SCAN_IN), .B1(P3_U3151), .Y(n12693));
  OAI21X1 g10905(.A0(n12598), .A1(n11299), .B0(n12693), .Y(n12694));
  NOR4X1  g10906(.A(n12692), .B(n12689), .C(n12688), .D(n12694), .Y(n12695));
  NAND2X1 g10907(.A(n12695), .B(n12687), .Y(P3_U3196));
  XOR2X1  g10908(.A(n11249), .B(P3_REG2_REG_13__SCAN_IN), .Y(n12697));
  XOR2X1  g10909(.A(n12697), .B(n12375), .Y(n12698));
  XOR2X1  g10910(.A(n11249), .B(n12502), .Y(n12699));
  XOR2X1  g10911(.A(n12699), .B(n12446), .Y(n12700));
  OAI22X1 g10912(.A0(n10589), .A1(n11249), .B0(n10587), .B1(n12700), .Y(n12701));
  AOI21X1 g10913(.A0(n12698), .A1(n12391), .B0(n12701), .Y(n12702));
  NOR2X1  g10914(.A(n12700), .B(n12469), .Y(n12703));
  INVX1   g10915(.A(n12698), .Y(n12704));
  NOR2X1  g10916(.A(n12704), .B(n12472), .Y(n12705));
  NOR2X1  g10917(.A(n12581), .B(n12508), .Y(n12706));
  XOR2X1  g10918(.A(n12504), .B(n12501), .Y(n12707));
  XOR2X1  g10919(.A(n12707), .B(n12706), .Y(n12708));
  OAI22X1 g10920(.A0(n1540), .A1(n12332), .B0(n11234), .B1(P3_STATE_REG_SCAN_IN), .Y(n12709));
  AOI21X1 g10921(.A0(n12599), .A1(n12501), .B0(n12709), .Y(n12710));
  OAI21X1 g10922(.A0(n12708), .A1(n12596), .B0(n12710), .Y(n12711));
  NOR3X1  g10923(.A(n12711), .B(n12705), .C(n12703), .Y(n12712));
  OAI21X1 g10924(.A0(n12702), .A1(n12605), .B0(n12712), .Y(P3_U3195));
  XOR2X1  g10925(.A(n11199), .B(P3_REG2_REG_12__SCAN_IN), .Y(n12714));
  XOR2X1  g10926(.A(n12714), .B(n12374), .Y(n12715));
  NOR2X1  g10927(.A(n12715), .B(n12392), .Y(n12716));
  XOR2X1  g10928(.A(n11199), .B(P3_REG1_REG_12__SCAN_IN), .Y(n12717));
  XOR2X1  g10929(.A(n12717), .B(n12445), .Y(n12718));
  OAI22X1 g10930(.A0(n10589), .A1(n11199), .B0(n10587), .B1(n12718), .Y(n12719));
  OAI21X1 g10931(.A0(n12719), .A1(n12716), .B0(n12334), .Y(n12720));
  NOR2X1  g10932(.A(n12718), .B(n12469), .Y(n12721));
  NOR2X1  g10933(.A(n12715), .B(n12472), .Y(n12722));
  XOR2X1  g10934(.A(n12507), .B(n11200), .Y(n12723));
  XOR2X1  g10935(.A(n12723), .B(n12580), .Y(n12724));
  OAI22X1 g10936(.A0(n1544), .A1(n12332), .B0(n11187), .B1(P3_STATE_REG_SCAN_IN), .Y(n12725));
  AOI21X1 g10937(.A0(n12599), .A1(n11200), .B0(n12725), .Y(n12726));
  OAI21X1 g10938(.A0(n12724), .A1(n12596), .B0(n12726), .Y(n12727));
  NOR3X1  g10939(.A(n12727), .B(n12722), .C(n12721), .Y(n12728));
  NAND2X1 g10940(.A(n12728), .B(n12720), .Y(P3_U3194));
  XOR2X1  g10941(.A(n11142), .B(P3_REG2_REG_11__SCAN_IN), .Y(n12730));
  XOR2X1  g10942(.A(n12730), .B(n12373), .Y(n12731));
  XOR2X1  g10943(.A(n11142), .B(n11123), .Y(n12732));
  XOR2X1  g10944(.A(n12732), .B(n12444), .Y(n12733));
  OAI22X1 g10945(.A0(n10589), .A1(n11142), .B0(n10587), .B1(n12733), .Y(n12734));
  AOI21X1 g10946(.A0(n12731), .A1(n12391), .B0(n12734), .Y(n12735));
  AOI21X1 g10947(.A0(n12577), .A1(n12575), .B0(n12520), .Y(n12736));
  OAI21X1 g10948(.A0(n12515), .A1(n11098), .B0(n12736), .Y(n12737));
  XOR2X1  g10949(.A(n12511), .B(n11143), .Y(n12738));
  AOI21X1 g10950(.A0(n12515), .A1(n11098), .B0(n12738), .Y(n12739));
  NAND2X1 g10951(.A(n12739), .B(n12737), .Y(n12740));
  INVX1   g10952(.A(n12517), .Y(n12741));
  NOR2X1  g10953(.A(n12741), .B(n12513), .Y(n12742));
  OAI21X1 g10954(.A0(n12736), .A1(n12576), .B0(n12742), .Y(n12743));
  AOI21X1 g10955(.A0(n12743), .A1(n12740), .B0(n12596), .Y(n12744));
  AOI22X1 g10956(.A0(P3_ADDR_REG_11__SCAN_IN), .A1(n12333), .B0(P3_REG3_REG_11__SCAN_IN), .B1(P3_U3151), .Y(n12745));
  OAI21X1 g10957(.A0(n12598), .A1(n11142), .B0(n12745), .Y(n12746));
  AOI21X1 g10958(.A0(n12731), .A1(n12471), .B0(n12746), .Y(n12747));
  OAI21X1 g10959(.A0(n12733), .A1(n12469), .B0(n12747), .Y(n12748));
  NOR2X1  g10960(.A(n12748), .B(n12744), .Y(n12749));
  OAI21X1 g10961(.A0(n12735), .A1(n12605), .B0(n12749), .Y(P3_U3193));
  XOR2X1  g10962(.A(n12515), .B(n11098), .Y(n12751));
  XOR2X1  g10963(.A(n12751), .B(n12736), .Y(n12752));
  XOR2X1  g10964(.A(n11097), .B(P3_REG2_REG_10__SCAN_IN), .Y(n12753));
  XOR2X1  g10965(.A(n12753), .B(n12372), .Y(n12754));
  NOR2X1  g10966(.A(n12754), .B(n12392), .Y(n12755));
  XOR2X1  g10967(.A(n11097), .B(P3_REG1_REG_10__SCAN_IN), .Y(n12756));
  XOR2X1  g10968(.A(n12756), .B(n12443), .Y(n12757));
  OAI22X1 g10969(.A0(n10589), .A1(n11097), .B0(n10587), .B1(n12757), .Y(n12758));
  NOR2X1  g10970(.A(n12758), .B(n12755), .Y(n12759));
  NOR2X1  g10971(.A(n12759), .B(n12605), .Y(n12760));
  NOR2X1  g10972(.A(n12757), .B(n12469), .Y(n12761));
  NOR2X1  g10973(.A(n12754), .B(n12472), .Y(n12762));
  AOI22X1 g10974(.A0(P3_ADDR_REG_10__SCAN_IN), .A1(n12333), .B0(P3_REG3_REG_10__SCAN_IN), .B1(P3_U3151), .Y(n12763));
  OAI21X1 g10975(.A0(n12598), .A1(n11097), .B0(n12763), .Y(n12764));
  NOR4X1  g10976(.A(n12762), .B(n12761), .C(n12760), .D(n12764), .Y(n12765));
  OAI21X1 g10977(.A0(n12752), .A1(n12596), .B0(n12765), .Y(P3_U3192));
  XOR2X1  g10978(.A(n12519), .B(n11047), .Y(n12767));
  XOR2X1  g10979(.A(n12767), .B(n12575), .Y(n12768));
  XOR2X1  g10980(.A(n11047), .B(P3_REG2_REG_9__SCAN_IN), .Y(n12769));
  XOR2X1  g10981(.A(n12769), .B(n12371), .Y(n12770));
  NAND2X1 g10982(.A(n12770), .B(n12391), .Y(n12771));
  XOR2X1  g10983(.A(n11047), .B(P3_REG1_REG_9__SCAN_IN), .Y(n12772));
  XOR2X1  g10984(.A(n12772), .B(n12442), .Y(n12773));
  AOI22X1 g10985(.A0(n11992), .A1(n11048), .B0(n10678), .B1(n12773), .Y(n12774));
  AOI21X1 g10986(.A0(n12774), .A1(n12771), .B0(n12605), .Y(n12775));
  NAND2X1 g10987(.A(n12773), .B(n12468), .Y(n12776));
  AOI22X1 g10988(.A0(P3_ADDR_REG_9__SCAN_IN), .A1(n12333), .B0(P3_REG3_REG_9__SCAN_IN), .B1(P3_U3151), .Y(n12777));
  OAI21X1 g10989(.A0(n12598), .A1(n11047), .B0(n12777), .Y(n12778));
  AOI21X1 g10990(.A0(n12770), .A1(n12471), .B0(n12778), .Y(n12779));
  NAND2X1 g10991(.A(n12779), .B(n12776), .Y(n12780));
  NOR2X1  g10992(.A(n12780), .B(n12775), .Y(n12781));
  OAI21X1 g10993(.A0(n12768), .A1(n12596), .B0(n12781), .Y(P3_U3191));
  INVX1   g10994(.A(n12596), .Y(n12783));
  NOR2X1  g10995(.A(n12570), .B(n10959), .Y(n12784));
  AOI21X1 g10996(.A0(n12570), .A1(n10959), .B0(n12563), .Y(n12785));
  XOR2X1  g10997(.A(n12566), .B(n11004), .Y(n12786));
  NOR3X1  g10998(.A(n12786), .B(n12785), .C(n12784), .Y(n12787));
  INVX1   g10999(.A(n12784), .Y(n12788));
  OAI21X1 g11000(.A0(n12569), .A1(n10960), .B0(n12786), .Y(n12789));
  AOI21X1 g11001(.A0(n12788), .A1(n12563), .B0(n12789), .Y(n12790));
  OAI21X1 g11002(.A0(n12790), .A1(n12787), .B0(n12783), .Y(n12791));
  XOR2X1  g11003(.A(n11003), .B(P3_REG2_REG_8__SCAN_IN), .Y(n12792));
  XOR2X1  g11004(.A(n12792), .B(n12370), .Y(n12793));
  NOR2X1  g11005(.A(n12793), .B(n12392), .Y(n12794));
  XOR2X1  g11006(.A(n11003), .B(P3_REG1_REG_8__SCAN_IN), .Y(n12795));
  XOR2X1  g11007(.A(n12795), .B(n12441), .Y(n12796));
  OAI22X1 g11008(.A0(n10589), .A1(n11003), .B0(n10587), .B1(n12796), .Y(n12797));
  OAI21X1 g11009(.A0(n12797), .A1(n12794), .B0(n12334), .Y(n12798));
  NOR2X1  g11010(.A(n12796), .B(n12469), .Y(n12799));
  NOR2X1  g11011(.A(n12793), .B(n12472), .Y(n12800));
  AOI22X1 g11012(.A0(P3_ADDR_REG_8__SCAN_IN), .A1(n12333), .B0(P3_REG3_REG_8__SCAN_IN), .B1(P3_U3151), .Y(n12801));
  OAI21X1 g11013(.A0(n12598), .A1(n11003), .B0(n12801), .Y(n12802));
  NOR3X1  g11014(.A(n12802), .B(n12800), .C(n12799), .Y(n12803));
  NAND3X1 g11015(.A(n12803), .B(n12798), .C(n12791), .Y(P3_U3190));
  XOR2X1  g11016(.A(n12569), .B(n10960), .Y(n12805));
  XOR2X1  g11017(.A(n12805), .B(n12563), .Y(n12806));
  NAND2X1 g11018(.A(n12806), .B(n12783), .Y(n12807));
  NOR3X1  g11019(.A(n4574), .B(n10959), .C(n10589), .Y(n12808));
  XOR2X1  g11020(.A(n10959), .B(n10955), .Y(n12809));
  XOR2X1  g11021(.A(n12809), .B(n12440), .Y(n12810));
  XOR2X1  g11022(.A(n10959), .B(n10952), .Y(n12811));
  XOR2X1  g11023(.A(n12811), .B(n12369), .Y(n12812));
  OAI22X1 g11024(.A0(n12810), .A1(n10587), .B0(n12392), .B1(n12812), .Y(n12813));
  OAI21X1 g11025(.A0(n12813), .A1(n12808), .B0(n12334), .Y(n12814));
  NOR2X1  g11026(.A(n12598), .B(n10959), .Y(n12815));
  NOR2X1  g11027(.A(n12810), .B(n12469), .Y(n12816));
  AOI22X1 g11028(.A0(P3_ADDR_REG_7__SCAN_IN), .A1(n12333), .B0(P3_REG3_REG_7__SCAN_IN), .B1(P3_U3151), .Y(n12817));
  OAI21X1 g11029(.A0(n12812), .A1(n12472), .B0(n12817), .Y(n12818));
  NOR3X1  g11030(.A(n12818), .B(n12816), .C(n12815), .Y(n12819));
  NAND3X1 g11031(.A(n12819), .B(n12814), .C(n12807), .Y(P3_U3189));
  NOR2X1  g11032(.A(n12535), .B(n10801), .Y(n12821));
  AOI21X1 g11033(.A0(n12561), .A1(n12559), .B0(n12821), .Y(n12822));
  OAI21X1 g11034(.A0(n12530), .A1(n10853), .B0(n12822), .Y(n12823));
  XOR2X1  g11035(.A(n12525), .B(n10917), .Y(n12824));
  AOI21X1 g11036(.A0(n12530), .A1(n10853), .B0(n12824), .Y(n12825));
  NOR2X1  g11037(.A(n12822), .B(n12537), .Y(n12826));
  NOR3X1  g11038(.A(n12826), .B(n12533), .C(n12527), .Y(n12827));
  AOI21X1 g11039(.A0(n12825), .A1(n12823), .B0(n12827), .Y(n12828));
  XOR2X1  g11040(.A(n10916), .B(n10912), .Y(n12829));
  XOR2X1  g11041(.A(n12829), .B(n12439), .Y(n12830));
  XOR2X1  g11042(.A(n10916), .B(n10909), .Y(n12831));
  XOR2X1  g11043(.A(n12831), .B(n12368), .Y(n12832));
  AOI22X1 g11044(.A0(n12830), .A1(n10678), .B0(n12391), .B1(n12832), .Y(n12833));
  OAI21X1 g11045(.A0(n10589), .A1(n10916), .B0(n12833), .Y(n12834));
  NAND2X1 g11046(.A(n12599), .B(n10917), .Y(n12835));
  NAND2X1 g11047(.A(n12830), .B(n12468), .Y(n12836));
  OAI22X1 g11048(.A0(n1559), .A1(n12332), .B0(n10892), .B1(P3_STATE_REG_SCAN_IN), .Y(n12837));
  AOI21X1 g11049(.A0(n12832), .A1(n12471), .B0(n12837), .Y(n12838));
  NAND3X1 g11050(.A(n12838), .B(n12836), .C(n12835), .Y(n12839));
  AOI21X1 g11051(.A0(n12834), .A1(n12334), .B0(n12839), .Y(n12840));
  OAI21X1 g11052(.A0(n12828), .A1(n12596), .B0(n12840), .Y(P3_U3188));
  XOR2X1  g11053(.A(n12530), .B(n10853), .Y(n12842));
  XOR2X1  g11054(.A(n12842), .B(n12822), .Y(n12843));
  NAND2X1 g11055(.A(n11992), .B(n10853), .Y(n12844));
  XOR2X1  g11056(.A(n10852), .B(P3_REG1_REG_5__SCAN_IN), .Y(n12845));
  XOR2X1  g11057(.A(n12845), .B(n12438), .Y(n12846));
  XOR2X1  g11058(.A(n10852), .B(P3_REG2_REG_5__SCAN_IN), .Y(n12847));
  XOR2X1  g11059(.A(n12847), .B(n12367), .Y(n12848));
  AOI22X1 g11060(.A0(n12846), .A1(n10678), .B0(n12391), .B1(n12848), .Y(n12849));
  AOI21X1 g11061(.A0(n12849), .A1(n12844), .B0(n12605), .Y(n12850));
  NOR2X1  g11062(.A(n12598), .B(n10852), .Y(n12851));
  NAND2X1 g11063(.A(n12846), .B(n12468), .Y(n12852));
  OAI22X1 g11064(.A0(n1561), .A1(n12332), .B0(n10839), .B1(P3_STATE_REG_SCAN_IN), .Y(n12853));
  AOI21X1 g11065(.A0(n12848), .A1(n12471), .B0(n12853), .Y(n12854));
  NAND2X1 g11066(.A(n12854), .B(n12852), .Y(n12855));
  NOR3X1  g11067(.A(n12855), .B(n12851), .C(n12850), .Y(n12856));
  OAI21X1 g11068(.A0(n12843), .A1(n12596), .B0(n12856), .Y(P3_U3187));
  INVX1   g11069(.A(n10801), .Y(n12858));
  NOR3X1  g11070(.A(n4574), .B(n12858), .C(n10589), .Y(n12859));
  XOR2X1  g11071(.A(n10801), .B(n10814), .Y(n12860));
  XOR2X1  g11072(.A(n12860), .B(n12437), .Y(n12861));
  XOR2X1  g11073(.A(n10801), .B(n10811), .Y(n12862));
  XOR2X1  g11074(.A(n12862), .B(n12366), .Y(n12863));
  OAI22X1 g11075(.A0(n12861), .A1(n10587), .B0(n12392), .B1(n12863), .Y(n12864));
  OAI21X1 g11076(.A0(n12864), .A1(n12859), .B0(n12334), .Y(n12865));
  XOR2X1  g11077(.A(n12535), .B(n10801), .Y(n12866));
  XOR2X1  g11078(.A(n12866), .B(n12559), .Y(n12867));
  NOR2X1  g11079(.A(n12861), .B(n12469), .Y(n12868));
  AOI22X1 g11080(.A0(P3_ADDR_REG_4__SCAN_IN), .A1(n12333), .B0(P3_REG3_REG_4__SCAN_IN), .B1(P3_U3151), .Y(n12869));
  OAI21X1 g11081(.A0(n12863), .A1(n12472), .B0(n12869), .Y(n12870));
  NOR2X1  g11082(.A(n12870), .B(n12868), .Y(n12871));
  OAI21X1 g11083(.A0(n12598), .A1(n12858), .B0(n12871), .Y(n12872));
  AOI21X1 g11084(.A0(n12867), .A1(n12783), .B0(n12872), .Y(n12873));
  NAND2X1 g11085(.A(n12873), .B(n12865), .Y(P3_U3186));
  NOR3X1  g11086(.A(n4574), .B(n10750), .C(n10589), .Y(n12875));
  NOR2X1  g11087(.A(n10703), .B(n10689), .Y(n12876));
  NOR2X1  g11088(.A(n12434), .B(n12433), .Y(n12877));
  OAI21X1 g11089(.A0(n12877), .A1(n12876), .B0(n12431), .Y(n12878));
  XOR2X1  g11090(.A(n10750), .B(n10759), .Y(n12879));
  XOR2X1  g11091(.A(n12879), .B(n12878), .Y(n12880));
  NOR2X1  g11092(.A(n10703), .B(n10685), .Y(n12881));
  NOR2X1  g11093(.A(n12363), .B(n12362), .Y(n12882));
  OAI21X1 g11094(.A0(n12882), .A1(n12881), .B0(n12360), .Y(n12883));
  XOR2X1  g11095(.A(n10750), .B(n10756), .Y(n12884));
  XOR2X1  g11096(.A(n12884), .B(n12883), .Y(n12885));
  OAI22X1 g11097(.A0(n12880), .A1(n10587), .B0(n12392), .B1(n12885), .Y(n12886));
  OAI21X1 g11098(.A0(n12886), .A1(n12875), .B0(n12334), .Y(n12887));
  NOR2X1  g11099(.A(n12554), .B(n10702), .Y(n12888));
  NOR2X1  g11100(.A(n12553), .B(n10703), .Y(n12889));
  NOR3X1  g11101(.A(n12889), .B(n12547), .C(n12544), .Y(n12890));
  XOR2X1  g11102(.A(n12550), .B(n10751), .Y(n12891));
  NOR3X1  g11103(.A(n12891), .B(n12890), .C(n12888), .Y(n12892));
  NOR2X1  g11104(.A(n12888), .B(n12548), .Y(n12893));
  OAI21X1 g11105(.A0(n12553), .A1(n10703), .B0(n12891), .Y(n12894));
  NOR2X1  g11106(.A(n12894), .B(n12893), .Y(n12895));
  OAI21X1 g11107(.A0(n12895), .A1(n12892), .B0(n12783), .Y(n12896));
  NOR2X1  g11108(.A(n12598), .B(n10750), .Y(n12897));
  NOR2X1  g11109(.A(n12880), .B(n12469), .Y(n12898));
  AOI22X1 g11110(.A0(P3_ADDR_REG_3__SCAN_IN), .A1(n12333), .B0(P3_REG3_REG_3__SCAN_IN), .B1(P3_U3151), .Y(n12899));
  OAI21X1 g11111(.A0(n12885), .A1(n12472), .B0(n12899), .Y(n12900));
  NOR3X1  g11112(.A(n12900), .B(n12898), .C(n12897), .Y(n12901));
  NAND3X1 g11113(.A(n12901), .B(n12896), .C(n12887), .Y(P3_U3185));
  NOR3X1  g11114(.A(n4574), .B(n10702), .C(n10589), .Y(n12903));
  XOR2X1  g11115(.A(n10702), .B(P3_REG1_REG_2__SCAN_IN), .Y(n12904));
  XOR2X1  g11116(.A(n12904), .B(n12877), .Y(n12905));
  XOR2X1  g11117(.A(n10702), .B(P3_REG2_REG_2__SCAN_IN), .Y(n12906));
  XOR2X1  g11118(.A(n12906), .B(n12882), .Y(n12907));
  OAI22X1 g11119(.A0(n12905), .A1(n10587), .B0(n12392), .B1(n12907), .Y(n12908));
  OAI21X1 g11120(.A0(n12908), .A1(n12903), .B0(n12334), .Y(n12909));
  NOR2X1  g11121(.A(n12905), .B(n12469), .Y(n12910));
  AOI22X1 g11122(.A0(P3_ADDR_REG_2__SCAN_IN), .A1(n12333), .B0(P3_REG3_REG_2__SCAN_IN), .B1(P3_U3151), .Y(n12911));
  OAI21X1 g11123(.A0(n12907), .A1(n12472), .B0(n12911), .Y(n12912));
  NOR2X1  g11124(.A(n12912), .B(n12910), .Y(n12913));
  XOR2X1  g11125(.A(n12553), .B(n10702), .Y(n12914));
  XOR2X1  g11126(.A(n12914), .B(n12548), .Y(n12915));
  AOI22X1 g11127(.A0(n12599), .A1(n10703), .B0(n12783), .B1(n12915), .Y(n12916));
  NAND3X1 g11128(.A(n12916), .B(n12913), .C(n12909), .Y(P3_U3184));
  NOR3X1  g11129(.A(n4574), .B(n10664), .C(n10589), .Y(n12918));
  XOR2X1  g11130(.A(n12432), .B(n10643), .Y(n12919));
  XOR2X1  g11131(.A(n12919), .B(n10665), .Y(n12920));
  XOR2X1  g11132(.A(n12361), .B(n10640), .Y(n12921));
  XOR2X1  g11133(.A(n12921), .B(n10665), .Y(n12922));
  OAI22X1 g11134(.A0(n12920), .A1(n10587), .B0(n12392), .B1(n12922), .Y(n12923));
  OAI21X1 g11135(.A0(n12923), .A1(n12918), .B0(n12334), .Y(n12924));
  NOR2X1  g11136(.A(n12598), .B(n10664), .Y(n12925));
  NOR2X1  g11137(.A(n12920), .B(n12469), .Y(n12926));
  NOR2X1  g11138(.A(n12922), .B(n12472), .Y(n12927));
  XOR2X1  g11139(.A(n12541), .B(n10664), .Y(n12928));
  XOR2X1  g11140(.A(n12928), .B(n12545), .Y(n12929));
  AOI22X1 g11141(.A0(P3_ADDR_REG_1__SCAN_IN), .A1(n12333), .B0(P3_REG3_REG_1__SCAN_IN), .B1(P3_U3151), .Y(n12930));
  OAI21X1 g11142(.A0(n12929), .A1(n12596), .B0(n12930), .Y(n12931));
  NOR4X1  g11143(.A(n12927), .B(n12926), .C(n12925), .D(n12931), .Y(n12932));
  NAND2X1 g11144(.A(n12932), .B(n12924), .Y(P3_U3183));
  AOI21X1 g11145(.A0(n10592), .A1(n10591), .B0(n10589), .Y(n12934));
  XOR2X1  g11146(.A(n10593), .B(n10609), .Y(n12935));
  XOR2X1  g11147(.A(n10593), .B(n10596), .Y(n12936));
  OAI22X1 g11148(.A0(n12935), .A1(n10587), .B0(n12392), .B1(n12936), .Y(n12937));
  OAI21X1 g11149(.A0(n12937), .A1(n12934), .B0(n12334), .Y(n12938));
  NAND2X1 g11150(.A(n12599), .B(n10593), .Y(n12939));
  NOR2X1  g11151(.A(n12935), .B(n12469), .Y(n12940));
  NOR2X1  g11152(.A(n12936), .B(n12472), .Y(n12941));
  NOR2X1  g11153(.A(n12332), .B(n1579), .Y(n12942));
  XOR2X1  g11154(.A(n12543), .B(n10593), .Y(n12943));
  OAI22X1 g11155(.A0(n12596), .A1(n12943), .B0(n10608), .B1(P3_STATE_REG_SCAN_IN), .Y(n12944));
  NOR4X1  g11156(.A(n12942), .B(n12941), .C(n12940), .D(n12944), .Y(n12945));
  NAND3X1 g11157(.A(n12945), .B(n12939), .C(n12938), .Y(P3_U3182));
  NAND2X1 g11158(.A(n12594), .B(P3_DATAO_REG_0__SCAN_IN), .Y(n12947));
  OAI21X1 g11159(.A0(n12594), .A1(n10615), .B0(n12947), .Y(P3_U3491));
  NAND2X1 g11160(.A(n12594), .B(P3_DATAO_REG_1__SCAN_IN), .Y(n12949));
  OAI21X1 g11161(.A0(n12594), .A1(n10645), .B0(n12949), .Y(P3_U3492));
  NAND2X1 g11162(.A(n12594), .B(P3_DATAO_REG_2__SCAN_IN), .Y(n12951));
  OAI21X1 g11163(.A0(n12594), .A1(n10691), .B0(n12951), .Y(P3_U3493));
  NAND2X1 g11164(.A(n12594), .B(P3_DATAO_REG_3__SCAN_IN), .Y(n12953));
  OAI21X1 g11165(.A0(n12594), .A1(n10761), .B0(n12953), .Y(P3_U3494));
  NAND2X1 g11166(.A(n12594), .B(P3_DATAO_REG_4__SCAN_IN), .Y(n12955));
  OAI21X1 g11167(.A0(n12594), .A1(n10816), .B0(n12955), .Y(P3_U3495));
  NAND2X1 g11168(.A(n12594), .B(P3_DATAO_REG_5__SCAN_IN), .Y(n12957));
  OAI21X1 g11169(.A0(n12594), .A1(n10859), .B0(n12957), .Y(P3_U3496));
  NAND2X1 g11170(.A(n12594), .B(P3_DATAO_REG_6__SCAN_IN), .Y(n12959));
  OAI21X1 g11171(.A0(n12594), .A1(n10914), .B0(n12959), .Y(P3_U3497));
  NAND2X1 g11172(.A(n12594), .B(P3_DATAO_REG_7__SCAN_IN), .Y(n12961));
  OAI21X1 g11173(.A0(n12594), .A1(n10957), .B0(n12961), .Y(P3_U3498));
  NAND2X1 g11174(.A(n12594), .B(P3_DATAO_REG_8__SCAN_IN), .Y(n12963));
  OAI21X1 g11175(.A0(n12594), .A1(n11061), .B0(n12963), .Y(P3_U3499));
  NAND2X1 g11176(.A(n12594), .B(P3_DATAO_REG_9__SCAN_IN), .Y(n12965));
  OAI21X1 g11177(.A0(n12594), .A1(n11045), .B0(n12965), .Y(P3_U3500));
  NAND2X1 g11178(.A(n12594), .B(P3_DATAO_REG_10__SCAN_IN), .Y(n12967));
  OAI21X1 g11179(.A0(n12594), .A1(n11095), .B0(n12967), .Y(P3_U3501));
  NAND2X1 g11180(.A(n12594), .B(P3_DATAO_REG_11__SCAN_IN), .Y(n12969));
  OAI21X1 g11181(.A0(n12594), .A1(n11140), .B0(n12969), .Y(P3_U3502));
  NAND2X1 g11182(.A(n12594), .B(P3_DATAO_REG_12__SCAN_IN), .Y(n12971));
  OAI21X1 g11183(.A0(n12594), .A1(n11207), .B0(n12971), .Y(P3_U3503));
  NAND2X1 g11184(.A(n12594), .B(P3_DATAO_REG_13__SCAN_IN), .Y(n12973));
  OAI21X1 g11185(.A0(n12594), .A1(n11266), .B0(n12973), .Y(P3_U3504));
  NAND2X1 g11186(.A(n12594), .B(P3_DATAO_REG_14__SCAN_IN), .Y(n12975));
  OAI21X1 g11187(.A0(n12594), .A1(n11344), .B0(n12975), .Y(P3_U3505));
  NAND2X1 g11188(.A(n12594), .B(P3_DATAO_REG_15__SCAN_IN), .Y(n12977));
  OAI21X1 g11189(.A0(n12594), .A1(n11337), .B0(n12977), .Y(P3_U3506));
  NAND2X1 g11190(.A(n12594), .B(P3_DATAO_REG_16__SCAN_IN), .Y(n12979));
  OAI21X1 g11191(.A0(n12594), .A1(n11377), .B0(n12979), .Y(P3_U3507));
  NAND2X1 g11192(.A(n12594), .B(P3_DATAO_REG_17__SCAN_IN), .Y(n12981));
  OAI21X1 g11193(.A0(n12594), .A1(n11485), .B0(n12981), .Y(P3_U3508));
  NAND2X1 g11194(.A(n12594), .B(P3_DATAO_REG_18__SCAN_IN), .Y(n12983));
  OAI21X1 g11195(.A0(n12594), .A1(n11498), .B0(n12983), .Y(P3_U3509));
  NAND2X1 g11196(.A(n12594), .B(P3_DATAO_REG_19__SCAN_IN), .Y(n12985));
  OAI21X1 g11197(.A0(n12594), .A1(n11521), .B0(n12985), .Y(P3_U3510));
  NAND2X1 g11198(.A(n12594), .B(P3_DATAO_REG_20__SCAN_IN), .Y(n12987));
  OAI21X1 g11199(.A0(n12594), .A1(n11562), .B0(n12987), .Y(P3_U3511));
  NAND2X1 g11200(.A(n12594), .B(P3_DATAO_REG_21__SCAN_IN), .Y(n12989));
  OAI21X1 g11201(.A0(n12594), .A1(n11607), .B0(n12989), .Y(P3_U3512));
  NAND2X1 g11202(.A(n12594), .B(P3_DATAO_REG_22__SCAN_IN), .Y(n12991));
  OAI21X1 g11203(.A0(n12594), .A1(n11645), .B0(n12991), .Y(P3_U3513));
  NAND2X1 g11204(.A(n12594), .B(P3_DATAO_REG_23__SCAN_IN), .Y(n12993));
  OAI21X1 g11205(.A0(n12594), .A1(n11736), .B0(n12993), .Y(P3_U3514));
  NAND2X1 g11206(.A(n12594), .B(P3_DATAO_REG_24__SCAN_IN), .Y(n12995));
  OAI21X1 g11207(.A0(n12594), .A1(n11731), .B0(n12995), .Y(P3_U3515));
  NAND2X1 g11208(.A(n12594), .B(P3_DATAO_REG_25__SCAN_IN), .Y(n12997));
  OAI21X1 g11209(.A0(n12594), .A1(n11777), .B0(n12997), .Y(P3_U3516));
  NAND2X1 g11210(.A(n12594), .B(P3_DATAO_REG_26__SCAN_IN), .Y(n12999));
  OAI21X1 g11211(.A0(n12594), .A1(n11820), .B0(n12999), .Y(P3_U3517));
  NAND2X1 g11212(.A(n12594), .B(P3_DATAO_REG_27__SCAN_IN), .Y(n13001));
  OAI21X1 g11213(.A0(n12594), .A1(n11910), .B0(n13001), .Y(P3_U3518));
  NAND2X1 g11214(.A(n12594), .B(P3_DATAO_REG_28__SCAN_IN), .Y(n13003));
  OAI21X1 g11215(.A0(n12594), .A1(n11903), .B0(n13003), .Y(P3_U3519));
  NAND2X1 g11216(.A(n12594), .B(P3_DATAO_REG_29__SCAN_IN), .Y(n13005));
  OAI21X1 g11217(.A0(n12594), .A1(n11949), .B0(n13005), .Y(P3_U3520));
  INVX1   g11218(.A(n11990), .Y(n13007));
  NAND2X1 g11219(.A(n12594), .B(P3_DATAO_REG_30__SCAN_IN), .Y(n13008));
  OAI21X1 g11220(.A0(n12594), .A1(n13007), .B0(n13008), .Y(P3_U3521));
  NAND2X1 g11221(.A(n12594), .B(P3_DATAO_REG_31__SCAN_IN), .Y(n13010));
  OAI21X1 g11222(.A0(n12594), .A1(n12010), .B0(n13010), .Y(P3_U3522));
  NOR2X1  g11223(.A(n10560), .B(n10445), .Y(n13013));
  NAND3X1 g11224(.A(n13013), .B(n10571), .C(n10562), .Y(n13014));
  OAI21X1 g11225(.A0(n10577), .A1(n10560), .B0(n13014), .Y(n13015));
  INVX1   g11226(.A(n13015), .Y(n13016));
  OAI22X1 g11227(.A0(n11991), .A1(n12010), .B0(n12326), .B1(n13016), .Y(n13017));
  OAI22X1 g11228(.A0(n11991), .A1(n12326), .B0(n12010), .B1(n13016), .Y(n13018));
  XOR2X1  g11229(.A(n13018), .B(n13017), .Y(n13019));
  OAI22X1 g11230(.A0(n11991), .A1(n12321), .B0(n13007), .B1(n13016), .Y(n13020));
  INVX1   g11231(.A(n11991), .Y(n13021));
  AOI22X1 g11232(.A0(n13021), .A1(n11990), .B0(n12016), .B1(n13015), .Y(n13022));
  AOI21X1 g11233(.A0(n13022), .A1(n13020), .B0(n13019), .Y(n13023));
  AOI21X1 g11234(.A0(n13021), .A1(n11950), .B0(n10445), .Y(n13024));
  OAI21X1 g11235(.A0(n13016), .A1(n11957), .B0(n13024), .Y(n13025));
  INVX1   g11236(.A(n10396), .Y(n13026));
  AOI21X1 g11237(.A0(n10403), .A1(n10402), .B0(n10398), .Y(n13027));
  NOR3X1  g11238(.A(n10400), .B(n10399), .C(n10397), .Y(n13028));
  OAI21X1 g11239(.A0(n13028), .A1(n13027), .B0(n1790), .Y(n13029));
  AOI21X1 g11240(.A0(n13029), .A1(n13026), .B0(n10590), .Y(n13030));
  NAND2X1 g11241(.A(n13021), .B(n13030), .Y(n13031));
  AOI22X1 g11242(.A0(n11950), .A1(n13015), .B0(n11902), .B1(n10445), .Y(n13032));
  AOI21X1 g11243(.A0(n13032), .A1(n13031), .B0(n13025), .Y(n13033));
  AOI22X1 g11244(.A0(n11902), .A1(n13015), .B0(n11863), .B1(n10445), .Y(n13034));
  INVX1   g11245(.A(n13034), .Y(n13035));
  AOI21X1 g11246(.A0(n13021), .A1(n11941), .B0(n13035), .Y(n13036));
  AOI21X1 g11247(.A0(n13021), .A1(n11902), .B0(n10445), .Y(n13037));
  OAI21X1 g11248(.A0(n13016), .A1(n11908), .B0(n13037), .Y(n13038));
  NOR2X1  g11249(.A(n13038), .B(n13036), .Y(n13039));
  AOI22X1 g11250(.A0(n11863), .A1(n13015), .B0(n11814), .B1(n10445), .Y(n13040));
  OAI21X1 g11251(.A0(n11991), .A1(n11869), .B0(n13040), .Y(n13041));
  AOI21X1 g11252(.A0(n13021), .A1(n11863), .B0(n10445), .Y(n13042));
  INVX1   g11253(.A(n13042), .Y(n13043));
  AOI21X1 g11254(.A0(n13015), .A1(n11915), .B0(n13043), .Y(n13044));
  AOI22X1 g11255(.A0(n11814), .A1(n13015), .B0(n11778), .B1(n10445), .Y(n13045));
  INVX1   g11256(.A(n13045), .Y(n13046));
  AOI21X1 g11257(.A0(n13021), .A1(n11821), .B0(n13046), .Y(n13047));
  INVX1   g11258(.A(n13047), .Y(n13048));
  AOI21X1 g11259(.A0(n13021), .A1(n11814), .B0(n10445), .Y(n13049));
  INVX1   g11260(.A(n13049), .Y(n13050));
  AOI21X1 g11261(.A0(n13015), .A1(n11821), .B0(n13050), .Y(n13051));
  AOI22X1 g11262(.A0(n13048), .A1(n13051), .B0(n13044), .B1(n13041), .Y(n13052));
  AOI22X1 g11263(.A0(n11778), .A1(n13015), .B0(n11730), .B1(n10445), .Y(n13053));
  OAI21X1 g11264(.A0(n11991), .A1(n11789), .B0(n13053), .Y(n13054));
  AOI21X1 g11265(.A0(n13021), .A1(n11778), .B0(n10445), .Y(n13055));
  INVX1   g11266(.A(n13055), .Y(n13056));
  AOI21X1 g11267(.A0(n13015), .A1(n11808), .B0(n13056), .Y(n13057));
  NAND2X1 g11268(.A(n13057), .B(n13054), .Y(n13058));
  AOI21X1 g11269(.A0(n13021), .A1(n11730), .B0(n10445), .Y(n13059));
  OAI21X1 g11270(.A0(n13016), .A1(n12280), .B0(n13059), .Y(n13060));
  OAI22X1 g11271(.A0(n11731), .A1(n13016), .B0(n11736), .B1(n10446), .Y(n13061));
  AOI21X1 g11272(.A0(n13021), .A1(n11737), .B0(n13061), .Y(n13062));
  NAND2X1 g11273(.A(n13062), .B(n13060), .Y(n13063));
  AOI22X1 g11274(.A0(n11473), .A1(n13015), .B0(n11424), .B1(n10445), .Y(n13064));
  OAI21X1 g11275(.A0(n11991), .A1(n11483), .B0(n13064), .Y(n13065));
  OAI21X1 g11276(.A0(n11991), .A1(n11498), .B0(n10446), .Y(n13066));
  AOI21X1 g11277(.A0(n13015), .A1(n11508), .B0(n13066), .Y(n13067));
  AOI22X1 g11278(.A0(n11424), .A1(n13015), .B0(n11369), .B1(n10445), .Y(n13068));
  OAI21X1 g11279(.A0(n11991), .A1(n11435), .B0(n13068), .Y(n13069));
  OAI21X1 g11280(.A0(n11991), .A1(n11485), .B0(n10446), .Y(n13070));
  AOI21X1 g11281(.A0(n13015), .A1(n11436), .B0(n13070), .Y(n13071));
  NAND2X1 g11282(.A(n13071), .B(n13069), .Y(n13072));
  AOI22X1 g11283(.A0(n11369), .A1(n13015), .B0(n11331), .B1(n10445), .Y(n13073));
  OAI21X1 g11284(.A0(n11991), .A1(n11391), .B0(n13073), .Y(n13074));
  OAI21X1 g11285(.A0(n11991), .A1(n11377), .B0(n10446), .Y(n13075));
  AOI21X1 g11286(.A0(n13015), .A1(n11382), .B0(n13075), .Y(n13076));
  AOI21X1 g11287(.A0(n13015), .A1(n11006), .B0(n10445), .Y(n13077));
  OAI21X1 g11288(.A0(n11991), .A1(n11061), .B0(n13077), .Y(n13078));
  OAI22X1 g11289(.A0(n12176), .A1(n11991), .B0(n10957), .B1(n10446), .Y(n13079));
  AOI21X1 g11290(.A0(n13015), .A1(n10996), .B0(n13079), .Y(n13080));
  NAND2X1 g11291(.A(n13080), .B(n13078), .Y(n13081));
  OAI21X1 g11292(.A0(n10956), .A1(n10954), .B0(n13021), .Y(n13082));
  AOI21X1 g11293(.A0(n13015), .A1(n10962), .B0(n10445), .Y(n13083));
  AOI22X1 g11294(.A0(n10962), .A1(n13021), .B0(n10897), .B1(n10445), .Y(n13084));
  OAI21X1 g11295(.A0(n13016), .A1(n10957), .B0(n13084), .Y(n13085));
  AOI21X1 g11296(.A0(n13083), .A1(n13082), .B0(n13085), .Y(n13086));
  OAI22X1 g11297(.A0(n10705), .A1(n11991), .B0(n10645), .B1(n10446), .Y(n13087));
  AOI21X1 g11298(.A0(n13015), .A1(n10709), .B0(n13087), .Y(n13088));
  AOI21X1 g11299(.A0(n13015), .A1(n10711), .B0(n10445), .Y(n13089));
  OAI21X1 g11300(.A0(n11991), .A1(n10691), .B0(n13089), .Y(n13090));
  AOI22X1 g11301(.A0(n10788), .A1(n13021), .B0(n10709), .B1(n10445), .Y(n13091));
  OAI21X1 g11302(.A0(n13016), .A1(n10761), .B0(n13091), .Y(n13092));
  OAI21X1 g11303(.A0(n13016), .A1(n10753), .B0(n10446), .Y(n13093));
  AOI21X1 g11304(.A0(n13021), .A1(n10738), .B0(n13093), .Y(n13094));
  NAND2X1 g11305(.A(n13094), .B(n13092), .Y(n13095));
  OAI21X1 g11306(.A0(n13090), .A1(n13088), .B0(n13095), .Y(n13096));
  AOI21X1 g11307(.A0(n13015), .A1(n10720), .B0(n10445), .Y(n13097));
  OAI21X1 g11308(.A0(n11991), .A1(n10645), .B0(n13097), .Y(n13098));
  OAI22X1 g11309(.A0(n10667), .A1(n11991), .B0(n10615), .B1(n10446), .Y(n13099));
  AOI21X1 g11310(.A0(n13015), .A1(n10662), .B0(n13099), .Y(n13100));
  NOR2X1  g11311(.A(n13100), .B(n13098), .Y(n13101));
  OAI21X1 g11312(.A0(n10614), .A1(n10607), .B0(n13021), .Y(n13102));
  AOI21X1 g11313(.A0(n13015), .A1(n10595), .B0(n10445), .Y(n13103));
  NAND4X1 g11314(.A(n13102), .B(n13013), .C(n10563), .D(n13103), .Y(n13104));
  AOI22X1 g11315(.A0(n13021), .A1(n10595), .B0(n10658), .B1(n13015), .Y(n13105));
  AOI22X1 g11316(.A0(n13102), .A1(n13103), .B0(n13013), .B1(n10563), .Y(n13106));
  OAI21X1 g11317(.A0(n13106), .A1(n13105), .B0(n13104), .Y(n13107));
  NOR3X1  g11318(.A(n13107), .B(n13101), .C(n13096), .Y(n13108));
  AOI22X1 g11319(.A0(n13098), .A1(n13100), .B0(n13090), .B1(n13088), .Y(n13109));
  NOR2X1  g11320(.A(n13109), .B(n13096), .Y(n13110));
  AOI21X1 g11321(.A0(n13015), .A1(n10919), .B0(n10445), .Y(n13111));
  OAI21X1 g11322(.A0(n11991), .A1(n10914), .B0(n13111), .Y(n13112));
  OAI22X1 g11323(.A0(n10932), .A1(n11991), .B0(n10859), .B1(n10446), .Y(n13113));
  AOI21X1 g11324(.A0(n13015), .A1(n10897), .B0(n13113), .Y(n13114));
  NAND2X1 g11325(.A(n13114), .B(n13112), .Y(n13115));
  OAI21X1 g11326(.A0(n13016), .A1(n10861), .B0(n10446), .Y(n13116));
  AOI21X1 g11327(.A0(n13021), .A1(n10844), .B0(n13116), .Y(n13117));
  AOI22X1 g11328(.A0(n10855), .A1(n13021), .B0(n10793), .B1(n10445), .Y(n13118));
  OAI21X1 g11329(.A0(n13016), .A1(n10859), .B0(n13118), .Y(n13119));
  OAI21X1 g11330(.A0(n13119), .A1(n13117), .B0(n13115), .Y(n13120));
  OAI21X1 g11331(.A0(n13016), .A1(n10803), .B0(n10446), .Y(n13121));
  AOI21X1 g11332(.A0(n13021), .A1(n10793), .B0(n13121), .Y(n13122));
  AOI22X1 g11333(.A0(n10835), .A1(n13021), .B0(n10738), .B1(n10445), .Y(n13123));
  OAI21X1 g11334(.A0(n13016), .A1(n10816), .B0(n13123), .Y(n13124));
  OAI22X1 g11335(.A0(n13122), .A1(n13124), .B0(n13094), .B1(n13092), .Y(n13125));
  NOR4X1  g11336(.A(n13120), .B(n13110), .C(n13108), .D(n13125), .Y(n13126));
  NAND2X1 g11337(.A(n13124), .B(n13122), .Y(n13127));
  NOR2X1  g11338(.A(n13127), .B(n13120), .Y(n13128));
  NAND2X1 g11339(.A(n13119), .B(n13117), .Y(n13129));
  AOI21X1 g11340(.A0(n13114), .A1(n13112), .B0(n13129), .Y(n13130));
  NAND3X1 g11341(.A(n13085), .B(n13083), .C(n13082), .Y(n13131));
  OAI21X1 g11342(.A0(n13114), .A1(n13112), .B0(n13131), .Y(n13132));
  NOR4X1  g11343(.A(n13130), .B(n13128), .C(n13126), .D(n13132), .Y(n13133));
  OAI22X1 g11344(.A0(n13086), .A1(n13133), .B0(n13080), .B1(n13078), .Y(n13134));
  AOI22X1 g11345(.A0(n11050), .A1(n13021), .B0(n10996), .B1(n10445), .Y(n13135));
  OAI21X1 g11346(.A0(n13016), .A1(n11045), .B0(n13135), .Y(n13136));
  INVX1   g11347(.A(n13136), .Y(n13137));
  AOI21X1 g11348(.A0(n13015), .A1(n11050), .B0(n10445), .Y(n13138));
  OAI21X1 g11349(.A0(n11991), .A1(n11045), .B0(n13138), .Y(n13139));
  NOR2X1  g11350(.A(n13139), .B(n13137), .Y(n13140));
  AOI21X1 g11351(.A0(n13134), .A1(n13081), .B0(n13140), .Y(n13141));
  OAI21X1 g11352(.A0(n11991), .A1(n11207), .B0(n10446), .Y(n13142));
  AOI21X1 g11353(.A0(n13015), .A1(n11232), .B0(n13142), .Y(n13143));
  AOI22X1 g11354(.A0(n11232), .A1(n13021), .B0(n11131), .B1(n10445), .Y(n13144));
  OAI21X1 g11355(.A0(n13016), .A1(n11207), .B0(n13144), .Y(n13145));
  NOR2X1  g11356(.A(n13145), .B(n13143), .Y(n13146));
  AOI21X1 g11357(.A0(n13021), .A1(n11131), .B0(n10445), .Y(n13147));
  OAI21X1 g11358(.A0(n13016), .A1(n11150), .B0(n13147), .Y(n13148));
  AOI22X1 g11359(.A0(n11145), .A1(n13021), .B0(n11086), .B1(n10445), .Y(n13149));
  OAI21X1 g11360(.A0(n13016), .A1(n11140), .B0(n13149), .Y(n13150));
  INVX1   g11361(.A(n13150), .Y(n13151));
  AOI21X1 g11362(.A0(n13151), .A1(n13148), .B0(n13146), .Y(n13152));
  AOI21X1 g11363(.A0(n13021), .A1(n11086), .B0(n10445), .Y(n13153));
  OAI21X1 g11364(.A0(n13016), .A1(n11100), .B0(n13153), .Y(n13154));
  AOI22X1 g11365(.A0(n11102), .A1(n13021), .B0(n11036), .B1(n10445), .Y(n13155));
  OAI21X1 g11366(.A0(n13016), .A1(n11095), .B0(n13155), .Y(n13156));
  INVX1   g11367(.A(n13156), .Y(n13157));
  AOI22X1 g11368(.A0(n13154), .A1(n13157), .B0(n13139), .B1(n13137), .Y(n13158));
  NAND2X1 g11369(.A(n13158), .B(n13152), .Y(n13159));
  OAI22X1 g11370(.A0(n11337), .A1(n13016), .B0(n11344), .B1(n10446), .Y(n13160));
  AOI21X1 g11371(.A0(n13021), .A1(n11342), .B0(n13160), .Y(n13161));
  AOI21X1 g11372(.A0(n13021), .A1(n11331), .B0(n10445), .Y(n13162));
  OAI21X1 g11373(.A0(n13016), .A1(n11390), .B0(n13162), .Y(n13163));
  OAI22X1 g11374(.A0(n11344), .A1(n13016), .B0(n11266), .B1(n10446), .Y(n13164));
  AOI21X1 g11375(.A0(n13021), .A1(n11323), .B0(n13164), .Y(n13165));
  AOI21X1 g11376(.A0(n13021), .A1(n11292), .B0(n10445), .Y(n13166));
  OAI21X1 g11377(.A0(n13016), .A1(n11302), .B0(n13166), .Y(n13167));
  OAI22X1 g11378(.A0(n13165), .A1(n13167), .B0(n13163), .B1(n13161), .Y(n13168));
  NOR2X1  g11379(.A(n13157), .B(n13154), .Y(n13169));
  NAND2X1 g11380(.A(n13169), .B(n13152), .Y(n13170));
  NOR2X1  g11381(.A(n13151), .B(n13148), .Y(n13171));
  OAI21X1 g11382(.A0(n13145), .A1(n13143), .B0(n13171), .Y(n13172));
  AOI22X1 g11383(.A0(n11251), .A1(n13021), .B0(n11191), .B1(n10445), .Y(n13173));
  OAI21X1 g11384(.A0(n13016), .A1(n11266), .B0(n13173), .Y(n13174));
  OAI21X1 g11385(.A0(n11991), .A1(n11266), .B0(n10446), .Y(n13175));
  AOI21X1 g11386(.A0(n13015), .A1(n11251), .B0(n13175), .Y(n13176));
  AOI22X1 g11387(.A0(n13174), .A1(n13176), .B0(n13145), .B1(n13143), .Y(n13177));
  NAND3X1 g11388(.A(n13177), .B(n13172), .C(n13170), .Y(n13178));
  NOR2X1  g11389(.A(n13178), .B(n13168), .Y(n13179));
  OAI21X1 g11390(.A0(n13159), .A1(n13141), .B0(n13179), .Y(n13180));
  NOR3X1  g11391(.A(n13176), .B(n13174), .C(n13168), .Y(n13181));
  NOR2X1  g11392(.A(n13076), .B(n13074), .Y(n13182));
  NOR2X1  g11393(.A(n13163), .B(n13161), .Y(n13183));
  NAND2X1 g11394(.A(n13163), .B(n13161), .Y(n13184));
  NAND2X1 g11395(.A(n13167), .B(n13165), .Y(n13185));
  OAI21X1 g11396(.A0(n13185), .A1(n13183), .B0(n13184), .Y(n13186));
  NOR3X1  g11397(.A(n13186), .B(n13182), .C(n13181), .Y(n13187));
  AOI22X1 g11398(.A0(n13180), .A1(n13187), .B0(n13076), .B1(n13074), .Y(n13188));
  NOR2X1  g11399(.A(n13071), .B(n13069), .Y(n13189));
  OAI21X1 g11400(.A0(n13189), .A1(n13188), .B0(n13072), .Y(n13190));
  OAI21X1 g11401(.A0(n13190), .A1(n13067), .B0(n13065), .Y(n13191));
  INVX1   g11402(.A(n11608), .Y(n13192));
  AOI21X1 g11403(.A0(n13021), .A1(n11601), .B0(n10445), .Y(n13193));
  OAI21X1 g11404(.A0(n13016), .A1(n13192), .B0(n13193), .Y(n13194));
  AOI22X1 g11405(.A0(n11601), .A1(n13015), .B0(n11554), .B1(n10445), .Y(n13195));
  OAI21X1 g11406(.A0(n11991), .A1(n13192), .B0(n13195), .Y(n13196));
  INVX1   g11407(.A(n13196), .Y(n13197));
  AOI21X1 g11408(.A0(n13021), .A1(n11554), .B0(n10445), .Y(n13198));
  INVX1   g11409(.A(n13198), .Y(n13199));
  AOI21X1 g11410(.A0(n13015), .A1(n11560), .B0(n13199), .Y(n13200));
  AOI22X1 g11411(.A0(n11554), .A1(n13015), .B0(n11515), .B1(n10445), .Y(n13201));
  OAI21X1 g11412(.A0(n11991), .A1(n11563), .B0(n13201), .Y(n13202));
  AOI21X1 g11413(.A0(n13021), .A1(n11515), .B0(n10445), .Y(n13203));
  INVX1   g11414(.A(n13203), .Y(n13204));
  AOI21X1 g11415(.A0(n13015), .A1(n11523), .B0(n13204), .Y(n13205));
  AOI22X1 g11416(.A0(n11515), .A1(n13015), .B0(n11473), .B1(n10445), .Y(n13206));
  OAI21X1 g11417(.A0(n11991), .A1(n11585), .B0(n13206), .Y(n13207));
  AOI22X1 g11418(.A0(n13205), .A1(n13207), .B0(n13202), .B1(n13200), .Y(n13208));
  OAI21X1 g11419(.A0(n13197), .A1(n13194), .B0(n13208), .Y(n13209));
  AOI21X1 g11420(.A0(n13190), .A1(n13067), .B0(n13209), .Y(n13210));
  NAND2X1 g11421(.A(n13210), .B(n13191), .Y(n13211));
  INVX1   g11422(.A(n11699), .Y(n13212));
  OAI21X1 g11423(.A0(n11991), .A1(n11736), .B0(n10446), .Y(n13213));
  AOI21X1 g11424(.A0(n13015), .A1(n13212), .B0(n13213), .Y(n13214));
  AOI22X1 g11425(.A0(n11691), .A1(n13015), .B0(n11639), .B1(n10445), .Y(n13215));
  OAI21X1 g11426(.A0(n11991), .A1(n11699), .B0(n13215), .Y(n13216));
  NOR2X1  g11427(.A(n13216), .B(n13214), .Y(n13217));
  OAI21X1 g11428(.A0(n11991), .A1(n11645), .B0(n10446), .Y(n13218));
  AOI21X1 g11429(.A0(n13015), .A1(n11646), .B0(n13218), .Y(n13219));
  AOI22X1 g11430(.A0(n11639), .A1(n13015), .B0(n11601), .B1(n10445), .Y(n13220));
  OAI21X1 g11431(.A0(n11991), .A1(n11704), .B0(n13220), .Y(n13221));
  NOR2X1  g11432(.A(n13221), .B(n13219), .Y(n13222));
  NAND2X1 g11433(.A(n13197), .B(n13194), .Y(n13223));
  NAND2X1 g11434(.A(n13202), .B(n13200), .Y(n13224));
  NOR2X1  g11435(.A(n13207), .B(n13205), .Y(n13225));
  NAND2X1 g11436(.A(n13225), .B(n13224), .Y(n13226));
  OAI21X1 g11437(.A0(n13202), .A1(n13200), .B0(n13226), .Y(n13227));
  OAI21X1 g11438(.A0(n13197), .A1(n13194), .B0(n13227), .Y(n13228));
  NAND2X1 g11439(.A(n13228), .B(n13223), .Y(n13229));
  NOR3X1  g11440(.A(n13229), .B(n13222), .C(n13217), .Y(n13230));
  NAND3X1 g11441(.A(n13230), .B(n13211), .C(n13063), .Y(n13231));
  NOR2X1  g11442(.A(n13062), .B(n13060), .Y(n13232));
  AOI22X1 g11443(.A0(n13219), .A1(n13221), .B0(n13216), .B1(n13214), .Y(n13233));
  NOR2X1  g11444(.A(n13233), .B(n13217), .Y(n13234));
  AOI21X1 g11445(.A0(n13234), .A1(n13063), .B0(n13232), .Y(n13235));
  NAND4X1 g11446(.A(n13231), .B(n13058), .C(n13052), .D(n13235), .Y(n13236));
  NOR3X1  g11447(.A(n13236), .B(n13039), .C(n13033), .Y(n13237));
  NAND2X1 g11448(.A(n13237), .B(n13023), .Y(n13238));
  INVX1   g11449(.A(n13024), .Y(n13239));
  AOI21X1 g11450(.A0(n13015), .A1(n13030), .B0(n13239), .Y(n13240));
  OAI21X1 g11451(.A0(n11991), .A1(n11957), .B0(n13032), .Y(n13241));
  OAI21X1 g11452(.A0(n11991), .A1(n11908), .B0(n13034), .Y(n13242));
  INVX1   g11453(.A(n13037), .Y(n13243));
  AOI21X1 g11454(.A0(n13015), .A1(n11941), .B0(n13243), .Y(n13244));
  NAND2X1 g11455(.A(n13244), .B(n13242), .Y(n13245));
  NOR2X1  g11456(.A(n13244), .B(n13242), .Y(n13246));
  NOR2X1  g11457(.A(n13044), .B(n13041), .Y(n13247));
  AOI21X1 g11458(.A0(n13247), .A1(n13245), .B0(n13246), .Y(n13248));
  AOI21X1 g11459(.A0(n13248), .A1(n13240), .B0(n13241), .Y(n13249));
  NAND2X1 g11460(.A(n13241), .B(n13240), .Y(n13250));
  NAND2X1 g11461(.A(n13038), .B(n13036), .Y(n13251));
  INVX1   g11462(.A(n13040), .Y(n13252));
  AOI21X1 g11463(.A0(n13021), .A1(n11915), .B0(n13252), .Y(n13253));
  OAI21X1 g11464(.A0(n13016), .A1(n11869), .B0(n13042), .Y(n13254));
  NAND2X1 g11465(.A(n13254), .B(n13253), .Y(n13255));
  OAI21X1 g11466(.A0(n13255), .A1(n13039), .B0(n13251), .Y(n13256));
  INVX1   g11467(.A(n13051), .Y(n13257));
  OAI22X1 g11468(.A0(n13047), .A1(n13257), .B0(n13254), .B1(n13253), .Y(n13258));
  NOR2X1  g11469(.A(n13057), .B(n13054), .Y(n13259));
  AOI21X1 g11470(.A0(n13257), .A1(n13047), .B0(n13259), .Y(n13260));
  NOR3X1  g11471(.A(n13260), .B(n13258), .C(n13039), .Y(n13261));
  AOI22X1 g11472(.A0(n13256), .A1(n13025), .B0(n13250), .B1(n13261), .Y(n13262));
  OAI21X1 g11473(.A0(n13022), .A1(n13020), .B0(n13262), .Y(n13263));
  OAI21X1 g11474(.A0(n13263), .A1(n13249), .B0(n13023), .Y(n13264));
  AOI22X1 g11475(.A0(n13021), .A1(n12025), .B0(n12009), .B1(n13015), .Y(n13265));
  NOR3X1  g11476(.A(n10580), .B(n10560), .C(n10446), .Y(n13266));
  NOR3X1  g11477(.A(n13266), .B(n13265), .C(n13017), .Y(n13267));
  AOI21X1 g11478(.A0(n13266), .A1(n13017), .B0(n13267), .Y(n13269));
  XOR2X1  g11479(.A(n11991), .B(n10571), .Y(n13270));
  INVX1   g11480(.A(n13270), .Y(n13271));
  NAND4X1 g11481(.A(n13269), .B(n13264), .C(n13238), .D(n13271), .Y(n13272));
  XOR2X1  g11482(.A(n13265), .B(n13017), .Y(n13273));
  AOI22X1 g11483(.A0(n13021), .A1(n12016), .B0(n11990), .B1(n13015), .Y(n13274));
  OAI22X1 g11484(.A0(n11991), .A1(n13007), .B0(n12321), .B1(n13016), .Y(n13275));
  OAI21X1 g11485(.A0(n13275), .A1(n13274), .B0(n13273), .Y(n13276));
  NOR4X1  g11486(.A(n13039), .B(n13033), .C(n13276), .D(n13236), .Y(n13277));
  NOR2X1  g11487(.A(n13022), .B(n13020), .Y(n13278));
  OAI22X1 g11488(.A0(n13054), .A1(n13057), .B0(n13051), .B1(n13048), .Y(n13279));
  NAND3X1 g11489(.A(n13279), .B(n13052), .C(n13245), .Y(n13280));
  OAI22X1 g11490(.A0(n13248), .A1(n13240), .B0(n13033), .B1(n13280), .Y(n13281));
  NOR3X1  g11491(.A(n13281), .B(n13278), .C(n13249), .Y(n13282));
  OAI21X1 g11492(.A0(n13282), .A1(n13276), .B0(n13269), .Y(n13283));
  OAI21X1 g11493(.A0(n13283), .A1(n13277), .B0(n13270), .Y(n13284));
  NAND3X1 g11494(.A(n13284), .B(n13272), .C(n10575), .Y(n13285));
  NAND4X1 g11495(.A(n10678), .B(n10581), .C(n10528), .D(n10589), .Y(n13286));
  NOR3X1  g11496(.A(n13286), .B(n13283), .C(n13277), .Y(n13287));
  NAND2X1 g11497(.A(n12009), .B(n11990), .Y(n13290));
  AOI22X1 g11498(.A0(n12009), .A1(n12326), .B0(n12016), .B1(n13290), .Y(n13291));
  AOI22X1 g11499(.A0(n11903), .A1(n11941), .B0(n11915), .B1(n11910), .Y(n13294));
  OAI21X1 g11500(.A0(n11950), .A1(n11957), .B0(n13294), .Y(n13295));
  NOR2X1  g11501(.A(n11884), .B(n13295), .Y(n13297));
  NAND2X1 g11502(.A(n13297), .B(n13291), .Y(n13298));
  NOR4X1  g11503(.A(n12016), .B(n12010), .C(n13007), .D(n12326), .Y(n13300));
  AOI21X1 g11504(.A0(n12010), .A1(n12025), .B0(n13300), .Y(n13301));
  NAND2X1 g11505(.A(n11869), .B(n11863), .Y(n13302));
  NOR2X1  g11506(.A(n13302), .B(n13295), .Y(n13303));
  AOI21X1 g11507(.A0(n11949), .A1(n13030), .B0(n11960), .Y(n13305));
  OAI21X1 g11508(.A0(n13305), .A1(n13303), .B0(n13291), .Y(n13306));
  NOR2X1  g11509(.A(n13030), .B(n11949), .Y(n13307));
  NAND2X1 g11510(.A(n11789), .B(n11778), .Y(n13309));
  NAND2X1 g11511(.A(n11699), .B(n11691), .Y(n13311));
  AOI22X1 g11512(.A0(n11645), .A1(n11646), .B0(n11608), .B1(n11607), .Y(n13312));
  NAND2X1 g11513(.A(n11625), .B(n13312), .Y(n13314));
  NOR2X1  g11514(.A(n11646), .B(n11645), .Y(n13317));
  AOI21X1 g11515(.A0(n11648), .A1(n11755), .B0(n13317), .Y(n13318));
  NAND3X1 g11516(.A(n13318), .B(n13314), .C(n13311), .Y(n13319));
  AOI22X1 g11517(.A0(n11515), .A1(n11585), .B0(n11483), .B1(n11473), .Y(n13320));
  NOR2X1  g11518(.A(n11435), .B(n11424), .Y(n13321));
  NAND2X1 g11519(.A(n13321), .B(n13320), .Y(n13322));
  NOR2X1  g11520(.A(n11483), .B(n11473), .Y(n13324));
  OAI22X1 g11521(.A0(n11554), .A1(n11563), .B0(n11585), .B1(n11515), .Y(n13325));
  AOI21X1 g11522(.A0(n13324), .A1(n11584), .B0(n13325), .Y(n13326));
  NAND3X1 g11523(.A(n13326), .B(n13322), .C(n13312), .Y(n13327));
  NAND2X1 g11524(.A(n11302), .B(n11292), .Y(n13329));
  AOI22X1 g11525(.A0(n10816), .A1(n10835), .B0(n10788), .B1(n10761), .Y(n13330));
  OAI22X1 g11526(.A0(n10761), .A1(n10788), .B0(n10711), .B1(n10691), .Y(n13331));
  NAND2X1 g11527(.A(n13331), .B(n13330), .Y(n13332));
  AOI22X1 g11528(.A0(n10946), .A1(n10977), .B0(n10932), .B1(n10897), .Y(n13333));
  AOI22X1 g11529(.A0(n10844), .A1(n10861), .B0(n10803), .B1(n10793), .Y(n13334));
  NAND3X1 g11530(.A(n13334), .B(n13333), .C(n13332), .Y(n13335));
  NAND2X1 g11531(.A(n10870), .B(n13333), .Y(n13337));
  OAI22X1 g11532(.A0(n11086), .A1(n11100), .B0(n11092), .B1(n11036), .Y(n13338));
  NOR2X1  g11533(.A(n11063), .B(n13338), .Y(n13340));
  OAI21X1 g11534(.A0(n10957), .A1(n10962), .B0(n10933), .Y(n13343));
  NAND4X1 g11535(.A(n13340), .B(n13337), .C(n13335), .D(n13343), .Y(n13344));
  AOI22X1 g11536(.A0(n10691), .A1(n10711), .B0(n10720), .B1(n10645), .Y(n13345));
  NAND2X1 g11537(.A(n13345), .B(n13343), .Y(n13346));
  NAND2X1 g11538(.A(n10615), .B(n10595), .Y(n13348));
  OAI21X1 g11539(.A0(n13348), .A1(n10721), .B0(n13330), .Y(n13349));
  NOR2X1  g11540(.A(n13349), .B(n13346), .Y(n13350));
  NAND3X1 g11541(.A(n13350), .B(n13340), .C(n13337), .Y(n13351));
  NAND2X1 g11542(.A(n12176), .B(n10996), .Y(n13352));
  NOR2X1  g11543(.A(n13352), .B(n13338), .Y(n13353));
  NAND2X1 g11544(.A(n11092), .B(n11036), .Y(n13355));
  NOR2X1  g11545(.A(n13355), .B(n11139), .Y(n13356));
  AOI22X1 g11546(.A0(n11239), .A1(n11261), .B0(n11202), .B1(n11191), .Y(n13357));
  AOI22X1 g11547(.A0(n11131), .A1(n11150), .B0(n11100), .B1(n11086), .Y(n13358));
  NAND2X1 g11548(.A(n13358), .B(n13357), .Y(n13359));
  NOR3X1  g11549(.A(n13359), .B(n13356), .C(n13353), .Y(n13360));
  NAND3X1 g11550(.A(n13360), .B(n13351), .C(n13344), .Y(n13361));
  NAND2X1 g11551(.A(n11151), .B(n13357), .Y(n13363));
  NOR2X1  g11552(.A(n11202), .B(n11191), .Y(n13365));
  OAI22X1 g11553(.A0(n11292), .A1(n11302), .B0(n11261), .B1(n11239), .Y(n13366));
  AOI21X1 g11554(.A0(n13365), .A1(n11315), .B0(n13366), .Y(n13367));
  NAND3X1 g11555(.A(n13367), .B(n13363), .C(n13361), .Y(n13368));
  AOI21X1 g11556(.A0(n13368), .A1(n13329), .B0(n11387), .Y(n13370));
  OAI21X1 g11557(.A0(n13370), .A1(n11375), .B0(n11388), .Y(n13372));
  INVX1   g11558(.A(n13320), .Y(n13373));
  OAI22X1 g11559(.A0(n11485), .A1(n11436), .B0(n11382), .B1(n11377), .Y(n13374));
  NOR2X1  g11560(.A(n13374), .B(n13373), .Y(n13375));
  AOI21X1 g11561(.A0(n13375), .A1(n13372), .B0(n13327), .Y(n13376));
  NOR3X1  g11562(.A(n13376), .B(n13319), .C(n11800), .Y(n13377));
  NAND2X1 g11563(.A(n13377), .B(n13309), .Y(n13378));
  AOI22X1 g11564(.A0(n11731), .A1(n11737), .B0(n13212), .B1(n11736), .Y(n13380));
  NOR2X1  g11565(.A(n13380), .B(n11800), .Y(n13381));
  NAND2X1 g11566(.A(n13381), .B(n13309), .Y(n13382));
  NAND3X1 g11567(.A(n13382), .B(n11825), .C(n13378), .Y(n13383));
  NOR3X1  g11568(.A(n13383), .B(n11888), .C(n13295), .Y(n13384));
  OAI21X1 g11569(.A0(n13384), .A1(n13307), .B0(n13291), .Y(n13385));
  NAND4X1 g11570(.A(n13306), .B(n13301), .C(n13298), .D(n13385), .Y(n13386));
  NAND2X1 g11571(.A(n13386), .B(n10622), .Y(n13387));
  NAND4X1 g11572(.A(n12321), .B(n12009), .C(n11990), .D(n12025), .Y(n13388));
  OAI21X1 g11573(.A0(n12009), .A1(n12326), .B0(n13388), .Y(n13389));
  AOI21X1 g11574(.A0(n13297), .A1(n13291), .B0(n13389), .Y(n13390));
  NAND4X1 g11575(.A(n13306), .B(n13390), .C(n10626), .D(n13385), .Y(n13391));
  NOR2X1  g11576(.A(n11992), .B(n10587), .Y(n13392));
  AOI21X1 g11577(.A0(n13392), .A1(n10581), .B0(n10446), .Y(n13393));
  OAI21X1 g11578(.A0(n10563), .A1(n10445), .B0(n12329), .Y(n13394));
  OAI21X1 g11579(.A0(n13394), .A1(n13393), .B0(P3_B_REG_SCAN_IN), .Y(n13395));
  XOR2X1  g11580(.A(n12321), .B(n13007), .Y(n13396));
  XOR2X1  g11581(.A(n12326), .B(n12010), .Y(n13397));
  XOR2X1  g11582(.A(n11699), .B(n11736), .Y(n13401));
  XOR2X1  g11583(.A(n11646), .B(n11639), .Y(n13402));
  XOR2X1  g11584(.A(n11435), .B(n11485), .Y(n13405));
  XOR2X1  g11585(.A(n10705), .B(n10691), .Y(n13406));
  NOR2X1  g11586(.A(n13406), .B(n10672), .Y(n13407));
  XOR2X1  g11587(.A(n11102), .B(n11086), .Y(n13408));
  NOR4X1  g11588(.A(n11166), .B(n10817), .C(n10762), .D(n13408), .Y(n13409));
  NAND2X1 g11589(.A(n13409), .B(n13407), .Y(n13410));
  XOR2X1  g11590(.A(n11302), .B(n11344), .Y(n13411));
  XOR2X1  g11591(.A(n10615), .B(n10635), .Y(n13412));
  NOR2X1  g11592(.A(n13412), .B(n11208), .Y(n13413));
  NAND3X1 g11593(.A(n10877), .B(n13413), .C(n10920), .Y(n13415));
  INVX1   g11594(.A(n11007), .Y(n13416));
  NAND4X1 g11595(.A(n11267), .B(n11051), .C(n13416), .D(n10963), .Y(n13419));
  NOR4X1  g11596(.A(n13415), .B(n13411), .C(n13410), .D(n13419), .Y(n13420));
  OAI21X1 g11597(.A0(n11399), .A1(n11398), .B0(n13420), .Y(n13421));
  NOR4X1  g11598(.A(n13405), .B(n11499), .C(n11404), .D(n13421), .Y(n13422));
  NAND4X1 g11599(.A(n11570), .B(n11609), .C(n11524), .D(n13422), .Y(n13423));
  NOR4X1  g11600(.A(n13402), .B(n13401), .C(n11739), .D(n13423), .Y(n13424));
  NAND3X1 g11601(.A(n13424), .B(n11822), .C(n11790), .Y(n13425));
  AOI21X1 g11602(.A0(n11916), .A1(n11911), .B0(n13425), .Y(n13426));
  NAND3X1 g11603(.A(n13426), .B(n11909), .C(n11965), .Y(n13427));
  NOR3X1  g11604(.A(n13427), .B(n13397), .C(n13396), .Y(n13428));
  XOR2X1  g11605(.A(n13428), .B(n10576), .Y(n13429));
  NAND2X1 g11606(.A(n10566), .B(n10560), .Y(n13430));
  INVX1   g11607(.A(n13430), .Y(n13431));
  NAND2X1 g11608(.A(n13431), .B(n13429), .Y(n13432));
  NAND4X1 g11609(.A(n13395), .B(n13391), .C(n13387), .D(n13432), .Y(n13433));
  NOR2X1  g11610(.A(n13433), .B(n13287), .Y(n13434));
  NAND2X1 g11611(.A(n13395), .B(n10445), .Y(n13435));
  NAND2X1 g11612(.A(n13395), .B(P3_U3151), .Y(n13436));
  OAI21X1 g11613(.A0(n13435), .A1(n13287), .B0(n13436), .Y(n13437));
  AOI21X1 g11614(.A0(n13434), .A1(n13285), .B0(n13437), .Y(P3_U3296));
  AOI21X1 g11615(.A0(n10576), .A1(n10560), .B0(n10566), .Y(n13439));
  INVX1   g11616(.A(n13439), .Y(n13440));
  OAI21X1 g11617(.A0(n13430), .A1(n12105), .B0(n13440), .Y(n13441));
  XOR2X1  g11618(.A(n13441), .B(n10705), .Y(n13442));
  XOR2X1  g11619(.A(n13441), .B(n10753), .Y(n13443));
  AOI22X1 g11620(.A0(n13442), .A1(n10691), .B0(n10761), .B1(n13443), .Y(n13444));
  AOI21X1 g11621(.A0(n13431), .A1(n10557), .B0(n13439), .Y(n13445));
  XOR2X1  g11622(.A(n13445), .B(n10667), .Y(n13446));
  AOI21X1 g11623(.A0(n13445), .A1(n10635), .B0(n10615), .Y(n13447));
  OAI21X1 g11624(.A0(n13446), .A1(n10662), .B0(n13447), .Y(n13448));
  XOR2X1  g11625(.A(n13441), .B(n10667), .Y(n13449));
  NAND2X1 g11626(.A(n13441), .B(n10635), .Y(n13450));
  AOI21X1 g11627(.A0(n13449), .A1(n10645), .B0(n13450), .Y(n13451));
  NOR2X1  g11628(.A(n13449), .B(n10645), .Y(n13452));
  NOR2X1  g11629(.A(n13452), .B(n13451), .Y(n13453));
  NAND2X1 g11630(.A(n13453), .B(n13448), .Y(n13454));
  NOR2X1  g11631(.A(n13442), .B(n10691), .Y(n13455));
  NAND2X1 g11632(.A(n13455), .B(n10738), .Y(n13456));
  INVX1   g11633(.A(n13443), .Y(n13457));
  OAI21X1 g11634(.A0(n13455), .A1(n10738), .B0(n13457), .Y(n13458));
  NAND2X1 g11635(.A(n13458), .B(n13456), .Y(n13459));
  AOI21X1 g11636(.A0(n13454), .A1(n13444), .B0(n13459), .Y(n13460));
  XOR2X1  g11637(.A(n13441), .B(n10803), .Y(n13461));
  NOR2X1  g11638(.A(n13461), .B(n10816), .Y(n13462));
  NOR2X1  g11639(.A(n13461), .B(n13460), .Y(n13463));
  NOR2X1  g11640(.A(n13463), .B(n13462), .Y(n13464));
  OAI21X1 g11641(.A0(n13460), .A1(n10816), .B0(n13464), .Y(n13465));
  XOR2X1  g11642(.A(n13445), .B(n11006), .Y(n13466));
  INVX1   g11643(.A(n13466), .Y(n13467));
  NOR2X1  g11644(.A(n13467), .B(n10996), .Y(n13468));
  INVX1   g11645(.A(n13468), .Y(n13469));
  XOR2X1  g11646(.A(n13445), .B(n10919), .Y(n13470));
  XOR2X1  g11647(.A(n13445), .B(n10962), .Y(n13471));
  AOI22X1 g11648(.A0(n13470), .A1(n10914), .B0(n10957), .B1(n13471), .Y(n13472));
  INVX1   g11649(.A(n13472), .Y(n13473));
  XOR2X1  g11650(.A(n13441), .B(n10861), .Y(n13474));
  AOI21X1 g11651(.A0(n13474), .A1(n10859), .B0(n13473), .Y(n13475));
  NAND2X1 g11652(.A(n13475), .B(n13469), .Y(n13476));
  INVX1   g11653(.A(n13476), .Y(n13477));
  INVX1   g11654(.A(n13471), .Y(n13478));
  NOR2X1  g11655(.A(n13470), .B(n10914), .Y(n13479));
  OAI21X1 g11656(.A0(n13479), .A1(n10946), .B0(n13478), .Y(n13480));
  NOR2X1  g11657(.A(n13474), .B(n10859), .Y(n13481));
  AOI22X1 g11658(.A0(n13479), .A1(n10946), .B0(n13472), .B1(n13481), .Y(n13482));
  NAND2X1 g11659(.A(n13482), .B(n13480), .Y(n13483));
  NOR2X1  g11660(.A(n13466), .B(n11061), .Y(n13484));
  AOI21X1 g11661(.A0(n13483), .A1(n13469), .B0(n13484), .Y(n13485));
  INVX1   g11662(.A(n13485), .Y(n13486));
  AOI21X1 g11663(.A0(n13477), .A1(n13465), .B0(n13486), .Y(n13487));
  NOR2X1  g11664(.A(n13487), .B(n11045), .Y(n13488));
  XOR2X1  g11665(.A(n13445), .B(n11050), .Y(n13489));
  AOI21X1 g11666(.A0(n13487), .A1(n11045), .B0(n13489), .Y(n13490));
  XOR2X1  g11667(.A(n13441), .B(n11302), .Y(n13491));
  INVX1   g11668(.A(n13491), .Y(n13492));
  NOR2X1  g11669(.A(n13492), .B(n11292), .Y(n13493));
  XOR2X1  g11670(.A(n13441), .B(n11202), .Y(n13494));
  XOR2X1  g11671(.A(n13445), .B(n11251), .Y(n13495));
  AOI22X1 g11672(.A0(n13494), .A1(n11207), .B0(n11266), .B1(n13495), .Y(n13496));
  INVX1   g11673(.A(n13496), .Y(n13497));
  XOR2X1  g11674(.A(n13445), .B(n11145), .Y(n13498));
  INVX1   g11675(.A(n13498), .Y(n13499));
  NOR2X1  g11676(.A(n13499), .B(n11131), .Y(n13500));
  XOR2X1  g11677(.A(n13445), .B(n11102), .Y(n13501));
  INVX1   g11678(.A(n13501), .Y(n13502));
  NOR2X1  g11679(.A(n13502), .B(n11086), .Y(n13503));
  NOR4X1  g11680(.A(n13500), .B(n13497), .C(n13493), .D(n13503), .Y(n13504));
  OAI21X1 g11681(.A0(n13490), .A1(n13488), .B0(n13504), .Y(n13505));
  NOR4X1  g11682(.A(n13500), .B(n13497), .C(n11095), .D(n13501), .Y(n13506));
  INVX1   g11683(.A(n13495), .Y(n13507));
  NOR2X1  g11684(.A(n13507), .B(n11239), .Y(n13508));
  NOR2X1  g11685(.A(n13498), .B(n11140), .Y(n13509));
  NAND2X1 g11686(.A(n13509), .B(n13496), .Y(n13510));
  NOR2X1  g11687(.A(n13494), .B(n11207), .Y(n13511));
  AOI21X1 g11688(.A0(n13507), .A1(n11239), .B0(n13511), .Y(n13512));
  AOI21X1 g11689(.A0(n13512), .A1(n13510), .B0(n13508), .Y(n13513));
  NOR2X1  g11690(.A(n13513), .B(n13506), .Y(n13514));
  NOR2X1  g11691(.A(n13514), .B(n13493), .Y(n13515));
  AOI21X1 g11692(.A0(n13492), .A1(n11292), .B0(n13515), .Y(n13516));
  NAND2X1 g11693(.A(n13516), .B(n13505), .Y(n13517));
  XOR2X1  g11694(.A(n13445), .B(n11342), .Y(n13518));
  XOR2X1  g11695(.A(n13518), .B(n11331), .Y(n13519));
  XOR2X1  g11696(.A(n13519), .B(n13517), .Y(n13520));
  NOR3X1  g11697(.A(n10557), .B(n10553), .C(n10550), .Y(n13521));
  INVX1   g11698(.A(n13521), .Y(n13522));
  NOR3X1  g11699(.A(n10579), .B(n10575), .C(n13522), .Y(n13523));
  NAND2X1 g11700(.A(n10564), .B(n10563), .Y(n13524));
  INVX1   g11701(.A(n13524), .Y(n13525));
  NOR3X1  g11702(.A(n10577), .B(n10566), .C(n10564), .Y(n13526));
  NOR4X1  g11703(.A(n13525), .B(n12033), .C(n10629), .D(n13526), .Y(n13527));
  NOR4X1  g11704(.A(n12105), .B(n10552), .C(n10550), .D(n13527), .Y(n13528));
  OAI21X1 g11705(.A0(n13528), .A1(n13523), .B0(n10528), .Y(n13529));
  NOR3X1  g11706(.A(n12105), .B(n10552), .C(n10550), .Y(n13530));
  INVX1   g11707(.A(n13530), .Y(n13531));
  NOR4X1  g11708(.A(n10454), .B(n10446), .C(P3_U3151), .D(n12120), .Y(n13532));
  NOR2X1  g11709(.A(n13527), .B(n13530), .Y(n13533));
  NOR3X1  g11710(.A(n10579), .B(n10575), .C(n13521), .Y(n13534));
  NOR2X1  g11711(.A(n10454), .B(n10446), .Y(n13535));
  NAND3X1 g11712(.A(n10576), .B(n10564), .C(n10562), .Y(n13536));
  NAND3X1 g11713(.A(n10566), .B(n10564), .C(n10562), .Y(n13537));
  NAND3X1 g11714(.A(n13537), .B(n13536), .C(n13535), .Y(n13538));
  NOR3X1  g11715(.A(n13538), .B(n13534), .C(n13533), .Y(n13539));
  INVX1   g11716(.A(n13539), .Y(n13540));
  AOI22X1 g11717(.A0(n13532), .A1(n13531), .B0(P3_STATE_REG_SCAN_IN), .B1(n13540), .Y(n13541));
  INVX1   g11718(.A(n13541), .Y(n13542));
  NOR2X1  g11719(.A(n10582), .B(n10529), .Y(n13543));
  NOR4X1  g11720(.A(n10557), .B(n10553), .C(n10550), .D(n10636), .Y(n13544));
  INVX1   g11721(.A(n13544), .Y(n13545));
  NOR2X1  g11722(.A(n13545), .B(n11377), .Y(n13546));
  NOR4X1  g11723(.A(n10557), .B(n10553), .C(n10550), .D(n10679), .Y(n13547));
  INVX1   g11724(.A(n13547), .Y(n13548));
  OAI22X1 g11725(.A0(n12223), .A1(n13521), .B0(n11344), .B1(n13548), .Y(n13549));
  OAI21X1 g11726(.A0(n13549), .A1(n13546), .B0(n13543), .Y(n13550));
  AOI22X1 g11727(.A0(n12103), .A1(n10528), .B0(n13530), .B1(n13532), .Y(n13551));
  AOI22X1 g11728(.A0(n11342), .A1(n13627), .B0(P3_REG3_REG_15__SCAN_IN), .B1(P3_U3151), .Y(n13553));
  NAND2X1 g11729(.A(n13553), .B(n13550), .Y(n13554));
  AOI21X1 g11730(.A0(n13542), .A1(n11329), .B0(n13554), .Y(n13555));
  OAI21X1 g11731(.A0(n13529), .A1(n13520), .B0(n13555), .Y(P3_U3181));
  XOR2X1  g11732(.A(n13445), .B(n11737), .Y(n13557));
  INVX1   g11733(.A(n13557), .Y(n13558));
  NOR2X1  g11734(.A(n13558), .B(n11730), .Y(n13559));
  INVX1   g11735(.A(n13559), .Y(n13560));
  XOR2X1  g11736(.A(n13441), .B(n11699), .Y(n13561));
  NOR2X1  g11737(.A(n13561), .B(n11736), .Y(n13562));
  INVX1   g11738(.A(n13562), .Y(n13563));
  NAND2X1 g11739(.A(n13561), .B(n11736), .Y(n13564));
  INVX1   g11740(.A(n13564), .Y(n13565));
  XOR2X1  g11741(.A(n13445), .B(n11646), .Y(n13566));
  NOR2X1  g11742(.A(n13566), .B(n11645), .Y(n13567));
  INVX1   g11743(.A(n13566), .Y(n13568));
  NOR2X1  g11744(.A(n13568), .B(n11639), .Y(n13569));
  INVX1   g11745(.A(n13569), .Y(n13570));
  XOR2X1  g11746(.A(n13445), .B(n11608), .Y(n13571));
  INVX1   g11747(.A(n13571), .Y(n13572));
  XOR2X1  g11748(.A(n13445), .B(n11523), .Y(n13573));
  XOR2X1  g11749(.A(n13445), .B(n11560), .Y(n13574));
  AOI22X1 g11750(.A0(n13571), .A1(n11607), .B0(n11562), .B1(n13574), .Y(n13575));
  INVX1   g11751(.A(n13575), .Y(n13576));
  NOR3X1  g11752(.A(n13576), .B(n13573), .C(n11521), .Y(n13577));
  NOR2X1  g11753(.A(n13574), .B(n11562), .Y(n13578));
  AOI21X1 g11754(.A0(n13572), .A1(n11601), .B0(n13578), .Y(n13579));
  INVX1   g11755(.A(n13579), .Y(n13580));
  OAI22X1 g11756(.A0(n13577), .A1(n13580), .B0(n13572), .B1(n11601), .Y(n13581));
  XOR2X1  g11757(.A(n13441), .B(n11483), .Y(n13582));
  NOR2X1  g11758(.A(n13582), .B(n11498), .Y(n13583));
  INVX1   g11759(.A(n13582), .Y(n13584));
  NOR2X1  g11760(.A(n13584), .B(n11473), .Y(n13585));
  INVX1   g11761(.A(n13585), .Y(n13586));
  XOR2X1  g11762(.A(n13445), .B(n11382), .Y(n13587));
  XOR2X1  g11763(.A(n13441), .B(n11435), .Y(n13588));
  AOI22X1 g11764(.A0(n13587), .A1(n11377), .B0(n11485), .B1(n13588), .Y(n13589));
  INVX1   g11765(.A(n13589), .Y(n13590));
  INVX1   g11766(.A(n13518), .Y(n13591));
  NOR2X1  g11767(.A(n13591), .B(n11331), .Y(n13592));
  AOI21X1 g11768(.A0(n13516), .A1(n13505), .B0(n13592), .Y(n13593));
  AOI21X1 g11769(.A0(n13591), .A1(n11331), .B0(n13593), .Y(n13594));
  NOR2X1  g11770(.A(n13587), .B(n11377), .Y(n13595));
  INVX1   g11771(.A(n13595), .Y(n13596));
  AOI21X1 g11772(.A0(n13596), .A1(n11485), .B0(n13588), .Y(n13597));
  AOI21X1 g11773(.A0(n13595), .A1(n11424), .B0(n13597), .Y(n13598));
  OAI21X1 g11774(.A0(n13594), .A1(n13590), .B0(n13598), .Y(n13599));
  AOI21X1 g11775(.A0(n13599), .A1(n13586), .B0(n13583), .Y(n13600));
  AOI21X1 g11776(.A0(n13573), .A1(n11521), .B0(n13576), .Y(n13601));
  INVX1   g11777(.A(n13601), .Y(n13602));
  OAI21X1 g11778(.A0(n13602), .A1(n13600), .B0(n13581), .Y(n13603));
  AOI21X1 g11779(.A0(n13603), .A1(n13570), .B0(n13567), .Y(n13604));
  OAI21X1 g11780(.A0(n13604), .A1(n13565), .B0(n13563), .Y(n13605));
  NAND2X1 g11781(.A(n13605), .B(n13560), .Y(n13606));
  XOR2X1  g11782(.A(n13441), .B(n11789), .Y(n13607));
  INVX1   g11783(.A(n13607), .Y(n13608));
  XOR2X1  g11784(.A(n13445), .B(n11821), .Y(n13609));
  INVX1   g11785(.A(n13609), .Y(n13610));
  OAI22X1 g11786(.A0(n13608), .A1(n11778), .B0(n11814), .B1(n13610), .Y(n13611));
  NOR2X1  g11787(.A(n13609), .B(n11820), .Y(n13612));
  NOR3X1  g11788(.A(n13612), .B(n13611), .C(n13606), .Y(n13613));
  XOR2X1  g11789(.A(n13609), .B(n11814), .Y(n13614));
  NOR2X1  g11790(.A(n13557), .B(n11731), .Y(n13615));
  AOI21X1 g11791(.A0(n13608), .A1(n11778), .B0(n13615), .Y(n13616));
  NAND3X1 g11792(.A(n13616), .B(n13614), .C(n13606), .Y(n13617));
  INVX1   g11793(.A(n13615), .Y(n13618));
  NOR3X1  g11794(.A(n13618), .B(n13612), .C(n13611), .Y(n13619));
  NOR2X1  g11795(.A(n13619), .B(n13529), .Y(n13620));
  NOR2X1  g11796(.A(n13608), .B(n11778), .Y(n13621));
  NAND2X1 g11797(.A(n13608), .B(n11778), .Y(n13622));
  NOR3X1  g11798(.A(n13622), .B(n13612), .C(n13611), .Y(n13623));
  AOI21X1 g11799(.A0(n13614), .A1(n13621), .B0(n13623), .Y(n13624));
  NAND3X1 g11800(.A(n13624), .B(n13620), .C(n13617), .Y(n13625));
  NAND4X1 g11801(.A(n10557), .B(n10553), .C(n10549), .D(n12393), .Y(n13626));
  AOI21X1 g11802(.A0(n13626), .A1(n12148), .B0(n10529), .Y(n13627));
  NOR2X1  g11803(.A(n11810), .B(n13521), .Y(n13630));
  AOI21X1 g11804(.A0(n13547), .A1(n11778), .B0(n13630), .Y(n13631));
  OAI21X1 g11805(.A0(n13545), .A1(n11910), .B0(n13631), .Y(n13632));
  AOI22X1 g11806(.A0(n13543), .A1(n13632), .B0(P3_REG3_REG_26__SCAN_IN), .B1(P3_U3151), .Y(n13633));
  OAI21X1 g11807(.A0(n13541), .A1(n11810), .B0(n13633), .Y(n13634));
  AOI21X1 g11808(.A0(n13627), .A1(n11821), .B0(n13634), .Y(n13635));
  OAI21X1 g11809(.A0(n13625), .A1(n13613), .B0(n13635), .Y(P3_U3180));
  XOR2X1  g11810(.A(n13470), .B(n10914), .Y(n13637));
  NAND2X1 g11811(.A(n13474), .B(n10859), .Y(n13638));
  AOI21X1 g11812(.A0(n13638), .A1(n13465), .B0(n13481), .Y(n13639));
  NOR2X1  g11813(.A(n13637), .B(n13639), .Y(n13641));
  AOI21X1 g11814(.A0(n13639), .A1(n13637), .B0(n13641), .Y(n13642));
  NOR2X1  g11815(.A(n13545), .B(n10957), .Y(n13643));
  OAI22X1 g11816(.A0(n10894), .A1(n13521), .B0(n10859), .B1(n13548), .Y(n13644));
  OAI21X1 g11817(.A0(n13644), .A1(n13643), .B0(n13543), .Y(n13645));
  AOI22X1 g11818(.A0(n10919), .A1(n13627), .B0(P3_REG3_REG_6__SCAN_IN), .B1(P3_U3151), .Y(n13646));
  NAND2X1 g11819(.A(n13646), .B(n13645), .Y(n13647));
  AOI21X1 g11820(.A0(n13542), .A1(n10895), .B0(n13647), .Y(n13648));
  OAI21X1 g11821(.A0(n13642), .A1(n13529), .B0(n13648), .Y(P3_U3179));
  XOR2X1  g11822(.A(n13582), .B(n11473), .Y(n13650));
  XOR2X1  g11823(.A(n13650), .B(n13599), .Y(n13651));
  INVX1   g11824(.A(n13543), .Y(n13652));
  OAI22X1 g11825(.A0(n11470), .A1(n13521), .B0(n11485), .B1(n13548), .Y(n13653));
  AOI21X1 g11826(.A0(n13544), .A1(n11515), .B0(n13653), .Y(n13654));
  AOI22X1 g11827(.A0(n11508), .A1(n13627), .B0(P3_REG3_REG_18__SCAN_IN), .B1(P3_U3151), .Y(n13655));
  OAI21X1 g11828(.A0(n13654), .A1(n13652), .B0(n13655), .Y(n13656));
  AOI21X1 g11829(.A0(n13542), .A1(n11471), .B0(n13656), .Y(n13657));
  OAI21X1 g11830(.A0(n13651), .A1(n13529), .B0(n13657), .Y(P3_U3178));
  INVX1   g11831(.A(n13529), .Y(n13659));
  XOR2X1  g11832(.A(n13442), .B(n10709), .Y(n13660));
  INVX1   g11833(.A(n13442), .Y(n13661));
  NOR2X1  g11834(.A(n13661), .B(n10709), .Y(n13662));
  OAI21X1 g11835(.A0(n13455), .A1(n13662), .B0(n13454), .Y(n13663));
  OAI21X1 g11836(.A0(n13660), .A1(n13454), .B0(n13663), .Y(n13664));
  NAND2X1 g11837(.A(n13664), .B(n13659), .Y(n13665));
  NAND2X1 g11838(.A(n13542), .B(P3_REG3_REG_2__SCAN_IN), .Y(n13666));
  AOI22X1 g11839(.A0(n10662), .A1(n13547), .B0(n13522), .B1(P3_REG3_REG_2__SCAN_IN), .Y(n13667));
  OAI21X1 g11840(.A0(n13545), .A1(n10761), .B0(n13667), .Y(n13668));
  OAI22X1 g11841(.A0(n10705), .A1(n13551), .B0(n10688), .B1(P3_STATE_REG_SCAN_IN), .Y(n13669));
  AOI21X1 g11842(.A0(n13668), .A1(n13543), .B0(n13669), .Y(n13670));
  NAND3X1 g11843(.A(n13670), .B(n13666), .C(n13665), .Y(P3_U3177));
  NOR2X1  g11844(.A(n13501), .B(n11095), .Y(n13672));
  NOR2X1  g11845(.A(n13490), .B(n13488), .Y(n13673));
  NOR2X1  g11846(.A(n13503), .B(n13673), .Y(n13674));
  NOR2X1  g11847(.A(n13674), .B(n13672), .Y(n13675));
  XOR2X1  g11848(.A(n13498), .B(n11140), .Y(n13676));
  INVX1   g11849(.A(n13500), .Y(n13677));
  INVX1   g11850(.A(n13509), .Y(n13678));
  AOI21X1 g11851(.A0(n13678), .A1(n13677), .B0(n13675), .Y(n13679));
  AOI21X1 g11852(.A0(n13676), .A1(n13675), .B0(n13679), .Y(n13680));
  NOR2X1  g11853(.A(n13545), .B(n11207), .Y(n13681));
  OAI22X1 g11854(.A0(n11128), .A1(n13521), .B0(n11095), .B1(n13548), .Y(n13682));
  OAI21X1 g11855(.A0(n13682), .A1(n13681), .B0(n13543), .Y(n13683));
  AOI22X1 g11856(.A0(n11145), .A1(n13627), .B0(P3_REG3_REG_11__SCAN_IN), .B1(P3_U3151), .Y(n13684));
  NAND2X1 g11857(.A(n13684), .B(n13683), .Y(n13685));
  AOI21X1 g11858(.A0(n13542), .A1(n12195), .B0(n13685), .Y(n13686));
  OAI21X1 g11859(.A0(n13680), .A1(n13529), .B0(n13686), .Y(P3_U3176));
  XOR2X1  g11860(.A(n13566), .B(n11639), .Y(n13688));
  XOR2X1  g11861(.A(n13688), .B(n13603), .Y(n13689));
  AOI22X1 g11862(.A0(n11637), .A1(n13522), .B0(n11601), .B1(n13547), .Y(n13690));
  OAI21X1 g11863(.A0(n13545), .A1(n11736), .B0(n13690), .Y(n13691));
  AOI22X1 g11864(.A0(n13543), .A1(n13691), .B0(P3_REG3_REG_22__SCAN_IN), .B1(P3_U3151), .Y(n13692));
  OAI21X1 g11865(.A0(n13541), .A1(n11636), .B0(n13692), .Y(n13693));
  AOI21X1 g11866(.A0(n13627), .A1(n11646), .B0(n13693), .Y(n13694));
  OAI21X1 g11867(.A0(n13689), .A1(n13529), .B0(n13694), .Y(P3_U3175));
  OAI21X1 g11868(.A0(n13674), .A1(n13672), .B0(n13677), .Y(n13696));
  NAND2X1 g11869(.A(n13696), .B(n13678), .Y(n13697));
  NOR2X1  g11870(.A(n13697), .B(n13511), .Y(n13698));
  OAI21X1 g11871(.A0(n13495), .A1(n11266), .B0(n13496), .Y(n13699));
  NOR2X1  g11872(.A(n13699), .B(n13698), .Y(n13700));
  AOI22X1 g11873(.A0(n13678), .A1(n13696), .B0(n13494), .B1(n11207), .Y(n13701));
  AOI21X1 g11874(.A0(n13507), .A1(n11266), .B0(n13511), .Y(n13702));
  OAI21X1 g11875(.A0(n13507), .A1(n11266), .B0(n13702), .Y(n13703));
  OAI21X1 g11876(.A0(n13703), .A1(n13701), .B0(n13659), .Y(n13704));
  INVX1   g11877(.A(n11237), .Y(n13705));
  OAI22X1 g11878(.A0(n13705), .A1(n13521), .B0(n11207), .B1(n13548), .Y(n13706));
  AOI21X1 g11879(.A0(n13544), .A1(n11292), .B0(n13706), .Y(n13707));
  AOI22X1 g11880(.A0(n11251), .A1(n13627), .B0(P3_REG3_REG_13__SCAN_IN), .B1(P3_U3151), .Y(n13708));
  OAI21X1 g11881(.A0(n13707), .A1(n13652), .B0(n13708), .Y(n13709));
  AOI21X1 g11882(.A0(n13542), .A1(n11237), .B0(n13709), .Y(n13710));
  OAI21X1 g11883(.A0(n13704), .A1(n13700), .B0(n13710), .Y(P3_U3174));
  XOR2X1  g11884(.A(n13574), .B(n11562), .Y(n13712));
  NOR2X1  g11885(.A(n13573), .B(n11521), .Y(n13713));
  AOI21X1 g11886(.A0(n13573), .A1(n11521), .B0(n13600), .Y(n13714));
  NOR2X1  g11887(.A(n13714), .B(n13713), .Y(n13715));
  NOR2X1  g11888(.A(n13712), .B(n13715), .Y(n13717));
  AOI21X1 g11889(.A0(n13715), .A1(n13712), .B0(n13717), .Y(n13718));
  AOI22X1 g11890(.A0(n11552), .A1(n13522), .B0(n11515), .B1(n13547), .Y(n13719));
  OAI21X1 g11891(.A0(n13545), .A1(n11607), .B0(n13719), .Y(n13720));
  AOI22X1 g11892(.A0(n13543), .A1(n13720), .B0(P3_REG3_REG_20__SCAN_IN), .B1(P3_U3151), .Y(n13721));
  OAI21X1 g11893(.A0(n13541), .A1(n11551), .B0(n13721), .Y(n13722));
  AOI21X1 g11894(.A0(n13627), .A1(n11560), .B0(n13722), .Y(n13723));
  OAI21X1 g11895(.A0(n13718), .A1(n13529), .B0(n13723), .Y(P3_U3173));
  AOI21X1 g11896(.A0(n13543), .A1(n13522), .B0(n13542), .Y(n13725));
  NOR3X1  g11897(.A(n10645), .B(n10582), .C(n10529), .Y(n13727));
  AOI22X1 g11898(.A0(n13544), .A1(n13727), .B0(P3_REG3_REG_0__SCAN_IN), .B1(P3_U3151), .Y(n13728));
  OAI21X1 g11899(.A0(n13551), .A1(n10635), .B0(n13728), .Y(n13729));
  AOI21X1 g11900(.A0(n13412), .A1(n13659), .B0(n13729), .Y(n13730));
  OAI21X1 g11901(.A0(n13725), .A1(n10608), .B0(n13730), .Y(P3_U3172));
  XOR2X1  g11902(.A(n13489), .B(n11045), .Y(n13732));
  XOR2X1  g11903(.A(n13732), .B(n13487), .Y(n13733));
  NOR2X1  g11904(.A(n13545), .B(n11095), .Y(n13734));
  OAI22X1 g11905(.A0(n11033), .A1(n13521), .B0(n11061), .B1(n13548), .Y(n13735));
  OAI21X1 g11906(.A0(n13735), .A1(n13734), .B0(n13543), .Y(n13736));
  AOI22X1 g11907(.A0(n11050), .A1(n13627), .B0(P3_REG3_REG_9__SCAN_IN), .B1(P3_U3151), .Y(n13737));
  NAND2X1 g11908(.A(n13737), .B(n13736), .Y(n13738));
  AOI21X1 g11909(.A0(n13542), .A1(n11032), .B0(n13738), .Y(n13739));
  OAI21X1 g11910(.A0(n13733), .A1(n13529), .B0(n13739), .Y(P3_U3171));
  XOR2X1  g11911(.A(n13461), .B(n10816), .Y(n13741));
  XOR2X1  g11912(.A(n13741), .B(n13460), .Y(n13742));
  OAI22X1 g11913(.A0(n10790), .A1(n13521), .B0(n10761), .B1(n13548), .Y(n13743));
  AOI21X1 g11914(.A0(n13544), .A1(n10844), .B0(n13743), .Y(n13744));
  AOI22X1 g11915(.A0(n10835), .A1(n13627), .B0(P3_REG3_REG_4__SCAN_IN), .B1(P3_U3151), .Y(n13745));
  OAI21X1 g11916(.A0(n13744), .A1(n13652), .B0(n13745), .Y(n13746));
  AOI21X1 g11917(.A0(n13542), .A1(n10791), .B0(n13746), .Y(n13747));
  OAI21X1 g11918(.A0(n13742), .A1(n13529), .B0(n13747), .Y(P3_U3170));
  NOR2X1  g11919(.A(n13604), .B(n13565), .Y(n13749));
  NOR2X1  g11920(.A(n13749), .B(n13562), .Y(n13750));
  XOR2X1  g11921(.A(n13557), .B(n11731), .Y(n13751));
  AOI21X1 g11922(.A0(n13618), .A1(n13560), .B0(n13750), .Y(n13752));
  AOI21X1 g11923(.A0(n13751), .A1(n13750), .B0(n13752), .Y(n13753));
  AOI22X1 g11924(.A0(n11728), .A1(n13522), .B0(n11691), .B1(n13547), .Y(n13754));
  OAI21X1 g11925(.A0(n13545), .A1(n11777), .B0(n13754), .Y(n13755));
  AOI22X1 g11926(.A0(n13543), .A1(n13755), .B0(P3_REG3_REG_24__SCAN_IN), .B1(P3_U3151), .Y(n13756));
  OAI21X1 g11927(.A0(n13541), .A1(n11727), .B0(n13756), .Y(n13757));
  AOI21X1 g11928(.A0(n13627), .A1(n11737), .B0(n13757), .Y(n13758));
  OAI21X1 g11929(.A0(n13753), .A1(n13529), .B0(n13758), .Y(P3_U3169));
  OAI21X1 g11930(.A0(n13588), .A1(n11485), .B0(n13589), .Y(n13760));
  AOI21X1 g11931(.A0(n13596), .A1(n13594), .B0(n13760), .Y(n13761));
  AOI21X1 g11932(.A0(n13587), .A1(n11377), .B0(n13594), .Y(n13762));
  INVX1   g11933(.A(n13588), .Y(n13763));
  AOI21X1 g11934(.A0(n13763), .A1(n11485), .B0(n13595), .Y(n13764));
  OAI21X1 g11935(.A0(n13763), .A1(n11485), .B0(n13764), .Y(n13765));
  OAI21X1 g11936(.A0(n13765), .A1(n13762), .B0(n13659), .Y(n13766));
  INVX1   g11937(.A(n11422), .Y(n13767));
  OAI22X1 g11938(.A0(n13767), .A1(n13521), .B0(n11377), .B1(n13548), .Y(n13768));
  AOI21X1 g11939(.A0(n13544), .A1(n11473), .B0(n13768), .Y(n13769));
  AOI22X1 g11940(.A0(n11436), .A1(n13627), .B0(P3_REG3_REG_17__SCAN_IN), .B1(P3_U3151), .Y(n13770));
  OAI21X1 g11941(.A0(n13769), .A1(n13652), .B0(n13770), .Y(n13771));
  AOI21X1 g11942(.A0(n13542), .A1(n11422), .B0(n13771), .Y(n13772));
  OAI21X1 g11943(.A0(n13766), .A1(n13761), .B0(n13772), .Y(P3_U3168));
  XOR2X1  g11944(.A(n13474), .B(n10844), .Y(n13774));
  XOR2X1  g11945(.A(n13774), .B(n13465), .Y(n13775));
  NOR2X1  g11946(.A(n13545), .B(n10914), .Y(n13776));
  OAI22X1 g11947(.A0(n10841), .A1(n13521), .B0(n10816), .B1(n13548), .Y(n13777));
  OAI21X1 g11948(.A0(n13777), .A1(n13776), .B0(n13543), .Y(n13778));
  AOI22X1 g11949(.A0(n10855), .A1(n13627), .B0(P3_REG3_REG_5__SCAN_IN), .B1(P3_U3151), .Y(n13779));
  NAND2X1 g11950(.A(n13779), .B(n13778), .Y(n13780));
  AOI21X1 g11951(.A0(n13542), .A1(n10842), .B0(n13780), .Y(n13781));
  OAI21X1 g11952(.A0(n13775), .A1(n13529), .B0(n13781), .Y(P3_U3167));
  XOR2X1  g11953(.A(n13587), .B(n11377), .Y(n13783));
  NOR2X1  g11954(.A(n13783), .B(n13594), .Y(n13785));
  AOI21X1 g11955(.A0(n13783), .A1(n13594), .B0(n13785), .Y(n13786));
  NOR2X1  g11956(.A(n13545), .B(n11485), .Y(n13787));
  OAI22X1 g11957(.A0(n11366), .A1(n13521), .B0(n11337), .B1(n13548), .Y(n13788));
  OAI21X1 g11958(.A0(n13788), .A1(n13787), .B0(n13543), .Y(n13789));
  AOI22X1 g11959(.A0(n11382), .A1(n13627), .B0(P3_REG3_REG_16__SCAN_IN), .B1(P3_U3151), .Y(n13790));
  NAND2X1 g11960(.A(n13790), .B(n13789), .Y(n13791));
  AOI21X1 g11961(.A0(n13542), .A1(n11367), .B0(n13791), .Y(n13792));
  OAI21X1 g11962(.A0(n13786), .A1(n13529), .B0(n13792), .Y(P3_U3166));
  AOI21X1 g11963(.A0(n13605), .A1(n13560), .B0(n13615), .Y(n13794));
  XOR2X1  g11964(.A(n13607), .B(n11777), .Y(n13795));
  NOR2X1  g11965(.A(n13795), .B(n13794), .Y(n13797));
  AOI21X1 g11966(.A0(n13795), .A1(n13794), .B0(n13797), .Y(n13798));
  AOI22X1 g11967(.A0(n12288), .A1(n13522), .B0(n11730), .B1(n13547), .Y(n13799));
  OAI21X1 g11968(.A0(n13545), .A1(n11820), .B0(n13799), .Y(n13800));
  AOI22X1 g11969(.A0(n13543), .A1(n13800), .B0(P3_REG3_REG_25__SCAN_IN), .B1(P3_U3151), .Y(n13801));
  OAI21X1 g11970(.A0(n13541), .A1(n11770), .B0(n13801), .Y(n13802));
  AOI21X1 g11971(.A0(n13627), .A1(n11808), .B0(n13802), .Y(n13803));
  OAI21X1 g11972(.A0(n13798), .A1(n13529), .B0(n13803), .Y(P3_U3165));
  XOR2X1  g11973(.A(n13494), .B(n11191), .Y(n13805));
  NOR2X1  g11974(.A(n13805), .B(n13697), .Y(n13806));
  AOI21X1 g11975(.A0(n13805), .A1(n13697), .B0(n13806), .Y(n13808));
  NOR2X1  g11976(.A(n13545), .B(n11266), .Y(n13809));
  OAI22X1 g11977(.A0(n11188), .A1(n13521), .B0(n11140), .B1(n13548), .Y(n13810));
  OAI21X1 g11978(.A0(n13810), .A1(n13809), .B0(n13543), .Y(n13811));
  AOI22X1 g11979(.A0(n11232), .A1(n13627), .B0(P3_REG3_REG_12__SCAN_IN), .B1(P3_U3151), .Y(n13812));
  NAND2X1 g11980(.A(n13812), .B(n13811), .Y(n13813));
  AOI21X1 g11981(.A0(n13542), .A1(n11189), .B0(n13813), .Y(n13814));
  OAI21X1 g11982(.A0(n13808), .A1(n13529), .B0(n13814), .Y(P3_U3164));
  NOR3X1  g11983(.A(n13714), .B(n13578), .C(n13713), .Y(n13816));
  OAI21X1 g11984(.A0(n13571), .A1(n11607), .B0(n13575), .Y(n13817));
  NOR2X1  g11985(.A(n13817), .B(n13816), .Y(n13818));
  AOI21X1 g11986(.A0(n13574), .A1(n11562), .B0(n13715), .Y(n13819));
  AOI21X1 g11987(.A0(n13572), .A1(n11607), .B0(n13578), .Y(n13820));
  OAI21X1 g11988(.A0(n13572), .A1(n11607), .B0(n13820), .Y(n13821));
  OAI21X1 g11989(.A0(n13821), .A1(n13819), .B0(n13659), .Y(n13822));
  AOI22X1 g11990(.A0(n11599), .A1(n13522), .B0(n11554), .B1(n13547), .Y(n13823));
  OAI21X1 g11991(.A0(n13545), .A1(n11645), .B0(n13823), .Y(n13824));
  AOI22X1 g11992(.A0(n13543), .A1(n13824), .B0(P3_REG3_REG_21__SCAN_IN), .B1(P3_U3151), .Y(n13825));
  OAI21X1 g11993(.A0(n13541), .A1(n12260), .B0(n13825), .Y(n13826));
  AOI21X1 g11994(.A0(n13627), .A1(n11608), .B0(n13826), .Y(n13827));
  OAI21X1 g11995(.A0(n13822), .A1(n13818), .B0(n13827), .Y(P3_U3163));
  AOI21X1 g11996(.A0(n13441), .A1(n10635), .B0(n13447), .Y(n13829));
  XOR2X1  g11997(.A(n13446), .B(n10645), .Y(n13830));
  XOR2X1  g11998(.A(n13830), .B(n13829), .Y(n13831));
  NOR2X1  g11999(.A(n13545), .B(n10691), .Y(n13832));
  OAI22X1 g12000(.A0(n10615), .A1(n13548), .B0(n13521), .B1(n10642), .Y(n13833));
  OAI21X1 g12001(.A0(n13833), .A1(n13832), .B0(n13543), .Y(n13834));
  AOI22X1 g12002(.A0(n10720), .A1(n13627), .B0(P3_REG3_REG_1__SCAN_IN), .B1(P3_U3151), .Y(n13835));
  NAND2X1 g12003(.A(n13835), .B(n13834), .Y(n13836));
  AOI21X1 g12004(.A0(n13831), .A1(n13659), .B0(n13836), .Y(n13837));
  OAI21X1 g12005(.A0(n13541), .A1(n10642), .B0(n13837), .Y(P3_U3162));
  AOI21X1 g12006(.A0(n13475), .A1(n13465), .B0(n13483), .Y(n13839));
  XOR2X1  g12007(.A(n13466), .B(n11061), .Y(n13840));
  XOR2X1  g12008(.A(n13840), .B(n13839), .Y(n13841));
  NOR2X1  g12009(.A(n13545), .B(n11045), .Y(n13842));
  OAI22X1 g12010(.A0(n10993), .A1(n13521), .B0(n10957), .B1(n13548), .Y(n13843));
  OAI21X1 g12011(.A0(n13843), .A1(n13842), .B0(n13543), .Y(n13844));
  AOI22X1 g12012(.A0(n11006), .A1(n13627), .B0(P3_REG3_REG_8__SCAN_IN), .B1(P3_U3151), .Y(n13845));
  NAND2X1 g12013(.A(n13845), .B(n13844), .Y(n13846));
  AOI21X1 g12014(.A0(n13542), .A1(n10994), .B0(n13846), .Y(n13847));
  OAI21X1 g12015(.A0(n13841), .A1(n13529), .B0(n13847), .Y(P3_U3161));
  XOR2X1  g12016(.A(n13445), .B(n11869), .Y(n13849));
  NOR2X1  g12017(.A(n13849), .B(n11863), .Y(n13850));
  AOI21X1 g12018(.A0(n13607), .A1(n11777), .B0(n11820), .Y(n13851));
  AOI22X1 g12019(.A0(n13557), .A1(n11731), .B0(n11777), .B1(n13607), .Y(n13852));
  AOI22X1 g12020(.A0(n13610), .A1(n13852), .B0(n13851), .B1(n13560), .Y(n13853));
  NOR3X1  g12021(.A(n13853), .B(n13850), .C(n13750), .Y(n13854));
  INVX1   g12022(.A(n13612), .Y(n13855));
  OAI21X1 g12023(.A0(n13609), .A1(n11820), .B0(n13616), .Y(n13856));
  OAI21X1 g12024(.A0(n13849), .A1(n11863), .B0(n13856), .Y(n13857));
  AOI21X1 g12025(.A0(n13855), .A1(n13611), .B0(n13857), .Y(n13858));
  INVX1   g12026(.A(n13849), .Y(n13859));
  XOR2X1  g12027(.A(n13445), .B(n11902), .Y(n13860));
  XOR2X1  g12028(.A(n13860), .B(n11941), .Y(n13861));
  INVX1   g12029(.A(n13861), .Y(n13862));
  OAI21X1 g12030(.A0(n13859), .A1(n11910), .B0(n13862), .Y(n13863));
  NOR3X1  g12031(.A(n13863), .B(n13858), .C(n13854), .Y(n13864));
  OAI21X1 g12032(.A0(n13616), .A1(n13611), .B0(n13855), .Y(n13865));
  AOI21X1 g12033(.A0(n13849), .A1(n11863), .B0(n13865), .Y(n13866));
  OAI21X1 g12034(.A0(n13853), .A1(n13750), .B0(n13866), .Y(n13867));
  NOR2X1  g12035(.A(n13862), .B(n13850), .Y(n13868));
  AOI21X1 g12036(.A0(n13868), .A1(n13867), .B0(n13864), .Y(n13869));
  NOR2X1  g12037(.A(n11898), .B(n13521), .Y(n13870));
  AOI21X1 g12038(.A0(n13547), .A1(n11863), .B0(n13870), .Y(n13871));
  OAI21X1 g12039(.A0(n13545), .A1(n11949), .B0(n13871), .Y(n13872));
  AOI22X1 g12040(.A0(n13543), .A1(n13872), .B0(P3_REG3_REG_28__SCAN_IN), .B1(P3_U3151), .Y(n13873));
  OAI21X1 g12041(.A0(n13541), .A1(n11898), .B0(n13873), .Y(n13874));
  AOI21X1 g12042(.A0(n13627), .A1(n11941), .B0(n13874), .Y(n13875));
  OAI21X1 g12043(.A0(n13869), .A1(n13529), .B0(n13875), .Y(P3_U3160));
  XOR2X1  g12044(.A(n13573), .B(n11521), .Y(n13877));
  NOR2X1  g12045(.A(n13877), .B(n13600), .Y(n13879));
  AOI21X1 g12046(.A0(n13877), .A1(n13600), .B0(n13879), .Y(n13880));
  NAND2X1 g12047(.A(n13544), .B(n11554), .Y(n13881));
  AOI22X1 g12048(.A0(n11513), .A1(n13522), .B0(n11473), .B1(n13547), .Y(n13882));
  AOI21X1 g12049(.A0(n13882), .A1(n13881), .B0(n13652), .Y(n13883));
  AOI21X1 g12050(.A0(P3_REG3_REG_19__SCAN_IN), .A1(P3_U3151), .B0(n13883), .Y(n13884));
  OAI21X1 g12051(.A0(n13551), .A1(n11585), .B0(n13884), .Y(n13885));
  AOI21X1 g12052(.A0(n13542), .A1(n11513), .B0(n13885), .Y(n13886));
  OAI21X1 g12053(.A0(n13880), .A1(n13529), .B0(n13886), .Y(P3_U3159));
  NOR2X1  g12054(.A(n13455), .B(n13454), .Y(n13888));
  OAI21X1 g12055(.A0(n13443), .A1(n10761), .B0(n13444), .Y(n13889));
  OAI21X1 g12056(.A0(n13661), .A1(n10709), .B0(n13454), .Y(n13890));
  OAI22X1 g12057(.A0(n13442), .A1(n10691), .B0(n10738), .B1(n13443), .Y(n13891));
  AOI21X1 g12058(.A0(n13443), .A1(n10738), .B0(n13891), .Y(n13892));
  AOI21X1 g12059(.A0(n13892), .A1(n13890), .B0(n13529), .Y(n13893));
  OAI21X1 g12060(.A0(n13889), .A1(n13888), .B0(n13893), .Y(n13894));
  NAND2X1 g12061(.A(n13542), .B(n10736), .Y(n13895));
  AOI22X1 g12062(.A0(n10709), .A1(n13547), .B0(n13522), .B1(n10736), .Y(n13896));
  OAI21X1 g12063(.A0(n13545), .A1(n10816), .B0(n13896), .Y(n13897));
  OAI22X1 g12064(.A0(n10753), .A1(n13551), .B0(n10736), .B1(P3_STATE_REG_SCAN_IN), .Y(n13898));
  AOI21X1 g12065(.A0(n13897), .A1(n13543), .B0(n13898), .Y(n13899));
  NAND3X1 g12066(.A(n13899), .B(n13895), .C(n13894), .Y(P3_U3158));
  XOR2X1  g12067(.A(n13501), .B(n11095), .Y(n13901));
  XOR2X1  g12068(.A(n13901), .B(n13673), .Y(n13902));
  NOR2X1  g12069(.A(n13545), .B(n11140), .Y(n13903));
  OAI22X1 g12070(.A0(n11083), .A1(n13521), .B0(n11045), .B1(n13548), .Y(n13904));
  OAI21X1 g12071(.A0(n13904), .A1(n13903), .B0(n13543), .Y(n13905));
  AOI22X1 g12072(.A0(n11102), .A1(n13627), .B0(P3_REG3_REG_10__SCAN_IN), .B1(P3_U3151), .Y(n13906));
  NAND2X1 g12073(.A(n13906), .B(n13905), .Y(n13907));
  AOI21X1 g12074(.A0(n13542), .A1(n11084), .B0(n13907), .Y(n13908));
  OAI21X1 g12075(.A0(n13902), .A1(n13529), .B0(n13908), .Y(P3_U3157));
  XOR2X1  g12076(.A(n13561), .B(n11736), .Y(n13910));
  XOR2X1  g12077(.A(n13910), .B(n13604), .Y(n13911));
  NOR2X1  g12078(.A(n12274), .B(n13521), .Y(n13912));
  AOI21X1 g12079(.A0(n13547), .A1(n11639), .B0(n13912), .Y(n13913));
  OAI21X1 g12080(.A0(n13545), .A1(n11731), .B0(n13913), .Y(n13914));
  AOI22X1 g12081(.A0(n13543), .A1(n13914), .B0(P3_REG3_REG_23__SCAN_IN), .B1(P3_U3151), .Y(n13915));
  OAI21X1 g12082(.A0(n13541), .A1(n12274), .B0(n13915), .Y(n13916));
  AOI21X1 g12083(.A0(n13627), .A1(n13212), .B0(n13916), .Y(n13917));
  OAI21X1 g12084(.A0(n13911), .A1(n13529), .B0(n13917), .Y(P3_U3156));
  NOR3X1  g12085(.A(n13503), .B(n13500), .C(n13497), .Y(n13919));
  OAI21X1 g12086(.A0(n13490), .A1(n13488), .B0(n13919), .Y(n13920));
  NAND2X1 g12087(.A(n13920), .B(n13514), .Y(n13921));
  XOR2X1  g12088(.A(n13491), .B(n11292), .Y(n13922));
  XOR2X1  g12089(.A(n13922), .B(n13921), .Y(n13923));
  NOR2X1  g12090(.A(n13545), .B(n11337), .Y(n13924));
  OAI22X1 g12091(.A0(n11289), .A1(n13521), .B0(n11266), .B1(n13548), .Y(n13925));
  OAI21X1 g12092(.A0(n13925), .A1(n13924), .B0(n13543), .Y(n13926));
  AOI22X1 g12093(.A0(n11323), .A1(n13627), .B0(P3_REG3_REG_14__SCAN_IN), .B1(P3_U3151), .Y(n13927));
  NAND2X1 g12094(.A(n13927), .B(n13926), .Y(n13928));
  AOI21X1 g12095(.A0(n13542), .A1(n11290), .B0(n13928), .Y(n13929));
  OAI21X1 g12096(.A0(n13923), .A1(n13529), .B0(n13929), .Y(P3_U3155));
  INVX1   g12097(.A(n13853), .Y(n13931));
  AOI21X1 g12098(.A0(n13931), .A1(n13605), .B0(n13865), .Y(n13932));
  XOR2X1  g12099(.A(n13849), .B(n11863), .Y(n13933));
  XOR2X1  g12100(.A(n13933), .B(n13932), .Y(n13934));
  AOI22X1 g12101(.A0(n11858), .A1(n13522), .B0(n11814), .B1(n13547), .Y(n13935));
  OAI21X1 g12102(.A0(n13545), .A1(n11903), .B0(n13935), .Y(n13936));
  AOI22X1 g12103(.A0(n13543), .A1(n13936), .B0(P3_REG3_REG_27__SCAN_IN), .B1(P3_U3151), .Y(n13937));
  OAI21X1 g12104(.A0(n13541), .A1(n11859), .B0(n13937), .Y(n13938));
  AOI21X1 g12105(.A0(n13627), .A1(n11915), .B0(n13938), .Y(n13939));
  OAI21X1 g12106(.A0(n13934), .A1(n13529), .B0(n13939), .Y(P3_U3154));
  INVX1   g12107(.A(n13479), .Y(n13941));
  OAI21X1 g12108(.A0(n13471), .A1(n10957), .B0(n13472), .Y(n13942));
  AOI21X1 g12109(.A0(n13639), .A1(n13941), .B0(n13942), .Y(n13943));
  AOI21X1 g12110(.A0(n13470), .A1(n10914), .B0(n13639), .Y(n13944));
  AOI21X1 g12111(.A0(n13478), .A1(n10957), .B0(n13479), .Y(n13945));
  OAI21X1 g12112(.A0(n13478), .A1(n10957), .B0(n13945), .Y(n13946));
  OAI21X1 g12113(.A0(n13946), .A1(n13944), .B0(n13659), .Y(n13947));
  NOR2X1  g12114(.A(n13545), .B(n11061), .Y(n13948));
  OAI22X1 g12115(.A0(n10943), .A1(n13521), .B0(n10914), .B1(n13548), .Y(n13949));
  OAI21X1 g12116(.A0(n13949), .A1(n13948), .B0(n13543), .Y(n13950));
  AOI22X1 g12117(.A0(n10962), .A1(n13627), .B0(P3_REG3_REG_7__SCAN_IN), .B1(P3_U3151), .Y(n13951));
  NAND2X1 g12118(.A(n13951), .B(n13950), .Y(n13952));
  AOI21X1 g12119(.A0(n13542), .A1(n10944), .B0(n13952), .Y(n13953));
  OAI21X1 g12120(.A0(n13947), .A1(n13943), .B0(n13953), .Y(P3_U3153));
  INVX1   g12121(.A(n13535), .Y(n13955));
  AOI21X1 g12122(.A0(n11247), .A1(n10446), .B0(P3_U3151), .Y(n13956));
  OAI21X1 g12123(.A0(n12331), .A1(n13955), .B0(n13956), .Y(P3_U3150));
endmodule


