//Converted to Combinational (Partial output: n6131) , Module name: s38417_n6131 , Timestamp: 2018-12-03T15:51:14.374125 
module s38417_n6131 ( g2116, g1905, g1918, g2006, g2039, g2108, g2110, g2112, g2109, g2009, g2003, g2040, g2020, g2013, g2111, g2113, g2072, g2033, g2052, g2046, g2066, g2059, g2026, g2106, g2105, g2107, g2085, g2084, g2086, g2094, g2093, g2095, g2097, g2096, g2098, g2103, g2102, g2104, g2100, g2099, g2101, g2088, g2087, g2089, g2091, g2090, g2092, g2079, g2078, g2080, g2082, g2081, g2083, n6131 );
input g2116, g1905, g1918, g2006, g2039, g2108, g2110, g2112, g2109, g2009, g2003, g2040, g2020, g2013, g2111, g2113, g2072, g2033, g2052, g2046, g2066, g2059, g2026, g2106, g2105, g2107, g2085, g2084, g2086, g2094, g2093, g2095, g2097, g2096, g2098, g2103, g2102, g2104, g2100, g2099, g2101, g2088, g2087, g2089, g2091, g2090, g2092, g2079, g2078, g2080, g2082, g2081, g2083;
output n6131;
wire n8254, n8347, n8210, n8346, n8340, n8344, n8345, n8213, n8296, n8339, n8312, n8321, n8330, n8343, n8294, n8334, n8338, n8311, n8299, n8303, n8307, n8316, n8320, n8325, n8329, n8342, n8341, n8282, n8333, n8221_1, n8337, n8234, n8310, n8237, n8298, n8245, n8302, n8241, n8306, n8225, n8315, n8319, n8324, n8328, n8331, n8332, n8335, n8336, n8308, n8309, n8295, n8297, n8300, n8301, n8304, n8305, n8313, n8314, n8317, n8318, n8322, n8323, n8326, n8327;
MX2X1    g3304(.A(n8347), .B(g2116), .S0(n8254), .Y(n6131));
NAND4X1  g3209(.A(g2006), .B(g1918), .C(g1905), .D(n8210), .Y(n8254));
NOR4X1   g3302(.A(n8345), .B(n8344), .C(n8340), .D(n8346), .Y(n8347));
INVX1    g3165(.A(g2039), .Y(n8210));
OAI22X1  g3301(.A0(g2110), .A1(n8296), .B0(n8213), .B1(g2108), .Y(n8346));
NOR4X1   g3295(.A(n8330), .B(n8321), .C(n8312), .D(n8339), .Y(n8340));
OAI21X1  g3299(.A0(g2112), .A1(n8294), .B0(n8343), .Y(n8344));
NOR2X1   g3300(.A(g2109), .B(n8294), .Y(n8345));
INVX1    g3168(.A(g2009), .Y(n8213));
INVX1    g3251(.A(g2006), .Y(n8296));
OR2X1    g3294(.A(n8338), .B(n8334), .Y(n8339));
OR4X1    g3267(.A(n8307), .B(n8303), .C(n8299), .D(n8311), .Y(n8312));
NAND2X1  g3276(.A(n8320), .B(n8316), .Y(n8321));
NAND2X1  g3285(.A(n8329), .B(n8325), .Y(n8330));
AOI22X1  g3298(.A0(n8341), .A1(g2006), .B0(g2009), .B1(n8342), .Y(n8343));
INVX1    g3249(.A(g2003), .Y(n8294));
XOR2X1   g3289(.A(n8333), .B(n8282), .Y(n8334));
XOR2X1   g3293(.A(n8337), .B(n8221_1), .Y(n8338));
XOR2X1   g3266(.A(n8310), .B(n8234), .Y(n8311));
XOR2X1   g3254(.A(n8298), .B(n8237), .Y(n8299));
XOR2X1   g3258(.A(n8302), .B(n8245), .Y(n8303));
XOR2X1   g3262(.A(n8306), .B(n8241), .Y(n8307));
XOR2X1   g3271(.A(n8315), .B(n8225), .Y(n8316));
XOR2X1   g3275(.A(n8319), .B(g2040), .Y(n8320));
XOR2X1   g3280(.A(n8324), .B(g2020), .Y(n8325));
XOR2X1   g3284(.A(n8328), .B(g2013), .Y(n8329));
INVX1    g3297(.A(g2111), .Y(n8342));
INVX1    g3296(.A(g2113), .Y(n8341));
INVX1    g3237(.A(g2072), .Y(n8282));
NOR2X1   g3288(.A(n8332), .B(n8331), .Y(n8333));
INVX1    g3176(.A(g2033), .Y(n8221_1));
NOR2X1   g3292(.A(n8336), .B(n8335), .Y(n8337));
INVX1    g3189(.A(g2052), .Y(n8234));
NOR2X1   g3265(.A(n8309), .B(n8308), .Y(n8310));
INVX1    g3192(.A(g2046), .Y(n8237));
NOR2X1   g3253(.A(n8297), .B(n8295), .Y(n8298));
INVX1    g3200(.A(g2066), .Y(n8245));
NOR2X1   g3257(.A(n8301), .B(n8300), .Y(n8302));
INVX1    g3196(.A(g2059), .Y(n8241));
NOR2X1   g3261(.A(n8305), .B(n8304), .Y(n8306));
INVX1    g3180(.A(g2026), .Y(n8225));
OR2X1    g3270(.A(n8314), .B(n8313), .Y(n8315));
NOR2X1   g3274(.A(n8318), .B(n8317), .Y(n8319));
NOR2X1   g3279(.A(n8323), .B(n8322), .Y(n8324));
NOR2X1   g3283(.A(n8327), .B(n8326), .Y(n8328));
NOR2X1   g3286(.A(g2106), .B(n8294), .Y(n8331));
OAI22X1  g3287(.A0(g2107), .A1(n8296), .B0(n8213), .B1(g2105), .Y(n8332));
NOR2X1   g3290(.A(g2085), .B(n8294), .Y(n8335));
OAI22X1  g3291(.A0(g2086), .A1(n8296), .B0(n8213), .B1(g2084), .Y(n8336));
NOR2X1   g3263(.A(g2094), .B(n8294), .Y(n8308));
OAI22X1  g3264(.A0(g2095), .A1(n8296), .B0(n8213), .B1(g2093), .Y(n8309));
NOR2X1   g3250(.A(g2097), .B(n8294), .Y(n8295));
OAI22X1  g3252(.A0(g2098), .A1(n8296), .B0(n8213), .B1(g2096), .Y(n8297));
NOR2X1   g3255(.A(g2103), .B(n8294), .Y(n8300));
OAI22X1  g3256(.A0(g2104), .A1(n8296), .B0(n8213), .B1(g2102), .Y(n8301));
NOR2X1   g3259(.A(g2100), .B(n8294), .Y(n8304));
OAI22X1  g3260(.A0(g2101), .A1(n8296), .B0(n8213), .B1(g2099), .Y(n8305));
NOR2X1   g3268(.A(g2088), .B(n8294), .Y(n8313));
OAI22X1  g3269(.A0(g2089), .A1(n8296), .B0(n8213), .B1(g2087), .Y(n8314));
NOR2X1   g3272(.A(g2091), .B(n8294), .Y(n8317));
OAI22X1  g3273(.A0(g2092), .A1(n8296), .B0(n8213), .B1(g2090), .Y(n8318));
NOR2X1   g3277(.A(g2079), .B(n8294), .Y(n8322));
OAI22X1  g3278(.A0(g2080), .A1(n8296), .B0(n8213), .B1(g2078), .Y(n8323));
NOR2X1   g3281(.A(g2082), .B(n8294), .Y(n8326));
OAI22X1  g3282(.A0(g2083), .A1(n8296), .B0(n8213), .B1(g2081), .Y(n8327));

endmodule
