// Benchmark "b21_C" written by ABC on Wed Aug 05 14:44:42 2020

module b21_C ( 
    P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
    SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_, SI_17_,
    SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_, SI_8_,
    SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
    P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
    P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
    P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
    P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
    P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
    P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
    P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
    P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
    P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
    P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN,
    P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN,
    P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN,
    P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN,
    P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN,
    P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
    P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
    P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
    P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
    P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
    P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
    P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
    P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
    P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
    P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
    P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
    P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
    P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
    P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
    P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
    P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
    P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
    P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
    P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
    P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
    P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
    P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
    P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
    P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
    P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
    P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
    P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
    P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
    P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
    P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
    P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
    P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
    P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
    P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
    P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
    P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
    P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
    P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
    P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
    P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
    P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
    P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
    P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
    P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
    P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
    P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
    P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
    P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
    P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
    P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
    P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
    P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
    P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
    P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
    P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
    P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
    P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
    P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
    P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
    P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
    P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
    P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
    P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
    P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
    P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
    P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
    P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
    P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
    P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
    P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
    P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
    P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
    P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
    P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
    P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
    P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
    P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
    P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
    P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
    P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
    P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
    P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
    P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
    P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
    P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
    P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
    P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
    P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
    P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
    P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
    P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
    P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
    P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
    P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
    P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
    P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
    P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
    P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
    P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
    P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
    P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
    P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
    P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
    P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
    P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
    P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
    P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
    P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
    P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
    P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
    P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
    P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
    P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
    P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
    P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
    P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
    P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
    P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
    P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
    P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
    P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
    P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
    P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
    P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
    P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
    P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
    P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
    P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
    P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
    P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
    P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
    P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
    P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
    P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
    P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
    P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
    P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
    P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
    P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
    P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
    P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
    P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
    P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
    P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
    P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
    P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
    P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
    P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
    P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
    P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
    P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
    P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
    P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
    P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
    P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
    P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
    P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
    P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
    P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
    P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
    P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
    P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
    P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
    P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
    P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
    P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
    P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
    P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
    P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
    P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
    P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
    P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
    P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
    P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
    P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
    P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
    P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
    P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
    P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
    P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
    P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
    P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
    P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
    P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
    P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
    P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
    P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
    P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
    P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
    P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
    P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
    P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
    P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
    P2_DATAO_REG_5__SCAN_IN,
    ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
    ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
    ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
    ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
    U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348,
    P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341,
    P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334,
    P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327,
    P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440, P1_U3441,
    P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315,
    P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308,
    P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301,
    P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294,
    P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463, P1_U3466,
    P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484, P1_U3487,
    P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505, P1_U3508,
    P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516,
    P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523,
    P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530,
    P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537,
    P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544,
    P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551,
    P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289, P1_U3288,
    P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281,
    P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274,
    P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267,
    P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262, P1_U3261,
    P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254,
    P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247,
    P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241, P1_U3555,
    P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562,
    P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569,
    P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576,
    P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583,
    P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238, P1_U3237,
    P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230,
    P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223,
    P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216,
    P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084, P1_U3083,
    P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354, P2_U3353,
    P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347, P2_U3346,
    P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340, P2_U3339,
    P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333, P2_U3332,
    P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437, P2_U3438,
    P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320,
    P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313,
    P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306,
    P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299,
    P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
    P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
    P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502, P2_U3505,
    P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
    P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
    P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
    P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533, P2_U3534,
    P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541,
    P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548,
    P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294, P2_U3293,
    P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286,
    P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279,
    P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272,
    P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265,
    P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
    P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
    P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3552,
    P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
    P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565, P2_U3566,
    P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573,
    P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580,
    P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
    P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
    P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
    P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
    P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152, P2_U3151,
    P2_U3966  );
  input  P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_,
    SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
    SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
    SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
    P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
    P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
    P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
    P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
    P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
    P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
    P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
    P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
    P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
    P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN,
    P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN,
    P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN,
    P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN,
    P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN,
    P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
    P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
    P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
    P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
    P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
    P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
    P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
    P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
    P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
    P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
    P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
    P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
    P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
    P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
    P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
    P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
    P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
    P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
    P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
    P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
    P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
    P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
    P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
    P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
    P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
    P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
    P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
    P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
    P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
    P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
    P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
    P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
    P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
    P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
    P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
    P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
    P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
    P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
    P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
    P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
    P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
    P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
    P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
    P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
    P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
    P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
    P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
    P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
    P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
    P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
    P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
    P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
    P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
    P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
    P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
    P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
    P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
    P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
    P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
    P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
    P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
    P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
    P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
    P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
    P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
    P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
    P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
    P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
    P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
    P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
    P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
    P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
    P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
    P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
    P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
    P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
    P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
    P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
    P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
    P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
    P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
    P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
    P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
    P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
    P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
    P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
    P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
    P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
    P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
    P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
    P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
    P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
    P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
    P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
    P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
    P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
    P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
    P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
    P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
    P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
    P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
    P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
    P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
    P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
    P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
    P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
    P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
    P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
    P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
    P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
    P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
    P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
    P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
    P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
    P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
    P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
    P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
    P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
    P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
    P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
    P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
    P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
    P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
    P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
    P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
    P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
    P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
    P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
    P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
    P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
    P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
    P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
    P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
    P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
    P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
    P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
    P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
    P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
    P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
    P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
    P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
    P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
    P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
    P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
    P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
    P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
    P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
    P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
    P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
    P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
    P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
    P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
    P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
    P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
    P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
    P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
    P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
    P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
    P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
    P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
    P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
    P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
    P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
    P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
    P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
    P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
    P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
    P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
    P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
    P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
    P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
    P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
    P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
    P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
    P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
    P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
    P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
    P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
    P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
    P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
    P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
    P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
    P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
    P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
    P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
    P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
    P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
    P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
    P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
    P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
    P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
    P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
    P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
    P2_DATAO_REG_5__SCAN_IN;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
    ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
    ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
    ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
    U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348,
    P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341,
    P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334,
    P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327,
    P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440, P1_U3441,
    P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315,
    P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308,
    P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301,
    P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294,
    P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463, P1_U3466,
    P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484, P1_U3487,
    P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505, P1_U3508,
    P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515, P1_U3516,
    P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523,
    P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530,
    P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537,
    P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544,
    P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551,
    P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289, P1_U3288,
    P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281,
    P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274,
    P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267,
    P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262, P1_U3261,
    P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254,
    P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247,
    P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241, P1_U3555,
    P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561, P1_U3562,
    P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569,
    P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576,
    P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583,
    P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238, P1_U3237,
    P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230,
    P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223,
    P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216,
    P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084, P1_U3083,
    P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354, P2_U3353,
    P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347, P2_U3346,
    P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340, P2_U3339,
    P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333, P2_U3332,
    P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437, P2_U3438,
    P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320,
    P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313,
    P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306,
    P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299,
    P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
    P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
    P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502, P2_U3505,
    P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
    P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
    P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
    P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533, P2_U3534,
    P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541,
    P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548,
    P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294, P2_U3293,
    P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286,
    P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279,
    P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272,
    P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3265,
    P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258,
    P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251,
    P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3552,
    P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
    P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565, P2_U3566,
    P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572, P2_U3573,
    P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579, P2_U3580,
    P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
    P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
    P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
    P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
    P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152, P2_U3151,
    P2_U3966;
  wire n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
    n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
    n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
    n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
    n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
    n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
    n1094, n1095, n1096, n1098, n1100, n1101, n1103, n1104, n1106, n1108,
    n1110, n1112, n1114, n1116, n1118, n1120, n1122, n1124, n1126, n1128,
    n1130, n1132, n1134, n1135, n1136, n1137, n1138, n1139, n1142, n1144,
    n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
    n1156, n1157, n1158, n1159, n1160, n1162, n1163, n1165, n1166, n1167,
    n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
    n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1188,
    n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
    n1199, n1200, n1201, n1202, n1204, n1205, n1206, n1207, n1208, n1209,
    n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1219, n1220,
    n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
    n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
    n1241, n1242, n1243, n1244, n1246, n1247, n1248, n1249, n1250, n1251,
    n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
    n1262, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
    n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
    n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
    n1293, n1294, n1295, n1296, n1298, n1299, n1300, n1301, n1302, n1303,
    n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
    n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1322, n1323, n1324,
    n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
    n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
    n1345, n1346, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
    n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
    n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
    n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
    n1387, n1388, n1389, n1390, n1392, n1393, n1394, n1395, n1396, n1397,
    n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
    n1408, n1409, n1410, n1411, n1413, n1414, n1415, n1416, n1417, n1418,
    n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
    n1429, n1430, n1431, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
    n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
    n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
    n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
    n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
    n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
    n1492, n1493, n1494, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
    n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
    n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
    n1523, n1524, n1525, n1526, n1528, n1529, n1530, n1531, n1532, n1533,
    n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
    n1544, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
    n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
    n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1574, n1575,
    n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
    n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
    n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
    n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
    n1617, n1618, n1619, n1620, n1622, n1623, n1624, n1625, n1626, n1627,
    n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
    n1638, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
    n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
    n1659, n1660, n1661, n1662, n1664, n1665, n1666, n1667, n1668, n1669,
    n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
    n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1690,
    n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
    n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
    n1711, n1712, n1713, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
    n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
    n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
    n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
    n1753, n1754, n1755, n1756, n1757, n1759, n1760, n1761, n1762, n1763,
    n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
    n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1783, n1784,
    n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
    n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
    n1805, n1806, n1807, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
    n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
    n1826, n1827, n1828, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
    n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
    n1847, n1848, n1849, n1850, n1852, n1853, n1854, n1855, n1856, n1857,
    n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
    n1868, n1869, n1870, n1871, n1873, n1874, n1875, n1876, n1877, n1878,
    n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
    n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1897, n1898, n1900,
    n1902, n1904, n1906, n1908, n1910, n1912, n1914, n1916, n1918, n1920,
    n1922, n1924, n1926, n1928, n1930, n1932, n1934, n1936, n1938, n1940,
    n1942, n1944, n1946, n1948, n1950, n1952, n1954, n1956, n1958, n1960,
    n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
    n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
    n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
    n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
    n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
    n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
    n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
    n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
    n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
    n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
    n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
    n2071, n2072, n2073, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
    n2082, n2083, n2084, n2085, n2086, n2087, n2089, n2090, n2091, n2092,
    n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
    n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
    n2113, n2114, n2115, n2116, n2118, n2119, n2120, n2121, n2122, n2123,
    n2124, n2125, n2126, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
    n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
    n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
    n2155, n2156, n2157, n2158, n2159, n2161, n2162, n2163, n2164, n2165,
    n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
    n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
    n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
    n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
    n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2216,
    n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2227, n2228,
    n2229, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
    n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
    n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
    n2264, n2265, n2266, n2267, n2268, n2270, n2271, n2272, n2273, n2274,
    n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
    n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
    n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
    n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
    n2315, n2316, n2317, n2318, n2319, n2320, n2322, n2323, n2324, n2325,
    n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
    n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
    n2346, n2347, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
    n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
    n2367, n2368, n2369, n2370, n2371, n2373, n2374, n2375, n2376, n2377,
    n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
    n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
    n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
    n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2418,
    n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2428, n2429,
    n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
    n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
    n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
    n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
    n2471, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
    n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
    n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
    n2502, n2503, n2504, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
    n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
    n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
    n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
    n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2553,
    n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
    n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
    n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
    n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
    n2594, n2595, n2596, n2597, n2598, n2599, n2601, n2602, n2603, n2604,
    n2605, n2606, n2607, n2608, n2609, n2611, n2612, n2613, n2614, n2615,
    n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
    n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
    n2636, n2637, n2638, n2639, n2640, n2642, n2643, n2644, n2645, n2646,
    n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
    n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
    n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
    n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
    n2687, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
    n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
    n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
    n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
    n2728, n2729, n2730, n2731, n2733, n2734, n2735, n2736, n2737, n2738,
    n2739, n2740, n2741, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
    n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
    n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
    n2770, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
    n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
    n2791, n2792, n2793, n2794, n2796, n2797, n2798, n2799, n2800, n2801,
    n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
    n2812, n2813, n2814, n2815, n2816, n2817, n2819, n2820, n2821, n2822,
    n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
    n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
    n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
    n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
    n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2871, n2872, n2873,
    n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2883, n2884, n2885,
    n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
    n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
    n2906, n2907, n2908, n2909, n2910, n2911, n2913, n2914, n2915, n2916,
    n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
    n2927, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
    n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
    n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2956, n2957, n2958,
    n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
    n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
    n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
    n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
    n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
    n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
    n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
    n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
    n3040, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
    n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
    n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
    n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3079, n3080, n3081,
    n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
    n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
    n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
    n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
    n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
    n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
    n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
    n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
    n3163, n3164, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
    n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
    n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
    n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
    n3204, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
    n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
    n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
    n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
    n3245, n3246, n3247, n3249, n3250, n3252, n3253, n3254, n3255, n3256,
    n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
    n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
    n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
    n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3297,
    n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
    n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
    n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
    n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3336, n3337, n3338,
    n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
    n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3358, n3359,
    n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
    n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3379, n3380,
    n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3391,
    n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
    n3403, n3404, n3405, n3407, n3409, n3411, n3413, n3415, n3417, n3419,
    n3421, n3423, n3425, n3427, n3429, n3431, n3433, n3435, n3437, n3439,
    n3441, n3443, n3445, n3447, n3449, n3451, n3453, n3455, n3457, n3459,
    n3461, n3463, n3465, n3467, n3469, n3470, n3471, n3472, n3473, n3474,
    n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
    n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3494, n3495,
    n3496, n3497, n3498, n3500, n3501, n3502, n3503, n3504, n3505, n3507,
    n3508, n3509, n3510, n3511, n3512, n3514, n3515, n3516, n3517, n3518,
    n3519, n3520, n3521, n3522, n3523, n3524, n3526, n3527, n3528, n3529,
    n3530, n3531, n3533, n3534, n3535, n3536, n3537, n3538, n3540, n3541,
    n3542, n3543, n3544, n3545, n3547, n3548, n3549, n3550, n3551, n3552,
    n3553, n3554, n3556, n3557, n3558, n3559, n3560, n3561, n3563, n3564,
    n3565, n3566, n3567, n3568, n3570, n3571, n3572, n3573, n3574, n3575,
    n3576, n3577, n3578, n3580, n3581, n3582, n3583, n3584, n3585, n3587,
    n3588, n3589, n3590, n3591, n3592, n3594, n3595, n3596, n3597, n3598,
    n3599, n3601, n3602, n3603, n3604, n3605, n3607, n3608, n3609, n3610,
    n3611, n3612, n3614, n3615, n3616, n3617, n3618, n3619, n3621, n3622,
    n3623, n3624, n3625, n3626, n3628, n3629, n3630, n3631, n3632, n3633,
    n3634, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3644, n3645,
    n3646, n3647, n3648, n3649, n3650, n3652, n3653, n3654, n3655, n3656,
    n3657, n3658, n3659, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
    n3668, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3679,
    n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3689, n3690,
    n3691, n3692, n3693, n3694, n3695, n3697, n3698, n3699, n3700, n3701,
    n3702, n3703, n3704, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
    n3713, n3714, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3724,
    n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3733, n3734, n3735,
    n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
    n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
    n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
    n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
    n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
    n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
    n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
    n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
    n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
    n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
    n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
    n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
    n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
    n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
    n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
    n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
    n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
    n3910, n3912, n3913, n3914, n3915, n3916, n3918, n3919, n3920, n3921,
    n3922, n3923, n3924, n3925, n3926, n3927, n3929, n3930, n3931, n3932,
    n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
    n3945, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
    n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
    n3966, n3967, n3968, n3970, n3971, n3972, n3973, n3974, n3976, n3977,
    n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3986, n3987, n3988,
    n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3999,
    n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
    n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
    n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
    n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4042, n4043,
    n4044, n4045, n4046, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
    n4055, n4057, n4058, n4059, n4060, n4061, n4063, n4064, n4065, n4066,
    n4067, n4068, n4069, n4070, n4072, n4073, n4074, n4075, n4076, n4077,
    n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087,
    n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097,
    n4099, n4101, n4102, n4103, n4104, n4106, n4107, n4108, n4109, n4110,
    n4111, n4112, n4113, n4115, n4116, n4117, n4119, n4120, n4121, n4123,
    n4124, n4125, n4126, n4127, n4128, n4129, n4131, n4132, n4133, n4134,
    n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
    n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4153, n4154, n4156,
    n4157, n4158, n4159, n4160, n4162, n4163, n4164, n4165, n4166, n4168,
    n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
    n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
    n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
    n4199, n4200, n4201, n4204, n4205, n4206, n4207, n4208, n4209, n4210,
    n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
    n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4229, n4230, n4231,
    n4232, n4233, n4234, n4236, n4237, n4238, n4239, n4240, n4241, n4243,
    n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
    n4254, n4255, n4256, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
    n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
    n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
    n4286, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4297,
    n4299, n4301, n4303, n4305, n4307, n4309, n4311, n4313, n4315, n4317,
    n4319, n4321, n4323, n4325, n4327, n4329, n4331, n4333, n4335, n4337,
    n4339, n4341, n4343, n4345, n4347, n4349, n4351, n4353, n4355, n4357,
    n4358, n4360, n4361, n4363, n4364, n4365, n4366, n4372, n4374, n4375,
    n4377, n4378, n4380, n4383, n4387, n4388, n4389, n4390, n4391, n4392,
    n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4404,
    n4405, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
    n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
    n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
    n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
    n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
    n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
    n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
    n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
    n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
    n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
    n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4514, n4515, n4516,
    n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526,
    n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4535, n4536, n4537,
    n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
    n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
    n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
    n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
    n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
    n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
    n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
    n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
    n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
    n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
    n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
    n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
    n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
    n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
    n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
    n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
    n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
    n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
    n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
    n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4738,
    n4741, n4742, n4744, n4745, n4747, n4749, n4752, n4753, n4754, n4755,
    n4757, n4760, n4761, n4762, n4763, n4767, n4768, n4770, n4771, n4772,
    n4774, n4777, n4778, n4779, n4780, n4782, n4784, n4785, n4786, n4787,
    n4788, n4790, n4791, n4792, n4793, n4794, n4796, n4799, n4800, n4801,
    n4802, n4803, n4804, n4805, n4806, n4808, n4809, n4811, n4812, n4813,
    n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
    n4824, n4825, n4826, n4827, n4828, n4831, n4832, n4833, n4834, n4835,
    n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
    n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
    n4856, n4857, n4858, n4859, n4860, n4861, n4863, n4864, n4865, n4866,
    n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876,
    n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886,
    n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896,
    n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906,
    n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916,
    n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926,
    n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936,
    n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946,
    n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956,
    n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966,
    n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976,
    n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986,
    n4987, n4988, n4989, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
    n4998, n5000, n5001, n5002, n5004, n5005, n5006, n5007, n5008, n5009,
    n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
    n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
    n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
    n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
    n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
    n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
    n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
    n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
    n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
    n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
    n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
    n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
    n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
    n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
    n5150, n5151, n5152, n5153, n5155, n5156, n5157, n5158, n5159, n5160,
    n5161, n5162, n5163, n5164, n5165, n5166, n5168, n5169, n5170, n5171,
    n5172, n5173, n5174, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
    n5183, n5184, n5185, n5186, n5187, n5189, n5190, n5191, n5192, n5193,
    n5194, n5195, n5196, n5197, n5198, n5200, n5201, n5202, n5203, n5204,
    n5205, n5206, n5207, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
    n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5225, n5226,
    n5227, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5237, n5238,
    n5239, n5240, n5241, n5242, n5243, n5245, n5246, n5247, n5248, n5249,
    n5250, n5251, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
    n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5272,
    n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
    n5283, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5294,
    n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
    n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5316,
    n5317, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
    n5328, n5329, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
    n5339, n5340, n5341, n5342, n5343, n5345, n5346, n5347, n5348, n5349,
    n5350, n5351, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5361,
    n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
    n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
    n5382, n5383, n5384, n5385, n5386, n5388, n5389, n5390, n5391, n5392,
    n5393, n5394, n5395, n5396, n5397, n5399, n5400, n5401, n5402, n5403,
    n5404, n5405, n5406, n5407, n5408, n5409, n5411, n5412, n5413, n5414,
    n5415, n5416, n5417, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
    n5426, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5436, n5437,
    n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
    n5448, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
    n5459, n5460, n5462, n5463, n5464, n5466, n5467, n5469, n5470, n5471,
    n5472, n5473, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5483,
    n5484, n5485, n5486, n5487, n5488, n5490, n5491, n5492, n5493, n5494,
    n5495, n5497, n5498, n5499, n5500, n5501, n5503, n5504, n5505, n5506,
    n5507, n5508, n5509, n5510, n5511, n5513, n5514, n5515, n5516, n5517,
    n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5528, n5529,
    n5530, n5531, n5532, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
    n5541, n5543, n5544, n5545, n5546, n5547, n5549, n5550, n5551, n5552,
    n5553, n5554, n5555, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
    n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5573, n5574, n5575,
    n5576, n5577, n5578, n5580, n5581, n5582, n5583, n5584, n5585, n5587,
    n5588, n5590, n5591, n5592, n5593, n5594, n5596, n5597, n5598, n5599,
    n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
    n5610, n5611, n5612, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
    n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5631, n5632,
    n5633, n5636, n5637, n5638, n5639, n5641, n5642, n5643, n5644, n5645,
    n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5654, n5655, n5656,
    n5657, n5658, n5659, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
    n5668, n5669, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5679,
    n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5690,
    n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
    n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5710, n5711, n5712,
    n5713, n5714, n5715, n5716, n5718, n5719, n5720, n5721, n5722, n5723,
    n5724, n5726, n5727, n5728, n5729, n5730, n5731, n5733, n5734, n5735,
    n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
    n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5754, n5755, n5756,
    n5758, n5760, n5762, n5764, n5766, n5768, n5770, n5772, n5774, n5776,
    n5778, n5780, n5782, n5784, n5786, n5788, n5790, n5792, n5794, n5796,
    n5798, n5800, n5802, n5804, n5806, n5808, n5810, n5812, n5814, n5816,
    n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
    n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
    n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
    n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
    n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
    n5868, n5869, n5870, n5871, n5875, n5876, n5877, n5878, n5879, n5880,
    n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
    n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5900, n5901,
    n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
    n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
    n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
    n5932, n5933, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
    n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
    n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
    n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
    n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5981, n5982, n5983,
    n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
    n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
    n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
    n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6022, n6023, n6024,
    n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
    n6035, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
    n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
    n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
    n6066, n6067, n6068, n6069, n6071, n6072, n6073, n6074, n6075, n6076,
    n6077, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
    n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
    n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
    n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
    n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6128, n6129,
    n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
    n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
    n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
    n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
    n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6179, n6180,
    n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
    n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
    n6201, n6202, n6203, n6204, n6206, n6207, n6208, n6209, n6210, n6211,
    n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
    n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6230, n6231, n6232,
    n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
    n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
    n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
    n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
    n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6282, n6283,
    n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
    n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
    n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
    n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
    n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6334, n6335,
    n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
    n6346, n6347, n6348, n6349, n6351, n6352, n6353, n6354, n6355, n6356,
    n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366,
    n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376,
    n6377, n6378, n6379, n6381, n6382, n6383, n6384, n6385, n6386, n6387,
    n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397,
    n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407,
    n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417,
    n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427,
    n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6437, n6438,
    n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
    n6449, n6450, n6451, n6452, n6453, n6454, n6456, n6457, n6458, n6459,
    n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6470,
    n6471, n6472, n6473, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
    n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
    n6496, n6497, n6498, n6499, n6501, n6502, n6503, n6504, n6505, n6506,
    n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516,
    n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6525, n6526, n6527,
    n6528, n6529, n6530, n6532, n6534, n6535, n6536, n6537, n6538, n6539,
    n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
    n6550, n6551, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
    n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6573,
    n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
    n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
    n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6604,
    n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
    n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6626,
    n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636,
    n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646,
    n6647, n6648, n6649, n6650, n6651, n6653, n6654, n6655, n6656, n6657,
    n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667,
    n6668, n6669, n6670, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
    n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
    n6690, n6691, n6692, n6693, n6694, n6695, n6697, n6698, n6699, n6700,
    n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
    n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6723, n6724,
    n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
    n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
    n6745, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
    n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
    n6766, n6771, n6772, n6773, n6774, n6776, n6778, n6779, n6780, n6781,
    n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
    n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
    n6802, n6803, n6804, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
    n6813, n6814, n6815, n6816, n6817, n6818, n6821, n6822, n6826, n6827,
    n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837,
    n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847,
    n6848, n6849, n6850, n6851, n6853, n6854, n6855, n6856, n6857, n6858,
    n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
    n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6879, n6880, n6881,
    n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
    n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6901, n6902,
    n6903, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
    n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
    n6924, n6925, n6926, n6931, n6932, n6933, n6934, n6935, n6936, n6937,
    n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947,
    n6948, n6949, n6950, n6951, n6952, n6954, n6955, n6956, n6957, n6958,
    n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
    n6969, n6970, n6971, n6972, n6973, n6977, n6978, n6979, n6980, n6981,
    n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
    n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7002,
    n7003, n7004, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
    n7014, n7015, n7016, n7017, n7018, n7022, n7023, n7024, n7025, n7026,
    n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
    n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7045, n7046, n7047,
    n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
    n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7070,
    n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
    n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7090, n7091,
    n7092, n7094, n7095, n7096, n7098, n7099, n7100, n7101, n7102, n7103,
    n7104, n7107, n7108, n7109, n7113, n7114, n7115, n7116, n7117, n7118,
    n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
    n7129, n7130, n7131, n7132, n7134, n7135, n7136, n7138, n7139, n7140,
    n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7151,
    n7152, n7153, n7154, n7155, n7159, n7160, n7161, n7162, n7163, n7164,
    n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
    n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7183, n7184, n7185,
    n7186, n7187, n7188, n7190, n7191, n7192, n7193, n7194, n7195, n7196,
    n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206,
    n7207, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
    n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
    n7231, n7232, n7233, n7235, n7236, n7238, n7240, n7241, n7242, n7243,
    n7244, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
    n7255, n7256, n7257, n7258, n7259, n7265, n7266, n7267, n7268, n7269,
    n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
    n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7290,
    n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300,
    n7301, n7302, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
    n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
    n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7332, n7333, n7334,
    n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
    n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
    n7355, n7356, n7357, n7358, n7360, n7361, n7362, n7363, n7364, n7365,
    n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
    n7376, n7377, n7378, n7381, n7382, n7383, n7384, n7385, n7386, n7387,
    n7388, n7389, n7390, n7391, n7393, n7394, n7395, n7396, n7397, n7398,
    n7399, n7400, n7401, n7402, n7403, n7404, n7406, n7407, n7408, n7409,
    n7410, n7411, n7412, n7413, n7415, n7416, n7417, n7419, n7421, n7423,
    n7425, n7427, n7429, n7431, n7433, n7435, n7437, n7439, n7441, n7443,
    n7445, n7447, n7449, n7451, n7453, n7455, n7457, n7459, n7461, n7463,
    n7465, n7467, n7469, n7471, n7473, n7475, n7477, n7479, n7481, n7482,
    n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
    n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7502, n7503,
    n7504, n7505, n7506, n7508, n7509, n7510, n7511, n7513, n7514, n7515,
    n7516, n7517, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
    n7527, n7528, n7530, n7531, n7532, n7533, n7534, n7536, n7537, n7538,
    n7539, n7540, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7550,
    n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7560, n7561,
    n7562, n7563, n7564, n7565, n7566, n7568, n7569, n7570, n7571, n7572,
    n7573, n7574, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
    n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7594, n7595,
    n7596, n7597, n7598, n7599, n7600, n7601, n7603, n7604, n7605, n7606,
    n7607, n7608, n7609, n7611, n7612, n7613, n7614, n7615, n7616, n7617,
    n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7628, n7629,
    n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7638, n7639, n7640,
    n7641, n7642, n7643, n7644, n7645, n7647, n7648, n7649, n7650, n7651,
    n7652, n7653, n7654, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
    n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7673, n7674,
    n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7683, n7684, n7685,
    n7686, n7687, n7688, n7689, n7691, n7692, n7693, n7694, n7695, n7696,
    n7697, n7699, n7700, n7701, n7702, n7703, n7704, n7706, n7707, n7708,
    n7709, n7710, n7711, n7712, n7714, n7715, n7716, n7717, n7718, n7719,
    n7720, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7731,
    n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7740, n7741, n7742,
    n7743, n7745, n7746, n7747, n7748, n7750, n7751, n7752, n7753, n7754,
    n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
    n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
    n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
    n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
    n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
    n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
    n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
    n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
    n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
    n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
    n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
    n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
    n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
    n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
    n7895, n7896, n7897, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
    n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7915, n7916,
    n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926,
    n7927, n7928, n7929, n7931, n7932, n7933, n7934, n7935, n7936, n7937,
    n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947,
    n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7956, n7957, n7959,
    n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
    n7970, n7971, n7972, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
    n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7990, n7991,
    n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001,
    n8002, n8003, n8004, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
    n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
    n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
    n8033, n8034, n8035, n8036, n8037, n8039, n8041, n8042, n8043, n8044,
    n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
    n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
    n8066, n8067, n8068, n8069, n8070, n8072, n8073, n8074, n8075, n8076,
    n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086,
    n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096,
    n8097, n8099, n8101, n8102, n8103, n8104, n8106, n8107, n8108, n8109,
    n8110, n8111, n8112, n8113, n8114, n8115, n8117, n8118, n8120, n8121,
    n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
    n8132, n8133, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
    n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
    n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8163,
    n8164, n8166, n8167, n8168, n8169, n8171, n8172, n8173, n8174, n8175,
    n8176, n8177, n8178, n8179, n8181, n8182, n8183, n8184, n8185, n8186,
    n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196,
    n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206,
    n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216,
    n8217, n8218, n8220, n8222, n8223, n8224, n8225, n8227, n8228, n8229,
    n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8238, n8239, n8240,
    n8241, n8242, n8243, n8244, n8245, n8246, n8248, n8249, n8250, n8251,
    n8252, n8253, n8254, n8255, n8256, n8257, n8259, n8260, n8261, n8262,
    n8263, n8264, n8265, n8266, n8268, n8269, n8270, n8271, n8272, n8273,
    n8274, n8275, n8276, n8277, n8278, n8280, n8281, n8282, n8283, n8284,
    n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
    n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
    n8306, n8307, n8308, n8310, n8312, n8314, n8316, n8318, n8320, n8322,
    n8324, n8326, n8328, n8330, n8332, n8334, n8336, n8338, n8340, n8342,
    n8344, n8346, n8348, n8350, n8352, n8354, n8356, n8358, n8360, n8362,
    n8364, n8366, n8368, n8370, n8372, n8374, n8375, n8376, n8377, n8378,
    n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
    n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
    n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
    n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
    n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
    n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
    n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
    n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
    n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
    n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
    n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
    n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
    n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
    n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
    n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
    n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
    n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
    n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
    n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
    n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
    n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
    n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
    n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
    n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
    n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
    n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8639, n8640,
    n8642, n8645, n8647, n8648, n8649, n8650, n8651, n8652, n8655, n8656,
    n8659, n8660, n8671, n8672, n8673, n8674, n8679, n8681, n8682, n8683,
    n8684, n8685, n8686, n8687, n8688, n8689, n8691, n8692, n8693, n8694,
    n8695, n8697, n8698, n8699, n8700, n8701, n8702, n8704, n8705, n8706,
    n8707, n8710, n8711, n8713, n8714, n8715, n8716, n8718, n8720, n8721,
    n8722, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
    n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8747, n8750, n8752,
    n8756, n8758, n8762, n8764, n8766, n8774, n8782, n8786, n8789, n8790,
    n8792, n8793, n8795, n8796, n8797, n8798, n8804, n8808, n8809, n8811,
    n8812, n8813, n8823, n8824, n8827, n8828, n8834, n8838, n8839, n8840,
    n8842, n8843, n8848, n8852, n8854, n8855, n8856, n8857, n8861, n8862,
    n8864, n8865, n8866, n8869, n8870, n8876, n8877, n8878, n8879, n8880,
    n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
    n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
    n8901, n8904, n8908, n8909, n8911, n8912, n8913, n8916, n8918, n8919,
    n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
    n8933, n8934, n8935, n8936, n8938, n8939, n8940, n8941, n8942, n8943,
    n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
    n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963,
    n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973,
    n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
    n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
    n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
    n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
    n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
    n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
    n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
    n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
    n9055, n9056, n9057, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
    n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
    n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
    n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
    n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
    n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
    n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
    n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
    n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
    n9146, n9148, n9149, n9150, n9151, n9152, n9153, n9155, n9156, n9158,
    n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9167, n9168, n9169,
    n9170, n9171, n9172, n9173, n9175, n9176, n9177, n9178, n9179, n9180,
    n9181, n9183, n9184, n9186, n9187, n9188, n9190, n9191, n9192, n9193,
    n9194, n9195, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9205,
    n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
    n9216, n9217, n9219, n9220, n9221, n9223, n9224, n9225, n9226, n9227,
    n9228, n9229, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
    n9239, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9249, n9250,
    n9251, n9252, n9253, n9254, n9255, n9256, n9258, n9259, n9260, n9261,
    n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9270, n9271, n9272,
    n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9283,
    n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9294,
    n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9304, n9306, n9307,
    n9308, n9309, n9310, n9311, n9312, n9314, n9316, n9317, n9318, n9319,
    n9320, n9321, n9322, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
    n9331, n9332, n9333, n9334, n9335, n9337, n9338, n9339, n9340, n9341,
    n9342, n9343, n9344, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
    n9353, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
    n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
    n9374, n9375, n9376, n9377, n9378, n9380, n9382, n9383, n9384, n9385,
    n9386, n9387, n9388, n9390, n9391, n9392, n9393, n9394, n9395, n9396,
    n9397, n9398, n9399, n9400, n9401, n9402, n9404, n9405, n9406, n9407,
    n9408, n9409, n9410, n9411, n9413, n9414, n9415, n9416, n9417, n9418,
    n9419, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9430,
    n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
    n9441, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451,
    n9452, n9453, n9454, n9455, n9456, n9458, n9459, n9460;
  NAND2X1 g0000(.A(P2_ADDR_REG_17__SCAN_IN), .B(P1_ADDR_REG_17__SCAN_IN), .Y(n1034));
  NOR2X1  g0001(.A(P2_ADDR_REG_17__SCAN_IN), .B(P1_ADDR_REG_17__SCAN_IN), .Y(n1035));
  NOR2X1  g0002(.A(P2_ADDR_REG_16__SCAN_IN), .B(P1_ADDR_REG_16__SCAN_IN), .Y(n1036));
  NAND2X1 g0003(.A(P2_ADDR_REG_15__SCAN_IN), .B(P1_ADDR_REG_15__SCAN_IN), .Y(n1037));
  NAND2X1 g0004(.A(P2_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), .Y(n1038));
  NAND2X1 g0005(.A(P2_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), .Y(n1039));
  NAND2X1 g0006(.A(P2_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), .Y(n1040));
  INVX1   g0007(.A(P1_ADDR_REG_11__SCAN_IN), .Y(n1041));
  INVX1   g0008(.A(P2_ADDR_REG_11__SCAN_IN), .Y(n1042));
  NAND2X1 g0009(.A(P2_ADDR_REG_10__SCAN_IN), .B(P1_ADDR_REG_10__SCAN_IN), .Y(n1043));
  INVX1   g0010(.A(P1_ADDR_REG_9__SCAN_IN), .Y(n1044));
  INVX1   g0011(.A(P2_ADDR_REG_9__SCAN_IN), .Y(n1045));
  NAND2X1 g0012(.A(P2_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), .Y(n1046));
  INVX1   g0013(.A(P1_ADDR_REG_7__SCAN_IN), .Y(n1047));
  INVX1   g0014(.A(P2_ADDR_REG_7__SCAN_IN), .Y(n1048));
  NAND2X1 g0015(.A(P2_ADDR_REG_6__SCAN_IN), .B(P1_ADDR_REG_6__SCAN_IN), .Y(n1049));
  NAND2X1 g0016(.A(P2_ADDR_REG_5__SCAN_IN), .B(P1_ADDR_REG_5__SCAN_IN), .Y(n1050));
  NAND2X1 g0017(.A(P2_ADDR_REG_4__SCAN_IN), .B(P1_ADDR_REG_4__SCAN_IN), .Y(n1051));
  INVX1   g0018(.A(P1_ADDR_REG_3__SCAN_IN), .Y(n1052));
  INVX1   g0019(.A(P2_ADDR_REG_3__SCAN_IN), .Y(n1053));
  NAND2X1 g0020(.A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Y(n1054));
  INVX1   g0021(.A(P2_ADDR_REG_1__SCAN_IN), .Y(n1055));
  NAND3X1 g0022(.A(P2_ADDR_REG_0__SCAN_IN), .B(P1_ADDR_REG_0__SCAN_IN), .C(P1_ADDR_REG_1__SCAN_IN), .Y(n1056));
  AOI21X1 g0023(.A0(P2_ADDR_REG_0__SCAN_IN), .A1(P1_ADDR_REG_0__SCAN_IN), .B0(P1_ADDR_REG_1__SCAN_IN), .Y(n1057));
  OAI21X1 g0024(.A0(n1057), .A1(n1055), .B0(n1056), .Y(n1058));
  OAI21X1 g0025(.A0(P2_ADDR_REG_2__SCAN_IN), .A1(P1_ADDR_REG_2__SCAN_IN), .B0(n1058), .Y(n1059));
  NAND2X1 g0026(.A(n1059), .B(n1054), .Y(n1060));
  OAI21X1 g0027(.A0(P2_ADDR_REG_3__SCAN_IN), .A1(P1_ADDR_REG_3__SCAN_IN), .B0(n1060), .Y(n1061));
  OAI21X1 g0028(.A0(n1053), .A1(n1052), .B0(n1061), .Y(n1062));
  OAI21X1 g0029(.A0(P2_ADDR_REG_4__SCAN_IN), .A1(P1_ADDR_REG_4__SCAN_IN), .B0(n1062), .Y(n1063));
  NAND2X1 g0030(.A(n1063), .B(n1051), .Y(n1064));
  OAI21X1 g0031(.A0(P2_ADDR_REG_5__SCAN_IN), .A1(P1_ADDR_REG_5__SCAN_IN), .B0(n1064), .Y(n1065));
  NAND2X1 g0032(.A(n1065), .B(n1050), .Y(n1066));
  OAI21X1 g0033(.A0(P2_ADDR_REG_6__SCAN_IN), .A1(P1_ADDR_REG_6__SCAN_IN), .B0(n1066), .Y(n1067));
  NAND2X1 g0034(.A(n1067), .B(n1049), .Y(n1068));
  OAI21X1 g0035(.A0(P2_ADDR_REG_7__SCAN_IN), .A1(P1_ADDR_REG_7__SCAN_IN), .B0(n1068), .Y(n1069));
  OAI21X1 g0036(.A0(n1048), .A1(n1047), .B0(n1069), .Y(n1070));
  OAI21X1 g0037(.A0(P2_ADDR_REG_8__SCAN_IN), .A1(P1_ADDR_REG_8__SCAN_IN), .B0(n1070), .Y(n1071));
  NAND2X1 g0038(.A(n1071), .B(n1046), .Y(n1072));
  OAI21X1 g0039(.A0(P2_ADDR_REG_9__SCAN_IN), .A1(P1_ADDR_REG_9__SCAN_IN), .B0(n1072), .Y(n1073));
  OAI21X1 g0040(.A0(n1045), .A1(n1044), .B0(n1073), .Y(n1074));
  OAI21X1 g0041(.A0(P2_ADDR_REG_10__SCAN_IN), .A1(P1_ADDR_REG_10__SCAN_IN), .B0(n1074), .Y(n1075));
  NAND2X1 g0042(.A(n1075), .B(n1043), .Y(n1076));
  OAI21X1 g0043(.A0(P2_ADDR_REG_11__SCAN_IN), .A1(P1_ADDR_REG_11__SCAN_IN), .B0(n1076), .Y(n1077));
  OAI21X1 g0044(.A0(n1042), .A1(n1041), .B0(n1077), .Y(n1078));
  OAI21X1 g0045(.A0(P2_ADDR_REG_12__SCAN_IN), .A1(P1_ADDR_REG_12__SCAN_IN), .B0(n1078), .Y(n1079));
  NAND2X1 g0046(.A(n1079), .B(n1040), .Y(n1080));
  OAI21X1 g0047(.A0(P2_ADDR_REG_13__SCAN_IN), .A1(P1_ADDR_REG_13__SCAN_IN), .B0(n1080), .Y(n1081));
  NAND2X1 g0048(.A(n1081), .B(n1039), .Y(n1082));
  OAI21X1 g0049(.A0(P2_ADDR_REG_14__SCAN_IN), .A1(P1_ADDR_REG_14__SCAN_IN), .B0(n1082), .Y(n1083));
  NAND2X1 g0050(.A(n1083), .B(n1038), .Y(n1084));
  OAI21X1 g0051(.A0(P2_ADDR_REG_15__SCAN_IN), .A1(P1_ADDR_REG_15__SCAN_IN), .B0(n1084), .Y(n1085));
  AOI21X1 g0052(.A0(n1085), .A1(n1037), .B0(n1036), .Y(n1086));
  AOI21X1 g0053(.A0(P2_ADDR_REG_16__SCAN_IN), .A1(P1_ADDR_REG_16__SCAN_IN), .B0(n1086), .Y(n1087));
  OAI21X1 g0054(.A0(n1087), .A1(n1035), .B0(n1034), .Y(n1088));
  AOI21X1 g0055(.A0(P2_ADDR_REG_18__SCAN_IN), .A1(P1_ADDR_REG_18__SCAN_IN), .B0(n1088), .Y(n1089));
  INVX1   g0056(.A(P1_ADDR_REG_19__SCAN_IN), .Y(n1090));
  XOR2X1  g0057(.A(P2_ADDR_REG_19__SCAN_IN), .B(n1090), .Y(n1091));
  INVX1   g0058(.A(n1091), .Y(n1092));
  OAI21X1 g0059(.A0(P2_ADDR_REG_18__SCAN_IN), .A1(P1_ADDR_REG_18__SCAN_IN), .B0(n1092), .Y(n1093));
  NOR2X1  g0060(.A(n1093), .B(n1089), .Y(n1094));
  OAI21X1 g0061(.A0(P2_ADDR_REG_18__SCAN_IN), .A1(P1_ADDR_REG_18__SCAN_IN), .B0(n1088), .Y(n1095));
  AOI21X1 g0062(.A0(P2_ADDR_REG_18__SCAN_IN), .A1(P1_ADDR_REG_18__SCAN_IN), .B0(n1092), .Y(n1096));
  AOI21X1 g0063(.A0(n1096), .A1(n1095), .B0(n1094), .Y(ADD_1071_U4));
  XOR2X1  g0064(.A(P2_ADDR_REG_18__SCAN_IN), .B(P1_ADDR_REG_18__SCAN_IN), .Y(n1098));
  XOR2X1  g0065(.A(n1098), .B(n1088), .Y(ADD_1071_U55));
  INVX1   g0066(.A(P1_ADDR_REG_17__SCAN_IN), .Y(n1100));
  XOR2X1  g0067(.A(P2_ADDR_REG_17__SCAN_IN), .B(n1100), .Y(n1101));
  XOR2X1  g0068(.A(n1101), .B(n1087), .Y(ADD_1071_U56));
  NAND2X1 g0069(.A(n1085), .B(n1037), .Y(n1103));
  XOR2X1  g0070(.A(P2_ADDR_REG_16__SCAN_IN), .B(P1_ADDR_REG_16__SCAN_IN), .Y(n1104));
  XOR2X1  g0071(.A(n1104), .B(n1103), .Y(ADD_1071_U57));
  XOR2X1  g0072(.A(P2_ADDR_REG_15__SCAN_IN), .B(P1_ADDR_REG_15__SCAN_IN), .Y(n1106));
  XOR2X1  g0073(.A(n1106), .B(n1084), .Y(ADD_1071_U58));
  XOR2X1  g0074(.A(P2_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), .Y(n1108));
  XOR2X1  g0075(.A(n1108), .B(n1082), .Y(ADD_1071_U59));
  XOR2X1  g0076(.A(P2_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), .Y(n1110));
  XOR2X1  g0077(.A(n1110), .B(n1080), .Y(ADD_1071_U60));
  XOR2X1  g0078(.A(P2_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), .Y(n1112));
  XOR2X1  g0079(.A(n1112), .B(n1078), .Y(ADD_1071_U61));
  XOR2X1  g0080(.A(P2_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), .Y(n1114));
  XOR2X1  g0081(.A(n1114), .B(n1076), .Y(ADD_1071_U62));
  XOR2X1  g0082(.A(P2_ADDR_REG_10__SCAN_IN), .B(P1_ADDR_REG_10__SCAN_IN), .Y(n1116));
  XOR2X1  g0083(.A(n1116), .B(n1074), .Y(ADD_1071_U63));
  XOR2X1  g0084(.A(P2_ADDR_REG_9__SCAN_IN), .B(P1_ADDR_REG_9__SCAN_IN), .Y(n1118));
  XOR2X1  g0085(.A(n1118), .B(n1072), .Y(ADD_1071_U47));
  XOR2X1  g0086(.A(P2_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), .Y(n1120));
  XOR2X1  g0087(.A(n1120), .B(n1070), .Y(ADD_1071_U48));
  XOR2X1  g0088(.A(P2_ADDR_REG_7__SCAN_IN), .B(P1_ADDR_REG_7__SCAN_IN), .Y(n1122));
  XOR2X1  g0089(.A(n1122), .B(n1068), .Y(ADD_1071_U49));
  XOR2X1  g0090(.A(P2_ADDR_REG_6__SCAN_IN), .B(P1_ADDR_REG_6__SCAN_IN), .Y(n1124));
  XOR2X1  g0091(.A(n1124), .B(n1066), .Y(ADD_1071_U50));
  XOR2X1  g0092(.A(P2_ADDR_REG_5__SCAN_IN), .B(P1_ADDR_REG_5__SCAN_IN), .Y(n1126));
  XOR2X1  g0093(.A(n1126), .B(n1064), .Y(ADD_1071_U51));
  XOR2X1  g0094(.A(P2_ADDR_REG_4__SCAN_IN), .B(P1_ADDR_REG_4__SCAN_IN), .Y(n1128));
  XOR2X1  g0095(.A(n1128), .B(n1062), .Y(ADD_1071_U52));
  XOR2X1  g0096(.A(P2_ADDR_REG_3__SCAN_IN), .B(P1_ADDR_REG_3__SCAN_IN), .Y(n1130));
  XOR2X1  g0097(.A(n1130), .B(n1060), .Y(ADD_1071_U53));
  XOR2X1  g0098(.A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Y(n1132));
  XOR2X1  g0099(.A(n1132), .B(n1058), .Y(ADD_1071_U54));
  NAND2X1 g0100(.A(P2_ADDR_REG_0__SCAN_IN), .B(P1_ADDR_REG_0__SCAN_IN), .Y(n1134));
  XOR2X1  g0101(.A(n1134), .B(P2_ADDR_REG_1__SCAN_IN), .Y(n1135));
  NOR2X1  g0102(.A(n1056), .B(n1055), .Y(n1136));
  INVX1   g0103(.A(P1_ADDR_REG_1__SCAN_IN), .Y(n1137));
  NOR2X1  g0104(.A(P2_ADDR_REG_1__SCAN_IN), .B(n1137), .Y(n1138));
  AOI21X1 g0105(.A0(n1138), .A1(n1134), .B0(n1136), .Y(n1139));
  OAI21X1 g0106(.A0(n1135), .A1(P1_ADDR_REG_1__SCAN_IN), .B0(n1139), .Y(ADD_1071_U5));
  XOR2X1  g0107(.A(P2_ADDR_REG_0__SCAN_IN), .B(P1_ADDR_REG_0__SCAN_IN), .Y(ADD_1071_U46));
  INVX1   g0108(.A(P2_RD_REG_SCAN_IN), .Y(n1142));
  XOR2X1  g0109(.A(P1_RD_REG_SCAN_IN), .B(n1142), .Y(U126));
  INVX1   g0110(.A(P2_WR_REG_SCAN_IN), .Y(n1144));
  XOR2X1  g0111(.A(P1_WR_REG_SCAN_IN), .B(n1144), .Y(U123));
  NAND3X1 g0112(.A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), .C(n1142), .Y(n1146));
  NOR2X1  g0113(.A(P2_ADDR_REG_19__SCAN_IN), .B(P1_RD_REG_SCAN_IN), .Y(n1147));
  NAND2X1 g0114(.A(n1147), .B(n1090), .Y(n1148));
  NAND2X1 g0115(.A(n1148), .B(n1146), .Y(n1149));
  INVX1   g0116(.A(P2_DATAO_REG_0__SCAN_IN), .Y(n1150));
  INVX1   g0117(.A(P2_ADDR_REG_19__SCAN_IN), .Y(n1151));
  NOR3X1  g0118(.A(n1151), .B(n1090), .C(P2_RD_REG_SCAN_IN), .Y(n1152));
  NOR3X1  g0119(.A(P2_ADDR_REG_19__SCAN_IN), .B(P1_RD_REG_SCAN_IN), .C(P1_ADDR_REG_19__SCAN_IN), .Y(n1153));
  NOR3X1  g0120(.A(n1153), .B(n1152), .C(n1150), .Y(n1154));
  INVX1   g0121(.A(SI_0_), .Y(n1155));
  NOR2X1  g0122(.A(n1153), .B(n1152), .Y(n1156));
  AOI21X1 g0123(.A0(n1148), .A1(n1146), .B0(n1150), .Y(n1157));
  AOI21X1 g0124(.A0(n1156), .A1(P1_DATAO_REG_0__SCAN_IN), .B0(n1157), .Y(n1158));
  XOR2X1  g0125(.A(n1158), .B(n1155), .Y(n1159));
  AOI21X1 g0126(.A0(n1159), .A1(n1149), .B0(n1154), .Y(n1160));
  INVX1   g0127(.A(P1_STATE_REG_SCAN_IN), .Y(P1_U3084));
  NOR2X1  g0128(.A(P1_U3084), .B(P1_IR_REG_31__SCAN_IN), .Y(n1162));
  OAI21X1 g0129(.A0(n1162), .A1(P1_STATE_REG_SCAN_IN), .B0(P1_IR_REG_0__SCAN_IN), .Y(n1163));
  OAI21X1 g0130(.A0(n1160), .A1(P1_STATE_REG_SCAN_IN), .B0(n1163), .Y(P1_U3353));
  INVX1   g0131(.A(P2_DATAO_REG_1__SCAN_IN), .Y(n1165));
  NOR3X1  g0132(.A(n1153), .B(n1152), .C(n1165), .Y(n1166));
  INVX1   g0133(.A(SI_1_), .Y(n1167));
  INVX1   g0134(.A(P1_DATAO_REG_1__SCAN_IN), .Y(n1168));
  OAI21X1 g0135(.A0(n1153), .A1(n1152), .B0(P2_DATAO_REG_1__SCAN_IN), .Y(n1169));
  OAI21X1 g0136(.A0(n1149), .A1(n1168), .B0(n1169), .Y(n1170));
  NOR2X1  g0137(.A(n1158), .B(n1155), .Y(n1171));
  XOR2X1  g0138(.A(n1171), .B(n1170), .Y(n1172));
  NAND2X1 g0139(.A(n1172), .B(n1167), .Y(n1173));
  INVX1   g0140(.A(P1_DATAO_REG_0__SCAN_IN), .Y(n1174));
  OAI21X1 g0141(.A0(n1153), .A1(n1152), .B0(P2_DATAO_REG_0__SCAN_IN), .Y(n1175));
  OAI21X1 g0142(.A0(n1149), .A1(n1174), .B0(n1175), .Y(n1176));
  NOR2X1  g0143(.A(n1155), .B(n1167), .Y(n1177));
  NAND3X1 g0144(.A(n1177), .B(n1170), .C(n1176), .Y(n1178));
  NOR2X1  g0145(.A(n1170), .B(n1167), .Y(n1179));
  OAI21X1 g0146(.A0(n1158), .A1(n1155), .B0(n1179), .Y(n1180));
  NAND3X1 g0147(.A(n1180), .B(n1178), .C(n1173), .Y(n1181));
  AOI21X1 g0148(.A0(n1181), .A1(n1149), .B0(n1166), .Y(n1182));
  INVX1   g0149(.A(P1_IR_REG_31__SCAN_IN), .Y(n1183));
  NOR2X1  g0150(.A(P1_U3084), .B(n1183), .Y(n1184));
  XOR2X1  g0151(.A(P1_IR_REG_1__SCAN_IN), .B(P1_IR_REG_0__SCAN_IN), .Y(n1185));
  AOI22X1 g0152(.A0(n1184), .A1(n1185), .B0(n1162), .B1(P1_IR_REG_1__SCAN_IN), .Y(n1186));
  OAI21X1 g0153(.A0(n1182), .A1(P1_STATE_REG_SCAN_IN), .B0(n1186), .Y(P1_U3352));
  INVX1   g0154(.A(P2_DATAO_REG_2__SCAN_IN), .Y(n1188));
  NOR3X1  g0155(.A(n1153), .B(n1152), .C(n1188), .Y(n1189));
  NAND3X1 g0156(.A(n1170), .B(n1176), .C(SI_0_), .Y(n1190));
  AOI22X1 g0157(.A0(n1170), .A1(SI_1_), .B0(n1176), .B1(n1177), .Y(n1191));
  NAND2X1 g0158(.A(n1191), .B(n1190), .Y(n1192));
  INVX1   g0159(.A(SI_2_), .Y(n1193));
  AOI21X1 g0160(.A0(n1148), .A1(n1146), .B0(n1188), .Y(n1194));
  AOI21X1 g0161(.A0(n1156), .A1(P1_DATAO_REG_2__SCAN_IN), .B0(n1194), .Y(n1195));
  XOR2X1  g0162(.A(n1195), .B(n1193), .Y(n1196));
  XOR2X1  g0163(.A(n1196), .B(n1192), .Y(n1197));
  AOI21X1 g0164(.A0(n1197), .A1(n1149), .B0(n1189), .Y(n1198));
  INVX1   g0165(.A(P1_IR_REG_2__SCAN_IN), .Y(n1199));
  NOR2X1  g0166(.A(P1_IR_REG_1__SCAN_IN), .B(P1_IR_REG_0__SCAN_IN), .Y(n1200));
  XOR2X1  g0167(.A(n1200), .B(n1199), .Y(n1201));
  AOI22X1 g0168(.A0(n1184), .A1(n1201), .B0(n1162), .B1(P1_IR_REG_2__SCAN_IN), .Y(n1202));
  OAI21X1 g0169(.A0(n1198), .A1(P1_STATE_REG_SCAN_IN), .B0(n1202), .Y(P1_U3351));
  INVX1   g0170(.A(P2_DATAO_REG_3__SCAN_IN), .Y(n1204));
  NOR3X1  g0171(.A(n1153), .B(n1152), .C(n1204), .Y(n1205));
  NOR2X1  g0172(.A(n1195), .B(n1193), .Y(n1206));
  AOI22X1 g0173(.A0(n1191), .A1(n1190), .B0(n1193), .B1(n1195), .Y(n1207));
  NOR2X1  g0174(.A(n1207), .B(n1206), .Y(n1208));
  AOI21X1 g0175(.A0(n1148), .A1(n1146), .B0(n1204), .Y(n1209));
  AOI21X1 g0176(.A0(n1156), .A1(P1_DATAO_REG_3__SCAN_IN), .B0(n1209), .Y(n1210));
  XOR2X1  g0177(.A(n1210), .B(SI_3_), .Y(n1211));
  XOR2X1  g0178(.A(n1211), .B(n1208), .Y(n1212));
  AOI21X1 g0179(.A0(n1212), .A1(n1149), .B0(n1205), .Y(n1213));
  INVX1   g0180(.A(P1_IR_REG_3__SCAN_IN), .Y(n1214));
  NOR3X1  g0181(.A(P1_IR_REG_2__SCAN_IN), .B(P1_IR_REG_1__SCAN_IN), .C(P1_IR_REG_0__SCAN_IN), .Y(n1215));
  XOR2X1  g0182(.A(n1215), .B(n1214), .Y(n1216));
  AOI22X1 g0183(.A0(n1184), .A1(n1216), .B0(n1162), .B1(P1_IR_REG_3__SCAN_IN), .Y(n1217));
  OAI21X1 g0184(.A0(n1213), .A1(P1_STATE_REG_SCAN_IN), .B0(n1217), .Y(P1_U3350));
  INVX1   g0185(.A(P2_DATAO_REG_4__SCAN_IN), .Y(n1219));
  NOR3X1  g0186(.A(n1153), .B(n1152), .C(n1219), .Y(n1220));
  INVX1   g0187(.A(P1_DATAO_REG_2__SCAN_IN), .Y(n1221));
  OAI21X1 g0188(.A0(n1153), .A1(n1152), .B0(P2_DATAO_REG_2__SCAN_IN), .Y(n1222));
  OAI21X1 g0189(.A0(n1149), .A1(n1221), .B0(n1222), .Y(n1223));
  INVX1   g0190(.A(P1_DATAO_REG_3__SCAN_IN), .Y(n1224));
  OAI21X1 g0191(.A0(n1153), .A1(n1152), .B0(P2_DATAO_REG_3__SCAN_IN), .Y(n1225));
  OAI21X1 g0192(.A0(n1149), .A1(n1224), .B0(n1225), .Y(n1226));
  OAI22X1 g0193(.A0(n1223), .A1(SI_2_), .B0(SI_3_), .B1(n1226), .Y(n1227));
  AOI21X1 g0194(.A0(n1191), .A1(n1190), .B0(n1227), .Y(n1228));
  NAND2X1 g0195(.A(n1223), .B(SI_2_), .Y(n1229));
  NOR2X1  g0196(.A(n1226), .B(SI_3_), .Y(n1230));
  NAND2X1 g0197(.A(n1226), .B(SI_3_), .Y(n1231));
  OAI21X1 g0198(.A0(n1230), .A1(n1229), .B0(n1231), .Y(n1232));
  NOR2X1  g0199(.A(n1232), .B(n1228), .Y(n1233));
  INVX1   g0200(.A(P1_DATAO_REG_4__SCAN_IN), .Y(n1234));
  NOR3X1  g0201(.A(n1153), .B(n1152), .C(n1234), .Y(n1235));
  AOI21X1 g0202(.A0(n1148), .A1(n1146), .B0(n1219), .Y(n1236));
  NOR2X1  g0203(.A(n1236), .B(n1235), .Y(n1237));
  XOR2X1  g0204(.A(n1237), .B(SI_4_), .Y(n1238));
  XOR2X1  g0205(.A(n1238), .B(n1233), .Y(n1239));
  AOI21X1 g0206(.A0(n1239), .A1(n1149), .B0(n1220), .Y(n1240));
  NAND2X1 g0207(.A(n1215), .B(n1214), .Y(n1241));
  NOR2X1  g0208(.A(P1_IR_REG_4__SCAN_IN), .B(P1_IR_REG_3__SCAN_IN), .Y(n1242));
  AOI22X1 g0209(.A0(n1241), .A1(P1_IR_REG_4__SCAN_IN), .B0(n1215), .B1(n1242), .Y(n1243));
  AOI22X1 g0210(.A0(n1184), .A1(n1243), .B0(n1162), .B1(P1_IR_REG_4__SCAN_IN), .Y(n1244));
  OAI21X1 g0211(.A0(n1240), .A1(P1_STATE_REG_SCAN_IN), .B0(n1244), .Y(P1_U3349));
  INVX1   g0212(.A(P2_DATAO_REG_5__SCAN_IN), .Y(n1246));
  NOR3X1  g0213(.A(n1153), .B(n1152), .C(n1246), .Y(n1247));
  NOR3X1  g0214(.A(n1236), .B(n1235), .C(SI_4_), .Y(n1248));
  OAI21X1 g0215(.A0(n1236), .A1(n1235), .B0(SI_4_), .Y(n1249));
  OAI21X1 g0216(.A0(n1248), .A1(n1233), .B0(n1249), .Y(n1250));
  INVX1   g0217(.A(SI_5_), .Y(n1251));
  INVX1   g0218(.A(P1_DATAO_REG_5__SCAN_IN), .Y(n1252));
  NOR3X1  g0219(.A(n1153), .B(n1152), .C(n1252), .Y(n1253));
  AOI21X1 g0220(.A0(n1148), .A1(n1146), .B0(n1246), .Y(n1254));
  NOR2X1  g0221(.A(n1254), .B(n1253), .Y(n1255));
  XOR2X1  g0222(.A(n1255), .B(n1251), .Y(n1256));
  XOR2X1  g0223(.A(n1256), .B(n1250), .Y(n1257));
  AOI21X1 g0224(.A0(n1257), .A1(n1149), .B0(n1247), .Y(n1258));
  INVX1   g0225(.A(P1_IR_REG_4__SCAN_IN), .Y(n1259));
  NAND3X1 g0226(.A(n1215), .B(n1259), .C(n1214), .Y(n1260));
  XOR2X1  g0227(.A(n1260), .B(P1_IR_REG_5__SCAN_IN), .Y(n1261));
  AOI22X1 g0228(.A0(n1184), .A1(n1261), .B0(n1162), .B1(P1_IR_REG_5__SCAN_IN), .Y(n1262));
  OAI21X1 g0229(.A0(n1258), .A1(P1_STATE_REG_SCAN_IN), .B0(n1262), .Y(P1_U3348));
  INVX1   g0230(.A(P2_DATAO_REG_6__SCAN_IN), .Y(n1264));
  NOR3X1  g0231(.A(n1153), .B(n1152), .C(n1264), .Y(n1265));
  AOI21X1 g0232(.A0(n1148), .A1(n1146), .B0(n1165), .Y(n1266));
  AOI21X1 g0233(.A0(n1156), .A1(P1_DATAO_REG_1__SCAN_IN), .B0(n1266), .Y(n1267));
  NOR3X1  g0234(.A(n1267), .B(n1158), .C(n1155), .Y(n1268));
  INVX1   g0235(.A(n1177), .Y(n1269));
  OAI22X1 g0236(.A0(n1267), .A1(n1167), .B0(n1158), .B1(n1269), .Y(n1270));
  INVX1   g0237(.A(SI_3_), .Y(n1271));
  AOI22X1 g0238(.A0(n1195), .A1(n1193), .B0(n1271), .B1(n1210), .Y(n1272));
  OAI21X1 g0239(.A0(n1270), .A1(n1268), .B0(n1272), .Y(n1273));
  NAND2X1 g0240(.A(n1210), .B(n1271), .Y(n1274));
  NOR2X1  g0241(.A(n1210), .B(n1271), .Y(n1275));
  AOI21X1 g0242(.A0(n1274), .A1(n1206), .B0(n1275), .Y(n1276));
  NAND2X1 g0243(.A(n1276), .B(n1273), .Y(n1277));
  NOR3X1  g0244(.A(n1254), .B(n1253), .C(SI_5_), .Y(n1278));
  OAI21X1 g0245(.A0(n1254), .A1(n1253), .B0(SI_5_), .Y(n1279));
  OAI21X1 g0246(.A0(n1278), .A1(n1249), .B0(n1279), .Y(n1280));
  NOR2X1  g0247(.A(n1278), .B(n1248), .Y(n1281));
  AOI21X1 g0248(.A0(n1281), .A1(n1277), .B0(n1280), .Y(n1282));
  INVX1   g0249(.A(P1_DATAO_REG_6__SCAN_IN), .Y(n1283));
  NOR3X1  g0250(.A(n1153), .B(n1152), .C(n1283), .Y(n1284));
  AOI21X1 g0251(.A0(n1148), .A1(n1146), .B0(n1264), .Y(n1285));
  NOR2X1  g0252(.A(n1285), .B(n1284), .Y(n1286));
  XOR2X1  g0253(.A(n1286), .B(SI_6_), .Y(n1287));
  XOR2X1  g0254(.A(n1287), .B(n1282), .Y(n1288));
  AOI21X1 g0255(.A0(n1288), .A1(n1149), .B0(n1265), .Y(n1289));
  INVX1   g0256(.A(P1_IR_REG_5__SCAN_IN), .Y(n1290));
  NAND3X1 g0257(.A(n1242), .B(n1215), .C(n1290), .Y(n1291));
  INVX1   g0258(.A(P1_IR_REG_6__SCAN_IN), .Y(n1292));
  NAND2X1 g0259(.A(n1292), .B(n1290), .Y(n1293));
  NOR2X1  g0260(.A(n1293), .B(n1260), .Y(n1294));
  AOI21X1 g0261(.A0(n1291), .A1(P1_IR_REG_6__SCAN_IN), .B0(n1294), .Y(n1295));
  AOI22X1 g0262(.A0(n1184), .A1(n1295), .B0(n1162), .B1(P1_IR_REG_6__SCAN_IN), .Y(n1296));
  OAI21X1 g0263(.A0(n1289), .A1(P1_STATE_REG_SCAN_IN), .B0(n1296), .Y(P1_U3347));
  INVX1   g0264(.A(P2_DATAO_REG_7__SCAN_IN), .Y(n1298));
  NOR3X1  g0265(.A(n1153), .B(n1152), .C(n1298), .Y(n1299));
  NOR3X1  g0266(.A(n1285), .B(n1284), .C(SI_6_), .Y(n1300));
  NOR3X1  g0267(.A(n1300), .B(n1278), .C(n1248), .Y(n1301));
  OAI21X1 g0268(.A0(n1232), .A1(n1228), .B0(n1301), .Y(n1302));
  INVX1   g0269(.A(SI_6_), .Y(n1303));
  NAND3X1 g0270(.A(n1148), .B(n1146), .C(P1_DATAO_REG_6__SCAN_IN), .Y(n1304));
  OAI21X1 g0271(.A0(n1153), .A1(n1152), .B0(P2_DATAO_REG_6__SCAN_IN), .Y(n1305));
  NAND3X1 g0272(.A(n1305), .B(n1304), .C(n1303), .Y(n1306));
  AOI21X1 g0273(.A0(n1305), .A1(n1304), .B0(n1303), .Y(n1307));
  AOI21X1 g0274(.A0(n1306), .A1(n1280), .B0(n1307), .Y(n1308));
  NAND2X1 g0275(.A(n1308), .B(n1302), .Y(n1309));
  INVX1   g0276(.A(SI_7_), .Y(n1310));
  INVX1   g0277(.A(P1_DATAO_REG_7__SCAN_IN), .Y(n1311));
  NOR3X1  g0278(.A(n1153), .B(n1152), .C(n1311), .Y(n1312));
  AOI21X1 g0279(.A0(n1148), .A1(n1146), .B0(n1298), .Y(n1313));
  NOR2X1  g0280(.A(n1313), .B(n1312), .Y(n1314));
  XOR2X1  g0281(.A(n1314), .B(n1310), .Y(n1315));
  XOR2X1  g0282(.A(n1315), .B(n1309), .Y(n1316));
  AOI21X1 g0283(.A0(n1316), .A1(n1149), .B0(n1299), .Y(n1317));
  INVX1   g0284(.A(P1_IR_REG_7__SCAN_IN), .Y(n1318));
  XOR2X1  g0285(.A(n1294), .B(n1318), .Y(n1319));
  AOI22X1 g0286(.A0(n1184), .A1(n1319), .B0(n1162), .B1(P1_IR_REG_7__SCAN_IN), .Y(n1320));
  OAI21X1 g0287(.A0(n1317), .A1(P1_STATE_REG_SCAN_IN), .B0(n1320), .Y(P1_U3346));
  INVX1   g0288(.A(P2_DATAO_REG_8__SCAN_IN), .Y(n1322));
  NOR3X1  g0289(.A(n1153), .B(n1152), .C(n1322), .Y(n1323));
  NAND2X1 g0290(.A(n1306), .B(n1281), .Y(n1324));
  AOI21X1 g0291(.A0(n1276), .A1(n1273), .B0(n1324), .Y(n1325));
  NAND2X1 g0292(.A(n1306), .B(n1280), .Y(n1326));
  OAI21X1 g0293(.A0(n1286), .A1(n1303), .B0(n1326), .Y(n1327));
  NAND3X1 g0294(.A(n1148), .B(n1146), .C(P1_DATAO_REG_7__SCAN_IN), .Y(n1328));
  OAI21X1 g0295(.A0(n1153), .A1(n1152), .B0(P2_DATAO_REG_7__SCAN_IN), .Y(n1329));
  NAND2X1 g0296(.A(n1329), .B(n1328), .Y(n1330));
  OAI22X1 g0297(.A0(n1327), .A1(n1325), .B0(SI_7_), .B1(n1330), .Y(n1331));
  OAI21X1 g0298(.A0(n1314), .A1(n1310), .B0(n1331), .Y(n1332));
  INVX1   g0299(.A(SI_8_), .Y(n1333));
  AOI21X1 g0300(.A0(n1148), .A1(n1146), .B0(n1322), .Y(n1334));
  AOI21X1 g0301(.A0(n1156), .A1(P1_DATAO_REG_8__SCAN_IN), .B0(n1334), .Y(n1335));
  XOR2X1  g0302(.A(n1335), .B(n1333), .Y(n1336));
  XOR2X1  g0303(.A(n1336), .B(n1332), .Y(n1337));
  AOI21X1 g0304(.A0(n1337), .A1(n1149), .B0(n1323), .Y(n1338));
  NOR2X1  g0305(.A(P1_IR_REG_6__SCAN_IN), .B(P1_IR_REG_5__SCAN_IN), .Y(n1339));
  NAND4X1 g0306(.A(n1242), .B(n1215), .C(n1318), .D(n1339), .Y(n1340));
  INVX1   g0307(.A(P1_IR_REG_8__SCAN_IN), .Y(n1341));
  NOR4X1  g0308(.A(P1_IR_REG_5__SCAN_IN), .B(P1_IR_REG_4__SCAN_IN), .C(P1_IR_REG_3__SCAN_IN), .D(P1_IR_REG_6__SCAN_IN), .Y(n1342));
  NAND4X1 g0309(.A(n1215), .B(n1341), .C(n1318), .D(n1342), .Y(n1343));
  INVX1   g0310(.A(n1343), .Y(n1344));
  AOI21X1 g0311(.A0(n1340), .A1(P1_IR_REG_8__SCAN_IN), .B0(n1344), .Y(n1345));
  AOI22X1 g0312(.A0(n1184), .A1(n1345), .B0(n1162), .B1(P1_IR_REG_8__SCAN_IN), .Y(n1346));
  OAI21X1 g0313(.A0(n1338), .A1(P1_STATE_REG_SCAN_IN), .B0(n1346), .Y(P1_U3345));
  INVX1   g0314(.A(P2_DATAO_REG_9__SCAN_IN), .Y(n1348));
  NOR3X1  g0315(.A(n1153), .B(n1152), .C(n1348), .Y(n1349));
  AOI21X1 g0316(.A0(n1329), .A1(n1328), .B0(n1310), .Y(n1350));
  NAND3X1 g0317(.A(n1148), .B(n1146), .C(P1_DATAO_REG_8__SCAN_IN), .Y(n1351));
  OAI21X1 g0318(.A0(n1153), .A1(n1152), .B0(P2_DATAO_REG_8__SCAN_IN), .Y(n1352));
  NAND3X1 g0319(.A(n1352), .B(n1351), .C(n1333), .Y(n1353));
  AOI21X1 g0320(.A0(n1352), .A1(n1351), .B0(n1333), .Y(n1354));
  AOI21X1 g0321(.A0(n1353), .A1(n1350), .B0(n1354), .Y(n1355));
  INVX1   g0322(.A(n1355), .Y(n1356));
  AOI22X1 g0323(.A0(n1314), .A1(n1310), .B0(n1333), .B1(n1335), .Y(n1357));
  AOI21X1 g0324(.A0(n1357), .A1(n1309), .B0(n1356), .Y(n1358));
  AOI21X1 g0325(.A0(n1148), .A1(n1146), .B0(n1348), .Y(n1359));
  AOI21X1 g0326(.A0(n1156), .A1(P1_DATAO_REG_9__SCAN_IN), .B0(n1359), .Y(n1360));
  XOR2X1  g0327(.A(n1360), .B(SI_9_), .Y(n1361));
  XOR2X1  g0328(.A(n1361), .B(n1358), .Y(n1362));
  AOI21X1 g0329(.A0(n1362), .A1(n1149), .B0(n1349), .Y(n1363));
  XOR2X1  g0330(.A(n1343), .B(P1_IR_REG_9__SCAN_IN), .Y(n1364));
  AOI22X1 g0331(.A0(n1184), .A1(n1364), .B0(n1162), .B1(P1_IR_REG_9__SCAN_IN), .Y(n1365));
  OAI21X1 g0332(.A0(n1363), .A1(P1_STATE_REG_SCAN_IN), .B0(n1365), .Y(P1_U3344));
  INVX1   g0333(.A(P2_DATAO_REG_10__SCAN_IN), .Y(n1367));
  NOR3X1  g0334(.A(n1153), .B(n1152), .C(n1367), .Y(n1368));
  INVX1   g0335(.A(P1_DATAO_REG_9__SCAN_IN), .Y(n1369));
  OAI21X1 g0336(.A0(n1153), .A1(n1152), .B0(P2_DATAO_REG_9__SCAN_IN), .Y(n1370));
  OAI21X1 g0337(.A0(n1149), .A1(n1369), .B0(n1370), .Y(n1371));
  NOR2X1  g0338(.A(n1371), .B(SI_9_), .Y(n1372));
  NAND2X1 g0339(.A(n1371), .B(SI_9_), .Y(n1373));
  OAI21X1 g0340(.A0(n1372), .A1(n1355), .B0(n1373), .Y(n1374));
  OAI21X1 g0341(.A0(n1330), .A1(SI_7_), .B0(n1353), .Y(n1375));
  NOR2X1  g0342(.A(n1372), .B(n1375), .Y(n1376));
  AOI21X1 g0343(.A0(n1376), .A1(n1309), .B0(n1374), .Y(n1377));
  AOI21X1 g0344(.A0(n1148), .A1(n1146), .B0(n1367), .Y(n1378));
  AOI21X1 g0345(.A0(n1156), .A1(P1_DATAO_REG_10__SCAN_IN), .B0(n1378), .Y(n1379));
  XOR2X1  g0346(.A(n1379), .B(SI_10_), .Y(n1380));
  XOR2X1  g0347(.A(n1380), .B(n1377), .Y(n1381));
  AOI21X1 g0348(.A0(n1381), .A1(n1149), .B0(n1368), .Y(n1382));
  INVX1   g0349(.A(P1_IR_REG_9__SCAN_IN), .Y(n1383));
  INVX1   g0350(.A(P1_IR_REG_10__SCAN_IN), .Y(n1384));
  AOI21X1 g0351(.A0(n1344), .A1(n1383), .B0(n1384), .Y(n1385));
  NOR2X1  g0352(.A(P1_IR_REG_10__SCAN_IN), .B(P1_IR_REG_9__SCAN_IN), .Y(n1386));
  INVX1   g0353(.A(n1386), .Y(n1387));
  NOR2X1  g0354(.A(n1387), .B(n1343), .Y(n1388));
  NOR2X1  g0355(.A(n1388), .B(n1385), .Y(n1389));
  AOI22X1 g0356(.A0(n1184), .A1(n1389), .B0(n1162), .B1(P1_IR_REG_10__SCAN_IN), .Y(n1390));
  OAI21X1 g0357(.A0(n1382), .A1(P1_STATE_REG_SCAN_IN), .B0(n1390), .Y(P1_U3343));
  INVX1   g0358(.A(P2_DATAO_REG_11__SCAN_IN), .Y(n1392));
  NOR3X1  g0359(.A(n1153), .B(n1152), .C(n1392), .Y(n1393));
  INVX1   g0360(.A(P1_DATAO_REG_10__SCAN_IN), .Y(n1394));
  NOR3X1  g0361(.A(n1153), .B(n1152), .C(n1394), .Y(n1395));
  NOR3X1  g0362(.A(n1378), .B(n1395), .C(SI_10_), .Y(n1396));
  INVX1   g0363(.A(n1396), .Y(n1397));
  NAND2X1 g0364(.A(n1397), .B(n1376), .Y(n1398));
  AOI21X1 g0365(.A0(n1308), .A1(n1302), .B0(n1398), .Y(n1399));
  INVX1   g0366(.A(SI_10_), .Y(n1400));
  NAND2X1 g0367(.A(n1397), .B(n1374), .Y(n1401));
  OAI21X1 g0368(.A0(n1379), .A1(n1400), .B0(n1401), .Y(n1402));
  NOR2X1  g0369(.A(n1402), .B(n1399), .Y(n1403));
  AOI21X1 g0370(.A0(n1148), .A1(n1146), .B0(n1392), .Y(n1404));
  AOI21X1 g0371(.A0(n1156), .A1(P1_DATAO_REG_11__SCAN_IN), .B0(n1404), .Y(n1405));
  XOR2X1  g0372(.A(n1405), .B(SI_11_), .Y(n1406));
  XOR2X1  g0373(.A(n1406), .B(n1403), .Y(n1407));
  AOI21X1 g0374(.A0(n1407), .A1(n1149), .B0(n1393), .Y(n1408));
  INVX1   g0375(.A(P1_IR_REG_11__SCAN_IN), .Y(n1409));
  XOR2X1  g0376(.A(n1388), .B(n1409), .Y(n1410));
  AOI22X1 g0377(.A0(n1184), .A1(n1410), .B0(n1162), .B1(P1_IR_REG_11__SCAN_IN), .Y(n1411));
  OAI21X1 g0378(.A0(n1408), .A1(P1_STATE_REG_SCAN_IN), .B0(n1411), .Y(P1_U3342));
  INVX1   g0379(.A(P2_DATAO_REG_12__SCAN_IN), .Y(n1413));
  NOR3X1  g0380(.A(n1153), .B(n1152), .C(n1413), .Y(n1414));
  INVX1   g0381(.A(SI_11_), .Y(n1415));
  INVX1   g0382(.A(P1_DATAO_REG_11__SCAN_IN), .Y(n1416));
  OAI21X1 g0383(.A0(n1153), .A1(n1152), .B0(P2_DATAO_REG_11__SCAN_IN), .Y(n1417));
  OAI21X1 g0384(.A0(n1149), .A1(n1416), .B0(n1417), .Y(n1418));
  OAI22X1 g0385(.A0(n1402), .A1(n1399), .B0(SI_11_), .B1(n1418), .Y(n1419));
  OAI21X1 g0386(.A0(n1405), .A1(n1415), .B0(n1419), .Y(n1420));
  INVX1   g0387(.A(SI_12_), .Y(n1421));
  AOI21X1 g0388(.A0(n1148), .A1(n1146), .B0(n1413), .Y(n1422));
  AOI21X1 g0389(.A0(n1156), .A1(P1_DATAO_REG_12__SCAN_IN), .B0(n1422), .Y(n1423));
  XOR2X1  g0390(.A(n1423), .B(n1421), .Y(n1424));
  XOR2X1  g0391(.A(n1424), .B(n1420), .Y(n1425));
  AOI21X1 g0392(.A0(n1425), .A1(n1149), .B0(n1414), .Y(n1426));
  INVX1   g0393(.A(P1_IR_REG_12__SCAN_IN), .Y(n1427));
  AOI21X1 g0394(.A0(n1388), .A1(n1409), .B0(n1427), .Y(n1428));
  NOR4X1  g0395(.A(n1343), .B(P1_IR_REG_12__SCAN_IN), .C(P1_IR_REG_11__SCAN_IN), .D(n1387), .Y(n1429));
  NOR2X1  g0396(.A(n1429), .B(n1428), .Y(n1430));
  AOI22X1 g0397(.A0(n1184), .A1(n1430), .B0(n1162), .B1(P1_IR_REG_12__SCAN_IN), .Y(n1431));
  OAI21X1 g0398(.A0(n1426), .A1(P1_STATE_REG_SCAN_IN), .B0(n1431), .Y(P1_U3341));
  INVX1   g0399(.A(P2_DATAO_REG_13__SCAN_IN), .Y(n1433));
  NOR3X1  g0400(.A(n1153), .B(n1152), .C(n1433), .Y(n1434));
  NOR2X1  g0401(.A(n1405), .B(n1415), .Y(n1435));
  NAND2X1 g0402(.A(n1423), .B(n1421), .Y(n1436));
  NOR2X1  g0403(.A(n1423), .B(n1421), .Y(n1437));
  AOI21X1 g0404(.A0(n1436), .A1(n1435), .B0(n1437), .Y(n1438));
  OAI21X1 g0405(.A0(n1418), .A1(SI_11_), .B0(n1436), .Y(n1439));
  OAI21X1 g0406(.A0(n1439), .A1(n1403), .B0(n1438), .Y(n1440));
  INVX1   g0407(.A(P1_DATAO_REG_13__SCAN_IN), .Y(n1441));
  OAI21X1 g0408(.A0(n1153), .A1(n1152), .B0(P2_DATAO_REG_13__SCAN_IN), .Y(n1442));
  OAI21X1 g0409(.A0(n1149), .A1(n1441), .B0(n1442), .Y(n1443));
  XOR2X1  g0410(.A(n1443), .B(SI_13_), .Y(n1444));
  XOR2X1  g0411(.A(n1444), .B(n1440), .Y(n1445));
  AOI21X1 g0412(.A0(n1445), .A1(n1149), .B0(n1434), .Y(n1446));
  INVX1   g0413(.A(P1_IR_REG_13__SCAN_IN), .Y(n1447));
  XOR2X1  g0414(.A(n1429), .B(n1447), .Y(n1448));
  AOI22X1 g0415(.A0(n1184), .A1(n1448), .B0(n1162), .B1(P1_IR_REG_13__SCAN_IN), .Y(n1449));
  OAI21X1 g0416(.A0(n1446), .A1(P1_STATE_REG_SCAN_IN), .B0(n1449), .Y(P1_U3340));
  INVX1   g0417(.A(P2_DATAO_REG_14__SCAN_IN), .Y(n1451));
  NOR3X1  g0418(.A(n1153), .B(n1152), .C(n1451), .Y(n1452));
  NOR2X1  g0419(.A(n1443), .B(SI_13_), .Y(n1453));
  NOR2X1  g0420(.A(n1453), .B(n1438), .Y(n1454));
  AOI21X1 g0421(.A0(n1443), .A1(SI_13_), .B0(n1454), .Y(n1455));
  AOI22X1 g0422(.A0(n1405), .A1(n1415), .B0(n1421), .B1(n1423), .Y(n1456));
  OAI21X1 g0423(.A0(n1443), .A1(SI_13_), .B0(n1456), .Y(n1457));
  OAI21X1 g0424(.A0(n1457), .A1(n1403), .B0(n1455), .Y(n1458));
  INVX1   g0425(.A(SI_14_), .Y(n1459));
  AOI21X1 g0426(.A0(n1148), .A1(n1146), .B0(n1451), .Y(n1460));
  AOI21X1 g0427(.A0(n1156), .A1(P1_DATAO_REG_14__SCAN_IN), .B0(n1460), .Y(n1461));
  XOR2X1  g0428(.A(n1461), .B(n1459), .Y(n1462));
  XOR2X1  g0429(.A(n1462), .B(n1458), .Y(n1463));
  AOI21X1 g0430(.A0(n1463), .A1(n1149), .B0(n1452), .Y(n1464));
  INVX1   g0431(.A(P1_IR_REG_14__SCAN_IN), .Y(n1465));
  AOI21X1 g0432(.A0(n1429), .A1(n1447), .B0(n1465), .Y(n1466));
  INVX1   g0433(.A(n1429), .Y(n1467));
  NOR3X1  g0434(.A(n1467), .B(P1_IR_REG_14__SCAN_IN), .C(P1_IR_REG_13__SCAN_IN), .Y(n1468));
  NOR2X1  g0435(.A(n1468), .B(n1466), .Y(n1469));
  AOI22X1 g0436(.A0(n1184), .A1(n1469), .B0(n1162), .B1(P1_IR_REG_14__SCAN_IN), .Y(n1470));
  OAI21X1 g0437(.A0(n1464), .A1(P1_STATE_REG_SCAN_IN), .B0(n1470), .Y(P1_U3339));
  INVX1   g0438(.A(P2_DATAO_REG_15__SCAN_IN), .Y(n1472));
  NOR3X1  g0439(.A(n1153), .B(n1152), .C(n1472), .Y(n1473));
  NOR3X1  g0440(.A(n1396), .B(n1372), .C(n1375), .Y(n1474));
  OAI21X1 g0441(.A0(n1327), .A1(n1325), .B0(n1474), .Y(n1475));
  NOR2X1  g0442(.A(n1379), .B(n1400), .Y(n1476));
  AOI21X1 g0443(.A0(n1397), .A1(n1374), .B0(n1476), .Y(n1477));
  NOR2X1  g0444(.A(n1453), .B(n1439), .Y(n1478));
  NAND2X1 g0445(.A(n1461), .B(n1459), .Y(n1479));
  NAND2X1 g0446(.A(n1479), .B(n1478), .Y(n1480));
  AOI21X1 g0447(.A0(n1477), .A1(n1475), .B0(n1480), .Y(n1481));
  INVX1   g0448(.A(n1479), .Y(n1482));
  NOR2X1  g0449(.A(n1461), .B(n1459), .Y(n1483));
  INVX1   g0450(.A(n1483), .Y(n1484));
  OAI21X1 g0451(.A0(n1482), .A1(n1455), .B0(n1484), .Y(n1485));
  NOR2X1  g0452(.A(n1485), .B(n1481), .Y(n1486));
  AOI21X1 g0453(.A0(n1148), .A1(n1146), .B0(n1472), .Y(n1487));
  AOI21X1 g0454(.A0(n1156), .A1(P1_DATAO_REG_15__SCAN_IN), .B0(n1487), .Y(n1488));
  XOR2X1  g0455(.A(n1488), .B(SI_15_), .Y(n1489));
  XOR2X1  g0456(.A(n1489), .B(n1486), .Y(n1490));
  AOI21X1 g0457(.A0(n1490), .A1(n1149), .B0(n1473), .Y(n1491));
  INVX1   g0458(.A(P1_IR_REG_15__SCAN_IN), .Y(n1492));
  XOR2X1  g0459(.A(n1468), .B(n1492), .Y(n1493));
  AOI22X1 g0460(.A0(n1184), .A1(n1493), .B0(n1162), .B1(P1_IR_REG_15__SCAN_IN), .Y(n1494));
  OAI21X1 g0461(.A0(n1491), .A1(P1_STATE_REG_SCAN_IN), .B0(n1494), .Y(P1_U3338));
  INVX1   g0462(.A(P2_DATAO_REG_16__SCAN_IN), .Y(n1496));
  NOR3X1  g0463(.A(n1153), .B(n1152), .C(n1496), .Y(n1497));
  INVX1   g0464(.A(SI_15_), .Y(n1498));
  NOR2X1  g0465(.A(n1488), .B(n1498), .Y(n1499));
  NOR2X1  g0466(.A(n1482), .B(n1457), .Y(n1500));
  OAI21X1 g0467(.A0(n1402), .A1(n1399), .B0(n1500), .Y(n1501));
  NAND2X1 g0468(.A(n1443), .B(SI_13_), .Y(n1502));
  OAI21X1 g0469(.A0(n1453), .A1(n1438), .B0(n1502), .Y(n1503));
  AOI21X1 g0470(.A0(n1479), .A1(n1503), .B0(n1483), .Y(n1504));
  AOI22X1 g0471(.A0(n1504), .A1(n1501), .B0(n1498), .B1(n1488), .Y(n1505));
  NOR2X1  g0472(.A(n1505), .B(n1499), .Y(n1506));
  AOI21X1 g0473(.A0(n1148), .A1(n1146), .B0(n1496), .Y(n1507));
  AOI21X1 g0474(.A0(n1156), .A1(P1_DATAO_REG_16__SCAN_IN), .B0(n1507), .Y(n1508));
  XOR2X1  g0475(.A(n1508), .B(SI_16_), .Y(n1509));
  XOR2X1  g0476(.A(n1509), .B(n1506), .Y(n1510));
  AOI21X1 g0477(.A0(n1510), .A1(n1149), .B0(n1497), .Y(n1511));
  INVX1   g0478(.A(P1_IR_REG_16__SCAN_IN), .Y(n1512));
  NOR4X1  g0479(.A(P1_IR_REG_15__SCAN_IN), .B(P1_IR_REG_14__SCAN_IN), .C(P1_IR_REG_13__SCAN_IN), .D(n1467), .Y(n1513));
  NOR4X1  g0480(.A(P1_IR_REG_12__SCAN_IN), .B(P1_IR_REG_11__SCAN_IN), .C(P1_IR_REG_10__SCAN_IN), .D(P1_IR_REG_13__SCAN_IN), .Y(n1514));
  NAND2X1 g0481(.A(n1514), .B(n1465), .Y(n1515));
  NOR2X1  g0482(.A(P1_IR_REG_16__SCAN_IN), .B(P1_IR_REG_15__SCAN_IN), .Y(n1516));
  NAND3X1 g0483(.A(n1516), .B(n1200), .C(n1290), .Y(n1517));
  NOR4X1  g0484(.A(P1_IR_REG_8__SCAN_IN), .B(P1_IR_REG_7__SCAN_IN), .C(P1_IR_REG_6__SCAN_IN), .D(P1_IR_REG_9__SCAN_IN), .Y(n1518));
  INVX1   g0485(.A(n1518), .Y(n1519));
  NOR2X1  g0486(.A(P1_IR_REG_3__SCAN_IN), .B(P1_IR_REG_2__SCAN_IN), .Y(n1520));
  NAND2X1 g0487(.A(n1520), .B(n1259), .Y(n1521));
  NOR4X1  g0488(.A(n1519), .B(n1517), .C(n1515), .D(n1521), .Y(n1522));
  INVX1   g0489(.A(n1522), .Y(n1523));
  OAI21X1 g0490(.A0(n1513), .A1(n1512), .B0(n1523), .Y(n1524));
  INVX1   g0491(.A(n1524), .Y(n1525));
  AOI22X1 g0492(.A0(n1184), .A1(n1525), .B0(n1162), .B1(P1_IR_REG_16__SCAN_IN), .Y(n1526));
  OAI21X1 g0493(.A0(n1511), .A1(P1_STATE_REG_SCAN_IN), .B0(n1526), .Y(P1_U3337));
  INVX1   g0494(.A(P2_DATAO_REG_17__SCAN_IN), .Y(n1528));
  NOR3X1  g0495(.A(n1153), .B(n1152), .C(n1528), .Y(n1529));
  INVX1   g0496(.A(SI_16_), .Y(n1530));
  NOR2X1  g0497(.A(n1508), .B(n1530), .Y(n1531));
  INVX1   g0498(.A(n1499), .Y(n1532));
  NAND2X1 g0499(.A(n1488), .B(n1498), .Y(n1533));
  OAI21X1 g0500(.A0(n1485), .A1(n1481), .B0(n1533), .Y(n1534));
  AOI22X1 g0501(.A0(n1534), .A1(n1532), .B0(n1530), .B1(n1508), .Y(n1535));
  NOR2X1  g0502(.A(n1535), .B(n1531), .Y(n1536));
  AOI21X1 g0503(.A0(n1148), .A1(n1146), .B0(n1528), .Y(n1537));
  AOI21X1 g0504(.A0(n1156), .A1(P1_DATAO_REG_17__SCAN_IN), .B0(n1537), .Y(n1538));
  XOR2X1  g0505(.A(n1538), .B(SI_17_), .Y(n1539));
  XOR2X1  g0506(.A(n1539), .B(n1536), .Y(n1540));
  AOI21X1 g0507(.A0(n1540), .A1(n1149), .B0(n1529), .Y(n1541));
  INVX1   g0508(.A(P1_IR_REG_17__SCAN_IN), .Y(n1542));
  XOR2X1  g0509(.A(n1522), .B(n1542), .Y(n1543));
  AOI22X1 g0510(.A0(n1184), .A1(n1543), .B0(n1162), .B1(P1_IR_REG_17__SCAN_IN), .Y(n1544));
  OAI21X1 g0511(.A0(n1541), .A1(P1_STATE_REG_SCAN_IN), .B0(n1544), .Y(P1_U3336));
  INVX1   g0512(.A(P2_DATAO_REG_18__SCAN_IN), .Y(n1546));
  NOR3X1  g0513(.A(n1153), .B(n1152), .C(n1546), .Y(n1547));
  INVX1   g0514(.A(SI_17_), .Y(n1548));
  NOR2X1  g0515(.A(n1538), .B(n1548), .Y(n1549));
  INVX1   g0516(.A(n1531), .Y(n1550));
  INVX1   g0517(.A(n1508), .Y(n1551));
  OAI22X1 g0518(.A0(n1505), .A1(n1499), .B0(SI_16_), .B1(n1551), .Y(n1552));
  AOI22X1 g0519(.A0(n1552), .A1(n1550), .B0(n1548), .B1(n1538), .Y(n1553));
  NOR2X1  g0520(.A(n1553), .B(n1549), .Y(n1554));
  AOI21X1 g0521(.A0(n1148), .A1(n1146), .B0(n1546), .Y(n1555));
  AOI21X1 g0522(.A0(n1156), .A1(P1_DATAO_REG_18__SCAN_IN), .B0(n1555), .Y(n1556));
  XOR2X1  g0523(.A(n1556), .B(SI_18_), .Y(n1557));
  XOR2X1  g0524(.A(n1557), .B(n1554), .Y(n1558));
  AOI21X1 g0525(.A0(n1558), .A1(n1149), .B0(n1547), .Y(n1559));
  OAI21X1 g0526(.A0(n1523), .A1(P1_IR_REG_17__SCAN_IN), .B0(P1_IR_REG_18__SCAN_IN), .Y(n1560));
  NOR3X1  g0527(.A(P1_IR_REG_12__SCAN_IN), .B(P1_IR_REG_11__SCAN_IN), .C(P1_IR_REG_10__SCAN_IN), .Y(n1561));
  NAND2X1 g0528(.A(n1561), .B(n1447), .Y(n1562));
  NOR2X1  g0529(.A(n1562), .B(P1_IR_REG_14__SCAN_IN), .Y(n1563));
  INVX1   g0530(.A(P1_IR_REG_1__SCAN_IN), .Y(n1564));
  INVX1   g0531(.A(P1_IR_REG_18__SCAN_IN), .Y(n1565));
  NAND4X1 g0532(.A(n1542), .B(n1290), .C(n1564), .D(n1565), .Y(n1566));
  NOR3X1  g0533(.A(n1566), .B(P1_IR_REG_16__SCAN_IN), .C(P1_IR_REG_15__SCAN_IN), .Y(n1567));
  NOR4X1  g0534(.A(P1_IR_REG_3__SCAN_IN), .B(P1_IR_REG_2__SCAN_IN), .C(P1_IR_REG_0__SCAN_IN), .D(P1_IR_REG_4__SCAN_IN), .Y(n1568));
  NAND4X1 g0535(.A(n1567), .B(n1518), .C(n1563), .D(n1568), .Y(n1569));
  NAND2X1 g0536(.A(n1569), .B(n1560), .Y(n1570));
  INVX1   g0537(.A(n1570), .Y(n1571));
  AOI22X1 g0538(.A0(n1184), .A1(n1571), .B0(n1162), .B1(P1_IR_REG_18__SCAN_IN), .Y(n1572));
  OAI21X1 g0539(.A0(n1559), .A1(P1_STATE_REG_SCAN_IN), .B0(n1572), .Y(P1_U3335));
  INVX1   g0540(.A(P2_DATAO_REG_19__SCAN_IN), .Y(n1574));
  NOR3X1  g0541(.A(n1153), .B(n1152), .C(n1574), .Y(n1575));
  INVX1   g0542(.A(SI_18_), .Y(n1576));
  NOR2X1  g0543(.A(n1556), .B(n1576), .Y(n1577));
  INVX1   g0544(.A(n1549), .Y(n1578));
  INVX1   g0545(.A(n1538), .Y(n1579));
  OAI22X1 g0546(.A0(n1535), .A1(n1531), .B0(SI_17_), .B1(n1579), .Y(n1580));
  AOI22X1 g0547(.A0(n1580), .A1(n1578), .B0(n1576), .B1(n1556), .Y(n1581));
  NOR2X1  g0548(.A(n1581), .B(n1577), .Y(n1582));
  AOI21X1 g0549(.A0(n1148), .A1(n1146), .B0(n1574), .Y(n1583));
  AOI21X1 g0550(.A0(n1156), .A1(P1_DATAO_REG_19__SCAN_IN), .B0(n1583), .Y(n1584));
  XOR2X1  g0551(.A(n1584), .B(SI_19_), .Y(n1585));
  XOR2X1  g0552(.A(n1585), .B(n1582), .Y(n1586));
  AOI21X1 g0553(.A0(n1586), .A1(n1149), .B0(n1575), .Y(n1587));
  NOR4X1  g0554(.A(P1_IR_REG_9__SCAN_IN), .B(P1_IR_REG_8__SCAN_IN), .C(P1_IR_REG_7__SCAN_IN), .D(n1293), .Y(n1588));
  INVX1   g0555(.A(P1_IR_REG_19__SCAN_IN), .Y(n1589));
  NAND4X1 g0556(.A(n1565), .B(n1512), .C(n1259), .D(n1589), .Y(n1590));
  NOR4X1  g0557(.A(n1241), .B(P1_IR_REG_17__SCAN_IN), .C(P1_IR_REG_15__SCAN_IN), .D(n1590), .Y(n1591));
  NAND2X1 g0558(.A(n1591), .B(n1588), .Y(n1592));
  NOR2X1  g0559(.A(n1592), .B(n1515), .Y(n1593));
  AOI21X1 g0560(.A0(n1569), .A1(P1_IR_REG_19__SCAN_IN), .B0(n1593), .Y(n1594));
  AOI22X1 g0561(.A0(n1184), .A1(n1594), .B0(n1162), .B1(P1_IR_REG_19__SCAN_IN), .Y(n1595));
  OAI21X1 g0562(.A0(n1587), .A1(P1_STATE_REG_SCAN_IN), .B0(n1595), .Y(P1_U3334));
  INVX1   g0563(.A(P2_DATAO_REG_20__SCAN_IN), .Y(n1597));
  NOR3X1  g0564(.A(n1153), .B(n1152), .C(n1597), .Y(n1598));
  INVX1   g0565(.A(SI_19_), .Y(n1599));
  NOR2X1  g0566(.A(n1584), .B(n1599), .Y(n1600));
  INVX1   g0567(.A(n1577), .Y(n1601));
  INVX1   g0568(.A(n1556), .Y(n1602));
  OAI22X1 g0569(.A0(n1553), .A1(n1549), .B0(SI_18_), .B1(n1602), .Y(n1603));
  AOI22X1 g0570(.A0(n1603), .A1(n1601), .B0(n1599), .B1(n1584), .Y(n1604));
  NOR2X1  g0571(.A(n1604), .B(n1600), .Y(n1605));
  AOI21X1 g0572(.A0(n1148), .A1(n1146), .B0(n1597), .Y(n1606));
  AOI21X1 g0573(.A0(n1156), .A1(P1_DATAO_REG_20__SCAN_IN), .B0(n1606), .Y(n1607));
  XOR2X1  g0574(.A(n1607), .B(SI_20_), .Y(n1608));
  XOR2X1  g0575(.A(n1608), .B(n1605), .Y(n1609));
  AOI21X1 g0576(.A0(n1609), .A1(n1149), .B0(n1598), .Y(n1610));
  NAND3X1 g0577(.A(n1591), .B(n1588), .C(n1563), .Y(n1611));
  NAND4X1 g0578(.A(n1492), .B(n1465), .C(n1447), .D(n1561), .Y(n1612));
  INVX1   g0579(.A(P1_IR_REG_20__SCAN_IN), .Y(n1613));
  NAND2X1 g0580(.A(n1568), .B(n1613), .Y(n1614));
  NAND3X1 g0581(.A(n1565), .B(n1542), .C(n1564), .Y(n1615));
  NOR3X1  g0582(.A(n1615), .B(P1_IR_REG_19__SCAN_IN), .C(P1_IR_REG_16__SCAN_IN), .Y(n1616));
  NAND2X1 g0583(.A(n1616), .B(n1588), .Y(n1617));
  NOR3X1  g0584(.A(n1617), .B(n1614), .C(n1612), .Y(n1618));
  AOI21X1 g0585(.A0(n1611), .A1(P1_IR_REG_20__SCAN_IN), .B0(n1618), .Y(n1619));
  AOI22X1 g0586(.A0(n1184), .A1(n1619), .B0(n1162), .B1(P1_IR_REG_20__SCAN_IN), .Y(n1620));
  OAI21X1 g0587(.A0(n1610), .A1(P1_STATE_REG_SCAN_IN), .B0(n1620), .Y(P1_U3333));
  INVX1   g0588(.A(P2_DATAO_REG_21__SCAN_IN), .Y(n1622));
  NOR3X1  g0589(.A(n1153), .B(n1152), .C(n1622), .Y(n1623));
  INVX1   g0590(.A(SI_20_), .Y(n1624));
  NOR2X1  g0591(.A(n1607), .B(n1624), .Y(n1625));
  INVX1   g0592(.A(n1600), .Y(n1626));
  INVX1   g0593(.A(n1584), .Y(n1627));
  OAI22X1 g0594(.A0(n1581), .A1(n1577), .B0(SI_19_), .B1(n1627), .Y(n1628));
  AOI22X1 g0595(.A0(n1628), .A1(n1626), .B0(n1624), .B1(n1607), .Y(n1629));
  NOR2X1  g0596(.A(n1629), .B(n1625), .Y(n1630));
  AOI21X1 g0597(.A0(n1148), .A1(n1146), .B0(n1622), .Y(n1631));
  AOI21X1 g0598(.A0(n1156), .A1(P1_DATAO_REG_21__SCAN_IN), .B0(n1631), .Y(n1632));
  XOR2X1  g0599(.A(n1632), .B(SI_21_), .Y(n1633));
  XOR2X1  g0600(.A(n1633), .B(n1630), .Y(n1634));
  AOI21X1 g0601(.A0(n1634), .A1(n1149), .B0(n1623), .Y(n1635));
  INVX1   g0602(.A(P1_IR_REG_21__SCAN_IN), .Y(n1636));
  XOR2X1  g0603(.A(n1618), .B(n1636), .Y(n1637));
  AOI22X1 g0604(.A0(n1184), .A1(n1637), .B0(n1162), .B1(P1_IR_REG_21__SCAN_IN), .Y(n1638));
  OAI21X1 g0605(.A0(n1635), .A1(P1_STATE_REG_SCAN_IN), .B0(n1638), .Y(P1_U3332));
  INVX1   g0606(.A(P2_DATAO_REG_22__SCAN_IN), .Y(n1640));
  NOR3X1  g0607(.A(n1153), .B(n1152), .C(n1640), .Y(n1641));
  INVX1   g0608(.A(SI_21_), .Y(n1642));
  NOR2X1  g0609(.A(n1632), .B(n1642), .Y(n1643));
  INVX1   g0610(.A(n1625), .Y(n1644));
  INVX1   g0611(.A(n1607), .Y(n1645));
  OAI22X1 g0612(.A0(n1604), .A1(n1600), .B0(SI_20_), .B1(n1645), .Y(n1646));
  AOI22X1 g0613(.A0(n1646), .A1(n1644), .B0(n1642), .B1(n1632), .Y(n1647));
  NOR2X1  g0614(.A(n1647), .B(n1643), .Y(n1648));
  AOI21X1 g0615(.A0(n1148), .A1(n1146), .B0(n1640), .Y(n1649));
  AOI21X1 g0616(.A0(n1156), .A1(P1_DATAO_REG_22__SCAN_IN), .B0(n1649), .Y(n1650));
  XOR2X1  g0617(.A(n1650), .B(SI_22_), .Y(n1651));
  XOR2X1  g0618(.A(n1651), .B(n1648), .Y(n1652));
  AOI21X1 g0619(.A0(n1652), .A1(n1149), .B0(n1641), .Y(n1653));
  NOR3X1  g0620(.A(P1_IR_REG_21__SCAN_IN), .B(P1_IR_REG_20__SCAN_IN), .C(P1_IR_REG_0__SCAN_IN), .Y(n1654));
  NAND3X1 g0621(.A(n1654), .B(n1520), .C(n1259), .Y(n1655));
  NOR2X1  g0622(.A(n1655), .B(n1612), .Y(n1656));
  NAND3X1 g0623(.A(n1656), .B(n1616), .C(n1588), .Y(n1657));
  INVX1   g0624(.A(P1_IR_REG_22__SCAN_IN), .Y(n1658));
  NAND4X1 g0625(.A(n1636), .B(n1613), .C(n1589), .D(n1658), .Y(n1659));
  NOR3X1  g0626(.A(n1659), .B(P1_IR_REG_18__SCAN_IN), .C(P1_IR_REG_17__SCAN_IN), .Y(n1660));
  AOI22X1 g0627(.A0(n1657), .A1(P1_IR_REG_22__SCAN_IN), .B0(n1522), .B1(n1660), .Y(n1661));
  AOI22X1 g0628(.A0(n1184), .A1(n1661), .B0(n1162), .B1(P1_IR_REG_22__SCAN_IN), .Y(n1662));
  OAI21X1 g0629(.A0(n1653), .A1(P1_STATE_REG_SCAN_IN), .B0(n1662), .Y(P1_U3331));
  INVX1   g0630(.A(P2_DATAO_REG_23__SCAN_IN), .Y(n1664));
  NOR3X1  g0631(.A(n1153), .B(n1152), .C(n1664), .Y(n1665));
  INVX1   g0632(.A(SI_22_), .Y(n1666));
  NOR2X1  g0633(.A(n1650), .B(n1666), .Y(n1667));
  INVX1   g0634(.A(n1643), .Y(n1668));
  INVX1   g0635(.A(n1632), .Y(n1669));
  OAI22X1 g0636(.A0(n1629), .A1(n1625), .B0(SI_21_), .B1(n1669), .Y(n1670));
  AOI22X1 g0637(.A0(n1670), .A1(n1668), .B0(n1666), .B1(n1650), .Y(n1671));
  NOR2X1  g0638(.A(n1671), .B(n1667), .Y(n1672));
  AOI21X1 g0639(.A0(n1148), .A1(n1146), .B0(n1664), .Y(n1673));
  AOI21X1 g0640(.A0(n1156), .A1(P1_DATAO_REG_23__SCAN_IN), .B0(n1673), .Y(n1674));
  XOR2X1  g0641(.A(n1674), .B(SI_23_), .Y(n1675));
  XOR2X1  g0642(.A(n1675), .B(n1672), .Y(n1676));
  AOI21X1 g0643(.A0(n1676), .A1(n1149), .B0(n1665), .Y(n1677));
  INVX1   g0644(.A(P1_IR_REG_23__SCAN_IN), .Y(n1678));
  AOI21X1 g0645(.A0(n1660), .A1(n1522), .B0(n1678), .Y(n1679));
  NAND3X1 g0646(.A(n1658), .B(n1636), .C(n1613), .Y(n1680));
  NAND3X1 g0647(.A(n1589), .B(n1565), .C(n1512), .Y(n1681));
  NOR3X1  g0648(.A(n1681), .B(n1680), .C(n1612), .Y(n1682));
  NOR3X1  g0649(.A(P1_IR_REG_9__SCAN_IN), .B(P1_IR_REG_8__SCAN_IN), .C(P1_IR_REG_7__SCAN_IN), .Y(n1683));
  NAND3X1 g0650(.A(n1683), .B(n1339), .C(n1259), .Y(n1684));
  NAND4X1 g0651(.A(n1200), .B(n1678), .C(n1542), .D(n1520), .Y(n1685));
  NOR2X1  g0652(.A(n1685), .B(n1684), .Y(n1686));
  AOI21X1 g0653(.A0(n1686), .A1(n1682), .B0(n1679), .Y(n1687));
  AOI22X1 g0654(.A0(n1184), .A1(n1687), .B0(n1162), .B1(P1_IR_REG_23__SCAN_IN), .Y(n1688));
  OAI21X1 g0655(.A0(n1677), .A1(P1_STATE_REG_SCAN_IN), .B0(n1688), .Y(P1_U3330));
  INVX1   g0656(.A(P2_DATAO_REG_24__SCAN_IN), .Y(n1690));
  NOR3X1  g0657(.A(n1153), .B(n1152), .C(n1690), .Y(n1691));
  INVX1   g0658(.A(SI_23_), .Y(n1692));
  NOR2X1  g0659(.A(n1674), .B(n1692), .Y(n1693));
  INVX1   g0660(.A(n1667), .Y(n1694));
  INVX1   g0661(.A(n1650), .Y(n1695));
  OAI22X1 g0662(.A0(n1647), .A1(n1643), .B0(SI_22_), .B1(n1695), .Y(n1696));
  AOI22X1 g0663(.A0(n1696), .A1(n1694), .B0(n1692), .B1(n1674), .Y(n1697));
  NOR2X1  g0664(.A(n1697), .B(n1693), .Y(n1698));
  AOI21X1 g0665(.A0(n1148), .A1(n1146), .B0(n1690), .Y(n1699));
  AOI21X1 g0666(.A0(n1156), .A1(P1_DATAO_REG_24__SCAN_IN), .B0(n1699), .Y(n1700));
  XOR2X1  g0667(.A(n1700), .B(SI_24_), .Y(n1701));
  XOR2X1  g0668(.A(n1701), .B(n1698), .Y(n1702));
  AOI21X1 g0669(.A0(n1702), .A1(n1149), .B0(n1691), .Y(n1703));
  INVX1   g0670(.A(P1_IR_REG_24__SCAN_IN), .Y(n1704));
  AOI21X1 g0671(.A0(n1686), .A1(n1682), .B0(n1704), .Y(n1705));
  NOR3X1  g0672(.A(P1_IR_REG_16__SCAN_IN), .B(P1_IR_REG_15__SCAN_IN), .C(P1_IR_REG_14__SCAN_IN), .Y(n1706));
  NOR4X1  g0673(.A(P1_IR_REG_19__SCAN_IN), .B(P1_IR_REG_18__SCAN_IN), .C(P1_IR_REG_17__SCAN_IN), .D(P1_IR_REG_20__SCAN_IN), .Y(n1707));
  NAND3X1 g0674(.A(n1707), .B(n1706), .C(n1200), .Y(n1708));
  NOR3X1  g0675(.A(P1_IR_REG_23__SCAN_IN), .B(P1_IR_REG_22__SCAN_IN), .C(P1_IR_REG_21__SCAN_IN), .Y(n1709));
  NAND3X1 g0676(.A(n1709), .B(n1520), .C(n1704), .Y(n1710));
  NOR4X1  g0677(.A(n1708), .B(n1684), .C(n1562), .D(n1710), .Y(n1711));
  NOR2X1  g0678(.A(n1711), .B(n1705), .Y(n1712));
  AOI22X1 g0679(.A0(n1184), .A1(n1712), .B0(n1162), .B1(P1_IR_REG_24__SCAN_IN), .Y(n1713));
  OAI21X1 g0680(.A0(n1703), .A1(P1_STATE_REG_SCAN_IN), .B0(n1713), .Y(P1_U3329));
  INVX1   g0681(.A(P2_DATAO_REG_25__SCAN_IN), .Y(n1715));
  NOR3X1  g0682(.A(n1153), .B(n1152), .C(n1715), .Y(n1716));
  INVX1   g0683(.A(SI_24_), .Y(n1717));
  NOR2X1  g0684(.A(n1700), .B(n1717), .Y(n1718));
  INVX1   g0685(.A(n1693), .Y(n1719));
  INVX1   g0686(.A(n1674), .Y(n1720));
  OAI22X1 g0687(.A0(n1671), .A1(n1667), .B0(SI_23_), .B1(n1720), .Y(n1721));
  AOI22X1 g0688(.A0(n1721), .A1(n1719), .B0(n1717), .B1(n1700), .Y(n1722));
  NOR2X1  g0689(.A(n1722), .B(n1718), .Y(n1723));
  AOI21X1 g0690(.A0(n1148), .A1(n1146), .B0(n1715), .Y(n1724));
  AOI21X1 g0691(.A0(n1156), .A1(P1_DATAO_REG_25__SCAN_IN), .B0(n1724), .Y(n1725));
  XOR2X1  g0692(.A(n1725), .B(SI_25_), .Y(n1726));
  XOR2X1  g0693(.A(n1726), .B(n1723), .Y(n1727));
  AOI21X1 g0694(.A0(n1727), .A1(n1149), .B0(n1716), .Y(n1728));
  INVX1   g0695(.A(P1_IR_REG_25__SCAN_IN), .Y(n1729));
  XOR2X1  g0696(.A(n1711), .B(n1729), .Y(n1730));
  AOI22X1 g0697(.A0(n1184), .A1(n1730), .B0(n1162), .B1(P1_IR_REG_25__SCAN_IN), .Y(n1731));
  OAI21X1 g0698(.A0(n1728), .A1(P1_STATE_REG_SCAN_IN), .B0(n1731), .Y(P1_U3328));
  INVX1   g0699(.A(P2_DATAO_REG_26__SCAN_IN), .Y(n1733));
  NOR3X1  g0700(.A(n1153), .B(n1152), .C(n1733), .Y(n1734));
  INVX1   g0701(.A(SI_25_), .Y(n1735));
  NOR2X1  g0702(.A(n1725), .B(n1735), .Y(n1736));
  INVX1   g0703(.A(n1718), .Y(n1737));
  INVX1   g0704(.A(n1700), .Y(n1738));
  OAI22X1 g0705(.A0(n1697), .A1(n1693), .B0(SI_24_), .B1(n1738), .Y(n1739));
  AOI22X1 g0706(.A0(n1739), .A1(n1737), .B0(n1735), .B1(n1725), .Y(n1740));
  NOR2X1  g0707(.A(n1740), .B(n1736), .Y(n1741));
  AOI21X1 g0708(.A0(n1148), .A1(n1146), .B0(n1733), .Y(n1742));
  AOI21X1 g0709(.A0(n1156), .A1(P1_DATAO_REG_26__SCAN_IN), .B0(n1742), .Y(n1743));
  XOR2X1  g0710(.A(n1743), .B(SI_26_), .Y(n1744));
  XOR2X1  g0711(.A(n1744), .B(n1741), .Y(n1745));
  AOI21X1 g0712(.A0(n1745), .A1(n1149), .B0(n1734), .Y(n1746));
  INVX1   g0713(.A(P1_IR_REG_26__SCAN_IN), .Y(n1747));
  NAND4X1 g0714(.A(n1520), .B(n1729), .C(n1704), .D(n1709), .Y(n1748));
  NOR4X1  g0715(.A(n1708), .B(n1684), .C(n1562), .D(n1748), .Y(n1749));
  NOR2X1  g0716(.A(n1749), .B(n1747), .Y(n1750));
  NOR4X1  g0717(.A(P1_IR_REG_18__SCAN_IN), .B(P1_IR_REG_17__SCAN_IN), .C(P1_IR_REG_1__SCAN_IN), .D(P1_IR_REG_19__SCAN_IN), .Y(n1751));
  NAND4X1 g0718(.A(n1706), .B(n1654), .C(n1514), .D(n1751), .Y(n1752));
  NOR4X1  g0719(.A(P1_IR_REG_24__SCAN_IN), .B(P1_IR_REG_23__SCAN_IN), .C(P1_IR_REG_22__SCAN_IN), .D(P1_IR_REG_25__SCAN_IN), .Y(n1753));
  NAND3X1 g0720(.A(n1753), .B(n1520), .C(n1747), .Y(n1754));
  NOR3X1  g0721(.A(n1754), .B(n1752), .C(n1684), .Y(n1755));
  NOR2X1  g0722(.A(n1755), .B(n1750), .Y(n1756));
  AOI22X1 g0723(.A0(n1184), .A1(n1756), .B0(n1162), .B1(P1_IR_REG_26__SCAN_IN), .Y(n1757));
  OAI21X1 g0724(.A0(n1746), .A1(P1_STATE_REG_SCAN_IN), .B0(n1757), .Y(P1_U3327));
  INVX1   g0725(.A(P2_DATAO_REG_27__SCAN_IN), .Y(n1759));
  NOR3X1  g0726(.A(n1153), .B(n1152), .C(n1759), .Y(n1760));
  INVX1   g0727(.A(SI_26_), .Y(n1761));
  NOR2X1  g0728(.A(n1743), .B(n1761), .Y(n1762));
  INVX1   g0729(.A(n1736), .Y(n1763));
  INVX1   g0730(.A(n1725), .Y(n1764));
  OAI22X1 g0731(.A0(n1722), .A1(n1718), .B0(SI_25_), .B1(n1764), .Y(n1765));
  AOI22X1 g0732(.A0(n1765), .A1(n1763), .B0(n1761), .B1(n1743), .Y(n1766));
  AOI21X1 g0733(.A0(n1148), .A1(n1146), .B0(n1759), .Y(n1767));
  AOI21X1 g0734(.A0(n1156), .A1(P1_DATAO_REG_27__SCAN_IN), .B0(n1767), .Y(n1768));
  XOR2X1  g0735(.A(n1768), .B(SI_27_), .Y(n1769));
  NOR3X1  g0736(.A(n1769), .B(n1766), .C(n1762), .Y(n1770));
  INVX1   g0737(.A(n1762), .Y(n1771));
  INVX1   g0738(.A(n1743), .Y(n1772));
  OAI22X1 g0739(.A0(n1740), .A1(n1736), .B0(SI_26_), .B1(n1772), .Y(n1773));
  INVX1   g0740(.A(n1769), .Y(n1774));
  AOI21X1 g0741(.A0(n1773), .A1(n1771), .B0(n1774), .Y(n1775));
  OAI21X1 g0742(.A0(n1775), .A1(n1770), .B0(n1149), .Y(n1776));
  INVX1   g0743(.A(n1776), .Y(n1777));
  OAI21X1 g0744(.A0(n1777), .A1(n1760), .B0(P1_U3084), .Y(n1778));
  INVX1   g0745(.A(P1_IR_REG_27__SCAN_IN), .Y(n1779));
  XOR2X1  g0746(.A(n1755), .B(n1779), .Y(n1780));
  AOI22X1 g0747(.A0(n1184), .A1(n1780), .B0(n1162), .B1(P1_IR_REG_27__SCAN_IN), .Y(n1781));
  NAND2X1 g0748(.A(n1781), .B(n1778), .Y(P1_U3326));
  INVX1   g0749(.A(P2_DATAO_REG_28__SCAN_IN), .Y(n1783));
  NOR3X1  g0750(.A(n1153), .B(n1152), .C(n1783), .Y(n1784));
  INVX1   g0751(.A(SI_27_), .Y(n1785));
  NOR2X1  g0752(.A(n1768), .B(n1785), .Y(n1786));
  AOI22X1 g0753(.A0(n1773), .A1(n1771), .B0(n1785), .B1(n1768), .Y(n1787));
  NOR2X1  g0754(.A(n1787), .B(n1786), .Y(n1788));
  AOI21X1 g0755(.A0(n1148), .A1(n1146), .B0(n1783), .Y(n1789));
  AOI21X1 g0756(.A0(n1156), .A1(P1_DATAO_REG_28__SCAN_IN), .B0(n1789), .Y(n1790));
  XOR2X1  g0757(.A(n1790), .B(SI_28_), .Y(n1791));
  XOR2X1  g0758(.A(n1791), .B(n1788), .Y(n1792));
  AOI21X1 g0759(.A0(n1792), .A1(n1149), .B0(n1784), .Y(n1793));
  INVX1   g0760(.A(P1_IR_REG_28__SCAN_IN), .Y(n1794));
  NAND2X1 g0761(.A(n1683), .B(n1342), .Y(n1795));
  NAND4X1 g0762(.A(n1779), .B(n1747), .C(n1199), .D(n1753), .Y(n1796));
  NOR3X1  g0763(.A(n1796), .B(n1795), .C(n1752), .Y(n1797));
  NAND4X1 g0764(.A(n1589), .B(n1565), .C(n1542), .D(n1200), .Y(n1798));
  NAND4X1 g0765(.A(n1658), .B(n1636), .C(n1613), .D(n1706), .Y(n1799));
  NOR3X1  g0766(.A(n1799), .B(n1798), .C(n1562), .Y(n1800));
  NAND4X1 g0767(.A(n1729), .B(n1704), .C(n1678), .D(n1747), .Y(n1801));
  NAND3X1 g0768(.A(n1794), .B(n1779), .C(n1199), .Y(n1802));
  NOR3X1  g0769(.A(n1802), .B(n1801), .C(n1795), .Y(n1803));
  NAND2X1 g0770(.A(n1803), .B(n1800), .Y(n1804));
  OAI21X1 g0771(.A0(n1797), .A1(n1794), .B0(n1804), .Y(n1805));
  NOR3X1  g0772(.A(n1805), .B(P1_U3084), .C(n1183), .Y(n1806));
  AOI21X1 g0773(.A0(n1162), .A1(P1_IR_REG_28__SCAN_IN), .B0(n1806), .Y(n1807));
  OAI21X1 g0774(.A0(n1793), .A1(P1_STATE_REG_SCAN_IN), .B0(n1807), .Y(P1_U3325));
  INVX1   g0775(.A(P2_DATAO_REG_29__SCAN_IN), .Y(n1809));
  NOR3X1  g0776(.A(n1153), .B(n1152), .C(n1809), .Y(n1810));
  INVX1   g0777(.A(SI_28_), .Y(n1811));
  NOR2X1  g0778(.A(n1790), .B(n1811), .Y(n1812));
  INVX1   g0779(.A(n1786), .Y(n1813));
  INVX1   g0780(.A(n1768), .Y(n1814));
  OAI22X1 g0781(.A0(n1766), .A1(n1762), .B0(SI_27_), .B1(n1814), .Y(n1815));
  AOI22X1 g0782(.A0(n1815), .A1(n1813), .B0(n1811), .B1(n1790), .Y(n1816));
  NOR2X1  g0783(.A(n1816), .B(n1812), .Y(n1817));
  AOI21X1 g0784(.A0(n1148), .A1(n1146), .B0(n1809), .Y(n1818));
  AOI21X1 g0785(.A0(n1156), .A1(P1_DATAO_REG_29__SCAN_IN), .B0(n1818), .Y(n1819));
  XOR2X1  g0786(.A(n1819), .B(SI_29_), .Y(n1820));
  XOR2X1  g0787(.A(n1820), .B(n1817), .Y(n1821));
  AOI21X1 g0788(.A0(n1821), .A1(n1149), .B0(n1810), .Y(n1822));
  NAND2X1 g0789(.A(n1804), .B(P1_IR_REG_29__SCAN_IN), .Y(n1823));
  NOR4X1  g0790(.A(n1801), .B(n1795), .C(P1_IR_REG_29__SCAN_IN), .D(n1802), .Y(n1824));
  NAND2X1 g0791(.A(n1824), .B(n1800), .Y(n1825));
  NAND2X1 g0792(.A(n1825), .B(n1823), .Y(n1826));
  NOR3X1  g0793(.A(n1826), .B(P1_U3084), .C(n1183), .Y(n1827));
  AOI21X1 g0794(.A0(n1162), .A1(P1_IR_REG_29__SCAN_IN), .B0(n1827), .Y(n1828));
  OAI21X1 g0795(.A0(n1822), .A1(P1_STATE_REG_SCAN_IN), .B0(n1828), .Y(P1_U3324));
  INVX1   g0796(.A(P2_DATAO_REG_30__SCAN_IN), .Y(n1830));
  NOR3X1  g0797(.A(n1153), .B(n1152), .C(n1830), .Y(n1831));
  INVX1   g0798(.A(SI_29_), .Y(n1832));
  NOR2X1  g0799(.A(n1819), .B(n1832), .Y(n1833));
  INVX1   g0800(.A(n1833), .Y(n1834));
  INVX1   g0801(.A(n1819), .Y(n1835));
  OAI22X1 g0802(.A0(n1816), .A1(n1812), .B0(SI_29_), .B1(n1835), .Y(n1836));
  AOI21X1 g0803(.A0(n1148), .A1(n1146), .B0(n1830), .Y(n1837));
  AOI21X1 g0804(.A0(n1156), .A1(P1_DATAO_REG_30__SCAN_IN), .B0(n1837), .Y(n1838));
  XOR2X1  g0805(.A(n1838), .B(SI_30_), .Y(n1839));
  INVX1   g0806(.A(n1839), .Y(n1840));
  NAND3X1 g0807(.A(n1840), .B(n1836), .C(n1834), .Y(n1841));
  INVX1   g0808(.A(n1812), .Y(n1842));
  INVX1   g0809(.A(n1790), .Y(n1843));
  OAI22X1 g0810(.A0(n1787), .A1(n1786), .B0(SI_28_), .B1(n1843), .Y(n1844));
  AOI22X1 g0811(.A0(n1844), .A1(n1842), .B0(n1832), .B1(n1819), .Y(n1845));
  OAI21X1 g0812(.A0(n1845), .A1(n1833), .B0(n1839), .Y(n1846));
  AOI21X1 g0813(.A0(n1846), .A1(n1841), .B0(n1156), .Y(n1847));
  NOR2X1  g0814(.A(n1847), .B(n1831), .Y(n1848));
  XOR2X1  g0815(.A(n1825), .B(P1_IR_REG_30__SCAN_IN), .Y(n1849));
  AOI22X1 g0816(.A0(n1184), .A1(n1849), .B0(n1162), .B1(P1_IR_REG_30__SCAN_IN), .Y(n1850));
  OAI21X1 g0817(.A0(n1848), .A1(P1_STATE_REG_SCAN_IN), .B0(n1850), .Y(P1_U3323));
  INVX1   g0818(.A(P2_DATAO_REG_31__SCAN_IN), .Y(n1852));
  NOR3X1  g0819(.A(n1153), .B(n1152), .C(n1852), .Y(n1853));
  INVX1   g0820(.A(SI_30_), .Y(n1854));
  AOI21X1 g0821(.A0(n1148), .A1(n1146), .B0(n1852), .Y(n1855));
  AOI21X1 g0822(.A0(n1156), .A1(P1_DATAO_REG_31__SCAN_IN), .B0(n1855), .Y(n1856));
  XOR2X1  g0823(.A(n1856), .B(SI_31_), .Y(n1857));
  AOI21X1 g0824(.A0(n1838), .A1(n1854), .B0(n1857), .Y(n1858));
  INVX1   g0825(.A(n1858), .Y(n1859));
  AOI21X1 g0826(.A0(n1836), .A1(n1834), .B0(n1859), .Y(n1860));
  NOR2X1  g0827(.A(n1838), .B(n1854), .Y(n1861));
  INVX1   g0828(.A(n1861), .Y(n1862));
  NAND3X1 g0829(.A(n1862), .B(n1857), .C(n1834), .Y(n1863));
  NAND3X1 g0830(.A(n1857), .B(n1838), .C(n1854), .Y(n1864));
  OAI21X1 g0831(.A0(n1862), .A1(n1857), .B0(n1864), .Y(n1865));
  INVX1   g0832(.A(n1865), .Y(n1866));
  OAI21X1 g0833(.A0(n1863), .A1(n1845), .B0(n1866), .Y(n1867));
  NOR3X1  g0834(.A(n1867), .B(n1860), .C(n1156), .Y(n1868));
  OAI21X1 g0835(.A0(n1868), .A1(n1853), .B0(P1_U3084), .Y(n1869));
  NOR2X1  g0836(.A(n1825), .B(P1_IR_REG_30__SCAN_IN), .Y(n1870));
  NAND3X1 g0837(.A(n1870), .B(P1_STATE_REG_SCAN_IN), .C(P1_IR_REG_31__SCAN_IN), .Y(n1871));
  NAND2X1 g0838(.A(n1871), .B(n1869), .Y(P1_U3322));
  NOR2X1  g0839(.A(P1_IR_REG_31__SCAN_IN), .B(n1678), .Y(n1873));
  AOI21X1 g0840(.A0(n1687), .A1(P1_IR_REG_31__SCAN_IN), .B0(n1873), .Y(n1874));
  INVX1   g0841(.A(n1874), .Y(n1875));
  NAND2X1 g0842(.A(n1712), .B(P1_IR_REG_31__SCAN_IN), .Y(n1876));
  OAI21X1 g0843(.A0(P1_IR_REG_31__SCAN_IN), .A1(n1704), .B0(n1876), .Y(n1877));
  INVX1   g0844(.A(n1877), .Y(n1878));
  NAND2X1 g0845(.A(n1756), .B(P1_IR_REG_31__SCAN_IN), .Y(n1879));
  OAI21X1 g0846(.A0(P1_IR_REG_31__SCAN_IN), .A1(n1747), .B0(n1879), .Y(n1880));
  INVX1   g0847(.A(n1880), .Y(n1881));
  NOR2X1  g0848(.A(P1_IR_REG_31__SCAN_IN), .B(n1729), .Y(n1882));
  AOI21X1 g0849(.A0(n1730), .A1(P1_IR_REG_31__SCAN_IN), .B0(n1882), .Y(n1883));
  NOR3X1  g0850(.A(n1883), .B(n1881), .C(n1878), .Y(n1884));
  INVX1   g0851(.A(P1_B_REG_SCAN_IN), .Y(n1885));
  INVX1   g0852(.A(n1883), .Y(n1886));
  NOR4X1  g0853(.A(n1881), .B(n1877), .C(n1885), .D(n1886), .Y(n1887));
  OAI21X1 g0854(.A0(n1878), .A1(P1_B_REG_SCAN_IN), .B0(n1880), .Y(n1888));
  NOR2X1  g0855(.A(n1888), .B(n1887), .Y(n1889));
  NOR4X1  g0856(.A(n1884), .B(n1875), .C(P1_U3084), .D(n1889), .Y(n1890));
  OAI21X1 g0857(.A0(n1886), .A1(n1881), .B0(n1878), .Y(n1891));
  NAND2X1 g0858(.A(n1891), .B(n1890), .Y(n1892));
  NOR3X1  g0859(.A(n1884), .B(n1875), .C(P1_U3084), .Y(n1893));
  INVX1   g0860(.A(n1893), .Y(n1894));
  OAI21X1 g0861(.A0(n1889), .A1(n1894), .B0(P1_D_REG_0__SCAN_IN), .Y(n1895));
  NAND2X1 g0862(.A(n1895), .B(n1892), .Y(P1_U3440));
  OAI21X1 g0863(.A0(n1886), .A1(n1880), .B0(n1890), .Y(n1897));
  OAI21X1 g0864(.A0(n1889), .A1(n1894), .B0(P1_D_REG_1__SCAN_IN), .Y(n1898));
  NAND2X1 g0865(.A(n1898), .B(n1897), .Y(P1_U3441));
  INVX1   g0866(.A(P1_D_REG_2__SCAN_IN), .Y(n1900));
  NOR2X1  g0867(.A(n1890), .B(n1900), .Y(P1_U3321));
  INVX1   g0868(.A(P1_D_REG_3__SCAN_IN), .Y(n1902));
  NOR2X1  g0869(.A(n1890), .B(n1902), .Y(P1_U3320));
  INVX1   g0870(.A(P1_D_REG_4__SCAN_IN), .Y(n1904));
  NOR2X1  g0871(.A(n1890), .B(n1904), .Y(P1_U3319));
  INVX1   g0872(.A(P1_D_REG_5__SCAN_IN), .Y(n1906));
  NOR2X1  g0873(.A(n1890), .B(n1906), .Y(P1_U3318));
  INVX1   g0874(.A(P1_D_REG_6__SCAN_IN), .Y(n1908));
  NOR2X1  g0875(.A(n1890), .B(n1908), .Y(P1_U3317));
  INVX1   g0876(.A(P1_D_REG_7__SCAN_IN), .Y(n1910));
  NOR2X1  g0877(.A(n1890), .B(n1910), .Y(P1_U3316));
  INVX1   g0878(.A(P1_D_REG_8__SCAN_IN), .Y(n1912));
  NOR2X1  g0879(.A(n1890), .B(n1912), .Y(P1_U3315));
  INVX1   g0880(.A(P1_D_REG_9__SCAN_IN), .Y(n1914));
  NOR2X1  g0881(.A(n1890), .B(n1914), .Y(P1_U3314));
  INVX1   g0882(.A(P1_D_REG_10__SCAN_IN), .Y(n1916));
  NOR2X1  g0883(.A(n1890), .B(n1916), .Y(P1_U3313));
  INVX1   g0884(.A(P1_D_REG_11__SCAN_IN), .Y(n1918));
  NOR2X1  g0885(.A(n1890), .B(n1918), .Y(P1_U3312));
  INVX1   g0886(.A(P1_D_REG_12__SCAN_IN), .Y(n1920));
  NOR2X1  g0887(.A(n1890), .B(n1920), .Y(P1_U3311));
  INVX1   g0888(.A(P1_D_REG_13__SCAN_IN), .Y(n1922));
  NOR2X1  g0889(.A(n1890), .B(n1922), .Y(P1_U3310));
  INVX1   g0890(.A(P1_D_REG_14__SCAN_IN), .Y(n1924));
  NOR2X1  g0891(.A(n1890), .B(n1924), .Y(P1_U3309));
  INVX1   g0892(.A(P1_D_REG_15__SCAN_IN), .Y(n1926));
  NOR2X1  g0893(.A(n1890), .B(n1926), .Y(P1_U3308));
  INVX1   g0894(.A(P1_D_REG_16__SCAN_IN), .Y(n1928));
  NOR2X1  g0895(.A(n1890), .B(n1928), .Y(P1_U3307));
  INVX1   g0896(.A(P1_D_REG_17__SCAN_IN), .Y(n1930));
  NOR2X1  g0897(.A(n1890), .B(n1930), .Y(P1_U3306));
  INVX1   g0898(.A(P1_D_REG_18__SCAN_IN), .Y(n1932));
  NOR2X1  g0899(.A(n1890), .B(n1932), .Y(P1_U3305));
  INVX1   g0900(.A(P1_D_REG_19__SCAN_IN), .Y(n1934));
  NOR2X1  g0901(.A(n1890), .B(n1934), .Y(P1_U3304));
  INVX1   g0902(.A(P1_D_REG_20__SCAN_IN), .Y(n1936));
  NOR2X1  g0903(.A(n1890), .B(n1936), .Y(P1_U3303));
  INVX1   g0904(.A(P1_D_REG_21__SCAN_IN), .Y(n1938));
  NOR2X1  g0905(.A(n1890), .B(n1938), .Y(P1_U3302));
  INVX1   g0906(.A(P1_D_REG_22__SCAN_IN), .Y(n1940));
  NOR2X1  g0907(.A(n1890), .B(n1940), .Y(P1_U3301));
  INVX1   g0908(.A(P1_D_REG_23__SCAN_IN), .Y(n1942));
  NOR2X1  g0909(.A(n1890), .B(n1942), .Y(P1_U3300));
  INVX1   g0910(.A(P1_D_REG_24__SCAN_IN), .Y(n1944));
  NOR2X1  g0911(.A(n1890), .B(n1944), .Y(P1_U3299));
  INVX1   g0912(.A(P1_D_REG_25__SCAN_IN), .Y(n1946));
  NOR2X1  g0913(.A(n1890), .B(n1946), .Y(P1_U3298));
  INVX1   g0914(.A(P1_D_REG_26__SCAN_IN), .Y(n1948));
  NOR2X1  g0915(.A(n1890), .B(n1948), .Y(P1_U3297));
  INVX1   g0916(.A(P1_D_REG_27__SCAN_IN), .Y(n1950));
  NOR2X1  g0917(.A(n1890), .B(n1950), .Y(P1_U3296));
  INVX1   g0918(.A(P1_D_REG_28__SCAN_IN), .Y(n1952));
  NOR2X1  g0919(.A(n1890), .B(n1952), .Y(P1_U3295));
  INVX1   g0920(.A(P1_D_REG_29__SCAN_IN), .Y(n1954));
  NOR2X1  g0921(.A(n1890), .B(n1954), .Y(P1_U3294));
  INVX1   g0922(.A(P1_D_REG_30__SCAN_IN), .Y(n1956));
  NOR2X1  g0923(.A(n1890), .B(n1956), .Y(P1_U3293));
  INVX1   g0924(.A(P1_D_REG_31__SCAN_IN), .Y(n1958));
  NOR2X1  g0925(.A(n1890), .B(n1958), .Y(P1_U3292));
  OAI21X1 g0926(.A0(P1_D_REG_7__SCAN_IN), .A1(P1_D_REG_3__SCAN_IN), .B0(n1889), .Y(n1960));
  OAI21X1 g0927(.A0(P1_D_REG_9__SCAN_IN), .A1(P1_D_REG_8__SCAN_IN), .B0(n1889), .Y(n1961));
  OAI21X1 g0928(.A0(P1_D_REG_10__SCAN_IN), .A1(P1_D_REG_5__SCAN_IN), .B0(n1889), .Y(n1962));
  OAI21X1 g0929(.A0(P1_D_REG_6__SCAN_IN), .A1(P1_D_REG_4__SCAN_IN), .B0(n1889), .Y(n1963));
  NAND4X1 g0930(.A(n1962), .B(n1961), .C(n1960), .D(n1963), .Y(n1964));
  OAI21X1 g0931(.A0(P1_D_REG_28__SCAN_IN), .A1(P1_D_REG_27__SCAN_IN), .B0(n1889), .Y(n1965));
  OAI21X1 g0932(.A0(P1_D_REG_26__SCAN_IN), .A1(P1_D_REG_25__SCAN_IN), .B0(n1889), .Y(n1966));
  OAI21X1 g0933(.A0(P1_D_REG_31__SCAN_IN), .A1(P1_D_REG_30__SCAN_IN), .B0(n1889), .Y(n1967));
  OAI21X1 g0934(.A0(P1_D_REG_29__SCAN_IN), .A1(P1_D_REG_2__SCAN_IN), .B0(n1889), .Y(n1968));
  NAND4X1 g0935(.A(n1967), .B(n1966), .C(n1965), .D(n1968), .Y(n1969));
  OAI21X1 g0936(.A0(P1_D_REG_21__SCAN_IN), .A1(P1_D_REG_20__SCAN_IN), .B0(n1889), .Y(n1970));
  OAI21X1 g0937(.A0(P1_D_REG_19__SCAN_IN), .A1(P1_D_REG_18__SCAN_IN), .B0(n1889), .Y(n1971));
  OAI21X1 g0938(.A0(P1_D_REG_23__SCAN_IN), .A1(P1_D_REG_22__SCAN_IN), .B0(n1889), .Y(n1972));
  NAND3X1 g0939(.A(n1972), .B(n1971), .C(n1970), .Y(n1973));
  OAI21X1 g0940(.A0(P1_D_REG_14__SCAN_IN), .A1(P1_D_REG_12__SCAN_IN), .B0(n1889), .Y(n1974));
  OAI21X1 g0941(.A0(P1_D_REG_13__SCAN_IN), .A1(P1_D_REG_11__SCAN_IN), .B0(n1889), .Y(n1975));
  OAI21X1 g0942(.A0(P1_D_REG_24__SCAN_IN), .A1(P1_D_REG_16__SCAN_IN), .B0(n1889), .Y(n1976));
  OAI21X1 g0943(.A0(P1_D_REG_17__SCAN_IN), .A1(P1_D_REG_15__SCAN_IN), .B0(n1889), .Y(n1977));
  NAND4X1 g0944(.A(n1976), .B(n1975), .C(n1974), .D(n1977), .Y(n1978));
  NOR4X1  g0945(.A(n1973), .B(n1969), .C(n1964), .D(n1978), .Y(n1979));
  INVX1   g0946(.A(n1979), .Y(n1980));
  AOI21X1 g0947(.A0(n1883), .A1(n1881), .B0(n1889), .Y(n1981));
  AOI21X1 g0948(.A0(n1889), .A1(P1_D_REG_1__SCAN_IN), .B0(n1981), .Y(n1982));
  NOR2X1  g0949(.A(P1_IR_REG_31__SCAN_IN), .B(n1658), .Y(n1983));
  AOI21X1 g0950(.A0(n1661), .A1(P1_IR_REG_31__SCAN_IN), .B0(n1983), .Y(n1984));
  INVX1   g0951(.A(n1984), .Y(n1985));
  NOR2X1  g0952(.A(P1_IR_REG_31__SCAN_IN), .B(n1613), .Y(n1986));
  AOI21X1 g0953(.A0(n1619), .A1(P1_IR_REG_31__SCAN_IN), .B0(n1986), .Y(n1987));
  NOR2X1  g0954(.A(P1_IR_REG_31__SCAN_IN), .B(n1636), .Y(n1988));
  AOI21X1 g0955(.A0(n1637), .A1(P1_IR_REG_31__SCAN_IN), .B0(n1988), .Y(n1989));
  AOI21X1 g0956(.A0(n1989), .A1(n1987), .B0(n1985), .Y(n1990));
  INVX1   g0957(.A(n1989), .Y(n1991));
  NOR2X1  g0958(.A(P1_IR_REG_31__SCAN_IN), .B(n1589), .Y(n1992));
  AOI21X1 g0959(.A0(n1594), .A1(P1_IR_REG_31__SCAN_IN), .B0(n1992), .Y(n1993));
  NAND2X1 g0960(.A(n1993), .B(n1987), .Y(n1994));
  OAI21X1 g0961(.A0(n1991), .A1(n1984), .B0(n1994), .Y(n1995));
  OAI21X1 g0962(.A0(n1995), .A1(n1990), .B0(n1982), .Y(n1996));
  NOR2X1  g0963(.A(n1996), .B(n1980), .Y(n1997));
  AOI21X1 g0964(.A0(n1881), .A1(n1878), .B0(n1889), .Y(n1998));
  AOI21X1 g0965(.A0(n1889), .A1(P1_D_REG_0__SCAN_IN), .B0(n1998), .Y(n1999));
  NAND3X1 g0966(.A(n1999), .B(n1997), .C(n1893), .Y(n2000));
  NAND2X1 g0967(.A(n1780), .B(P1_IR_REG_31__SCAN_IN), .Y(n2001));
  OAI21X1 g0968(.A0(P1_IR_REG_31__SCAN_IN), .A1(n1779), .B0(n2001), .Y(n2002));
  NOR2X1  g0969(.A(n1805), .B(n1183), .Y(n2003));
  NOR2X1  g0970(.A(P1_IR_REG_31__SCAN_IN), .B(n1794), .Y(n2004));
  NOR3X1  g0971(.A(n2004), .B(n2003), .C(n2002), .Y(n2005));
  NAND2X1 g0972(.A(P1_IR_REG_31__SCAN_IN), .B(P1_IR_REG_0__SCAN_IN), .Y(n2006));
  NAND2X1 g0973(.A(n1183), .B(P1_IR_REG_0__SCAN_IN), .Y(n2007));
  NAND2X1 g0974(.A(n2007), .B(n2006), .Y(n2008));
  NOR2X1  g0975(.A(n2005), .B(n1160), .Y(n2009));
  AOI21X1 g0976(.A0(n2008), .A1(n2005), .B0(n2009), .Y(n2010));
  INVX1   g0977(.A(P1_REG0_REG_0__SCAN_IN), .Y(n2011));
  INVX1   g0978(.A(P1_IR_REG_30__SCAN_IN), .Y(n2012));
  NAND2X1 g0979(.A(n1849), .B(P1_IR_REG_31__SCAN_IN), .Y(n2013));
  OAI21X1 g0980(.A0(P1_IR_REG_31__SCAN_IN), .A1(n2012), .B0(n2013), .Y(n2014));
  NAND2X1 g0981(.A(n1183), .B(P1_IR_REG_29__SCAN_IN), .Y(n2015));
  OAI21X1 g0982(.A0(n1826), .A1(n1183), .B0(n2015), .Y(n2016));
  NOR3X1  g0983(.A(n2016), .B(n2014), .C(n2011), .Y(n2017));
  INVX1   g0984(.A(P1_REG2_REG_0__SCAN_IN), .Y(n2018));
  NOR2X1  g0985(.A(P1_IR_REG_31__SCAN_IN), .B(n2012), .Y(n2019));
  AOI21X1 g0986(.A0(n1849), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2019), .Y(n2020));
  NOR3X1  g0987(.A(n2016), .B(n2020), .C(n2018), .Y(n2021));
  NOR2X1  g0988(.A(n2021), .B(n2017), .Y(n2022));
  NAND3X1 g0989(.A(n2016), .B(n2020), .C(P1_REG1_REG_0__SCAN_IN), .Y(n2023));
  NAND3X1 g0990(.A(n2016), .B(n2014), .C(P1_REG3_REG_0__SCAN_IN), .Y(n2024));
  NAND3X1 g0991(.A(n2024), .B(n2023), .C(n2022), .Y(n2025));
  XOR2X1  g0992(.A(n2025), .B(n2010), .Y(n2026));
  INVX1   g0993(.A(n1987), .Y(n2027));
  NOR3X1  g0994(.A(n1993), .B(n2027), .C(n1984), .Y(n2028));
  INVX1   g0995(.A(n2028), .Y(n2029));
  NOR2X1  g0996(.A(n2029), .B(n2026), .Y(n2030));
  INVX1   g0997(.A(n2030), .Y(n2031));
  NAND2X1 g0998(.A(n2024), .B(n2023), .Y(n2032));
  NOR4X1  g0999(.A(n2021), .B(n2017), .C(n2010), .D(n2032), .Y(n2033));
  NAND2X1 g1000(.A(n2008), .B(n2005), .Y(n2034));
  OAI21X1 g1001(.A0(n2005), .A1(n1160), .B0(n2034), .Y(n2035));
  INVX1   g1002(.A(n2025), .Y(n2036));
  NOR2X1  g1003(.A(n2036), .B(n2035), .Y(n2037));
  NOR3X1  g1004(.A(n1993), .B(n1989), .C(n1987), .Y(n2038));
  NAND2X1 g1005(.A(n1569), .B(P1_IR_REG_19__SCAN_IN), .Y(n2039));
  NAND3X1 g1006(.A(n1611), .B(n2039), .C(P1_IR_REG_31__SCAN_IN), .Y(n2040));
  OAI21X1 g1007(.A0(P1_IR_REG_31__SCAN_IN), .A1(n1589), .B0(n2040), .Y(n2041));
  NOR3X1  g1008(.A(n2041), .B(n1987), .C(n1984), .Y(n2042));
  OAI22X1 g1009(.A0(n2038), .A1(n2042), .B0(n2037), .B1(n2033), .Y(n2043));
  NOR3X1  g1010(.A(n1993), .B(n1987), .C(n1984), .Y(n2044));
  NOR3X1  g1011(.A(n2041), .B(n1989), .C(n1987), .Y(n2045));
  OAI22X1 g1012(.A0(n2044), .A1(n2045), .B0(n2037), .B1(n2033), .Y(n2046));
  NOR3X1  g1013(.A(n1994), .B(n1989), .C(n1985), .Y(n2047));
  NAND3X1 g1014(.A(n1993), .B(n1987), .C(n1985), .Y(n2048));
  NOR2X1  g1015(.A(n2048), .B(n1991), .Y(n2049));
  OAI22X1 g1016(.A0(n2047), .A1(n2049), .B0(n2037), .B1(n2033), .Y(n2050));
  NAND4X1 g1017(.A(n2046), .B(n2043), .C(n2031), .D(n2050), .Y(n2051));
  NOR3X1  g1018(.A(n1993), .B(n2027), .C(n1985), .Y(n2052));
  INVX1   g1019(.A(n2052), .Y(n2053));
  NOR4X1  g1020(.A(n2003), .B(n1989), .C(n1984), .D(n2004), .Y(n2054));
  INVX1   g1021(.A(P1_REG2_REG_1__SCAN_IN), .Y(n2055));
  NOR3X1  g1022(.A(n2016), .B(n2020), .C(n2055), .Y(n2056));
  INVX1   g1023(.A(P1_REG0_REG_1__SCAN_IN), .Y(n2057));
  NOR3X1  g1024(.A(n2016), .B(n2014), .C(n2057), .Y(n2058));
  NOR2X1  g1025(.A(n2058), .B(n2056), .Y(n2059));
  NAND3X1 g1026(.A(n2016), .B(n2020), .C(P1_REG1_REG_1__SCAN_IN), .Y(n2060));
  NAND3X1 g1027(.A(n2016), .B(n2014), .C(P1_REG3_REG_1__SCAN_IN), .Y(n2061));
  NAND3X1 g1028(.A(n2061), .B(n2060), .C(n2059), .Y(n2062));
  NOR3X1  g1029(.A(n1991), .B(n2027), .C(n1985), .Y(n2063));
  INVX1   g1030(.A(n2063), .Y(n2064));
  NOR2X1  g1031(.A(n2041), .B(n1987), .Y(n2065));
  NOR2X1  g1032(.A(n1993), .B(n1985), .Y(n2066));
  NOR2X1  g1033(.A(n1991), .B(n1985), .Y(n2067));
  AOI22X1 g1034(.A0(n2066), .A1(n1989), .B0(n2065), .B1(n2067), .Y(n2068));
  AOI21X1 g1035(.A0(n2068), .A1(n2064), .B0(n2010), .Y(n2069));
  AOI21X1 g1036(.A0(n2062), .A1(n2054), .B0(n2069), .Y(n2070));
  OAI21X1 g1037(.A0(n2053), .A1(n2026), .B0(n2070), .Y(n2071));
  NOR2X1  g1038(.A(n2071), .B(n2051), .Y(n2072));
  NAND2X1 g1039(.A(n2000), .B(P1_REG0_REG_0__SCAN_IN), .Y(n2073));
  OAI21X1 g1040(.A0(n2072), .A1(n2000), .B0(n2073), .Y(P1_U3454));
  NAND2X1 g1041(.A(n2061), .B(n2060), .Y(n2075));
  NOR3X1  g1042(.A(n2075), .B(n2058), .C(n2056), .Y(n2076));
  NOR2X1  g1043(.A(P1_IR_REG_31__SCAN_IN), .B(n1564), .Y(n2077));
  AOI21X1 g1044(.A0(n1185), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2077), .Y(n2078));
  NOR4X1  g1045(.A(n2004), .B(n2003), .C(n2002), .D(n2078), .Y(n2079));
  INVX1   g1046(.A(n2079), .Y(n2080));
  OAI21X1 g1047(.A0(n2005), .A1(n1182), .B0(n2080), .Y(n2081));
  XOR2X1  g1048(.A(n2081), .B(n2076), .Y(n2082));
  NAND2X1 g1049(.A(n2025), .B(n2035), .Y(n2083));
  INVX1   g1050(.A(n2083), .Y(n2084));
  XOR2X1  g1051(.A(n2084), .B(n2082), .Y(n2085));
  INVX1   g1052(.A(n2085), .Y(n2086));
  OAI21X1 g1053(.A0(n2049), .A1(n2042), .B0(n2086), .Y(n2087));
  XOR2X1  g1054(.A(n2082), .B(n2033), .Y(n2089));
  INVX1   g1055(.A(n2089), .Y(n2090));
  AOI22X1 g1056(.A0(n2086), .A1(n2047), .B0(n2038), .B1(n2090), .Y(n2091));
  NOR2X1  g1057(.A(n2004), .B(n2003), .Y(n2092));
  NOR3X1  g1058(.A(n2092), .B(n1989), .C(n1984), .Y(n2093));
  AOI22X1 g1059(.A0(n2090), .A1(n2045), .B0(n2025), .B1(n2093), .Y(n2094));
  OAI21X1 g1060(.A0(n2044), .A1(n2028), .B0(n2090), .Y(n2095));
  NAND4X1 g1061(.A(n2094), .B(n2091), .C(n2087), .D(n2095), .Y(n2096));
  INVX1   g1062(.A(n1166), .Y(n2097));
  NAND2X1 g1063(.A(n1180), .B(n1178), .Y(n2098));
  AOI21X1 g1064(.A0(n1172), .A1(n1167), .B0(n2098), .Y(n2099));
  OAI21X1 g1065(.A0(n2099), .A1(n1156), .B0(n2097), .Y(n2100));
  INVX1   g1066(.A(n2005), .Y(n2101));
  AOI21X1 g1067(.A0(n2101), .A1(n2100), .B0(n2079), .Y(n2102));
  XOR2X1  g1068(.A(n2102), .B(n2010), .Y(n2103));
  INVX1   g1069(.A(n2054), .Y(n2104));
  NOR2X1  g1070(.A(n2016), .B(n2014), .Y(n2105));
  NOR2X1  g1071(.A(n2016), .B(n2020), .Y(n2106));
  AOI22X1 g1072(.A0(n2105), .A1(P1_REG0_REG_2__SCAN_IN), .B0(P1_REG2_REG_2__SCAN_IN), .B1(n2106), .Y(n2107));
  NAND3X1 g1073(.A(n2016), .B(n2020), .C(P1_REG1_REG_2__SCAN_IN), .Y(n2108));
  NAND3X1 g1074(.A(n2016), .B(n2014), .C(P1_REG3_REG_2__SCAN_IN), .Y(n2109));
  NAND3X1 g1075(.A(n2109), .B(n2108), .C(n2107), .Y(n2110));
  INVX1   g1076(.A(n2110), .Y(n2111));
  OAI22X1 g1077(.A0(n2102), .A1(n2068), .B0(n2104), .B1(n2111), .Y(n2112));
  AOI21X1 g1078(.A0(n2103), .A1(n2063), .B0(n2112), .Y(n2113));
  OAI21X1 g1079(.A0(n2085), .A1(n2053), .B0(n2113), .Y(n2114));
  NOR2X1  g1080(.A(n2114), .B(n2096), .Y(n2115));
  NAND2X1 g1081(.A(n2000), .B(P1_REG0_REG_1__SCAN_IN), .Y(n2116));
  OAI21X1 g1082(.A0(n2115), .A1(n2000), .B0(n2116), .Y(P1_U3457));
  NOR2X1  g1083(.A(P1_IR_REG_31__SCAN_IN), .B(n1199), .Y(n2118));
  AOI21X1 g1084(.A0(n1201), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2118), .Y(n2119));
  INVX1   g1085(.A(n2119), .Y(n2120));
  NAND2X1 g1086(.A(n2120), .B(n2005), .Y(n2121));
  OAI21X1 g1087(.A0(n2005), .A1(n1198), .B0(n2121), .Y(n2122));
  XOR2X1  g1088(.A(n2122), .B(n2110), .Y(n2123));
  NAND2X1 g1089(.A(n2081), .B(n2062), .Y(n2124));
  NOR2X1  g1090(.A(n2081), .B(n2062), .Y(n2125));
  OAI21X1 g1091(.A0(n2083), .A1(n2125), .B0(n2124), .Y(n2126));
  NOR2X1  g1092(.A(n2123), .B(n2126), .Y(n2128));
  AOI21X1 g1093(.A0(n2126), .A1(n2123), .B0(n2128), .Y(n2129));
  AOI22X1 g1094(.A0(n2093), .A1(n2062), .B0(n2047), .B1(n2129), .Y(n2130));
  OAI21X1 g1095(.A0(n2049), .A1(n2042), .B0(n2129), .Y(n2131));
  NAND4X1 g1096(.A(n2023), .B(n2022), .C(n2035), .D(n2024), .Y(n2132));
  AOI21X1 g1097(.A0(n2076), .A1(n2033), .B0(n2081), .Y(n2133));
  AOI21X1 g1098(.A0(n2062), .A1(n2132), .B0(n2133), .Y(n2134));
  XOR2X1  g1099(.A(n2134), .B(n2123), .Y(n2135));
  OAI21X1 g1100(.A0(n2045), .A1(n2044), .B0(n2135), .Y(n2136));
  OAI21X1 g1101(.A0(n2038), .A1(n2028), .B0(n2135), .Y(n2137));
  NAND4X1 g1102(.A(n2136), .B(n2131), .C(n2130), .D(n2137), .Y(n2138));
  NAND2X1 g1103(.A(n2129), .B(n2052), .Y(n2139));
  NOR2X1  g1104(.A(n2005), .B(n1198), .Y(n2140));
  AOI21X1 g1105(.A0(n2120), .A1(n2005), .B0(n2140), .Y(n2141));
  NOR2X1  g1106(.A(n2081), .B(n2035), .Y(n2142));
  XOR2X1  g1107(.A(n2142), .B(n2141), .Y(n2143));
  INVX1   g1108(.A(P1_REG2_REG_3__SCAN_IN), .Y(n2144));
  NOR2X1  g1109(.A(n1826), .B(n1183), .Y(n2145));
  AOI21X1 g1110(.A0(n1183), .A1(P1_IR_REG_29__SCAN_IN), .B0(n2145), .Y(n2146));
  NAND2X1 g1111(.A(n2146), .B(n2014), .Y(n2147));
  NAND2X1 g1112(.A(n2105), .B(P1_REG0_REG_3__SCAN_IN), .Y(n2148));
  OAI21X1 g1113(.A0(n2147), .A1(n2144), .B0(n2148), .Y(n2149));
  INVX1   g1114(.A(P1_REG1_REG_3__SCAN_IN), .Y(n2150));
  NAND2X1 g1115(.A(n2016), .B(n2020), .Y(n2151));
  NAND2X1 g1116(.A(n2016), .B(n2014), .Y(n2152));
  OAI22X1 g1117(.A0(n2151), .A1(n2150), .B0(P1_REG3_REG_3__SCAN_IN), .B1(n2152), .Y(n2153));
  NOR2X1  g1118(.A(n2153), .B(n2149), .Y(n2154));
  OAI22X1 g1119(.A0(n2141), .A1(n2068), .B0(n2104), .B1(n2154), .Y(n2155));
  AOI21X1 g1120(.A0(n2143), .A1(n2063), .B0(n2155), .Y(n2156));
  NAND2X1 g1121(.A(n2156), .B(n2139), .Y(n2157));
  NOR2X1  g1122(.A(n2157), .B(n2138), .Y(n2158));
  NAND2X1 g1123(.A(n2000), .B(P1_REG0_REG_2__SCAN_IN), .Y(n2159));
  OAI21X1 g1124(.A0(n2158), .A1(n2000), .B0(n2159), .Y(P1_U3460));
  NAND2X1 g1125(.A(n2122), .B(n2110), .Y(n2161));
  NOR2X1  g1126(.A(n2122), .B(n2110), .Y(n2162));
  OAI21X1 g1127(.A0(n2162), .A1(n2124), .B0(n2161), .Y(n2163));
  NOR3X1  g1128(.A(n2162), .B(n2083), .C(n2125), .Y(n2164));
  AOI22X1 g1129(.A0(n2105), .A1(P1_REG0_REG_3__SCAN_IN), .B0(P1_REG2_REG_3__SCAN_IN), .B1(n2106), .Y(n2165));
  INVX1   g1130(.A(n2153), .Y(n2166));
  NAND2X1 g1131(.A(n2166), .B(n2165), .Y(n2167));
  NOR2X1  g1132(.A(P1_IR_REG_31__SCAN_IN), .B(n1214), .Y(n2168));
  AOI21X1 g1133(.A0(n1216), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2168), .Y(n2169));
  INVX1   g1134(.A(n2169), .Y(n2170));
  NAND2X1 g1135(.A(n2170), .B(n2005), .Y(n2171));
  OAI21X1 g1136(.A0(n2005), .A1(n1213), .B0(n2171), .Y(n2172));
  INVX1   g1137(.A(n2172), .Y(n2173));
  XOR2X1  g1138(.A(n2173), .B(n2167), .Y(n2174));
  NOR3X1  g1139(.A(n2174), .B(n2164), .C(n2163), .Y(n2175));
  NOR2X1  g1140(.A(n2164), .B(n2163), .Y(n2176));
  XOR2X1  g1141(.A(n2172), .B(n2167), .Y(n2177));
  NOR2X1  g1142(.A(n2177), .B(n2176), .Y(n2178));
  NOR2X1  g1143(.A(n2178), .B(n2175), .Y(n2179));
  INVX1   g1144(.A(n2179), .Y(n2180));
  AOI22X1 g1145(.A0(n2110), .A1(n2093), .B0(n2047), .B1(n2180), .Y(n2181));
  OAI22X1 g1146(.A0(n2175), .A1(n2178), .B0(n2049), .B1(n2042), .Y(n2182));
  INVX1   g1147(.A(n2044), .Y(n2183));
  INVX1   g1148(.A(n2045), .Y(n2184));
  NOR2X1  g1149(.A(n2122), .B(n2111), .Y(n2185));
  OAI21X1 g1150(.A0(n2062), .A1(n2132), .B0(n2102), .Y(n2186));
  OAI21X1 g1151(.A0(n2076), .A1(n2033), .B0(n2186), .Y(n2187));
  NAND4X1 g1152(.A(n2109), .B(n2108), .C(n2107), .D(n2122), .Y(n2188));
  INVX1   g1153(.A(n2188), .Y(n2189));
  NOR2X1  g1154(.A(n2174), .B(n2189), .Y(n2190));
  OAI21X1 g1155(.A0(n2187), .A1(n2185), .B0(n2190), .Y(n2191));
  NAND2X1 g1156(.A(n2141), .B(n2110), .Y(n2192));
  NAND2X1 g1157(.A(n2187), .B(n2188), .Y(n2193));
  NAND3X1 g1158(.A(n2193), .B(n2174), .C(n2192), .Y(n2194));
  AOI22X1 g1159(.A0(n2191), .A1(n2194), .B0(n2184), .B1(n2183), .Y(n2195));
  INVX1   g1160(.A(n2038), .Y(n2196));
  AOI22X1 g1161(.A0(n2191), .A1(n2194), .B0(n2196), .B1(n2029), .Y(n2197));
  NOR2X1  g1162(.A(n2197), .B(n2195), .Y(n2198));
  NAND3X1 g1163(.A(n2198), .B(n2182), .C(n2181), .Y(n2199));
  NOR3X1  g1164(.A(n2122), .B(n2081), .C(n2035), .Y(n2200));
  XOR2X1  g1165(.A(n2173), .B(n2200), .Y(n2201));
  AOI22X1 g1166(.A0(n2105), .A1(P1_REG0_REG_4__SCAN_IN), .B0(P1_REG2_REG_4__SCAN_IN), .B1(n2106), .Y(n2202));
  INVX1   g1167(.A(P1_REG1_REG_4__SCAN_IN), .Y(n2203));
  INVX1   g1168(.A(P1_REG3_REG_4__SCAN_IN), .Y(n2204));
  XOR2X1  g1169(.A(P1_REG3_REG_3__SCAN_IN), .B(n2204), .Y(n2205));
  OAI22X1 g1170(.A0(n2152), .A1(n2205), .B0(n2151), .B1(n2203), .Y(n2206));
  INVX1   g1171(.A(n2206), .Y(n2207));
  NAND2X1 g1172(.A(n2207), .B(n2202), .Y(n2208));
  INVX1   g1173(.A(n2208), .Y(n2209));
  OAI22X1 g1174(.A0(n2173), .A1(n2068), .B0(n2104), .B1(n2209), .Y(n2210));
  AOI21X1 g1175(.A0(n2201), .A1(n2063), .B0(n2210), .Y(n2211));
  OAI21X1 g1176(.A0(n2179), .A1(n2053), .B0(n2211), .Y(n2212));
  NOR2X1  g1177(.A(n2212), .B(n2199), .Y(n2213));
  NAND2X1 g1178(.A(n2000), .B(P1_REG0_REG_3__SCAN_IN), .Y(n2214));
  OAI21X1 g1179(.A0(n2213), .A1(n2000), .B0(n2214), .Y(P1_U3463));
  INVX1   g1180(.A(n2042), .Y(n2216));
  INVX1   g1181(.A(n2049), .Y(n2217));
  NOR2X1  g1182(.A(P1_IR_REG_31__SCAN_IN), .B(n1259), .Y(n2218));
  AOI21X1 g1183(.A0(n1243), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2218), .Y(n2219));
  INVX1   g1184(.A(n2219), .Y(n2220));
  NAND2X1 g1185(.A(n2220), .B(n2005), .Y(n2221));
  OAI21X1 g1186(.A0(n2005), .A1(n1240), .B0(n2221), .Y(n2222));
  INVX1   g1187(.A(n2222), .Y(n2223));
  XOR2X1  g1188(.A(n2223), .B(n2208), .Y(n2224));
  NOR3X1  g1189(.A(n2172), .B(n2153), .C(n2149), .Y(n2227));
  NOR2X1  g1190(.A(n2227), .B(n2162), .Y(n2228));
  OAI21X1 g1191(.A0(n2153), .A1(n2149), .B0(n2172), .Y(n2229));
  XOR2X1  g1192(.A(n2222), .B(n2208), .Y(n2235));
  NOR2X1  g1193(.A(n2235), .B(n2324), .Y(n2236));
  AOI21X1 g1194(.A0(n2324), .A1(n2235), .B0(n2236), .Y(n2237));
  AOI21X1 g1195(.A0(n2217), .A1(n2216), .B0(n2237), .Y(n2238));
  INVX1   g1196(.A(n2047), .Y(n2239));
  NAND3X1 g1197(.A(n2172), .B(n2166), .C(n2165), .Y(n2240));
  NAND2X1 g1198(.A(n2240), .B(n2188), .Y(n2241));
  NOR2X1  g1199(.A(n2241), .B(n2134), .Y(n2242));
  OAI21X1 g1200(.A0(n2167), .A1(n2185), .B0(n2173), .Y(n2243));
  OAI21X1 g1201(.A0(n2154), .A1(n2192), .B0(n2243), .Y(n2244));
  NOR2X1  g1202(.A(n2244), .B(n2242), .Y(n2245));
  XOR2X1  g1203(.A(n2245), .B(n2224), .Y(n2246));
  OAI22X1 g1204(.A0(n2237), .A1(n2239), .B0(n2196), .B1(n2246), .Y(n2247));
  INVX1   g1205(.A(n2246), .Y(n2248));
  AOI22X1 g1206(.A0(n2167), .A1(n2093), .B0(n2045), .B1(n2248), .Y(n2249));
  OAI21X1 g1207(.A0(n2044), .A1(n2028), .B0(n2248), .Y(n2250));
  NAND2X1 g1208(.A(n2250), .B(n2249), .Y(n2251));
  NAND2X1 g1209(.A(n2173), .B(n2200), .Y(n2252));
  XOR2X1  g1210(.A(n2222), .B(n2252), .Y(n2253));
  INVX1   g1211(.A(P1_REG2_REG_5__SCAN_IN), .Y(n2254));
  NAND2X1 g1212(.A(n2105), .B(P1_REG0_REG_5__SCAN_IN), .Y(n2255));
  OAI21X1 g1213(.A0(n2147), .A1(n2254), .B0(n2255), .Y(n2256));
  NAND3X1 g1214(.A(n2016), .B(n2020), .C(P1_REG1_REG_5__SCAN_IN), .Y(n2257));
  NAND2X1 g1215(.A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), .Y(n2258));
  XOR2X1  g1216(.A(n2258), .B(P1_REG3_REG_5__SCAN_IN), .Y(n2259));
  INVX1   g1217(.A(n2259), .Y(n2260));
  NAND3X1 g1218(.A(n2260), .B(n2016), .C(n2014), .Y(n2261));
  NAND2X1 g1219(.A(n2261), .B(n2257), .Y(n2262));
  NOR2X1  g1220(.A(n2262), .B(n2256), .Y(n2263));
  OAI22X1 g1221(.A0(n2223), .A1(n2068), .B0(n2104), .B1(n2263), .Y(n2264));
  AOI21X1 g1222(.A0(n2253), .A1(n2063), .B0(n2264), .Y(n2265));
  OAI21X1 g1223(.A0(n2237), .A1(n2053), .B0(n2265), .Y(n2266));
  NOR4X1  g1224(.A(n2251), .B(n2247), .C(n2238), .D(n2266), .Y(n2267));
  NAND2X1 g1225(.A(n2000), .B(P1_REG0_REG_4__SCAN_IN), .Y(n2268));
  OAI21X1 g1226(.A0(n2267), .A1(n2000), .B0(n2268), .Y(P1_U3466));
  INVX1   g1227(.A(n2324), .Y(n2270));
  INVX1   g1228(.A(n2202), .Y(n2271));
  OAI21X1 g1229(.A0(n2206), .A1(n2271), .B0(n2222), .Y(n2272));
  INVX1   g1230(.A(n2272), .Y(n2273));
  INVX1   g1231(.A(n2263), .Y(n2274));
  NOR2X1  g1232(.A(P1_IR_REG_31__SCAN_IN), .B(n1290), .Y(n2275));
  AOI21X1 g1233(.A0(n1261), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2275), .Y(n2276));
  NOR4X1  g1234(.A(n2004), .B(n2003), .C(n2002), .D(n2276), .Y(n2277));
  INVX1   g1235(.A(n2277), .Y(n2278));
  OAI21X1 g1236(.A0(n2005), .A1(n1258), .B0(n2278), .Y(n2279));
  OAI22X1 g1237(.A0(n2274), .A1(n2279), .B0(n2222), .B1(n2208), .Y(n2280));
  AOI21X1 g1238(.A0(n2279), .A1(n2274), .B0(n2280), .Y(n2281));
  OAI21X1 g1239(.A0(n2273), .A1(n2270), .B0(n2281), .Y(n2282));
  AOI21X1 g1240(.A0(n2223), .A1(n2209), .B0(n2324), .Y(n2283));
  INVX1   g1241(.A(n2279), .Y(n2284));
  NOR2X1  g1242(.A(n2284), .B(n2274), .Y(n2285));
  NOR2X1  g1243(.A(n2279), .B(n2263), .Y(n2286));
  NOR3X1  g1244(.A(n2286), .B(n2285), .C(n2273), .Y(n2287));
  INVX1   g1245(.A(n2287), .Y(n2288));
  OAI21X1 g1246(.A0(n2288), .A1(n2283), .B0(n2282), .Y(n2289));
  INVX1   g1247(.A(n2289), .Y(n2290));
  AOI22X1 g1248(.A0(n2208), .A1(n2093), .B0(n2047), .B1(n2290), .Y(n2291));
  OAI21X1 g1249(.A0(n2049), .A1(n2042), .B0(n2290), .Y(n2292));
  XOR2X1  g1250(.A(n2279), .B(n2263), .Y(n2293));
  AOI21X1 g1251(.A0(n2207), .A1(n2202), .B0(n2222), .Y(n2294));
  NOR2X1  g1252(.A(n2223), .B(n2208), .Y(n2295));
  NAND3X1 g1253(.A(n2240), .B(n2187), .C(n2188), .Y(n2296));
  AOI21X1 g1254(.A0(n2154), .A1(n2192), .B0(n2172), .Y(n2297));
  AOI21X1 g1255(.A0(n2167), .A1(n2185), .B0(n2297), .Y(n2298));
  AOI21X1 g1256(.A0(n2298), .A1(n2296), .B0(n2295), .Y(n2299));
  NOR2X1  g1257(.A(n2299), .B(n2294), .Y(n2300));
  XOR2X1  g1258(.A(n2300), .B(n2293), .Y(n2301));
  INVX1   g1259(.A(n2301), .Y(n2302));
  OAI21X1 g1260(.A0(n2045), .A1(n2044), .B0(n2302), .Y(n2303));
  OAI21X1 g1261(.A0(n2038), .A1(n2028), .B0(n2302), .Y(n2304));
  NAND4X1 g1262(.A(n2303), .B(n2292), .C(n2291), .D(n2304), .Y(n2305));
  NOR2X1  g1263(.A(n2289), .B(n2053), .Y(n2306));
  NOR2X1  g1264(.A(n2222), .B(n2252), .Y(n2307));
  XOR2X1  g1265(.A(n2279), .B(n2307), .Y(n2308));
  INVX1   g1266(.A(n2068), .Y(n2309));
  AOI22X1 g1267(.A0(n2105), .A1(P1_REG0_REG_6__SCAN_IN), .B0(P1_REG2_REG_6__SCAN_IN), .B1(n2106), .Y(n2310));
  INVX1   g1268(.A(P1_REG1_REG_6__SCAN_IN), .Y(n2311));
  NAND3X1 g1269(.A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_5__SCAN_IN), .C(P1_REG3_REG_4__SCAN_IN), .Y(n2312));
  XOR2X1  g1270(.A(n2312), .B(P1_REG3_REG_6__SCAN_IN), .Y(n2313));
  OAI22X1 g1271(.A0(n2152), .A1(n2313), .B0(n2151), .B1(n2311), .Y(n2314));
  INVX1   g1272(.A(n2314), .Y(n2315));
  NAND2X1 g1273(.A(n2315), .B(n2310), .Y(n2316));
  AOI22X1 g1274(.A0(n2279), .A1(n2309), .B0(n2054), .B1(n2316), .Y(n2317));
  OAI21X1 g1275(.A0(n2308), .A1(n2064), .B0(n2317), .Y(n2318));
  NOR3X1  g1276(.A(n2318), .B(n2306), .C(n2305), .Y(n2319));
  NAND2X1 g1277(.A(n2000), .B(P1_REG0_REG_5__SCAN_IN), .Y(n2320));
  OAI21X1 g1278(.A0(n2319), .A1(n2000), .B0(n2320), .Y(P1_U3469));
  INVX1   g1279(.A(n2093), .Y(n2322));
  OAI21X1 g1280(.A0(n2227), .A1(n2161), .B0(n2229), .Y(n2323));
  AOI21X1 g1281(.A0(n2228), .A1(n2126), .B0(n2323), .Y(n2324));
  AOI21X1 g1282(.A0(n2284), .A1(n2272), .B0(n2263), .Y(n2325));
  AOI21X1 g1283(.A0(n2279), .A1(n2273), .B0(n2325), .Y(n2326));
  OAI21X1 g1284(.A0(n2324), .A1(n2280), .B0(n2326), .Y(n2327));
  NOR2X1  g1285(.A(P1_IR_REG_31__SCAN_IN), .B(n1292), .Y(n2328));
  AOI21X1 g1286(.A0(n1295), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2328), .Y(n2329));
  INVX1   g1287(.A(n2329), .Y(n2330));
  NOR2X1  g1288(.A(n2005), .B(n1289), .Y(n2331));
  AOI21X1 g1289(.A0(n2330), .A1(n2005), .B0(n2331), .Y(n2332));
  NOR2X1  g1290(.A(n2332), .B(n2316), .Y(n2333));
  INVX1   g1291(.A(n2333), .Y(n2334));
  INVX1   g1292(.A(P1_REG2_REG_6__SCAN_IN), .Y(n2335));
  NAND2X1 g1293(.A(n2105), .B(P1_REG0_REG_6__SCAN_IN), .Y(n2336));
  OAI21X1 g1294(.A0(n2147), .A1(n2335), .B0(n2336), .Y(n2337));
  NOR2X1  g1295(.A(n2314), .B(n2337), .Y(n2338));
  NAND2X1 g1296(.A(n2330), .B(n2005), .Y(n2339));
  OAI21X1 g1297(.A0(n2005), .A1(n1289), .B0(n2339), .Y(n2340));
  NOR2X1  g1298(.A(n2340), .B(n2338), .Y(n2341));
  INVX1   g1299(.A(n2341), .Y(n2342));
  AOI21X1 g1300(.A0(n2342), .A1(n2334), .B0(n2327), .Y(n2343));
  XOR2X1  g1301(.A(n2340), .B(n2338), .Y(n2344));
  AOI21X1 g1302(.A0(n2344), .A1(n2327), .B0(n2343), .Y(n2345));
  OAI22X1 g1303(.A0(n2263), .A1(n2322), .B0(n2239), .B1(n2345), .Y(n2346));
  AOI21X1 g1304(.A0(n2217), .A1(n2216), .B0(n2345), .Y(n2347));
  NOR3X1  g1305(.A(n2299), .B(n2286), .C(n2294), .Y(n2349));
  NOR3X1  g1306(.A(n2349), .B(n2344), .C(n2285), .Y(n2350));
  NOR2X1  g1307(.A(n2300), .B(n2285), .Y(n2351));
  NOR4X1  g1308(.A(n2341), .B(n2333), .C(n2286), .D(n2351), .Y(n2352));
  OAI22X1 g1309(.A0(n2350), .A1(n2352), .B0(n2045), .B1(n2044), .Y(n2353));
  OAI22X1 g1310(.A0(n2350), .A1(n2352), .B0(n2038), .B1(n2028), .Y(n2354));
  NAND2X1 g1311(.A(n2354), .B(n2353), .Y(n2355));
  NAND4X1 g1312(.A(n2223), .B(n2173), .C(n2200), .D(n2284), .Y(n2356));
  XOR2X1  g1313(.A(n2340), .B(n2356), .Y(n2357));
  AOI22X1 g1314(.A0(n2105), .A1(P1_REG0_REG_7__SCAN_IN), .B0(P1_REG2_REG_7__SCAN_IN), .B1(n2106), .Y(n2358));
  INVX1   g1315(.A(n2151), .Y(n2359));
  INVX1   g1316(.A(n2152), .Y(n2360));
  NAND4X1 g1317(.A(P1_REG3_REG_5__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), .C(P1_REG3_REG_6__SCAN_IN), .D(P1_REG3_REG_3__SCAN_IN), .Y(n2361));
  XOR2X1  g1318(.A(n2361), .B(P1_REG3_REG_7__SCAN_IN), .Y(n2362));
  INVX1   g1319(.A(n2362), .Y(n2363));
  AOI22X1 g1320(.A0(n2360), .A1(n2363), .B0(n2359), .B1(P1_REG1_REG_7__SCAN_IN), .Y(n2364));
  NAND2X1 g1321(.A(n2364), .B(n2358), .Y(n2365));
  INVX1   g1322(.A(n2365), .Y(n2366));
  OAI22X1 g1323(.A0(n2332), .A1(n2068), .B0(n2104), .B1(n2366), .Y(n2367));
  AOI21X1 g1324(.A0(n2357), .A1(n2063), .B0(n2367), .Y(n2368));
  OAI21X1 g1325(.A0(n2345), .A1(n2053), .B0(n2368), .Y(n2369));
  NOR4X1  g1326(.A(n2355), .B(n2347), .C(n2346), .D(n2369), .Y(n2370));
  NAND2X1 g1327(.A(n2000), .B(P1_REG0_REG_6__SCAN_IN), .Y(n2371));
  OAI21X1 g1328(.A0(n2370), .A1(n2000), .B0(n2371), .Y(P1_U3472));
  NOR2X1  g1329(.A(n2332), .B(n2338), .Y(n2373));
  NOR2X1  g1330(.A(n2373), .B(n2327), .Y(n2374));
  NOR2X1  g1331(.A(P1_IR_REG_31__SCAN_IN), .B(n1318), .Y(n2375));
  AOI21X1 g1332(.A0(n1319), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2375), .Y(n2376));
  INVX1   g1333(.A(n2376), .Y(n2377));
  NOR2X1  g1334(.A(n2005), .B(n1317), .Y(n2378));
  AOI21X1 g1335(.A0(n2377), .A1(n2005), .B0(n2378), .Y(n2379));
  AOI22X1 g1336(.A0(n2366), .A1(n2379), .B0(n2332), .B1(n2338), .Y(n2380));
  OAI21X1 g1337(.A0(n2379), .A1(n2366), .B0(n2380), .Y(n2381));
  NAND2X1 g1338(.A(n2340), .B(n2316), .Y(n2382));
  OAI21X1 g1339(.A0(n2340), .A1(n2316), .B0(n2327), .Y(n2383));
  NAND2X1 g1340(.A(n2377), .B(n2005), .Y(n2384));
  OAI21X1 g1341(.A0(n2005), .A1(n1317), .B0(n2384), .Y(n2385));
  XOR2X1  g1342(.A(n2385), .B(n2366), .Y(n2386));
  NAND3X1 g1343(.A(n2386), .B(n2383), .C(n2382), .Y(n2387));
  OAI21X1 g1344(.A0(n2381), .A1(n2374), .B0(n2387), .Y(n2388));
  OAI22X1 g1345(.A0(n2338), .A1(n2322), .B0(n2239), .B1(n2388), .Y(n2389));
  AOI21X1 g1346(.A0(n2217), .A1(n2216), .B0(n2388), .Y(n2390));
  AOI22X1 g1347(.A0(n2338), .A1(n2340), .B0(n2279), .B1(n2263), .Y(n2391));
  NOR2X1  g1348(.A(n2341), .B(n2286), .Y(n2392));
  NAND2X1 g1349(.A(n2391), .B(n2294), .Y(n2393));
  AOI21X1 g1350(.A0(n2393), .A1(n2392), .B0(n2333), .Y(n2394));
  AOI21X1 g1351(.A0(n2391), .A1(n2299), .B0(n2394), .Y(n2395));
  XOR2X1  g1352(.A(n2395), .B(n2386), .Y(n2396));
  INVX1   g1353(.A(n2396), .Y(n2397));
  OAI21X1 g1354(.A0(n2045), .A1(n2044), .B0(n2397), .Y(n2398));
  OAI21X1 g1355(.A0(n2038), .A1(n2028), .B0(n2397), .Y(n2399));
  NAND2X1 g1356(.A(n2399), .B(n2398), .Y(n2400));
  NAND3X1 g1357(.A(n2332), .B(n2284), .C(n2307), .Y(n2401));
  XOR2X1  g1358(.A(n2385), .B(n2401), .Y(n2402));
  AOI22X1 g1359(.A0(n2105), .A1(P1_REG0_REG_8__SCAN_IN), .B0(P1_REG2_REG_8__SCAN_IN), .B1(n2106), .Y(n2403));
  INVX1   g1360(.A(P1_REG3_REG_8__SCAN_IN), .Y(n2404));
  INVX1   g1361(.A(P1_REG3_REG_7__SCAN_IN), .Y(n2405));
  NOR2X1  g1362(.A(n2361), .B(n2405), .Y(n2406));
  XOR2X1  g1363(.A(n2406), .B(n2404), .Y(n2407));
  INVX1   g1364(.A(n2407), .Y(n2408));
  AOI22X1 g1365(.A0(n2360), .A1(n2408), .B0(n2359), .B1(P1_REG1_REG_8__SCAN_IN), .Y(n2409));
  NAND2X1 g1366(.A(n2409), .B(n2403), .Y(n2410));
  INVX1   g1367(.A(n2410), .Y(n2411));
  OAI22X1 g1368(.A0(n2379), .A1(n2068), .B0(n2104), .B1(n2411), .Y(n2412));
  AOI21X1 g1369(.A0(n2402), .A1(n2063), .B0(n2412), .Y(n2413));
  OAI21X1 g1370(.A0(n2388), .A1(n2053), .B0(n2413), .Y(n2414));
  NOR4X1  g1371(.A(n2400), .B(n2390), .C(n2389), .D(n2414), .Y(n2415));
  NAND2X1 g1372(.A(n2000), .B(P1_REG0_REG_7__SCAN_IN), .Y(n2416));
  OAI21X1 g1373(.A0(n2415), .A1(n2000), .B0(n2416), .Y(P1_U3475));
  OAI21X1 g1374(.A0(n2385), .A1(n2373), .B0(n2365), .Y(n2418));
  OAI21X1 g1375(.A0(n2379), .A1(n2382), .B0(n2418), .Y(n2419));
  AOI21X1 g1376(.A0(n2380), .A1(n2327), .B0(n2419), .Y(n2420));
  NOR2X1  g1377(.A(P1_IR_REG_31__SCAN_IN), .B(n1341), .Y(n2421));
  AOI21X1 g1378(.A0(n1345), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2421), .Y(n2422));
  INVX1   g1379(.A(n2422), .Y(n2423));
  NAND2X1 g1380(.A(n2423), .B(n2005), .Y(n2424));
  OAI21X1 g1381(.A0(n2005), .A1(n1338), .B0(n2424), .Y(n2425));
  XOR2X1  g1382(.A(n2425), .B(n2411), .Y(n2426));
  XOR2X1  g1383(.A(n2425), .B(n2410), .Y(n2428));
  NOR2X1  g1384(.A(n2428), .B(n2420), .Y(n2429));
  AOI21X1 g1385(.A0(n2428), .A1(n2420), .B0(n2429), .Y(n2430));
  OAI22X1 g1386(.A0(n2366), .A1(n2322), .B0(n2239), .B1(n2430), .Y(n2431));
  AOI21X1 g1387(.A0(n2217), .A1(n2216), .B0(n2430), .Y(n2432));
  AOI21X1 g1388(.A0(n2364), .A1(n2358), .B0(n2385), .Y(n2433));
  INVX1   g1389(.A(n2395), .Y(n2434));
  NOR2X1  g1390(.A(n2379), .B(n2365), .Y(n2435));
  NOR2X1  g1391(.A(n2426), .B(n2435), .Y(n2436));
  OAI21X1 g1392(.A0(n2434), .A1(n2433), .B0(n2436), .Y(n2437));
  NOR2X1  g1393(.A(n2428), .B(n2433), .Y(n2438));
  OAI21X1 g1394(.A0(n2395), .A1(n2435), .B0(n2438), .Y(n2439));
  NAND2X1 g1395(.A(n2439), .B(n2437), .Y(n2440));
  OAI21X1 g1396(.A0(n2045), .A1(n2044), .B0(n2440), .Y(n2441));
  OAI21X1 g1397(.A0(n2038), .A1(n2028), .B0(n2440), .Y(n2442));
  NAND2X1 g1398(.A(n2442), .B(n2441), .Y(n2443));
  NOR3X1  g1399(.A(n2385), .B(n2340), .C(n2356), .Y(n2444));
  INVX1   g1400(.A(n2425), .Y(n2445));
  XOR2X1  g1401(.A(n2445), .B(n2444), .Y(n2446));
  INVX1   g1402(.A(P1_REG3_REG_9__SCAN_IN), .Y(n2447));
  NOR3X1  g1403(.A(n2361), .B(n2405), .C(n2404), .Y(n2448));
  XOR2X1  g1404(.A(n2448), .B(n2447), .Y(n2449));
  INVX1   g1405(.A(n2449), .Y(n2450));
  AOI22X1 g1406(.A0(n2360), .A1(n2450), .B0(n2105), .B1(P1_REG0_REG_9__SCAN_IN), .Y(n2451));
  AOI22X1 g1407(.A0(n2106), .A1(P1_REG2_REG_9__SCAN_IN), .B0(P1_REG1_REG_9__SCAN_IN), .B1(n2359), .Y(n2452));
  NAND2X1 g1408(.A(n2452), .B(n2451), .Y(n2453));
  INVX1   g1409(.A(n2453), .Y(n2454));
  OAI22X1 g1410(.A0(n2445), .A1(n2068), .B0(n2104), .B1(n2454), .Y(n2455));
  AOI21X1 g1411(.A0(n2446), .A1(n2063), .B0(n2455), .Y(n2456));
  OAI21X1 g1412(.A0(n2430), .A1(n2053), .B0(n2456), .Y(n2457));
  NOR4X1  g1413(.A(n2443), .B(n2432), .C(n2431), .D(n2457), .Y(n2458));
  NAND2X1 g1414(.A(n2000), .B(P1_REG0_REG_8__SCAN_IN), .Y(n2459));
  OAI21X1 g1415(.A0(n2458), .A1(n2000), .B0(n2459), .Y(P1_U3478));
  NOR2X1  g1416(.A(n2425), .B(n2410), .Y(n2461));
  NOR2X1  g1417(.A(n2445), .B(n2411), .Y(n2462));
  INVX1   g1418(.A(n2462), .Y(n2463));
  OAI21X1 g1419(.A0(n2461), .A1(n2420), .B0(n2463), .Y(n2464));
  NOR2X1  g1420(.A(P1_IR_REG_31__SCAN_IN), .B(n1383), .Y(n2465));
  AOI21X1 g1421(.A0(n1364), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2465), .Y(n2466));
  INVX1   g1422(.A(n2466), .Y(n2467));
  NAND2X1 g1423(.A(n2467), .B(n2005), .Y(n2468));
  OAI21X1 g1424(.A0(n2005), .A1(n1363), .B0(n2468), .Y(n2469));
  XOR2X1  g1425(.A(n2469), .B(n2454), .Y(n2470));
  NOR2X1  g1426(.A(n2464), .B(n2470), .Y(n2471));
  AOI21X1 g1427(.A0(n2470), .A1(n2464), .B0(n2471), .Y(n2473));
  INVX1   g1428(.A(n2473), .Y(n2474));
  OAI21X1 g1429(.A0(n2049), .A1(n2042), .B0(n2474), .Y(n2475));
  AOI22X1 g1430(.A0(n2411), .A1(n2425), .B0(n2385), .B1(n2366), .Y(n2476));
  INVX1   g1431(.A(n2476), .Y(n2477));
  NOR2X1  g1432(.A(n2477), .B(n2395), .Y(n2478));
  OAI21X1 g1433(.A0(n2410), .A1(n2433), .B0(n2445), .Y(n2479));
  NAND2X1 g1434(.A(n2410), .B(n2433), .Y(n2480));
  NAND2X1 g1435(.A(n2480), .B(n2479), .Y(n2481));
  NOR2X1  g1436(.A(n2481), .B(n2478), .Y(n2482));
  XOR2X1  g1437(.A(n2482), .B(n2470), .Y(n2483));
  INVX1   g1438(.A(n2483), .Y(n2484));
  AOI22X1 g1439(.A0(n2474), .A1(n2047), .B0(n2038), .B1(n2484), .Y(n2485));
  AOI22X1 g1440(.A0(n2410), .A1(n2093), .B0(n2045), .B1(n2484), .Y(n2486));
  OAI21X1 g1441(.A0(n2044), .A1(n2028), .B0(n2484), .Y(n2487));
  NAND4X1 g1442(.A(n2486), .B(n2485), .C(n2475), .D(n2487), .Y(n2488));
  NAND2X1 g1443(.A(n2445), .B(n2444), .Y(n2489));
  XOR2X1  g1444(.A(n2469), .B(n2489), .Y(n2490));
  INVX1   g1445(.A(n2469), .Y(n2491));
  INVX1   g1446(.A(P1_REG3_REG_10__SCAN_IN), .Y(n2492));
  NOR4X1  g1447(.A(n2405), .B(n2404), .C(n2447), .D(n2361), .Y(n2493));
  XOR2X1  g1448(.A(n2493), .B(n2492), .Y(n2494));
  INVX1   g1449(.A(n2494), .Y(n2495));
  AOI22X1 g1450(.A0(n2360), .A1(n2495), .B0(n2105), .B1(P1_REG0_REG_10__SCAN_IN), .Y(n2496));
  AOI22X1 g1451(.A0(n2106), .A1(P1_REG2_REG_10__SCAN_IN), .B0(P1_REG1_REG_10__SCAN_IN), .B1(n2359), .Y(n2497));
  NAND2X1 g1452(.A(n2497), .B(n2496), .Y(n2498));
  INVX1   g1453(.A(n2498), .Y(n2499));
  OAI22X1 g1454(.A0(n2491), .A1(n2068), .B0(n2104), .B1(n2499), .Y(n2500));
  AOI21X1 g1455(.A0(n2490), .A1(n2063), .B0(n2500), .Y(n2501));
  OAI21X1 g1456(.A0(n2473), .A1(n2053), .B0(n2501), .Y(n2502));
  NOR2X1  g1457(.A(n2502), .B(n2488), .Y(n2503));
  NAND2X1 g1458(.A(n2000), .B(P1_REG0_REG_9__SCAN_IN), .Y(n2504));
  OAI21X1 g1459(.A0(n2503), .A1(n2000), .B0(n2504), .Y(P1_U3481));
  AOI21X1 g1460(.A0(n2469), .A1(n2453), .B0(n2464), .Y(n2506));
  NOR2X1  g1461(.A(P1_IR_REG_31__SCAN_IN), .B(n1384), .Y(n2507));
  AOI21X1 g1462(.A0(n1389), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2507), .Y(n2508));
  INVX1   g1463(.A(n2508), .Y(n2509));
  NAND2X1 g1464(.A(n2509), .B(n2005), .Y(n2510));
  OAI21X1 g1465(.A0(n2005), .A1(n1382), .B0(n2510), .Y(n2511));
  INVX1   g1466(.A(n2511), .Y(n2512));
  NOR2X1  g1467(.A(n2512), .B(n2499), .Y(n2513));
  NOR2X1  g1468(.A(n2511), .B(n2498), .Y(n2514));
  AOI21X1 g1469(.A0(n2491), .A1(n2454), .B0(n2514), .Y(n2515));
  INVX1   g1470(.A(n2515), .Y(n2516));
  NOR3X1  g1471(.A(n2516), .B(n2513), .C(n2506), .Y(n2517));
  OAI21X1 g1472(.A0(n2469), .A1(n2453), .B0(n2464), .Y(n2518));
  XOR2X1  g1473(.A(n2511), .B(n2499), .Y(n2519));
  INVX1   g1474(.A(n2519), .Y(n2520));
  AOI21X1 g1475(.A0(n2469), .A1(n2453), .B0(n2520), .Y(n2521));
  AOI21X1 g1476(.A0(n2521), .A1(n2518), .B0(n2517), .Y(n2522));
  INVX1   g1477(.A(n2522), .Y(n2523));
  OAI22X1 g1478(.A0(n2454), .A1(n2322), .B0(n2239), .B1(n2523), .Y(n2524));
  AOI21X1 g1479(.A0(n2217), .A1(n2216), .B0(n2523), .Y(n2525));
  NOR2X1  g1480(.A(n2491), .B(n2453), .Y(n2526));
  NOR2X1  g1481(.A(n2469), .B(n2454), .Y(n2527));
  INVX1   g1482(.A(n2527), .Y(n2528));
  OAI21X1 g1483(.A0(n2482), .A1(n2526), .B0(n2528), .Y(n2529));
  XOR2X1  g1484(.A(n2529), .B(n2520), .Y(n2530));
  INVX1   g1485(.A(n2530), .Y(n2531));
  OAI21X1 g1486(.A0(n2045), .A1(n2044), .B0(n2531), .Y(n2532));
  OAI21X1 g1487(.A0(n2038), .A1(n2028), .B0(n2531), .Y(n2533));
  NAND2X1 g1488(.A(n2533), .B(n2532), .Y(n2534));
  NOR4X1  g1489(.A(n2425), .B(n2385), .C(n2401), .D(n2469), .Y(n2535));
  NOR2X1  g1490(.A(n2512), .B(n2535), .Y(n2536));
  NOR3X1  g1491(.A(n2511), .B(n2469), .C(n2489), .Y(n2537));
  NOR2X1  g1492(.A(n2537), .B(n2536), .Y(n2538));
  NAND2X1 g1493(.A(n2493), .B(P1_REG3_REG_10__SCAN_IN), .Y(n2539));
  XOR2X1  g1494(.A(n2539), .B(P1_REG3_REG_11__SCAN_IN), .Y(n2540));
  INVX1   g1495(.A(n2540), .Y(n2541));
  NAND3X1 g1496(.A(n2541), .B(n2016), .C(n2014), .Y(n2542));
  NAND2X1 g1497(.A(n2105), .B(P1_REG0_REG_11__SCAN_IN), .Y(n2543));
  AOI22X1 g1498(.A0(n2106), .A1(P1_REG2_REG_11__SCAN_IN), .B0(P1_REG1_REG_11__SCAN_IN), .B1(n2359), .Y(n2544));
  NAND3X1 g1499(.A(n2544), .B(n2543), .C(n2542), .Y(n2545));
  INVX1   g1500(.A(n2545), .Y(n2546));
  OAI22X1 g1501(.A0(n2512), .A1(n2068), .B0(n2104), .B1(n2546), .Y(n2547));
  AOI21X1 g1502(.A0(n2538), .A1(n2063), .B0(n2547), .Y(n2548));
  OAI21X1 g1503(.A0(n2523), .A1(n2053), .B0(n2548), .Y(n2549));
  NOR4X1  g1504(.A(n2534), .B(n2525), .C(n2524), .D(n2549), .Y(n2550));
  NAND2X1 g1505(.A(n2000), .B(P1_REG0_REG_10__SCAN_IN), .Y(n2551));
  OAI21X1 g1506(.A0(n2550), .A1(n2000), .B0(n2551), .Y(P1_U3484));
  NOR2X1  g1507(.A(n2511), .B(n2499), .Y(n2553));
  NOR2X1  g1508(.A(n2529), .B(n2553), .Y(n2554));
  INVX1   g1509(.A(n2554), .Y(n2555));
  NAND2X1 g1510(.A(n2511), .B(n2499), .Y(n2556));
  INVX1   g1511(.A(n2556), .Y(n2557));
  NOR2X1  g1512(.A(P1_IR_REG_31__SCAN_IN), .B(n1409), .Y(n2558));
  AOI21X1 g1513(.A0(n1410), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2558), .Y(n2559));
  INVX1   g1514(.A(n2559), .Y(n2560));
  NAND2X1 g1515(.A(n2560), .B(n2005), .Y(n2561));
  OAI21X1 g1516(.A0(n2005), .A1(n1408), .B0(n2561), .Y(n2562));
  NAND2X1 g1517(.A(n2562), .B(n2546), .Y(n2563));
  NOR2X1  g1518(.A(n2562), .B(n2546), .Y(n2564));
  INVX1   g1519(.A(n2564), .Y(n2565));
  AOI21X1 g1520(.A0(n2565), .A1(n2563), .B0(n2557), .Y(n2566));
  NAND2X1 g1521(.A(n2529), .B(n2556), .Y(n2567));
  INVX1   g1522(.A(n2563), .Y(n2568));
  NOR3X1  g1523(.A(n2564), .B(n2568), .C(n2553), .Y(n2569));
  AOI22X1 g1524(.A0(n2567), .A1(n2569), .B0(n2566), .B1(n2555), .Y(n2570));
  OAI22X1 g1525(.A0(n2499), .A1(n2512), .B0(n2491), .B1(n2454), .Y(n2571));
  AOI21X1 g1526(.A0(n2515), .A1(n2462), .B0(n2571), .Y(n2572));
  OAI21X1 g1527(.A0(n2425), .A1(n2410), .B0(n2515), .Y(n2573));
  OAI22X1 g1528(.A0(n2572), .A1(n2514), .B0(n2420), .B1(n2573), .Y(n2574));
  AOI21X1 g1529(.A0(n2565), .A1(n2563), .B0(n2574), .Y(n2575));
  XOR2X1  g1530(.A(n2562), .B(n2545), .Y(n2576));
  INVX1   g1531(.A(n2576), .Y(n2577));
  AOI21X1 g1532(.A0(n2577), .A1(n2574), .B0(n2575), .Y(n2578));
  OAI22X1 g1533(.A0(n2499), .A1(n2322), .B0(n2239), .B1(n2578), .Y(n2579));
  NOR2X1  g1534(.A(n2578), .B(n2217), .Y(n2580));
  NOR2X1  g1535(.A(n2578), .B(n2216), .Y(n2581));
  NOR3X1  g1536(.A(n2581), .B(n2580), .C(n2579), .Y(n2582));
  OAI21X1 g1537(.A0(n2570), .A1(n2184), .B0(n2582), .Y(n2583));
  NOR2X1  g1538(.A(n2570), .B(n2196), .Y(n2584));
  AOI21X1 g1539(.A0(n2183), .A1(n2029), .B0(n2570), .Y(n2585));
  INVX1   g1540(.A(n2562), .Y(n2586));
  XOR2X1  g1541(.A(n2586), .B(n2537), .Y(n2587));
  NAND3X1 g1542(.A(n2493), .B(P1_REG3_REG_10__SCAN_IN), .C(P1_REG3_REG_11__SCAN_IN), .Y(n2588));
  XOR2X1  g1543(.A(n2588), .B(P1_REG3_REG_12__SCAN_IN), .Y(n2589));
  INVX1   g1544(.A(n2589), .Y(n2590));
  AOI22X1 g1545(.A0(n2360), .A1(n2590), .B0(n2105), .B1(P1_REG0_REG_12__SCAN_IN), .Y(n2591));
  AOI22X1 g1546(.A0(n2106), .A1(P1_REG2_REG_12__SCAN_IN), .B0(P1_REG1_REG_12__SCAN_IN), .B1(n2359), .Y(n2592));
  NAND2X1 g1547(.A(n2592), .B(n2591), .Y(n2593));
  INVX1   g1548(.A(n2593), .Y(n2594));
  OAI22X1 g1549(.A0(n2586), .A1(n2068), .B0(n2104), .B1(n2594), .Y(n2595));
  AOI21X1 g1550(.A0(n2587), .A1(n2063), .B0(n2595), .Y(n2596));
  OAI21X1 g1551(.A0(n2578), .A1(n2053), .B0(n2596), .Y(n2597));
  NOR4X1  g1552(.A(n2585), .B(n2584), .C(n2583), .D(n2597), .Y(n2598));
  NAND2X1 g1553(.A(n2000), .B(P1_REG0_REG_11__SCAN_IN), .Y(n2599));
  OAI21X1 g1554(.A0(n2598), .A1(n2000), .B0(n2599), .Y(P1_U3487));
  OAI21X1 g1555(.A0(n2562), .A1(n2545), .B0(n2574), .Y(n2601));
  OAI21X1 g1556(.A0(n2586), .A1(n2546), .B0(n2601), .Y(n2602));
  NOR2X1  g1557(.A(P1_IR_REG_31__SCAN_IN), .B(n1427), .Y(n2603));
  AOI21X1 g1558(.A0(n1430), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2603), .Y(n2604));
  INVX1   g1559(.A(n2604), .Y(n2605));
  NAND2X1 g1560(.A(n2605), .B(n2005), .Y(n2606));
  OAI21X1 g1561(.A0(n2005), .A1(n1426), .B0(n2606), .Y(n2607));
  XOR2X1  g1562(.A(n2607), .B(n2594), .Y(n2608));
  NOR2X1  g1563(.A(n2602), .B(n2608), .Y(n2609));
  AOI21X1 g1564(.A0(n2608), .A1(n2602), .B0(n2609), .Y(n2611));
  INVX1   g1565(.A(n2611), .Y(n2612));
  OAI21X1 g1566(.A0(n2049), .A1(n2042), .B0(n2612), .Y(n2613));
  NOR2X1  g1567(.A(n2564), .B(n2553), .Y(n2614));
  NAND3X1 g1568(.A(n2563), .B(n2556), .C(n2527), .Y(n2615));
  AOI21X1 g1569(.A0(n2615), .A1(n2614), .B0(n2568), .Y(n2616));
  INVX1   g1570(.A(n2616), .Y(n2617));
  NOR3X1  g1571(.A(n2568), .B(n2557), .C(n2526), .Y(n2618));
  OAI21X1 g1572(.A0(n2481), .A1(n2478), .B0(n2618), .Y(n2619));
  NAND2X1 g1573(.A(n2619), .B(n2617), .Y(n2620));
  XOR2X1  g1574(.A(n2620), .B(n2608), .Y(n2621));
  AOI22X1 g1575(.A0(n2612), .A1(n2047), .B0(n2038), .B1(n2621), .Y(n2622));
  AOI22X1 g1576(.A0(n2545), .A1(n2093), .B0(n2045), .B1(n2621), .Y(n2623));
  OAI21X1 g1577(.A0(n2044), .A1(n2028), .B0(n2621), .Y(n2624));
  NAND4X1 g1578(.A(n2623), .B(n2622), .C(n2613), .D(n2624), .Y(n2625));
  NOR4X1  g1579(.A(n2511), .B(n2469), .C(n2489), .D(n2562), .Y(n2626));
  INVX1   g1580(.A(n2607), .Y(n2627));
  XOR2X1  g1581(.A(n2627), .B(n2626), .Y(n2628));
  NAND4X1 g1582(.A(P1_REG3_REG_10__SCAN_IN), .B(P1_REG3_REG_12__SCAN_IN), .C(P1_REG3_REG_11__SCAN_IN), .D(n2493), .Y(n2629));
  XOR2X1  g1583(.A(n2629), .B(P1_REG3_REG_13__SCAN_IN), .Y(n2630));
  INVX1   g1584(.A(n2630), .Y(n2631));
  AOI22X1 g1585(.A0(n2360), .A1(n2631), .B0(n2105), .B1(P1_REG0_REG_13__SCAN_IN), .Y(n2632));
  AOI22X1 g1586(.A0(n2106), .A1(P1_REG2_REG_13__SCAN_IN), .B0(P1_REG1_REG_13__SCAN_IN), .B1(n2359), .Y(n2633));
  NAND2X1 g1587(.A(n2633), .B(n2632), .Y(n2634));
  INVX1   g1588(.A(n2634), .Y(n2635));
  OAI22X1 g1589(.A0(n2627), .A1(n2068), .B0(n2104), .B1(n2635), .Y(n2636));
  AOI21X1 g1590(.A0(n2628), .A1(n2063), .B0(n2636), .Y(n2637));
  OAI21X1 g1591(.A0(n2611), .A1(n2053), .B0(n2637), .Y(n2638));
  NOR2X1  g1592(.A(n2638), .B(n2625), .Y(n2639));
  NAND2X1 g1593(.A(n2000), .B(P1_REG0_REG_12__SCAN_IN), .Y(n2640));
  OAI21X1 g1594(.A0(n2639), .A1(n2000), .B0(n2640), .Y(P1_U3490));
  NOR2X1  g1595(.A(n2627), .B(n2594), .Y(n2642));
  NOR2X1  g1596(.A(n2642), .B(n2602), .Y(n2643));
  INVX1   g1597(.A(n2643), .Y(n2644));
  NOR2X1  g1598(.A(P1_IR_REG_31__SCAN_IN), .B(n1447), .Y(n2645));
  AOI21X1 g1599(.A0(n1448), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2645), .Y(n2646));
  INVX1   g1600(.A(n2646), .Y(n2647));
  NAND2X1 g1601(.A(n2647), .B(n2005), .Y(n2648));
  OAI21X1 g1602(.A0(n2005), .A1(n1446), .B0(n2648), .Y(n2649));
  OAI22X1 g1603(.A0(n2634), .A1(n2649), .B0(n2607), .B1(n2593), .Y(n2650));
  AOI21X1 g1604(.A0(n2649), .A1(n2634), .B0(n2650), .Y(n2651));
  OAI21X1 g1605(.A0(n2607), .A1(n2593), .B0(n2602), .Y(n2652));
  INVX1   g1606(.A(n2649), .Y(n2653));
  NOR2X1  g1607(.A(n2653), .B(n2634), .Y(n2654));
  NOR2X1  g1608(.A(n2649), .B(n2635), .Y(n2655));
  NOR3X1  g1609(.A(n2655), .B(n2654), .C(n2642), .Y(n2656));
  AOI22X1 g1610(.A0(n2652), .A1(n2656), .B0(n2651), .B1(n2644), .Y(n2657));
  INVX1   g1611(.A(n2657), .Y(n2658));
  OAI22X1 g1612(.A0(n2594), .A1(n2322), .B0(n2239), .B1(n2658), .Y(n2659));
  AOI21X1 g1613(.A0(n2217), .A1(n2216), .B0(n2658), .Y(n2660));
  XOR2X1  g1614(.A(n2649), .B(n2635), .Y(n2661));
  NOR2X1  g1615(.A(n2607), .B(n2594), .Y(n2662));
  AOI22X1 g1616(.A0(n2617), .A1(n2619), .B0(n2607), .B1(n2594), .Y(n2663));
  NOR2X1  g1617(.A(n2663), .B(n2662), .Y(n2664));
  XOR2X1  g1618(.A(n2664), .B(n2661), .Y(n2665));
  INVX1   g1619(.A(n2665), .Y(n2666));
  OAI21X1 g1620(.A0(n2045), .A1(n2044), .B0(n2666), .Y(n2667));
  OAI21X1 g1621(.A0(n2038), .A1(n2028), .B0(n2666), .Y(n2668));
  NAND2X1 g1622(.A(n2668), .B(n2667), .Y(n2669));
  INVX1   g1623(.A(n2626), .Y(n2670));
  NOR2X1  g1624(.A(n2607), .B(n2670), .Y(n2671));
  XOR2X1  g1625(.A(n2653), .B(n2671), .Y(n2672));
  INVX1   g1626(.A(P1_REG3_REG_14__SCAN_IN), .Y(n2673));
  INVX1   g1627(.A(P1_REG3_REG_13__SCAN_IN), .Y(n2674));
  NOR2X1  g1628(.A(n2629), .B(n2674), .Y(n2675));
  XOR2X1  g1629(.A(n2675), .B(n2673), .Y(n2676));
  INVX1   g1630(.A(n2676), .Y(n2677));
  NAND3X1 g1631(.A(n2677), .B(n2016), .C(n2014), .Y(n2678));
  NAND3X1 g1632(.A(n2016), .B(n2020), .C(P1_REG1_REG_14__SCAN_IN), .Y(n2679));
  AOI22X1 g1633(.A0(n2105), .A1(P1_REG0_REG_14__SCAN_IN), .B0(P1_REG2_REG_14__SCAN_IN), .B1(n2106), .Y(n2680));
  NAND3X1 g1634(.A(n2680), .B(n2679), .C(n2678), .Y(n2681));
  INVX1   g1635(.A(n2681), .Y(n2682));
  OAI22X1 g1636(.A0(n2653), .A1(n2068), .B0(n2104), .B1(n2682), .Y(n2683));
  AOI21X1 g1637(.A0(n2672), .A1(n2063), .B0(n2683), .Y(n2684));
  OAI21X1 g1638(.A0(n2658), .A1(n2053), .B0(n2684), .Y(n2685));
  NOR4X1  g1639(.A(n2669), .B(n2660), .C(n2659), .D(n2685), .Y(n2686));
  NAND2X1 g1640(.A(n2000), .B(P1_REG0_REG_13__SCAN_IN), .Y(n2687));
  OAI21X1 g1641(.A0(n2686), .A1(n2000), .B0(n2687), .Y(P1_U3493));
  NOR2X1  g1642(.A(P1_IR_REG_31__SCAN_IN), .B(n1465), .Y(n2689));
  AOI21X1 g1643(.A0(n1469), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2689), .Y(n2690));
  INVX1   g1644(.A(n2690), .Y(n2691));
  NOR2X1  g1645(.A(n2005), .B(n1464), .Y(n2692));
  AOI21X1 g1646(.A0(n2691), .A1(n2005), .B0(n2692), .Y(n2693));
  XOR2X1  g1647(.A(n2693), .B(n2681), .Y(n2694));
  INVX1   g1648(.A(n2694), .Y(n2695));
  INVX1   g1649(.A(n2655), .Y(n2696));
  OAI22X1 g1650(.A0(n2653), .A1(n2634), .B0(n2662), .B1(n2663), .Y(n2697));
  NAND2X1 g1651(.A(n2697), .B(n2696), .Y(n2698));
  XOR2X1  g1652(.A(n2698), .B(n2695), .Y(n2699));
  NOR2X1  g1653(.A(n2699), .B(n2184), .Y(n2700));
  NOR3X1  g1654(.A(n2650), .B(n2586), .C(n2546), .Y(n2701));
  OAI22X1 g1655(.A0(n2635), .A1(n2653), .B0(n2627), .B1(n2594), .Y(n2702));
  OAI22X1 g1656(.A0(n2701), .A1(n2702), .B0(n2649), .B1(n2634), .Y(n2703));
  OAI21X1 g1657(.A0(n2650), .A1(n2601), .B0(n2703), .Y(n2704));
  XOR2X1  g1658(.A(n2704), .B(n2694), .Y(n2705));
  INVX1   g1659(.A(n2705), .Y(n2706));
  AOI22X1 g1660(.A0(n2634), .A1(n2093), .B0(n2047), .B1(n2706), .Y(n2707));
  OAI21X1 g1661(.A0(n2049), .A1(n2042), .B0(n2706), .Y(n2708));
  NAND2X1 g1662(.A(n2708), .B(n2707), .Y(n2709));
  NOR2X1  g1663(.A(n2699), .B(n2196), .Y(n2710));
  AOI21X1 g1664(.A0(n2183), .A1(n2029), .B0(n2699), .Y(n2711));
  NOR4X1  g1665(.A(n2710), .B(n2709), .C(n2700), .D(n2711), .Y(n2712));
  INVX1   g1666(.A(n2712), .Y(n2713));
  NOR2X1  g1667(.A(n2705), .B(n2053), .Y(n2714));
  NOR3X1  g1668(.A(n2649), .B(n2607), .C(n2670), .Y(n2715));
  NAND4X1 g1669(.A(n2653), .B(n2627), .C(n2626), .D(n2693), .Y(n2716));
  OAI21X1 g1670(.A0(n2693), .A1(n2715), .B0(n2716), .Y(n2717));
  INVX1   g1671(.A(n2693), .Y(n2718));
  INVX1   g1672(.A(P1_REG3_REG_15__SCAN_IN), .Y(n2719));
  NOR3X1  g1673(.A(n2629), .B(n2673), .C(n2674), .Y(n2720));
  XOR2X1  g1674(.A(n2720), .B(n2719), .Y(n2721));
  INVX1   g1675(.A(n2721), .Y(n2722));
  INVX1   g1676(.A(P1_REG1_REG_15__SCAN_IN), .Y(n2723));
  AOI22X1 g1677(.A0(n2105), .A1(P1_REG0_REG_15__SCAN_IN), .B0(P1_REG2_REG_15__SCAN_IN), .B1(n2106), .Y(n2724));
  OAI21X1 g1678(.A0(n2151), .A1(n2723), .B0(n2724), .Y(n2725));
  AOI21X1 g1679(.A0(n2722), .A1(n2360), .B0(n2725), .Y(n2726));
  INVX1   g1680(.A(n2726), .Y(n2727));
  AOI22X1 g1681(.A0(n2718), .A1(n2309), .B0(n2054), .B1(n2727), .Y(n2728));
  OAI21X1 g1682(.A0(n2717), .A1(n2064), .B0(n2728), .Y(n2729));
  NOR3X1  g1683(.A(n2729), .B(n2714), .C(n2713), .Y(n2730));
  NAND2X1 g1684(.A(n2000), .B(P1_REG0_REG_14__SCAN_IN), .Y(n2731));
  OAI21X1 g1685(.A0(n2730), .A1(n2000), .B0(n2731), .Y(P1_U3496));
  NOR2X1  g1686(.A(P1_IR_REG_31__SCAN_IN), .B(n1492), .Y(n2733));
  AOI21X1 g1687(.A0(n1493), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2733), .Y(n2734));
  INVX1   g1688(.A(n2734), .Y(n2735));
  NOR2X1  g1689(.A(n2005), .B(n1491), .Y(n2736));
  AOI21X1 g1690(.A0(n2735), .A1(n2005), .B0(n2736), .Y(n2737));
  XOR2X1  g1691(.A(n2737), .B(n2727), .Y(n2738));
  NOR2X1  g1692(.A(n2693), .B(n2681), .Y(n2739));
  INVX1   g1693(.A(n2739), .Y(n2740));
  NOR2X1  g1694(.A(n2718), .B(n2682), .Y(n2741));
  XOR2X1  g1695(.A(n4814), .B(n2738), .Y(n2743));
  NOR2X1  g1696(.A(n2743), .B(n2184), .Y(n2744));
  NOR2X1  g1697(.A(n2693), .B(n2682), .Y(n2745));
  NAND2X1 g1698(.A(n2693), .B(n2682), .Y(n2746));
  AOI21X1 g1699(.A0(n2746), .A1(n2704), .B0(n2745), .Y(n2747));
  XOR2X1  g1700(.A(n2747), .B(n2738), .Y(n2748));
  AOI22X1 g1701(.A0(n2681), .A1(n2093), .B0(n2047), .B1(n2748), .Y(n2749));
  OAI21X1 g1702(.A0(n2049), .A1(n2042), .B0(n2748), .Y(n2750));
  NAND2X1 g1703(.A(n2750), .B(n2749), .Y(n2751));
  NOR2X1  g1704(.A(n2743), .B(n2196), .Y(n2752));
  AOI21X1 g1705(.A0(n2183), .A1(n2029), .B0(n2743), .Y(n2753));
  NOR4X1  g1706(.A(n2752), .B(n2751), .C(n2744), .D(n2753), .Y(n2754));
  INVX1   g1707(.A(n2754), .Y(n2755));
  NAND2X1 g1708(.A(n2748), .B(n2052), .Y(n2756));
  INVX1   g1709(.A(n2737), .Y(n2757));
  XOR2X1  g1710(.A(n2757), .B(n2716), .Y(n2758));
  NOR4X1  g1711(.A(n2673), .B(n2674), .C(n2719), .D(n2629), .Y(n2759));
  XOR2X1  g1712(.A(n2759), .B(P1_REG3_REG_16__SCAN_IN), .Y(n2760));
  NAND3X1 g1713(.A(n2760), .B(n2016), .C(n2014), .Y(n2761));
  NAND3X1 g1714(.A(n2016), .B(n2020), .C(P1_REG1_REG_16__SCAN_IN), .Y(n2762));
  AOI22X1 g1715(.A0(n2105), .A1(P1_REG0_REG_16__SCAN_IN), .B0(P1_REG2_REG_16__SCAN_IN), .B1(n2106), .Y(n2763));
  NAND3X1 g1716(.A(n2763), .B(n2762), .C(n2761), .Y(n2764));
  INVX1   g1717(.A(n2764), .Y(n2765));
  OAI22X1 g1718(.A0(n2737), .A1(n2068), .B0(n2104), .B1(n2765), .Y(n2766));
  AOI21X1 g1719(.A0(n2758), .A1(n2063), .B0(n2766), .Y(n2767));
  NAND2X1 g1720(.A(n2767), .B(n2756), .Y(n2768));
  NOR2X1  g1721(.A(n2768), .B(n2755), .Y(n2769));
  NAND2X1 g1722(.A(n2000), .B(P1_REG0_REG_15__SCAN_IN), .Y(n2770));
  OAI21X1 g1723(.A0(n2769), .A1(n2000), .B0(n2770), .Y(P1_U3499));
  NOR2X1  g1724(.A(n2757), .B(n2726), .Y(n2772));
  INVX1   g1725(.A(n4814), .Y(n2773));
  NOR2X1  g1726(.A(n2737), .B(n2727), .Y(n2774));
  NOR2X1  g1727(.A(P1_IR_REG_31__SCAN_IN), .B(n1512), .Y(n2775));
  AOI21X1 g1728(.A0(n1525), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2775), .Y(n2776));
  INVX1   g1729(.A(n2776), .Y(n2777));
  NOR2X1  g1730(.A(n2005), .B(n1511), .Y(n2778));
  AOI21X1 g1731(.A0(n2777), .A1(n2005), .B0(n2778), .Y(n2779));
  XOR2X1  g1732(.A(n2779), .B(n2764), .Y(n2780));
  NOR2X1  g1733(.A(n2780), .B(n2774), .Y(n2781));
  OAI21X1 g1734(.A0(n2773), .A1(n2772), .B0(n2781), .Y(n2782));
  NOR2X1  g1735(.A(n2779), .B(n2764), .Y(n2783));
  INVX1   g1736(.A(n2779), .Y(n2784));
  OAI22X1 g1737(.A0(n2765), .A1(n2784), .B0(n2757), .B1(n2726), .Y(n2785));
  NOR2X1  g1738(.A(n2785), .B(n2783), .Y(n2786));
  OAI21X1 g1739(.A0(n4814), .A1(n2774), .B0(n2786), .Y(n2787));
  AOI21X1 g1740(.A0(n2787), .A1(n2782), .B0(n2184), .Y(n2788));
  INVX1   g1741(.A(n2788), .Y(n2789));
  NAND2X1 g1742(.A(n2757), .B(n2727), .Y(n2790));
  NOR2X1  g1743(.A(n2757), .B(n2727), .Y(n2791));
  OAI21X1 g1744(.A0(n2791), .A1(n2747), .B0(n2790), .Y(n2792));
  NOR2X1  g1745(.A(n2792), .B(n2780), .Y(n2793));
  XOR2X1  g1746(.A(n2779), .B(n2765), .Y(n2794));
  AOI21X1 g1747(.A0(n2780), .A1(n2792), .B0(n2793), .Y(n2796));
  INVX1   g1748(.A(n2796), .Y(n2797));
  AOI22X1 g1749(.A0(n2727), .A1(n2093), .B0(n2047), .B1(n2797), .Y(n2798));
  OAI21X1 g1750(.A0(n2049), .A1(n2042), .B0(n2797), .Y(n2799));
  NAND3X1 g1751(.A(n2799), .B(n2798), .C(n2789), .Y(n2800));
  AOI21X1 g1752(.A0(n2787), .A1(n2782), .B0(n2196), .Y(n2801));
  AOI22X1 g1753(.A0(n2782), .A1(n2787), .B0(n2183), .B1(n2029), .Y(n2802));
  NOR2X1  g1754(.A(n2757), .B(n2716), .Y(n2803));
  XOR2X1  g1755(.A(n2779), .B(n2803), .Y(n2804));
  NAND2X1 g1756(.A(n2759), .B(P1_REG3_REG_16__SCAN_IN), .Y(n2805));
  XOR2X1  g1757(.A(n2805), .B(P1_REG3_REG_17__SCAN_IN), .Y(n2806));
  INVX1   g1758(.A(n2806), .Y(n2807));
  NAND3X1 g1759(.A(n2807), .B(n2016), .C(n2014), .Y(n2808));
  NAND3X1 g1760(.A(n2016), .B(n2020), .C(P1_REG1_REG_17__SCAN_IN), .Y(n2809));
  AOI22X1 g1761(.A0(n2105), .A1(P1_REG0_REG_17__SCAN_IN), .B0(P1_REG2_REG_17__SCAN_IN), .B1(n2106), .Y(n2810));
  NAND3X1 g1762(.A(n2810), .B(n2809), .C(n2808), .Y(n2811));
  INVX1   g1763(.A(n2811), .Y(n2812));
  OAI22X1 g1764(.A0(n2779), .A1(n2068), .B0(n2104), .B1(n2812), .Y(n2813));
  AOI21X1 g1765(.A0(n2804), .A1(n2063), .B0(n2813), .Y(n2814));
  OAI21X1 g1766(.A0(n2796), .A1(n2053), .B0(n2814), .Y(n2815));
  NOR4X1  g1767(.A(n2802), .B(n2801), .C(n2800), .D(n2815), .Y(n2816));
  NAND2X1 g1768(.A(n2000), .B(P1_REG0_REG_16__SCAN_IN), .Y(n2817));
  OAI21X1 g1769(.A0(n2816), .A1(n2000), .B0(n2817), .Y(P1_U3502));
  NOR2X1  g1770(.A(n2779), .B(n2765), .Y(n2819));
  NOR2X1  g1771(.A(P1_IR_REG_31__SCAN_IN), .B(n1542), .Y(n2820));
  AOI21X1 g1772(.A0(n1543), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2820), .Y(n2821));
  INVX1   g1773(.A(n2821), .Y(n2822));
  NOR2X1  g1774(.A(n2005), .B(n1541), .Y(n2823));
  AOI21X1 g1775(.A0(n2822), .A1(n2005), .B0(n2823), .Y(n2824));
  INVX1   g1776(.A(n2824), .Y(n2825));
  AOI22X1 g1777(.A0(n2812), .A1(n2824), .B0(n2779), .B1(n2765), .Y(n2826));
  INVX1   g1778(.A(n2826), .Y(n2827));
  AOI21X1 g1779(.A0(n2825), .A1(n2811), .B0(n2827), .Y(n2828));
  OAI21X1 g1780(.A0(n2819), .A1(n2792), .B0(n2828), .Y(n2829));
  INVX1   g1781(.A(n2792), .Y(n2830));
  NOR2X1  g1782(.A(n2784), .B(n2764), .Y(n2831));
  NOR2X1  g1783(.A(n2824), .B(n2811), .Y(n2832));
  NOR2X1  g1784(.A(n2825), .B(n2812), .Y(n2833));
  NOR3X1  g1785(.A(n2833), .B(n2832), .C(n2819), .Y(n2834));
  OAI21X1 g1786(.A0(n2831), .A1(n2830), .B0(n2834), .Y(n2835));
  NAND2X1 g1787(.A(n2835), .B(n2829), .Y(n2836));
  AOI21X1 g1788(.A0(n2217), .A1(n2216), .B0(n2836), .Y(n2837));
  XOR2X1  g1789(.A(n2824), .B(n2811), .Y(n2838));
  INVX1   g1790(.A(n2783), .Y(n2839));
  NOR3X1  g1791(.A(n2774), .B(n2718), .C(n2682), .Y(n2840));
  OAI21X1 g1792(.A0(n2840), .A1(n2785), .B0(n2839), .Y(n2841));
  INVX1   g1793(.A(n2841), .Y(n2842));
  NOR3X1  g1794(.A(n2783), .B(n2774), .C(n2739), .Y(n2843));
  INVX1   g1795(.A(n2843), .Y(n2844));
  AOI21X1 g1796(.A0(n2697), .A1(n2696), .B0(n2844), .Y(n2845));
  NOR2X1  g1797(.A(n2845), .B(n2842), .Y(n2846));
  XOR2X1  g1798(.A(n2846), .B(n2838), .Y(n2847));
  OAI22X1 g1799(.A0(n2836), .A1(n2239), .B0(n2196), .B1(n2847), .Y(n2848));
  OAI22X1 g1800(.A0(n2765), .A1(n2322), .B0(n2184), .B1(n2847), .Y(n2849));
  INVX1   g1801(.A(n2847), .Y(n2850));
  OAI21X1 g1802(.A0(n2044), .A1(n2028), .B0(n2850), .Y(n2851));
  INVX1   g1803(.A(n2851), .Y(n2852));
  NOR4X1  g1804(.A(n2849), .B(n2848), .C(n2837), .D(n2852), .Y(n2853));
  INVX1   g1805(.A(n2853), .Y(n2854));
  NOR3X1  g1806(.A(n2784), .B(n2757), .C(n2716), .Y(n2855));
  XOR2X1  g1807(.A(n2824), .B(n2855), .Y(n2856));
  NAND3X1 g1808(.A(n2759), .B(P1_REG3_REG_16__SCAN_IN), .C(P1_REG3_REG_17__SCAN_IN), .Y(n2857));
  XOR2X1  g1809(.A(n2857), .B(P1_REG3_REG_18__SCAN_IN), .Y(n2858));
  INVX1   g1810(.A(n2858), .Y(n2859));
  NAND3X1 g1811(.A(n2859), .B(n2016), .C(n2014), .Y(n2860));
  NAND3X1 g1812(.A(n2016), .B(n2020), .C(P1_REG1_REG_18__SCAN_IN), .Y(n2861));
  AOI22X1 g1813(.A0(n2105), .A1(P1_REG0_REG_18__SCAN_IN), .B0(P1_REG2_REG_18__SCAN_IN), .B1(n2106), .Y(n2862));
  NAND3X1 g1814(.A(n2862), .B(n2861), .C(n2860), .Y(n2863));
  INVX1   g1815(.A(n2863), .Y(n2864));
  OAI22X1 g1816(.A0(n2824), .A1(n2068), .B0(n2104), .B1(n2864), .Y(n2865));
  AOI21X1 g1817(.A0(n2856), .A1(n2063), .B0(n2865), .Y(n2866));
  OAI21X1 g1818(.A0(n2836), .A1(n2053), .B0(n2866), .Y(n2867));
  NOR2X1  g1819(.A(n2867), .B(n2854), .Y(n2868));
  NAND2X1 g1820(.A(n2000), .B(P1_REG0_REG_17__SCAN_IN), .Y(n2869));
  OAI21X1 g1821(.A0(n2868), .A1(n2000), .B0(n2869), .Y(P1_U3505));
  INVX1   g1822(.A(n2819), .Y(n2871));
  AOI21X1 g1823(.A0(n2824), .A1(n2871), .B0(n2812), .Y(n2872));
  AOI21X1 g1824(.A0(n2825), .A1(n2819), .B0(n2872), .Y(n2873));
  INVX1   g1825(.A(n2873), .Y(n2874));
  AOI21X1 g1826(.A0(n2826), .A1(n2792), .B0(n2874), .Y(n2875));
  NOR2X1  g1827(.A(P1_IR_REG_31__SCAN_IN), .B(n1565), .Y(n2876));
  AOI21X1 g1828(.A0(n1571), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2876), .Y(n2877));
  INVX1   g1829(.A(n2877), .Y(n2878));
  NOR2X1  g1830(.A(n2005), .B(n1559), .Y(n2879));
  AOI21X1 g1831(.A0(n2878), .A1(n2005), .B0(n2879), .Y(n2880));
  XOR2X1  g1832(.A(n2880), .B(n2864), .Y(n2883));
  NOR2X1  g1833(.A(n2883), .B(n2875), .Y(n2884));
  AOI21X1 g1834(.A0(n2883), .A1(n2875), .B0(n2884), .Y(n2885));
  INVX1   g1835(.A(n2885), .Y(n2886));
  AOI22X1 g1836(.A0(n2811), .A1(n2093), .B0(n2047), .B1(n2886), .Y(n2887));
  OAI21X1 g1837(.A0(n2049), .A1(n2042), .B0(n2886), .Y(n2888));
  INVX1   g1838(.A(n2833), .Y(n2889));
  OAI22X1 g1839(.A0(n2842), .A1(n2845), .B0(n2824), .B1(n2811), .Y(n2890));
  NAND2X1 g1840(.A(n2890), .B(n2889), .Y(n2891));
  XOR2X1  g1841(.A(n2891), .B(n2883), .Y(n2892));
  INVX1   g1842(.A(n2892), .Y(n2893));
  OAI21X1 g1843(.A0(n2045), .A1(n2044), .B0(n2893), .Y(n2894));
  OAI21X1 g1844(.A0(n2038), .A1(n2028), .B0(n2893), .Y(n2895));
  NAND4X1 g1845(.A(n2894), .B(n2888), .C(n2887), .D(n2895), .Y(n2896));
  NAND2X1 g1846(.A(n2824), .B(n2855), .Y(n2897));
  INVX1   g1847(.A(n2880), .Y(n2898));
  XOR2X1  g1848(.A(n2898), .B(n2897), .Y(n2899));
  NAND4X1 g1849(.A(P1_REG3_REG_16__SCAN_IN), .B(P1_REG3_REG_17__SCAN_IN), .C(P1_REG3_REG_18__SCAN_IN), .D(n2759), .Y(n2900));
  XOR2X1  g1850(.A(n2900), .B(P1_REG3_REG_19__SCAN_IN), .Y(n2901));
  INVX1   g1851(.A(n2901), .Y(n2902));
  NAND3X1 g1852(.A(n2016), .B(n2020), .C(P1_REG1_REG_19__SCAN_IN), .Y(n2903));
  AOI22X1 g1853(.A0(n2105), .A1(P1_REG0_REG_19__SCAN_IN), .B0(P1_REG2_REG_19__SCAN_IN), .B1(n2106), .Y(n2904));
  NAND2X1 g1854(.A(n2904), .B(n2903), .Y(n2905));
  AOI21X1 g1855(.A0(n2902), .A1(n2360), .B0(n2905), .Y(n2906));
  OAI22X1 g1856(.A0(n2880), .A1(n2068), .B0(n2104), .B1(n2906), .Y(n2907));
  AOI21X1 g1857(.A0(n2899), .A1(n2063), .B0(n2907), .Y(n2908));
  OAI21X1 g1858(.A0(n2885), .A1(n2053), .B0(n2908), .Y(n2909));
  NOR2X1  g1859(.A(n2909), .B(n2896), .Y(n2910));
  NAND2X1 g1860(.A(n2000), .B(P1_REG0_REG_18__SCAN_IN), .Y(n2911));
  OAI21X1 g1861(.A0(n2910), .A1(n2000), .B0(n2911), .Y(P1_U3508));
  NAND2X1 g1862(.A(n2005), .B(n2041), .Y(n2913));
  OAI21X1 g1863(.A0(n2005), .A1(n1587), .B0(n2913), .Y(n2914));
  XOR2X1  g1864(.A(n2914), .B(n2906), .Y(n2915));
  AOI21X1 g1865(.A0(n2890), .A1(n2889), .B0(n2864), .Y(n2916));
  NAND3X1 g1866(.A(n2890), .B(n2864), .C(n2889), .Y(n2917));
  AOI21X1 g1867(.A0(n2917), .A1(n2880), .B0(n2916), .Y(n2918));
  XOR2X1  g1868(.A(n2918), .B(n2915), .Y(n2919));
  NOR2X1  g1869(.A(n2919), .B(n2184), .Y(n2920));
  NOR2X1  g1870(.A(n2898), .B(n2863), .Y(n2921));
  NOR2X1  g1871(.A(n2880), .B(n2864), .Y(n2922));
  INVX1   g1872(.A(n2922), .Y(n2923));
  OAI21X1 g1873(.A0(n2921), .A1(n2875), .B0(n2923), .Y(n2924));
  NOR2X1  g1874(.A(n2924), .B(n2915), .Y(n2925));
  INVX1   g1875(.A(n2906), .Y(n2926));
  XOR2X1  g1876(.A(n2914), .B(n2926), .Y(n2927));
  AOI21X1 g1877(.A0(n2915), .A1(n2924), .B0(n2925), .Y(n2929));
  OAI22X1 g1878(.A0(n2864), .A1(n2322), .B0(n2239), .B1(n2929), .Y(n2930));
  AOI21X1 g1879(.A0(n2217), .A1(n2216), .B0(n2929), .Y(n2931));
  NOR3X1  g1880(.A(n2931), .B(n2930), .C(n2920), .Y(n2932));
  NOR2X1  g1881(.A(n2919), .B(n2196), .Y(n2933));
  AOI21X1 g1882(.A0(n2183), .A1(n2029), .B0(n2919), .Y(n2934));
  NOR2X1  g1883(.A(n2934), .B(n2933), .Y(n2935));
  NAND2X1 g1884(.A(n2935), .B(n2932), .Y(n2936));
  NOR2X1  g1885(.A(n2898), .B(n2897), .Y(n2937));
  NOR2X1  g1886(.A(n2005), .B(n1587), .Y(n2938));
  AOI21X1 g1887(.A0(n2005), .A1(n2041), .B0(n2938), .Y(n2939));
  XOR2X1  g1888(.A(n2939), .B(n2937), .Y(n2940));
  INVX1   g1889(.A(P1_REG3_REG_20__SCAN_IN), .Y(n2941));
  INVX1   g1890(.A(P1_REG3_REG_19__SCAN_IN), .Y(n2942));
  NOR2X1  g1891(.A(n2900), .B(n2942), .Y(n2943));
  XOR2X1  g1892(.A(n2943), .B(n2941), .Y(n2944));
  AOI22X1 g1893(.A0(n2105), .A1(P1_REG0_REG_20__SCAN_IN), .B0(P1_REG2_REG_20__SCAN_IN), .B1(n2106), .Y(n2945));
  INVX1   g1894(.A(n2945), .Y(n2946));
  AOI21X1 g1895(.A0(n2359), .A1(P1_REG1_REG_20__SCAN_IN), .B0(n2946), .Y(n2947));
  OAI21X1 g1896(.A0(n2944), .A1(n2152), .B0(n2947), .Y(n2948));
  INVX1   g1897(.A(n2948), .Y(n2949));
  OAI22X1 g1898(.A0(n2939), .A1(n2068), .B0(n2104), .B1(n2949), .Y(n2950));
  AOI21X1 g1899(.A0(n2940), .A1(n2063), .B0(n2950), .Y(n2951));
  OAI21X1 g1900(.A0(n2929), .A1(n2053), .B0(n2951), .Y(n2952));
  NOR2X1  g1901(.A(n2952), .B(n2936), .Y(n2953));
  NAND2X1 g1902(.A(n2000), .B(P1_REG0_REG_19__SCAN_IN), .Y(n2954));
  OAI21X1 g1903(.A0(n2953), .A1(n2000), .B0(n2954), .Y(P1_U3510));
  NOR2X1  g1904(.A(n2005), .B(n1610), .Y(n2956));
  XOR2X1  g1905(.A(n2956), .B(n2949), .Y(n2957));
  NOR2X1  g1906(.A(n2914), .B(n2906), .Y(n2958));
  NAND2X1 g1907(.A(n2914), .B(n2906), .Y(n2959));
  INVX1   g1908(.A(n2959), .Y(n2960));
  NOR2X1  g1909(.A(n2918), .B(n2960), .Y(n2961));
  NOR2X1  g1910(.A(n2961), .B(n2958), .Y(n2962));
  XOR2X1  g1911(.A(n2962), .B(n2957), .Y(n2963));
  NOR2X1  g1912(.A(n2963), .B(n2184), .Y(n2964));
  INVX1   g1913(.A(n2964), .Y(n2965));
  NOR2X1  g1914(.A(n2939), .B(n2906), .Y(n2966));
  NOR2X1  g1915(.A(n2966), .B(n2924), .Y(n2967));
  INVX1   g1916(.A(n2956), .Y(n2968));
  OAI22X1 g1917(.A0(n2948), .A1(n2956), .B0(n2914), .B1(n2926), .Y(n2969));
  INVX1   g1918(.A(n2969), .Y(n2970));
  OAI21X1 g1919(.A0(n2968), .A1(n2949), .B0(n2970), .Y(n2971));
  INVX1   g1920(.A(n2924), .Y(n2972));
  AOI21X1 g1921(.A0(n2939), .A1(n2906), .B0(n2972), .Y(n2973));
  OAI21X1 g1922(.A0(n2939), .A1(n2906), .B0(n2957), .Y(n2974));
  OAI22X1 g1923(.A0(n2973), .A1(n2974), .B0(n2971), .B1(n2967), .Y(n2975));
  INVX1   g1924(.A(n2975), .Y(n2976));
  AOI22X1 g1925(.A0(n2926), .A1(n2093), .B0(n2047), .B1(n2976), .Y(n2977));
  OAI21X1 g1926(.A0(n2049), .A1(n2042), .B0(n2976), .Y(n2978));
  NOR2X1  g1927(.A(n2963), .B(n2196), .Y(n2979));
  AOI21X1 g1928(.A0(n2183), .A1(n2029), .B0(n2963), .Y(n2980));
  NOR2X1  g1929(.A(n2980), .B(n2979), .Y(n2981));
  NAND4X1 g1930(.A(n2978), .B(n2977), .C(n2965), .D(n2981), .Y(n2982));
  NOR2X1  g1931(.A(n2975), .B(n2053), .Y(n2983));
  NAND4X1 g1932(.A(n2880), .B(n2824), .C(n2855), .D(n2939), .Y(n2984));
  XOR2X1  g1933(.A(n2968), .B(n2984), .Y(n2985));
  INVX1   g1934(.A(P1_REG3_REG_21__SCAN_IN), .Y(n2986));
  NOR3X1  g1935(.A(n2900), .B(n2942), .C(n2941), .Y(n2987));
  XOR2X1  g1936(.A(n2987), .B(n2986), .Y(n2988));
  INVX1   g1937(.A(n2988), .Y(n2989));
  NAND3X1 g1938(.A(n2016), .B(n2020), .C(P1_REG1_REG_21__SCAN_IN), .Y(n2990));
  AOI22X1 g1939(.A0(n2105), .A1(P1_REG0_REG_21__SCAN_IN), .B0(P1_REG2_REG_21__SCAN_IN), .B1(n2106), .Y(n2991));
  NAND2X1 g1940(.A(n2991), .B(n2990), .Y(n2992));
  AOI21X1 g1941(.A0(n2989), .A1(n2360), .B0(n2992), .Y(n2993));
  INVX1   g1942(.A(n2993), .Y(n2994));
  AOI22X1 g1943(.A0(n2956), .A1(n2309), .B0(n2054), .B1(n2994), .Y(n2995));
  OAI21X1 g1944(.A0(n2985), .A1(n2064), .B0(n2995), .Y(n2996));
  NOR3X1  g1945(.A(n2996), .B(n2983), .C(n2982), .Y(n2997));
  NAND2X1 g1946(.A(n2000), .B(P1_REG0_REG_20__SCAN_IN), .Y(n2998));
  OAI21X1 g1947(.A0(n2997), .A1(n2000), .B0(n2998), .Y(P1_U3511));
  NOR2X1  g1948(.A(n2005), .B(n1635), .Y(n3000));
  XOR2X1  g1949(.A(n3000), .B(n2993), .Y(n3001));
  NOR3X1  g1950(.A(n2948), .B(n2005), .C(n1610), .Y(n3002));
  INVX1   g1951(.A(n3002), .Y(n3003));
  NOR2X1  g1952(.A(n2956), .B(n2949), .Y(n3004));
  INVX1   g1953(.A(n2958), .Y(n3005));
  OAI21X1 g1954(.A0(n2918), .A1(n2960), .B0(n3005), .Y(n3006));
  AOI21X1 g1955(.A0(n3006), .A1(n3003), .B0(n3004), .Y(n3007));
  XOR2X1  g1956(.A(n3007), .B(n3001), .Y(n3008));
  NOR2X1  g1957(.A(n3008), .B(n2184), .Y(n3009));
  AOI21X1 g1958(.A0(n2914), .A1(n2926), .B0(n2956), .Y(n3010));
  AOI21X1 g1959(.A0(n2956), .A1(n2966), .B0(n2948), .Y(n3011));
  NOR2X1  g1960(.A(n3011), .B(n3010), .Y(n3012));
  AOI21X1 g1961(.A0(n2970), .A1(n2924), .B0(n3012), .Y(n3013));
  NOR3X1  g1962(.A(n2994), .B(n2005), .C(n1635), .Y(n3014));
  OAI21X1 g1963(.A0(n2005), .A1(n1635), .B0(n2994), .Y(n3015));
  INVX1   g1964(.A(n3015), .Y(n3016));
  NOR3X1  g1965(.A(n3012), .B(n3016), .C(n3014), .Y(n3017));
  OAI21X1 g1966(.A0(n2969), .A1(n2972), .B0(n3017), .Y(n3018));
  OAI21X1 g1967(.A0(n3013), .A1(n3001), .B0(n3018), .Y(n3019));
  OAI22X1 g1968(.A0(n2949), .A1(n2322), .B0(n2239), .B1(n3019), .Y(n3020));
  AOI21X1 g1969(.A0(n2217), .A1(n2216), .B0(n3019), .Y(n3021));
  NOR3X1  g1970(.A(n3021), .B(n3020), .C(n3009), .Y(n3022));
  INVX1   g1971(.A(n3008), .Y(n3023));
  AOI21X1 g1972(.A0(n2183), .A1(n2029), .B0(n3008), .Y(n3024));
  AOI21X1 g1973(.A0(n3023), .A1(n2038), .B0(n3024), .Y(n3025));
  NAND2X1 g1974(.A(n3025), .B(n3022), .Y(n3026));
  NOR2X1  g1975(.A(n2956), .B(n2984), .Y(n3027));
  INVX1   g1976(.A(n3000), .Y(n3028));
  XOR2X1  g1977(.A(n3028), .B(n3027), .Y(n3029));
  NOR4X1  g1978(.A(n2942), .B(n2986), .C(n2941), .D(n2900), .Y(n3030));
  XOR2X1  g1979(.A(n3030), .B(P1_REG3_REG_22__SCAN_IN), .Y(n3031));
  NAND3X1 g1980(.A(n2016), .B(n2020), .C(P1_REG1_REG_22__SCAN_IN), .Y(n3032));
  AOI22X1 g1981(.A0(n2105), .A1(P1_REG0_REG_22__SCAN_IN), .B0(P1_REG2_REG_22__SCAN_IN), .B1(n2106), .Y(n3033));
  NAND2X1 g1982(.A(n3033), .B(n3032), .Y(n3034));
  AOI21X1 g1983(.A0(n3031), .A1(n2360), .B0(n3034), .Y(n3035));
  OAI22X1 g1984(.A0(n3028), .A1(n2068), .B0(n2104), .B1(n3035), .Y(n3036));
  AOI21X1 g1985(.A0(n3029), .A1(n2063), .B0(n3036), .Y(n3037));
  OAI21X1 g1986(.A0(n3019), .A1(n2053), .B0(n3037), .Y(n3038));
  NOR2X1  g1987(.A(n3038), .B(n3026), .Y(n3039));
  NAND2X1 g1988(.A(n2000), .B(P1_REG0_REG_21__SCAN_IN), .Y(n3040));
  OAI21X1 g1989(.A0(n3039), .A1(n2000), .B0(n3040), .Y(P1_U3512));
  NOR2X1  g1990(.A(n2005), .B(n1653), .Y(n3042));
  XOR2X1  g1991(.A(n3042), .B(n3035), .Y(n3043));
  INVX1   g1992(.A(n3014), .Y(n3044));
  INVX1   g1993(.A(n3004), .Y(n3045));
  OAI21X1 g1994(.A0(n2962), .A1(n3002), .B0(n3045), .Y(n3046));
  AOI21X1 g1995(.A0(n3046), .A1(n3044), .B0(n3016), .Y(n3047));
  XOR2X1  g1996(.A(n3047), .B(n3043), .Y(n3048));
  OAI21X1 g1997(.A0(n2005), .A1(n1635), .B0(n2993), .Y(n3049));
  NOR2X1  g1998(.A(n2969), .B(n2921), .Y(n3050));
  NAND2X1 g1999(.A(n3050), .B(n3049), .Y(n3051));
  OAI22X1 g2000(.A0(n3010), .A1(n3011), .B0(n2969), .B1(n2923), .Y(n3052));
  NOR3X1  g2001(.A(n2993), .B(n2005), .C(n1635), .Y(n3053));
  AOI21X1 g2002(.A0(n3052), .A1(n3049), .B0(n3053), .Y(n3054));
  OAI21X1 g2003(.A0(n3051), .A1(n2875), .B0(n3054), .Y(n3055));
  XOR2X1  g2004(.A(n3055), .B(n3043), .Y(n3056));
  OAI22X1 g2005(.A0(n2993), .A1(n2322), .B0(n2239), .B1(n3056), .Y(n3057));
  AOI21X1 g2006(.A0(n2217), .A1(n2216), .B0(n3056), .Y(n3058));
  NOR2X1  g2007(.A(n3058), .B(n3057), .Y(n3059));
  OAI21X1 g2008(.A0(n3048), .A1(n2184), .B0(n3059), .Y(n3060));
  NOR2X1  g2009(.A(n3048), .B(n2196), .Y(n3061));
  AOI21X1 g2010(.A0(n2183), .A1(n2029), .B0(n3048), .Y(n3062));
  NOR3X1  g2011(.A(n3000), .B(n2956), .C(n2984), .Y(n3063));
  INVX1   g2012(.A(n3042), .Y(n3064));
  XOR2X1  g2013(.A(n3064), .B(n3063), .Y(n3065));
  NAND2X1 g2014(.A(n3030), .B(P1_REG3_REG_22__SCAN_IN), .Y(n3066));
  XOR2X1  g2015(.A(n3066), .B(P1_REG3_REG_23__SCAN_IN), .Y(n3067));
  AOI22X1 g2016(.A0(n2105), .A1(P1_REG0_REG_23__SCAN_IN), .B0(P1_REG2_REG_23__SCAN_IN), .B1(n2106), .Y(n3068));
  INVX1   g2017(.A(n3068), .Y(n3069));
  AOI21X1 g2018(.A0(n2359), .A1(P1_REG1_REG_23__SCAN_IN), .B0(n3069), .Y(n3070));
  OAI21X1 g2019(.A0(n3067), .A1(n2152), .B0(n3070), .Y(n3071));
  INVX1   g2020(.A(n3071), .Y(n3072));
  OAI22X1 g2021(.A0(n3064), .A1(n2068), .B0(n2104), .B1(n3072), .Y(n3073));
  AOI21X1 g2022(.A0(n3065), .A1(n2063), .B0(n3073), .Y(n3074));
  OAI21X1 g2023(.A0(n3056), .A1(n2053), .B0(n3074), .Y(n3075));
  NOR4X1  g2024(.A(n3062), .B(n3061), .C(n3060), .D(n3075), .Y(n3076));
  NAND2X1 g2025(.A(n2000), .B(P1_REG0_REG_22__SCAN_IN), .Y(n3077));
  OAI21X1 g2026(.A0(n3076), .A1(n2000), .B0(n3077), .Y(P1_U3513));
  OAI21X1 g2027(.A0(n3042), .A1(n3035), .B0(n3047), .Y(n3079));
  INVX1   g2028(.A(n3035), .Y(n3080));
  NOR3X1  g2029(.A(n3080), .B(n2005), .C(n1653), .Y(n3081));
  NAND2X1 g2030(.A(n1696), .B(n1694), .Y(n3082));
  XOR2X1  g2031(.A(n1675), .B(n3082), .Y(n3083));
  NOR2X1  g2032(.A(n3083), .B(n1156), .Y(n3084));
  OAI21X1 g2033(.A0(n3084), .A1(n1665), .B0(n2101), .Y(n3085));
  XOR2X1  g2034(.A(n3085), .B(n3071), .Y(n3086));
  NOR2X1  g2035(.A(n3086), .B(n3081), .Y(n3087));
  NAND2X1 g2036(.A(n3087), .B(n3079), .Y(n3088));
  NOR3X1  g2037(.A(n3071), .B(n2005), .C(n1677), .Y(n3089));
  NOR2X1  g2038(.A(n3042), .B(n3035), .Y(n3090));
  AOI21X1 g2039(.A0(n3085), .A1(n3071), .B0(n3090), .Y(n3091));
  INVX1   g2040(.A(n3091), .Y(n3092));
  NOR2X1  g2041(.A(n3092), .B(n3089), .Y(n3093));
  OAI21X1 g2042(.A0(n3047), .A1(n3081), .B0(n3093), .Y(n3094));
  AOI21X1 g2043(.A0(n3094), .A1(n3088), .B0(n2184), .Y(n3095));
  INVX1   g2044(.A(n3086), .Y(n3096));
  NOR3X1  g2045(.A(n3035), .B(n2005), .C(n1653), .Y(n3097));
  OAI21X1 g2046(.A0(n2005), .A1(n1653), .B0(n3035), .Y(n3098));
  AOI21X1 g2047(.A0(n3098), .A1(n3055), .B0(n3097), .Y(n3099));
  XOR2X1  g2048(.A(n3099), .B(n3096), .Y(n3100));
  OAI22X1 g2049(.A0(n3035), .A1(n2322), .B0(n2239), .B1(n3100), .Y(n3101));
  AOI21X1 g2050(.A0(n2217), .A1(n2216), .B0(n3100), .Y(n3102));
  NOR3X1  g2051(.A(n3102), .B(n3101), .C(n3095), .Y(n3103));
  AOI21X1 g2052(.A0(n3094), .A1(n3088), .B0(n2196), .Y(n3104));
  AOI22X1 g2053(.A0(n3088), .A1(n3094), .B0(n2183), .B1(n2029), .Y(n3105));
  NOR2X1  g2054(.A(n3105), .B(n3104), .Y(n3106));
  NAND2X1 g2055(.A(n3106), .B(n3103), .Y(n3107));
  NOR2X1  g2056(.A(n3100), .B(n2053), .Y(n3108));
  OAI21X1 g2057(.A0(n2005), .A1(n1653), .B0(n3063), .Y(n3109));
  XOR2X1  g2058(.A(n3085), .B(n3109), .Y(n3110));
  INVX1   g2059(.A(n3085), .Y(n3111));
  NAND3X1 g2060(.A(n3030), .B(P1_REG3_REG_23__SCAN_IN), .C(P1_REG3_REG_22__SCAN_IN), .Y(n3112));
  XOR2X1  g2061(.A(n3112), .B(P1_REG3_REG_24__SCAN_IN), .Y(n3113));
  AOI22X1 g2062(.A0(n2105), .A1(P1_REG0_REG_24__SCAN_IN), .B0(P1_REG2_REG_24__SCAN_IN), .B1(n2106), .Y(n3114));
  INVX1   g2063(.A(n3114), .Y(n3115));
  AOI21X1 g2064(.A0(n2359), .A1(P1_REG1_REG_24__SCAN_IN), .B0(n3115), .Y(n3116));
  OAI21X1 g2065(.A0(n3113), .A1(n2152), .B0(n3116), .Y(n3117));
  AOI22X1 g2066(.A0(n3111), .A1(n2309), .B0(n2054), .B1(n3117), .Y(n3118));
  OAI21X1 g2067(.A0(n3110), .A1(n2064), .B0(n3118), .Y(n3119));
  NOR3X1  g2068(.A(n3119), .B(n3108), .C(n3107), .Y(n3120));
  NAND2X1 g2069(.A(n2000), .B(P1_REG0_REG_23__SCAN_IN), .Y(n3121));
  OAI21X1 g2070(.A0(n3120), .A1(n2000), .B0(n3121), .Y(P1_U3514));
  INVX1   g2071(.A(n3117), .Y(n3123));
  NOR2X1  g2072(.A(n2005), .B(n1703), .Y(n3124));
  XOR2X1  g2073(.A(n3124), .B(n3123), .Y(n3125));
  INVX1   g2074(.A(n3089), .Y(n3126));
  OAI21X1 g2075(.A0(n3081), .A1(n3015), .B0(n3091), .Y(n3127));
  NAND2X1 g2076(.A(n3127), .B(n3126), .Y(n3128));
  NOR3X1  g2077(.A(n3089), .B(n3081), .C(n3014), .Y(n3129));
  INVX1   g2078(.A(n3129), .Y(n3130));
  OAI21X1 g2079(.A0(n3130), .A1(n3007), .B0(n3128), .Y(n3131));
  XOR2X1  g2080(.A(n3131), .B(n3125), .Y(n3132));
  NAND2X1 g2081(.A(n3132), .B(n2045), .Y(n3133));
  INVX1   g2082(.A(n3133), .Y(n3134));
  NOR3X1  g2083(.A(n3072), .B(n2005), .C(n1677), .Y(n3135));
  AOI21X1 g2084(.A0(n3085), .A1(n3072), .B0(n3099), .Y(n3136));
  NOR2X1  g2085(.A(n3136), .B(n3135), .Y(n3137));
  NOR3X1  g2086(.A(n3117), .B(n2005), .C(n1703), .Y(n3138));
  NOR2X1  g2087(.A(n3124), .B(n3123), .Y(n3139));
  OAI21X1 g2088(.A0(n3139), .A1(n3138), .B0(n3137), .Y(n3140));
  XOR2X1  g2089(.A(n3124), .B(n3117), .Y(n3141));
  OAI21X1 g2090(.A0(n3141), .A1(n3137), .B0(n3140), .Y(n3142));
  AOI22X1 g2091(.A0(n3071), .A1(n2093), .B0(n2047), .B1(n3142), .Y(n3143));
  OAI21X1 g2092(.A0(n2049), .A1(n2042), .B0(n3142), .Y(n3144));
  NAND2X1 g2093(.A(n3144), .B(n3143), .Y(n3145));
  NAND2X1 g2094(.A(n3132), .B(n2038), .Y(n3146));
  OAI21X1 g2095(.A0(n2044), .A1(n2028), .B0(n3132), .Y(n3147));
  NAND2X1 g2096(.A(n3147), .B(n3146), .Y(n3148));
  NAND2X1 g2097(.A(n3142), .B(n2052), .Y(n3149));
  NOR2X1  g2098(.A(n3111), .B(n3109), .Y(n3150));
  INVX1   g2099(.A(n3124), .Y(n3151));
  XOR2X1  g2100(.A(n3151), .B(n3150), .Y(n3152));
  NAND4X1 g2101(.A(P1_REG3_REG_23__SCAN_IN), .B(P1_REG3_REG_24__SCAN_IN), .C(P1_REG3_REG_22__SCAN_IN), .D(n3030), .Y(n3153));
  XOR2X1  g2102(.A(n3153), .B(P1_REG3_REG_25__SCAN_IN), .Y(n3154));
  AOI22X1 g2103(.A0(n2105), .A1(P1_REG0_REG_25__SCAN_IN), .B0(P1_REG2_REG_25__SCAN_IN), .B1(n2106), .Y(n3155));
  INVX1   g2104(.A(n3155), .Y(n3156));
  AOI21X1 g2105(.A0(n2359), .A1(P1_REG1_REG_25__SCAN_IN), .B0(n3156), .Y(n3157));
  OAI21X1 g2106(.A0(n3154), .A1(n2152), .B0(n3157), .Y(n3158));
  INVX1   g2107(.A(n3158), .Y(n3159));
  OAI22X1 g2108(.A0(n3151), .A1(n2068), .B0(n2104), .B1(n3159), .Y(n3160));
  AOI21X1 g2109(.A0(n3152), .A1(n2063), .B0(n3160), .Y(n3161));
  NAND2X1 g2110(.A(n3161), .B(n3149), .Y(n3162));
  NOR4X1  g2111(.A(n3148), .B(n3145), .C(n3134), .D(n3162), .Y(n3163));
  NAND2X1 g2112(.A(n2000), .B(P1_REG0_REG_24__SCAN_IN), .Y(n3164));
  OAI21X1 g2113(.A0(n3163), .A1(n2000), .B0(n3164), .Y(P1_U3515));
  NOR2X1  g2114(.A(n2005), .B(n1728), .Y(n3166));
  XOR2X1  g2115(.A(n3166), .B(n3159), .Y(n3167));
  INVX1   g2116(.A(n3138), .Y(n3168));
  AOI21X1 g2117(.A0(n3131), .A1(n3168), .B0(n3139), .Y(n3169));
  XOR2X1  g2118(.A(n3169), .B(n3167), .Y(n3170));
  NOR3X1  g2119(.A(n3123), .B(n2005), .C(n1703), .Y(n3171));
  INVX1   g2120(.A(n3171), .Y(n3172));
  OAI22X1 g2121(.A0(n3135), .A1(n3136), .B0(n3124), .B1(n3117), .Y(n3173));
  NAND2X1 g2122(.A(n3173), .B(n3172), .Y(n3174));
  NOR2X1  g2123(.A(n3174), .B(n3167), .Y(n3175));
  NAND2X1 g2124(.A(n1739), .B(n1737), .Y(n3176));
  XOR2X1  g2125(.A(n1726), .B(n3176), .Y(n3177));
  NOR2X1  g2126(.A(n3177), .B(n1156), .Y(n3178));
  OAI21X1 g2127(.A0(n3178), .A1(n1716), .B0(n2101), .Y(n3179));
  XOR2X1  g2128(.A(n3179), .B(n3159), .Y(n3180));
  AOI21X1 g2129(.A0(n3173), .A1(n3172), .B0(n3180), .Y(n3181));
  NOR2X1  g2130(.A(n3181), .B(n3175), .Y(n3182));
  OAI22X1 g2131(.A0(n3123), .A1(n2322), .B0(n2239), .B1(n3182), .Y(n3183));
  AOI21X1 g2132(.A0(n2217), .A1(n2216), .B0(n3182), .Y(n3184));
  NOR2X1  g2133(.A(n3184), .B(n3183), .Y(n3185));
  OAI21X1 g2134(.A0(n3170), .A1(n2184), .B0(n3185), .Y(n3186));
  NOR2X1  g2135(.A(n3170), .B(n2196), .Y(n3187));
  AOI21X1 g2136(.A0(n2183), .A1(n2029), .B0(n3170), .Y(n3188));
  NAND2X1 g2137(.A(n3151), .B(n3150), .Y(n3189));
  XOR2X1  g2138(.A(n3166), .B(n3189), .Y(n3190));
  INVX1   g2139(.A(P1_REG3_REG_26__SCAN_IN), .Y(n3191));
  INVX1   g2140(.A(P1_REG3_REG_25__SCAN_IN), .Y(n3192));
  NOR2X1  g2141(.A(n3153), .B(n3192), .Y(n3193));
  XOR2X1  g2142(.A(n3193), .B(n3191), .Y(n3194));
  AOI22X1 g2143(.A0(n2105), .A1(P1_REG0_REG_26__SCAN_IN), .B0(P1_REG2_REG_26__SCAN_IN), .B1(n2106), .Y(n3195));
  INVX1   g2144(.A(n3195), .Y(n3196));
  AOI21X1 g2145(.A0(n2359), .A1(P1_REG1_REG_26__SCAN_IN), .B0(n3196), .Y(n3197));
  OAI21X1 g2146(.A0(n3194), .A1(n2152), .B0(n3197), .Y(n3198));
  INVX1   g2147(.A(n3198), .Y(n3199));
  OAI22X1 g2148(.A0(n3179), .A1(n2068), .B0(n2104), .B1(n3199), .Y(n3200));
  AOI21X1 g2149(.A0(n3190), .A1(n2063), .B0(n3200), .Y(n3201));
  OAI21X1 g2150(.A0(n3182), .A1(n2053), .B0(n3201), .Y(n3202));
  NOR4X1  g2151(.A(n3188), .B(n3187), .C(n3186), .D(n3202), .Y(n3203));
  NAND2X1 g2152(.A(n2000), .B(P1_REG0_REG_25__SCAN_IN), .Y(n3204));
  OAI21X1 g2153(.A0(n3203), .A1(n2000), .B0(n3204), .Y(P1_U3516));
  NOR2X1  g2154(.A(n2005), .B(n1746), .Y(n3206));
  XOR2X1  g2155(.A(n3206), .B(n3199), .Y(n3207));
  INVX1   g2156(.A(n3207), .Y(n3208));
  NOR3X1  g2157(.A(n3158), .B(n2005), .C(n1728), .Y(n3209));
  NOR2X1  g2158(.A(n3166), .B(n3159), .Y(n3210));
  INVX1   g2159(.A(n3210), .Y(n3211));
  OAI21X1 g2160(.A0(n3169), .A1(n3209), .B0(n3211), .Y(n3212));
  XOR2X1  g2161(.A(n3212), .B(n3208), .Y(n3213));
  NOR2X1  g2162(.A(n3213), .B(n2184), .Y(n3214));
  NOR3X1  g2163(.A(n3159), .B(n2005), .C(n1728), .Y(n3215));
  INVX1   g2164(.A(n3215), .Y(n3216));
  NAND3X1 g2165(.A(n3216), .B(n3173), .C(n3172), .Y(n3217));
  OAI21X1 g2166(.A0(n2005), .A1(n1728), .B0(n3159), .Y(n3218));
  OAI21X1 g2167(.A0(n3206), .A1(n3198), .B0(n3218), .Y(n3219));
  NOR3X1  g2168(.A(n3199), .B(n2005), .C(n1746), .Y(n3220));
  NOR2X1  g2169(.A(n3220), .B(n3219), .Y(n3221));
  NAND2X1 g2170(.A(n3218), .B(n3174), .Y(n3222));
  NOR2X1  g2171(.A(n3208), .B(n3215), .Y(n3223));
  AOI22X1 g2172(.A0(n3222), .A1(n3223), .B0(n3221), .B1(n3217), .Y(n3224));
  AOI22X1 g2173(.A0(n3158), .A1(n2093), .B0(n2047), .B1(n3224), .Y(n3225));
  OAI21X1 g2174(.A0(n2049), .A1(n2042), .B0(n3224), .Y(n3226));
  NAND2X1 g2175(.A(n3226), .B(n3225), .Y(n3227));
  NOR2X1  g2176(.A(n3227), .B(n3214), .Y(n3228));
  NOR2X1  g2177(.A(n3213), .B(n2196), .Y(n3229));
  AOI21X1 g2178(.A0(n2183), .A1(n2029), .B0(n3213), .Y(n3230));
  NOR2X1  g2179(.A(n3230), .B(n3229), .Y(n3231));
  NAND2X1 g2180(.A(n3231), .B(n3228), .Y(n3232));
  INVX1   g2181(.A(n3224), .Y(n3233));
  NOR2X1  g2182(.A(n3233), .B(n2053), .Y(n3234));
  NOR4X1  g2183(.A(n3124), .B(n3111), .C(n3109), .D(n3166), .Y(n3235));
  XOR2X1  g2184(.A(n3206), .B(n3235), .Y(n3236));
  INVX1   g2185(.A(P1_REG3_REG_27__SCAN_IN), .Y(n3237));
  NOR3X1  g2186(.A(n3153), .B(n3192), .C(n3191), .Y(n3238));
  XOR2X1  g2187(.A(n3238), .B(n3237), .Y(n3239));
  AOI22X1 g2188(.A0(n2105), .A1(P1_REG0_REG_27__SCAN_IN), .B0(P1_REG2_REG_27__SCAN_IN), .B1(n2106), .Y(n3240));
  INVX1   g2189(.A(n3240), .Y(n3241));
  AOI21X1 g2190(.A0(n2359), .A1(P1_REG1_REG_27__SCAN_IN), .B0(n3241), .Y(n3242));
  OAI21X1 g2191(.A0(n3239), .A1(n2152), .B0(n3242), .Y(n3243));
  AOI22X1 g2192(.A0(n3206), .A1(n2309), .B0(n2054), .B1(n3243), .Y(n3244));
  OAI21X1 g2193(.A0(n3236), .A1(n2064), .B0(n3244), .Y(n3245));
  NOR3X1  g2194(.A(n3245), .B(n3234), .C(n3232), .Y(n3246));
  NAND2X1 g2195(.A(n2000), .B(P1_REG0_REG_26__SCAN_IN), .Y(n3247));
  OAI21X1 g2196(.A0(n3246), .A1(n2000), .B0(n3247), .Y(P1_U3517));
  OAI21X1 g2197(.A0(n2005), .A1(n1746), .B0(n3198), .Y(n3249));
  INVX1   g2198(.A(n3249), .Y(n3250));
  NAND2X1 g2199(.A(n3206), .B(n3199), .Y(n3252));
  INVX1   g2200(.A(n3243), .Y(n3253));
  INVX1   g2201(.A(n1760), .Y(n3254));
  AOI21X1 g2202(.A0(n1776), .A1(n3254), .B0(n2005), .Y(n3255));
  XOR2X1  g2203(.A(n3255), .B(n3253), .Y(n3256));
  INVX1   g2204(.A(n3256), .Y(n3257));
  NAND2X1 g2205(.A(n3257), .B(n3252), .Y(n3258));
  NOR2X1  g2206(.A(n3258), .B(n4824), .Y(n3259));
  NAND2X1 g2207(.A(n3256), .B(n3249), .Y(n3260));
  AOI21X1 g2208(.A0(n3212), .A1(n3252), .B0(n3260), .Y(n3261));
  OAI21X1 g2209(.A0(n3261), .A1(n3259), .B0(n2045), .Y(n3262));
  NAND2X1 g2210(.A(n1765), .B(n1763), .Y(n3263));
  XOR2X1  g2211(.A(n1744), .B(n3263), .Y(n3264));
  NOR2X1  g2212(.A(n3264), .B(n1156), .Y(n3265));
  OAI21X1 g2213(.A0(n3265), .A1(n1734), .B0(n2101), .Y(n3266));
  AOI22X1 g2214(.A0(n3199), .A1(n3266), .B0(n3179), .B1(n3159), .Y(n3267));
  OAI21X1 g2215(.A0(n3215), .A1(n3171), .B0(n3267), .Y(n3268));
  NOR2X1  g2216(.A(n3219), .B(n3173), .Y(n3269));
  NOR2X1  g2217(.A(n3269), .B(n3220), .Y(n3270));
  NAND2X1 g2218(.A(n3270), .B(n3268), .Y(n3271));
  XOR2X1  g2219(.A(n3271), .B(n3257), .Y(n3272));
  AOI22X1 g2220(.A0(n3198), .A1(n2093), .B0(n2047), .B1(n3272), .Y(n3273));
  OAI21X1 g2221(.A0(n2049), .A1(n2042), .B0(n3272), .Y(n3274));
  NAND3X1 g2222(.A(n3274), .B(n3273), .C(n3262), .Y(n3275));
  NOR2X1  g2223(.A(n3261), .B(n3259), .Y(n3276));
  NOR2X1  g2224(.A(n3276), .B(n2196), .Y(n3277));
  AOI21X1 g2225(.A0(n2183), .A1(n2029), .B0(n3276), .Y(n3278));
  NAND2X1 g2226(.A(n3272), .B(n2052), .Y(n3279));
  NOR3X1  g2227(.A(n3206), .B(n3166), .C(n3189), .Y(n3280));
  INVX1   g2228(.A(n3255), .Y(n3281));
  XOR2X1  g2229(.A(n3281), .B(n3280), .Y(n3282));
  INVX1   g2230(.A(P1_REG3_REG_28__SCAN_IN), .Y(n3283));
  NOR4X1  g2231(.A(n3237), .B(n3192), .C(n3191), .D(n3153), .Y(n3284));
  XOR2X1  g2232(.A(n3284), .B(n3283), .Y(n3285));
  AOI22X1 g2233(.A0(n2105), .A1(P1_REG0_REG_28__SCAN_IN), .B0(P1_REG2_REG_28__SCAN_IN), .B1(n2106), .Y(n3286));
  INVX1   g2234(.A(n3286), .Y(n3287));
  AOI21X1 g2235(.A0(n2359), .A1(P1_REG1_REG_28__SCAN_IN), .B0(n3287), .Y(n3288));
  OAI21X1 g2236(.A0(n3285), .A1(n2152), .B0(n3288), .Y(n3289));
  INVX1   g2237(.A(n3289), .Y(n3290));
  OAI22X1 g2238(.A0(n3281), .A1(n2068), .B0(n2104), .B1(n3290), .Y(n3291));
  AOI21X1 g2239(.A0(n3282), .A1(n2063), .B0(n3291), .Y(n3292));
  NAND2X1 g2240(.A(n3292), .B(n3279), .Y(n3293));
  NOR4X1  g2241(.A(n3278), .B(n3277), .C(n3275), .D(n3293), .Y(n3294));
  NAND2X1 g2242(.A(n2000), .B(P1_REG0_REG_27__SCAN_IN), .Y(n3295));
  OAI21X1 g2243(.A0(n3294), .A1(n2000), .B0(n3295), .Y(P1_U3518));
  NOR2X1  g2244(.A(n2005), .B(n1793), .Y(n3297));
  XOR2X1  g2245(.A(n3297), .B(n3290), .Y(n3298));
  AOI21X1 g2246(.A0(n3253), .A1(n3249), .B0(n3255), .Y(n3299));
  AOI21X1 g2247(.A0(n3243), .A1(n3250), .B0(n3299), .Y(n3300));
  NAND2X1 g2248(.A(n3255), .B(n3253), .Y(n3301));
  NAND3X1 g2249(.A(n3301), .B(n3212), .C(n3252), .Y(n3302));
  NAND2X1 g2250(.A(n3302), .B(n3300), .Y(n3303));
  XOR2X1  g2251(.A(n3303), .B(n3298), .Y(n3304));
  NAND2X1 g2252(.A(n3304), .B(n2045), .Y(n3305));
  AOI21X1 g2253(.A0(n3281), .A1(n3253), .B0(n3268), .Y(n3306));
  AOI21X1 g2254(.A0(n3255), .A1(n3243), .B0(n3306), .Y(n3307));
  OAI22X1 g2255(.A0(n3255), .A1(n3243), .B0(n3220), .B1(n3269), .Y(n3308));
  NAND2X1 g2256(.A(n3308), .B(n3307), .Y(n3309));
  XOR2X1  g2257(.A(n3309), .B(n3298), .Y(n3310));
  OAI22X1 g2258(.A0(n3253), .A1(n2322), .B0(n2239), .B1(n3310), .Y(n3311));
  AOI21X1 g2259(.A0(n2217), .A1(n2216), .B0(n3310), .Y(n3312));
  NOR2X1  g2260(.A(n3312), .B(n3311), .Y(n3313));
  NAND2X1 g2261(.A(n3313), .B(n3305), .Y(n3314));
  NAND2X1 g2262(.A(n3304), .B(n2038), .Y(n3315));
  OAI21X1 g2263(.A0(n2044), .A1(n2028), .B0(n3304), .Y(n3316));
  NAND2X1 g2264(.A(n3316), .B(n3315), .Y(n3317));
  NAND2X1 g2265(.A(n3281), .B(n3280), .Y(n3318));
  XOR2X1  g2266(.A(n3297), .B(n3318), .Y(n3319));
  INVX1   g2267(.A(n1784), .Y(n3320));
  NAND2X1 g2268(.A(n1815), .B(n1813), .Y(n3321));
  XOR2X1  g2269(.A(n1791), .B(n3321), .Y(n3322));
  OAI21X1 g2270(.A0(n3322), .A1(n1156), .B0(n3320), .Y(n3323));
  NAND2X1 g2271(.A(n2101), .B(n3323), .Y(n3324));
  NAND4X1 g2272(.A(n2360), .B(P1_REG3_REG_27__SCAN_IN), .C(P1_REG3_REG_28__SCAN_IN), .D(n3238), .Y(n3325));
  NAND2X1 g2273(.A(n2105), .B(P1_REG0_REG_29__SCAN_IN), .Y(n3326));
  AOI22X1 g2274(.A0(n2106), .A1(P1_REG2_REG_29__SCAN_IN), .B0(P1_REG1_REG_29__SCAN_IN), .B1(n2359), .Y(n3327));
  NAND3X1 g2275(.A(n3327), .B(n3326), .C(n3325), .Y(n3328));
  INVX1   g2276(.A(n3328), .Y(n3329));
  OAI22X1 g2277(.A0(n3324), .A1(n2068), .B0(n2104), .B1(n3329), .Y(n3330));
  AOI21X1 g2278(.A0(n3319), .A1(n2063), .B0(n3330), .Y(n3331));
  OAI21X1 g2279(.A0(n3310), .A1(n2053), .B0(n3331), .Y(n3332));
  NOR3X1  g2280(.A(n3332), .B(n3317), .C(n3314), .Y(n3333));
  NAND2X1 g2281(.A(n2000), .B(P1_REG0_REG_28__SCAN_IN), .Y(n3334));
  OAI21X1 g2282(.A0(n3333), .A1(n2000), .B0(n3334), .Y(P1_U3519));
  AOI21X1 g2283(.A0(n3308), .A1(n3307), .B0(n3324), .Y(n3336));
  NOR3X1  g2284(.A(n3290), .B(n2005), .C(n1793), .Y(n3337));
  AOI21X1 g2285(.A0(n3308), .A1(n3307), .B0(n3290), .Y(n3338));
  NOR3X1  g2286(.A(n3338), .B(n3337), .C(n3336), .Y(n3339));
  INVX1   g2287(.A(n1810), .Y(n3340));
  NOR3X1  g2288(.A(n1820), .B(n1816), .C(n1812), .Y(n3341));
  INVX1   g2289(.A(n1820), .Y(n3342));
  AOI21X1 g2290(.A0(n1844), .A1(n1842), .B0(n3342), .Y(n3343));
  OAI21X1 g2291(.A0(n3343), .A1(n3341), .B0(n1149), .Y(n3344));
  AOI21X1 g2292(.A0(n3344), .A1(n3340), .B0(n2005), .Y(n3345));
  XOR2X1  g2293(.A(n3345), .B(n3329), .Y(n3346));
  XOR2X1  g2294(.A(n3346), .B(n3339), .Y(n3347));
  NAND2X1 g2295(.A(n3347), .B(n2047), .Y(n3348));
  AOI21X1 g2296(.A0(n2092), .A1(n1885), .B0(n2005), .Y(n3349));
  NOR3X1  g2297(.A(n3349), .B(n1989), .C(n1984), .Y(n3350));
  NAND3X1 g2298(.A(n2016), .B(n2020), .C(P1_REG1_REG_30__SCAN_IN), .Y(n3351));
  AOI22X1 g2299(.A0(n2105), .A1(P1_REG0_REG_30__SCAN_IN), .B0(P1_REG2_REG_30__SCAN_IN), .B1(n2106), .Y(n3352));
  NAND2X1 g2300(.A(n3352), .B(n3351), .Y(n3353));
  AOI22X1 g2301(.A0(n3350), .A1(n3353), .B0(n3289), .B1(n2093), .Y(n3354));
  OAI21X1 g2302(.A0(n2049), .A1(n2042), .B0(n3347), .Y(n3355));
  NAND3X1 g2303(.A(n3355), .B(n3354), .C(n3348), .Y(n3356));
  OAI21X1 g2304(.A0(n3324), .A1(n3289), .B0(n4365), .Y(n3358));
  AOI21X1 g2305(.A0(n3302), .A1(n3300), .B0(n3358), .Y(n3359));
  OAI21X1 g2306(.A0(n2005), .A1(n1793), .B0(n3289), .Y(n3360));
  NAND4X1 g2307(.A(n3302), .B(n3300), .C(n3360), .D(n3346), .Y(n3361));
  NOR3X1  g2308(.A(n3289), .B(n2005), .C(n1793), .Y(n3362));
  NOR2X1  g2309(.A(n3346), .B(n3360), .Y(n3363));
  AOI21X1 g2310(.A0(n3346), .A1(n3362), .B0(n3363), .Y(n3364));
  NAND2X1 g2311(.A(n3364), .B(n3361), .Y(n3365));
  OAI22X1 g2312(.A0(n3359), .A1(n3365), .B0(n2045), .B1(n2044), .Y(n3366));
  OAI22X1 g2313(.A0(n3359), .A1(n3365), .B0(n2038), .B1(n2028), .Y(n3367));
  NAND2X1 g2314(.A(n3367), .B(n3366), .Y(n3368));
  XOR2X1  g2315(.A(n4365), .B(n3339), .Y(n3369));
  NOR2X1  g2316(.A(n3369), .B(n2053), .Y(n3370));
  NAND2X1 g2317(.A(n3344), .B(n3340), .Y(n3371));
  NAND2X1 g2318(.A(n2101), .B(n3371), .Y(n3372));
  NOR2X1  g2319(.A(n3297), .B(n3318), .Y(n3373));
  XOR2X1  g2320(.A(n3345), .B(n3373), .Y(n3374));
  OAI22X1 g2321(.A0(n3372), .A1(n2068), .B0(n2064), .B1(n3374), .Y(n3375));
  NOR4X1  g2322(.A(n3370), .B(n3368), .C(n3356), .D(n3375), .Y(n3376));
  NAND2X1 g2323(.A(n2000), .B(P1_REG0_REG_29__SCAN_IN), .Y(n3377));
  OAI21X1 g2324(.A0(n3376), .A1(n2000), .B0(n3377), .Y(P1_U3520));
  NAND2X1 g2325(.A(n3372), .B(n3373), .Y(n3379));
  NOR2X1  g2326(.A(n2005), .B(n1848), .Y(n3380));
  XOR2X1  g2327(.A(n3380), .B(n3379), .Y(n3381));
  OAI21X1 g2328(.A0(n1847), .A1(n1831), .B0(n2101), .Y(n3382));
  NAND3X1 g2329(.A(n2016), .B(n2020), .C(P1_REG1_REG_31__SCAN_IN), .Y(n3383));
  AOI22X1 g2330(.A0(n2105), .A1(P1_REG0_REG_31__SCAN_IN), .B0(P1_REG2_REG_31__SCAN_IN), .B1(n2106), .Y(n3384));
  NAND2X1 g2331(.A(n3384), .B(n3383), .Y(n3385));
  NAND2X1 g2332(.A(n3385), .B(n3350), .Y(n3386));
  OAI21X1 g2333(.A0(n3382), .A1(n2068), .B0(n3386), .Y(n3387));
  AOI21X1 g2334(.A0(n3381), .A1(n2063), .B0(n3387), .Y(n3388));
  NAND2X1 g2335(.A(n2000), .B(P1_REG0_REG_30__SCAN_IN), .Y(n3389));
  OAI21X1 g2336(.A0(n3388), .A1(n2000), .B0(n3389), .Y(P1_U3521));
  NAND3X1 g2337(.A(n3382), .B(n3372), .C(n3373), .Y(n3391));
  INVX1   g2338(.A(n1853), .Y(n3392));
  OAI21X1 g2339(.A0(n1845), .A1(n1833), .B0(n1858), .Y(n3393));
  NAND4X1 g2340(.A(n1857), .B(n1836), .C(n1834), .D(n1862), .Y(n3394));
  NAND4X1 g2341(.A(n3394), .B(n3393), .C(n1149), .D(n1866), .Y(n3395));
  AOI21X1 g2342(.A0(n3395), .A1(n3392), .B0(n2005), .Y(n3396));
  XOR2X1  g2343(.A(n3396), .B(n3391), .Y(n3397));
  OAI21X1 g2344(.A0(n1868), .A1(n1853), .B0(n2101), .Y(n3398));
  OAI21X1 g2345(.A0(n3398), .A1(n2068), .B0(n3386), .Y(n3399));
  AOI21X1 g2346(.A0(n3397), .A1(n2063), .B0(n3399), .Y(n3400));
  NAND2X1 g2347(.A(n2000), .B(P1_REG0_REG_31__SCAN_IN), .Y(n3401));
  OAI21X1 g2348(.A0(n3400), .A1(n2000), .B0(n3401), .Y(P1_U3522));
  INVX1   g2349(.A(n1999), .Y(n3403));
  NAND3X1 g2350(.A(n3403), .B(n1997), .C(n1893), .Y(n3404));
  NAND2X1 g2351(.A(n3404), .B(P1_REG1_REG_0__SCAN_IN), .Y(n3405));
  OAI21X1 g2352(.A0(n3404), .A1(n2072), .B0(n3405), .Y(P1_U3523));
  NAND2X1 g2353(.A(n3404), .B(P1_REG1_REG_1__SCAN_IN), .Y(n3407));
  OAI21X1 g2354(.A0(n3404), .A1(n2115), .B0(n3407), .Y(P1_U3524));
  NAND2X1 g2355(.A(n3404), .B(P1_REG1_REG_2__SCAN_IN), .Y(n3409));
  OAI21X1 g2356(.A0(n3404), .A1(n2158), .B0(n3409), .Y(P1_U3525));
  NAND2X1 g2357(.A(n3404), .B(P1_REG1_REG_3__SCAN_IN), .Y(n3411));
  OAI21X1 g2358(.A0(n3404), .A1(n2213), .B0(n3411), .Y(P1_U3526));
  NAND2X1 g2359(.A(n3404), .B(P1_REG1_REG_4__SCAN_IN), .Y(n3413));
  OAI21X1 g2360(.A0(n3404), .A1(n2267), .B0(n3413), .Y(P1_U3527));
  NAND2X1 g2361(.A(n3404), .B(P1_REG1_REG_5__SCAN_IN), .Y(n3415));
  OAI21X1 g2362(.A0(n3404), .A1(n2319), .B0(n3415), .Y(P1_U3528));
  NAND2X1 g2363(.A(n3404), .B(P1_REG1_REG_6__SCAN_IN), .Y(n3417));
  OAI21X1 g2364(.A0(n3404), .A1(n2370), .B0(n3417), .Y(P1_U3529));
  NAND2X1 g2365(.A(n3404), .B(P1_REG1_REG_7__SCAN_IN), .Y(n3419));
  OAI21X1 g2366(.A0(n3404), .A1(n2415), .B0(n3419), .Y(P1_U3530));
  NAND2X1 g2367(.A(n3404), .B(P1_REG1_REG_8__SCAN_IN), .Y(n3421));
  OAI21X1 g2368(.A0(n3404), .A1(n2458), .B0(n3421), .Y(P1_U3531));
  NAND2X1 g2369(.A(n3404), .B(P1_REG1_REG_9__SCAN_IN), .Y(n3423));
  OAI21X1 g2370(.A0(n3404), .A1(n2503), .B0(n3423), .Y(P1_U3532));
  NAND2X1 g2371(.A(n3404), .B(P1_REG1_REG_10__SCAN_IN), .Y(n3425));
  OAI21X1 g2372(.A0(n3404), .A1(n2550), .B0(n3425), .Y(P1_U3533));
  NAND2X1 g2373(.A(n3404), .B(P1_REG1_REG_11__SCAN_IN), .Y(n3427));
  OAI21X1 g2374(.A0(n3404), .A1(n2598), .B0(n3427), .Y(P1_U3534));
  NAND2X1 g2375(.A(n3404), .B(P1_REG1_REG_12__SCAN_IN), .Y(n3429));
  OAI21X1 g2376(.A0(n3404), .A1(n2639), .B0(n3429), .Y(P1_U3535));
  NAND2X1 g2377(.A(n3404), .B(P1_REG1_REG_13__SCAN_IN), .Y(n3431));
  OAI21X1 g2378(.A0(n3404), .A1(n2686), .B0(n3431), .Y(P1_U3536));
  NAND2X1 g2379(.A(n3404), .B(P1_REG1_REG_14__SCAN_IN), .Y(n3433));
  OAI21X1 g2380(.A0(n3404), .A1(n2730), .B0(n3433), .Y(P1_U3537));
  NAND2X1 g2381(.A(n3404), .B(P1_REG1_REG_15__SCAN_IN), .Y(n3435));
  OAI21X1 g2382(.A0(n3404), .A1(n2769), .B0(n3435), .Y(P1_U3538));
  NAND2X1 g2383(.A(n3404), .B(P1_REG1_REG_16__SCAN_IN), .Y(n3437));
  OAI21X1 g2384(.A0(n3404), .A1(n2816), .B0(n3437), .Y(P1_U3539));
  NAND2X1 g2385(.A(n3404), .B(P1_REG1_REG_17__SCAN_IN), .Y(n3439));
  OAI21X1 g2386(.A0(n3404), .A1(n2868), .B0(n3439), .Y(P1_U3540));
  NAND2X1 g2387(.A(n3404), .B(P1_REG1_REG_18__SCAN_IN), .Y(n3441));
  OAI21X1 g2388(.A0(n3404), .A1(n2910), .B0(n3441), .Y(P1_U3541));
  NAND2X1 g2389(.A(n3404), .B(P1_REG1_REG_19__SCAN_IN), .Y(n3443));
  OAI21X1 g2390(.A0(n3404), .A1(n2953), .B0(n3443), .Y(P1_U3542));
  NAND2X1 g2391(.A(n3404), .B(P1_REG1_REG_20__SCAN_IN), .Y(n3445));
  OAI21X1 g2392(.A0(n3404), .A1(n2997), .B0(n3445), .Y(P1_U3543));
  NAND2X1 g2393(.A(n3404), .B(P1_REG1_REG_21__SCAN_IN), .Y(n3447));
  OAI21X1 g2394(.A0(n3404), .A1(n3039), .B0(n3447), .Y(P1_U3544));
  NAND2X1 g2395(.A(n3404), .B(P1_REG1_REG_22__SCAN_IN), .Y(n3449));
  OAI21X1 g2396(.A0(n3404), .A1(n3076), .B0(n3449), .Y(P1_U3545));
  NAND2X1 g2397(.A(n3404), .B(P1_REG1_REG_23__SCAN_IN), .Y(n3451));
  OAI21X1 g2398(.A0(n3404), .A1(n3120), .B0(n3451), .Y(P1_U3546));
  NAND2X1 g2399(.A(n3404), .B(P1_REG1_REG_24__SCAN_IN), .Y(n3453));
  OAI21X1 g2400(.A0(n3404), .A1(n3163), .B0(n3453), .Y(P1_U3547));
  NAND2X1 g2401(.A(n3404), .B(P1_REG1_REG_25__SCAN_IN), .Y(n3455));
  OAI21X1 g2402(.A0(n3404), .A1(n3203), .B0(n3455), .Y(P1_U3548));
  NAND2X1 g2403(.A(n3404), .B(P1_REG1_REG_26__SCAN_IN), .Y(n3457));
  OAI21X1 g2404(.A0(n3404), .A1(n3246), .B0(n3457), .Y(P1_U3549));
  NAND2X1 g2405(.A(n3404), .B(P1_REG1_REG_27__SCAN_IN), .Y(n3459));
  OAI21X1 g2406(.A0(n3404), .A1(n3294), .B0(n3459), .Y(P1_U3550));
  NAND2X1 g2407(.A(n3404), .B(P1_REG1_REG_28__SCAN_IN), .Y(n3461));
  OAI21X1 g2408(.A0(n3404), .A1(n3333), .B0(n3461), .Y(P1_U3551));
  NAND2X1 g2409(.A(n3404), .B(P1_REG1_REG_29__SCAN_IN), .Y(n3463));
  OAI21X1 g2410(.A0(n3404), .A1(n3376), .B0(n3463), .Y(P1_U3552));
  NAND2X1 g2411(.A(n3404), .B(P1_REG1_REG_30__SCAN_IN), .Y(n3465));
  OAI21X1 g2412(.A0(n3404), .A1(n3388), .B0(n3465), .Y(P1_U3553));
  NAND2X1 g2413(.A(n3404), .B(P1_REG1_REG_31__SCAN_IN), .Y(n3467));
  OAI21X1 g2414(.A0(n3404), .A1(n3400), .B0(n3467), .Y(P1_U3554));
  NOR4X1  g2415(.A(n1991), .B(n2027), .C(n1985), .D(n1993), .Y(n3469));
  INVX1   g2416(.A(n3469), .Y(n3470));
  INVX1   g2417(.A(n1982), .Y(n3471));
  NOR2X1  g2418(.A(n1989), .B(n1984), .Y(n3472));
  INVX1   g2419(.A(n3472), .Y(n3473));
  AOI21X1 g2420(.A0(n1993), .A1(n1987), .B0(n3473), .Y(n3474));
  INVX1   g2421(.A(n3474), .Y(n3475));
  NAND4X1 g2422(.A(n1999), .B(n3471), .C(n1979), .D(n3475), .Y(n3476));
  NAND2X1 g2423(.A(n3476), .B(n3470), .Y(n3477));
  NAND4X1 g2424(.A(n2062), .B(n2054), .C(n1893), .D(n3477), .Y(n3478));
  NAND2X1 g2425(.A(n3477), .B(n1893), .Y(n3479));
  INVX1   g2426(.A(n3479), .Y(n3480));
  AOI21X1 g2427(.A0(n3477), .A1(n1893), .B0(n2018), .Y(n3481));
  AOI21X1 g2428(.A0(n3480), .A1(n2051), .B0(n3481), .Y(n3482));
  INVX1   g2429(.A(n2026), .Y(n3483));
  NAND3X1 g2430(.A(n1989), .B(n2027), .C(n1984), .Y(n3484));
  NOR2X1  g2431(.A(n3484), .B(n3479), .Y(n3485));
  NOR4X1  g2432(.A(n1993), .B(n1989), .C(n2027), .D(n3479), .Y(n3486));
  AOI22X1 g2433(.A0(n3485), .A1(n2035), .B0(n3483), .B1(n3486), .Y(n3487));
  NOR4X1  g2434(.A(n1991), .B(n2027), .C(n1985), .D(n2041), .Y(n3488));
  INVX1   g2435(.A(n3488), .Y(n3489));
  NOR2X1  g2436(.A(n3489), .B(n3479), .Y(n3490));
  NOR2X1  g2437(.A(n3479), .B(n3470), .Y(n3491));
  AOI22X1 g2438(.A0(n3490), .A1(n2035), .B0(P1_REG3_REG_0__SCAN_IN), .B1(n3491), .Y(n3492));
  NAND4X1 g2439(.A(n3487), .B(n3482), .C(n3478), .D(n3492), .Y(P1_U3291));
  NAND4X1 g2440(.A(n2110), .B(n2054), .C(n1893), .D(n3477), .Y(n3494));
  AOI21X1 g2441(.A0(n3477), .A1(n1893), .B0(n2055), .Y(n3495));
  AOI21X1 g2442(.A0(n3480), .A1(n2096), .B0(n3495), .Y(n3496));
  AOI22X1 g2443(.A0(n3485), .A1(n2081), .B0(n2086), .B1(n3486), .Y(n3497));
  AOI22X1 g2444(.A0(n3490), .A1(n2103), .B0(P1_REG3_REG_1__SCAN_IN), .B1(n3491), .Y(n3498));
  NAND4X1 g2445(.A(n3497), .B(n3496), .C(n3494), .D(n3498), .Y(P1_U3290));
  NAND4X1 g2446(.A(n2167), .B(n2054), .C(n1893), .D(n3477), .Y(n3500));
  AOI22X1 g2447(.A0(n3485), .A1(n2122), .B0(n2143), .B1(n3490), .Y(n3501));
  INVX1   g2448(.A(P1_REG2_REG_2__SCAN_IN), .Y(n3502));
  AOI21X1 g2449(.A0(n3477), .A1(n1893), .B0(n3502), .Y(n3503));
  AOI21X1 g2450(.A0(n3480), .A1(n2138), .B0(n3503), .Y(n3504));
  AOI22X1 g2451(.A0(n3486), .A1(n2129), .B0(P1_REG3_REG_2__SCAN_IN), .B1(n3491), .Y(n3505));
  NAND4X1 g2452(.A(n3504), .B(n3501), .C(n3500), .D(n3505), .Y(P1_U3289));
  INVX1   g2453(.A(P1_REG3_REG_3__SCAN_IN), .Y(n3507));
  AOI22X1 g2454(.A0(n3486), .A1(n2180), .B0(n3507), .B1(n3491), .Y(n3508));
  AOI22X1 g2455(.A0(n3485), .A1(n2172), .B0(n2201), .B1(n3490), .Y(n3509));
  NAND2X1 g2456(.A(n3480), .B(n2199), .Y(n3510));
  NOR2X1  g2457(.A(n3479), .B(n2104), .Y(n3511));
  AOI22X1 g2458(.A0(n3479), .A1(P1_REG2_REG_3__SCAN_IN), .B0(n2208), .B1(n3511), .Y(n3512));
  NAND4X1 g2459(.A(n3510), .B(n3509), .C(n3508), .D(n3512), .Y(P1_U3288));
  NOR3X1  g2460(.A(n2251), .B(n2247), .C(n2238), .Y(n3514));
  INVX1   g2461(.A(P1_REG2_REG_4__SCAN_IN), .Y(n3515));
  INVX1   g2462(.A(n3511), .Y(n3516));
  OAI22X1 g2463(.A0(n3480), .A1(n3515), .B0(n2263), .B1(n3516), .Y(n3517));
  INVX1   g2464(.A(n3486), .Y(n3518));
  INVX1   g2465(.A(n3491), .Y(n3519));
  OAI22X1 g2466(.A0(n3518), .A1(n2237), .B0(n2205), .B1(n3519), .Y(n3520));
  INVX1   g2467(.A(n3485), .Y(n3521));
  NAND4X1 g2468(.A(n3477), .B(n2253), .C(n1893), .D(n3488), .Y(n3522));
  OAI21X1 g2469(.A0(n3521), .A1(n2223), .B0(n3522), .Y(n3523));
  NOR3X1  g2470(.A(n3523), .B(n3520), .C(n3517), .Y(n3524));
  OAI21X1 g2471(.A0(n3479), .A1(n3514), .B0(n3524), .Y(P1_U3287));
  NAND2X1 g2472(.A(n3480), .B(n2305), .Y(n3526));
  OAI22X1 g2473(.A0(n3480), .A1(n2254), .B0(n2338), .B1(n3516), .Y(n3527));
  OAI22X1 g2474(.A0(n3518), .A1(n2289), .B0(n2259), .B1(n3519), .Y(n3528));
  INVX1   g2475(.A(n3490), .Y(n3529));
  OAI22X1 g2476(.A0(n3521), .A1(n2284), .B0(n2308), .B1(n3529), .Y(n3530));
  NOR3X1  g2477(.A(n3530), .B(n3528), .C(n3527), .Y(n3531));
  NAND2X1 g2478(.A(n3531), .B(n3526), .Y(P1_U3286));
  NOR3X1  g2479(.A(n2355), .B(n2347), .C(n2346), .Y(n3533));
  OAI22X1 g2480(.A0(n3480), .A1(n2335), .B0(n2366), .B1(n3516), .Y(n3534));
  OAI22X1 g2481(.A0(n3518), .A1(n2345), .B0(n2313), .B1(n3519), .Y(n3535));
  NAND4X1 g2482(.A(n3477), .B(n2357), .C(n1893), .D(n3488), .Y(n3536));
  OAI21X1 g2483(.A0(n3521), .A1(n2332), .B0(n3536), .Y(n3537));
  NOR3X1  g2484(.A(n3537), .B(n3535), .C(n3534), .Y(n3538));
  OAI21X1 g2485(.A0(n3479), .A1(n3533), .B0(n3538), .Y(P1_U3285));
  NOR3X1  g2486(.A(n2400), .B(n2390), .C(n2389), .Y(n3540));
  AOI22X1 g2487(.A0(n3490), .A1(n2402), .B0(n2363), .B1(n3491), .Y(n3541));
  OAI21X1 g2488(.A0(n3521), .A1(n2379), .B0(n3541), .Y(n3542));
  AOI22X1 g2489(.A0(n3479), .A1(P1_REG2_REG_7__SCAN_IN), .B0(n2410), .B1(n3511), .Y(n3543));
  OAI21X1 g2490(.A0(n3518), .A1(n2388), .B0(n3543), .Y(n3544));
  NOR2X1  g2491(.A(n3544), .B(n3542), .Y(n3545));
  OAI21X1 g2492(.A0(n3479), .A1(n3540), .B0(n3545), .Y(P1_U3284));
  NOR3X1  g2493(.A(n2443), .B(n2432), .C(n2431), .Y(n3547));
  NOR2X1  g2494(.A(n3518), .B(n2430), .Y(n3548));
  AOI22X1 g2495(.A0(n3479), .A1(P1_REG2_REG_8__SCAN_IN), .B0(n2453), .B1(n3511), .Y(n3549));
  INVX1   g2496(.A(n3484), .Y(n3550));
  NAND4X1 g2497(.A(n3477), .B(n2425), .C(n1893), .D(n3550), .Y(n3551));
  AOI22X1 g2498(.A0(n3490), .A1(n2446), .B0(n2408), .B1(n3491), .Y(n3552));
  NAND3X1 g2499(.A(n3552), .B(n3551), .C(n3549), .Y(n3553));
  NOR2X1  g2500(.A(n3553), .B(n3548), .Y(n3554));
  OAI21X1 g2501(.A0(n3479), .A1(n3547), .B0(n3554), .Y(P1_U3283));
  NAND2X1 g2502(.A(n3480), .B(n2488), .Y(n3556));
  AOI22X1 g2503(.A0(n3479), .A1(P1_REG2_REG_9__SCAN_IN), .B0(n2469), .B1(n3485), .Y(n3557));
  NAND4X1 g2504(.A(n3469), .B(n2450), .C(n1893), .D(n3477), .Y(n3558));
  AOI22X1 g2505(.A0(n3511), .A1(n2498), .B0(n2490), .B1(n3490), .Y(n3559));
  NAND3X1 g2506(.A(n3559), .B(n3558), .C(n3557), .Y(n3560));
  AOI21X1 g2507(.A0(n3486), .A1(n2474), .B0(n3560), .Y(n3561));
  NAND2X1 g2508(.A(n3561), .B(n3556), .Y(P1_U3282));
  NOR3X1  g2509(.A(n2534), .B(n2525), .C(n2524), .Y(n3563));
  NAND2X1 g2510(.A(n3490), .B(n2538), .Y(n3564));
  AOI22X1 g2511(.A0(n3479), .A1(P1_REG2_REG_10__SCAN_IN), .B0(n2511), .B1(n3485), .Y(n3565));
  AOI22X1 g2512(.A0(n3511), .A1(n2545), .B0(n2495), .B1(n3491), .Y(n3566));
  NAND3X1 g2513(.A(n3566), .B(n3565), .C(n3564), .Y(n3567));
  AOI21X1 g2514(.A0(n3486), .A1(n2522), .B0(n3567), .Y(n3568));
  OAI21X1 g2515(.A0(n3479), .A1(n3563), .B0(n3568), .Y(P1_U3281));
  NOR2X1  g2516(.A(n2570), .B(n2184), .Y(n3570));
  INVX1   g2517(.A(n2582), .Y(n3571));
  NOR4X1  g2518(.A(n2584), .B(n3571), .C(n3570), .D(n2585), .Y(n3572));
  NOR2X1  g2519(.A(n3518), .B(n2578), .Y(n3573));
  NAND2X1 g2520(.A(n3490), .B(n2587), .Y(n3574));
  AOI22X1 g2521(.A0(n3479), .A1(P1_REG2_REG_11__SCAN_IN), .B0(n2593), .B1(n3511), .Y(n3575));
  AOI22X1 g2522(.A0(n3485), .A1(n2562), .B0(n2541), .B1(n3491), .Y(n3576));
  NAND3X1 g2523(.A(n3576), .B(n3575), .C(n3574), .Y(n3577));
  NOR2X1  g2524(.A(n3577), .B(n3573), .Y(n3578));
  OAI21X1 g2525(.A0(n3479), .A1(n3572), .B0(n3578), .Y(P1_U3280));
  NAND2X1 g2526(.A(n3480), .B(n2625), .Y(n3580));
  NAND2X1 g2527(.A(n3490), .B(n2628), .Y(n3581));
  AOI22X1 g2528(.A0(n3479), .A1(P1_REG2_REG_12__SCAN_IN), .B0(n2634), .B1(n3511), .Y(n3582));
  AOI22X1 g2529(.A0(n3485), .A1(n2607), .B0(n2590), .B1(n3491), .Y(n3583));
  NAND3X1 g2530(.A(n3583), .B(n3582), .C(n3581), .Y(n3584));
  AOI21X1 g2531(.A0(n3486), .A1(n2612), .B0(n3584), .Y(n3585));
  NAND2X1 g2532(.A(n3585), .B(n3580), .Y(P1_U3279));
  NOR3X1  g2533(.A(n2669), .B(n2660), .C(n2659), .Y(n3587));
  NAND2X1 g2534(.A(n3490), .B(n2672), .Y(n3588));
  AOI22X1 g2535(.A0(n3479), .A1(P1_REG2_REG_13__SCAN_IN), .B0(n2681), .B1(n3511), .Y(n3589));
  AOI22X1 g2536(.A0(n3485), .A1(n2649), .B0(n2631), .B1(n3491), .Y(n3590));
  NAND3X1 g2537(.A(n3590), .B(n3589), .C(n3588), .Y(n3591));
  AOI21X1 g2538(.A0(n3486), .A1(n2657), .B0(n3591), .Y(n3592));
  OAI21X1 g2539(.A0(n3479), .A1(n3587), .B0(n3592), .Y(P1_U3278));
  INVX1   g2540(.A(P1_REG2_REG_14__SCAN_IN), .Y(n3594));
  OAI22X1 g2541(.A0(n3480), .A1(n3594), .B0(n2726), .B1(n3516), .Y(n3595));
  OAI22X1 g2542(.A0(n3521), .A1(n2693), .B0(n2676), .B1(n3519), .Y(n3596));
  NOR2X1  g2543(.A(n3596), .B(n3595), .Y(n3597));
  OAI21X1 g2544(.A0(n3529), .A1(n2717), .B0(n3597), .Y(n3598));
  AOI21X1 g2545(.A0(n3486), .A1(n2706), .B0(n3598), .Y(n3599));
  OAI21X1 g2546(.A0(n3479), .A1(n2712), .B0(n3599), .Y(P1_U3277));
  NAND2X1 g2547(.A(n3490), .B(n2758), .Y(n3601));
  AOI22X1 g2548(.A0(n3479), .A1(P1_REG2_REG_15__SCAN_IN), .B0(n2757), .B1(n3485), .Y(n3602));
  AOI22X1 g2549(.A0(n3511), .A1(n2764), .B0(n2722), .B1(n3491), .Y(n3603));
  NAND3X1 g2550(.A(n3603), .B(n3602), .C(n3601), .Y(n3604));
  AOI21X1 g2551(.A0(n3486), .A1(n2748), .B0(n3604), .Y(n3605));
  OAI21X1 g2552(.A0(n3479), .A1(n2754), .B0(n3605), .Y(P1_U3276));
  NOR3X1  g2553(.A(n2802), .B(n2801), .C(n2800), .Y(n3607));
  NAND2X1 g2554(.A(n3490), .B(n2804), .Y(n3608));
  AOI22X1 g2555(.A0(n3479), .A1(P1_REG2_REG_16__SCAN_IN), .B0(n2784), .B1(n3485), .Y(n3609));
  AOI22X1 g2556(.A0(n3511), .A1(n2811), .B0(n2760), .B1(n3491), .Y(n3610));
  NAND3X1 g2557(.A(n3610), .B(n3609), .C(n3608), .Y(n3611));
  AOI21X1 g2558(.A0(n3486), .A1(n2797), .B0(n3611), .Y(n3612));
  OAI21X1 g2559(.A0(n3479), .A1(n3607), .B0(n3612), .Y(P1_U3275));
  NAND2X1 g2560(.A(n3480), .B(n2854), .Y(n3614));
  NAND3X1 g2561(.A(n3486), .B(n2835), .C(n2829), .Y(n3615));
  NAND2X1 g2562(.A(n3490), .B(n2856), .Y(n3616));
  AOI22X1 g2563(.A0(n3479), .A1(P1_REG2_REG_17__SCAN_IN), .B0(n2863), .B1(n3511), .Y(n3617));
  OAI21X1 g2564(.A0(n3519), .A1(n2806), .B0(n3617), .Y(n3618));
  AOI21X1 g2565(.A0(n3485), .A1(n2825), .B0(n3618), .Y(n3619));
  NAND4X1 g2566(.A(n3616), .B(n3615), .C(n3614), .D(n3619), .Y(P1_U3274));
  NAND2X1 g2567(.A(n3480), .B(n2896), .Y(n3621));
  NAND2X1 g2568(.A(n3486), .B(n2886), .Y(n3622));
  NAND2X1 g2569(.A(n3490), .B(n2899), .Y(n3623));
  AOI22X1 g2570(.A0(n3479), .A1(P1_REG2_REG_18__SCAN_IN), .B0(n2926), .B1(n3511), .Y(n3624));
  OAI21X1 g2571(.A0(n3519), .A1(n2858), .B0(n3624), .Y(n3625));
  AOI21X1 g2572(.A0(n3485), .A1(n2898), .B0(n3625), .Y(n3626));
  NAND4X1 g2573(.A(n3623), .B(n3622), .C(n3621), .D(n3626), .Y(P1_U3273));
  NAND2X1 g2574(.A(n3480), .B(n2936), .Y(n3628));
  NOR2X1  g2575(.A(n2927), .B(n2972), .Y(n3629));
  OAI21X1 g2576(.A0(n3629), .A1(n2925), .B0(n3486), .Y(n3630));
  NAND2X1 g2577(.A(n3490), .B(n2940), .Y(n3631));
  AOI22X1 g2578(.A0(n3479), .A1(P1_REG2_REG_19__SCAN_IN), .B0(n2902), .B1(n3491), .Y(n3632));
  OAI21X1 g2579(.A0(n3516), .A1(n2949), .B0(n3632), .Y(n3633));
  AOI21X1 g2580(.A0(n3485), .A1(n2914), .B0(n3633), .Y(n3634));
  NAND4X1 g2581(.A(n3631), .B(n3630), .C(n3628), .D(n3634), .Y(P1_U3272));
  NAND2X1 g2582(.A(n3480), .B(n2982), .Y(n3636));
  INVX1   g2583(.A(n2944), .Y(n3637));
  AOI22X1 g2584(.A0(n3479), .A1(P1_REG2_REG_20__SCAN_IN), .B0(n3637), .B1(n3491), .Y(n3638));
  OAI21X1 g2585(.A0(n3516), .A1(n2993), .B0(n3638), .Y(n3639));
  AOI21X1 g2586(.A0(n3485), .A1(n2956), .B0(n3639), .Y(n3640));
  OAI21X1 g2587(.A0(n3529), .A1(n2985), .B0(n3640), .Y(n3641));
  AOI21X1 g2588(.A0(n3486), .A1(n2976), .B0(n3641), .Y(n3642));
  NAND2X1 g2589(.A(n3642), .B(n3636), .Y(P1_U3271));
  NAND2X1 g2590(.A(n3480), .B(n3026), .Y(n3644));
  INVX1   g2591(.A(n3019), .Y(n3645));
  NAND2X1 g2592(.A(n3486), .B(n3645), .Y(n3646));
  NAND2X1 g2593(.A(n3490), .B(n3029), .Y(n3647));
  AOI22X1 g2594(.A0(n3479), .A1(P1_REG2_REG_21__SCAN_IN), .B0(n2989), .B1(n3491), .Y(n3648));
  OAI21X1 g2595(.A0(n3516), .A1(n3035), .B0(n3648), .Y(n3649));
  AOI21X1 g2596(.A0(n3485), .A1(n3000), .B0(n3649), .Y(n3650));
  NAND4X1 g2597(.A(n3647), .B(n3646), .C(n3644), .D(n3650), .Y(P1_U3270));
  NOR3X1  g2598(.A(n3062), .B(n3061), .C(n3060), .Y(n3652));
  NOR2X1  g2599(.A(n3518), .B(n3056), .Y(n3653));
  NAND2X1 g2600(.A(n3490), .B(n3065), .Y(n3654));
  AOI22X1 g2601(.A0(n3479), .A1(P1_REG2_REG_22__SCAN_IN), .B0(n3031), .B1(n3491), .Y(n3655));
  OAI21X1 g2602(.A0(n3516), .A1(n3072), .B0(n3655), .Y(n3656));
  AOI21X1 g2603(.A0(n3485), .A1(n3042), .B0(n3656), .Y(n3657));
  NAND2X1 g2604(.A(n3657), .B(n3654), .Y(n3658));
  NOR2X1  g2605(.A(n3658), .B(n3653), .Y(n3659));
  OAI21X1 g2606(.A0(n3479), .A1(n3652), .B0(n3659), .Y(P1_U3269));
  NAND2X1 g2607(.A(n3480), .B(n3107), .Y(n3661));
  NOR2X1  g2608(.A(n3518), .B(n3100), .Y(n3662));
  INVX1   g2609(.A(n3067), .Y(n3663));
  AOI22X1 g2610(.A0(n3479), .A1(P1_REG2_REG_23__SCAN_IN), .B0(n3663), .B1(n3491), .Y(n3664));
  OAI21X1 g2611(.A0(n3516), .A1(n3123), .B0(n3664), .Y(n3665));
  AOI21X1 g2612(.A0(n3485), .A1(n3111), .B0(n3665), .Y(n3666));
  OAI21X1 g2613(.A0(n3529), .A1(n3110), .B0(n3666), .Y(n3667));
  NOR2X1  g2614(.A(n3667), .B(n3662), .Y(n3668));
  NAND2X1 g2615(.A(n3668), .B(n3661), .Y(P1_U3268));
  NOR3X1  g2616(.A(n3148), .B(n3145), .C(n3134), .Y(n3670));
  NAND2X1 g2617(.A(n3490), .B(n3152), .Y(n3671));
  INVX1   g2618(.A(n3113), .Y(n3672));
  AOI22X1 g2619(.A0(n3479), .A1(P1_REG2_REG_24__SCAN_IN), .B0(n3672), .B1(n3491), .Y(n3673));
  OAI21X1 g2620(.A0(n3516), .A1(n3159), .B0(n3673), .Y(n3674));
  AOI21X1 g2621(.A0(n3485), .A1(n3124), .B0(n3674), .Y(n3675));
  NAND2X1 g2622(.A(n3675), .B(n3671), .Y(n3676));
  AOI21X1 g2623(.A0(n3486), .A1(n3142), .B0(n3676), .Y(n3677));
  OAI21X1 g2624(.A0(n3479), .A1(n3670), .B0(n3677), .Y(P1_U3267));
  NOR3X1  g2625(.A(n3188), .B(n3187), .C(n3186), .Y(n3679));
  NOR2X1  g2626(.A(n3518), .B(n3182), .Y(n3680));
  NAND2X1 g2627(.A(n3490), .B(n3190), .Y(n3681));
  INVX1   g2628(.A(n3154), .Y(n3682));
  AOI22X1 g2629(.A0(n3479), .A1(P1_REG2_REG_25__SCAN_IN), .B0(n3682), .B1(n3491), .Y(n3683));
  OAI21X1 g2630(.A0(n3516), .A1(n3199), .B0(n3683), .Y(n3684));
  AOI21X1 g2631(.A0(n3485), .A1(n3166), .B0(n3684), .Y(n3685));
  NAND2X1 g2632(.A(n3685), .B(n3681), .Y(n3686));
  NOR2X1  g2633(.A(n3686), .B(n3680), .Y(n3687));
  OAI21X1 g2634(.A0(n3479), .A1(n3679), .B0(n3687), .Y(P1_U3266));
  NOR4X1  g2635(.A(n3229), .B(n3227), .C(n3214), .D(n3230), .Y(n3689));
  INVX1   g2636(.A(n3194), .Y(n3690));
  AOI22X1 g2637(.A0(n3479), .A1(P1_REG2_REG_26__SCAN_IN), .B0(n3690), .B1(n3491), .Y(n3691));
  OAI21X1 g2638(.A0(n3516), .A1(n3253), .B0(n3691), .Y(n3692));
  AOI21X1 g2639(.A0(n3485), .A1(n3206), .B0(n3692), .Y(n3693));
  OAI21X1 g2640(.A0(n3529), .A1(n3236), .B0(n3693), .Y(n3694));
  AOI21X1 g2641(.A0(n3486), .A1(n3224), .B0(n3694), .Y(n3695));
  OAI21X1 g2642(.A0(n3479), .A1(n3689), .B0(n3695), .Y(P1_U3265));
  NOR3X1  g2643(.A(n3278), .B(n3277), .C(n3275), .Y(n3697));
  NAND2X1 g2644(.A(n3490), .B(n3282), .Y(n3698));
  INVX1   g2645(.A(n3239), .Y(n3699));
  AOI22X1 g2646(.A0(n3479), .A1(P1_REG2_REG_27__SCAN_IN), .B0(n3699), .B1(n3491), .Y(n3700));
  OAI21X1 g2647(.A0(n3516), .A1(n3290), .B0(n3700), .Y(n3701));
  AOI21X1 g2648(.A0(n3485), .A1(n3255), .B0(n3701), .Y(n3702));
  NAND2X1 g2649(.A(n3702), .B(n3698), .Y(n3703));
  AOI21X1 g2650(.A0(n3486), .A1(n3272), .B0(n3703), .Y(n3704));
  OAI21X1 g2651(.A0(n3479), .A1(n3697), .B0(n3704), .Y(P1_U3264));
  OAI21X1 g2652(.A0(n3317), .A1(n3314), .B0(n3480), .Y(n3706));
  NOR2X1  g2653(.A(n3518), .B(n3310), .Y(n3707));
  NAND2X1 g2654(.A(n3490), .B(n3319), .Y(n3708));
  INVX1   g2655(.A(n3285), .Y(n3709));
  AOI22X1 g2656(.A0(n3479), .A1(P1_REG2_REG_28__SCAN_IN), .B0(n3709), .B1(n3491), .Y(n3710));
  OAI21X1 g2657(.A0(n3516), .A1(n3329), .B0(n3710), .Y(n3711));
  AOI21X1 g2658(.A0(n3485), .A1(n3297), .B0(n3711), .Y(n3712));
  NAND2X1 g2659(.A(n3712), .B(n3708), .Y(n3713));
  NOR2X1  g2660(.A(n3713), .B(n3707), .Y(n3714));
  NAND2X1 g2661(.A(n3714), .B(n3706), .Y(P1_U3263));
  OAI21X1 g2662(.A0(n3368), .A1(n3356), .B0(n3480), .Y(n3716));
  NAND2X1 g2663(.A(n3479), .B(P1_REG2_REG_29__SCAN_IN), .Y(n3717));
  NAND4X1 g2664(.A(n3238), .B(P1_REG3_REG_27__SCAN_IN), .C(P1_REG3_REG_28__SCAN_IN), .D(n3491), .Y(n3718));
  NAND2X1 g2665(.A(n3718), .B(n3717), .Y(n3719));
  AOI21X1 g2666(.A0(n3485), .A1(n3345), .B0(n3719), .Y(n3720));
  OAI21X1 g2667(.A0(n3529), .A1(n3374), .B0(n3720), .Y(n3721));
  AOI21X1 g2668(.A0(n3486), .A1(n3347), .B0(n3721), .Y(n3722));
  NAND2X1 g2669(.A(n3722), .B(n3716), .Y(P1_U3355));
  NAND2X1 g2670(.A(n3490), .B(n3381), .Y(n3724));
  INVX1   g2671(.A(n1831), .Y(n3725));
  NAND2X1 g2672(.A(n1836), .B(n1834), .Y(n3726));
  XOR2X1  g2673(.A(n1839), .B(n3726), .Y(n3727));
  OAI21X1 g2674(.A0(n3727), .A1(n1156), .B0(n3725), .Y(n3728));
  NAND3X1 g2675(.A(n3485), .B(n2101), .C(n3728), .Y(n3729));
  NAND4X1 g2676(.A(n3385), .B(n3350), .C(n1893), .D(n3477), .Y(n3730));
  NAND2X1 g2677(.A(n3479), .B(P1_REG2_REG_30__SCAN_IN), .Y(n3731));
  NAND4X1 g2678(.A(n3730), .B(n3729), .C(n3724), .D(n3731), .Y(P1_U3262));
  NAND2X1 g2679(.A(n3490), .B(n3397), .Y(n3733));
  NAND2X1 g2680(.A(n3485), .B(n3396), .Y(n3734));
  NAND2X1 g2681(.A(n3479), .B(P1_REG2_REG_31__SCAN_IN), .Y(n3735));
  NAND4X1 g2682(.A(n3734), .B(n3733), .C(n3730), .D(n3735), .Y(P1_U3261));
  OAI21X1 g2683(.A0(n3472), .A1(n1884), .B0(n1874), .Y(n3737));
  NAND2X1 g2684(.A(n3737), .B(n2101), .Y(n3738));
  NOR4X1  g2685(.A(n1884), .B(n1875), .C(P1_U3084), .D(n3738), .Y(n3739));
  INVX1   g2686(.A(P1_REG2_REG_18__SCAN_IN), .Y(n3740));
  INVX1   g2687(.A(P1_REG2_REG_16__SCAN_IN), .Y(n3741));
  INVX1   g2688(.A(P1_REG2_REG_17__SCAN_IN), .Y(n3742));
  AOI22X1 g2689(.A0(n2776), .A1(n3741), .B0(n3742), .B1(n2821), .Y(n3743));
  NOR2X1  g2690(.A(n2735), .B(P1_REG2_REG_15__SCAN_IN), .Y(n3744));
  INVX1   g2691(.A(P1_REG2_REG_13__SCAN_IN), .Y(n3745));
  NAND2X1 g2692(.A(n2646), .B(n3745), .Y(n3746));
  INVX1   g2693(.A(P1_REG2_REG_11__SCAN_IN), .Y(n3747));
  NOR2X1  g2694(.A(n2559), .B(n3747), .Y(n3748));
  INVX1   g2695(.A(n3748), .Y(n3749));
  INVX1   g2696(.A(P1_REG2_REG_12__SCAN_IN), .Y(n3750));
  AOI22X1 g2697(.A0(n2604), .A1(n3750), .B0(n3745), .B1(n2646), .Y(n3751));
  INVX1   g2698(.A(n3751), .Y(n3752));
  NOR2X1  g2699(.A(n2604), .B(n3750), .Y(n3753));
  AOI21X1 g2700(.A0(n2647), .A1(P1_REG2_REG_13__SCAN_IN), .B0(n3753), .Y(n3754));
  OAI21X1 g2701(.A0(n3752), .A1(n3749), .B0(n3754), .Y(n3755));
  INVX1   g2702(.A(P1_REG2_REG_10__SCAN_IN), .Y(n3756));
  INVX1   g2703(.A(P1_REG2_REG_8__SCAN_IN), .Y(n3757));
  NOR2X1  g2704(.A(n2422), .B(n3757), .Y(n3758));
  INVX1   g2705(.A(P1_REG2_REG_9__SCAN_IN), .Y(n3759));
  AOI22X1 g2706(.A0(n2466), .A1(n3759), .B0(n3756), .B1(n2508), .Y(n3760));
  NAND2X1 g2707(.A(n2467), .B(P1_REG2_REG_9__SCAN_IN), .Y(n3761));
  OAI21X1 g2708(.A0(n2508), .A1(n3756), .B0(n3761), .Y(n3762));
  AOI21X1 g2709(.A0(n3760), .A1(n3758), .B0(n3762), .Y(n3763));
  AOI21X1 g2710(.A0(n2508), .A1(n3756), .B0(n3763), .Y(n3764));
  OAI22X1 g2711(.A0(n2330), .A1(P1_REG2_REG_6__SCAN_IN), .B0(P1_REG2_REG_7__SCAN_IN), .B1(n2377), .Y(n3765));
  AOI22X1 g2712(.A0(n2219), .A1(n3515), .B0(n2254), .B1(n2276), .Y(n3766));
  AOI22X1 g2713(.A0(n2119), .A1(n3502), .B0(n2144), .B1(n2169), .Y(n3767));
  INVX1   g2714(.A(n2078), .Y(n3768));
  AOI21X1 g2715(.A0(n2007), .A1(n2006), .B0(n2018), .Y(n3769));
  OAI21X1 g2716(.A0(n3768), .A1(P1_REG2_REG_1__SCAN_IN), .B0(n3769), .Y(n3770));
  INVX1   g2717(.A(n3770), .Y(n3771));
  NOR2X1  g2718(.A(n2078), .B(n2055), .Y(n3772));
  OAI21X1 g2719(.A0(n3772), .A1(n3771), .B0(n3767), .Y(n3773));
  NOR2X1  g2720(.A(n2169), .B(n2144), .Y(n3774));
  INVX1   g2721(.A(n3774), .Y(n3775));
  NOR2X1  g2722(.A(n2119), .B(n3502), .Y(n3776));
  OAI21X1 g2723(.A0(n2170), .A1(P1_REG2_REG_3__SCAN_IN), .B0(n3776), .Y(n3777));
  NAND3X1 g2724(.A(n3777), .B(n3775), .C(n3773), .Y(n3778));
  NAND2X1 g2725(.A(n3778), .B(n3766), .Y(n3779));
  NOR2X1  g2726(.A(n2219), .B(n3515), .Y(n3780));
  INVX1   g2727(.A(n3780), .Y(n3781));
  AOI21X1 g2728(.A0(n3781), .A1(n2254), .B0(n2276), .Y(n3782));
  AOI21X1 g2729(.A0(n3780), .A1(P1_REG2_REG_5__SCAN_IN), .B0(n3782), .Y(n3783));
  NAND2X1 g2730(.A(n3783), .B(n3779), .Y(n3784));
  INVX1   g2731(.A(n3784), .Y(n3785));
  NOR2X1  g2732(.A(n2329), .B(n2335), .Y(n3786));
  INVX1   g2733(.A(P1_REG2_REG_7__SCAN_IN), .Y(n3787));
  INVX1   g2734(.A(n3786), .Y(n3788));
  AOI21X1 g2735(.A0(n3788), .A1(n3787), .B0(n2376), .Y(n3789));
  AOI21X1 g2736(.A0(n3786), .A1(P1_REG2_REG_7__SCAN_IN), .B0(n3789), .Y(n3790));
  OAI21X1 g2737(.A0(n3785), .A1(n3765), .B0(n3790), .Y(n3791));
  NOR2X1  g2738(.A(n2423), .B(P1_REG2_REG_8__SCAN_IN), .Y(n3792));
  INVX1   g2739(.A(n3792), .Y(n3793));
  NAND3X1 g2740(.A(n3793), .B(n3791), .C(n3760), .Y(n3794));
  INVX1   g2741(.A(n3794), .Y(n3795));
  NOR2X1  g2742(.A(n3795), .B(n3764), .Y(n3796));
  NOR2X1  g2743(.A(n2560), .B(P1_REG2_REG_11__SCAN_IN), .Y(n3797));
  NOR3X1  g2744(.A(n3797), .B(n3796), .C(n3752), .Y(n3798));
  AOI21X1 g2745(.A0(n3755), .A1(n3746), .B0(n3798), .Y(n3799));
  AOI21X1 g2746(.A0(n2690), .A1(n3594), .B0(n3799), .Y(n3800));
  AOI21X1 g2747(.A0(n2691), .A1(P1_REG2_REG_14__SCAN_IN), .B0(n3800), .Y(n3801));
  NOR2X1  g2748(.A(n3801), .B(n3744), .Y(n3802));
  AOI21X1 g2749(.A0(n2735), .A1(P1_REG2_REG_15__SCAN_IN), .B0(n3802), .Y(n3803));
  INVX1   g2750(.A(n3803), .Y(n3804));
  NOR2X1  g2751(.A(n2776), .B(n3741), .Y(n3805));
  INVX1   g2752(.A(n3805), .Y(n3806));
  AOI21X1 g2753(.A0(n3806), .A1(n3742), .B0(n2821), .Y(n3807));
  AOI21X1 g2754(.A0(n3805), .A1(P1_REG2_REG_17__SCAN_IN), .B0(n3807), .Y(n3808));
  INVX1   g2755(.A(n3808), .Y(n3809));
  AOI21X1 g2756(.A0(n3804), .A1(n3743), .B0(n3809), .Y(n3810));
  OAI21X1 g2757(.A0(n2877), .A1(n3740), .B0(n3810), .Y(n3811));
  XOR2X1  g2758(.A(n1993), .B(P1_REG2_REG_19__SCAN_IN), .Y(n3812));
  AOI21X1 g2759(.A0(n2877), .A1(n3740), .B0(n3812), .Y(n3813));
  NAND2X1 g2760(.A(n3813), .B(n3811), .Y(n3814));
  AOI21X1 g2761(.A0(n2877), .A1(n3740), .B0(n3810), .Y(n3815));
  OAI21X1 g2762(.A0(n2877), .A1(n3740), .B0(n3812), .Y(n3816));
  OAI21X1 g2763(.A0(n3816), .A1(n3815), .B0(n3814), .Y(n3817));
  NOR4X1  g2764(.A(n2044), .B(n2042), .C(n2028), .D(n3488), .Y(n3818));
  NOR2X1  g2765(.A(n1994), .B(n1984), .Y(n3819));
  NOR4X1  g2766(.A(n3819), .B(n2045), .C(n2038), .D(n3469), .Y(n3820));
  NAND2X1 g2767(.A(n1991), .B(n1987), .Y(n3821));
  NAND4X1 g2768(.A(n3820), .B(n3818), .C(n3484), .D(n3821), .Y(n3822));
  INVX1   g2769(.A(n3822), .Y(n3823));
  INVX1   g2770(.A(n2002), .Y(n3824));
  NOR2X1  g2771(.A(n2092), .B(n3824), .Y(n3825));
  INVX1   g2772(.A(n3825), .Y(n3826));
  INVX1   g2773(.A(P1_REG1_REG_16__SCAN_IN), .Y(n3829));
  INVX1   g2774(.A(P1_REG1_REG_17__SCAN_IN), .Y(n3830));
  AOI22X1 g2775(.A0(n2776), .A1(n3829), .B0(n3830), .B1(n2821), .Y(n3831));
  NOR2X1  g2776(.A(n2691), .B(P1_REG1_REG_14__SCAN_IN), .Y(n3832));
  NOR2X1  g2777(.A(n2647), .B(P1_REG1_REG_13__SCAN_IN), .Y(n3833));
  INVX1   g2778(.A(P1_REG1_REG_11__SCAN_IN), .Y(n3834));
  NOR2X1  g2779(.A(n2559), .B(n3834), .Y(n3835));
  INVX1   g2780(.A(P1_REG1_REG_12__SCAN_IN), .Y(n3836));
  INVX1   g2781(.A(P1_REG1_REG_13__SCAN_IN), .Y(n3837));
  AOI22X1 g2782(.A0(n2604), .A1(n3836), .B0(n3837), .B1(n2646), .Y(n3838));
  NAND2X1 g2783(.A(n3838), .B(n3835), .Y(n3839));
  NOR2X1  g2784(.A(n2604), .B(n3836), .Y(n3840));
  AOI21X1 g2785(.A0(n2647), .A1(P1_REG1_REG_13__SCAN_IN), .B0(n3840), .Y(n3841));
  AOI21X1 g2786(.A0(n3841), .A1(n3839), .B0(n3833), .Y(n3842));
  NOR2X1  g2787(.A(n2605), .B(P1_REG1_REG_12__SCAN_IN), .Y(n3843));
  INVX1   g2788(.A(P1_REG1_REG_10__SCAN_IN), .Y(n3844));
  NAND2X1 g2789(.A(n2508), .B(n3844), .Y(n3845));
  INVX1   g2790(.A(P1_REG1_REG_8__SCAN_IN), .Y(n3846));
  NOR2X1  g2791(.A(n2422), .B(n3846), .Y(n3847));
  INVX1   g2792(.A(P1_REG1_REG_9__SCAN_IN), .Y(n3848));
  AOI22X1 g2793(.A0(n2466), .A1(n3848), .B0(n3844), .B1(n2508), .Y(n3849));
  NAND2X1 g2794(.A(n3849), .B(n3847), .Y(n3850));
  AOI22X1 g2795(.A0(n2467), .A1(P1_REG1_REG_9__SCAN_IN), .B0(P1_REG1_REG_10__SCAN_IN), .B1(n2509), .Y(n3851));
  NAND2X1 g2796(.A(n3851), .B(n3850), .Y(n3852));
  INVX1   g2797(.A(P1_REG1_REG_7__SCAN_IN), .Y(n3853));
  AOI22X1 g2798(.A0(n2329), .A1(n2311), .B0(n3853), .B1(n2376), .Y(n3854));
  INVX1   g2799(.A(n3854), .Y(n3855));
  INVX1   g2800(.A(P1_REG1_REG_5__SCAN_IN), .Y(n3856));
  AOI22X1 g2801(.A0(n2219), .A1(n2203), .B0(n3856), .B1(n2276), .Y(n3857));
  INVX1   g2802(.A(P1_REG1_REG_2__SCAN_IN), .Y(n3858));
  AOI22X1 g2803(.A0(n2119), .A1(n3858), .B0(n2150), .B1(n2169), .Y(n3859));
  INVX1   g2804(.A(P1_REG1_REG_1__SCAN_IN), .Y(n3860));
  NAND2X1 g2805(.A(n2008), .B(P1_REG1_REG_0__SCAN_IN), .Y(n3861));
  AOI21X1 g2806(.A0(n2078), .A1(n3860), .B0(n3861), .Y(n3862));
  NOR2X1  g2807(.A(n2078), .B(n3860), .Y(n3863));
  OAI21X1 g2808(.A0(n3863), .A1(n3862), .B0(n3859), .Y(n3864));
  NOR2X1  g2809(.A(n2169), .B(n2150), .Y(n3865));
  INVX1   g2810(.A(n3865), .Y(n3866));
  NOR2X1  g2811(.A(n2119), .B(n3858), .Y(n3867));
  OAI21X1 g2812(.A0(n2170), .A1(P1_REG1_REG_3__SCAN_IN), .B0(n3867), .Y(n3868));
  NAND3X1 g2813(.A(n3868), .B(n3866), .C(n3864), .Y(n3869));
  NAND2X1 g2814(.A(n3869), .B(n3857), .Y(n3870));
  NOR2X1  g2815(.A(n2219), .B(n2203), .Y(n3871));
  INVX1   g2816(.A(n3871), .Y(n3872));
  AOI21X1 g2817(.A0(n3872), .A1(n3856), .B0(n2276), .Y(n3873));
  AOI21X1 g2818(.A0(n3871), .A1(P1_REG1_REG_5__SCAN_IN), .B0(n3873), .Y(n3874));
  NAND2X1 g2819(.A(n3874), .B(n3870), .Y(n3875));
  INVX1   g2820(.A(n3875), .Y(n3876));
  NOR3X1  g2821(.A(n2329), .B(n3853), .C(n2311), .Y(n3877));
  OAI21X1 g2822(.A0(n2329), .A1(n2311), .B0(n3853), .Y(n3878));
  AOI21X1 g2823(.A0(n3878), .A1(n2377), .B0(n3877), .Y(n3879));
  OAI21X1 g2824(.A0(n3876), .A1(n3855), .B0(n3879), .Y(n3880));
  INVX1   g2825(.A(n3849), .Y(n3881));
  NOR2X1  g2826(.A(n2423), .B(P1_REG1_REG_8__SCAN_IN), .Y(n3882));
  NOR2X1  g2827(.A(n3882), .B(n3881), .Y(n3883));
  AOI22X1 g2828(.A0(n3880), .A1(n3883), .B0(n3852), .B1(n3845), .Y(n3884));
  NOR2X1  g2829(.A(n2560), .B(P1_REG1_REG_11__SCAN_IN), .Y(n3885));
  NOR4X1  g2830(.A(n3884), .B(n3843), .C(n3833), .D(n3885), .Y(n3886));
  NOR2X1  g2831(.A(n3886), .B(n3842), .Y(n3887));
  NOR2X1  g2832(.A(n3887), .B(n3832), .Y(n3888));
  AOI21X1 g2833(.A0(n2691), .A1(P1_REG1_REG_14__SCAN_IN), .B0(n3888), .Y(n3889));
  AOI21X1 g2834(.A0(n2734), .A1(n2723), .B0(n3889), .Y(n3890));
  AOI21X1 g2835(.A0(n2735), .A1(P1_REG1_REG_15__SCAN_IN), .B0(n3890), .Y(n3891));
  INVX1   g2836(.A(n3891), .Y(n3892));
  NOR2X1  g2837(.A(n2776), .B(n3829), .Y(n3893));
  INVX1   g2838(.A(n3893), .Y(n3894));
  AOI21X1 g2839(.A0(n3894), .A1(n3830), .B0(n2821), .Y(n3895));
  AOI21X1 g2840(.A0(n3893), .A1(P1_REG1_REG_17__SCAN_IN), .B0(n3895), .Y(n3896));
  INVX1   g2841(.A(n3896), .Y(n3897));
  AOI21X1 g2842(.A0(n3892), .A1(n3831), .B0(n3897), .Y(n3898));
  INVX1   g2843(.A(n3898), .Y(n3899));
  INVX1   g2844(.A(P1_REG1_REG_18__SCAN_IN), .Y(n3900));
  NOR2X1  g2845(.A(n2877), .B(n3900), .Y(n3901));
  XOR2X1  g2846(.A(n1993), .B(P1_REG1_REG_19__SCAN_IN), .Y(n3902));
  AOI21X1 g2847(.A0(n2877), .A1(n3900), .B0(n3902), .Y(n3903));
  OAI21X1 g2848(.A0(n3901), .A1(n3899), .B0(n3903), .Y(n3904));
  AOI21X1 g2849(.A0(n2877), .A1(n3900), .B0(n3898), .Y(n3905));
  OAI21X1 g2850(.A0(n2877), .A1(n3900), .B0(n3902), .Y(n3906));
  OAI21X1 g2851(.A0(n3906), .A1(n3905), .B0(n3904), .Y(n3907));
  INVX1   g2852(.A(n3907), .Y(n3908));
  INVX1   g2853(.A(n2092), .Y(n3910));
  AOI22X1 g2854(.A0(n3824), .A1(n3908), .B0(n2041), .B1(n2092), .Y(n3912));
  OAI21X1 g2855(.A0(n3826), .A1(n3817), .B0(n3912), .Y(n3913));
  NAND2X1 g2856(.A(n3913), .B(n3739), .Y(n3914));
  NAND3X1 g2857(.A(n1886), .B(n1880), .C(n1877), .Y(n3915));
  NOR2X1  g2858(.A(n3915), .B(n1875), .Y(n3916));
  NAND2X1 g2859(.A(n3738), .B(P1_STATE_REG_SCAN_IN), .Y(P1_U3083));
  NOR2X1  g2860(.A(P1_U3083), .B(n3916), .Y(n3918));
  NOR4X1  g2861(.A(n2002), .B(n1874), .C(P1_U3084), .D(n3918), .Y(n3919));
  NOR4X1  g2862(.A(n3918), .B(n1874), .C(P1_U3084), .D(n3826), .Y(n3920));
  INVX1   g2863(.A(n3920), .Y(n3921));
  NOR4X1  g2864(.A(n3910), .B(n1874), .C(P1_U3084), .D(n3918), .Y(n3922));
  INVX1   g2865(.A(n3918), .Y(n3923));
  OAI22X1 g2866(.A0(P1_STATE_REG_SCAN_IN), .A1(n2942), .B0(n1090), .B1(n3923), .Y(n3924));
  AOI21X1 g2867(.A0(n3922), .A1(n2041), .B0(n3924), .Y(n3925));
  OAI21X1 g2868(.A0(n3921), .A1(n3817), .B0(n3925), .Y(n3926));
  AOI21X1 g2869(.A0(n3919), .A1(n3908), .B0(n3926), .Y(n3927));
  NAND2X1 g2870(.A(n3927), .B(n3914), .Y(P1_U3260));
  XOR2X1  g2871(.A(n2877), .B(P1_REG2_REG_18__SCAN_IN), .Y(n3929));
  INVX1   g2872(.A(n3929), .Y(n3930));
  XOR2X1  g2873(.A(n3930), .B(n3810), .Y(n3931));
  NOR2X1  g2874(.A(n3931), .B(n3826), .Y(n3932));
  XOR2X1  g2875(.A(n2877), .B(n3900), .Y(n3935));
  XOR2X1  g2876(.A(n3935), .B(n3898), .Y(n3936));
  OAI22X1 g2877(.A0(n3910), .A1(n2877), .B0(n2002), .B1(n3936), .Y(n3937));
  OAI21X1 g2878(.A0(n3937), .A1(n3932), .B0(n3739), .Y(n3938));
  INVX1   g2879(.A(n3919), .Y(n3939));
  NOR2X1  g2880(.A(n3936), .B(n3939), .Y(n3940));
  NOR2X1  g2881(.A(n3931), .B(n3921), .Y(n3941));
  INVX1   g2882(.A(n3922), .Y(n3942));
  AOI22X1 g2883(.A0(P1_U3084), .A1(P1_REG3_REG_18__SCAN_IN), .B0(P1_ADDR_REG_18__SCAN_IN), .B1(n3918), .Y(n3943));
  OAI21X1 g2884(.A0(n3942), .A1(n2877), .B0(n3943), .Y(n3944));
  NOR3X1  g2885(.A(n3944), .B(n3941), .C(n3940), .Y(n3945));
  NAND2X1 g2886(.A(n3945), .B(n3938), .Y(P1_U3259));
  INVX1   g2887(.A(n3739), .Y(n3947));
  OAI21X1 g2888(.A0(n2821), .A1(n3742), .B0(n3743), .Y(n3948));
  AOI21X1 g2889(.A0(n3806), .A1(n3803), .B0(n3948), .Y(n3949));
  NOR2X1  g2890(.A(n2777), .B(P1_REG2_REG_16__SCAN_IN), .Y(n3950));
  INVX1   g2891(.A(n3950), .Y(n3951));
  XOR2X1  g2892(.A(n2821), .B(P1_REG2_REG_17__SCAN_IN), .Y(n3952));
  OAI21X1 g2893(.A0(n2776), .A1(n3741), .B0(n3952), .Y(n3953));
  AOI21X1 g2894(.A0(n3804), .A1(n3951), .B0(n3953), .Y(n3954));
  NOR3X1  g2895(.A(n3954), .B(n3949), .C(n3826), .Y(n3955));
  OAI21X1 g2896(.A0(n2821), .A1(n3830), .B0(n3831), .Y(n3956));
  AOI21X1 g2897(.A0(n3894), .A1(n3891), .B0(n3956), .Y(n3957));
  AOI21X1 g2898(.A0(n2776), .A1(n3829), .B0(n3891), .Y(n3958));
  XOR2X1  g2899(.A(n2821), .B(n3830), .Y(n3959));
  NOR3X1  g2900(.A(n3959), .B(n3958), .C(n3893), .Y(n3960));
  NOR3X1  g2901(.A(n3960), .B(n3957), .C(n2002), .Y(n3961));
  NOR3X1  g2902(.A(n3823), .B(n2821), .C(n3910), .Y(n3962));
  NOR3X1  g2903(.A(n3962), .B(n3961), .C(n3955), .Y(n3963));
  NOR3X1  g2904(.A(n3960), .B(n3957), .C(n3939), .Y(n3964));
  NOR3X1  g2905(.A(n3954), .B(n3949), .C(n3921), .Y(n3965));
  AOI22X1 g2906(.A0(P1_U3084), .A1(P1_REG3_REG_17__SCAN_IN), .B0(P1_ADDR_REG_17__SCAN_IN), .B1(n3918), .Y(n3966));
  OAI21X1 g2907(.A0(n3942), .A1(n2821), .B0(n3966), .Y(n3967));
  NOR3X1  g2908(.A(n3967), .B(n3965), .C(n3964), .Y(n3968));
  OAI21X1 g2909(.A0(n3963), .A1(n3947), .B0(n3968), .Y(P1_U3258));
  XOR2X1  g2910(.A(n2776), .B(n3741), .Y(n3970));
  AOI21X1 g2911(.A0(n3806), .A1(n3951), .B0(n3803), .Y(n3971));
  AOI21X1 g2912(.A0(n3970), .A1(n3803), .B0(n3971), .Y(n3972));
  NOR2X1  g2913(.A(n3972), .B(n3826), .Y(n3973));
  XOR2X1  g2914(.A(n2776), .B(n3829), .Y(n3974));
  NOR2X1  g2915(.A(n3974), .B(n3891), .Y(n3976));
  AOI21X1 g2916(.A0(n3974), .A1(n3891), .B0(n3976), .Y(n3977));
  OAI22X1 g2917(.A0(n3910), .A1(n2776), .B0(n2002), .B1(n3977), .Y(n3978));
  OAI21X1 g2918(.A0(n3978), .A1(n3973), .B0(n3739), .Y(n3979));
  NOR2X1  g2919(.A(n3977), .B(n3939), .Y(n3980));
  NOR2X1  g2920(.A(n3972), .B(n3921), .Y(n3981));
  AOI22X1 g2921(.A0(P1_U3084), .A1(P1_REG3_REG_16__SCAN_IN), .B0(P1_ADDR_REG_16__SCAN_IN), .B1(n3918), .Y(n3982));
  OAI21X1 g2922(.A0(n3942), .A1(n2776), .B0(n3982), .Y(n3983));
  NOR3X1  g2923(.A(n3983), .B(n3981), .C(n3980), .Y(n3984));
  NAND2X1 g2924(.A(n3984), .B(n3979), .Y(P1_U3257));
  XOR2X1  g2925(.A(n2734), .B(P1_REG2_REG_15__SCAN_IN), .Y(n3986));
  XOR2X1  g2926(.A(n3986), .B(n3801), .Y(n3987));
  XOR2X1  g2927(.A(n2734), .B(n2723), .Y(n3988));
  XOR2X1  g2928(.A(n3988), .B(n3889), .Y(n3989));
  OAI22X1 g2929(.A0(n3910), .A1(n2734), .B0(n2002), .B1(n3989), .Y(n3990));
  AOI21X1 g2930(.A0(n3987), .A1(n3825), .B0(n3990), .Y(n3991));
  NOR2X1  g2931(.A(n3989), .B(n3939), .Y(n3992));
  NAND2X1 g2932(.A(n3987), .B(n3920), .Y(n3993));
  NAND2X1 g2933(.A(n3922), .B(n2735), .Y(n3994));
  AOI22X1 g2934(.A0(P1_U3084), .A1(P1_REG3_REG_15__SCAN_IN), .B0(P1_ADDR_REG_15__SCAN_IN), .B1(n3918), .Y(n3995));
  NAND3X1 g2935(.A(n3995), .B(n3994), .C(n3993), .Y(n3996));
  NOR2X1  g2936(.A(n3996), .B(n3992), .Y(n3997));
  OAI21X1 g2937(.A0(n3991), .A1(n3947), .B0(n3997), .Y(P1_U3256));
  XOR2X1  g2938(.A(n2690), .B(P1_REG2_REG_14__SCAN_IN), .Y(n3999));
  XOR2X1  g2939(.A(n3999), .B(n3799), .Y(n4000));
  NAND2X1 g2940(.A(n4000), .B(n3825), .Y(n4001));
  XOR2X1  g2941(.A(n2690), .B(P1_REG1_REG_14__SCAN_IN), .Y(n4002));
  XOR2X1  g2942(.A(n4002), .B(n3887), .Y(n4003));
  AOI22X1 g2943(.A0(n2092), .A1(n2691), .B0(n3824), .B1(n4003), .Y(n4004));
  NAND2X1 g2944(.A(n4004), .B(n4001), .Y(n4005));
  NAND2X1 g2945(.A(n4005), .B(n3739), .Y(n4006));
  NAND2X1 g2946(.A(n4000), .B(n3920), .Y(n4007));
  AOI22X1 g2947(.A0(P1_U3084), .A1(P1_REG3_REG_14__SCAN_IN), .B0(P1_ADDR_REG_14__SCAN_IN), .B1(n3918), .Y(n4008));
  AOI22X1 g2948(.A0(n3922), .A1(n2691), .B0(n3919), .B1(n4003), .Y(n4009));
  NAND4X1 g2949(.A(n4008), .B(n4007), .C(n4006), .D(n4009), .Y(P1_U3255));
  INVX1   g2950(.A(n3753), .Y(n4011));
  INVX1   g2951(.A(n3796), .Y(n4012));
  INVX1   g2952(.A(n3797), .Y(n4013));
  AOI21X1 g2953(.A0(n4013), .A1(n4012), .B0(n3748), .Y(n4014));
  OAI21X1 g2954(.A0(n2646), .A1(n3745), .B0(n3751), .Y(n4015));
  AOI21X1 g2955(.A0(n4014), .A1(n4011), .B0(n4015), .Y(n4016));
  NOR2X1  g2956(.A(n2605), .B(P1_REG2_REG_12__SCAN_IN), .Y(n4017));
  NOR2X1  g2957(.A(n4014), .B(n4017), .Y(n4018));
  XOR2X1  g2958(.A(n2646), .B(n3745), .Y(n4019));
  NOR3X1  g2959(.A(n4019), .B(n4018), .C(n3753), .Y(n4020));
  NOR3X1  g2960(.A(n4020), .B(n4016), .C(n3826), .Y(n4021));
  INVX1   g2961(.A(n3884), .Y(n4022));
  INVX1   g2962(.A(n3885), .Y(n4023));
  AOI21X1 g2963(.A0(n4023), .A1(n4022), .B0(n3835), .Y(n4024));
  INVX1   g2964(.A(n4024), .Y(n4025));
  NOR2X1  g2965(.A(n4025), .B(n3840), .Y(n4026));
  OAI21X1 g2966(.A0(n2646), .A1(n3837), .B0(n3838), .Y(n4027));
  XOR2X1  g2967(.A(n2646), .B(n3837), .Y(n4028));
  NOR2X1  g2968(.A(n4028), .B(n3840), .Y(n4029));
  OAI21X1 g2969(.A0(n4024), .A1(n3843), .B0(n4029), .Y(n4030));
  OAI21X1 g2970(.A0(n4027), .A1(n4026), .B0(n4030), .Y(n4031));
  OAI22X1 g2971(.A0(n3910), .A1(n2646), .B0(n2002), .B1(n4031), .Y(n4032));
  OAI21X1 g2972(.A0(n4032), .A1(n4021), .B0(n3739), .Y(n4033));
  NOR2X1  g2973(.A(n4031), .B(n3939), .Y(n4034));
  NOR3X1  g2974(.A(n4020), .B(n4016), .C(n3921), .Y(n4035));
  AOI22X1 g2975(.A0(P1_U3084), .A1(P1_REG3_REG_13__SCAN_IN), .B0(P1_ADDR_REG_13__SCAN_IN), .B1(n3918), .Y(n4036));
  OAI21X1 g2976(.A0(n3942), .A1(n2646), .B0(n4036), .Y(n4037));
  NOR3X1  g2977(.A(n4037), .B(n4035), .C(n4034), .Y(n4038));
  NAND2X1 g2978(.A(n4038), .B(n4033), .Y(P1_U3254));
  XOR2X1  g2979(.A(n2604), .B(n3750), .Y(n4042));
  NOR2X1  g2980(.A(n4042), .B(n4014), .Y(n4043));
  AOI21X1 g2981(.A0(n4042), .A1(n4014), .B0(n4043), .Y(n4044));
  NOR2X1  g2982(.A(n4044), .B(n3826), .Y(n4045));
  XOR2X1  g2983(.A(n2604), .B(n3836), .Y(n4046));
  NOR2X1  g2984(.A(n4046), .B(n4024), .Y(n4048));
  AOI21X1 g2985(.A0(n4046), .A1(n4024), .B0(n4048), .Y(n4049));
  OAI22X1 g2986(.A0(n3910), .A1(n2604), .B0(n2002), .B1(n4049), .Y(n4050));
  OAI21X1 g2987(.A0(n4050), .A1(n4045), .B0(n3739), .Y(n4051));
  AOI22X1 g2988(.A0(P1_U3084), .A1(P1_REG3_REG_12__SCAN_IN), .B0(P1_ADDR_REG_12__SCAN_IN), .B1(n3918), .Y(n4052));
  OAI21X1 g2989(.A0(n4044), .A1(n3921), .B0(n4052), .Y(n4053));
  OAI22X1 g2990(.A0(n3942), .A1(n2604), .B0(n3939), .B1(n4049), .Y(n4054));
  NOR2X1  g2991(.A(n4054), .B(n4053), .Y(n4055));
  NAND2X1 g2992(.A(n4055), .B(n4051), .Y(P1_U3253));
  XOR2X1  g2993(.A(n2559), .B(n3747), .Y(n4057));
  AOI21X1 g2994(.A0(n4013), .A1(n3749), .B0(n3796), .Y(n4058));
  AOI21X1 g2995(.A0(n4057), .A1(n3796), .B0(n4058), .Y(n4059));
  NOR2X1  g2996(.A(n4059), .B(n3826), .Y(n4060));
  XOR2X1  g2997(.A(n2559), .B(n3834), .Y(n4061));
  NOR2X1  g2998(.A(n4061), .B(n3884), .Y(n4063));
  AOI21X1 g2999(.A0(n4061), .A1(n3884), .B0(n4063), .Y(n4064));
  OAI22X1 g3000(.A0(n3910), .A1(n2559), .B0(n2002), .B1(n4064), .Y(n4065));
  OAI21X1 g3001(.A0(n4065), .A1(n4060), .B0(n3739), .Y(n4066));
  AOI22X1 g3002(.A0(P1_U3084), .A1(P1_REG3_REG_11__SCAN_IN), .B0(P1_ADDR_REG_11__SCAN_IN), .B1(n3918), .Y(n4067));
  OAI21X1 g3003(.A0(n4059), .A1(n3921), .B0(n4067), .Y(n4068));
  OAI22X1 g3004(.A0(n3942), .A1(n2559), .B0(n3939), .B1(n4064), .Y(n4069));
  NOR2X1  g3005(.A(n4069), .B(n4068), .Y(n4070));
  NAND2X1 g3006(.A(n4070), .B(n4066), .Y(P1_U3252));
  AOI21X1 g3007(.A0(n3793), .A1(n3791), .B0(n3758), .Y(n4072));
  OAI21X1 g3008(.A0(n2508), .A1(n3756), .B0(n3760), .Y(n4073));
  AOI21X1 g3009(.A0(n4072), .A1(n3761), .B0(n4073), .Y(n4074));
  AOI21X1 g3010(.A0(n2466), .A1(n3759), .B0(n4072), .Y(n4075));
  AOI22X1 g3011(.A0(n2467), .A1(P1_REG2_REG_9__SCAN_IN), .B0(n3756), .B1(n2509), .Y(n4076));
  OAI21X1 g3012(.A0(n2509), .A1(n3756), .B0(n4076), .Y(n4077));
  NOR2X1  g3013(.A(n4077), .B(n4075), .Y(n4078));
  NOR3X1  g3014(.A(n4078), .B(n4074), .C(n3826), .Y(n4079));
  NAND2X1 g3015(.A(n2467), .B(P1_REG1_REG_9__SCAN_IN), .Y(n4080));
  INVX1   g3016(.A(n3882), .Y(n4081));
  AOI21X1 g3017(.A0(n4081), .A1(n3880), .B0(n3847), .Y(n4082));
  OAI21X1 g3018(.A0(n2508), .A1(n3844), .B0(n3849), .Y(n4083));
  AOI21X1 g3019(.A0(n4082), .A1(n4080), .B0(n4083), .Y(n4084));
  AOI21X1 g3020(.A0(n2466), .A1(n3848), .B0(n4082), .Y(n4085));
  AOI22X1 g3021(.A0(n2467), .A1(P1_REG1_REG_9__SCAN_IN), .B0(n3844), .B1(n2509), .Y(n4086));
  OAI21X1 g3022(.A0(n2509), .A1(n3844), .B0(n4086), .Y(n4087));
  NOR2X1  g3023(.A(n4087), .B(n4085), .Y(n4088));
  NOR3X1  g3024(.A(n4088), .B(n4084), .C(n2002), .Y(n4089));
  NOR3X1  g3025(.A(n3823), .B(n2508), .C(n3910), .Y(n4090));
  NOR3X1  g3026(.A(n4090), .B(n4089), .C(n4079), .Y(n4091));
  NOR3X1  g3027(.A(n4078), .B(n4074), .C(n3921), .Y(n4092));
  NAND2X1 g3028(.A(n3918), .B(P1_ADDR_REG_10__SCAN_IN), .Y(n4093));
  OAI21X1 g3029(.A0(P1_STATE_REG_SCAN_IN), .A1(n2492), .B0(n4093), .Y(n4094));
  NOR3X1  g3030(.A(n4088), .B(n4084), .C(n3939), .Y(n4095));
  NOR2X1  g3031(.A(n3942), .B(n2508), .Y(n4096));
  NOR4X1  g3032(.A(n4095), .B(n4094), .C(n4092), .D(n4096), .Y(n4097));
  OAI21X1 g3033(.A0(n4091), .A1(n3947), .B0(n4097), .Y(P1_U3251));
  XOR2X1  g3034(.A(n2466), .B(n3759), .Y(n4099));
  NOR2X1  g3035(.A(n4099), .B(n4072), .Y(n4101));
  AOI21X1 g3036(.A0(n4099), .A1(n4072), .B0(n4101), .Y(n4102));
  NOR2X1  g3037(.A(n4102), .B(n3826), .Y(n4103));
  XOR2X1  g3038(.A(n2466), .B(n3848), .Y(n4104));
  NOR2X1  g3039(.A(n4104), .B(n4082), .Y(n4106));
  AOI21X1 g3040(.A0(n4104), .A1(n4082), .B0(n4106), .Y(n4107));
  OAI22X1 g3041(.A0(n3910), .A1(n2466), .B0(n2002), .B1(n4107), .Y(n4108));
  OAI21X1 g3042(.A0(n4108), .A1(n4103), .B0(n3739), .Y(n4109));
  AOI22X1 g3043(.A0(P1_U3084), .A1(P1_REG3_REG_9__SCAN_IN), .B0(P1_ADDR_REG_9__SCAN_IN), .B1(n3918), .Y(n4110));
  OAI21X1 g3044(.A0(n4102), .A1(n3921), .B0(n4110), .Y(n4111));
  OAI22X1 g3045(.A0(n3942), .A1(n2466), .B0(n3939), .B1(n4107), .Y(n4112));
  NOR2X1  g3046(.A(n4112), .B(n4111), .Y(n4113));
  NAND2X1 g3047(.A(n4113), .B(n4109), .Y(P1_U3250));
  NOR3X1  g3048(.A(n3823), .B(n2422), .C(n3910), .Y(n4115));
  XOR2X1  g3049(.A(n2422), .B(P1_REG1_REG_8__SCAN_IN), .Y(n4116));
  NOR2X1  g3050(.A(n4116), .B(n3880), .Y(n4117));
  AOI21X1 g3051(.A0(n4116), .A1(n3880), .B0(n4117), .Y(n4119));
  XOR2X1  g3052(.A(n2422), .B(P1_REG2_REG_8__SCAN_IN), .Y(n4120));
  NOR2X1  g3053(.A(n4120), .B(n3791), .Y(n4121));
  AOI21X1 g3054(.A0(n4120), .A1(n3791), .B0(n4121), .Y(n4123));
  OAI22X1 g3055(.A0(n4119), .A1(n2002), .B0(n3826), .B1(n4123), .Y(n4124));
  OAI21X1 g3056(.A0(n4124), .A1(n4115), .B0(n3739), .Y(n4125));
  AOI22X1 g3057(.A0(P1_U3084), .A1(P1_REG3_REG_8__SCAN_IN), .B0(P1_ADDR_REG_8__SCAN_IN), .B1(n3918), .Y(n4126));
  NOR2X1  g3058(.A(n4123), .B(n3921), .Y(n4127));
  OAI22X1 g3059(.A0(n3942), .A1(n2422), .B0(n3939), .B1(n4119), .Y(n4128));
  NOR2X1  g3060(.A(n4128), .B(n4127), .Y(n4129));
  NAND3X1 g3061(.A(n4129), .B(n4126), .C(n4125), .Y(P1_U3249));
  NOR2X1  g3062(.A(n2329), .B(n2311), .Y(n4131));
  AOI21X1 g3063(.A0(n2377), .A1(P1_REG1_REG_7__SCAN_IN), .B0(n3855), .Y(n4132));
  OAI21X1 g3064(.A0(n4131), .A1(n3875), .B0(n4132), .Y(n4133));
  AOI22X1 g3065(.A0(n3870), .A1(n3874), .B0(n2329), .B1(n2311), .Y(n4134));
  AOI21X1 g3066(.A0(n2377), .A1(n3853), .B0(n4131), .Y(n4135));
  OAI21X1 g3067(.A0(n2377), .A1(n3853), .B0(n4135), .Y(n4136));
  OAI21X1 g3068(.A0(n4136), .A1(n4134), .B0(n4133), .Y(n4137));
  INVX1   g3069(.A(n4137), .Y(n4138));
  NAND3X1 g3070(.A(n3788), .B(n3783), .C(n3779), .Y(n4139));
  AOI21X1 g3071(.A0(n2377), .A1(P1_REG2_REG_7__SCAN_IN), .B0(n3765), .Y(n4140));
  AOI22X1 g3072(.A0(n3779), .A1(n3783), .B0(n2329), .B1(n2335), .Y(n4141));
  AOI21X1 g3073(.A0(n2377), .A1(n3787), .B0(n3786), .Y(n4142));
  OAI21X1 g3074(.A0(n2377), .A1(n3787), .B0(n4142), .Y(n4143));
  NOR2X1  g3075(.A(n4143), .B(n4141), .Y(n4144));
  AOI21X1 g3076(.A0(n4140), .A1(n4139), .B0(n4144), .Y(n4145));
  AOI22X1 g3077(.A0(n4138), .A1(n3824), .B0(n3825), .B1(n4145), .Y(n4146));
  OAI21X1 g3078(.A0(n3910), .A1(n2376), .B0(n4146), .Y(n4147));
  OAI22X1 g3079(.A0(P1_STATE_REG_SCAN_IN), .A1(n2405), .B0(n1047), .B1(n3923), .Y(n4148));
  AOI21X1 g3080(.A0(n4147), .A1(n3739), .B0(n4148), .Y(n4149));
  NAND2X1 g3081(.A(n4145), .B(n3920), .Y(n4150));
  AOI22X1 g3082(.A0(n3922), .A1(n2377), .B0(n3919), .B1(n4138), .Y(n4151));
  NAND3X1 g3083(.A(n4151), .B(n4150), .C(n4149), .Y(P1_U3248));
  XOR2X1  g3084(.A(n2329), .B(n2335), .Y(n4153));
  NAND3X1 g3085(.A(n4153), .B(n3783), .C(n3779), .Y(n4154));
  OAI21X1 g3086(.A0(n4153), .A1(n3785), .B0(n4154), .Y(n4156));
  NAND2X1 g3087(.A(n4156), .B(n3920), .Y(n4157));
  AOI22X1 g3088(.A0(P1_U3084), .A1(P1_REG3_REG_6__SCAN_IN), .B0(P1_ADDR_REG_6__SCAN_IN), .B1(n3918), .Y(n4158));
  XOR2X1  g3089(.A(n2329), .B(n2311), .Y(n4159));
  NAND3X1 g3090(.A(n4159), .B(n3874), .C(n3870), .Y(n4160));
  OAI21X1 g3091(.A0(n4159), .A1(n3876), .B0(n4160), .Y(n4162));
  NAND2X1 g3092(.A(n4162), .B(n3919), .Y(n4163));
  AOI22X1 g3093(.A0(n4156), .A1(n3825), .B0(n3824), .B1(n4162), .Y(n4164));
  OAI21X1 g3094(.A0(n3910), .A1(n2329), .B0(n4164), .Y(n4165));
  AOI22X1 g3095(.A0(n3922), .A1(n2330), .B0(n3739), .B1(n4165), .Y(n4166));
  NAND4X1 g3096(.A(n4163), .B(n4158), .C(n4157), .D(n4166), .Y(P1_U3247));
  NOR2X1  g3097(.A(n2170), .B(P1_REG2_REG_3__SCAN_IN), .Y(n4168));
  NOR2X1  g3098(.A(n2120), .B(P1_REG2_REG_2__SCAN_IN), .Y(n4169));
  NOR3X1  g3099(.A(n3770), .B(n4169), .C(n4168), .Y(n4170));
  NOR3X1  g3100(.A(n4169), .B(n2078), .C(n2055), .Y(n4171));
  NOR2X1  g3101(.A(n4171), .B(n3776), .Y(n4172));
  OAI21X1 g3102(.A0(n4172), .A1(n4168), .B0(n3775), .Y(n4173));
  NOR2X1  g3103(.A(n4173), .B(n4170), .Y(n4174));
  OAI21X1 g3104(.A0(n2276), .A1(n2254), .B0(n3766), .Y(n4175));
  AOI21X1 g3105(.A0(n4174), .A1(n3781), .B0(n4175), .Y(n4176));
  OAI22X1 g3106(.A0(n4170), .A1(n4173), .B0(n2220), .B1(P1_REG2_REG_4__SCAN_IN), .Y(n4177));
  OAI22X1 g3107(.A0(n2219), .A1(n3515), .B0(P1_REG2_REG_5__SCAN_IN), .B1(n2276), .Y(n4178));
  AOI21X1 g3108(.A0(n2276), .A1(P1_REG2_REG_5__SCAN_IN), .B0(n4178), .Y(n4179));
  AOI21X1 g3109(.A0(n4179), .A1(n4177), .B0(n4176), .Y(n4180));
  NAND2X1 g3110(.A(n4180), .B(n3920), .Y(n4181));
  AOI22X1 g3111(.A0(P1_U3084), .A1(P1_REG3_REG_5__SCAN_IN), .B0(P1_ADDR_REG_5__SCAN_IN), .B1(n3918), .Y(n4182));
  NOR2X1  g3112(.A(n2170), .B(P1_REG1_REG_3__SCAN_IN), .Y(n4183));
  NOR2X1  g3113(.A(n2120), .B(P1_REG1_REG_2__SCAN_IN), .Y(n4184));
  INVX1   g3114(.A(n3862), .Y(n4185));
  NOR3X1  g3115(.A(n4185), .B(n4184), .C(n4183), .Y(n4186));
  NOR3X1  g3116(.A(n4184), .B(n2078), .C(n3860), .Y(n4187));
  NOR2X1  g3117(.A(n4187), .B(n3867), .Y(n4188));
  OAI21X1 g3118(.A0(n4188), .A1(n4183), .B0(n3866), .Y(n4189));
  NOR2X1  g3119(.A(n4189), .B(n4186), .Y(n4190));
  OAI21X1 g3120(.A0(n2276), .A1(n3856), .B0(n3857), .Y(n4191));
  AOI21X1 g3121(.A0(n4190), .A1(n3872), .B0(n4191), .Y(n4192));
  OAI22X1 g3122(.A0(n4186), .A1(n4189), .B0(n2220), .B1(P1_REG1_REG_4__SCAN_IN), .Y(n4193));
  OAI22X1 g3123(.A0(n2219), .A1(n2203), .B0(P1_REG1_REG_5__SCAN_IN), .B1(n2276), .Y(n4194));
  AOI21X1 g3124(.A0(n2276), .A1(P1_REG1_REG_5__SCAN_IN), .B0(n4194), .Y(n4195));
  AOI21X1 g3125(.A0(n4195), .A1(n4193), .B0(n4192), .Y(n4196));
  NAND2X1 g3126(.A(n4196), .B(n3919), .Y(n4197));
  INVX1   g3127(.A(n2276), .Y(n4198));
  AOI22X1 g3128(.A0(n4180), .A1(n3825), .B0(n3824), .B1(n4196), .Y(n4199));
  OAI21X1 g3129(.A0(n3910), .A1(n2276), .B0(n4199), .Y(n4200));
  AOI22X1 g3130(.A0(n3922), .A1(n4198), .B0(n3739), .B1(n4200), .Y(n4201));
  NAND4X1 g3131(.A(n4197), .B(n4182), .C(n4181), .D(n4201), .Y(P1_U3246));
  NOR3X1  g3132(.A(n3915), .B(n1875), .C(P1_U3084), .Y(P1_U4006));
  INVX1   g3133(.A(P1_U4006), .Y(n4204));
  NAND2X1 g3134(.A(n2041), .B(n1989), .Y(n4205));
  OAI21X1 g3135(.A0(n1989), .A1(n1987), .B0(n4205), .Y(n4206));
  OAI21X1 g3136(.A0(n4206), .A1(n2067), .B0(n3915), .Y(n4207));
  NOR3X1  g3137(.A(n3819), .B(n2065), .C(n2038), .Y(n4208));
  AOI21X1 g3138(.A0(n4208), .A1(n4205), .B0(n1884), .Y(n4209));
  INVX1   g3139(.A(n2008), .Y(n4210));
  NAND3X1 g3140(.A(n1991), .B(n1987), .C(n3915), .Y(n4211));
  OAI22X1 g3141(.A0(n2010), .A1(n4211), .B0(n4210), .B1(n3915), .Y(n4212));
  AOI21X1 g3142(.A0(n4209), .A1(n2025), .B0(n4212), .Y(n4213));
  XOR2X1  g3143(.A(n4213), .B(n4207), .Y(n4214));
  INVX1   g3144(.A(n4207), .Y(n4215));
  AOI21X1 g3145(.A0(n2067), .A1(n3915), .B0(n4209), .Y(n4216));
  INVX1   g3146(.A(n4211), .Y(n4217));
  AOI22X1 g3147(.A0(n2025), .A1(n4217), .B0(n1884), .B1(P1_REG1_REG_0__SCAN_IN), .Y(n4218));
  OAI21X1 g3148(.A0(n4216), .A1(n2010), .B0(n4218), .Y(n4219));
  XOR2X1  g3149(.A(n4219), .B(n4215), .Y(n4220));
  XOR2X1  g3150(.A(n4220), .B(n4214), .Y(n4221));
  NOR2X1  g3151(.A(n2092), .B(n2002), .Y(n4222));
  NAND3X1 g3152(.A(n3825), .B(n4210), .C(P1_REG2_REG_0__SCAN_IN), .Y(n4223));
  AOI21X1 g3153(.A0(n2002), .A1(n2018), .B0(n2092), .Y(n4224));
  OAI21X1 g3154(.A0(n4224), .A1(n4210), .B0(n4223), .Y(n4225));
  AOI21X1 g3155(.A0(n4222), .A1(n4221), .B0(n4225), .Y(n4226));
  XOR2X1  g3156(.A(n2219), .B(n3515), .Y(n4227));
  NOR2X1  g3157(.A(n4227), .B(n4174), .Y(n4229));
  AOI21X1 g3158(.A0(n4227), .A1(n4174), .B0(n4229), .Y(n4230));
  AOI22X1 g3159(.A0(P1_U3084), .A1(P1_REG3_REG_4__SCAN_IN), .B0(P1_ADDR_REG_4__SCAN_IN), .B1(n3918), .Y(n4231));
  OAI21X1 g3160(.A0(n4230), .A1(n3921), .B0(n4231), .Y(n4232));
  NOR2X1  g3161(.A(n3942), .B(n2219), .Y(n4233));
  XOR2X1  g3162(.A(n2219), .B(n2203), .Y(n4234));
  NOR2X1  g3163(.A(n4234), .B(n4190), .Y(n4236));
  AOI21X1 g3164(.A0(n4234), .A1(n4190), .B0(n4236), .Y(n4237));
  OAI22X1 g3165(.A0(n4230), .A1(n3826), .B0(n2002), .B1(n4237), .Y(n4238));
  AOI21X1 g3166(.A0(n2092), .A1(n2220), .B0(n4238), .Y(n4239));
  OAI22X1 g3167(.A0(n4237), .A1(n3939), .B0(n3947), .B1(n4239), .Y(n4240));
  NOR3X1  g3168(.A(n4240), .B(n4233), .C(n4232), .Y(n4241));
  OAI21X1 g3169(.A0(n4226), .A1(n4204), .B0(n4241), .Y(P1_U3245));
  OAI21X1 g3170(.A0(n3770), .A1(n4169), .B0(n4172), .Y(n4243));
  XOR2X1  g3171(.A(n2169), .B(P1_REG2_REG_3__SCAN_IN), .Y(n4244));
  OAI21X1 g3172(.A0(n3774), .A1(n4168), .B0(n4243), .Y(n4245));
  OAI21X1 g3173(.A0(n4244), .A1(n4243), .B0(n4245), .Y(n4246));
  OAI22X1 g3174(.A0(P1_STATE_REG_SCAN_IN), .A1(n3507), .B0(n1052), .B1(n3923), .Y(n4247));
  AOI21X1 g3175(.A0(n4246), .A1(n3920), .B0(n4247), .Y(n4248));
  OAI21X1 g3176(.A0(n4185), .A1(n4184), .B0(n4188), .Y(n4249));
  XOR2X1  g3177(.A(n2169), .B(P1_REG1_REG_3__SCAN_IN), .Y(n4250));
  OAI21X1 g3178(.A0(n3865), .A1(n4183), .B0(n4249), .Y(n4251));
  OAI21X1 g3179(.A0(n4250), .A1(n4249), .B0(n4251), .Y(n4252));
  NAND2X1 g3180(.A(n4252), .B(n3919), .Y(n4253));
  AOI22X1 g3181(.A0(n4246), .A1(n3825), .B0(n3824), .B1(n4252), .Y(n4254));
  OAI21X1 g3182(.A0(n3910), .A1(n2169), .B0(n4254), .Y(n4255));
  AOI22X1 g3183(.A0(n3922), .A1(n2170), .B0(n3739), .B1(n4255), .Y(n4256));
  NAND3X1 g3184(.A(n4256), .B(n4253), .C(n4248), .Y(P1_U3244));
  NOR2X1  g3185(.A(n3772), .B(n3771), .Y(n4258));
  NOR3X1  g3186(.A(n3776), .B(n4258), .C(n4169), .Y(n4259));
  XOR2X1  g3187(.A(n2119), .B(P1_REG2_REG_2__SCAN_IN), .Y(n4260));
  AOI21X1 g3188(.A0(n4260), .A1(n4258), .B0(n4259), .Y(n4261));
  NAND2X1 g3189(.A(n4261), .B(n3920), .Y(n4262));
  AOI22X1 g3190(.A0(P1_U3084), .A1(P1_REG3_REG_2__SCAN_IN), .B0(P1_ADDR_REG_2__SCAN_IN), .B1(n3918), .Y(n4263));
  NAND2X1 g3191(.A(n4263), .B(n4262), .Y(n4264));
  NOR2X1  g3192(.A(n3863), .B(n3862), .Y(n4265));
  NOR3X1  g3193(.A(n3867), .B(n4265), .C(n4184), .Y(n4266));
  XOR2X1  g3194(.A(n2119), .B(P1_REG1_REG_2__SCAN_IN), .Y(n4267));
  AOI21X1 g3195(.A0(n4267), .A1(n4265), .B0(n4266), .Y(n4268));
  NAND3X1 g3196(.A(n3822), .B(n2120), .C(n2092), .Y(n4269));
  AOI22X1 g3197(.A0(n4261), .A1(n3825), .B0(n3824), .B1(n4268), .Y(n4270));
  AOI21X1 g3198(.A0(n4270), .A1(n4269), .B0(n3947), .Y(n4271));
  AOI21X1 g3199(.A0(n4268), .A1(n3919), .B0(n4271), .Y(n4272));
  OAI21X1 g3200(.A0(n3942), .A1(n2119), .B0(n4272), .Y(n4273));
  NOR2X1  g3201(.A(n4273), .B(n4264), .Y(n4274));
  OAI21X1 g3202(.A0(n4226), .A1(n4204), .B0(n4274), .Y(P1_U3243));
  XOR2X1  g3203(.A(n2078), .B(n2055), .Y(n4276));
  XOR2X1  g3204(.A(n4276), .B(n3769), .Y(n4277));
  INVX1   g3205(.A(P1_REG3_REG_1__SCAN_IN), .Y(n4278));
  OAI22X1 g3206(.A0(P1_STATE_REG_SCAN_IN), .A1(n4278), .B0(n1137), .B1(n3923), .Y(n4279));
  AOI21X1 g3207(.A0(n4277), .A1(n3920), .B0(n4279), .Y(n4280));
  XOR2X1  g3208(.A(n2078), .B(P1_REG1_REG_1__SCAN_IN), .Y(n4281));
  XOR2X1  g3209(.A(n4281), .B(n3861), .Y(n4282));
  NAND2X1 g3210(.A(n4282), .B(n3919), .Y(n4283));
  AOI22X1 g3211(.A0(n4277), .A1(n3825), .B0(n3824), .B1(n4282), .Y(n4284));
  OAI21X1 g3212(.A0(n3910), .A1(n2078), .B0(n4284), .Y(n4285));
  AOI22X1 g3213(.A0(n3922), .A1(n3768), .B0(n3739), .B1(n4285), .Y(n4286));
  NAND3X1 g3214(.A(n4286), .B(n4283), .C(n4280), .Y(P1_U3242));
  XOR2X1  g3215(.A(n2008), .B(P1_REG2_REG_0__SCAN_IN), .Y(n4288));
  NAND2X1 g3216(.A(n4288), .B(n3920), .Y(n4289));
  AOI22X1 g3217(.A0(P1_U3084), .A1(P1_REG3_REG_0__SCAN_IN), .B0(P1_ADDR_REG_0__SCAN_IN), .B1(n3918), .Y(n4290));
  XOR2X1  g3218(.A(n2008), .B(P1_REG1_REG_0__SCAN_IN), .Y(n4291));
  NAND2X1 g3219(.A(n4291), .B(n3919), .Y(n4292));
  AOI22X1 g3220(.A0(n4288), .A1(n3825), .B0(n3824), .B1(n4291), .Y(n4293));
  OAI21X1 g3221(.A0(n3910), .A1(n4210), .B0(n4293), .Y(n4294));
  AOI22X1 g3222(.A0(n3922), .A1(n2008), .B0(n3739), .B1(n4294), .Y(n4295));
  NAND4X1 g3223(.A(n4292), .B(n4290), .C(n4289), .D(n4295), .Y(P1_U3241));
  NAND2X1 g3224(.A(n4204), .B(P1_DATAO_REG_0__SCAN_IN), .Y(n4297));
  OAI21X1 g3225(.A0(n4204), .A1(n2036), .B0(n4297), .Y(P1_U3555));
  NAND2X1 g3226(.A(n4204), .B(P1_DATAO_REG_1__SCAN_IN), .Y(n4299));
  OAI21X1 g3227(.A0(n4204), .A1(n2076), .B0(n4299), .Y(P1_U3556));
  NAND2X1 g3228(.A(n4204), .B(P1_DATAO_REG_2__SCAN_IN), .Y(n4301));
  OAI21X1 g3229(.A0(n4204), .A1(n2111), .B0(n4301), .Y(P1_U3557));
  NAND2X1 g3230(.A(n4204), .B(P1_DATAO_REG_3__SCAN_IN), .Y(n4303));
  OAI21X1 g3231(.A0(n4204), .A1(n2154), .B0(n4303), .Y(P1_U3558));
  OAI21X1 g3232(.A0(n2206), .A1(n2271), .B0(P1_U4006), .Y(n4305));
  OAI21X1 g3233(.A0(P1_U4006), .A1(n1234), .B0(n4305), .Y(P1_U3559));
  NAND2X1 g3234(.A(n4204), .B(P1_DATAO_REG_5__SCAN_IN), .Y(n4307));
  OAI21X1 g3235(.A0(n4204), .A1(n2263), .B0(n4307), .Y(P1_U3560));
  NAND2X1 g3236(.A(n4204), .B(P1_DATAO_REG_6__SCAN_IN), .Y(n4309));
  OAI21X1 g3237(.A0(n4204), .A1(n2338), .B0(n4309), .Y(P1_U3561));
  NAND2X1 g3238(.A(n4204), .B(P1_DATAO_REG_7__SCAN_IN), .Y(n4311));
  OAI21X1 g3239(.A0(n4204), .A1(n2366), .B0(n4311), .Y(P1_U3562));
  NAND2X1 g3240(.A(n4204), .B(P1_DATAO_REG_8__SCAN_IN), .Y(n4313));
  OAI21X1 g3241(.A0(n4204), .A1(n2411), .B0(n4313), .Y(P1_U3563));
  NAND2X1 g3242(.A(n4204), .B(P1_DATAO_REG_9__SCAN_IN), .Y(n4315));
  OAI21X1 g3243(.A0(n4204), .A1(n2454), .B0(n4315), .Y(P1_U3564));
  NAND2X1 g3244(.A(n4204), .B(P1_DATAO_REG_10__SCAN_IN), .Y(n4317));
  OAI21X1 g3245(.A0(n4204), .A1(n2499), .B0(n4317), .Y(P1_U3565));
  NAND2X1 g3246(.A(n4204), .B(P1_DATAO_REG_11__SCAN_IN), .Y(n4319));
  OAI21X1 g3247(.A0(n4204), .A1(n2546), .B0(n4319), .Y(P1_U3566));
  NAND2X1 g3248(.A(n4204), .B(P1_DATAO_REG_12__SCAN_IN), .Y(n4321));
  OAI21X1 g3249(.A0(n4204), .A1(n2594), .B0(n4321), .Y(P1_U3567));
  NAND2X1 g3250(.A(n4204), .B(P1_DATAO_REG_13__SCAN_IN), .Y(n4323));
  OAI21X1 g3251(.A0(n4204), .A1(n2635), .B0(n4323), .Y(P1_U3568));
  NAND2X1 g3252(.A(n4204), .B(P1_DATAO_REG_14__SCAN_IN), .Y(n4325));
  OAI21X1 g3253(.A0(n4204), .A1(n2682), .B0(n4325), .Y(P1_U3569));
  NAND2X1 g3254(.A(n4204), .B(P1_DATAO_REG_15__SCAN_IN), .Y(n4327));
  OAI21X1 g3255(.A0(n4204), .A1(n2726), .B0(n4327), .Y(P1_U3570));
  NAND2X1 g3256(.A(n4204), .B(P1_DATAO_REG_16__SCAN_IN), .Y(n4329));
  OAI21X1 g3257(.A0(n4204), .A1(n2765), .B0(n4329), .Y(P1_U3571));
  NAND2X1 g3258(.A(n4204), .B(P1_DATAO_REG_17__SCAN_IN), .Y(n4331));
  OAI21X1 g3259(.A0(n4204), .A1(n2812), .B0(n4331), .Y(P1_U3572));
  NAND2X1 g3260(.A(n4204), .B(P1_DATAO_REG_18__SCAN_IN), .Y(n4333));
  OAI21X1 g3261(.A0(n4204), .A1(n2864), .B0(n4333), .Y(P1_U3573));
  NAND2X1 g3262(.A(n4204), .B(P1_DATAO_REG_19__SCAN_IN), .Y(n4335));
  OAI21X1 g3263(.A0(n4204), .A1(n2906), .B0(n4335), .Y(P1_U3574));
  NAND2X1 g3264(.A(n4204), .B(P1_DATAO_REG_20__SCAN_IN), .Y(n4337));
  OAI21X1 g3265(.A0(n4204), .A1(n2949), .B0(n4337), .Y(P1_U3575));
  NAND2X1 g3266(.A(n4204), .B(P1_DATAO_REG_21__SCAN_IN), .Y(n4339));
  OAI21X1 g3267(.A0(n4204), .A1(n2993), .B0(n4339), .Y(P1_U3576));
  NAND2X1 g3268(.A(n4204), .B(P1_DATAO_REG_22__SCAN_IN), .Y(n4341));
  OAI21X1 g3269(.A0(n4204), .A1(n3035), .B0(n4341), .Y(P1_U3577));
  NAND2X1 g3270(.A(n4204), .B(P1_DATAO_REG_23__SCAN_IN), .Y(n4343));
  OAI21X1 g3271(.A0(n4204), .A1(n3072), .B0(n4343), .Y(P1_U3578));
  NAND2X1 g3272(.A(n4204), .B(P1_DATAO_REG_24__SCAN_IN), .Y(n4345));
  OAI21X1 g3273(.A0(n4204), .A1(n3123), .B0(n4345), .Y(P1_U3579));
  NAND2X1 g3274(.A(n4204), .B(P1_DATAO_REG_25__SCAN_IN), .Y(n4347));
  OAI21X1 g3275(.A0(n4204), .A1(n3159), .B0(n4347), .Y(P1_U3580));
  NAND2X1 g3276(.A(n4204), .B(P1_DATAO_REG_26__SCAN_IN), .Y(n4349));
  OAI21X1 g3277(.A0(n4204), .A1(n3199), .B0(n4349), .Y(P1_U3581));
  NAND2X1 g3278(.A(n4204), .B(P1_DATAO_REG_27__SCAN_IN), .Y(n4351));
  OAI21X1 g3279(.A0(n4204), .A1(n3253), .B0(n4351), .Y(P1_U3582));
  NAND2X1 g3280(.A(n4204), .B(P1_DATAO_REG_28__SCAN_IN), .Y(n4353));
  OAI21X1 g3281(.A0(n4204), .A1(n3290), .B0(n4353), .Y(P1_U3583));
  NAND2X1 g3282(.A(n4204), .B(P1_DATAO_REG_29__SCAN_IN), .Y(n4355));
  OAI21X1 g3283(.A0(n4204), .A1(n3329), .B0(n4355), .Y(P1_U3584));
  INVX1   g3284(.A(n3353), .Y(n4357));
  NAND2X1 g3285(.A(n4204), .B(P1_DATAO_REG_30__SCAN_IN), .Y(n4358));
  OAI21X1 g3286(.A0(n4204), .A1(n4357), .B0(n4358), .Y(P1_U3585));
  INVX1   g3287(.A(n3385), .Y(n4360));
  NAND2X1 g3288(.A(n4204), .B(P1_DATAO_REG_31__SCAN_IN), .Y(n4361));
  OAI21X1 g3289(.A0(n4204), .A1(n4360), .B0(n4361), .Y(P1_U3586));
  XOR2X1  g3290(.A(n3382), .B(n4357), .Y(n4363));
  XOR2X1  g3291(.A(n3398), .B(n3385), .Y(n4364));
  XOR2X1  g3292(.A(n3345), .B(n3328), .Y(n4365));
  XOR2X1  g3293(.A(n3324), .B(n3290), .Y(n4366));
  XOR2X1  g3294(.A(n2956), .B(n2948), .Y(n4372));
  XOR2X1  g3295(.A(n2385), .B(n2365), .Y(n4374));
  INVX1   g3296(.A(n2123), .Y(n4375));
  NAND3X1 g3297(.A(n2026), .B(n4375), .C(n2082), .Y(n4377));
  NOR4X1  g3298(.A(n4374), .B(n2235), .C(n2177), .D(n4377), .Y(n4378));
  NAND4X1 g3299(.A(n4378), .B(n2470), .C(n2344), .D(n2293), .Y(n4380));
  NAND3X1 g3300(.A(n2519), .B(n2577), .C(n2426), .Y(n4383));
  NAND4X1 g3301(.A(n2738), .B(n2661), .C(n2608), .D(n2694), .Y(n4387));
  NOR4X1  g3302(.A(n4383), .B(n4380), .C(n2794), .D(n4387), .Y(n4388));
  NAND2X1 g3303(.A(n4388), .B(n2838), .Y(n4389));
  NOR4X1  g3304(.A(n4372), .B(n2927), .C(n2883), .D(n4389), .Y(n4390));
  NAND4X1 g3305(.A(n3001), .B(n3043), .C(n3086), .D(n4390), .Y(n4391));
  NOR3X1  g3306(.A(n4391), .B(n3180), .C(n3141), .Y(n4392));
  NAND3X1 g3307(.A(n4392), .B(n3207), .C(n3256), .Y(n4393));
  NOR3X1  g3308(.A(n4393), .B(n4366), .C(n4365), .Y(n4394));
  NAND2X1 g3309(.A(n4394), .B(n4364), .Y(n4395));
  NOR2X1  g3310(.A(n4395), .B(n4363), .Y(n4396));
  NOR3X1  g3311(.A(n4396), .B(n1993), .C(n1874), .Y(n4397));
  NOR4X1  g3312(.A(n4363), .B(n2041), .C(n1874), .D(n4395), .Y(n4398));
  OAI21X1 g3313(.A0(n4398), .A1(n4397), .B0(n1989), .Y(n4399));
  OAI21X1 g3314(.A0(n1993), .A1(n1985), .B0(n1875), .Y(n4400));
  INVX1   g3315(.A(n4400), .Y(n4401));
  AOI22X1 g3316(.A0(n4401), .A1(n3385), .B0(n3396), .B1(n2066), .Y(n4404));
  INVX1   g3317(.A(n2066), .Y(n4405));
  OAI22X1 g3318(.A0(n4400), .A1(n3398), .B0(n4405), .B1(n4360), .Y(n4407));
  XOR2X1  g3319(.A(n4407), .B(n4404), .Y(n4408));
  NAND3X1 g3320(.A(n3385), .B(n3353), .C(n2066), .Y(n4409));
  OAI21X1 g3321(.A0(n4400), .A1(n3382), .B0(n4409), .Y(n4410));
  NAND3X1 g3322(.A(n2066), .B(n2101), .C(n3728), .Y(n4411));
  NAND3X1 g3323(.A(n4401), .B(n3385), .C(n3353), .Y(n4412));
  NAND3X1 g3324(.A(n4412), .B(n4411), .C(n4410), .Y(n4413));
  AOI22X1 g3325(.A0(n3289), .A1(n1874), .B0(n2066), .B1(n3328), .Y(n4414));
  INVX1   g3326(.A(n4414), .Y(n4415));
  AOI21X1 g3327(.A0(n4401), .A1(n3345), .B0(n4415), .Y(n4416));
  NOR3X1  g3328(.A(n4405), .B(n2005), .C(n1822), .Y(n4417));
  OAI21X1 g3329(.A0(n4400), .A1(n3329), .B0(n1875), .Y(n4418));
  NOR3X1  g3330(.A(n4418), .B(n4417), .C(n4416), .Y(n4419));
  AOI22X1 g3331(.A0(n3243), .A1(n1874), .B0(n2066), .B1(n3289), .Y(n4420));
  INVX1   g3332(.A(n4420), .Y(n4421));
  AOI21X1 g3333(.A0(n4401), .A1(n3297), .B0(n4421), .Y(n4422));
  NAND3X1 g3334(.A(n2066), .B(n2101), .C(n3323), .Y(n4423));
  AOI21X1 g3335(.A0(n4401), .A1(n3289), .B0(n1874), .Y(n4424));
  NAND2X1 g3336(.A(n4424), .B(n4423), .Y(n4425));
  NOR2X1  g3337(.A(n4425), .B(n4422), .Y(n4426));
  AOI22X1 g3338(.A0(n3198), .A1(n1874), .B0(n2066), .B1(n3243), .Y(n4427));
  INVX1   g3339(.A(n4427), .Y(n4428));
  AOI21X1 g3340(.A0(n4401), .A1(n3255), .B0(n4428), .Y(n4429));
  INVX1   g3341(.A(n4429), .Y(n4430));
  AOI21X1 g3342(.A0(n4401), .A1(n3243), .B0(n1874), .Y(n4431));
  INVX1   g3343(.A(n4431), .Y(n4432));
  AOI21X1 g3344(.A0(n3255), .A1(n2066), .B0(n4432), .Y(n4433));
  NOR2X1  g3345(.A(n4433), .B(n4430), .Y(n4434));
  AOI21X1 g3346(.A0(n4425), .A1(n4422), .B0(n4434), .Y(n4435));
  NOR3X1  g3347(.A(n4435), .B(n4426), .C(n4419), .Y(n4436));
  NAND3X1 g3348(.A(n4436), .B(n4413), .C(n4408), .Y(n4437));
  NOR4X1  g3349(.A(n4404), .B(n2066), .C(n1875), .D(n4407), .Y(n4438));
  OAI22X1 g3350(.A0(n4400), .A1(n4360), .B0(n3398), .B1(n4405), .Y(n4439));
  AOI21X1 g3351(.A0(n4405), .A1(n1874), .B0(n4439), .Y(n4440));
  AOI21X1 g3352(.A0(n4440), .A1(n4407), .B0(n4438), .Y(n4441));
  XOR2X1  g3353(.A(n4407), .B(n4439), .Y(n4442));
  NAND3X1 g3354(.A(n4401), .B(n2101), .C(n3728), .Y(n4443));
  OAI21X1 g3355(.A0(n3382), .A1(n4405), .B0(n4412), .Y(n4444));
  AOI21X1 g3356(.A0(n4443), .A1(n4409), .B0(n4444), .Y(n4445));
  OAI21X1 g3357(.A0(n4400), .A1(n3324), .B0(n4420), .Y(n4446));
  NAND3X1 g3358(.A(n4424), .B(n4423), .C(n4446), .Y(n4447));
  NAND2X1 g3359(.A(n4433), .B(n4430), .Y(n4448));
  NOR3X1  g3360(.A(n4405), .B(n2005), .C(n1728), .Y(n4449));
  OAI21X1 g3361(.A0(n4400), .A1(n3159), .B0(n1875), .Y(n4450));
  AOI22X1 g3362(.A0(n3117), .A1(n1874), .B0(n2066), .B1(n3158), .Y(n4451));
  INVX1   g3363(.A(n4451), .Y(n4452));
  AOI21X1 g3364(.A0(n4401), .A1(n3166), .B0(n4452), .Y(n4453));
  OAI21X1 g3365(.A0(n4450), .A1(n4449), .B0(n4453), .Y(n4454));
  NOR3X1  g3366(.A(n4405), .B(n2005), .C(n1746), .Y(n4455));
  OAI21X1 g3367(.A0(n4400), .A1(n3199), .B0(n1875), .Y(n4456));
  NOR2X1  g3368(.A(n4456), .B(n4455), .Y(n4457));
  AOI22X1 g3369(.A0(n3158), .A1(n1874), .B0(n2066), .B1(n3198), .Y(n4458));
  OAI21X1 g3370(.A0(n4400), .A1(n3266), .B0(n4458), .Y(n4459));
  OAI21X1 g3371(.A0(n4459), .A1(n4457), .B0(n4454), .Y(n4460));
  NAND2X1 g3372(.A(n4459), .B(n4457), .Y(n4461));
  NAND4X1 g3373(.A(n4460), .B(n4448), .C(n4447), .D(n4461), .Y(n4462));
  NOR4X1  g3374(.A(n4419), .B(n4445), .C(n4442), .D(n4462), .Y(n4463));
  OAI21X1 g3375(.A0(n4400), .A1(n3123), .B0(n1875), .Y(n4464));
  AOI21X1 g3376(.A0(n3124), .A1(n2066), .B0(n4464), .Y(n4465));
  AOI22X1 g3377(.A0(n3071), .A1(n1874), .B0(n2066), .B1(n3117), .Y(n4466));
  OAI21X1 g3378(.A0(n4400), .A1(n3151), .B0(n4466), .Y(n4467));
  OAI21X1 g3379(.A0(n4400), .A1(n3072), .B0(n1875), .Y(n4468));
  AOI21X1 g3380(.A0(n3111), .A1(n2066), .B0(n4468), .Y(n4469));
  AOI22X1 g3381(.A0(n3080), .A1(n1874), .B0(n2066), .B1(n3071), .Y(n4470));
  OAI21X1 g3382(.A0(n4400), .A1(n3085), .B0(n4470), .Y(n4471));
  OAI22X1 g3383(.A0(n4469), .A1(n4471), .B0(n4467), .B1(n4465), .Y(n4472));
  AOI21X1 g3384(.A0(n4401), .A1(n2948), .B0(n1874), .Y(n4473));
  OAI21X1 g3385(.A0(n2968), .A1(n4405), .B0(n4473), .Y(n4474));
  OAI22X1 g3386(.A0(n2906), .A1(n1875), .B0(n4405), .B1(n2949), .Y(n4475));
  AOI21X1 g3387(.A0(n4401), .A1(n2956), .B0(n4475), .Y(n4476));
  NAND2X1 g3388(.A(n4476), .B(n4474), .Y(n4477));
  OAI21X1 g3389(.A0(n4400), .A1(n2906), .B0(n1875), .Y(n4478));
  AOI21X1 g3390(.A0(n2914), .A1(n2066), .B0(n4478), .Y(n4479));
  AOI22X1 g3391(.A0(n2863), .A1(n1874), .B0(n2066), .B1(n2926), .Y(n4480));
  OAI21X1 g3392(.A0(n4400), .A1(n2939), .B0(n4480), .Y(n4481));
  NOR2X1  g3393(.A(n4481), .B(n4479), .Y(n4482));
  OAI21X1 g3394(.A0(n4400), .A1(n2682), .B0(n1875), .Y(n4483));
  AOI21X1 g3395(.A0(n2718), .A1(n2066), .B0(n4483), .Y(n4484));
  AOI22X1 g3396(.A0(n2634), .A1(n1874), .B0(n2066), .B1(n2681), .Y(n4485));
  OAI21X1 g3397(.A0(n4400), .A1(n2693), .B0(n4485), .Y(n4486));
  NOR2X1  g3398(.A(n4486), .B(n4484), .Y(n4487));
  OAI21X1 g3399(.A0(n4400), .A1(n2635), .B0(n1875), .Y(n4488));
  AOI21X1 g3400(.A0(n2649), .A1(n2066), .B0(n4488), .Y(n4489));
  AOI22X1 g3401(.A0(n2593), .A1(n1874), .B0(n2066), .B1(n2634), .Y(n4490));
  OAI21X1 g3402(.A0(n4400), .A1(n2653), .B0(n4490), .Y(n4491));
  NOR2X1  g3403(.A(n4491), .B(n4489), .Y(n4492));
  OAI21X1 g3404(.A0(n2206), .A1(n2271), .B0(n4401), .Y(n4493));
  AOI21X1 g3405(.A0(n2222), .A1(n2066), .B0(n1874), .Y(n4494));
  NAND2X1 g3406(.A(n4494), .B(n4493), .Y(n4495));
  OAI21X1 g3407(.A0(n2206), .A1(n2271), .B0(n2066), .Y(n4496));
  AOI22X1 g3408(.A0(n2222), .A1(n4401), .B0(n2167), .B1(n1874), .Y(n4497));
  NAND3X1 g3409(.A(n4497), .B(n4496), .C(n4495), .Y(n4498));
  OAI21X1 g3410(.A0(n2153), .A1(n2149), .B0(n4401), .Y(n4499));
  AOI21X1 g3411(.A0(n2172), .A1(n2066), .B0(n1874), .Y(n4500));
  OAI21X1 g3412(.A0(n2153), .A1(n2149), .B0(n2066), .Y(n4501));
  AOI22X1 g3413(.A0(n2172), .A1(n4401), .B0(n2110), .B1(n1874), .Y(n4502));
  NAND2X1 g3414(.A(n4502), .B(n4501), .Y(n4503));
  AOI21X1 g3415(.A0(n4500), .A1(n4499), .B0(n4503), .Y(n4504));
  NAND2X1 g3416(.A(n4401), .B(n2110), .Y(n4505));
  AOI21X1 g3417(.A0(n2122), .A1(n2066), .B0(n1874), .Y(n4506));
  NAND2X1 g3418(.A(n4506), .B(n4505), .Y(n4507));
  NAND2X1 g3419(.A(n2110), .B(n2066), .Y(n4508));
  AOI22X1 g3420(.A0(n2122), .A1(n4401), .B0(n2062), .B1(n1874), .Y(n4509));
  NAND3X1 g3421(.A(n4509), .B(n4508), .C(n4507), .Y(n4510));
  NAND2X1 g3422(.A(n4509), .B(n4508), .Y(n4511));
  NAND3X1 g3423(.A(n4511), .B(n4506), .C(n4505), .Y(n4512));
  AOI21X1 g3424(.A0(n2081), .A1(n2066), .B0(n1874), .Y(n4514));
  OAI21X1 g3425(.A0(n2076), .A1(n4400), .B0(n4514), .Y(n4515));
  NOR2X1  g3426(.A(n2076), .B(n4405), .Y(n4516));
  OAI22X1 g3427(.A0(n2102), .A1(n4400), .B0(n2036), .B1(n1875), .Y(n4517));
  NOR2X1  g3428(.A(n4517), .B(n4516), .Y(n4518));
  NAND3X1 g3429(.A(n4518), .B(n4515), .C(n4512), .Y(n4519));
  NAND2X1 g3430(.A(n4500), .B(n4499), .Y(n4520));
  AOI21X1 g3431(.A0(n4502), .A1(n4501), .B0(n4520), .Y(n4521));
  AOI21X1 g3432(.A0(n4519), .A1(n4510), .B0(n4521), .Y(n4522));
  AOI21X1 g3433(.A0(n4497), .A1(n4496), .B0(n4495), .Y(n4523));
  INVX1   g3434(.A(n4523), .Y(n4524));
  OAI21X1 g3435(.A0(n4522), .A1(n4504), .B0(n4524), .Y(n4525));
  NAND2X1 g3436(.A(n4401), .B(n2279), .Y(n4526));
  AOI22X1 g3437(.A0(n2208), .A1(n1874), .B0(n2066), .B1(n2274), .Y(n4527));
  AOI21X1 g3438(.A0(n4401), .A1(n2274), .B0(n1874), .Y(n4528));
  OAI21X1 g3439(.A0(n2284), .A1(n4405), .B0(n4528), .Y(n4529));
  AOI21X1 g3440(.A0(n4527), .A1(n4526), .B0(n4529), .Y(n4530));
  AOI21X1 g3441(.A0(n4525), .A1(n4498), .B0(n4530), .Y(n4531));
  OAI21X1 g3442(.A0(n4518), .A1(n4515), .B0(n4512), .Y(n4532));
  OAI22X1 g3443(.A0(n4405), .A1(n2036), .B0(n2010), .B1(n4400), .Y(n4533));
  OAI21X1 g3444(.A0(n4405), .A1(n2010), .B0(n1875), .Y(n4535));
  AOI21X1 g3445(.A0(n2025), .A1(n4401), .B0(n4535), .Y(n4536));
  NOR3X1  g3446(.A(n1993), .B(n1985), .C(n1874), .Y(n4537));
  OAI21X1 g3447(.A0(n4537), .A1(n4536), .B0(n4533), .Y(n4538));
  AOI21X1 g3448(.A0(n4537), .A1(n4536), .B0(n4521), .Y(n4539));
  NAND2X1 g3449(.A(n4539), .B(n4538), .Y(n4540));
  NOR4X1  g3450(.A(n4532), .B(n4530), .C(n4523), .D(n4540), .Y(n4541));
  AOI22X1 g3451(.A0(n2274), .A1(n1874), .B0(n2066), .B1(n2316), .Y(n4542));
  OAI21X1 g3452(.A0(n4400), .A1(n2332), .B0(n4542), .Y(n4543));
  OAI21X1 g3453(.A0(n4400), .A1(n2338), .B0(n1875), .Y(n4544));
  AOI21X1 g3454(.A0(n2340), .A1(n2066), .B0(n4544), .Y(n4545));
  NAND3X1 g3455(.A(n4529), .B(n4527), .C(n4526), .Y(n4546));
  OAI21X1 g3456(.A0(n4545), .A1(n4543), .B0(n4546), .Y(n4547));
  NOR3X1  g3457(.A(n4547), .B(n4541), .C(n4531), .Y(n4548));
  NAND2X1 g3458(.A(n4401), .B(n2469), .Y(n4549));
  AOI22X1 g3459(.A0(n2410), .A1(n1874), .B0(n2066), .B1(n2453), .Y(n4550));
  NAND2X1 g3460(.A(n4550), .B(n4549), .Y(n4551));
  AOI21X1 g3461(.A0(n4401), .A1(n2453), .B0(n1874), .Y(n4552));
  INVX1   g3462(.A(n4552), .Y(n4553));
  AOI21X1 g3463(.A0(n2469), .A1(n2066), .B0(n4553), .Y(n4554));
  NAND2X1 g3464(.A(n4554), .B(n4551), .Y(n4555));
  AOI22X1 g3465(.A0(n2365), .A1(n1874), .B0(n2066), .B1(n2410), .Y(n4556));
  OAI21X1 g3466(.A0(n4400), .A1(n2445), .B0(n4556), .Y(n4557));
  OAI21X1 g3467(.A0(n4400), .A1(n2411), .B0(n1875), .Y(n4558));
  AOI21X1 g3468(.A0(n2425), .A1(n2066), .B0(n4558), .Y(n4559));
  NAND2X1 g3469(.A(n4559), .B(n4557), .Y(n4560));
  AOI22X1 g3470(.A0(n2316), .A1(n1874), .B0(n2066), .B1(n2365), .Y(n4561));
  OAI21X1 g3471(.A0(n4400), .A1(n2379), .B0(n4561), .Y(n4562));
  OAI21X1 g3472(.A0(n4400), .A1(n2366), .B0(n1875), .Y(n4563));
  AOI21X1 g3473(.A0(n2385), .A1(n2066), .B0(n4563), .Y(n4564));
  AOI22X1 g3474(.A0(n4562), .A1(n4564), .B0(n4545), .B1(n4543), .Y(n4565));
  NAND3X1 g3475(.A(n4565), .B(n4560), .C(n4555), .Y(n4566));
  OAI21X1 g3476(.A0(n4400), .A1(n2594), .B0(n1875), .Y(n4567));
  AOI21X1 g3477(.A0(n2607), .A1(n2066), .B0(n4567), .Y(n4568));
  AOI22X1 g3478(.A0(n2545), .A1(n1874), .B0(n2066), .B1(n2593), .Y(n4569));
  OAI21X1 g3479(.A0(n4400), .A1(n2627), .B0(n4569), .Y(n4570));
  OAI21X1 g3480(.A0(n4400), .A1(n2546), .B0(n1875), .Y(n4571));
  AOI21X1 g3481(.A0(n2562), .A1(n2066), .B0(n4571), .Y(n4572));
  AOI22X1 g3482(.A0(n2498), .A1(n1874), .B0(n2066), .B1(n2545), .Y(n4573));
  OAI21X1 g3483(.A0(n4400), .A1(n2586), .B0(n4573), .Y(n4574));
  OAI22X1 g3484(.A0(n4572), .A1(n4574), .B0(n4570), .B1(n4568), .Y(n4575));
  NAND2X1 g3485(.A(n4560), .B(n4555), .Y(n4576));
  NOR3X1  g3486(.A(n4564), .B(n4562), .C(n4576), .Y(n4577));
  INVX1   g3487(.A(n4555), .Y(n4578));
  NOR3X1  g3488(.A(n4559), .B(n4557), .C(n4578), .Y(n4579));
  AOI21X1 g3489(.A0(n4401), .A1(n2498), .B0(n1874), .Y(n4580));
  OAI21X1 g3490(.A0(n2512), .A1(n4405), .B0(n4580), .Y(n4581));
  OAI22X1 g3491(.A0(n2454), .A1(n1875), .B0(n4405), .B1(n2499), .Y(n4582));
  AOI21X1 g3492(.A0(n4401), .A1(n2511), .B0(n4582), .Y(n4583));
  NAND2X1 g3493(.A(n4583), .B(n4581), .Y(n4584));
  OAI21X1 g3494(.A0(n4554), .A1(n4551), .B0(n4584), .Y(n4585));
  NOR4X1  g3495(.A(n4579), .B(n4577), .C(n4575), .D(n4585), .Y(n4586));
  OAI21X1 g3496(.A0(n4566), .A1(n4548), .B0(n4586), .Y(n4587));
  NOR3X1  g3497(.A(n4583), .B(n4581), .C(n4575), .Y(n4588));
  NOR2X1  g3498(.A(n4570), .B(n4568), .Y(n4589));
  NAND2X1 g3499(.A(n4574), .B(n4572), .Y(n4590));
  AOI22X1 g3500(.A0(n4568), .A1(n4570), .B0(n4491), .B1(n4489), .Y(n4591));
  OAI21X1 g3501(.A0(n4590), .A1(n4589), .B0(n4591), .Y(n4592));
  NOR2X1  g3502(.A(n4592), .B(n4588), .Y(n4593));
  AOI21X1 g3503(.A0(n4593), .A1(n4587), .B0(n4492), .Y(n4594));
  AOI21X1 g3504(.A0(n4486), .A1(n4484), .B0(n4594), .Y(n4595));
  AOI22X1 g3505(.A0(n2681), .A1(n1874), .B0(n2066), .B1(n2727), .Y(n4596));
  OAI21X1 g3506(.A0(n4400), .A1(n2737), .B0(n4596), .Y(n4597));
  AOI21X1 g3507(.A0(n4401), .A1(n2727), .B0(n1874), .Y(n4598));
  OAI21X1 g3508(.A0(n2737), .A1(n4405), .B0(n4598), .Y(n4599));
  INVX1   g3509(.A(n4599), .Y(n4600));
  NAND2X1 g3510(.A(n4600), .B(n4597), .Y(n4601));
  OAI21X1 g3511(.A0(n4595), .A1(n4487), .B0(n4601), .Y(n4602));
  AOI21X1 g3512(.A0(n4401), .A1(n2863), .B0(n1874), .Y(n4603));
  OAI21X1 g3513(.A0(n2880), .A1(n4405), .B0(n4603), .Y(n4604));
  OAI22X1 g3514(.A0(n2812), .A1(n1875), .B0(n4405), .B1(n2864), .Y(n4605));
  AOI21X1 g3515(.A0(n4401), .A1(n2898), .B0(n4605), .Y(n4606));
  NAND2X1 g3516(.A(n4606), .B(n4604), .Y(n4607));
  AOI21X1 g3517(.A0(n4401), .A1(n2811), .B0(n1874), .Y(n4608));
  OAI21X1 g3518(.A0(n2824), .A1(n4405), .B0(n4608), .Y(n4609));
  AOI22X1 g3519(.A0(n2764), .A1(n1874), .B0(n2066), .B1(n2811), .Y(n4610));
  INVX1   g3520(.A(n4610), .Y(n4611));
  AOI21X1 g3521(.A0(n4401), .A1(n2825), .B0(n4611), .Y(n4612));
  NAND2X1 g3522(.A(n4612), .B(n4609), .Y(n4613));
  NAND2X1 g3523(.A(n4613), .B(n4607), .Y(n4614));
  OAI21X1 g3524(.A0(n4400), .A1(n2765), .B0(n1875), .Y(n4615));
  AOI21X1 g3525(.A0(n2784), .A1(n2066), .B0(n4615), .Y(n4616));
  AOI22X1 g3526(.A0(n2727), .A1(n1874), .B0(n2066), .B1(n2764), .Y(n4617));
  OAI21X1 g3527(.A0(n4400), .A1(n2779), .B0(n4617), .Y(n4618));
  OAI22X1 g3528(.A0(n4616), .A1(n4618), .B0(n4600), .B1(n4597), .Y(n4619));
  NOR2X1  g3529(.A(n4619), .B(n4614), .Y(n4620));
  NAND4X1 g3530(.A(n4616), .B(n4613), .C(n4607), .D(n4618), .Y(n4621));
  NAND2X1 g3531(.A(n4481), .B(n4479), .Y(n4622));
  NOR2X1  g3532(.A(n4606), .B(n4604), .Y(n4623));
  NOR2X1  g3533(.A(n4612), .B(n4609), .Y(n4624));
  AOI21X1 g3534(.A0(n4624), .A1(n4607), .B0(n4623), .Y(n4625));
  NAND3X1 g3535(.A(n4625), .B(n4622), .C(n4621), .Y(n4626));
  AOI21X1 g3536(.A0(n4620), .A1(n4602), .B0(n4626), .Y(n4627));
  OAI22X1 g3537(.A0(n4482), .A1(n4627), .B0(n4476), .B1(n4474), .Y(n4628));
  OAI21X1 g3538(.A0(n4400), .A1(n2993), .B0(n1875), .Y(n4629));
  AOI21X1 g3539(.A0(n3000), .A1(n2066), .B0(n4629), .Y(n4630));
  AOI22X1 g3540(.A0(n2948), .A1(n1874), .B0(n2066), .B1(n2994), .Y(n4631));
  OAI21X1 g3541(.A0(n4400), .A1(n3028), .B0(n4631), .Y(n4632));
  AOI22X1 g3542(.A0(n4630), .A1(n4632), .B0(n4628), .B1(n4477), .Y(n4633));
  AOI21X1 g3543(.A0(n4401), .A1(n3080), .B0(n1874), .Y(n4634));
  OAI21X1 g3544(.A0(n3064), .A1(n4405), .B0(n4634), .Y(n4635));
  AOI22X1 g3545(.A0(n2994), .A1(n1874), .B0(n2066), .B1(n3080), .Y(n4636));
  INVX1   g3546(.A(n4636), .Y(n4637));
  AOI21X1 g3547(.A0(n4401), .A1(n3042), .B0(n4637), .Y(n4638));
  NAND2X1 g3548(.A(n4638), .B(n4635), .Y(n4639));
  OAI21X1 g3549(.A0(n4632), .A1(n4630), .B0(n4639), .Y(n4640));
  NOR3X1  g3550(.A(n4640), .B(n4633), .C(n4472), .Y(n4641));
  NOR2X1  g3551(.A(n4467), .B(n4465), .Y(n4642));
  NAND2X1 g3552(.A(n4467), .B(n4465), .Y(n4643));
  NAND2X1 g3553(.A(n4471), .B(n4469), .Y(n4644));
  OAI21X1 g3554(.A0(n4644), .A1(n4642), .B0(n4643), .Y(n4645));
  NOR3X1  g3555(.A(n4453), .B(n4450), .C(n4449), .Y(n4646));
  NOR3X1  g3556(.A(n4638), .B(n4635), .C(n4472), .Y(n4647));
  NOR4X1  g3557(.A(n4646), .B(n4645), .C(n4641), .D(n4647), .Y(n4648));
  NAND4X1 g3558(.A(n4461), .B(n4448), .C(n4447), .D(n4648), .Y(n4649));
  NOR4X1  g3559(.A(n4419), .B(n4445), .C(n4442), .D(n4649), .Y(n4650));
  NAND3X1 g3560(.A(n4444), .B(n4443), .C(n4409), .Y(n4651));
  NOR2X1  g3561(.A(n4651), .B(n4442), .Y(n4652));
  OAI21X1 g3562(.A0(n4418), .A1(n4417), .B0(n4416), .Y(n4653));
  NOR3X1  g3563(.A(n4653), .B(n4445), .C(n4442), .Y(n4654));
  NOR4X1  g3564(.A(n4652), .B(n4650), .C(n4463), .D(n4654), .Y(n4655));
  NOR3X1  g3565(.A(n1989), .B(n1985), .C(n1874), .Y(n4656));
  NAND4X1 g3566(.A(n4655), .B(n4441), .C(n4437), .D(n4656), .Y(n4657));
  AOI21X1 g3567(.A0(n4657), .A1(n4399), .B0(n1987), .Y(n4658));
  AOI21X1 g3568(.A0(n2101), .A1(n3323), .B0(n3290), .Y(n4659));
  NOR4X1  g3569(.A(n3260), .B(n3179), .C(n3158), .D(n4659), .Y(n4660));
  OAI21X1 g3570(.A0(n3398), .A1(n3385), .B0(n4660), .Y(n4661));
  NOR4X1  g3571(.A(n3089), .B(n3042), .C(n3035), .D(n3138), .Y(n4662));
  NOR3X1  g3572(.A(n3138), .B(n3111), .C(n3072), .Y(n4663));
  NOR4X1  g3573(.A(n4662), .B(n3210), .C(n3139), .D(n4663), .Y(n4664));
  NAND4X1 g3574(.A(n3360), .B(n3256), .C(n3249), .D(n4664), .Y(n4665));
  NOR2X1  g3575(.A(n4659), .B(n3301), .Y(n4666));
  OAI21X1 g3576(.A0(n3398), .A1(n3385), .B0(n4666), .Y(n4667));
  NOR3X1  g3577(.A(n4659), .B(n3260), .C(n3252), .Y(n4668));
  OAI22X1 g3578(.A0(n3398), .A1(n3385), .B0(n3362), .B1(n4668), .Y(n4669));
  NAND4X1 g3579(.A(n4667), .B(n4665), .C(n4661), .D(n4669), .Y(n4670));
  AOI22X1 g3580(.A0(n3353), .A1(n3382), .B0(n3372), .B1(n3328), .Y(n4671));
  NOR3X1  g3581(.A(n3328), .B(n2005), .C(n1822), .Y(n4672));
  OAI21X1 g3582(.A0(n3380), .A1(n4357), .B0(n4672), .Y(n4673));
  NAND2X1 g3583(.A(n3396), .B(n4360), .Y(n4674));
  NOR2X1  g3584(.A(n3382), .B(n3353), .Y(n4675));
  NAND2X1 g3585(.A(n4675), .B(n4674), .Y(n4676));
  NAND2X1 g3586(.A(n3398), .B(n3385), .Y(n4677));
  NAND3X1 g3587(.A(n4677), .B(n4676), .C(n4673), .Y(n4678));
  AOI21X1 g3588(.A0(n4671), .A1(n4670), .B0(n4678), .Y(n4679));
  OAI21X1 g3589(.A0(n3398), .A1(n3385), .B0(n3362), .Y(n4680));
  NAND2X1 g3590(.A(n3382), .B(n3353), .Y(n4681));
  AOI22X1 g3591(.A0(n4666), .A1(n4674), .B0(n4672), .B1(n4681), .Y(n4682));
  NAND4X1 g3592(.A(n3256), .B(n3206), .C(n3199), .D(n3360), .Y(n4683));
  AOI21X1 g3593(.A0(n3396), .A1(n4360), .B0(n4683), .Y(n4684));
  NOR2X1  g3594(.A(n3396), .B(n4360), .Y(n4685));
  INVX1   g3595(.A(n2741), .Y(n4686));
  NOR3X1  g3596(.A(n2527), .B(n2433), .C(n2341), .Y(n4687));
  OAI21X1 g3597(.A0(n2425), .A1(n2411), .B0(n4687), .Y(n4688));
  INVX1   g3598(.A(n2286), .Y(n4689));
  AOI21X1 g3599(.A0(n2132), .A1(n1989), .B0(n2037), .Y(n4690));
  AOI21X1 g3600(.A0(n4690), .A1(n2081), .B0(n2076), .Y(n4691));
  NOR2X1  g3601(.A(n4690), .B(n2081), .Y(n4692));
  OAI21X1 g3602(.A0(n2172), .A1(n2154), .B0(n2192), .Y(n4693));
  NOR4X1  g3603(.A(n4692), .B(n4691), .C(n2294), .D(n4693), .Y(n4694));
  OAI21X1 g3604(.A0(n2333), .A1(n4689), .B0(n4694), .Y(n4695));
  AOI22X1 g3605(.A0(n2499), .A1(n2511), .B0(n2469), .B1(n2454), .Y(n4696));
  OAI21X1 g3606(.A0(n4695), .A1(n4688), .B0(n4696), .Y(n4697));
  NAND2X1 g3607(.A(n2425), .B(n2411), .Y(n4698));
  OAI21X1 g3608(.A0(n2425), .A1(n2411), .B0(n2435), .Y(n4699));
  AOI21X1 g3609(.A0(n4699), .A1(n4698), .B0(n2527), .Y(n4700));
  NAND2X1 g3610(.A(n2607), .B(n2594), .Y(n4701));
  NAND2X1 g3611(.A(n4701), .B(n2563), .Y(n4702));
  NOR2X1  g3612(.A(n2333), .B(n4689), .Y(n4703));
  OAI21X1 g3613(.A0(n2172), .A1(n2154), .B0(n2189), .Y(n4704));
  AOI21X1 g3614(.A0(n4704), .A1(n2240), .B0(n2294), .Y(n4705));
  NOR4X1  g3615(.A(n2333), .B(n2285), .C(n2295), .D(n4705), .Y(n4706));
  NOR3X1  g3616(.A(n4706), .B(n4703), .C(n4688), .Y(n4707));
  NOR4X1  g3617(.A(n4702), .B(n4700), .C(n4697), .D(n4707), .Y(n4708));
  NAND3X1 g3618(.A(n4701), .B(n2563), .C(n2553), .Y(n4709));
  OAI22X1 g3619(.A0(n2635), .A1(n2649), .B0(n2607), .B1(n2594), .Y(n4710));
  AOI21X1 g3620(.A0(n4701), .A1(n2564), .B0(n4710), .Y(n4711));
  NAND2X1 g3621(.A(n4711), .B(n4709), .Y(n4712));
  OAI22X1 g3622(.A0(n4708), .A1(n4712), .B0(n2653), .B1(n2634), .Y(n4713));
  AOI21X1 g3623(.A0(n4713), .A1(n4686), .B0(n2739), .Y(n4714));
  NOR2X1  g3624(.A(n2880), .B(n2863), .Y(n4715));
  NOR4X1  g3625(.A(n2832), .B(n2783), .C(n2774), .D(n4715), .Y(n4716));
  OAI21X1 g3626(.A0(n4714), .A1(n2772), .B0(n4716), .Y(n4717));
  NOR2X1  g3627(.A(n2898), .B(n2864), .Y(n4718));
  NOR4X1  g3628(.A(n2832), .B(n2784), .C(n2765), .D(n4715), .Y(n4719));
  NOR3X1  g3629(.A(n4715), .B(n2825), .C(n2812), .Y(n4720));
  NOR4X1  g3630(.A(n4719), .B(n2958), .C(n4718), .D(n4720), .Y(n4721));
  AOI21X1 g3631(.A0(n4721), .A1(n4717), .B0(n2960), .Y(n4722));
  NOR3X1  g3632(.A(n4722), .B(n3016), .C(n3004), .Y(n4723));
  OAI21X1 g3633(.A0(n3016), .A1(n3003), .B0(n3044), .Y(n4724));
  NOR3X1  g3634(.A(n4724), .B(n4723), .C(n3081), .Y(n4725));
  NAND3X1 g3635(.A(n4725), .B(n3168), .C(n3126), .Y(n4726));
  NOR3X1  g3636(.A(n4726), .B(n4685), .C(n4684), .Y(n4727));
  OAI21X1 g3637(.A0(n4675), .A1(n4660), .B0(n4674), .Y(n4728));
  NAND4X1 g3638(.A(n4727), .B(n4682), .C(n4680), .D(n4728), .Y(n4729));
  NAND2X1 g3639(.A(n4729), .B(n4674), .Y(n4730));
  NOR2X1  g3640(.A(n4730), .B(n4679), .Y(n4731));
  NAND3X1 g3641(.A(n2041), .B(n1987), .C(n1875), .Y(n4732));
  AOI21X1 g3642(.A0(n3385), .A1(n3353), .B0(n3382), .Y(n4733));
  AOI21X1 g3643(.A0(n3385), .A1(n3398), .B0(n4733), .Y(n4734));
  NOR2X1  g3644(.A(n3345), .B(n3329), .Y(n4735));
  NAND2X1 g3645(.A(n4735), .B(n4734), .Y(n4736));
  NOR3X1  g3646(.A(n3198), .B(n2005), .C(n1746), .Y(n4738));
  AOI22X1 g3647(.A0(n3158), .A1(n3179), .B0(n3151), .B1(n3117), .Y(n4741));
  NOR2X1  g3648(.A(n4741), .B(n3209), .Y(n4742));
  NOR2X1  g3649(.A(n3111), .B(n3072), .Y(n4744));
  NAND2X1 g3650(.A(n4744), .B(n3168), .Y(n4745));
  OAI22X1 g3651(.A0(n3035), .A1(n3042), .B0(n3000), .B1(n2993), .Y(n4747));
  NOR2X1  g3652(.A(n3003), .B(n4747), .Y(n4749));
  NAND2X1 g3653(.A(n3042), .B(n3035), .Y(n4752));
  OAI21X1 g3654(.A0(n3044), .A1(n3090), .B0(n4752), .Y(n4753));
  NOR3X1  g3655(.A(n4753), .B(n4749), .C(n3089), .Y(n4754));
  AOI22X1 g3656(.A0(n2906), .A1(n2914), .B0(n2898), .B1(n2864), .Y(n4755));
  NAND2X1 g3657(.A(n2833), .B(n4755), .Y(n4757));
  OAI22X1 g3658(.A0(n2949), .A1(n2956), .B0(n2914), .B1(n2906), .Y(n4760));
  AOI21X1 g3659(.A0(n4718), .A1(n2959), .B0(n4760), .Y(n4761));
  NAND2X1 g3660(.A(n4761), .B(n4757), .Y(n4762));
  NOR2X1  g3661(.A(n4762), .B(n4747), .Y(n4763));
  INVX1   g3662(.A(n2553), .Y(n4767));
  NAND2X1 g3663(.A(n2469), .B(n2454), .Y(n4768));
  NOR2X1  g3664(.A(n2445), .B(n2410), .Y(n4770));
  NAND2X1 g3665(.A(n2279), .B(n2263), .Y(n4771));
  OAI22X1 g3666(.A0(n2365), .A1(n2379), .B0(n2332), .B1(n2316), .Y(n4772));
  NAND3X1 g3667(.A(n2222), .B(n2207), .C(n2202), .Y(n4774));
  OAI21X1 g3668(.A0(n2240), .A1(n2294), .B0(n4774), .Y(n4777));
  AOI21X1 g3669(.A0(n4777), .A1(n4689), .B0(n4772), .Y(n4778));
  NAND2X1 g3670(.A(n4778), .B(n4771), .Y(n4779));
  NOR2X1  g3671(.A(n2425), .B(n2411), .Y(n4780));
  NAND2X1 g3672(.A(n2379), .B(n2365), .Y(n4782));
  OAI21X1 g3673(.A0(n2342), .A1(n2435), .B0(n4782), .Y(n4784));
  NOR2X1  g3674(.A(n4784), .B(n4780), .Y(n4785));
  AOI21X1 g3675(.A0(n4785), .A1(n4779), .B0(n4770), .Y(n4786));
  OAI21X1 g3676(.A0(n4786), .A1(n2527), .B0(n4768), .Y(n4787));
  NAND3X1 g3677(.A(n2385), .B(n2364), .C(n2358), .Y(n4788));
  NAND2X1 g3678(.A(n2341), .B(n4788), .Y(n4790));
  AOI22X1 g3679(.A0(n2208), .A1(n2223), .B0(n2173), .B1(n2167), .Y(n4791));
  NAND3X1 g3680(.A(n4791), .B(n4790), .C(n4782), .Y(n4792));
  OAI21X1 g3681(.A0(n4689), .A1(n4772), .B0(n4767), .Y(n4793));
  NOR4X1  g3682(.A(n4792), .B(n4780), .C(n2527), .D(n4793), .Y(n4794));
  AOI21X1 g3683(.A0(n2033), .A1(n2081), .B0(n2076), .Y(n4796));
  OAI22X1 g3684(.A0(n2111), .A1(n2122), .B0(n2081), .B1(n2033), .Y(n4799));
  NOR2X1  g3685(.A(n4799), .B(n4796), .Y(n4800));
  NAND2X1 g3686(.A(n4800), .B(n4794), .Y(n4801));
  NAND3X1 g3687(.A(n4794), .B(n2111), .C(n2122), .Y(n4802));
  AOI22X1 g3688(.A0(n2635), .A1(n2649), .B0(n2607), .B1(n2594), .Y(n4803));
  AOI22X1 g3689(.A0(n2546), .A1(n2562), .B0(n2511), .B1(n2499), .Y(n4804));
  NAND4X1 g3690(.A(n4803), .B(n4802), .C(n4801), .D(n4804), .Y(n4805));
  AOI21X1 g3691(.A0(n4787), .A1(n4767), .B0(n4805), .Y(n4806));
  NAND2X1 g3692(.A(n2564), .B(n4803), .Y(n4808));
  NAND2X1 g3693(.A(n2649), .B(n2635), .Y(n4809));
  NAND2X1 g3694(.A(n2662), .B(n4809), .Y(n4811));
  AOI22X1 g3695(.A0(n2681), .A1(n2693), .B0(n2653), .B1(n2634), .Y(n4812));
  NAND3X1 g3696(.A(n4812), .B(n4811), .C(n4808), .Y(n4813));
  OAI21X1 g3697(.A0(n4813), .A1(n4806), .B0(n2740), .Y(n4814));
  NAND2X1 g3698(.A(n2737), .B(n2727), .Y(n4815));
  AOI21X1 g3699(.A0(n4815), .A1(n4814), .B0(n2774), .Y(n4816));
  NOR2X1  g3700(.A(n2784), .B(n2765), .Y(n4817));
  NOR2X1  g3701(.A(n4817), .B(n4816), .Y(n4818));
  AOI22X1 g3702(.A0(n2812), .A1(n2825), .B0(n2784), .B1(n2765), .Y(n4819));
  NAND2X1 g3703(.A(n4819), .B(n4755), .Y(n4820));
  OAI21X1 g3704(.A0(n4820), .A1(n4818), .B0(n4763), .Y(n4821));
  NAND3X1 g3705(.A(n4821), .B(n4754), .C(n3168), .Y(n4822));
  AOI21X1 g3706(.A0(n4822), .A1(n4745), .B0(n3209), .Y(n4823));
  NOR3X1  g3707(.A(n4823), .B(n4742), .C(n3250), .Y(n4824));
  NAND2X1 g3708(.A(n3281), .B(n3243), .Y(n4825));
  OAI21X1 g3709(.A0(n4824), .A1(n4738), .B0(n4825), .Y(n4826));
  AOI22X1 g3710(.A0(n3253), .A1(n3255), .B0(n2101), .B1(n3323), .Y(n4827));
  AOI21X1 g3711(.A0(n4827), .A1(n4826), .B0(n3289), .Y(n4828));
  AOI21X1 g3712(.A0(n3301), .A1(n4826), .B0(n3324), .Y(n4831));
  NOR3X1  g3713(.A(n4831), .B(n4672), .C(n4828), .Y(n4832));
  NAND4X1 g3714(.A(n3385), .B(n3382), .C(n3353), .D(n3396), .Y(n4833));
  NAND4X1 g3715(.A(n1993), .B(n2027), .C(n1875), .D(n3472), .Y(n4834));
  AOI21X1 g3716(.A0(n4360), .A1(n3396), .B0(n4834), .Y(n4835));
  NAND2X1 g3717(.A(n4835), .B(n4833), .Y(n4836));
  AOI21X1 g3718(.A0(n4832), .A1(n4734), .B0(n4836), .Y(n4837));
  NOR2X1  g3719(.A(n1984), .B(n1874), .Y(n4838));
  NOR3X1  g3720(.A(n1994), .B(n1989), .C(n1984), .Y(n4839));
  AOI21X1 g3721(.A0(n4839), .A1(n3825), .B0(n1875), .Y(n4840));
  NOR4X1  g3722(.A(n4838), .B(n3916), .C(P1_U3084), .D(n4840), .Y(n4841));
  NOR2X1  g3723(.A(n4841), .B(n1885), .Y(n4842));
  AOI21X1 g3724(.A0(n4837), .A1(n4736), .B0(n4842), .Y(n4843));
  OAI21X1 g3725(.A0(n4732), .A1(n4731), .B0(n4843), .Y(n4844));
  NAND3X1 g3726(.A(n4655), .B(n4441), .C(n4437), .Y(n4845));
  NAND3X1 g3727(.A(n4839), .B(n3825), .C(n1893), .Y(n4846));
  NOR2X1  g3728(.A(n4846), .B(n4845), .Y(n4847));
  NAND2X1 g3729(.A(n4441), .B(n4437), .Y(n4848));
  AOI21X1 g3730(.A0(n4401), .A1(n3328), .B0(n1874), .Y(n4849));
  OAI21X1 g3731(.A0(n3372), .A1(n4405), .B0(n4849), .Y(n4850));
  NAND3X1 g3732(.A(n4850), .B(n4416), .C(n4413), .Y(n4851));
  AOI21X1 g3733(.A0(n4851), .A1(n4651), .B0(n4442), .Y(n4852));
  NOR4X1  g3734(.A(n4650), .B(n4463), .C(n4848), .D(n4852), .Y(n4853));
  NAND2X1 g3735(.A(n4671), .B(n4670), .Y(n4854));
  NAND4X1 g3736(.A(n4676), .B(n4673), .C(n4854), .D(n4677), .Y(n4855));
  NAND3X1 g3737(.A(n4729), .B(n4855), .C(n4674), .Y(n4856));
  NAND2X1 g3738(.A(n4838), .B(n2038), .Y(n4857));
  NAND3X1 g3739(.A(n1993), .B(n1987), .C(n1875), .Y(n4858));
  OAI22X1 g3740(.A0(n4857), .A1(n4853), .B0(n4856), .B1(n4858), .Y(n4859));
  NOR4X1  g3741(.A(n4847), .B(n4844), .C(n4658), .D(n4859), .Y(n4860));
  NOR2X1  g3742(.A(P1_STATE_REG_SCAN_IN), .B(P1_B_REG_SCAN_IN), .Y(n4861));
  NOR2X1  g3743(.A(n4861), .B(n4860), .Y(P1_U3240));
  AOI22X1 g3744(.A0(n4209), .A1(n2681), .B0(n2718), .B1(n4217), .Y(n4863));
  OAI22X1 g3745(.A0(n4211), .A1(n2682), .B0(n2693), .B1(n4216), .Y(n4864));
  XOR2X1  g3746(.A(n4864), .B(n4207), .Y(n4865));
  NOR2X1  g3747(.A(n4865), .B(n4863), .Y(n4866));
  NAND2X1 g3748(.A(n4865), .B(n4863), .Y(n4867));
  INVX1   g3749(.A(n2067), .Y(n4868));
  NOR2X1  g3750(.A(n2065), .B(n2038), .Y(n4869));
  AOI21X1 g3751(.A0(n4869), .A1(n2048), .B0(n1884), .Y(n4870));
  NOR2X1  g3752(.A(n4205), .B(n1884), .Y(n4871));
  NOR2X1  g3753(.A(n4871), .B(n4870), .Y(n4872));
  OAI21X1 g3754(.A0(n4868), .A1(n1884), .B0(n4872), .Y(n4873));
  AOI22X1 g3755(.A0(n4217), .A1(n2634), .B0(n2649), .B1(n4873), .Y(n4874));
  XOR2X1  g3756(.A(n4874), .B(n4215), .Y(n4875));
  AOI22X1 g3757(.A0(n4209), .A1(n2634), .B0(n2649), .B1(n4217), .Y(n4876));
  NAND2X1 g3758(.A(n4876), .B(n4875), .Y(n4877));
  INVX1   g3759(.A(n4877), .Y(n4878));
  AOI22X1 g3760(.A0(n4209), .A1(n2545), .B0(n2562), .B1(n4217), .Y(n4879));
  AOI22X1 g3761(.A0(n4217), .A1(n2545), .B0(n2562), .B1(n4873), .Y(n4880));
  XOR2X1  g3762(.A(n4880), .B(n4215), .Y(n4881));
  NOR2X1  g3763(.A(n4881), .B(n4879), .Y(n4882));
  AOI22X1 g3764(.A0(n4209), .A1(n2593), .B0(n2607), .B1(n4217), .Y(n4883));
  AOI22X1 g3765(.A0(n4217), .A1(n2593), .B0(n2607), .B1(n4873), .Y(n4884));
  XOR2X1  g3766(.A(n4884), .B(n4215), .Y(n4885));
  AOI22X1 g3767(.A0(n4883), .A1(n4885), .B0(n4876), .B1(n4875), .Y(n4886));
  OAI22X1 g3768(.A0(n4883), .A1(n4885), .B0(n4876), .B1(n4875), .Y(n4887));
  AOI21X1 g3769(.A0(n4886), .A1(n4882), .B0(n4887), .Y(n4888));
  AOI22X1 g3770(.A0(n4209), .A1(n2498), .B0(n2511), .B1(n4217), .Y(n4889));
  AOI22X1 g3771(.A0(n4217), .A1(n2498), .B0(n2511), .B1(n4873), .Y(n4890));
  XOR2X1  g3772(.A(n4890), .B(n4215), .Y(n4891));
  NOR2X1  g3773(.A(n4891), .B(n4889), .Y(n4892));
  NAND2X1 g3774(.A(n4891), .B(n4889), .Y(n4893));
  AOI22X1 g3775(.A0(n4217), .A1(n2453), .B0(n2469), .B1(n4873), .Y(n4894));
  XOR2X1  g3776(.A(n4894), .B(n4215), .Y(n4895));
  INVX1   g3777(.A(n4895), .Y(n4896));
  AOI22X1 g3778(.A0(n4209), .A1(n2453), .B0(n2469), .B1(n4217), .Y(n4897));
  INVX1   g3779(.A(n4897), .Y(n4898));
  NOR2X1  g3780(.A(n4898), .B(n4896), .Y(n4899));
  AOI22X1 g3781(.A0(n4209), .A1(n2410), .B0(n2425), .B1(n4217), .Y(n4900));
  AOI22X1 g3782(.A0(n4217), .A1(n2410), .B0(n2425), .B1(n4873), .Y(n4901));
  XOR2X1  g3783(.A(n4901), .B(n4215), .Y(n4902));
  NOR2X1  g3784(.A(n4902), .B(n4900), .Y(n4903));
  NAND2X1 g3785(.A(n4902), .B(n4900), .Y(n4904));
  AOI22X1 g3786(.A0(n4209), .A1(n2316), .B0(n2340), .B1(n4217), .Y(n4905));
  AOI22X1 g3787(.A0(n4217), .A1(n2316), .B0(n2340), .B1(n4873), .Y(n4906));
  XOR2X1  g3788(.A(n4906), .B(n4215), .Y(n4907));
  AOI22X1 g3789(.A0(n4209), .A1(n2365), .B0(n2385), .B1(n4217), .Y(n4908));
  AOI22X1 g3790(.A0(n4217), .A1(n2365), .B0(n2385), .B1(n4873), .Y(n4909));
  XOR2X1  g3791(.A(n4909), .B(n4215), .Y(n4910));
  AOI22X1 g3792(.A0(n4908), .A1(n4910), .B0(n4907), .B1(n4905), .Y(n4911));
  INVX1   g3793(.A(n4911), .Y(n4912));
  AOI22X1 g3794(.A0(n4209), .A1(n2274), .B0(n2279), .B1(n4217), .Y(n4913));
  AOI22X1 g3795(.A0(n4217), .A1(n2274), .B0(n2279), .B1(n4873), .Y(n4914));
  XOR2X1  g3796(.A(n4914), .B(n4215), .Y(n4915));
  NOR2X1  g3797(.A(n4915), .B(n4913), .Y(n4916));
  NAND2X1 g3798(.A(n4915), .B(n4913), .Y(n4917));
  AOI22X1 g3799(.A0(n4217), .A1(n2208), .B0(n2222), .B1(n4873), .Y(n4918));
  XOR2X1  g3800(.A(n4918), .B(n4215), .Y(n4919));
  AOI22X1 g3801(.A0(n4209), .A1(n2208), .B0(n2222), .B1(n4217), .Y(n4920));
  NAND2X1 g3802(.A(n4920), .B(n4919), .Y(n4921));
  INVX1   g3803(.A(n4921), .Y(n4922));
  AOI22X1 g3804(.A0(n4209), .A1(n2110), .B0(n2122), .B1(n4217), .Y(n4923));
  AOI22X1 g3805(.A0(n4217), .A1(n2110), .B0(n2122), .B1(n4873), .Y(n4924));
  XOR2X1  g3806(.A(n4924), .B(n4215), .Y(n4925));
  AOI22X1 g3807(.A0(n4209), .A1(n2167), .B0(n2172), .B1(n4217), .Y(n4926));
  AOI22X1 g3808(.A0(n4217), .A1(n2167), .B0(n2172), .B1(n4873), .Y(n4927));
  XOR2X1  g3809(.A(n4927), .B(n4215), .Y(n4928));
  AOI22X1 g3810(.A0(n4926), .A1(n4928), .B0(n4925), .B1(n4923), .Y(n4929));
  AOI22X1 g3811(.A0(n4209), .A1(n2062), .B0(n2081), .B1(n4217), .Y(n4930));
  INVX1   g3812(.A(n4930), .Y(n4931));
  AOI22X1 g3813(.A0(n4217), .A1(n2062), .B0(n2081), .B1(n4873), .Y(n4932));
  XOR2X1  g3814(.A(n4932), .B(n4207), .Y(n4933));
  NAND2X1 g3815(.A(n4933), .B(n4931), .Y(n4934));
  NOR2X1  g3816(.A(n4933), .B(n4931), .Y(n4935));
  NOR2X1  g3817(.A(n4213), .B(n4207), .Y(n4936));
  NAND2X1 g3818(.A(n4213), .B(n4207), .Y(n4937));
  AOI21X1 g3819(.A0(n4937), .A1(n4220), .B0(n4936), .Y(n4938));
  OAI21X1 g3820(.A0(n4938), .A1(n4935), .B0(n4934), .Y(n4939));
  INVX1   g3821(.A(n4923), .Y(n4940));
  XOR2X1  g3822(.A(n4924), .B(n4207), .Y(n4941));
  INVX1   g3823(.A(n4926), .Y(n4942));
  NAND3X1 g3824(.A(n4942), .B(n4941), .C(n4940), .Y(n4943));
  AOI21X1 g3825(.A0(n4941), .A1(n4940), .B0(n4942), .Y(n4944));
  OAI21X1 g3826(.A0(n4944), .A1(n4928), .B0(n4943), .Y(n4945));
  AOI21X1 g3827(.A0(n4939), .A1(n4929), .B0(n4945), .Y(n4946));
  NOR2X1  g3828(.A(n4920), .B(n4919), .Y(n4947));
  INVX1   g3829(.A(n4947), .Y(n4948));
  OAI21X1 g3830(.A0(n4946), .A1(n4922), .B0(n4948), .Y(n4949));
  AOI21X1 g3831(.A0(n4949), .A1(n4917), .B0(n4916), .Y(n4950));
  NOR2X1  g3832(.A(n4907), .B(n4905), .Y(n4951));
  INVX1   g3833(.A(n4951), .Y(n4952));
  INVX1   g3834(.A(n4908), .Y(n4953));
  INVX1   g3835(.A(n4910), .Y(n4954));
  OAI21X1 g3836(.A0(n4951), .A1(n4953), .B0(n4954), .Y(n4955));
  OAI21X1 g3837(.A0(n4952), .A1(n4908), .B0(n4955), .Y(n4956));
  INVX1   g3838(.A(n4956), .Y(n4957));
  OAI21X1 g3839(.A0(n4950), .A1(n4912), .B0(n4957), .Y(n4958));
  AOI21X1 g3840(.A0(n4958), .A1(n4904), .B0(n4903), .Y(n4959));
  NOR2X1  g3841(.A(n4897), .B(n4895), .Y(n4960));
  INVX1   g3842(.A(n4960), .Y(n4961));
  OAI21X1 g3843(.A0(n4959), .A1(n4899), .B0(n4961), .Y(n4962));
  AOI21X1 g3844(.A0(n4962), .A1(n4893), .B0(n4892), .Y(n4963));
  NAND2X1 g3845(.A(n4885), .B(n4883), .Y(n4964));
  INVX1   g3846(.A(n4964), .Y(n4965));
  NAND2X1 g3847(.A(n4881), .B(n4879), .Y(n4966));
  INVX1   g3848(.A(n4966), .Y(n4967));
  NOR3X1  g3849(.A(n4967), .B(n4965), .C(n4878), .Y(n4968));
  INVX1   g3850(.A(n4968), .Y(n4969));
  OAI22X1 g3851(.A0(n4963), .A1(n4969), .B0(n4888), .B1(n4878), .Y(n4970));
  AOI21X1 g3852(.A0(n4970), .A1(n4867), .B0(n4866), .Y(n4971));
  OAI22X1 g3853(.A0(n4211), .A1(n2726), .B0(n2737), .B1(n4216), .Y(n4972));
  XOR2X1  g3854(.A(n4972), .B(n4207), .Y(n4973));
  AOI22X1 g3855(.A0(n4209), .A1(n2727), .B0(n2757), .B1(n4217), .Y(n4974));
  XOR2X1  g3856(.A(n4974), .B(n4973), .Y(n4975));
  XOR2X1  g3857(.A(n4975), .B(n4971), .Y(n4976));
  NOR3X1  g3858(.A(n1999), .B(n1982), .C(n1980), .Y(n4977));
  OAI21X1 g3859(.A0(n2041), .A1(n2027), .B0(n1985), .Y(n4978));
  OAI21X1 g3860(.A0(n2041), .A1(n2027), .B0(n1991), .Y(n4979));
  NOR2X1  g3861(.A(n4979), .B(n1985), .Y(n4980));
  NOR4X1  g3862(.A(n3488), .B(n2049), .C(n2047), .D(n4980), .Y(n4981));
  OAI21X1 g3863(.A0(n4978), .A1(n1991), .B0(n4981), .Y(n4982));
  NAND3X1 g3864(.A(n4982), .B(n4977), .C(n1893), .Y(n4983));
  INVX1   g3865(.A(n4977), .Y(n4984));
  NOR4X1  g3866(.A(n1884), .B(n1875), .C(P1_U3084), .D(n3484), .Y(n4985));
  NAND3X1 g3867(.A(n3475), .B(n3915), .C(n1874), .Y(n4986));
  AOI21X1 g3868(.A0(n4982), .A1(n4984), .B0(n4986), .Y(n4987));
  NOR2X1  g3869(.A(n4987), .B(P1_U3084), .Y(n4988));
  AOI21X1 g3870(.A0(n4985), .A1(n4984), .B0(n4988), .Y(n4989));
  NOR4X1  g3871(.A(n1989), .B(n1984), .C(n1894), .D(n1994), .Y(n4991));
  INVX1   g3872(.A(n4991), .Y(n4992));
  NOR4X1  g3873(.A(n1999), .B(n1982), .C(n1980), .D(n2092), .Y(n4993));
  NOR4X1  g3874(.A(n1999), .B(n1982), .C(n1980), .D(n3910), .Y(n4994));
  INVX1   g3875(.A(n4994), .Y(n4995));
  OAI22X1 g3876(.A0(n4977), .A1(n2721), .B0(n2765), .B1(n4995), .Y(n4996));
  AOI21X1 g3877(.A0(n4993), .A1(n2681), .B0(n4996), .Y(n4997));
  AOI22X1 g3878(.A0(n4977), .A1(n4985), .B0(n3469), .B1(n1893), .Y(n4998));
  AOI22X1 g3879(.A0(n2757), .A1(n5145), .B0(P1_U3084), .B1(P1_REG3_REG_15__SCAN_IN), .Y(n5000));
  OAI21X1 g3880(.A0(n4997), .A1(n4992), .B0(n5000), .Y(n5001));
  AOI21X1 g3881(.A0(n5152), .A1(n2722), .B0(n5001), .Y(n5002));
  OAI21X1 g3882(.A0(n4983), .A1(n4976), .B0(n5002), .Y(P1_U3239));
  AOI22X1 g3883(.A0(n4209), .A1(n3117), .B0(n3124), .B1(n4217), .Y(n5004));
  INVX1   g3884(.A(n5004), .Y(n5005));
  AOI22X1 g3885(.A0(n4217), .A1(n3117), .B0(n3124), .B1(n4873), .Y(n5006));
  XOR2X1  g3886(.A(n5006), .B(n4207), .Y(n5007));
  NOR2X1  g3887(.A(n5007), .B(n5005), .Y(n5008));
  AOI22X1 g3888(.A0(n4209), .A1(n3071), .B0(n3111), .B1(n4217), .Y(n5009));
  OAI22X1 g3889(.A0(n4211), .A1(n3072), .B0(n3085), .B1(n4216), .Y(n5010));
  XOR2X1  g3890(.A(n5010), .B(n4207), .Y(n5011));
  NOR2X1  g3891(.A(n5011), .B(n5009), .Y(n5012));
  NAND2X1 g3892(.A(n5011), .B(n5009), .Y(n5013));
  AOI22X1 g3893(.A0(n4209), .A1(n3080), .B0(n3042), .B1(n4217), .Y(n5014));
  AOI22X1 g3894(.A0(n4217), .A1(n3080), .B0(n3042), .B1(n4873), .Y(n5015));
  XOR2X1  g3895(.A(n5015), .B(n4215), .Y(n5016));
  NOR2X1  g3896(.A(n5016), .B(n5014), .Y(n5017));
  INVX1   g3897(.A(n5017), .Y(n5018));
  NAND2X1 g3898(.A(n5016), .B(n5014), .Y(n5019));
  INVX1   g3899(.A(n5019), .Y(n5020));
  AOI22X1 g3900(.A0(n4217), .A1(n2994), .B0(n3000), .B1(n4873), .Y(n5021));
  XOR2X1  g3901(.A(n5021), .B(n4215), .Y(n5022));
  AOI22X1 g3902(.A0(n4209), .A1(n2994), .B0(n3000), .B1(n4217), .Y(n5023));
  NAND2X1 g3903(.A(n5023), .B(n5022), .Y(n5024));
  AOI22X1 g3904(.A0(n4209), .A1(n2926), .B0(n2914), .B1(n4217), .Y(n5025));
  AOI22X1 g3905(.A0(n4217), .A1(n2926), .B0(n2914), .B1(n4873), .Y(n5026));
  XOR2X1  g3906(.A(n5026), .B(n4215), .Y(n5027));
  NOR2X1  g3907(.A(n5027), .B(n5025), .Y(n5028));
  INVX1   g3908(.A(n5028), .Y(n5029));
  AOI22X1 g3909(.A0(n4209), .A1(n2948), .B0(n2956), .B1(n4217), .Y(n5030));
  AOI22X1 g3910(.A0(n4217), .A1(n2948), .B0(n2956), .B1(n4873), .Y(n5031));
  XOR2X1  g3911(.A(n5031), .B(n4215), .Y(n5032));
  NAND2X1 g3912(.A(n5032), .B(n5030), .Y(n5033));
  NAND2X1 g3913(.A(n5033), .B(n5024), .Y(n5034));
  INVX1   g3914(.A(n5022), .Y(n5035));
  INVX1   g3915(.A(n5023), .Y(n5036));
  NOR2X1  g3916(.A(n5032), .B(n5030), .Y(n5037));
  AOI21X1 g3917(.A0(n5036), .A1(n5035), .B0(n5037), .Y(n5038));
  OAI21X1 g3918(.A0(n5034), .A1(n5029), .B0(n5038), .Y(n5039));
  AOI22X1 g3919(.A0(n4209), .A1(n2863), .B0(n2898), .B1(n4217), .Y(n5040));
  OAI22X1 g3920(.A0(n4211), .A1(n2864), .B0(n2880), .B1(n4216), .Y(n5041));
  XOR2X1  g3921(.A(n5041), .B(n4207), .Y(n5042));
  NOR2X1  g3922(.A(n5042), .B(n5040), .Y(n5043));
  INVX1   g3923(.A(n5043), .Y(n5044));
  NAND2X1 g3924(.A(n5042), .B(n5040), .Y(n5045));
  INVX1   g3925(.A(n5045), .Y(n5046));
  AOI22X1 g3926(.A0(n4209), .A1(n2764), .B0(n2784), .B1(n4217), .Y(n5047));
  OAI22X1 g3927(.A0(n4211), .A1(n2765), .B0(n2779), .B1(n4216), .Y(n5048));
  XOR2X1  g3928(.A(n5048), .B(n4207), .Y(n5049));
  AOI22X1 g3929(.A0(n4209), .A1(n2811), .B0(n2825), .B1(n4217), .Y(n5050));
  AOI22X1 g3930(.A0(n4217), .A1(n2811), .B0(n2825), .B1(n4873), .Y(n5051));
  XOR2X1  g3931(.A(n5051), .B(n4215), .Y(n5052));
  AOI22X1 g3932(.A0(n5050), .A1(n5052), .B0(n5049), .B1(n5047), .Y(n5053));
  NOR2X1  g3933(.A(n4974), .B(n4973), .Y(n5054));
  INVX1   g3934(.A(n5054), .Y(n5055));
  NAND2X1 g3935(.A(n4974), .B(n4973), .Y(n5056));
  INVX1   g3936(.A(n5056), .Y(n5057));
  OAI21X1 g3937(.A0(n5057), .A1(n4971), .B0(n5055), .Y(n5058));
  NOR3X1  g3938(.A(n5050), .B(n5049), .C(n5047), .Y(n5059));
  NOR2X1  g3939(.A(n5049), .B(n5047), .Y(n5060));
  INVX1   g3940(.A(n5060), .Y(n5061));
  AOI21X1 g3941(.A0(n5061), .A1(n5050), .B0(n5052), .Y(n5062));
  NOR2X1  g3942(.A(n5062), .B(n5059), .Y(n5063));
  INVX1   g3943(.A(n5063), .Y(n5064));
  AOI21X1 g3944(.A0(n5058), .A1(n5053), .B0(n5064), .Y(n5065));
  OAI21X1 g3945(.A0(n5065), .A1(n5046), .B0(n5044), .Y(n5066));
  NAND2X1 g3946(.A(n5027), .B(n5025), .Y(n5067));
  INVX1   g3947(.A(n5067), .Y(n5068));
  NOR2X1  g3948(.A(n5068), .B(n5034), .Y(n5069));
  AOI22X1 g3949(.A0(n5066), .A1(n5069), .B0(n5039), .B1(n5024), .Y(n5070));
  OAI21X1 g3950(.A0(n5070), .A1(n5020), .B0(n5018), .Y(n5071));
  AOI21X1 g3951(.A0(n5071), .A1(n5013), .B0(n5012), .Y(n5072));
  AOI22X1 g3952(.A0(n4209), .A1(n3158), .B0(n3166), .B1(n4217), .Y(n5073));
  INVX1   g3953(.A(n5073), .Y(n5074));
  OAI22X1 g3954(.A0(n4211), .A1(n3159), .B0(n3179), .B1(n4216), .Y(n5075));
  XOR2X1  g3955(.A(n5075), .B(n4207), .Y(n5076));
  INVX1   g3956(.A(n5076), .Y(n5077));
  NAND2X1 g3957(.A(n5007), .B(n5005), .Y(n5078));
  INVX1   g3958(.A(n5078), .Y(n5079));
  AOI21X1 g3959(.A0(n5077), .A1(n5074), .B0(n5079), .Y(n5080));
  OAI21X1 g3960(.A0(n5072), .A1(n5008), .B0(n5080), .Y(n5081));
  OAI22X1 g3961(.A0(n4211), .A1(n3199), .B0(n3266), .B1(n4216), .Y(n5082));
  XOR2X1  g3962(.A(n5082), .B(n4207), .Y(n5083));
  OAI22X1 g3963(.A0(n4872), .A1(n3199), .B0(n3266), .B1(n4211), .Y(n5084));
  INVX1   g3964(.A(n5084), .Y(n5085));
  NOR2X1  g3965(.A(n5085), .B(n5083), .Y(n5086));
  INVX1   g3966(.A(n5086), .Y(n5087));
  AOI22X1 g3967(.A0(n5083), .A1(n5085), .B0(n5076), .B1(n5073), .Y(n5088));
  NAND3X1 g3968(.A(n5088), .B(n5087), .C(n5081), .Y(n5089));
  INVX1   g3969(.A(n5008), .Y(n5090));
  INVX1   g3970(.A(n5012), .Y(n5091));
  INVX1   g3971(.A(n5013), .Y(n5092));
  NAND2X1 g3972(.A(n5039), .B(n5024), .Y(n5093));
  INVX1   g3973(.A(n5053), .Y(n5094));
  INVX1   g3974(.A(n4866), .Y(n5095));
  INVX1   g3975(.A(n4867), .Y(n5096));
  NOR2X1  g3976(.A(n4888), .B(n4878), .Y(n5097));
  INVX1   g3977(.A(n4892), .Y(n5098));
  INVX1   g3978(.A(n4893), .Y(n5099));
  INVX1   g3979(.A(n4899), .Y(n5100));
  INVX1   g3980(.A(n4903), .Y(n5101));
  INVX1   g3981(.A(n4904), .Y(n5102));
  INVX1   g3982(.A(n4916), .Y(n5103));
  INVX1   g3983(.A(n4917), .Y(n5104));
  XOR2X1  g3984(.A(n4927), .B(n4207), .Y(n5105));
  OAI22X1 g3985(.A0(n4942), .A1(n5105), .B0(n4941), .B1(n4940), .Y(n5106));
  XOR2X1  g3986(.A(n4932), .B(n4215), .Y(n5107));
  NOR2X1  g3987(.A(n5107), .B(n4930), .Y(n5108));
  NAND2X1 g3988(.A(n5107), .B(n4930), .Y(n5109));
  XOR2X1  g3989(.A(n4219), .B(n4207), .Y(n5110));
  INVX1   g3990(.A(n4212), .Y(n5111));
  OAI21X1 g3991(.A0(n4872), .A1(n2036), .B0(n5111), .Y(n5112));
  NAND2X1 g3992(.A(n5112), .B(n4215), .Y(n5113));
  NOR2X1  g3993(.A(n5112), .B(n4215), .Y(n5114));
  OAI21X1 g3994(.A0(n5114), .A1(n5110), .B0(n5113), .Y(n5115));
  AOI21X1 g3995(.A0(n5115), .A1(n5109), .B0(n5108), .Y(n5116));
  NOR3X1  g3996(.A(n4926), .B(n4925), .C(n4923), .Y(n5117));
  OAI21X1 g3997(.A0(n4925), .A1(n4923), .B0(n4926), .Y(n5118));
  AOI21X1 g3998(.A0(n5118), .A1(n5105), .B0(n5117), .Y(n5119));
  OAI21X1 g3999(.A0(n5116), .A1(n5106), .B0(n5119), .Y(n5120));
  AOI21X1 g4000(.A0(n5120), .A1(n4921), .B0(n4947), .Y(n5121));
  OAI21X1 g4001(.A0(n5121), .A1(n5104), .B0(n5103), .Y(n5122));
  AOI21X1 g4002(.A0(n5122), .A1(n4911), .B0(n4956), .Y(n5123));
  OAI21X1 g4003(.A0(n5123), .A1(n5102), .B0(n5101), .Y(n5124));
  AOI21X1 g4004(.A0(n5124), .A1(n5100), .B0(n4960), .Y(n5125));
  OAI21X1 g4005(.A0(n5125), .A1(n5099), .B0(n5098), .Y(n5126));
  AOI21X1 g4006(.A0(n4968), .A1(n5126), .B0(n5097), .Y(n5127));
  OAI21X1 g4007(.A0(n5127), .A1(n5096), .B0(n5095), .Y(n5128));
  AOI21X1 g4008(.A0(n5056), .A1(n5128), .B0(n5054), .Y(n5129));
  OAI21X1 g4009(.A0(n5129), .A1(n5094), .B0(n5063), .Y(n5130));
  AOI21X1 g4010(.A0(n5130), .A1(n5045), .B0(n5043), .Y(n5131));
  INVX1   g4011(.A(n5069), .Y(n5132));
  OAI21X1 g4012(.A0(n5132), .A1(n5131), .B0(n5093), .Y(n5133));
  AOI21X1 g4013(.A0(n5133), .A1(n5019), .B0(n5017), .Y(n5134));
  OAI21X1 g4014(.A0(n5134), .A1(n5092), .B0(n5091), .Y(n5135));
  AOI21X1 g4015(.A0(n5135), .A1(n5090), .B0(n5079), .Y(n5136));
  XOR2X1  g4016(.A(n5085), .B(n5083), .Y(n5137));
  AOI21X1 g4017(.A0(n5077), .A1(n5074), .B0(n5137), .Y(n5138));
  INVX1   g4018(.A(n4983), .Y(n5139));
  NAND2X1 g4019(.A(n5076), .B(n5073), .Y(n5140));
  OAI21X1 g4020(.A0(n5137), .A1(n5140), .B0(n5139), .Y(n5141));
  AOI21X1 g4021(.A0(n5138), .A1(n5136), .B0(n5141), .Y(n5142));
  NAND2X1 g4022(.A(n5142), .B(n5089), .Y(n5143));
  NAND4X1 g4023(.A(n3403), .B(n3471), .C(n1979), .D(n3550), .Y(n5144));
  AOI21X1 g4024(.A0(n5144), .A1(n3470), .B0(n1894), .Y(n5145));
  NAND2X1 g4025(.A(n5145), .B(n3206), .Y(n5146));
  NOR2X1  g4026(.A(n4995), .B(n3253), .Y(n5147));
  INVX1   g4027(.A(n4993), .Y(n5148));
  OAI22X1 g4028(.A0(n4977), .A1(n3194), .B0(n3159), .B1(n5148), .Y(n5149));
  OAI21X1 g4029(.A0(n5149), .A1(n5147), .B0(n4991), .Y(n5150));
  NAND2X1 g4030(.A(n4984), .B(n3550), .Y(n5151));
  AOI21X1 g4031(.A0(n5151), .A1(n4987), .B0(P1_U3084), .Y(n5152));
  AOI22X1 g4032(.A0(n3690), .A1(n5152), .B0(P1_U3084), .B1(P1_REG3_REG_26__SCAN_IN), .Y(n5153));
  NAND4X1 g4033(.A(n5150), .B(n5146), .C(n5143), .D(n5153), .Y(P1_U3238));
  INVX1   g4034(.A(n4905), .Y(n5155));
  XOR2X1  g4035(.A(n4907), .B(n5155), .Y(n5156));
  NOR2X1  g4036(.A(n5156), .B(n5122), .Y(n5157));
  XOR2X1  g4037(.A(n4907), .B(n4905), .Y(n5158));
  NOR2X1  g4038(.A(n5158), .B(n4950), .Y(n5159));
  OAI21X1 g4039(.A0(n5159), .A1(n5157), .B0(n5139), .Y(n5160));
  NOR2X1  g4040(.A(n4989), .B(n2313), .Y(n5161));
  OAI22X1 g4041(.A0(n4977), .A1(n2313), .B0(n2263), .B1(n5148), .Y(n5162));
  AOI21X1 g4042(.A0(n4994), .A1(n2365), .B0(n5162), .Y(n5163));
  AOI22X1 g4043(.A0(n2340), .A1(n5145), .B0(P1_U3084), .B1(P1_REG3_REG_6__SCAN_IN), .Y(n5164));
  OAI21X1 g4044(.A0(n5163), .A1(n4992), .B0(n5164), .Y(n5165));
  NOR2X1  g4045(.A(n5165), .B(n5161), .Y(n5166));
  NAND2X1 g4046(.A(n5166), .B(n5160), .Y(P1_U3237));
  XOR2X1  g4047(.A(n5042), .B(n5040), .Y(n5168));
  XOR2X1  g4048(.A(n5168), .B(n5065), .Y(n5169));
  AOI22X1 g4049(.A0(n4984), .A1(n2859), .B0(n2926), .B1(n4994), .Y(n5170));
  OAI21X1 g4050(.A0(n5148), .A1(n2812), .B0(n5170), .Y(n5171));
  AOI22X1 g4051(.A0(n4991), .A1(n5171), .B0(P1_U3084), .B1(P1_REG3_REG_18__SCAN_IN), .Y(n5172));
  OAI21X1 g4052(.A0(n4989), .A1(n2858), .B0(n5172), .Y(n5173));
  AOI21X1 g4053(.A0(n5145), .A1(n2898), .B0(n5173), .Y(n5174));
  OAI21X1 g4054(.A0(n5169), .A1(n4983), .B0(n5174), .Y(P1_U3236));
  XOR2X1  g4055(.A(n4941), .B(n4923), .Y(n5176));
  NOR2X1  g4056(.A(n4941), .B(n4940), .Y(n5177));
  NOR2X1  g4057(.A(n4925), .B(n4923), .Y(n5178));
  OAI21X1 g4058(.A0(n5178), .A1(n5177), .B0(n4939), .Y(n5179));
  OAI21X1 g4059(.A0(n5176), .A1(n4939), .B0(n5179), .Y(n5180));
  NAND2X1 g4060(.A(n5180), .B(n5139), .Y(n5181));
  INVX1   g4061(.A(P1_REG3_REG_2__SCAN_IN), .Y(n5182));
  OAI22X1 g4062(.A0(n4977), .A1(n5182), .B0(n2076), .B1(n5148), .Y(n5183));
  AOI21X1 g4063(.A0(n4994), .A1(n2167), .B0(n5183), .Y(n5184));
  AOI22X1 g4064(.A0(n2122), .A1(n5145), .B0(P1_U3084), .B1(P1_REG3_REG_2__SCAN_IN), .Y(n5185));
  OAI21X1 g4065(.A0(n5184), .A1(n4992), .B0(n5185), .Y(n5186));
  AOI21X1 g4066(.A0(n5152), .A1(P1_REG3_REG_2__SCAN_IN), .B0(n5186), .Y(n5187));
  NAND2X1 g4067(.A(n5187), .B(n5181), .Y(P1_U3235));
  INVX1   g4068(.A(n4879), .Y(n5189));
  XOR2X1  g4069(.A(n4881), .B(n5189), .Y(n5190));
  OAI21X1 g4070(.A0(n4967), .A1(n4882), .B0(n5126), .Y(n5191));
  OAI21X1 g4071(.A0(n5190), .A1(n5126), .B0(n5191), .Y(n5192));
  NAND2X1 g4072(.A(n5192), .B(n5139), .Y(n5193));
  OAI22X1 g4073(.A0(n4977), .A1(n2540), .B0(n2499), .B1(n5148), .Y(n5194));
  AOI21X1 g4074(.A0(n4994), .A1(n2593), .B0(n5194), .Y(n5195));
  AOI22X1 g4075(.A0(n2562), .A1(n5145), .B0(P1_U3084), .B1(P1_REG3_REG_11__SCAN_IN), .Y(n5196));
  OAI21X1 g4076(.A0(n5195), .A1(n4992), .B0(n5196), .Y(n5197));
  AOI21X1 g4077(.A0(n5152), .A1(n2541), .B0(n5197), .Y(n5198));
  NAND2X1 g4078(.A(n5198), .B(n5193), .Y(P1_U3234));
  XOR2X1  g4079(.A(n5016), .B(n5014), .Y(n5200));
  XOR2X1  g4080(.A(n5200), .B(n5070), .Y(n5201));
  NAND2X1 g4081(.A(n5152), .B(n3031), .Y(n5202));
  AOI22X1 g4082(.A0(n4984), .A1(n3031), .B0(n2994), .B1(n4993), .Y(n5203));
  OAI21X1 g4083(.A0(n4995), .A1(n3072), .B0(n5203), .Y(n5204));
  AOI22X1 g4084(.A0(n4991), .A1(n5204), .B0(P1_U3084), .B1(P1_REG3_REG_22__SCAN_IN), .Y(n5205));
  NAND2X1 g4085(.A(n5205), .B(n5202), .Y(n5206));
  AOI21X1 g4086(.A0(n5145), .A1(n3042), .B0(n5206), .Y(n5207));
  OAI21X1 g4087(.A0(n5201), .A1(n4983), .B0(n5207), .Y(P1_U3233));
  NOR2X1  g4088(.A(n4885), .B(n4883), .Y(n5209));
  INVX1   g4089(.A(n5209), .Y(n5210));
  AOI21X1 g4090(.A0(n4966), .A1(n5126), .B0(n4882), .Y(n5211));
  OAI21X1 g4091(.A0(n4876), .A1(n4875), .B0(n4886), .Y(n5212));
  AOI21X1 g4092(.A0(n5211), .A1(n5210), .B0(n5212), .Y(n5213));
  INVX1   g4093(.A(n4876), .Y(n5214));
  OAI22X1 g4094(.A0(n4883), .A1(n4885), .B0(n5214), .B1(n4875), .Y(n5215));
  AOI21X1 g4095(.A0(n5214), .A1(n4875), .B0(n5215), .Y(n5216));
  OAI21X1 g4096(.A0(n5211), .A1(n4965), .B0(n5216), .Y(n5217));
  NAND2X1 g4097(.A(n5217), .B(n5139), .Y(n5218));
  OAI22X1 g4098(.A0(n4977), .A1(n2630), .B0(n2682), .B1(n4995), .Y(n5219));
  AOI21X1 g4099(.A0(n4993), .A1(n2593), .B0(n5219), .Y(n5220));
  AOI22X1 g4100(.A0(n2649), .A1(n5145), .B0(P1_U3084), .B1(P1_REG3_REG_13__SCAN_IN), .Y(n5221));
  OAI21X1 g4101(.A0(n5220), .A1(n4992), .B0(n5221), .Y(n5222));
  AOI21X1 g4102(.A0(n5152), .A1(n2631), .B0(n5222), .Y(n5223));
  OAI21X1 g4103(.A0(n5218), .A1(n5213), .B0(n5223), .Y(P1_U3232));
  AOI21X1 g4104(.A0(n5067), .A1(n5066), .B0(n5028), .Y(n5225));
  XOR2X1  g4105(.A(n5032), .B(n5030), .Y(n5226));
  NAND2X1 g4106(.A(n5225), .B(n5226), .Y(n5227));
  OAI21X1 g4107(.A0(n5226), .A1(n5225), .B0(n5227), .Y(n5229));
  NAND2X1 g4108(.A(n5229), .B(n5139), .Y(n5230));
  NAND2X1 g4109(.A(n5145), .B(n2956), .Y(n5231));
  OAI22X1 g4110(.A0(n4977), .A1(n2944), .B0(n2993), .B1(n4995), .Y(n5232));
  AOI21X1 g4111(.A0(n4993), .A1(n2926), .B0(n5232), .Y(n5233));
  OAI22X1 g4112(.A0(n4992), .A1(n5233), .B0(P1_STATE_REG_SCAN_IN), .B1(n2941), .Y(n5234));
  AOI21X1 g4113(.A0(n5152), .A1(n3637), .B0(n5234), .Y(n5235));
  NAND3X1 g4114(.A(n5235), .B(n5231), .C(n5230), .Y(P1_U3231));
  OAI21X1 g4115(.A0(n4991), .A1(n4985), .B0(n4984), .Y(n5237));
  OAI21X1 g4116(.A0(n4987), .A1(P1_U3084), .B0(n5237), .Y(n5238));
  NAND2X1 g4117(.A(n5238), .B(P1_REG3_REG_0__SCAN_IN), .Y(n5239));
  NAND4X1 g4118(.A(n4977), .B(n4221), .C(n1893), .D(n4982), .Y(n5240));
  NAND2X1 g4119(.A(n5145), .B(n2035), .Y(n5241));
  NOR2X1  g4120(.A(n4992), .B(n2076), .Y(n5242));
  AOI22X1 g4121(.A0(n4994), .A1(n5242), .B0(P1_U3084), .B1(P1_REG3_REG_0__SCAN_IN), .Y(n5243));
  NAND4X1 g4122(.A(n5241), .B(n5240), .C(n5239), .D(n5243), .Y(P1_U3230));
  XOR2X1  g4123(.A(n4897), .B(n4895), .Y(n5245));
  XOR2X1  g4124(.A(n5245), .B(n4959), .Y(n5246));
  OAI22X1 g4125(.A0(n4977), .A1(n2449), .B0(n2411), .B1(n5148), .Y(n5247));
  AOI21X1 g4126(.A0(n4994), .A1(n2498), .B0(n5247), .Y(n5248));
  AOI22X1 g4127(.A0(n2469), .A1(n5145), .B0(P1_U3084), .B1(P1_REG3_REG_9__SCAN_IN), .Y(n5249));
  OAI21X1 g4128(.A0(n5248), .A1(n4992), .B0(n5249), .Y(n5250));
  AOI21X1 g4129(.A0(n5152), .A1(n2450), .B0(n5250), .Y(n5251));
  OAI21X1 g4130(.A0(n5246), .A1(n4983), .B0(n5251), .Y(P1_U3229));
  XOR2X1  g4131(.A(n4920), .B(n4919), .Y(n5253));
  XOR2X1  g4132(.A(n5253), .B(n4946), .Y(n5254));
  NOR2X1  g4133(.A(n4989), .B(n2205), .Y(n5255));
  OAI22X1 g4134(.A0(n4977), .A1(n2205), .B0(n2154), .B1(n5148), .Y(n5256));
  AOI21X1 g4135(.A0(n4994), .A1(n2274), .B0(n5256), .Y(n5257));
  AOI22X1 g4136(.A0(n2222), .A1(n5145), .B0(P1_U3084), .B1(P1_REG3_REG_4__SCAN_IN), .Y(n5258));
  OAI21X1 g4137(.A0(n5257), .A1(n4992), .B0(n5258), .Y(n5259));
  NOR2X1  g4138(.A(n5259), .B(n5255), .Y(n5260));
  OAI21X1 g4139(.A0(n5254), .A1(n4983), .B0(n5260), .Y(P1_U3228));
  XOR2X1  g4140(.A(n5007), .B(n5004), .Y(n5262));
  NOR2X1  g4141(.A(n5262), .B(n5135), .Y(n5263));
  AOI21X1 g4142(.A0(n5078), .A1(n5090), .B0(n5072), .Y(n5264));
  OAI21X1 g4143(.A0(n5264), .A1(n5263), .B0(n5139), .Y(n5265));
  NAND2X1 g4144(.A(n5145), .B(n3124), .Y(n5266));
  NOR2X1  g4145(.A(n4995), .B(n3159), .Y(n5267));
  OAI22X1 g4146(.A0(n4977), .A1(n3113), .B0(n3072), .B1(n5148), .Y(n5268));
  OAI21X1 g4147(.A0(n5268), .A1(n5267), .B0(n4991), .Y(n5269));
  AOI22X1 g4148(.A0(n3672), .A1(n5152), .B0(P1_U3084), .B1(P1_REG3_REG_24__SCAN_IN), .Y(n5270));
  NAND4X1 g4149(.A(n5269), .B(n5266), .C(n5265), .D(n5270), .Y(P1_U3227));
  OAI21X1 g4150(.A0(n5052), .A1(n5050), .B0(n5053), .Y(n5272));
  AOI21X1 g4151(.A0(n5061), .A1(n5129), .B0(n5272), .Y(n5273));
  AOI21X1 g4152(.A0(n5049), .A1(n5047), .B0(n5129), .Y(n5274));
  INVX1   g4153(.A(n5052), .Y(n5275));
  AOI21X1 g4154(.A0(n5275), .A1(n5050), .B0(n5060), .Y(n5276));
  OAI21X1 g4155(.A0(n5275), .A1(n5050), .B0(n5276), .Y(n5277));
  OAI21X1 g4156(.A0(n5277), .A1(n5274), .B0(n5139), .Y(n5278));
  AOI22X1 g4157(.A0(n4984), .A1(n2807), .B0(n2863), .B1(n4994), .Y(n5279));
  OAI21X1 g4158(.A0(n5148), .A1(n2765), .B0(n5279), .Y(n5280));
  AOI22X1 g4159(.A0(n4991), .A1(n5280), .B0(P1_U3084), .B1(P1_REG3_REG_17__SCAN_IN), .Y(n5281));
  OAI21X1 g4160(.A0(n4989), .A1(n2806), .B0(n5281), .Y(n5282));
  AOI21X1 g4161(.A0(n5145), .A1(n2825), .B0(n5282), .Y(n5283));
  OAI21X1 g4162(.A0(n5278), .A1(n5273), .B0(n5283), .Y(P1_U3226));
  XOR2X1  g4163(.A(n4915), .B(n4913), .Y(n5285));
  XOR2X1  g4164(.A(n5285), .B(n5121), .Y(n5286));
  NAND2X1 g4165(.A(n4994), .B(n2316), .Y(n5287));
  AOI22X1 g4166(.A0(n4984), .A1(n2260), .B0(n2208), .B1(n4993), .Y(n5288));
  AOI21X1 g4167(.A0(n5288), .A1(n5287), .B0(n4992), .Y(n5289));
  AOI22X1 g4168(.A0(n2279), .A1(n5145), .B0(P1_U3084), .B1(P1_REG3_REG_5__SCAN_IN), .Y(n5290));
  OAI21X1 g4169(.A0(n4989), .A1(n2259), .B0(n5290), .Y(n5291));
  NOR2X1  g4170(.A(n5291), .B(n5289), .Y(n5292));
  OAI21X1 g4171(.A0(n5286), .A1(n4983), .B0(n5292), .Y(P1_U3225));
  INVX1   g4172(.A(n5047), .Y(n5294));
  XOR2X1  g4173(.A(n5049), .B(n5294), .Y(n5295));
  NOR2X1  g4174(.A(n5295), .B(n5058), .Y(n5296));
  XOR2X1  g4175(.A(n5049), .B(n5047), .Y(n5297));
  NOR2X1  g4176(.A(n5297), .B(n5129), .Y(n5298));
  OAI21X1 g4177(.A0(n5298), .A1(n5296), .B0(n5139), .Y(n5299));
  NAND2X1 g4178(.A(n5152), .B(n2760), .Y(n5300));
  AOI22X1 g4179(.A0(n4984), .A1(n2760), .B0(n2811), .B1(n4994), .Y(n5301));
  OAI21X1 g4180(.A0(n5148), .A1(n2726), .B0(n5301), .Y(n5302));
  NAND2X1 g4181(.A(n5302), .B(n4991), .Y(n5303));
  AOI22X1 g4182(.A0(n2784), .A1(n5145), .B0(P1_U3084), .B1(P1_REG3_REG_16__SCAN_IN), .Y(n5304));
  NAND4X1 g4183(.A(n5303), .B(n5300), .C(n5299), .D(n5304), .Y(P1_U3224));
  OAI21X1 g4184(.A0(n5072), .A1(n5008), .B0(n5078), .Y(n5306));
  XOR2X1  g4185(.A(n5076), .B(n5074), .Y(n5307));
  NOR2X1  g4186(.A(n5307), .B(n5306), .Y(n5308));
  XOR2X1  g4187(.A(n5076), .B(n5073), .Y(n5309));
  NOR2X1  g4188(.A(n5309), .B(n5136), .Y(n5310));
  OAI21X1 g4189(.A0(n5310), .A1(n5308), .B0(n5139), .Y(n5311));
  NAND2X1 g4190(.A(n5145), .B(n3166), .Y(n5312));
  AOI22X1 g4191(.A0(n4984), .A1(n3682), .B0(n3117), .B1(n4993), .Y(n5313));
  OAI21X1 g4192(.A0(n4995), .A1(n3199), .B0(n5313), .Y(n5314));
  OAI22X1 g4193(.A0(n3154), .A1(n4989), .B0(P1_STATE_REG_SCAN_IN), .B1(n3192), .Y(n5316));
  AOI21X1 g4194(.A0(n5314), .A1(n4991), .B0(n5316), .Y(n5317));
  NAND3X1 g4195(.A(n5317), .B(n5312), .C(n5311), .Y(P1_U3223));
  NOR2X1  g4196(.A(n4967), .B(n4963), .Y(n5319));
  INVX1   g4197(.A(n4883), .Y(n5320));
  XOR2X1  g4198(.A(n4885), .B(n5320), .Y(n5321));
  NOR3X1  g4199(.A(n5321), .B(n5319), .C(n4882), .Y(n5322));
  AOI21X1 g4200(.A0(n5210), .A1(n4964), .B0(n5211), .Y(n5323));
  OAI21X1 g4201(.A0(n5323), .A1(n5322), .B0(n5139), .Y(n5324));
  OAI22X1 g4202(.A0(n4977), .A1(n2589), .B0(n2635), .B1(n4995), .Y(n5325));
  AOI21X1 g4203(.A0(n4993), .A1(n2545), .B0(n5325), .Y(n5326));
  AOI22X1 g4204(.A0(n2607), .A1(n5145), .B0(P1_U3084), .B1(P1_REG3_REG_12__SCAN_IN), .Y(n5327));
  OAI21X1 g4205(.A0(n5326), .A1(n4992), .B0(n5327), .Y(n5328));
  AOI21X1 g4206(.A0(n5152), .A1(n2590), .B0(n5328), .Y(n5329));
  NAND2X1 g4207(.A(n5329), .B(n5324), .Y(P1_U3222));
  INVX1   g4208(.A(n5225), .Y(n5331));
  AOI21X1 g4209(.A0(n5036), .A1(n5035), .B0(n5034), .Y(n5332));
  OAI21X1 g4210(.A0(n5331), .A1(n5037), .B0(n5332), .Y(n5333));
  AOI21X1 g4211(.A0(n5023), .A1(n5035), .B0(n5037), .Y(n5334));
  OAI21X1 g4212(.A0(n5023), .A1(n5035), .B0(n5334), .Y(n5335));
  AOI21X1 g4213(.A0(n5331), .A1(n5033), .B0(n5335), .Y(n5336));
  NOR2X1  g4214(.A(n5336), .B(n4983), .Y(n5337));
  NAND2X1 g4215(.A(n5337), .B(n5333), .Y(n5338));
  NAND2X1 g4216(.A(n5145), .B(n3000), .Y(n5339));
  OAI22X1 g4217(.A0(n4977), .A1(n2988), .B0(n3035), .B1(n4995), .Y(n5340));
  AOI21X1 g4218(.A0(n4993), .A1(n2948), .B0(n5340), .Y(n5341));
  OAI22X1 g4219(.A0(n4992), .A1(n5341), .B0(P1_STATE_REG_SCAN_IN), .B1(n2986), .Y(n5342));
  AOI21X1 g4220(.A0(n5152), .A1(n2989), .B0(n5342), .Y(n5343));
  NAND3X1 g4221(.A(n5343), .B(n5339), .C(n5338), .Y(P1_U3221));
  AOI22X1 g4222(.A0(n4984), .A1(P1_REG3_REG_1__SCAN_IN), .B0(n2025), .B1(n4993), .Y(n5345));
  OAI21X1 g4223(.A0(n4995), .A1(n2111), .B0(n5345), .Y(n5346));
  OAI22X1 g4224(.A0(n2102), .A1(n4998), .B0(P1_STATE_REG_SCAN_IN), .B1(n4278), .Y(n5347));
  AOI21X1 g4225(.A0(n5346), .A1(n4991), .B0(n5347), .Y(n5348));
  XOR2X1  g4226(.A(n5107), .B(n4930), .Y(n5349));
  XOR2X1  g4227(.A(n5349), .B(n5115), .Y(n5350));
  AOI22X1 g4228(.A0(n5152), .A1(P1_REG3_REG_1__SCAN_IN), .B0(n5139), .B1(n5350), .Y(n5351));
  NAND2X1 g4229(.A(n5351), .B(n5348), .Y(P1_U3220));
  XOR2X1  g4230(.A(n4902), .B(n4900), .Y(n5353));
  XOR2X1  g4231(.A(n5353), .B(n5123), .Y(n5354));
  OAI22X1 g4232(.A0(n4977), .A1(n2407), .B0(n2366), .B1(n5148), .Y(n5355));
  AOI21X1 g4233(.A0(n4994), .A1(n2453), .B0(n5355), .Y(n5356));
  AOI22X1 g4234(.A0(n2425), .A1(n5145), .B0(P1_U3084), .B1(P1_REG3_REG_8__SCAN_IN), .Y(n5357));
  OAI21X1 g4235(.A0(n5356), .A1(n4992), .B0(n5357), .Y(n5358));
  AOI21X1 g4236(.A0(n5152), .A1(n2408), .B0(n5358), .Y(n5359));
  OAI21X1 g4237(.A0(n5354), .A1(n4983), .B0(n5359), .Y(P1_U3219));
  INVX1   g4238(.A(n5088), .Y(n5361));
  OAI22X1 g4239(.A0(n4211), .A1(n3253), .B0(n3281), .B1(n4216), .Y(n5362));
  XOR2X1  g4240(.A(n5362), .B(n4207), .Y(n5363));
  AOI22X1 g4241(.A0(n4209), .A1(n3243), .B0(n3255), .B1(n4217), .Y(n5364));
  NAND2X1 g4242(.A(n5364), .B(n5363), .Y(n5365));
  INVX1   g4243(.A(n5365), .Y(n5366));
  NOR4X1  g4244(.A(n5361), .B(n5072), .C(n5008), .D(n5366), .Y(n5367));
  OAI22X1 g4245(.A0(n4872), .A1(n3290), .B0(n3324), .B1(n4211), .Y(n5368));
  XOR2X1  g4246(.A(n5368), .B(n4207), .Y(n5369));
  OAI22X1 g4247(.A0(n4211), .A1(n3290), .B0(n3324), .B1(n4216), .Y(n5370));
  XOR2X1  g4248(.A(n5370), .B(n5369), .Y(n5371));
  NOR2X1  g4249(.A(n5361), .B(n5080), .Y(n5372));
  NOR2X1  g4250(.A(n5364), .B(n5363), .Y(n5373));
  AOI21X1 g4251(.A0(n5372), .A1(n5365), .B0(n5373), .Y(n5374));
  OAI21X1 g4252(.A0(n5366), .A1(n5087), .B0(n5374), .Y(n5375));
  NOR3X1  g4253(.A(n5375), .B(n5371), .C(n5367), .Y(n5376));
  NAND3X1 g4254(.A(n5088), .B(n5135), .C(n5090), .Y(n5377));
  NOR3X1  g4255(.A(n5373), .B(n5372), .C(n5086), .Y(n5378));
  NAND2X1 g4256(.A(n5371), .B(n5365), .Y(n5379));
  AOI21X1 g4257(.A0(n5378), .A1(n5377), .B0(n5379), .Y(n5380));
  OAI21X1 g4258(.A0(n5380), .A1(n5376), .B0(n5139), .Y(n5381));
  NAND3X1 g4259(.A(n5145), .B(n2101), .C(n3323), .Y(n5382));
  AOI22X1 g4260(.A0(n4984), .A1(n3709), .B0(n3328), .B1(n4994), .Y(n5383));
  OAI21X1 g4261(.A0(n5148), .A1(n3253), .B0(n5383), .Y(n5384));
  OAI22X1 g4262(.A0(n3285), .A1(n4989), .B0(P1_STATE_REG_SCAN_IN), .B1(n3283), .Y(n5385));
  AOI21X1 g4263(.A0(n5384), .A1(n4991), .B0(n5385), .Y(n5386));
  NAND3X1 g4264(.A(n5386), .B(n5382), .C(n5381), .Y(P1_U3218));
  INVX1   g4265(.A(n5025), .Y(n5388));
  XOR2X1  g4266(.A(n5027), .B(n5388), .Y(n5389));
  NOR2X1  g4267(.A(n5389), .B(n5066), .Y(n5390));
  AOI21X1 g4268(.A0(n5067), .A1(n5029), .B0(n5131), .Y(n5391));
  OAI21X1 g4269(.A0(n5391), .A1(n5390), .B0(n5139), .Y(n5392));
  AOI22X1 g4270(.A0(n4984), .A1(n2902), .B0(n2948), .B1(n4994), .Y(n5393));
  OAI21X1 g4271(.A0(n5148), .A1(n2864), .B0(n5393), .Y(n5394));
  AOI22X1 g4272(.A0(n4991), .A1(n5394), .B0(P1_U3084), .B1(P1_REG3_REG_19__SCAN_IN), .Y(n5395));
  OAI21X1 g4273(.A0(n4989), .A1(n2901), .B0(n5395), .Y(n5396));
  AOI21X1 g4274(.A0(n5145), .A1(n2914), .B0(n5396), .Y(n5397));
  NAND2X1 g4275(.A(n5397), .B(n5392), .Y(P1_U3217));
  AOI21X1 g4276(.A0(n5105), .A1(n4942), .B0(n5106), .Y(n5399));
  OAI21X1 g4277(.A0(n5178), .A1(n4939), .B0(n5399), .Y(n5400));
  OAI22X1 g4278(.A0(n4942), .A1(n4928), .B0(n4925), .B1(n4923), .Y(n5401));
  AOI21X1 g4279(.A0(n4928), .A1(n4942), .B0(n5401), .Y(n5402));
  OAI21X1 g4280(.A0(n5116), .A1(n5177), .B0(n5402), .Y(n5403));
  NAND3X1 g4281(.A(n5403), .B(n5400), .C(n5139), .Y(n5404));
  OAI22X1 g4282(.A0(n4977), .A1(P1_REG3_REG_3__SCAN_IN), .B0(n2111), .B1(n5148), .Y(n5405));
  AOI21X1 g4283(.A0(n4994), .A1(n2208), .B0(n5405), .Y(n5406));
  AOI22X1 g4284(.A0(n2172), .A1(n5145), .B0(P1_U3084), .B1(P1_REG3_REG_3__SCAN_IN), .Y(n5407));
  OAI21X1 g4285(.A0(n5406), .A1(n4992), .B0(n5407), .Y(n5408));
  AOI21X1 g4286(.A0(n5152), .A1(n3507), .B0(n5408), .Y(n5409));
  NAND2X1 g4287(.A(n5409), .B(n5404), .Y(P1_U3216));
  XOR2X1  g4288(.A(n4891), .B(n4889), .Y(n5411));
  XOR2X1  g4289(.A(n5411), .B(n5125), .Y(n5412));
  OAI22X1 g4290(.A0(n4977), .A1(n2494), .B0(n2454), .B1(n5148), .Y(n5413));
  AOI21X1 g4291(.A0(n4994), .A1(n2545), .B0(n5413), .Y(n5414));
  AOI22X1 g4292(.A0(n2511), .A1(n5145), .B0(P1_U3084), .B1(P1_REG3_REG_10__SCAN_IN), .Y(n5415));
  OAI21X1 g4293(.A0(n5414), .A1(n4992), .B0(n5415), .Y(n5416));
  AOI21X1 g4294(.A0(n5152), .A1(n2495), .B0(n5416), .Y(n5417));
  OAI21X1 g4295(.A0(n5412), .A1(n4983), .B0(n5417), .Y(P1_U3215));
  XOR2X1  g4296(.A(n5011), .B(n5009), .Y(n5419));
  XOR2X1  g4297(.A(n5419), .B(n5134), .Y(n5420));
  NOR2X1  g4298(.A(n4995), .B(n3123), .Y(n5421));
  OAI22X1 g4299(.A0(n4977), .A1(n3067), .B0(n3035), .B1(n5148), .Y(n5422));
  OAI21X1 g4300(.A0(n5422), .A1(n5421), .B0(n4991), .Y(n5423));
  AOI22X1 g4301(.A0(n3663), .A1(n5152), .B0(P1_U3084), .B1(P1_REG3_REG_23__SCAN_IN), .Y(n5424));
  NAND2X1 g4302(.A(n5424), .B(n5423), .Y(n5425));
  AOI21X1 g4303(.A0(n5145), .A1(n3111), .B0(n5425), .Y(n5426));
  OAI21X1 g4304(.A0(n5420), .A1(n4983), .B0(n5426), .Y(P1_U3214));
  XOR2X1  g4305(.A(n4865), .B(n4863), .Y(n5428));
  XOR2X1  g4306(.A(n5428), .B(n5127), .Y(n5429));
  OAI22X1 g4307(.A0(n4977), .A1(n2676), .B0(n2726), .B1(n4995), .Y(n5430));
  AOI21X1 g4308(.A0(n4993), .A1(n2634), .B0(n5430), .Y(n5431));
  AOI22X1 g4309(.A0(n2718), .A1(n5145), .B0(P1_U3084), .B1(P1_REG3_REG_14__SCAN_IN), .Y(n5432));
  OAI21X1 g4310(.A0(n5431), .A1(n4992), .B0(n5432), .Y(n5433));
  AOI21X1 g4311(.A0(n5152), .A1(n2677), .B0(n5433), .Y(n5434));
  OAI21X1 g4312(.A0(n5429), .A1(n4983), .B0(n5434), .Y(P1_U3213));
  NOR3X1  g4313(.A(n5361), .B(n5072), .C(n5008), .Y(n5436));
  INVX1   g4314(.A(n5364), .Y(n5437));
  XOR2X1  g4315(.A(n5437), .B(n5363), .Y(n5438));
  NOR4X1  g4316(.A(n5436), .B(n5372), .C(n5086), .D(n5438), .Y(n5439));
  NOR2X1  g4317(.A(n5372), .B(n5086), .Y(n5440));
  INVX1   g4318(.A(n5438), .Y(n5441));
  AOI21X1 g4319(.A0(n5440), .A1(n5377), .B0(n5441), .Y(n5442));
  OAI21X1 g4320(.A0(n5442), .A1(n5439), .B0(n5139), .Y(n5443));
  NAND2X1 g4321(.A(n5145), .B(n3255), .Y(n5444));
  AOI22X1 g4322(.A0(n4984), .A1(n3699), .B0(n3198), .B1(n4993), .Y(n5445));
  OAI21X1 g4323(.A0(n4995), .A1(n3290), .B0(n5445), .Y(n5446));
  OAI22X1 g4324(.A0(n3239), .A1(n4989), .B0(P1_STATE_REG_SCAN_IN), .B1(n3237), .Y(n5447));
  AOI21X1 g4325(.A0(n5446), .A1(n4991), .B0(n5447), .Y(n5448));
  NAND3X1 g4326(.A(n5448), .B(n5444), .C(n5443), .Y(P1_U3212));
  OAI21X1 g4327(.A0(n4910), .A1(n4908), .B0(n4911), .Y(n5450));
  AOI21X1 g4328(.A0(n4952), .A1(n4950), .B0(n5450), .Y(n5451));
  AOI21X1 g4329(.A0(n4907), .A1(n4905), .B0(n4950), .Y(n5452));
  AOI21X1 g4330(.A0(n4954), .A1(n4908), .B0(n4951), .Y(n5453));
  OAI21X1 g4331(.A0(n4954), .A1(n4908), .B0(n5453), .Y(n5454));
  OAI21X1 g4332(.A0(n5454), .A1(n5452), .B0(n5139), .Y(n5455));
  OAI22X1 g4333(.A0(n4977), .A1(n2362), .B0(n2338), .B1(n5148), .Y(n5456));
  AOI21X1 g4334(.A0(n4994), .A1(n2410), .B0(n5456), .Y(n5457));
  AOI22X1 g4335(.A0(n2385), .A1(n5145), .B0(P1_U3084), .B1(P1_REG3_REG_7__SCAN_IN), .Y(n5458));
  OAI21X1 g4336(.A0(n5457), .A1(n4992), .B0(n5458), .Y(n5459));
  AOI21X1 g4337(.A0(n5152), .A1(n2363), .B0(n5459), .Y(n5460));
  OAI21X1 g4338(.A0(n5455), .A1(n5451), .B0(n5460), .Y(P1_U3211));
  AOI21X1 g4339(.A0(n1148), .A1(n1146), .B0(n1174), .Y(n5462));
  AOI21X1 g4340(.A0(n1159), .A1(n1156), .B0(n5462), .Y(n5463));
  NAND2X1 g4341(.A(P2_IR_REG_0__SCAN_IN), .B(P2_STATE_REG_SCAN_IN), .Y(n5464));
  OAI21X1 g4342(.A0(n5463), .A1(P2_STATE_REG_SCAN_IN), .B0(n5464), .Y(P2_U3358));
  AOI21X1 g4343(.A0(n1148), .A1(n1146), .B0(n1168), .Y(n5466));
  AOI21X1 g4344(.A0(n1181), .A1(n1156), .B0(n5466), .Y(n5467));
  INVX1   g4345(.A(P2_STATE_REG_SCAN_IN), .Y(P2_U3152));
  NOR2X1  g4346(.A(P2_IR_REG_31__SCAN_IN), .B(P2_U3152), .Y(n5469));
  INVX1   g4347(.A(P2_IR_REG_31__SCAN_IN), .Y(n5470));
  NOR2X1  g4348(.A(n5470), .B(P2_U3152), .Y(n5471));
  XOR2X1  g4349(.A(P2_IR_REG_1__SCAN_IN), .B(P2_IR_REG_0__SCAN_IN), .Y(n5472));
  AOI22X1 g4350(.A0(n5471), .A1(n5472), .B0(n5469), .B1(P2_IR_REG_1__SCAN_IN), .Y(n5473));
  OAI21X1 g4351(.A0(n5467), .A1(P2_STATE_REG_SCAN_IN), .B0(n5473), .Y(P2_U3357));
  AOI21X1 g4352(.A0(n1148), .A1(n1146), .B0(n1221), .Y(n5475));
  AOI21X1 g4353(.A0(n1197), .A1(n1156), .B0(n5475), .Y(n5476));
  INVX1   g4354(.A(P2_IR_REG_0__SCAN_IN), .Y(n5477));
  INVX1   g4355(.A(P2_IR_REG_1__SCAN_IN), .Y(n5478));
  NAND2X1 g4356(.A(n5478), .B(n5477), .Y(n5479));
  XOR2X1  g4357(.A(n5479), .B(P2_IR_REG_2__SCAN_IN), .Y(n5480));
  AOI22X1 g4358(.A0(n5471), .A1(n5480), .B0(n5469), .B1(P2_IR_REG_2__SCAN_IN), .Y(n5481));
  OAI21X1 g4359(.A0(n5476), .A1(P2_STATE_REG_SCAN_IN), .B0(n5481), .Y(P2_U3356));
  AOI21X1 g4360(.A0(n1148), .A1(n1146), .B0(n1224), .Y(n5483));
  AOI21X1 g4361(.A0(n1212), .A1(n1156), .B0(n5483), .Y(n5484));
  INVX1   g4362(.A(P2_IR_REG_3__SCAN_IN), .Y(n5485));
  NOR3X1  g4363(.A(P2_IR_REG_2__SCAN_IN), .B(P2_IR_REG_1__SCAN_IN), .C(P2_IR_REG_0__SCAN_IN), .Y(n5486));
  XOR2X1  g4364(.A(n5486), .B(n5485), .Y(n5487));
  AOI22X1 g4365(.A0(n5471), .A1(n5487), .B0(n5469), .B1(P2_IR_REG_3__SCAN_IN), .Y(n5488));
  OAI21X1 g4366(.A0(n5484), .A1(P2_STATE_REG_SCAN_IN), .B0(n5488), .Y(P2_U3355));
  AOI21X1 g4367(.A0(n1148), .A1(n1146), .B0(n1234), .Y(n5490));
  AOI21X1 g4368(.A0(n1239), .A1(n1156), .B0(n5490), .Y(n5491));
  INVX1   g4369(.A(P2_IR_REG_4__SCAN_IN), .Y(n5492));
  NOR4X1  g4370(.A(P2_IR_REG_2__SCAN_IN), .B(P2_IR_REG_1__SCAN_IN), .C(P2_IR_REG_0__SCAN_IN), .D(P2_IR_REG_3__SCAN_IN), .Y(n5493));
  XOR2X1  g4371(.A(n5493), .B(n5492), .Y(n5494));
  AOI22X1 g4372(.A0(n5471), .A1(n5494), .B0(n5469), .B1(P2_IR_REG_4__SCAN_IN), .Y(n5495));
  OAI21X1 g4373(.A0(n5491), .A1(P2_STATE_REG_SCAN_IN), .B0(n5495), .Y(P2_U3354));
  AOI21X1 g4374(.A0(n1148), .A1(n1146), .B0(n1252), .Y(n5497));
  AOI21X1 g4375(.A0(n1257), .A1(n1156), .B0(n5497), .Y(n5498));
  NAND2X1 g4376(.A(n5493), .B(n5492), .Y(n5499));
  XOR2X1  g4377(.A(n5499), .B(P2_IR_REG_5__SCAN_IN), .Y(n5500));
  AOI22X1 g4378(.A0(n5471), .A1(n5500), .B0(n5469), .B1(P2_IR_REG_5__SCAN_IN), .Y(n5501));
  OAI21X1 g4379(.A0(n5498), .A1(P2_STATE_REG_SCAN_IN), .B0(n5501), .Y(P2_U3353));
  AOI21X1 g4380(.A0(n1148), .A1(n1146), .B0(n1283), .Y(n5503));
  AOI21X1 g4381(.A0(n1288), .A1(n1156), .B0(n5503), .Y(n5504));
  INVX1   g4382(.A(P2_IR_REG_5__SCAN_IN), .Y(n5505));
  NAND3X1 g4383(.A(n5493), .B(n5505), .C(n5492), .Y(n5506));
  INVX1   g4384(.A(P2_IR_REG_6__SCAN_IN), .Y(n5507));
  NAND2X1 g4385(.A(n5507), .B(n5505), .Y(n5508));
  NOR2X1  g4386(.A(n5508), .B(n5499), .Y(n5509));
  AOI21X1 g4387(.A0(n5506), .A1(P2_IR_REG_6__SCAN_IN), .B0(n5509), .Y(n5510));
  AOI22X1 g4388(.A0(n5471), .A1(n5510), .B0(n5469), .B1(P2_IR_REG_6__SCAN_IN), .Y(n5511));
  OAI21X1 g4389(.A0(n5504), .A1(P2_STATE_REG_SCAN_IN), .B0(n5511), .Y(P2_U3352));
  AOI21X1 g4390(.A0(n1148), .A1(n1146), .B0(n1311), .Y(n5513));
  AOI21X1 g4391(.A0(n1316), .A1(n1156), .B0(n5513), .Y(n5514));
  INVX1   g4392(.A(P2_IR_REG_7__SCAN_IN), .Y(n5515));
  XOR2X1  g4393(.A(n5509), .B(n5515), .Y(n5516));
  AOI22X1 g4394(.A0(n5471), .A1(n5516), .B0(n5469), .B1(P2_IR_REG_7__SCAN_IN), .Y(n5517));
  OAI21X1 g4395(.A0(n5514), .A1(P2_STATE_REG_SCAN_IN), .B0(n5517), .Y(P2_U3351));
  INVX1   g4396(.A(P1_DATAO_REG_8__SCAN_IN), .Y(n5519));
  AOI21X1 g4397(.A0(n1148), .A1(n1146), .B0(n5519), .Y(n5520));
  AOI21X1 g4398(.A0(n1337), .A1(n1156), .B0(n5520), .Y(n5521));
  INVX1   g4399(.A(P2_IR_REG_8__SCAN_IN), .Y(n5522));
  AOI21X1 g4400(.A0(n5509), .A1(n5515), .B0(n5522), .Y(n5523));
  NOR4X1  g4401(.A(n5499), .B(P2_IR_REG_8__SCAN_IN), .C(P2_IR_REG_7__SCAN_IN), .D(n5508), .Y(n5524));
  NOR2X1  g4402(.A(n5524), .B(n5523), .Y(n5525));
  AOI22X1 g4403(.A0(n5471), .A1(n5525), .B0(n5469), .B1(P2_IR_REG_8__SCAN_IN), .Y(n5526));
  OAI21X1 g4404(.A0(n5521), .A1(P2_STATE_REG_SCAN_IN), .B0(n5526), .Y(P2_U3350));
  AOI21X1 g4405(.A0(n1148), .A1(n1146), .B0(n1369), .Y(n5528));
  AOI21X1 g4406(.A0(n1362), .A1(n1156), .B0(n5528), .Y(n5529));
  INVX1   g4407(.A(P2_IR_REG_9__SCAN_IN), .Y(n5530));
  XOR2X1  g4408(.A(n5524), .B(n5530), .Y(n5531));
  AOI22X1 g4409(.A0(n5471), .A1(n5531), .B0(n5469), .B1(P2_IR_REG_9__SCAN_IN), .Y(n5532));
  OAI21X1 g4410(.A0(n5529), .A1(P2_STATE_REG_SCAN_IN), .B0(n5532), .Y(P2_U3349));
  AOI21X1 g4411(.A0(n1148), .A1(n1146), .B0(n1394), .Y(n5534));
  AOI21X1 g4412(.A0(n1381), .A1(n1156), .B0(n5534), .Y(n5535));
  INVX1   g4413(.A(P2_IR_REG_10__SCAN_IN), .Y(n5536));
  AOI21X1 g4414(.A0(n5524), .A1(n5530), .B0(n5536), .Y(n5537));
  INVX1   g4415(.A(n5524), .Y(n5538));
  NOR3X1  g4416(.A(n5538), .B(P2_IR_REG_10__SCAN_IN), .C(P2_IR_REG_9__SCAN_IN), .Y(n5539));
  NOR2X1  g4417(.A(n5539), .B(n5537), .Y(n5540));
  AOI22X1 g4418(.A0(n5471), .A1(n5540), .B0(n5469), .B1(P2_IR_REG_10__SCAN_IN), .Y(n5541));
  OAI21X1 g4419(.A0(n5535), .A1(P2_STATE_REG_SCAN_IN), .B0(n5541), .Y(P2_U3348));
  AOI21X1 g4420(.A0(n1148), .A1(n1146), .B0(n1416), .Y(n5543));
  AOI21X1 g4421(.A0(n1407), .A1(n1156), .B0(n5543), .Y(n5544));
  INVX1   g4422(.A(P2_IR_REG_11__SCAN_IN), .Y(n5545));
  XOR2X1  g4423(.A(n5539), .B(n5545), .Y(n5546));
  AOI22X1 g4424(.A0(n5471), .A1(n5546), .B0(n5469), .B1(P2_IR_REG_11__SCAN_IN), .Y(n5547));
  OAI21X1 g4425(.A0(n5544), .A1(P2_STATE_REG_SCAN_IN), .B0(n5547), .Y(P2_U3347));
  OAI21X1 g4426(.A0(n1153), .A1(n1152), .B0(P1_DATAO_REG_12__SCAN_IN), .Y(n5549));
  INVX1   g4427(.A(n5549), .Y(n5550));
  AOI21X1 g4428(.A0(n1425), .A1(n1156), .B0(n5550), .Y(n5551));
  NAND4X1 g4429(.A(n5545), .B(n5536), .C(n5530), .D(n5524), .Y(n5552));
  NOR4X1  g4430(.A(P2_IR_REG_11__SCAN_IN), .B(P2_IR_REG_10__SCAN_IN), .C(P2_IR_REG_9__SCAN_IN), .D(P2_IR_REG_12__SCAN_IN), .Y(n5553));
  AOI22X1 g4431(.A0(n5552), .A1(P2_IR_REG_12__SCAN_IN), .B0(n5524), .B1(n5553), .Y(n5554));
  AOI22X1 g4432(.A0(n5471), .A1(n5554), .B0(n5469), .B1(P2_IR_REG_12__SCAN_IN), .Y(n5555));
  OAI21X1 g4433(.A0(n5551), .A1(P2_STATE_REG_SCAN_IN), .B0(n5555), .Y(P2_U3346));
  AOI21X1 g4434(.A0(n1148), .A1(n1146), .B0(n1441), .Y(n5557));
  AOI21X1 g4435(.A0(n1445), .A1(n1156), .B0(n5557), .Y(n5558));
  INVX1   g4436(.A(P2_IR_REG_13__SCAN_IN), .Y(n5559));
  INVX1   g4437(.A(n5553), .Y(n5560));
  NOR2X1  g4438(.A(n5560), .B(n5538), .Y(n5561));
  XOR2X1  g4439(.A(n5561), .B(n5559), .Y(n5562));
  AOI22X1 g4440(.A0(n5471), .A1(n5562), .B0(n5469), .B1(P2_IR_REG_13__SCAN_IN), .Y(n5563));
  OAI21X1 g4441(.A0(n5558), .A1(P2_STATE_REG_SCAN_IN), .B0(n5563), .Y(P2_U3345));
  INVX1   g4442(.A(P1_DATAO_REG_14__SCAN_IN), .Y(n5565));
  AOI21X1 g4443(.A0(n1148), .A1(n1146), .B0(n5565), .Y(n5566));
  AOI21X1 g4444(.A0(n1463), .A1(n1156), .B0(n5566), .Y(n5567));
  NAND3X1 g4445(.A(n5553), .B(n5524), .C(n5559), .Y(n5568));
  NOR4X1  g4446(.A(n5538), .B(P2_IR_REG_14__SCAN_IN), .C(P2_IR_REG_13__SCAN_IN), .D(n5560), .Y(n5569));
  AOI21X1 g4447(.A0(n5568), .A1(P2_IR_REG_14__SCAN_IN), .B0(n5569), .Y(n5570));
  AOI22X1 g4448(.A0(n5471), .A1(n5570), .B0(n5469), .B1(P2_IR_REG_14__SCAN_IN), .Y(n5571));
  OAI21X1 g4449(.A0(n5567), .A1(P2_STATE_REG_SCAN_IN), .B0(n5571), .Y(P2_U3344));
  OAI21X1 g4450(.A0(n1153), .A1(n1152), .B0(P1_DATAO_REG_15__SCAN_IN), .Y(n5573));
  INVX1   g4451(.A(n5573), .Y(n5574));
  AOI21X1 g4452(.A0(n1490), .A1(n1156), .B0(n5574), .Y(n5575));
  INVX1   g4453(.A(P2_IR_REG_15__SCAN_IN), .Y(n5576));
  XOR2X1  g4454(.A(n5569), .B(n5576), .Y(n5577));
  AOI22X1 g4455(.A0(n5471), .A1(n5577), .B0(n5469), .B1(P2_IR_REG_15__SCAN_IN), .Y(n5578));
  OAI21X1 g4456(.A0(n5575), .A1(P2_STATE_REG_SCAN_IN), .B0(n5578), .Y(P2_U3343));
  OAI21X1 g4457(.A0(n1153), .A1(n1152), .B0(P1_DATAO_REG_16__SCAN_IN), .Y(n5580));
  INVX1   g4458(.A(n5580), .Y(n5581));
  AOI21X1 g4459(.A0(n1510), .A1(n1156), .B0(n5581), .Y(n5582));
  NAND2X1 g4460(.A(n5569), .B(n5576), .Y(n5583));
  NOR4X1  g4461(.A(P2_IR_REG_15__SCAN_IN), .B(P2_IR_REG_14__SCAN_IN), .C(P2_IR_REG_13__SCAN_IN), .D(P2_IR_REG_16__SCAN_IN), .Y(n5584));
  NAND3X1 g4462(.A(n5584), .B(n5553), .C(n5524), .Y(n5585));
  AOI21X1 g4463(.A0(n5583), .A1(P2_IR_REG_16__SCAN_IN), .B0(n5617), .Y(n5587));
  AOI22X1 g4464(.A0(n5471), .A1(n5587), .B0(n5469), .B1(P2_IR_REG_16__SCAN_IN), .Y(n5588));
  OAI21X1 g4465(.A0(n5582), .A1(P2_STATE_REG_SCAN_IN), .B0(n5588), .Y(P2_U3342));
  OAI21X1 g4466(.A0(n1153), .A1(n1152), .B0(P1_DATAO_REG_17__SCAN_IN), .Y(n5590));
  INVX1   g4467(.A(n5590), .Y(n5591));
  AOI21X1 g4468(.A0(n1540), .A1(n1156), .B0(n5591), .Y(n5592));
  XOR2X1  g4469(.A(n5585), .B(P2_IR_REG_17__SCAN_IN), .Y(n5593));
  AOI22X1 g4470(.A0(n5471), .A1(n5593), .B0(n5469), .B1(P2_IR_REG_17__SCAN_IN), .Y(n5594));
  OAI21X1 g4471(.A0(n5592), .A1(P2_STATE_REG_SCAN_IN), .B0(n5594), .Y(P2_U3341));
  OAI21X1 g4472(.A0(n1153), .A1(n1152), .B0(P1_DATAO_REG_18__SCAN_IN), .Y(n5596));
  INVX1   g4473(.A(n5596), .Y(n5597));
  AOI21X1 g4474(.A0(n1558), .A1(n1156), .B0(n5597), .Y(n5598));
  INVX1   g4475(.A(P2_IR_REG_18__SCAN_IN), .Y(n5599));
  INVX1   g4476(.A(P2_IR_REG_2__SCAN_IN), .Y(n5600));
  NAND4X1 g4477(.A(n5492), .B(n5485), .C(n5600), .D(n5505), .Y(n5601));
  NOR3X1  g4478(.A(P2_IR_REG_12__SCAN_IN), .B(P2_IR_REG_11__SCAN_IN), .C(P2_IR_REG_10__SCAN_IN), .Y(n5602));
  NOR4X1  g4479(.A(P2_IR_REG_8__SCAN_IN), .B(P2_IR_REG_7__SCAN_IN), .C(P2_IR_REG_6__SCAN_IN), .D(P2_IR_REG_9__SCAN_IN), .Y(n5603));
  NAND3X1 g4480(.A(n5603), .B(n5602), .C(n5584), .Y(n5604));
  NOR4X1  g4481(.A(n5601), .B(n5479), .C(P2_IR_REG_17__SCAN_IN), .D(n5604), .Y(n5605));
  NOR2X1  g4482(.A(P2_IR_REG_18__SCAN_IN), .B(P2_IR_REG_17__SCAN_IN), .Y(n5606));
  INVX1   g4483(.A(n5606), .Y(n5607));
  NOR4X1  g4484(.A(n5604), .B(n5601), .C(n5479), .D(n5607), .Y(n5608));
  INVX1   g4485(.A(n5608), .Y(n5609));
  OAI21X1 g4486(.A0(n5605), .A1(n5599), .B0(n5609), .Y(n5610));
  INVX1   g4487(.A(n5610), .Y(n5611));
  AOI22X1 g4488(.A0(n5471), .A1(n5611), .B0(n5469), .B1(P2_IR_REG_18__SCAN_IN), .Y(n5612));
  OAI21X1 g4489(.A0(n5598), .A1(P2_STATE_REG_SCAN_IN), .B0(n5612), .Y(P2_U3340));
  OAI21X1 g4490(.A0(n1153), .A1(n1152), .B0(P1_DATAO_REG_19__SCAN_IN), .Y(n5614));
  INVX1   g4491(.A(n5614), .Y(n5615));
  AOI21X1 g4492(.A0(n1586), .A1(n1156), .B0(n5615), .Y(n5616));
  NOR3X1  g4493(.A(n5604), .B(n5601), .C(n5479), .Y(n5617));
  NOR3X1  g4494(.A(P2_IR_REG_19__SCAN_IN), .B(P2_IR_REG_18__SCAN_IN), .C(P2_IR_REG_17__SCAN_IN), .Y(n5618));
  AOI22X1 g4495(.A0(n5609), .A1(P2_IR_REG_19__SCAN_IN), .B0(n5617), .B1(n5618), .Y(n5619));
  AOI22X1 g4496(.A0(n5471), .A1(n5619), .B0(n5469), .B1(P2_IR_REG_19__SCAN_IN), .Y(n5620));
  OAI21X1 g4497(.A0(n5616), .A1(P2_STATE_REG_SCAN_IN), .B0(n5620), .Y(P2_U3339));
  OAI21X1 g4498(.A0(n1153), .A1(n1152), .B0(P1_DATAO_REG_20__SCAN_IN), .Y(n5622));
  INVX1   g4499(.A(n5622), .Y(n5623));
  AOI21X1 g4500(.A0(n1609), .A1(n1156), .B0(n5623), .Y(n5624));
  INVX1   g4501(.A(P2_IR_REG_20__SCAN_IN), .Y(n5625));
  AOI21X1 g4502(.A0(n5618), .A1(n5617), .B0(n5625), .Y(n5626));
  NOR4X1  g4503(.A(P2_IR_REG_19__SCAN_IN), .B(P2_IR_REG_18__SCAN_IN), .C(P2_IR_REG_17__SCAN_IN), .D(P2_IR_REG_20__SCAN_IN), .Y(n5627));
  AOI21X1 g4504(.A0(n5627), .A1(n5617), .B0(n5626), .Y(n5628));
  AOI22X1 g4505(.A0(n5471), .A1(n5628), .B0(n5469), .B1(P2_IR_REG_20__SCAN_IN), .Y(n5629));
  OAI21X1 g4506(.A0(n5624), .A1(P2_STATE_REG_SCAN_IN), .B0(n5629), .Y(P2_U3338));
  OAI21X1 g4507(.A0(n1153), .A1(n1152), .B0(P1_DATAO_REG_21__SCAN_IN), .Y(n5631));
  INVX1   g4508(.A(n5631), .Y(n5632));
  AOI21X1 g4509(.A0(n1634), .A1(n1156), .B0(n5632), .Y(n5633));
  NOR4X1  g4510(.A(n5585), .B(P2_IR_REG_20__SCAN_IN), .C(P2_IR_REG_19__SCAN_IN), .D(n5607), .Y(n5636));
  XOR2X1  g4511(.A(n5636), .B(P2_IR_REG_21__SCAN_IN), .Y(n5637));
  NOR3X1  g4512(.A(n5637), .B(n5470), .C(P2_U3152), .Y(n5638));
  AOI21X1 g4513(.A0(n5469), .A1(P2_IR_REG_21__SCAN_IN), .B0(n5638), .Y(n5639));
  OAI21X1 g4514(.A0(n5633), .A1(P2_STATE_REG_SCAN_IN), .B0(n5639), .Y(P2_U3337));
  OAI21X1 g4515(.A0(n1153), .A1(n1152), .B0(P1_DATAO_REG_22__SCAN_IN), .Y(n5641));
  INVX1   g4516(.A(n5641), .Y(n5642));
  AOI21X1 g4517(.A0(n1652), .A1(n1156), .B0(n5642), .Y(n5643));
  INVX1   g4518(.A(P2_IR_REG_22__SCAN_IN), .Y(n5644));
  INVX1   g4519(.A(P2_IR_REG_19__SCAN_IN), .Y(n5645));
  NOR2X1  g4520(.A(P2_IR_REG_22__SCAN_IN), .B(P2_IR_REG_21__SCAN_IN), .Y(n5646));
  NAND3X1 g4521(.A(n5646), .B(n5625), .C(n5645), .Y(n5647));
  NOR3X1  g4522(.A(n5647), .B(n5607), .C(n5585), .Y(n5648));
  AOI21X1 g4523(.A0(P2_IR_REG_22__SCAN_IN), .A1(P2_IR_REG_21__SCAN_IN), .B0(n5648), .Y(n5649));
  OAI21X1 g4524(.A0(n5636), .A1(n5644), .B0(n5649), .Y(n5650));
  NOR3X1  g4525(.A(n5650), .B(n5470), .C(P2_U3152), .Y(n5651));
  AOI21X1 g4526(.A0(n5469), .A1(P2_IR_REG_22__SCAN_IN), .B0(n5651), .Y(n5652));
  OAI21X1 g4527(.A0(n5643), .A1(P2_STATE_REG_SCAN_IN), .B0(n5652), .Y(P2_U3336));
  OAI21X1 g4528(.A0(n1153), .A1(n1152), .B0(P1_DATAO_REG_23__SCAN_IN), .Y(n5654));
  INVX1   g4529(.A(n5654), .Y(n5655));
  AOI21X1 g4530(.A0(n1676), .A1(n1156), .B0(n5655), .Y(n5656));
  INVX1   g4531(.A(P2_IR_REG_23__SCAN_IN), .Y(n5657));
  XOR2X1  g4532(.A(n5648), .B(n5657), .Y(n5658));
  AOI22X1 g4533(.A0(n5471), .A1(n5658), .B0(n5469), .B1(P2_IR_REG_23__SCAN_IN), .Y(n5659));
  OAI21X1 g4534(.A0(n5656), .A1(P2_STATE_REG_SCAN_IN), .B0(n5659), .Y(P2_U3335));
  NAND2X1 g4535(.A(n1721), .B(n1719), .Y(n5661));
  XOR2X1  g4536(.A(n1701), .B(n5661), .Y(n5662));
  OAI21X1 g4537(.A0(n1153), .A1(n1152), .B0(P1_DATAO_REG_24__SCAN_IN), .Y(n5663));
  OAI21X1 g4538(.A0(n5662), .A1(n1149), .B0(n5663), .Y(n5664));
  INVX1   g4539(.A(n5664), .Y(n5665));
  INVX1   g4540(.A(P2_IR_REG_24__SCAN_IN), .Y(n5666));
  NOR4X1  g4541(.A(n5607), .B(n5585), .C(P2_IR_REG_23__SCAN_IN), .D(n5647), .Y(n5667));
  XOR2X1  g4542(.A(n5667), .B(n5666), .Y(n5668));
  AOI22X1 g4543(.A0(n5471), .A1(n5668), .B0(n5469), .B1(P2_IR_REG_24__SCAN_IN), .Y(n5669));
  OAI21X1 g4544(.A0(n5665), .A1(P2_STATE_REG_SCAN_IN), .B0(n5669), .Y(P2_U3334));
  OAI21X1 g4545(.A0(n1153), .A1(n1152), .B0(P1_DATAO_REG_25__SCAN_IN), .Y(n5671));
  INVX1   g4546(.A(n5671), .Y(n5672));
  AOI21X1 g4547(.A0(n1727), .A1(n1156), .B0(n5672), .Y(n5673));
  NOR4X1  g4548(.A(P2_IR_REG_23__SCAN_IN), .B(P2_IR_REG_22__SCAN_IN), .C(P2_IR_REG_21__SCAN_IN), .D(P2_IR_REG_24__SCAN_IN), .Y(n5674));
  NAND3X1 g4549(.A(n5674), .B(n5627), .C(n5617), .Y(n5675));
  XOR2X1  g4550(.A(n5675), .B(P2_IR_REG_25__SCAN_IN), .Y(n5676));
  AOI22X1 g4551(.A0(n5471), .A1(n5676), .B0(n5469), .B1(P2_IR_REG_25__SCAN_IN), .Y(n5677));
  OAI21X1 g4552(.A0(n5673), .A1(P2_STATE_REG_SCAN_IN), .B0(n5677), .Y(P2_U3333));
  OAI21X1 g4553(.A0(n1153), .A1(n1152), .B0(P1_DATAO_REG_26__SCAN_IN), .Y(n5679));
  INVX1   g4554(.A(n5679), .Y(n5680));
  AOI21X1 g4555(.A0(n1745), .A1(n1156), .B0(n5680), .Y(n5681));
  OAI21X1 g4556(.A0(n5675), .A1(P2_IR_REG_25__SCAN_IN), .B0(P2_IR_REG_26__SCAN_IN), .Y(n5682));
  INVX1   g4557(.A(P2_IR_REG_25__SCAN_IN), .Y(n5683));
  INVX1   g4558(.A(P2_IR_REG_26__SCAN_IN), .Y(n5684));
  NAND2X1 g4559(.A(n5684), .B(n5683), .Y(n5685));
  OAI21X1 g4560(.A0(n5685), .A1(n5675), .B0(n5682), .Y(n5686));
  INVX1   g4561(.A(n5686), .Y(n5687));
  AOI22X1 g4562(.A0(n5471), .A1(n5687), .B0(n5469), .B1(P2_IR_REG_26__SCAN_IN), .Y(n5688));
  OAI21X1 g4563(.A0(n5681), .A1(P2_STATE_REG_SCAN_IN), .B0(n5688), .Y(P2_U3332));
  NAND3X1 g4564(.A(n1774), .B(n1773), .C(n1771), .Y(n5690));
  OAI21X1 g4565(.A0(n1766), .A1(n1762), .B0(n1769), .Y(n5691));
  AOI21X1 g4566(.A0(n5691), .A1(n5690), .B0(n1149), .Y(n5692));
  OAI21X1 g4567(.A0(n1153), .A1(n1152), .B0(P1_DATAO_REG_27__SCAN_IN), .Y(n5693));
  INVX1   g4568(.A(n5693), .Y(n5694));
  NOR2X1  g4569(.A(n5694), .B(n5692), .Y(n5695));
  INVX1   g4570(.A(P2_IR_REG_27__SCAN_IN), .Y(n5696));
  NAND2X1 g4571(.A(n5674), .B(n5627), .Y(n5697));
  NOR3X1  g4572(.A(n5685), .B(n5697), .C(n5585), .Y(n5698));
  XOR2X1  g4573(.A(n5698), .B(n5696), .Y(n5699));
  AOI22X1 g4574(.A0(n5471), .A1(n5699), .B0(n5469), .B1(P2_IR_REG_27__SCAN_IN), .Y(n5700));
  OAI21X1 g4575(.A0(n5695), .A1(P2_STATE_REG_SCAN_IN), .B0(n5700), .Y(P2_U3331));
  OAI21X1 g4576(.A0(n1153), .A1(n1152), .B0(P1_DATAO_REG_28__SCAN_IN), .Y(n5702));
  INVX1   g4577(.A(n5702), .Y(n5703));
  AOI21X1 g4578(.A0(n1792), .A1(n1156), .B0(n5703), .Y(n5704));
  INVX1   g4579(.A(P2_IR_REG_28__SCAN_IN), .Y(n5705));
  NOR4X1  g4580(.A(n5697), .B(n5585), .C(P2_IR_REG_27__SCAN_IN), .D(n5685), .Y(n5706));
  XOR2X1  g4581(.A(n5706), .B(n5705), .Y(n5707));
  AOI22X1 g4582(.A0(n5471), .A1(n5707), .B0(n5469), .B1(P2_IR_REG_28__SCAN_IN), .Y(n5708));
  OAI21X1 g4583(.A0(n5704), .A1(P2_STATE_REG_SCAN_IN), .B0(n5708), .Y(P2_U3330));
  OAI21X1 g4584(.A0(n1153), .A1(n1152), .B0(P1_DATAO_REG_29__SCAN_IN), .Y(n5710));
  INVX1   g4585(.A(n5710), .Y(n5711));
  AOI21X1 g4586(.A0(n1821), .A1(n1156), .B0(n5711), .Y(n5712));
  INVX1   g4587(.A(P2_IR_REG_29__SCAN_IN), .Y(n5713));
  NOR4X1  g4588(.A(n5675), .B(P2_IR_REG_28__SCAN_IN), .C(P2_IR_REG_27__SCAN_IN), .D(n5685), .Y(n5714));
  XOR2X1  g4589(.A(n5714), .B(n5713), .Y(n5715));
  AOI22X1 g4590(.A0(n5471), .A1(n5715), .B0(n5469), .B1(P2_IR_REG_29__SCAN_IN), .Y(n5716));
  OAI21X1 g4591(.A0(n5712), .A1(P2_STATE_REG_SCAN_IN), .B0(n5716), .Y(P2_U3329));
  AOI21X1 g4592(.A0(n1846), .A1(n1841), .B0(n1149), .Y(n5718));
  OAI21X1 g4593(.A0(n1153), .A1(n1152), .B0(P1_DATAO_REG_30__SCAN_IN), .Y(n5719));
  INVX1   g4594(.A(n5719), .Y(n5720));
  NOR2X1  g4595(.A(n5720), .B(n5718), .Y(n5721));
  NAND2X1 g4596(.A(n5714), .B(n5713), .Y(n5722));
  XOR2X1  g4597(.A(n5722), .B(P2_IR_REG_30__SCAN_IN), .Y(n5723));
  AOI22X1 g4598(.A0(n5471), .A1(n5723), .B0(n5469), .B1(P2_IR_REG_30__SCAN_IN), .Y(n5724));
  OAI21X1 g4599(.A0(n5721), .A1(P2_STATE_REG_SCAN_IN), .B0(n5724), .Y(P2_U3328));
  NAND4X1 g4600(.A(n3394), .B(n3393), .C(n1156), .D(n1866), .Y(n5726));
  OAI21X1 g4601(.A0(n1153), .A1(n1152), .B0(P1_DATAO_REG_31__SCAN_IN), .Y(n5727));
  NAND2X1 g4602(.A(n5727), .B(n5726), .Y(n5728));
  NAND2X1 g4603(.A(n5728), .B(P2_U3152), .Y(n5729));
  NOR2X1  g4604(.A(n5722), .B(P2_IR_REG_30__SCAN_IN), .Y(n5730));
  NAND3X1 g4605(.A(n5730), .B(P2_IR_REG_31__SCAN_IN), .C(P2_STATE_REG_SCAN_IN), .Y(n5731));
  NAND2X1 g4606(.A(n5731), .B(n5729), .Y(P2_U3327));
  NOR2X1  g4607(.A(P2_IR_REG_31__SCAN_IN), .B(n5657), .Y(n5733));
  AOI21X1 g4608(.A0(n5658), .A1(P2_IR_REG_31__SCAN_IN), .B0(n5733), .Y(n5734));
  INVX1   g4609(.A(n5734), .Y(n5735));
  NOR2X1  g4610(.A(P2_IR_REG_31__SCAN_IN), .B(n5684), .Y(n5736));
  AOI21X1 g4611(.A0(n5687), .A1(P2_IR_REG_31__SCAN_IN), .B0(n5736), .Y(n5737));
  NOR2X1  g4612(.A(P2_IR_REG_31__SCAN_IN), .B(n5666), .Y(n5738));
  AOI21X1 g4613(.A0(n5668), .A1(P2_IR_REG_31__SCAN_IN), .B0(n5738), .Y(n5739));
  NOR2X1  g4614(.A(P2_IR_REG_31__SCAN_IN), .B(n5683), .Y(n5740));
  AOI21X1 g4615(.A0(n5676), .A1(P2_IR_REG_31__SCAN_IN), .B0(n5740), .Y(n5741));
  NOR3X1  g4616(.A(n5741), .B(n5739), .C(n5737), .Y(n5742));
  NOR3X1  g4617(.A(n5742), .B(n5735), .C(P2_U3152), .Y(n5743));
  INVX1   g4618(.A(n5737), .Y(n5744));
  INVX1   g4619(.A(n5741), .Y(n5745));
  XOR2X1  g4620(.A(n5739), .B(P2_B_REG_SCAN_IN), .Y(n5746));
  OAI21X1 g4621(.A0(n5746), .A1(n5745), .B0(n5744), .Y(n5747));
  OAI21X1 g4622(.A0(n5745), .A1(n5737), .B0(n5739), .Y(n5748));
  NAND3X1 g4623(.A(n5748), .B(n5747), .C(n5743), .Y(n5749));
  INVX1   g4624(.A(n5743), .Y(n5750));
  INVX1   g4625(.A(n5747), .Y(n5751));
  OAI21X1 g4626(.A0(n5751), .A1(n5750), .B0(P2_D_REG_0__SCAN_IN), .Y(n5752));
  NAND2X1 g4627(.A(n5752), .B(n5749), .Y(P2_U3437));
  NAND2X1 g4628(.A(n5741), .B(n5737), .Y(n5754));
  NAND3X1 g4629(.A(n5754), .B(n5747), .C(n5743), .Y(n5755));
  OAI21X1 g4630(.A0(n5751), .A1(n5750), .B0(P2_D_REG_1__SCAN_IN), .Y(n5756));
  NAND2X1 g4631(.A(n5756), .B(n5755), .Y(P2_U3438));
  INVX1   g4632(.A(P2_D_REG_2__SCAN_IN), .Y(n5758));
  AOI21X1 g4633(.A0(n5747), .A1(n5743), .B0(n5758), .Y(P2_U3326));
  INVX1   g4634(.A(P2_D_REG_3__SCAN_IN), .Y(n5760));
  AOI21X1 g4635(.A0(n5747), .A1(n5743), .B0(n5760), .Y(P2_U3325));
  INVX1   g4636(.A(P2_D_REG_4__SCAN_IN), .Y(n5762));
  AOI21X1 g4637(.A0(n5747), .A1(n5743), .B0(n5762), .Y(P2_U3324));
  INVX1   g4638(.A(P2_D_REG_5__SCAN_IN), .Y(n5764));
  AOI21X1 g4639(.A0(n5747), .A1(n5743), .B0(n5764), .Y(P2_U3323));
  INVX1   g4640(.A(P2_D_REG_6__SCAN_IN), .Y(n5766));
  AOI21X1 g4641(.A0(n5747), .A1(n5743), .B0(n5766), .Y(P2_U3322));
  INVX1   g4642(.A(P2_D_REG_7__SCAN_IN), .Y(n5768));
  AOI21X1 g4643(.A0(n5747), .A1(n5743), .B0(n5768), .Y(P2_U3321));
  INVX1   g4644(.A(P2_D_REG_8__SCAN_IN), .Y(n5770));
  AOI21X1 g4645(.A0(n5747), .A1(n5743), .B0(n5770), .Y(P2_U3320));
  INVX1   g4646(.A(P2_D_REG_9__SCAN_IN), .Y(n5772));
  AOI21X1 g4647(.A0(n5747), .A1(n5743), .B0(n5772), .Y(P2_U3319));
  INVX1   g4648(.A(P2_D_REG_10__SCAN_IN), .Y(n5774));
  AOI21X1 g4649(.A0(n5747), .A1(n5743), .B0(n5774), .Y(P2_U3318));
  INVX1   g4650(.A(P2_D_REG_11__SCAN_IN), .Y(n5776));
  AOI21X1 g4651(.A0(n5747), .A1(n5743), .B0(n5776), .Y(P2_U3317));
  INVX1   g4652(.A(P2_D_REG_12__SCAN_IN), .Y(n5778));
  AOI21X1 g4653(.A0(n5747), .A1(n5743), .B0(n5778), .Y(P2_U3316));
  INVX1   g4654(.A(P2_D_REG_13__SCAN_IN), .Y(n5780));
  AOI21X1 g4655(.A0(n5747), .A1(n5743), .B0(n5780), .Y(P2_U3315));
  INVX1   g4656(.A(P2_D_REG_14__SCAN_IN), .Y(n5782));
  AOI21X1 g4657(.A0(n5747), .A1(n5743), .B0(n5782), .Y(P2_U3314));
  INVX1   g4658(.A(P2_D_REG_15__SCAN_IN), .Y(n5784));
  AOI21X1 g4659(.A0(n5747), .A1(n5743), .B0(n5784), .Y(P2_U3313));
  INVX1   g4660(.A(P2_D_REG_16__SCAN_IN), .Y(n5786));
  AOI21X1 g4661(.A0(n5747), .A1(n5743), .B0(n5786), .Y(P2_U3312));
  INVX1   g4662(.A(P2_D_REG_17__SCAN_IN), .Y(n5788));
  AOI21X1 g4663(.A0(n5747), .A1(n5743), .B0(n5788), .Y(P2_U3311));
  INVX1   g4664(.A(P2_D_REG_18__SCAN_IN), .Y(n5790));
  AOI21X1 g4665(.A0(n5747), .A1(n5743), .B0(n5790), .Y(P2_U3310));
  INVX1   g4666(.A(P2_D_REG_19__SCAN_IN), .Y(n5792));
  AOI21X1 g4667(.A0(n5747), .A1(n5743), .B0(n5792), .Y(P2_U3309));
  INVX1   g4668(.A(P2_D_REG_20__SCAN_IN), .Y(n5794));
  AOI21X1 g4669(.A0(n5747), .A1(n5743), .B0(n5794), .Y(P2_U3308));
  INVX1   g4670(.A(P2_D_REG_21__SCAN_IN), .Y(n5796));
  AOI21X1 g4671(.A0(n5747), .A1(n5743), .B0(n5796), .Y(P2_U3307));
  INVX1   g4672(.A(P2_D_REG_22__SCAN_IN), .Y(n5798));
  AOI21X1 g4673(.A0(n5747), .A1(n5743), .B0(n5798), .Y(P2_U3306));
  INVX1   g4674(.A(P2_D_REG_23__SCAN_IN), .Y(n5800));
  AOI21X1 g4675(.A0(n5747), .A1(n5743), .B0(n5800), .Y(P2_U3305));
  INVX1   g4676(.A(P2_D_REG_24__SCAN_IN), .Y(n5802));
  AOI21X1 g4677(.A0(n5747), .A1(n5743), .B0(n5802), .Y(P2_U3304));
  INVX1   g4678(.A(P2_D_REG_25__SCAN_IN), .Y(n5804));
  AOI21X1 g4679(.A0(n5747), .A1(n5743), .B0(n5804), .Y(P2_U3303));
  INVX1   g4680(.A(P2_D_REG_26__SCAN_IN), .Y(n5806));
  AOI21X1 g4681(.A0(n5747), .A1(n5743), .B0(n5806), .Y(P2_U3302));
  INVX1   g4682(.A(P2_D_REG_27__SCAN_IN), .Y(n5808));
  AOI21X1 g4683(.A0(n5747), .A1(n5743), .B0(n5808), .Y(P2_U3301));
  INVX1   g4684(.A(P2_D_REG_28__SCAN_IN), .Y(n5810));
  AOI21X1 g4685(.A0(n5747), .A1(n5743), .B0(n5810), .Y(P2_U3300));
  INVX1   g4686(.A(P2_D_REG_29__SCAN_IN), .Y(n5812));
  AOI21X1 g4687(.A0(n5747), .A1(n5743), .B0(n5812), .Y(P2_U3299));
  INVX1   g4688(.A(P2_D_REG_30__SCAN_IN), .Y(n5814));
  AOI21X1 g4689(.A0(n5747), .A1(n5743), .B0(n5814), .Y(P2_U3298));
  INVX1   g4690(.A(P2_D_REG_31__SCAN_IN), .Y(n5816));
  AOI21X1 g4691(.A0(n5747), .A1(n5743), .B0(n5816), .Y(P2_U3297));
  OAI21X1 g4692(.A0(P2_D_REG_7__SCAN_IN), .A1(P2_D_REG_3__SCAN_IN), .B0(n5751), .Y(n5818));
  OAI21X1 g4693(.A0(P2_D_REG_9__SCAN_IN), .A1(P2_D_REG_8__SCAN_IN), .B0(n5751), .Y(n5819));
  OAI21X1 g4694(.A0(P2_D_REG_10__SCAN_IN), .A1(P2_D_REG_5__SCAN_IN), .B0(n5751), .Y(n5820));
  OAI21X1 g4695(.A0(P2_D_REG_6__SCAN_IN), .A1(P2_D_REG_4__SCAN_IN), .B0(n5751), .Y(n5821));
  NAND4X1 g4696(.A(n5820), .B(n5819), .C(n5818), .D(n5821), .Y(n5822));
  OAI21X1 g4697(.A0(P2_D_REG_28__SCAN_IN), .A1(P2_D_REG_27__SCAN_IN), .B0(n5751), .Y(n5823));
  OAI21X1 g4698(.A0(P2_D_REG_26__SCAN_IN), .A1(P2_D_REG_25__SCAN_IN), .B0(n5751), .Y(n5824));
  OAI21X1 g4699(.A0(P2_D_REG_31__SCAN_IN), .A1(P2_D_REG_30__SCAN_IN), .B0(n5751), .Y(n5825));
  OAI21X1 g4700(.A0(P2_D_REG_29__SCAN_IN), .A1(P2_D_REG_2__SCAN_IN), .B0(n5751), .Y(n5826));
  NAND4X1 g4701(.A(n5825), .B(n5824), .C(n5823), .D(n5826), .Y(n5827));
  OAI21X1 g4702(.A0(P2_D_REG_21__SCAN_IN), .A1(P2_D_REG_20__SCAN_IN), .B0(n5751), .Y(n5828));
  OAI21X1 g4703(.A0(P2_D_REG_19__SCAN_IN), .A1(P2_D_REG_18__SCAN_IN), .B0(n5751), .Y(n5829));
  OAI21X1 g4704(.A0(P2_D_REG_23__SCAN_IN), .A1(P2_D_REG_22__SCAN_IN), .B0(n5751), .Y(n5830));
  NAND3X1 g4705(.A(n5830), .B(n5829), .C(n5828), .Y(n5831));
  OAI21X1 g4706(.A0(P2_D_REG_14__SCAN_IN), .A1(P2_D_REG_12__SCAN_IN), .B0(n5751), .Y(n5832));
  OAI21X1 g4707(.A0(P2_D_REG_13__SCAN_IN), .A1(P2_D_REG_11__SCAN_IN), .B0(n5751), .Y(n5833));
  OAI21X1 g4708(.A0(P2_D_REG_24__SCAN_IN), .A1(P2_D_REG_16__SCAN_IN), .B0(n5751), .Y(n5834));
  OAI21X1 g4709(.A0(P2_D_REG_17__SCAN_IN), .A1(P2_D_REG_15__SCAN_IN), .B0(n5751), .Y(n5835));
  NAND4X1 g4710(.A(n5834), .B(n5833), .C(n5832), .D(n5835), .Y(n5836));
  NOR4X1  g4711(.A(n5831), .B(n5827), .C(n5822), .D(n5836), .Y(n5837));
  INVX1   g4712(.A(P2_D_REG_1__SCAN_IN), .Y(n5838));
  NOR2X1  g4713(.A(n5747), .B(n5838), .Y(n5839));
  AOI21X1 g4714(.A0(n5754), .A1(n5747), .B0(n5839), .Y(n5840));
  INVX1   g4715(.A(n5840), .Y(n5841));
  NAND2X1 g4716(.A(n5470), .B(P2_IR_REG_22__SCAN_IN), .Y(n5842));
  OAI21X1 g4717(.A0(n5650), .A1(n5470), .B0(n5842), .Y(n5843));
  INVX1   g4718(.A(P2_IR_REG_21__SCAN_IN), .Y(n5844));
  NOR2X1  g4719(.A(P2_IR_REG_31__SCAN_IN), .B(n5844), .Y(n5845));
  INVX1   g4720(.A(n5845), .Y(n5846));
  OAI21X1 g4721(.A0(n5637), .A1(n5470), .B0(n5846), .Y(n5847));
  INVX1   g4722(.A(n5847), .Y(n5848));
  XOR2X1  g4723(.A(n5848), .B(n5843), .Y(n5849));
  INVX1   g4724(.A(n5843), .Y(n5850));
  NOR2X1  g4725(.A(P2_IR_REG_31__SCAN_IN), .B(n5625), .Y(n5851));
  AOI21X1 g4726(.A0(n5628), .A1(P2_IR_REG_31__SCAN_IN), .B0(n5851), .Y(n5852));
  INVX1   g4727(.A(n5852), .Y(n5853));
  NOR2X1  g4728(.A(P2_IR_REG_31__SCAN_IN), .B(n5645), .Y(n5854));
  AOI21X1 g4729(.A0(n5619), .A1(P2_IR_REG_31__SCAN_IN), .B0(n5854), .Y(n5855));
  INVX1   g4730(.A(n5855), .Y(n5856));
  NOR2X1  g4731(.A(n5856), .B(n5853), .Y(n5857));
  AOI21X1 g4732(.A0(n5853), .A1(n5850), .B0(n5857), .Y(n5858));
  AOI21X1 g4733(.A0(n5858), .A1(n5849), .B0(n5841), .Y(n5859));
  AOI21X1 g4734(.A0(n5739), .A1(n5737), .B0(n5751), .Y(n5860));
  AOI21X1 g4735(.A0(n5751), .A1(P2_D_REG_0__SCAN_IN), .B0(n5860), .Y(n5861));
  NAND4X1 g4736(.A(n5859), .B(n5837), .C(n5743), .D(n5861), .Y(n5862));
  NAND2X1 g4737(.A(n5699), .B(P2_IR_REG_31__SCAN_IN), .Y(n5863));
  OAI21X1 g4738(.A0(P2_IR_REG_31__SCAN_IN), .A1(n5696), .B0(n5863), .Y(n5864));
  NAND2X1 g4739(.A(n5707), .B(P2_IR_REG_31__SCAN_IN), .Y(n5865));
  OAI21X1 g4740(.A0(P2_IR_REG_31__SCAN_IN), .A1(n5705), .B0(n5865), .Y(n5866));
  NOR2X1  g4741(.A(n5866), .B(n5864), .Y(n5867));
  NOR2X1  g4742(.A(P2_IR_REG_31__SCAN_IN), .B(n5696), .Y(n5868));
  AOI21X1 g4743(.A0(n5699), .A1(P2_IR_REG_31__SCAN_IN), .B0(n5868), .Y(n5869));
  NOR2X1  g4744(.A(P2_IR_REG_31__SCAN_IN), .B(n5705), .Y(n5870));
  AOI21X1 g4745(.A0(n5707), .A1(P2_IR_REG_31__SCAN_IN), .B0(n5870), .Y(n5871));
  INVX1   g4746(.A(n5477), .Y(n5875));
  NAND3X1 g4747(.A(n5875), .B(n5871), .C(n5869), .Y(n5876));
  OAI21X1 g4748(.A0(n5867), .A1(n5463), .B0(n5876), .Y(n5877));
  INVX1   g4749(.A(P2_REG1_REG_0__SCAN_IN), .Y(n5878));
  INVX1   g4750(.A(P2_REG2_REG_0__SCAN_IN), .Y(n5879));
  NOR2X1  g4751(.A(P2_IR_REG_31__SCAN_IN), .B(n5713), .Y(n5880));
  AOI21X1 g4752(.A0(n5715), .A1(P2_IR_REG_31__SCAN_IN), .B0(n5880), .Y(n5881));
  INVX1   g4753(.A(P2_IR_REG_30__SCAN_IN), .Y(n5882));
  XOR2X1  g4754(.A(n5722), .B(n5882), .Y(n5883));
  NOR2X1  g4755(.A(P2_IR_REG_31__SCAN_IN), .B(n5882), .Y(n5884));
  INVX1   g4756(.A(n5884), .Y(n5885));
  OAI21X1 g4757(.A0(n5883), .A1(n5470), .B0(n5885), .Y(n5886));
  NAND2X1 g4758(.A(n5886), .B(n5881), .Y(n5887));
  NAND2X1 g4759(.A(n5715), .B(P2_IR_REG_31__SCAN_IN), .Y(n5888));
  OAI21X1 g4760(.A0(P2_IR_REG_31__SCAN_IN), .A1(n5713), .B0(n5888), .Y(n5889));
  AOI21X1 g4761(.A0(n5723), .A1(P2_IR_REG_31__SCAN_IN), .B0(n5884), .Y(n5890));
  NAND2X1 g4762(.A(n5890), .B(n5889), .Y(n5891));
  OAI22X1 g4763(.A0(n5887), .A1(n5879), .B0(n5878), .B1(n5891), .Y(n5892));
  INVX1   g4764(.A(P2_REG3_REG_0__SCAN_IN), .Y(n5893));
  NAND2X1 g4765(.A(n5886), .B(n5889), .Y(n5894));
  NAND3X1 g4766(.A(n5890), .B(n5881), .C(P2_REG0_REG_0__SCAN_IN), .Y(n5895));
  OAI21X1 g4767(.A0(n5894), .A1(n5893), .B0(n5895), .Y(n5896));
  NOR2X1  g4768(.A(n5896), .B(n5892), .Y(n5897));
  XOR2X1  g4769(.A(n5897), .B(n5877), .Y(n5898));
  NOR3X1  g4770(.A(n5855), .B(n5853), .C(n5850), .Y(n5900));
  NOR3X1  g4771(.A(n5855), .B(n5852), .C(n5848), .Y(n5901));
  INVX1   g4772(.A(n5901), .Y(n5902));
  NOR3X1  g4773(.A(n5856), .B(n5852), .C(n5850), .Y(n5903));
  INVX1   g4774(.A(n5903), .Y(n5904));
  AOI21X1 g4775(.A0(n5904), .A1(n5902), .B0(n5898), .Y(n5905));
  AOI21X1 g4776(.A0(n5900), .A1(n8912), .B0(n5905), .Y(n5906));
  NOR3X1  g4777(.A(n5855), .B(n5852), .C(n5850), .Y(n5907));
  NOR3X1  g4778(.A(n5856), .B(n5852), .C(n5848), .Y(n5908));
  OAI21X1 g4779(.A0(n5908), .A1(n5907), .B0(n8912), .Y(n5909));
  NOR4X1  g4780(.A(n5853), .B(n5848), .C(n5843), .D(n5856), .Y(n5910));
  NOR4X1  g4781(.A(n5853), .B(n5847), .C(n5850), .D(n5856), .Y(n5911));
  OAI21X1 g4782(.A0(n5911), .A1(n5910), .B0(n8912), .Y(n5912));
  NAND3X1 g4783(.A(n5912), .B(n5909), .C(n5906), .Y(n5913));
  NAND3X1 g4784(.A(n5856), .B(n5852), .C(n5850), .Y(n5914));
  NOR3X1  g4785(.A(n5866), .B(n5848), .C(n5850), .Y(n5915));
  NOR2X1  g4786(.A(n5890), .B(n5889), .Y(n5916));
  NOR2X1  g4787(.A(n5886), .B(n5881), .Y(n5917));
  AOI22X1 g4788(.A0(n5916), .A1(P2_REG2_REG_1__SCAN_IN), .B0(P2_REG1_REG_1__SCAN_IN), .B1(n5917), .Y(n5918));
  NOR2X1  g4789(.A(n5890), .B(n5881), .Y(n5919));
  NOR2X1  g4790(.A(n5886), .B(n5889), .Y(n5920));
  AOI22X1 g4791(.A0(n5919), .A1(P2_REG3_REG_1__SCAN_IN), .B0(P2_REG0_REG_1__SCAN_IN), .B1(n5920), .Y(n5921));
  NAND2X1 g4792(.A(n5921), .B(n5918), .Y(n5922));
  INVX1   g4793(.A(n5877), .Y(n5923));
  NOR3X1  g4794(.A(n5853), .B(n5847), .C(n5843), .Y(n5924));
  INVX1   g4795(.A(n5924), .Y(n5925));
  NOR2X1  g4796(.A(n5847), .B(n5843), .Y(n5926));
  NOR3X1  g4797(.A(n5856), .B(n5852), .C(n5847), .Y(n5927));
  AOI22X1 g4798(.A0(n5926), .A1(n5856), .B0(n5850), .B1(n5927), .Y(n5928));
  AOI21X1 g4799(.A0(n5928), .A1(n5925), .B0(n5923), .Y(n5929));
  AOI21X1 g4800(.A0(n5922), .A1(n5915), .B0(n5929), .Y(n5930));
  OAI21X1 g4801(.A0(n5914), .A1(n5898), .B0(n5930), .Y(n5931));
  NOR2X1  g4802(.A(n5931), .B(n5913), .Y(n5932));
  NAND2X1 g4803(.A(n5862), .B(P2_REG0_REG_0__SCAN_IN), .Y(n5933));
  OAI21X1 g4804(.A0(n5932), .A1(n5862), .B0(n5933), .Y(P2_U3451));
  NOR2X1  g4805(.A(P2_IR_REG_31__SCAN_IN), .B(n5478), .Y(n5935));
  AOI21X1 g4806(.A0(n5472), .A1(P2_IR_REG_31__SCAN_IN), .B0(n5935), .Y(n5936));
  INVX1   g4807(.A(n5936), .Y(n5937));
  NAND3X1 g4808(.A(n5937), .B(n5871), .C(n5869), .Y(n5938));
  OAI21X1 g4809(.A0(n5867), .A1(n5467), .B0(n5938), .Y(n5939));
  XOR2X1  g4810(.A(n5939), .B(n5922), .Y(n5940));
  OAI21X1 g4811(.A0(n5896), .A1(n5892), .B0(n5877), .Y(n5941));
  XOR2X1  g4812(.A(n5941), .B(n5940), .Y(n5942));
  INVX1   g4813(.A(n5942), .Y(n5943));
  OAI21X1 g4814(.A0(n5911), .A1(n5903), .B0(n5943), .Y(n5944));
  AOI22X1 g4815(.A0(n5916), .A1(P2_REG2_REG_0__SCAN_IN), .B0(P2_REG1_REG_0__SCAN_IN), .B1(n5917), .Y(n5945));
  AOI22X1 g4816(.A0(n5919), .A1(P2_REG3_REG_0__SCAN_IN), .B0(P2_REG0_REG_0__SCAN_IN), .B1(n5920), .Y(n5946));
  NAND3X1 g4817(.A(n5946), .B(n5945), .C(n5877), .Y(n5947));
  INVX1   g4818(.A(P2_REG1_REG_1__SCAN_IN), .Y(n5948));
  INVX1   g4819(.A(P2_REG2_REG_1__SCAN_IN), .Y(n5949));
  OAI22X1 g4820(.A0(n5887), .A1(n5949), .B0(n5948), .B1(n5891), .Y(n5950));
  INVX1   g4821(.A(P2_REG3_REG_1__SCAN_IN), .Y(n5951));
  NAND3X1 g4822(.A(n5890), .B(n5881), .C(P2_REG0_REG_1__SCAN_IN), .Y(n5952));
  OAI21X1 g4823(.A0(n5894), .A1(n5951), .B0(n5952), .Y(n5953));
  NOR2X1  g4824(.A(n5953), .B(n5950), .Y(n5954));
  XOR2X1  g4825(.A(n5939), .B(n5954), .Y(n5955));
  XOR2X1  g4826(.A(n5955), .B(n5947), .Y(n5956));
  AOI22X1 g4827(.A0(n5943), .A1(n5910), .B0(n5901), .B1(n5956), .Y(n5957));
  INVX1   g4828(.A(n5897), .Y(n5958));
  NOR3X1  g4829(.A(n5871), .B(n5848), .C(n5850), .Y(n5959));
  AOI22X1 g4830(.A0(n5956), .A1(n5908), .B0(n5958), .B1(n5959), .Y(n5960));
  OAI21X1 g4831(.A0(n5907), .A1(n5900), .B0(n5956), .Y(n5961));
  NAND4X1 g4832(.A(n5960), .B(n5957), .C(n5944), .D(n5961), .Y(n5962));
  XOR2X1  g4833(.A(n5939), .B(n5923), .Y(n5963));
  INVX1   g4834(.A(n5963), .Y(n5964));
  INVX1   g4835(.A(n5915), .Y(n5965));
  NOR2X1  g4836(.A(n5867), .B(n5467), .Y(n5966));
  AOI21X1 g4837(.A0(n5937), .A1(n5867), .B0(n5966), .Y(n5967));
  INVX1   g4838(.A(P2_REG1_REG_2__SCAN_IN), .Y(n5968));
  INVX1   g4839(.A(P2_REG2_REG_2__SCAN_IN), .Y(n5969));
  OAI22X1 g4840(.A0(n5887), .A1(n5969), .B0(n5968), .B1(n5891), .Y(n5970));
  INVX1   g4841(.A(P2_REG3_REG_2__SCAN_IN), .Y(n5971));
  NAND3X1 g4842(.A(n5890), .B(n5881), .C(P2_REG0_REG_2__SCAN_IN), .Y(n5972));
  OAI21X1 g4843(.A0(n5894), .A1(n5971), .B0(n5972), .Y(n5973));
  NOR2X1  g4844(.A(n5973), .B(n5970), .Y(n5974));
  OAI22X1 g4845(.A0(n5967), .A1(n5928), .B0(n5965), .B1(n5974), .Y(n5975));
  AOI21X1 g4846(.A0(n5964), .A1(n5924), .B0(n5975), .Y(n5976));
  OAI21X1 g4847(.A0(n5942), .A1(n5914), .B0(n5976), .Y(n5977));
  NOR2X1  g4848(.A(n5977), .B(n5962), .Y(n5978));
  NAND2X1 g4849(.A(n5862), .B(P2_REG0_REG_1__SCAN_IN), .Y(n5979));
  OAI21X1 g4850(.A0(n5978), .A1(n5862), .B0(n5979), .Y(P2_U3454));
  NOR2X1  g4851(.A(n5967), .B(n5954), .Y(n5981));
  AOI21X1 g4852(.A0(n5967), .A1(n5954), .B0(n5941), .Y(n5982));
  NOR2X1  g4853(.A(n5982), .B(n5981), .Y(n5983));
  AOI22X1 g4854(.A0(n5916), .A1(P2_REG2_REG_2__SCAN_IN), .B0(P2_REG1_REG_2__SCAN_IN), .B1(n5917), .Y(n5984));
  AOI22X1 g4855(.A0(n5919), .A1(P2_REG3_REG_2__SCAN_IN), .B0(P2_REG0_REG_2__SCAN_IN), .B1(n5920), .Y(n5985));
  NOR2X1  g4856(.A(P2_IR_REG_31__SCAN_IN), .B(n5600), .Y(n5986));
  AOI21X1 g4857(.A0(n5480), .A1(P2_IR_REG_31__SCAN_IN), .B0(n5986), .Y(n5987));
  INVX1   g4858(.A(n5987), .Y(n5988));
  AOI21X1 g4859(.A0(n5871), .A1(n5869), .B0(n5476), .Y(n5989));
  AOI21X1 g4860(.A0(n5988), .A1(n5867), .B0(n5989), .Y(n5990));
  AOI21X1 g4861(.A0(n5985), .A1(n5984), .B0(n5990), .Y(n5991));
  NAND3X1 g4862(.A(n5990), .B(n5985), .C(n5984), .Y(n5992));
  INVX1   g4863(.A(n5992), .Y(n5993));
  NOR3X1  g4864(.A(n5983), .B(n5993), .C(n5991), .Y(n5994));
  NAND2X1 g4865(.A(n5985), .B(n5984), .Y(n5995));
  XOR2X1  g4866(.A(n5990), .B(n5995), .Y(n5996));
  AOI21X1 g4867(.A0(n5996), .A1(n5983), .B0(n5994), .Y(n5997));
  AOI22X1 g4868(.A0(n5959), .A1(n5922), .B0(n5910), .B1(n5997), .Y(n5998));
  OAI21X1 g4869(.A0(n5911), .A1(n5903), .B0(n5997), .Y(n5999));
  NAND2X1 g4870(.A(n5922), .B(n5947), .Y(n6000));
  OAI21X1 g4871(.A0(n5922), .A1(n5947), .B0(n5967), .Y(n6001));
  NAND2X1 g4872(.A(n6001), .B(n6000), .Y(n6002));
  XOR2X1  g4873(.A(n6002), .B(n5996), .Y(n6003));
  OAI21X1 g4874(.A0(n5908), .A1(n5907), .B0(n6003), .Y(n6004));
  OAI21X1 g4875(.A0(n5901), .A1(n5900), .B0(n6003), .Y(n6005));
  NAND4X1 g4876(.A(n6004), .B(n5999), .C(n5998), .D(n6005), .Y(n6006));
  NAND4X1 g4877(.A(n5856), .B(n5852), .C(n5850), .D(n5997), .Y(n6007));
  NOR2X1  g4878(.A(n5939), .B(n5877), .Y(n6008));
  XOR2X1  g4879(.A(n6008), .B(n5990), .Y(n6009));
  INVX1   g4880(.A(P2_REG2_REG_3__SCAN_IN), .Y(n6010));
  NAND3X1 g4881(.A(n5890), .B(n5881), .C(P2_REG0_REG_3__SCAN_IN), .Y(n6011));
  OAI21X1 g4882(.A0(n5887), .A1(n6010), .B0(n6011), .Y(n6012));
  INVX1   g4883(.A(P2_REG1_REG_3__SCAN_IN), .Y(n6013));
  OAI22X1 g4884(.A0(n5891), .A1(n6013), .B0(P2_REG3_REG_3__SCAN_IN), .B1(n5894), .Y(n6014));
  NOR2X1  g4885(.A(n6014), .B(n6012), .Y(n6015));
  OAI22X1 g4886(.A0(n5990), .A1(n5928), .B0(n5965), .B1(n6015), .Y(n6016));
  AOI21X1 g4887(.A0(n6009), .A1(n5924), .B0(n6016), .Y(n6017));
  NAND2X1 g4888(.A(n6017), .B(n6007), .Y(n6018));
  NOR2X1  g4889(.A(n6018), .B(n6006), .Y(n6019));
  NAND2X1 g4890(.A(n5862), .B(P2_REG0_REG_2__SCAN_IN), .Y(n6020));
  OAI21X1 g4891(.A0(n6019), .A1(n5862), .B0(n6020), .Y(P2_U3457));
  AOI21X1 g4892(.A0(n5992), .A1(n5981), .B0(n5991), .Y(n6022));
  INVX1   g4893(.A(n6022), .Y(n6023));
  AOI21X1 g4894(.A0(n5982), .A1(n5992), .B0(n6023), .Y(n6024));
  AOI22X1 g4895(.A0(n5916), .A1(P2_REG2_REG_3__SCAN_IN), .B0(P2_REG0_REG_3__SCAN_IN), .B1(n5920), .Y(n6025));
  INVX1   g4896(.A(P2_REG3_REG_3__SCAN_IN), .Y(n6026));
  AOI22X1 g4897(.A0(n5917), .A1(P2_REG1_REG_3__SCAN_IN), .B0(n6026), .B1(n5919), .Y(n6027));
  NAND2X1 g4898(.A(n6027), .B(n6025), .Y(n6028));
  NOR2X1  g4899(.A(P2_IR_REG_31__SCAN_IN), .B(n5485), .Y(n6029));
  AOI21X1 g4900(.A0(n5487), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6029), .Y(n6030));
  INVX1   g4901(.A(n6030), .Y(n6031));
  NAND3X1 g4902(.A(n6031), .B(n5871), .C(n5869), .Y(n6032));
  OAI21X1 g4903(.A0(n5867), .A1(n5484), .B0(n6032), .Y(n6033));
  INVX1   g4904(.A(n6033), .Y(n6034));
  XOR2X1  g4905(.A(n6034), .B(n6028), .Y(n6035));
  XOR2X1  g4906(.A(n6034), .B(n6015), .Y(n6037));
  NOR2X1  g4907(.A(n6037), .B(n6024), .Y(n6038));
  AOI21X1 g4908(.A0(n6037), .A1(n6024), .B0(n6038), .Y(n6039));
  INVX1   g4909(.A(n6039), .Y(n6040));
  AOI22X1 g4910(.A0(n5995), .A1(n5959), .B0(n5910), .B1(n6040), .Y(n6041));
  OAI21X1 g4911(.A0(n5911), .A1(n5903), .B0(n6040), .Y(n6042));
  NOR3X1  g4912(.A(n5990), .B(n5973), .C(n5970), .Y(n6043));
  AOI21X1 g4913(.A0(n5921), .A1(n5918), .B0(n5939), .Y(n6044));
  NAND3X1 g4914(.A(n5988), .B(n5871), .C(n5869), .Y(n6045));
  OAI21X1 g4915(.A0(n5867), .A1(n5476), .B0(n6045), .Y(n6046));
  AOI21X1 g4916(.A0(n5985), .A1(n5984), .B0(n6046), .Y(n6047));
  AOI21X1 g4917(.A0(n5897), .A1(n5877), .B0(n5954), .Y(n6048));
  AOI21X1 g4918(.A0(n5897), .A1(n5877), .B0(n5939), .Y(n6049));
  NOR4X1  g4919(.A(n6048), .B(n6047), .C(n6044), .D(n6049), .Y(n6050));
  NOR3X1  g4920(.A(n6050), .B(n6035), .C(n6043), .Y(n6051));
  AOI21X1 g4921(.A0(n6001), .A1(n6000), .B0(n6043), .Y(n6052));
  NOR3X1  g4922(.A(n6052), .B(n6037), .C(n6047), .Y(n6053));
  OAI22X1 g4923(.A0(n6051), .A1(n6053), .B0(n5908), .B1(n5907), .Y(n6054));
  OAI22X1 g4924(.A0(n6051), .A1(n6053), .B0(n5901), .B1(n5900), .Y(n6055));
  NAND4X1 g4925(.A(n6054), .B(n6042), .C(n6041), .D(n6055), .Y(n6056));
  NOR2X1  g4926(.A(n6039), .B(n5914), .Y(n6057));
  NOR3X1  g4927(.A(n6046), .B(n5939), .C(n5877), .Y(n6058));
  XOR2X1  g4928(.A(n6033), .B(n6058), .Y(n6059));
  INVX1   g4929(.A(n5928), .Y(n6060));
  AOI22X1 g4930(.A0(n5916), .A1(P2_REG2_REG_4__SCAN_IN), .B0(P2_REG0_REG_4__SCAN_IN), .B1(n5920), .Y(n6061));
  XOR2X1  g4931(.A(P2_REG3_REG_4__SCAN_IN), .B(n6026), .Y(n6062));
  INVX1   g4932(.A(n6062), .Y(n6063));
  AOI22X1 g4933(.A0(n5919), .A1(n6063), .B0(n5917), .B1(P2_REG1_REG_4__SCAN_IN), .Y(n6064));
  NAND2X1 g4934(.A(n6064), .B(n6061), .Y(n6065));
  AOI22X1 g4935(.A0(n6033), .A1(n6060), .B0(n5915), .B1(n6065), .Y(n6066));
  OAI21X1 g4936(.A0(n6059), .A1(n5925), .B0(n6066), .Y(n6067));
  NOR3X1  g4937(.A(n6067), .B(n6057), .C(n6056), .Y(n6068));
  NAND2X1 g4938(.A(n5862), .B(P2_REG0_REG_3__SCAN_IN), .Y(n6069));
  OAI21X1 g4939(.A0(n6068), .A1(n5862), .B0(n6069), .Y(P2_U3460));
  INVX1   g4940(.A(n5910), .Y(n6071));
  INVX1   g4941(.A(n5959), .Y(n6072));
  NOR2X1  g4942(.A(P2_IR_REG_31__SCAN_IN), .B(n5492), .Y(n6073));
  AOI21X1 g4943(.A0(n5494), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6073), .Y(n6074));
  INVX1   g4944(.A(n6074), .Y(n6075));
  NOR2X1  g4945(.A(n5867), .B(n5491), .Y(n6076));
  AOI21X1 g4946(.A0(n6075), .A1(n5867), .B0(n6076), .Y(n6077));
  NOR2X1  g4947(.A(n6034), .B(n6015), .Y(n6080));
  NAND2X1 g4948(.A(n6034), .B(n6015), .Y(n6081));
  INVX1   g4949(.A(n6081), .Y(n6082));
  NOR2X1  g4950(.A(n6082), .B(n6022), .Y(n6083));
  INVX1   g4951(.A(n5982), .Y(n6084));
  NOR3X1  g4952(.A(n6082), .B(n6084), .C(n5993), .Y(n6085));
  NOR3X1  g4953(.A(n6085), .B(n6083), .C(n6080), .Y(n6086));
  INVX1   g4954(.A(P2_REG2_REG_4__SCAN_IN), .Y(n6087));
  NAND3X1 g4955(.A(n5890), .B(n5881), .C(P2_REG0_REG_4__SCAN_IN), .Y(n6088));
  OAI21X1 g4956(.A0(n5887), .A1(n6087), .B0(n6088), .Y(n6089));
  INVX1   g4957(.A(P2_REG1_REG_4__SCAN_IN), .Y(n6090));
  OAI22X1 g4958(.A0(n5894), .A1(n6062), .B0(n5891), .B1(n6090), .Y(n6091));
  NOR2X1  g4959(.A(n6091), .B(n6089), .Y(n6092));
  XOR2X1  g4960(.A(n6077), .B(n6092), .Y(n6093));
  NOR2X1  g4961(.A(n6093), .B(n6086), .Y(n6094));
  AOI21X1 g4962(.A0(n6086), .A1(n6093), .B0(n6094), .Y(n6095));
  OAI22X1 g4963(.A0(n6015), .A1(n6072), .B0(n6071), .B1(n6095), .Y(n6096));
  INVX1   g4964(.A(n5911), .Y(n6097));
  AOI21X1 g4965(.A0(n6097), .A1(n5904), .B0(n6095), .Y(n6098));
  NOR3X1  g4966(.A(n6049), .B(n6048), .C(n6044), .Y(n6099));
  OAI22X1 g4967(.A0(n6028), .A1(n6034), .B0(n5990), .B1(n5995), .Y(n6100));
  OAI21X1 g4968(.A0(n6046), .A1(n5974), .B0(n6015), .Y(n6101));
  NOR3X1  g4969(.A(n6015), .B(n6046), .C(n5974), .Y(n6102));
  AOI21X1 g4970(.A0(n6101), .A1(n6034), .B0(n6102), .Y(n6103));
  OAI21X1 g4971(.A0(n6100), .A1(n6099), .B0(n6103), .Y(n6104));
  XOR2X1  g4972(.A(n6104), .B(n6093), .Y(n6105));
  INVX1   g4973(.A(n6105), .Y(n6106));
  OAI21X1 g4974(.A0(n5908), .A1(n5907), .B0(n6106), .Y(n6107));
  OAI21X1 g4975(.A0(n5901), .A1(n5900), .B0(n6106), .Y(n6108));
  NAND2X1 g4976(.A(n6108), .B(n6107), .Y(n6109));
  NAND2X1 g4977(.A(n6034), .B(n6058), .Y(n6110));
  NAND3X1 g4978(.A(n6075), .B(n5871), .C(n5869), .Y(n6111));
  OAI21X1 g4979(.A0(n5867), .A1(n5491), .B0(n6111), .Y(n6112));
  XOR2X1  g4980(.A(n6112), .B(n6110), .Y(n6113));
  INVX1   g4981(.A(P2_REG2_REG_5__SCAN_IN), .Y(n6114));
  NAND3X1 g4982(.A(n5890), .B(n5881), .C(P2_REG0_REG_5__SCAN_IN), .Y(n6115));
  OAI21X1 g4983(.A0(n5887), .A1(n6114), .B0(n6115), .Y(n6116));
  INVX1   g4984(.A(P2_REG1_REG_5__SCAN_IN), .Y(n6117));
  NAND2X1 g4985(.A(P2_REG3_REG_4__SCAN_IN), .B(P2_REG3_REG_3__SCAN_IN), .Y(n6118));
  XOR2X1  g4986(.A(n6118), .B(P2_REG3_REG_5__SCAN_IN), .Y(n6119));
  OAI22X1 g4987(.A0(n5894), .A1(n6119), .B0(n5891), .B1(n6117), .Y(n6120));
  NOR2X1  g4988(.A(n6120), .B(n6116), .Y(n6121));
  OAI22X1 g4989(.A0(n6077), .A1(n5928), .B0(n5965), .B1(n6121), .Y(n6122));
  AOI21X1 g4990(.A0(n6113), .A1(n5924), .B0(n6122), .Y(n6123));
  OAI21X1 g4991(.A0(n6095), .A1(n5914), .B0(n6123), .Y(n6124));
  NOR4X1  g4992(.A(n6109), .B(n6098), .C(n6096), .D(n6124), .Y(n6125));
  NAND2X1 g4993(.A(n5862), .B(P2_REG0_REG_4__SCAN_IN), .Y(n6126));
  OAI21X1 g4994(.A0(n6125), .A1(n5862), .B0(n6126), .Y(P2_U3463));
  INVX1   g4995(.A(n5908), .Y(n6128));
  NOR2X1  g4996(.A(P2_IR_REG_31__SCAN_IN), .B(n5505), .Y(n6129));
  AOI21X1 g4997(.A0(n5500), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6129), .Y(n6130));
  NOR3X1  g4998(.A(n6130), .B(n5866), .C(n5864), .Y(n6131));
  INVX1   g4999(.A(n6131), .Y(n6132));
  OAI21X1 g5000(.A0(n5867), .A1(n5498), .B0(n6132), .Y(n6133));
  XOR2X1  g5001(.A(n6133), .B(n6121), .Y(n6134));
  NAND3X1 g5002(.A(n6112), .B(n6064), .C(n6061), .Y(n6135));
  AOI21X1 g5003(.A0(n6064), .A1(n6061), .B0(n6112), .Y(n6136));
  AOI21X1 g5004(.A0(n6104), .A1(n6135), .B0(n6136), .Y(n6137));
  XOR2X1  g5005(.A(n6137), .B(n6134), .Y(n6138));
  NOR2X1  g5006(.A(n6138), .B(n6128), .Y(n6139));
  NOR2X1  g5007(.A(n6077), .B(n6092), .Y(n6140));
  NOR4X1  g5008(.A(n6085), .B(n6083), .C(n6080), .D(n6140), .Y(n6141));
  INVX1   g5009(.A(n6133), .Y(n6142));
  AOI22X1 g5010(.A0(n5916), .A1(P2_REG2_REG_5__SCAN_IN), .B0(P2_REG0_REG_5__SCAN_IN), .B1(n5920), .Y(n6143));
  INVX1   g5011(.A(n6119), .Y(n6144));
  AOI22X1 g5012(.A0(n5919), .A1(n6144), .B0(n5917), .B1(P2_REG1_REG_5__SCAN_IN), .Y(n6145));
  NAND2X1 g5013(.A(n6145), .B(n6143), .Y(n6146));
  OAI22X1 g5014(.A0(n6146), .A1(n6133), .B0(n6112), .B1(n6065), .Y(n6147));
  INVX1   g5015(.A(n6147), .Y(n6148));
  OAI21X1 g5016(.A0(n6142), .A1(n6121), .B0(n6148), .Y(n6149));
  AOI21X1 g5017(.A0(n6077), .A1(n6092), .B0(n6086), .Y(n6150));
  OAI21X1 g5018(.A0(n6091), .A1(n6089), .B0(n6112), .Y(n6151));
  NAND2X1 g5019(.A(n6134), .B(n6151), .Y(n6152));
  OAI22X1 g5020(.A0(n6150), .A1(n6152), .B0(n6149), .B1(n6141), .Y(n6153));
  OAI22X1 g5021(.A0(n6092), .A1(n6072), .B0(n6071), .B1(n6153), .Y(n6154));
  AOI21X1 g5022(.A0(n6097), .A1(n5904), .B0(n6153), .Y(n6155));
  INVX1   g5023(.A(n6138), .Y(n6156));
  OAI21X1 g5024(.A0(n5907), .A1(n5900), .B0(n6156), .Y(n6157));
  OAI21X1 g5025(.A0(n6138), .A1(n5902), .B0(n6157), .Y(n6158));
  NOR4X1  g5026(.A(n6155), .B(n6154), .C(n6139), .D(n6158), .Y(n6159));
  INVX1   g5027(.A(n6159), .Y(n6160));
  NOR2X1  g5028(.A(n6112), .B(n6110), .Y(n6161));
  XOR2X1  g5029(.A(n6142), .B(n6161), .Y(n6162));
  INVX1   g5030(.A(P2_REG2_REG_6__SCAN_IN), .Y(n6163));
  NAND3X1 g5031(.A(n5890), .B(n5881), .C(P2_REG0_REG_6__SCAN_IN), .Y(n6164));
  OAI21X1 g5032(.A0(n5887), .A1(n6163), .B0(n6164), .Y(n6165));
  NAND3X1 g5033(.A(n5890), .B(n5889), .C(P2_REG1_REG_6__SCAN_IN), .Y(n6166));
  NAND3X1 g5034(.A(P2_REG3_REG_4__SCAN_IN), .B(P2_REG3_REG_5__SCAN_IN), .C(P2_REG3_REG_3__SCAN_IN), .Y(n6167));
  XOR2X1  g5035(.A(n6167), .B(P2_REG3_REG_6__SCAN_IN), .Y(n6168));
  INVX1   g5036(.A(n6168), .Y(n6169));
  NAND3X1 g5037(.A(n6169), .B(n5886), .C(n5889), .Y(n6170));
  NAND2X1 g5038(.A(n6170), .B(n6166), .Y(n6171));
  NOR2X1  g5039(.A(n6171), .B(n6165), .Y(n6172));
  OAI22X1 g5040(.A0(n6142), .A1(n5928), .B0(n5965), .B1(n6172), .Y(n6173));
  AOI21X1 g5041(.A0(n6162), .A1(n5924), .B0(n6173), .Y(n6174));
  OAI21X1 g5042(.A0(n6153), .A1(n5914), .B0(n6174), .Y(n6175));
  NOR2X1  g5043(.A(n6175), .B(n6160), .Y(n6176));
  NAND2X1 g5044(.A(n5862), .B(P2_REG0_REG_5__SCAN_IN), .Y(n6177));
  OAI21X1 g5045(.A0(n6176), .A1(n5862), .B0(n6177), .Y(P2_U3466));
  INVX1   g5046(.A(n6137), .Y(n6179));
  AOI21X1 g5047(.A0(n6142), .A1(n6146), .B0(n6179), .Y(n6180));
  NOR2X1  g5048(.A(P2_IR_REG_31__SCAN_IN), .B(n5507), .Y(n6181));
  AOI21X1 g5049(.A0(n5510), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6181), .Y(n6182));
  INVX1   g5050(.A(n6182), .Y(n6183));
  NAND3X1 g5051(.A(n6183), .B(n5871), .C(n5869), .Y(n6184));
  OAI21X1 g5052(.A0(n5867), .A1(n5504), .B0(n6184), .Y(n6185));
  XOR2X1  g5053(.A(n6185), .B(n6172), .Y(n6186));
  AOI21X1 g5054(.A0(n6133), .A1(n6121), .B0(n6186), .Y(n6187));
  INVX1   g5055(.A(n6187), .Y(n6188));
  NOR2X1  g5056(.A(n6142), .B(n6146), .Y(n6189));
  OAI22X1 g5057(.A0(n6172), .A1(n6185), .B0(n6133), .B1(n6121), .Y(n6190));
  AOI21X1 g5058(.A0(n6185), .A1(n6172), .B0(n6190), .Y(n6191));
  OAI21X1 g5059(.A0(n6137), .A1(n6189), .B0(n6191), .Y(n6192));
  OAI21X1 g5060(.A0(n6188), .A1(n6180), .B0(n6192), .Y(n6193));
  INVX1   g5061(.A(n6193), .Y(n6194));
  NOR2X1  g5062(.A(n6194), .B(n6128), .Y(n6195));
  AOI21X1 g5063(.A0(n6033), .A1(n6028), .B0(n5991), .Y(n6196));
  OAI21X1 g5064(.A0(n5983), .A1(n5993), .B0(n6196), .Y(n6197));
  AOI21X1 g5065(.A0(n6034), .A1(n6015), .B0(n6147), .Y(n6198));
  NAND3X1 g5066(.A(n6133), .B(n6112), .C(n6065), .Y(n6199));
  OAI21X1 g5067(.A0(n6133), .A1(n6140), .B0(n6146), .Y(n6200));
  NAND2X1 g5068(.A(n6200), .B(n6199), .Y(n6201));
  AOI21X1 g5069(.A0(n6198), .A1(n6197), .B0(n6201), .Y(n6202));
  INVX1   g5070(.A(n6202), .Y(n6203));
  NOR2X1  g5071(.A(n6203), .B(n6186), .Y(n6204));
  AOI21X1 g5072(.A0(n6186), .A1(n6203), .B0(n6204), .Y(n6206));
  OAI22X1 g5073(.A0(n6121), .A1(n6072), .B0(n6071), .B1(n6206), .Y(n6207));
  AOI21X1 g5074(.A0(n6097), .A1(n5904), .B0(n6206), .Y(n6208));
  OAI21X1 g5075(.A0(n5907), .A1(n5900), .B0(n6193), .Y(n6209));
  OAI21X1 g5076(.A0(n6194), .A1(n5902), .B0(n6209), .Y(n6210));
  NOR4X1  g5077(.A(n6208), .B(n6207), .C(n6195), .D(n6210), .Y(n6211));
  INVX1   g5078(.A(n6211), .Y(n6212));
  NAND4X1 g5079(.A(n6077), .B(n6034), .C(n6058), .D(n6142), .Y(n6213));
  XOR2X1  g5080(.A(n6185), .B(n6213), .Y(n6214));
  INVX1   g5081(.A(n6185), .Y(n6215));
  INVX1   g5082(.A(P2_REG2_REG_7__SCAN_IN), .Y(n6216));
  NAND3X1 g5083(.A(n5890), .B(n5881), .C(P2_REG0_REG_7__SCAN_IN), .Y(n6217));
  OAI21X1 g5084(.A0(n5887), .A1(n6216), .B0(n6217), .Y(n6218));
  INVX1   g5085(.A(P2_REG1_REG_7__SCAN_IN), .Y(n6219));
  NAND4X1 g5086(.A(P2_REG3_REG_4__SCAN_IN), .B(P2_REG3_REG_5__SCAN_IN), .C(P2_REG3_REG_3__SCAN_IN), .D(P2_REG3_REG_6__SCAN_IN), .Y(n6220));
  XOR2X1  g5087(.A(n6220), .B(P2_REG3_REG_7__SCAN_IN), .Y(n6221));
  OAI22X1 g5088(.A0(n5894), .A1(n6221), .B0(n5891), .B1(n6219), .Y(n6222));
  NOR2X1  g5089(.A(n6222), .B(n6218), .Y(n6223));
  OAI22X1 g5090(.A0(n6215), .A1(n5928), .B0(n5965), .B1(n6223), .Y(n6224));
  AOI21X1 g5091(.A0(n6214), .A1(n5924), .B0(n6224), .Y(n6225));
  OAI21X1 g5092(.A0(n6206), .A1(n5914), .B0(n6225), .Y(n6226));
  NOR2X1  g5093(.A(n6226), .B(n6212), .Y(n6227));
  NAND2X1 g5094(.A(n5862), .B(P2_REG0_REG_6__SCAN_IN), .Y(n6228));
  OAI21X1 g5095(.A0(n6227), .A1(n5862), .B0(n6228), .Y(P2_U3469));
  AOI22X1 g5096(.A0(n5916), .A1(P2_REG2_REG_6__SCAN_IN), .B0(P2_REG0_REG_6__SCAN_IN), .B1(n5920), .Y(n6230));
  NAND3X1 g5097(.A(n6170), .B(n6166), .C(n6230), .Y(n6231));
  NAND2X1 g5098(.A(n6185), .B(n6231), .Y(n6232));
  INVX1   g5099(.A(n6232), .Y(n6233));
  INVX1   g5100(.A(n6223), .Y(n6234));
  NOR2X1  g5101(.A(P2_IR_REG_31__SCAN_IN), .B(n5515), .Y(n6235));
  AOI21X1 g5102(.A0(n5516), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6235), .Y(n6236));
  INVX1   g5103(.A(n6236), .Y(n6237));
  NAND3X1 g5104(.A(n6237), .B(n5871), .C(n5869), .Y(n6238));
  OAI21X1 g5105(.A0(n5867), .A1(n5514), .B0(n6238), .Y(n6239));
  OAI22X1 g5106(.A0(n6234), .A1(n6239), .B0(n6185), .B1(n6231), .Y(n6240));
  AOI21X1 g5107(.A0(n6239), .A1(n6234), .B0(n6240), .Y(n6241));
  OAI21X1 g5108(.A0(n6233), .A1(n6203), .B0(n6241), .Y(n6242));
  AOI21X1 g5109(.A0(n6215), .A1(n6172), .B0(n6202), .Y(n6243));
  XOR2X1  g5110(.A(n6239), .B(n6223), .Y(n6244));
  NAND2X1 g5111(.A(n6244), .B(n6232), .Y(n6245));
  OAI21X1 g5112(.A0(n6245), .A1(n6243), .B0(n6242), .Y(n6246));
  AOI21X1 g5113(.A0(n6097), .A1(n5904), .B0(n6246), .Y(n6247));
  NAND2X1 g5114(.A(n6133), .B(n6121), .Y(n6248));
  AOI21X1 g5115(.A0(n6248), .A1(n6136), .B0(n6190), .Y(n6249));
  AOI21X1 g5116(.A0(n6185), .A1(n6172), .B0(n6249), .Y(n6250));
  AOI21X1 g5117(.A0(n6033), .A1(n6015), .B0(n6043), .Y(n6251));
  NAND2X1 g5118(.A(n6251), .B(n6002), .Y(n6252));
  NAND2X1 g5119(.A(n6185), .B(n6172), .Y(n6253));
  NAND3X1 g5120(.A(n6253), .B(n6248), .C(n6135), .Y(n6254));
  AOI21X1 g5121(.A0(n6103), .A1(n6252), .B0(n6254), .Y(n6255));
  NOR2X1  g5122(.A(n6255), .B(n6250), .Y(n6256));
  XOR2X1  g5123(.A(n6256), .B(n6244), .Y(n6257));
  OAI22X1 g5124(.A0(n6246), .A1(n6071), .B0(n5902), .B1(n6257), .Y(n6258));
  INVX1   g5125(.A(n6257), .Y(n6259));
  AOI22X1 g5126(.A0(n6231), .A1(n5959), .B0(n5908), .B1(n6259), .Y(n6260));
  OAI21X1 g5127(.A0(n5907), .A1(n5900), .B0(n6259), .Y(n6261));
  NAND2X1 g5128(.A(n6261), .B(n6260), .Y(n6262));
  NOR4X1  g5129(.A(n6133), .B(n6112), .C(n6110), .D(n6185), .Y(n6263));
  INVX1   g5130(.A(n6239), .Y(n6264));
  XOR2X1  g5131(.A(n6264), .B(n6263), .Y(n6265));
  INVX1   g5132(.A(P2_REG2_REG_8__SCAN_IN), .Y(n6266));
  NAND3X1 g5133(.A(n5890), .B(n5881), .C(P2_REG0_REG_8__SCAN_IN), .Y(n6267));
  OAI21X1 g5134(.A0(n5887), .A1(n6266), .B0(n6267), .Y(n6268));
  INVX1   g5135(.A(P2_REG1_REG_8__SCAN_IN), .Y(n6269));
  INVX1   g5136(.A(P2_REG3_REG_8__SCAN_IN), .Y(n6270));
  INVX1   g5137(.A(P2_REG3_REG_7__SCAN_IN), .Y(n6271));
  NOR2X1  g5138(.A(n6220), .B(n6271), .Y(n6272));
  XOR2X1  g5139(.A(n6272), .B(n6270), .Y(n6273));
  OAI22X1 g5140(.A0(n5894), .A1(n6273), .B0(n5891), .B1(n6269), .Y(n6274));
  NOR2X1  g5141(.A(n6274), .B(n6268), .Y(n6275));
  OAI22X1 g5142(.A0(n6264), .A1(n5928), .B0(n5965), .B1(n6275), .Y(n6276));
  AOI21X1 g5143(.A0(n6265), .A1(n5924), .B0(n6276), .Y(n6277));
  OAI21X1 g5144(.A0(n6246), .A1(n5914), .B0(n6277), .Y(n6278));
  NOR4X1  g5145(.A(n6262), .B(n6258), .C(n6247), .D(n6278), .Y(n6279));
  NAND2X1 g5146(.A(n5862), .B(P2_REG0_REG_7__SCAN_IN), .Y(n6280));
  OAI21X1 g5147(.A0(n6279), .A1(n5862), .B0(n6280), .Y(P2_U3472));
  AOI21X1 g5148(.A0(n6264), .A1(n6232), .B0(n6223), .Y(n6282));
  AOI21X1 g5149(.A0(n6239), .A1(n6233), .B0(n6282), .Y(n6283));
  OAI21X1 g5150(.A0(n6240), .A1(n6202), .B0(n6283), .Y(n6284));
  NOR2X1  g5151(.A(P2_IR_REG_31__SCAN_IN), .B(n5522), .Y(n6285));
  AOI21X1 g5152(.A0(n5525), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6285), .Y(n6286));
  INVX1   g5153(.A(n6286), .Y(n6287));
  NAND3X1 g5154(.A(n6287), .B(n5871), .C(n5869), .Y(n6288));
  OAI21X1 g5155(.A0(n5867), .A1(n5521), .B0(n6288), .Y(n6289));
  XOR2X1  g5156(.A(n6289), .B(n6275), .Y(n6290));
  NOR2X1  g5157(.A(n6290), .B(n6284), .Y(n6291));
  INVX1   g5158(.A(n6275), .Y(n6292));
  XOR2X1  g5159(.A(n6289), .B(n6292), .Y(n6293));
  AOI21X1 g5160(.A0(n6290), .A1(n6284), .B0(n6291), .Y(n6295));
  AOI21X1 g5161(.A0(n6097), .A1(n5904), .B0(n6295), .Y(n6296));
  NOR2X1  g5162(.A(n6239), .B(n6223), .Y(n6297));
  NOR3X1  g5163(.A(n6255), .B(n6250), .C(n6297), .Y(n6298));
  AOI21X1 g5164(.A0(n6239), .A1(n6223), .B0(n6290), .Y(n6299));
  INVX1   g5165(.A(n6299), .Y(n6300));
  NOR3X1  g5166(.A(n6189), .B(n6112), .C(n6092), .Y(n6301));
  OAI21X1 g5167(.A0(n6301), .A1(n6190), .B0(n6253), .Y(n6302));
  NAND4X1 g5168(.A(n6248), .B(n6104), .C(n6135), .D(n6253), .Y(n6303));
  AOI22X1 g5169(.A0(n6302), .A1(n6303), .B0(n6239), .B1(n6223), .Y(n6304));
  INVX1   g5170(.A(n6297), .Y(n6305));
  NAND2X1 g5171(.A(n6290), .B(n6305), .Y(n6306));
  OAI22X1 g5172(.A0(n6304), .A1(n6306), .B0(n6300), .B1(n6298), .Y(n6307));
  NAND2X1 g5173(.A(n6307), .B(n5901), .Y(n6308));
  OAI21X1 g5174(.A0(n6295), .A1(n6071), .B0(n6308), .Y(n6309));
  AOI22X1 g5175(.A0(n6234), .A1(n5959), .B0(n5908), .B1(n6307), .Y(n6310));
  OAI21X1 g5176(.A0(n5907), .A1(n5900), .B0(n6307), .Y(n6311));
  NAND2X1 g5177(.A(n6311), .B(n6310), .Y(n6312));
  NOR2X1  g5178(.A(n5867), .B(n5521), .Y(n6313));
  AOI21X1 g5179(.A0(n6287), .A1(n5867), .B0(n6313), .Y(n6314));
  AOI21X1 g5180(.A0(n6264), .A1(n6263), .B0(n6314), .Y(n6315));
  NOR4X1  g5181(.A(n6239), .B(n6185), .C(n6213), .D(n6289), .Y(n6316));
  NOR2X1  g5182(.A(n6316), .B(n6315), .Y(n6317));
  INVX1   g5183(.A(P2_REG2_REG_9__SCAN_IN), .Y(n6318));
  NAND3X1 g5184(.A(n5890), .B(n5881), .C(P2_REG0_REG_9__SCAN_IN), .Y(n6319));
  OAI21X1 g5185(.A0(n5887), .A1(n6318), .B0(n6319), .Y(n6320));
  INVX1   g5186(.A(P2_REG1_REG_9__SCAN_IN), .Y(n6321));
  NOR3X1  g5187(.A(n5886), .B(n5881), .C(n6321), .Y(n6322));
  INVX1   g5188(.A(P2_REG3_REG_9__SCAN_IN), .Y(n6323));
  NOR3X1  g5189(.A(n6220), .B(n6270), .C(n6271), .Y(n6324));
  XOR2X1  g5190(.A(n6324), .B(n6323), .Y(n6325));
  NOR3X1  g5191(.A(n6325), .B(n5890), .C(n5881), .Y(n6326));
  NOR3X1  g5192(.A(n6326), .B(n6322), .C(n6320), .Y(n6327));
  OAI22X1 g5193(.A0(n6314), .A1(n5928), .B0(n5965), .B1(n6327), .Y(n6328));
  AOI21X1 g5194(.A0(n6317), .A1(n5924), .B0(n6328), .Y(n6329));
  OAI21X1 g5195(.A0(n6295), .A1(n5914), .B0(n6329), .Y(n6330));
  NOR4X1  g5196(.A(n6312), .B(n6309), .C(n6296), .D(n6330), .Y(n6331));
  NAND2X1 g5197(.A(n5862), .B(P2_REG0_REG_8__SCAN_IN), .Y(n6332));
  OAI21X1 g5198(.A0(n6331), .A1(n5862), .B0(n6332), .Y(P2_U3475));
  NOR2X1  g5199(.A(P2_IR_REG_31__SCAN_IN), .B(n5530), .Y(n6334));
  AOI21X1 g5200(.A0(n5531), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6334), .Y(n6335));
  INVX1   g5201(.A(n6335), .Y(n6336));
  NAND3X1 g5202(.A(n6336), .B(n5871), .C(n5869), .Y(n6337));
  OAI21X1 g5203(.A0(n5867), .A1(n5529), .B0(n6337), .Y(n6338));
  XOR2X1  g5204(.A(n6338), .B(n6327), .Y(n6339));
  AOI22X1 g5205(.A0(n6275), .A1(n6289), .B0(n6239), .B1(n6223), .Y(n6340));
  INVX1   g5206(.A(n6340), .Y(n6341));
  AOI21X1 g5207(.A0(n6303), .A1(n6302), .B0(n6341), .Y(n6342));
  OAI21X1 g5208(.A0(n6292), .A1(n6297), .B0(n6314), .Y(n6343));
  OAI21X1 g5209(.A0(n6275), .A1(n6305), .B0(n6343), .Y(n6344));
  NOR2X1  g5210(.A(n6344), .B(n6342), .Y(n6345));
  XOR2X1  g5211(.A(n6345), .B(n6339), .Y(n6346));
  INVX1   g5212(.A(n6346), .Y(n6347));
  OAI21X1 g5213(.A0(n5907), .A1(n5900), .B0(n6347), .Y(n6348));
  OAI21X1 g5214(.A0(n6346), .A1(n5902), .B0(n6348), .Y(n6349));
  NAND2X1 g5215(.A(n6314), .B(n6275), .Y(n6351));
  NOR2X1  g5216(.A(n6314), .B(n6275), .Y(n6352));
  AOI21X1 g5217(.A0(n6351), .A1(n6284), .B0(n6352), .Y(n6353));
  INVX1   g5218(.A(n6327), .Y(n6354));
  XOR2X1  g5219(.A(n6338), .B(n6354), .Y(n6355));
  NOR2X1  g5220(.A(n6355), .B(n6353), .Y(n6356));
  AOI21X1 g5221(.A0(n6353), .A1(n6355), .B0(n6356), .Y(n6357));
  AOI22X1 g5222(.A0(n6292), .A1(n5959), .B0(n5908), .B1(n6347), .Y(n6358));
  OAI21X1 g5223(.A0(n6357), .A1(n5904), .B0(n6358), .Y(n6359));
  INVX1   g5224(.A(n6357), .Y(n6360));
  OAI21X1 g5225(.A0(n5911), .A1(n5910), .B0(n6360), .Y(n6361));
  INVX1   g5226(.A(n6361), .Y(n6362));
  NOR2X1  g5227(.A(n5867), .B(n5529), .Y(n6363));
  AOI21X1 g5228(.A0(n6336), .A1(n5867), .B0(n6363), .Y(n6364));
  XOR2X1  g5229(.A(n6364), .B(n6316), .Y(n6365));
  INVX1   g5230(.A(P2_REG2_REG_10__SCAN_IN), .Y(n6366));
  NAND3X1 g5231(.A(n5890), .B(n5881), .C(P2_REG0_REG_10__SCAN_IN), .Y(n6367));
  OAI21X1 g5232(.A0(n5887), .A1(n6366), .B0(n6367), .Y(n6368));
  INVX1   g5233(.A(P2_REG1_REG_10__SCAN_IN), .Y(n6369));
  INVX1   g5234(.A(P2_REG3_REG_10__SCAN_IN), .Y(n6370));
  NOR4X1  g5235(.A(n6323), .B(n6270), .C(n6271), .D(n6220), .Y(n6371));
  XOR2X1  g5236(.A(n6371), .B(n6370), .Y(n6372));
  OAI22X1 g5237(.A0(n5894), .A1(n6372), .B0(n5891), .B1(n6369), .Y(n6373));
  NOR2X1  g5238(.A(n6373), .B(n6368), .Y(n6374));
  OAI22X1 g5239(.A0(n6364), .A1(n5928), .B0(n5965), .B1(n6374), .Y(n6375));
  AOI21X1 g5240(.A0(n6365), .A1(n5924), .B0(n6375), .Y(n6376));
  OAI21X1 g5241(.A0(n6357), .A1(n5914), .B0(n6376), .Y(n6377));
  NOR4X1  g5242(.A(n6362), .B(n6359), .C(n6349), .D(n6377), .Y(n6378));
  NAND2X1 g5243(.A(n5862), .B(P2_REG0_REG_9__SCAN_IN), .Y(n6379));
  OAI21X1 g5244(.A0(n6378), .A1(n5862), .B0(n6379), .Y(P2_U3478));
  INVX1   g5245(.A(n6353), .Y(n6381));
  NOR2X1  g5246(.A(n6364), .B(n6327), .Y(n6382));
  AOI22X1 g5247(.A0(n5916), .A1(P2_REG2_REG_10__SCAN_IN), .B0(P2_REG0_REG_10__SCAN_IN), .B1(n5920), .Y(n6383));
  INVX1   g5248(.A(n6372), .Y(n6384));
  AOI22X1 g5249(.A0(n5919), .A1(n6384), .B0(n5917), .B1(P2_REG1_REG_10__SCAN_IN), .Y(n6385));
  NAND2X1 g5250(.A(n6385), .B(n6383), .Y(n6386));
  NOR2X1  g5251(.A(P2_IR_REG_31__SCAN_IN), .B(n5536), .Y(n6387));
  AOI21X1 g5252(.A0(n5540), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6387), .Y(n6388));
  INVX1   g5253(.A(n6388), .Y(n6389));
  NAND3X1 g5254(.A(n6389), .B(n5871), .C(n5869), .Y(n6390));
  OAI21X1 g5255(.A0(n5867), .A1(n5535), .B0(n6390), .Y(n6391));
  OAI22X1 g5256(.A0(n6386), .A1(n6391), .B0(n6338), .B1(n6354), .Y(n6392));
  AOI21X1 g5257(.A0(n6391), .A1(n6386), .B0(n6392), .Y(n6393));
  OAI21X1 g5258(.A0(n6382), .A1(n6381), .B0(n6393), .Y(n6394));
  NOR2X1  g5259(.A(n6338), .B(n6354), .Y(n6395));
  XOR2X1  g5260(.A(n6391), .B(n6374), .Y(n6396));
  INVX1   g5261(.A(n6396), .Y(n6397));
  NOR2X1  g5262(.A(n6397), .B(n6382), .Y(n6398));
  OAI21X1 g5263(.A0(n6395), .A1(n6353), .B0(n6398), .Y(n6399));
  NAND2X1 g5264(.A(n6399), .B(n6394), .Y(n6400));
  AOI21X1 g5265(.A0(n6097), .A1(n5904), .B0(n6400), .Y(n6401));
  NAND2X1 g5266(.A(n6338), .B(n6327), .Y(n6402));
  INVX1   g5267(.A(n6402), .Y(n6403));
  OAI21X1 g5268(.A0(n6255), .A1(n6250), .B0(n6340), .Y(n6404));
  AOI21X1 g5269(.A0(n6275), .A1(n6305), .B0(n6289), .Y(n6405));
  AOI21X1 g5270(.A0(n6292), .A1(n6297), .B0(n6405), .Y(n6406));
  AOI21X1 g5271(.A0(n6406), .A1(n6404), .B0(n6403), .Y(n6407));
  AOI21X1 g5272(.A0(n6364), .A1(n6354), .B0(n6407), .Y(n6408));
  XOR2X1  g5273(.A(n6408), .B(n6396), .Y(n6409));
  OAI22X1 g5274(.A0(n6400), .A1(n6071), .B0(n5902), .B1(n6409), .Y(n6410));
  INVX1   g5275(.A(n6409), .Y(n6411));
  AOI22X1 g5276(.A0(n6354), .A1(n5959), .B0(n5908), .B1(n6411), .Y(n6412));
  OAI21X1 g5277(.A0(n5907), .A1(n5900), .B0(n6411), .Y(n6413));
  NAND2X1 g5278(.A(n6413), .B(n6412), .Y(n6414));
  NAND4X1 g5279(.A(n6314), .B(n6264), .C(n6263), .D(n6364), .Y(n6415));
  NOR2X1  g5280(.A(n6391), .B(n6338), .Y(n6416));
  AOI22X1 g5281(.A0(n6391), .A1(n6415), .B0(n6316), .B1(n6416), .Y(n6417));
  NOR2X1  g5282(.A(n5867), .B(n5535), .Y(n6418));
  AOI21X1 g5283(.A0(n6389), .A1(n5867), .B0(n6418), .Y(n6419));
  INVX1   g5284(.A(P2_REG2_REG_11__SCAN_IN), .Y(n6420));
  NAND3X1 g5285(.A(n5890), .B(n5881), .C(P2_REG0_REG_11__SCAN_IN), .Y(n6421));
  OAI21X1 g5286(.A0(n5887), .A1(n6420), .B0(n6421), .Y(n6422));
  INVX1   g5287(.A(P2_REG1_REG_11__SCAN_IN), .Y(n6423));
  NOR3X1  g5288(.A(n5886), .B(n5881), .C(n6423), .Y(n6424));
  INVX1   g5289(.A(P2_REG3_REG_11__SCAN_IN), .Y(n6425));
  INVX1   g5290(.A(n6371), .Y(n6426));
  NOR2X1  g5291(.A(n6426), .B(n6370), .Y(n6427));
  XOR2X1  g5292(.A(n6427), .B(n6425), .Y(n6428));
  NOR3X1  g5293(.A(n6428), .B(n5890), .C(n5881), .Y(n6429));
  NOR3X1  g5294(.A(n6429), .B(n6424), .C(n6422), .Y(n6430));
  OAI22X1 g5295(.A0(n6419), .A1(n5928), .B0(n5965), .B1(n6430), .Y(n6431));
  AOI21X1 g5296(.A0(n6417), .A1(n5924), .B0(n6431), .Y(n6432));
  OAI21X1 g5297(.A0(n6400), .A1(n5914), .B0(n6432), .Y(n6433));
  NOR4X1  g5298(.A(n6414), .B(n6410), .C(n6401), .D(n6433), .Y(n6434));
  NAND2X1 g5299(.A(n5862), .B(P2_REG0_REG_10__SCAN_IN), .Y(n6435));
  OAI21X1 g5300(.A0(n6434), .A1(n5862), .B0(n6435), .Y(P2_U3481));
  INVX1   g5301(.A(n6408), .Y(n6437));
  AOI21X1 g5302(.A0(n6419), .A1(n6386), .B0(n6437), .Y(n6438));
  NOR2X1  g5303(.A(P2_IR_REG_31__SCAN_IN), .B(n5545), .Y(n6439));
  AOI21X1 g5304(.A0(n5546), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6439), .Y(n6440));
  INVX1   g5305(.A(n6440), .Y(n6441));
  NAND3X1 g5306(.A(n6441), .B(n5871), .C(n5869), .Y(n6442));
  OAI21X1 g5307(.A0(n5867), .A1(n5544), .B0(n6442), .Y(n6443));
  XOR2X1  g5308(.A(n6443), .B(n6430), .Y(n6444));
  AOI21X1 g5309(.A0(n6391), .A1(n6374), .B0(n6444), .Y(n6445));
  INVX1   g5310(.A(n6445), .Y(n6446));
  NAND2X1 g5311(.A(n6391), .B(n6374), .Y(n6447));
  INVX1   g5312(.A(n6447), .Y(n6448));
  NAND2X1 g5313(.A(n6443), .B(n6430), .Y(n6449));
  INVX1   g5314(.A(n6449), .Y(n6450));
  INVX1   g5315(.A(n6430), .Y(n6451));
  NOR2X1  g5316(.A(n5867), .B(n5544), .Y(n6452));
  AOI21X1 g5317(.A0(n6441), .A1(n5867), .B0(n6452), .Y(n6453));
  AOI22X1 g5318(.A0(n6451), .A1(n6453), .B0(n6419), .B1(n6386), .Y(n6454));
  NOR2X1  g5319(.A(n8699), .B(n6450), .Y(n6456));
  OAI21X1 g5320(.A0(n6408), .A1(n6448), .B0(n6456), .Y(n6457));
  OAI21X1 g5321(.A0(n6446), .A1(n6438), .B0(n6457), .Y(n6458));
  INVX1   g5322(.A(n6458), .Y(n6459));
  NAND2X1 g5323(.A(n6391), .B(n6386), .Y(n6460));
  NOR2X1  g5324(.A(n6391), .B(n6386), .Y(n6461));
  AOI21X1 g5325(.A0(n6364), .A1(n6327), .B0(n6461), .Y(n6462));
  NAND3X1 g5326(.A(n6462), .B(n6351), .C(n6284), .Y(n6463));
  INVX1   g5327(.A(n6461), .Y(n6464));
  NOR3X1  g5328(.A(n6392), .B(n6314), .C(n6275), .Y(n6465));
  OAI21X1 g5329(.A0(n6465), .A1(n6382), .B0(n6464), .Y(n6466));
  NAND3X1 g5330(.A(n6466), .B(n6463), .C(n6460), .Y(n6467));
  NOR2X1  g5331(.A(n6467), .B(n6444), .Y(n6468));
  AOI21X1 g5332(.A0(n6444), .A1(n6467), .B0(n6468), .Y(n6470));
  NOR2X1  g5333(.A(n6470), .B(n6071), .Y(n6471));
  NOR2X1  g5334(.A(n6374), .B(n6072), .Y(n6472));
  NOR2X1  g5335(.A(n6470), .B(n6097), .Y(n6473));
  NOR2X1  g5336(.A(n6470), .B(n5904), .Y(n6479));
  NOR4X1  g5337(.A(n6473), .B(n6472), .C(n6471), .D(n6479), .Y(n6480));
  OAI21X1 g5338(.A0(n6459), .A1(n6128), .B0(n6480), .Y(n6481));
  OAI21X1 g5339(.A0(n5907), .A1(n5900), .B0(n6458), .Y(n6482));
  OAI21X1 g5340(.A0(n6459), .A1(n5902), .B0(n6482), .Y(n6483));
  NAND3X1 g5341(.A(n6419), .B(n6364), .C(n6316), .Y(n6484));
  XOR2X1  g5342(.A(n6443), .B(n6484), .Y(n6485));
  AOI22X1 g5343(.A0(n5916), .A1(P2_REG2_REG_12__SCAN_IN), .B0(P2_REG0_REG_12__SCAN_IN), .B1(n5920), .Y(n6486));
  NAND3X1 g5344(.A(n5890), .B(n5889), .C(P2_REG1_REG_12__SCAN_IN), .Y(n6487));
  INVX1   g5345(.A(P2_REG3_REG_12__SCAN_IN), .Y(n6488));
  NOR3X1  g5346(.A(n6426), .B(n6425), .C(n6370), .Y(n6489));
  XOR2X1  g5347(.A(n6489), .B(n6488), .Y(n6490));
  INVX1   g5348(.A(n6490), .Y(n6491));
  NAND3X1 g5349(.A(n6491), .B(n5886), .C(n5889), .Y(n6492));
  NAND3X1 g5350(.A(n6492), .B(n6487), .C(n6486), .Y(n6493));
  INVX1   g5351(.A(n6493), .Y(n6494));
  OAI22X1 g5352(.A0(n6453), .A1(n5928), .B0(n5965), .B1(n6494), .Y(n6495));
  AOI21X1 g5353(.A0(n6485), .A1(n5924), .B0(n6495), .Y(n6496));
  OAI21X1 g5354(.A0(n6470), .A1(n5914), .B0(n6496), .Y(n6497));
  NOR3X1  g5355(.A(n6497), .B(n6483), .C(n6481), .Y(n6498));
  NAND2X1 g5356(.A(n5862), .B(P2_REG0_REG_11__SCAN_IN), .Y(n6499));
  OAI21X1 g5357(.A0(n6498), .A1(n5862), .B0(n6499), .Y(P2_U3484));
  INVX1   g5358(.A(P2_IR_REG_12__SCAN_IN), .Y(n6501));
  NOR2X1  g5359(.A(P2_IR_REG_31__SCAN_IN), .B(n6501), .Y(n6502));
  AOI21X1 g5360(.A0(n5554), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6502), .Y(n6503));
  INVX1   g5361(.A(n6503), .Y(n6504));
  NAND3X1 g5362(.A(n6504), .B(n5871), .C(n5869), .Y(n6505));
  OAI21X1 g5363(.A0(n5867), .A1(n5551), .B0(n6505), .Y(n6506));
  XOR2X1  g5364(.A(n6506), .B(n6494), .Y(n6507));
  NAND3X1 g5365(.A(n6447), .B(n6364), .C(n6354), .Y(n6508));
  AOI21X1 g5366(.A0(n6508), .A1(n6454), .B0(n6450), .Y(n6509));
  NAND3X1 g5367(.A(n6449), .B(n6447), .C(n6402), .Y(n6510));
  AOI21X1 g5368(.A0(n6406), .A1(n6404), .B0(n6510), .Y(n6511));
  NOR2X1  g5369(.A(n6511), .B(n6509), .Y(n6512));
  XOR2X1  g5370(.A(n6512), .B(n6507), .Y(n6513));
  INVX1   g5371(.A(n6513), .Y(n6514));
  OAI21X1 g5372(.A0(n5907), .A1(n5900), .B0(n6514), .Y(n6515));
  OAI21X1 g5373(.A0(n6513), .A1(n5902), .B0(n6515), .Y(n6516));
  NOR2X1  g5374(.A(n6443), .B(n6451), .Y(n6517));
  INVX1   g5375(.A(n6517), .Y(n6518));
  NAND2X1 g5376(.A(n6443), .B(n6451), .Y(n6519));
  INVX1   g5377(.A(n6519), .Y(n6520));
  AOI21X1 g5378(.A0(n6467), .A1(n6518), .B0(n6520), .Y(n6521));
  INVX1   g5379(.A(n6521), .Y(n6522));
  NOR2X1  g5380(.A(n6522), .B(n6507), .Y(n6523));
  AOI21X1 g5381(.A0(n6507), .A1(n6522), .B0(n6523), .Y(n6525));
  AOI22X1 g5382(.A0(n6451), .A1(n5959), .B0(n5908), .B1(n6514), .Y(n6526));
  OAI21X1 g5383(.A0(n6525), .A1(n5904), .B0(n6526), .Y(n6527));
  INVX1   g5384(.A(n6506), .Y(n6528));
  NOR2X1  g5385(.A(n6528), .B(n6493), .Y(n6529));
  NOR2X1  g5386(.A(n6506), .B(n6494), .Y(n6530));
  OAI21X1 g5387(.A0(n6530), .A1(n6529), .B0(n6521), .Y(n6532));
  NAND2X1 g5388(.A(n6522), .B(n6507), .Y(n6534));
  AOI22X1 g5389(.A0(n6532), .A1(n6534), .B0(n6097), .B1(n6071), .Y(n6535));
  NAND3X1 g5390(.A(n6453), .B(n6416), .C(n6316), .Y(n6536));
  XOR2X1  g5391(.A(n6506), .B(n6536), .Y(n6537));
  AOI22X1 g5392(.A0(n5916), .A1(P2_REG2_REG_13__SCAN_IN), .B0(P2_REG0_REG_13__SCAN_IN), .B1(n5920), .Y(n6538));
  INVX1   g5393(.A(P2_REG1_REG_13__SCAN_IN), .Y(n6539));
  NOR3X1  g5394(.A(n5886), .B(n5881), .C(n6539), .Y(n6540));
  NAND4X1 g5395(.A(P2_REG3_REG_11__SCAN_IN), .B(P2_REG3_REG_12__SCAN_IN), .C(P2_REG3_REG_10__SCAN_IN), .D(n6371), .Y(n6541));
  XOR2X1  g5396(.A(n6541), .B(P2_REG3_REG_13__SCAN_IN), .Y(n6542));
  NOR3X1  g5397(.A(n6542), .B(n5890), .C(n5881), .Y(n6543));
  NOR2X1  g5398(.A(n6543), .B(n6540), .Y(n6544));
  NAND2X1 g5399(.A(n6544), .B(n6538), .Y(n6545));
  INVX1   g5400(.A(n6545), .Y(n6546));
  OAI22X1 g5401(.A0(n6528), .A1(n5928), .B0(n5965), .B1(n6546), .Y(n6547));
  AOI21X1 g5402(.A0(n6537), .A1(n5924), .B0(n6547), .Y(n6548));
  OAI21X1 g5403(.A0(n6525), .A1(n5914), .B0(n6548), .Y(n6549));
  NOR4X1  g5404(.A(n6535), .B(n6527), .C(n6516), .D(n6549), .Y(n6550));
  NAND2X1 g5405(.A(n5862), .B(P2_REG0_REG_12__SCAN_IN), .Y(n6551));
  OAI21X1 g5406(.A0(n6550), .A1(n5862), .B0(n6551), .Y(P2_U3487));
  NOR2X1  g5407(.A(n6528), .B(n6494), .Y(n6553));
  NOR2X1  g5408(.A(P2_IR_REG_31__SCAN_IN), .B(n5559), .Y(n6554));
  AOI21X1 g5409(.A0(n5562), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6554), .Y(n6555));
  INVX1   g5410(.A(n6555), .Y(n6556));
  NAND3X1 g5411(.A(n6556), .B(n5871), .C(n5869), .Y(n6557));
  OAI21X1 g5412(.A0(n5867), .A1(n5558), .B0(n6557), .Y(n6558));
  INVX1   g5413(.A(n6558), .Y(n6559));
  AOI22X1 g5414(.A0(n6546), .A1(n6559), .B0(n6528), .B1(n6494), .Y(n6560));
  INVX1   g5415(.A(n6560), .Y(n6561));
  AOI21X1 g5416(.A0(n6558), .A1(n6545), .B0(n6561), .Y(n6562));
  OAI21X1 g5417(.A0(n6522), .A1(n6553), .B0(n6562), .Y(n6563));
  NOR2X1  g5418(.A(n6559), .B(n6545), .Y(n6564));
  NOR2X1  g5419(.A(n6558), .B(n6546), .Y(n6565));
  NOR3X1  g5420(.A(n6565), .B(n6564), .C(n6553), .Y(n6566));
  INVX1   g5421(.A(n6566), .Y(n6567));
  AOI21X1 g5422(.A0(n6528), .A1(n6494), .B0(n6521), .Y(n6568));
  OAI21X1 g5423(.A0(n6568), .A1(n6567), .B0(n6563), .Y(n6569));
  OAI22X1 g5424(.A0(n6569), .A1(n6097), .B0(n5904), .B1(n6569), .Y(n6573));
  XOR2X1  g5425(.A(n6558), .B(n6546), .Y(n6574));
  INVX1   g5426(.A(n6509), .Y(n6575));
  INVX1   g5427(.A(n6510), .Y(n6576));
  OAI21X1 g5428(.A0(n6344), .A1(n6342), .B0(n6576), .Y(n6577));
  AOI21X1 g5429(.A0(n6577), .A1(n6575), .B0(n6529), .Y(n6578));
  NOR2X1  g5430(.A(n6578), .B(n6530), .Y(n6579));
  XOR2X1  g5431(.A(n6579), .B(n6574), .Y(n6580));
  OAI22X1 g5432(.A0(n6569), .A1(n6071), .B0(n5902), .B1(n6580), .Y(n6581));
  INVX1   g5433(.A(n6580), .Y(n6582));
  AOI22X1 g5434(.A0(n6493), .A1(n5959), .B0(n5908), .B1(n6582), .Y(n6583));
  OAI21X1 g5435(.A0(n5907), .A1(n5900), .B0(n6582), .Y(n6584));
  NAND2X1 g5436(.A(n6584), .B(n6583), .Y(n6585));
  NOR2X1  g5437(.A(n6506), .B(n6536), .Y(n6586));
  XOR2X1  g5438(.A(n6559), .B(n6586), .Y(n6587));
  AOI22X1 g5439(.A0(n5916), .A1(P2_REG2_REG_14__SCAN_IN), .B0(P2_REG0_REG_14__SCAN_IN), .B1(n5920), .Y(n6588));
  INVX1   g5440(.A(n6588), .Y(n6589));
  INVX1   g5441(.A(P2_REG1_REG_14__SCAN_IN), .Y(n6590));
  NOR3X1  g5442(.A(n5886), .B(n5881), .C(n6590), .Y(n6591));
  INVX1   g5443(.A(P2_REG3_REG_14__SCAN_IN), .Y(n6592));
  INVX1   g5444(.A(P2_REG3_REG_13__SCAN_IN), .Y(n6593));
  NOR2X1  g5445(.A(n6541), .B(n6593), .Y(n6594));
  XOR2X1  g5446(.A(n6594), .B(n6592), .Y(n6595));
  NOR3X1  g5447(.A(n6595), .B(n5890), .C(n5881), .Y(n6596));
  NOR3X1  g5448(.A(n6596), .B(n6591), .C(n6589), .Y(n6597));
  OAI22X1 g5449(.A0(n6559), .A1(n5928), .B0(n5965), .B1(n6597), .Y(n6598));
  AOI21X1 g5450(.A0(n6587), .A1(n5924), .B0(n6598), .Y(n6599));
  OAI21X1 g5451(.A0(n6569), .A1(n5914), .B0(n6599), .Y(n6600));
  NOR4X1  g5452(.A(n6585), .B(n6581), .C(n6573), .D(n6600), .Y(n6601));
  NAND2X1 g5453(.A(n5862), .B(P2_REG0_REG_13__SCAN_IN), .Y(n6602));
  OAI21X1 g5454(.A0(n6601), .A1(n5862), .B0(n6602), .Y(P2_U3490));
  INVX1   g5455(.A(P2_IR_REG_14__SCAN_IN), .Y(n6604));
  NOR2X1  g5456(.A(P2_IR_REG_31__SCAN_IN), .B(n6604), .Y(n6605));
  AOI21X1 g5457(.A0(n5570), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6605), .Y(n6606));
  INVX1   g5458(.A(n6606), .Y(n6607));
  NAND3X1 g5459(.A(n6607), .B(n5871), .C(n5869), .Y(n6608));
  OAI21X1 g5460(.A0(n5867), .A1(n5567), .B0(n6608), .Y(n6609));
  XOR2X1  g5461(.A(n6609), .B(n6597), .Y(n6610));
  INVX1   g5462(.A(n6530), .Y(n6611));
  OAI22X1 g5463(.A0(n6509), .A1(n6511), .B0(n6528), .B1(n6493), .Y(n6612));
  AOI21X1 g5464(.A0(n6612), .A1(n6611), .B0(n6564), .Y(n6613));
  NOR2X1  g5465(.A(n6613), .B(n6565), .Y(n6614));
  XOR2X1  g5466(.A(n6614), .B(n6610), .Y(n6615));
  INVX1   g5467(.A(n6610), .Y(n6616));
  OAI22X1 g5468(.A0(n6546), .A1(n6559), .B0(n6528), .B1(n6494), .Y(n6617));
  AOI21X1 g5469(.A0(n6560), .A1(n6520), .B0(n6617), .Y(n6618));
  AOI21X1 g5470(.A0(n6559), .A1(n6546), .B0(n6618), .Y(n6619));
  NOR2X1  g5471(.A(n6561), .B(n6517), .Y(n6620));
  AOI21X1 g5472(.A0(n6620), .A1(n6467), .B0(n6619), .Y(n6621));
  XOR2X1  g5473(.A(n6621), .B(n6616), .Y(n6622));
  OAI22X1 g5474(.A0(n6546), .A1(n6072), .B0(n6071), .B1(n6622), .Y(n6623));
  OAI22X1 g5475(.A0(n6622), .A1(n6097), .B0(n5904), .B1(n6622), .Y(n6626));
  NOR2X1  g5476(.A(n6626), .B(n6623), .Y(n6627));
  OAI21X1 g5477(.A0(n6615), .A1(n6128), .B0(n6627), .Y(n6628));
  NOR2X1  g5478(.A(n6615), .B(n5902), .Y(n6629));
  INVX1   g5479(.A(n5900), .Y(n6630));
  INVX1   g5480(.A(n5907), .Y(n6631));
  AOI21X1 g5481(.A0(n6631), .A1(n6630), .B0(n6615), .Y(n6632));
  NOR3X1  g5482(.A(n6558), .B(n6506), .C(n6536), .Y(n6633));
  INVX1   g5483(.A(n6609), .Y(n6634));
  NOR4X1  g5484(.A(n6558), .B(n6506), .C(n6536), .D(n6609), .Y(n6635));
  INVX1   g5485(.A(n6635), .Y(n6636));
  OAI21X1 g5486(.A0(n6634), .A1(n6633), .B0(n6636), .Y(n6637));
  NOR2X1  g5487(.A(n6637), .B(n5925), .Y(n6638));
  AOI22X1 g5488(.A0(n5916), .A1(P2_REG2_REG_15__SCAN_IN), .B0(P2_REG0_REG_15__SCAN_IN), .B1(n5920), .Y(n6639));
  NAND3X1 g5489(.A(n5890), .B(n5889), .C(P2_REG1_REG_15__SCAN_IN), .Y(n6640));
  NAND2X1 g5490(.A(n6594), .B(P2_REG3_REG_14__SCAN_IN), .Y(n6641));
  XOR2X1  g5491(.A(n6641), .B(P2_REG3_REG_15__SCAN_IN), .Y(n6642));
  INVX1   g5492(.A(n6642), .Y(n6643));
  NAND3X1 g5493(.A(n6643), .B(n5886), .C(n5889), .Y(n6644));
  NAND3X1 g5494(.A(n6644), .B(n6640), .C(n6639), .Y(n6645));
  INVX1   g5495(.A(n6645), .Y(n6646));
  OAI22X1 g5496(.A0(n6634), .A1(n5928), .B0(n5965), .B1(n6646), .Y(n6647));
  NOR2X1  g5497(.A(n6647), .B(n6638), .Y(n6648));
  OAI21X1 g5498(.A0(n6622), .A1(n5914), .B0(n6648), .Y(n6649));
  NOR4X1  g5499(.A(n6632), .B(n6629), .C(n6628), .D(n6649), .Y(n6650));
  NAND2X1 g5500(.A(n5862), .B(P2_REG0_REG_14__SCAN_IN), .Y(n6651));
  OAI21X1 g5501(.A0(n6650), .A1(n5862), .B0(n6651), .Y(P2_U3493));
  NOR2X1  g5502(.A(P2_IR_REG_31__SCAN_IN), .B(n5576), .Y(n6653));
  AOI21X1 g5503(.A0(n5577), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6653), .Y(n6654));
  INVX1   g5504(.A(n6654), .Y(n6655));
  NAND3X1 g5505(.A(n6655), .B(n5871), .C(n5869), .Y(n6656));
  OAI21X1 g5506(.A0(n5867), .A1(n5575), .B0(n6656), .Y(n6657));
  XOR2X1  g5507(.A(n6657), .B(n6646), .Y(n6658));
  INVX1   g5508(.A(n6658), .Y(n6659));
  INVX1   g5509(.A(n6597), .Y(n6660));
  NOR2X1  g5510(.A(n6634), .B(n6660), .Y(n6661));
  NAND2X1 g5511(.A(n6634), .B(n6660), .Y(n6662));
  OAI21X1 g5512(.A0(n6614), .A1(n6661), .B0(n6662), .Y(n6663));
  XOR2X1  g5513(.A(n6663), .B(n6659), .Y(n6664));
  NOR2X1  g5514(.A(n6634), .B(n6597), .Y(n6665));
  INVX1   g5515(.A(n6665), .Y(n6666));
  NOR2X1  g5516(.A(n6609), .B(n6660), .Y(n6667));
  OAI21X1 g5517(.A0(n6667), .A1(n6621), .B0(n6666), .Y(n6668));
  XOR2X1  g5518(.A(n6668), .B(n6658), .Y(n6669));
  OAI22X1 g5519(.A0(n6597), .A1(n6072), .B0(n6071), .B1(n6669), .Y(n6670));
  OAI22X1 g5520(.A0(n6669), .A1(n6097), .B0(n5904), .B1(n6669), .Y(n6673));
  NOR2X1  g5521(.A(n6673), .B(n6670), .Y(n6674));
  OAI21X1 g5522(.A0(n6664), .A1(n6128), .B0(n6674), .Y(n6675));
  NOR2X1  g5523(.A(n6664), .B(n5902), .Y(n6676));
  AOI21X1 g5524(.A0(n6631), .A1(n6630), .B0(n6664), .Y(n6677));
  INVX1   g5525(.A(n6657), .Y(n6678));
  XOR2X1  g5526(.A(n6678), .B(n6635), .Y(n6679));
  NAND3X1 g5527(.A(n5886), .B(n5881), .C(P2_REG2_REG_16__SCAN_IN), .Y(n6680));
  NAND3X1 g5528(.A(n5890), .B(n5881), .C(P2_REG0_REG_16__SCAN_IN), .Y(n6681));
  NAND3X1 g5529(.A(n5890), .B(n5889), .C(P2_REG1_REG_16__SCAN_IN), .Y(n6682));
  INVX1   g5530(.A(P2_REG3_REG_16__SCAN_IN), .Y(n6683));
  INVX1   g5531(.A(P2_REG3_REG_15__SCAN_IN), .Y(n6684));
  NOR4X1  g5532(.A(n6684), .B(n6593), .C(n6592), .D(n6541), .Y(n6685));
  XOR2X1  g5533(.A(n6685), .B(n6683), .Y(n6686));
  INVX1   g5534(.A(n6686), .Y(n6687));
  NAND3X1 g5535(.A(n6687), .B(n5886), .C(n5889), .Y(n6688));
  NAND4X1 g5536(.A(n6682), .B(n6681), .C(n6680), .D(n6688), .Y(n6689));
  INVX1   g5537(.A(n6689), .Y(n6690));
  OAI22X1 g5538(.A0(n6678), .A1(n5928), .B0(n5965), .B1(n6690), .Y(n6691));
  AOI21X1 g5539(.A0(n6679), .A1(n5924), .B0(n6691), .Y(n6692));
  OAI21X1 g5540(.A0(n6669), .A1(n5914), .B0(n6692), .Y(n6693));
  NOR4X1  g5541(.A(n6677), .B(n6676), .C(n6675), .D(n6693), .Y(n6694));
  NAND2X1 g5542(.A(n5862), .B(P2_REG0_REG_15__SCAN_IN), .Y(n6695));
  OAI21X1 g5543(.A0(n6694), .A1(n5862), .B0(n6695), .Y(P2_U3496));
  NOR2X1  g5544(.A(n6678), .B(n6645), .Y(n6697));
  AOI21X1 g5545(.A0(n6678), .A1(n6645), .B0(n6663), .Y(n6698));
  NAND2X1 g5546(.A(n5470), .B(P2_IR_REG_16__SCAN_IN), .Y(n6699));
  INVX1   g5547(.A(n6699), .Y(n6700));
  AOI21X1 g5548(.A0(n5587), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6700), .Y(n6701));
  INVX1   g5549(.A(n6701), .Y(n6702));
  NAND2X1 g5550(.A(n6702), .B(n5867), .Y(n6703));
  OAI21X1 g5551(.A0(n5867), .A1(n5582), .B0(n6703), .Y(n6704));
  XOR2X1  g5552(.A(n6704), .B(n6690), .Y(n6705));
  NOR3X1  g5553(.A(n6705), .B(n6698), .C(n6697), .Y(n6706));
  OAI21X1 g5554(.A0(n6678), .A1(n6645), .B0(n6663), .Y(n6707));
  OAI22X1 g5555(.A0(n6690), .A1(n6704), .B0(n6657), .B1(n6646), .Y(n6708));
  AOI21X1 g5556(.A0(n6704), .A1(n6690), .B0(n6708), .Y(n6709));
  AOI21X1 g5557(.A0(n6709), .A1(n6707), .B0(n6706), .Y(n6710));
  NOR2X1  g5558(.A(n6678), .B(n6646), .Y(n6712));
  NOR2X1  g5559(.A(n6657), .B(n6645), .Y(n6713));
  INVX1   g5560(.A(n6713), .Y(n6714));
  AOI21X1 g5561(.A0(n6714), .A1(n6668), .B0(n6712), .Y(n6715));
  XOR2X1  g5562(.A(n6704), .B(n6689), .Y(n6716));
  NOR2X1  g5563(.A(n6716), .B(n6715), .Y(n6717));
  AOI21X1 g5564(.A0(n6715), .A1(n6716), .B0(n6717), .Y(n6718));
  OAI22X1 g5565(.A0(n6646), .A1(n6072), .B0(n6071), .B1(n6718), .Y(n6719));
  OAI22X1 g5566(.A0(n6718), .A1(n6097), .B0(n5904), .B1(n6718), .Y(n6723));
  NOR2X1  g5567(.A(n6723), .B(n6719), .Y(n6724));
  OAI21X1 g5568(.A0(n6710), .A1(n6128), .B0(n6724), .Y(n6725));
  NOR2X1  g5569(.A(n6710), .B(n5902), .Y(n6726));
  AOI21X1 g5570(.A0(n6631), .A1(n6630), .B0(n6710), .Y(n6727));
  NAND2X1 g5571(.A(n6678), .B(n6635), .Y(n6728));
  XOR2X1  g5572(.A(n6704), .B(n6728), .Y(n6729));
  NOR2X1  g5573(.A(n5867), .B(n5582), .Y(n6730));
  AOI21X1 g5574(.A0(n6702), .A1(n5867), .B0(n6730), .Y(n6731));
  INVX1   g5575(.A(P2_REG3_REG_17__SCAN_IN), .Y(n6732));
  NOR3X1  g5576(.A(n6641), .B(n6684), .C(n6683), .Y(n6733));
  XOR2X1  g5577(.A(n6733), .B(n6732), .Y(n6734));
  NOR3X1  g5578(.A(n6734), .B(n5890), .C(n5881), .Y(n6735));
  INVX1   g5579(.A(P2_REG0_REG_17__SCAN_IN), .Y(n6736));
  NOR3X1  g5580(.A(n5886), .B(n5889), .C(n6736), .Y(n6737));
  AOI22X1 g5581(.A0(n5916), .A1(P2_REG2_REG_17__SCAN_IN), .B0(P2_REG1_REG_17__SCAN_IN), .B1(n5917), .Y(n6738));
  INVX1   g5582(.A(n6738), .Y(n6739));
  NOR3X1  g5583(.A(n6739), .B(n6737), .C(n6735), .Y(n6740));
  OAI22X1 g5584(.A0(n6731), .A1(n5928), .B0(n5965), .B1(n6740), .Y(n6741));
  AOI21X1 g5585(.A0(n6729), .A1(n5924), .B0(n6741), .Y(n6742));
  OAI21X1 g5586(.A0(n6718), .A1(n5914), .B0(n6742), .Y(n6743));
  NOR4X1  g5587(.A(n6727), .B(n6726), .C(n6725), .D(n6743), .Y(n6744));
  NAND2X1 g5588(.A(n5862), .B(P2_REG0_REG_16__SCAN_IN), .Y(n6745));
  OAI21X1 g5589(.A0(n6744), .A1(n5862), .B0(n6745), .Y(P2_U3499));
  INVX1   g5590(.A(n6740), .Y(n6747));
  NAND2X1 g5591(.A(n5470), .B(P2_IR_REG_17__SCAN_IN), .Y(n6748));
  INVX1   g5592(.A(n6748), .Y(n6749));
  AOI21X1 g5593(.A0(n5593), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6749), .Y(n6750));
  INVX1   g5594(.A(n6750), .Y(n6751));
  NAND3X1 g5595(.A(n6751), .B(n5871), .C(n5869), .Y(n6752));
  OAI21X1 g5596(.A0(n5867), .A1(n5592), .B0(n6752), .Y(n6753));
  INVX1   g5597(.A(n6753), .Y(n6754));
  AOI22X1 g5598(.A0(n6740), .A1(n6754), .B0(n6731), .B1(n6690), .Y(n6755));
  INVX1   g5599(.A(n6755), .Y(n6756));
  AOI21X1 g5600(.A0(n6753), .A1(n6747), .B0(n6756), .Y(n6757));
  OAI21X1 g5601(.A0(n6731), .A1(n6690), .B0(n6715), .Y(n6758));
  NAND2X1 g5602(.A(n6758), .B(n6757), .Y(n6759));
  NOR2X1  g5603(.A(n6731), .B(n6690), .Y(n6760));
  NOR2X1  g5604(.A(n6754), .B(n6747), .Y(n6761));
  NOR2X1  g5605(.A(n6753), .B(n6740), .Y(n6762));
  NOR3X1  g5606(.A(n6762), .B(n6761), .C(n6760), .Y(n6763));
  INVX1   g5607(.A(n6763), .Y(n6764));
  AOI21X1 g5608(.A0(n6731), .A1(n6690), .B0(n6715), .Y(n6765));
  OAI21X1 g5609(.A0(n6765), .A1(n6764), .B0(n6759), .Y(n6766));
  OAI22X1 g5610(.A0(n6766), .A1(n6097), .B0(n5904), .B1(n6766), .Y(n6771));
  XOR2X1  g5611(.A(n6753), .B(n6740), .Y(n6772));
  NOR2X1  g5612(.A(n6697), .B(n6662), .Y(n6773));
  OAI22X1 g5613(.A0(n6708), .A1(n6773), .B0(n6731), .B1(n6689), .Y(n6774));
  INVX1   g5614(.A(n6565), .Y(n6776));
  OAI22X1 g5615(.A0(n6645), .A1(n6678), .B0(n6634), .B1(n6660), .Y(n6778));
  AOI21X1 g5616(.A0(n6704), .A1(n6690), .B0(n6778), .Y(n6779));
  INVX1   g5617(.A(n6779), .Y(n6780));
  AOI21X1 g5618(.A0(n8715), .A1(n6776), .B0(n6780), .Y(n6781));
  NOR2X1  g5619(.A(n6781), .B(n8865), .Y(n6782));
  XOR2X1  g5620(.A(n6782), .B(n6772), .Y(n6783));
  OAI22X1 g5621(.A0(n6766), .A1(n6071), .B0(n5902), .B1(n6783), .Y(n6784));
  INVX1   g5622(.A(n6783), .Y(n6785));
  AOI22X1 g5623(.A0(n6689), .A1(n5959), .B0(n5908), .B1(n6785), .Y(n6786));
  OAI21X1 g5624(.A0(n5907), .A1(n5900), .B0(n6785), .Y(n6787));
  NAND2X1 g5625(.A(n6787), .B(n6786), .Y(n6788));
  NAND3X1 g5626(.A(n6731), .B(n6678), .C(n6635), .Y(n6789));
  XOR2X1  g5627(.A(n6753), .B(n6789), .Y(n6790));
  NOR4X1  g5628(.A(n6684), .B(n6732), .C(n6683), .D(n6641), .Y(n6791));
  XOR2X1  g5629(.A(n6791), .B(P2_REG3_REG_18__SCAN_IN), .Y(n6792));
  INVX1   g5630(.A(n6792), .Y(n6793));
  NOR3X1  g5631(.A(n6793), .B(n5890), .C(n5881), .Y(n6794));
  INVX1   g5632(.A(P2_REG0_REG_18__SCAN_IN), .Y(n6795));
  NOR3X1  g5633(.A(n5886), .B(n5889), .C(n6795), .Y(n6796));
  AOI22X1 g5634(.A0(n5916), .A1(P2_REG2_REG_18__SCAN_IN), .B0(P2_REG1_REG_18__SCAN_IN), .B1(n5917), .Y(n6797));
  INVX1   g5635(.A(n6797), .Y(n6798));
  NOR3X1  g5636(.A(n6798), .B(n6796), .C(n6794), .Y(n6799));
  OAI22X1 g5637(.A0(n6754), .A1(n5928), .B0(n5965), .B1(n6799), .Y(n6800));
  AOI21X1 g5638(.A0(n6790), .A1(n5924), .B0(n6800), .Y(n6801));
  OAI21X1 g5639(.A0(n6766), .A1(n5914), .B0(n6801), .Y(n6802));
  NOR4X1  g5640(.A(n6788), .B(n6784), .C(n6771), .D(n6802), .Y(n6803));
  NAND2X1 g5641(.A(n5862), .B(P2_REG0_REG_17__SCAN_IN), .Y(n6804));
  OAI21X1 g5642(.A0(n6803), .A1(n5862), .B0(n6804), .Y(P2_U3502));
  NAND3X1 g5643(.A(n6753), .B(n6704), .C(n6689), .Y(n6806));
  AOI21X1 g5644(.A0(n6704), .A1(n6689), .B0(n6753), .Y(n6807));
  OAI21X1 g5645(.A0(n6807), .A1(n6740), .B0(n6806), .Y(n6808));
  INVX1   g5646(.A(n6808), .Y(n6809));
  OAI21X1 g5647(.A0(n6756), .A1(n6715), .B0(n6809), .Y(n6810));
  NOR2X1  g5648(.A(P2_IR_REG_31__SCAN_IN), .B(n5599), .Y(n6811));
  AOI21X1 g5649(.A0(n5611), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6811), .Y(n6812));
  INVX1   g5650(.A(n6812), .Y(n6813));
  NAND3X1 g5651(.A(n6813), .B(n5871), .C(n5869), .Y(n6814));
  OAI21X1 g5652(.A0(n5867), .A1(n5598), .B0(n6814), .Y(n6815));
  XOR2X1  g5653(.A(n6815), .B(n6799), .Y(n6816));
  NOR2X1  g5654(.A(n6810), .B(n6816), .Y(n6817));
  INVX1   g5655(.A(n6799), .Y(n6818));
  AOI21X1 g5656(.A0(n6816), .A1(n6810), .B0(n6817), .Y(n6821));
  OAI22X1 g5657(.A0(n6740), .A1(n6072), .B0(n6071), .B1(n6821), .Y(n6822));
  OAI22X1 g5658(.A0(n6821), .A1(n6097), .B0(n5904), .B1(n6821), .Y(n6826));
  INVX1   g5659(.A(n6762), .Y(n6827));
  OAI22X1 g5660(.A0(n8865), .A1(n6781), .B0(n6754), .B1(n6747), .Y(n6828));
  NAND2X1 g5661(.A(n6828), .B(n6827), .Y(n6829));
  XOR2X1  g5662(.A(n6829), .B(n6816), .Y(n6830));
  OAI21X1 g5663(.A0(n5908), .A1(n5907), .B0(n6830), .Y(n6831));
  OAI21X1 g5664(.A0(n5901), .A1(n5900), .B0(n6830), .Y(n6832));
  NAND2X1 g5665(.A(n6832), .B(n6831), .Y(n6833));
  NAND4X1 g5666(.A(n6731), .B(n6678), .C(n6635), .D(n6754), .Y(n6834));
  XOR2X1  g5667(.A(n6815), .B(n6834), .Y(n6835));
  NOR2X1  g5668(.A(n5867), .B(n5598), .Y(n6836));
  AOI21X1 g5669(.A0(n6813), .A1(n5867), .B0(n6836), .Y(n6837));
  NAND4X1 g5670(.A(P2_REG3_REG_18__SCAN_IN), .B(P2_REG3_REG_17__SCAN_IN), .C(P2_REG3_REG_16__SCAN_IN), .D(n6685), .Y(n6838));
  XOR2X1  g5671(.A(n6838), .B(P2_REG3_REG_19__SCAN_IN), .Y(n6839));
  NOR3X1  g5672(.A(n6839), .B(n5890), .C(n5881), .Y(n6840));
  INVX1   g5673(.A(P2_REG1_REG_19__SCAN_IN), .Y(n6841));
  NOR3X1  g5674(.A(n5886), .B(n5881), .C(n6841), .Y(n6842));
  NAND3X1 g5675(.A(n5886), .B(n5881), .C(P2_REG2_REG_19__SCAN_IN), .Y(n6843));
  NAND3X1 g5676(.A(n5890), .B(n5881), .C(P2_REG0_REG_19__SCAN_IN), .Y(n6844));
  NAND2X1 g5677(.A(n6844), .B(n6843), .Y(n6845));
  NOR3X1  g5678(.A(n6845), .B(n6842), .C(n6840), .Y(n6846));
  OAI22X1 g5679(.A0(n6837), .A1(n5928), .B0(n5965), .B1(n6846), .Y(n6847));
  AOI21X1 g5680(.A0(n6835), .A1(n5924), .B0(n6847), .Y(n6848));
  OAI21X1 g5681(.A0(n6821), .A1(n5914), .B0(n6848), .Y(n6849));
  NOR4X1  g5682(.A(n6833), .B(n6826), .C(n6822), .D(n6849), .Y(n6850));
  NAND2X1 g5683(.A(n5862), .B(P2_REG0_REG_18__SCAN_IN), .Y(n6851));
  OAI21X1 g5684(.A0(n6850), .A1(n5862), .B0(n6851), .Y(P2_U3505));
  NAND3X1 g5685(.A(n5871), .B(n5869), .C(n5856), .Y(n6853));
  OAI21X1 g5686(.A0(n5867), .A1(n5616), .B0(n6853), .Y(n6854));
  XOR2X1  g5687(.A(n6854), .B(n6846), .Y(n6855));
  NOR2X1  g5688(.A(n6815), .B(n6799), .Y(n6856));
  AOI21X1 g5689(.A0(n6828), .A1(n6827), .B0(n6799), .Y(n6857));
  AOI21X1 g5690(.A0(n6828), .A1(n6827), .B0(n6815), .Y(n6858));
  NOR3X1  g5691(.A(n6858), .B(n6857), .C(n6856), .Y(n6859));
  XOR2X1  g5692(.A(n6859), .B(n6855), .Y(n6860));
  NOR2X1  g5693(.A(n6860), .B(n6128), .Y(n6861));
  INVX1   g5694(.A(n6861), .Y(n6862));
  NOR2X1  g5695(.A(n6815), .B(n6818), .Y(n6863));
  INVX1   g5696(.A(n6863), .Y(n6864));
  NAND2X1 g5697(.A(n6815), .B(n6818), .Y(n6865));
  INVX1   g5698(.A(n6865), .Y(n6866));
  AOI21X1 g5699(.A0(n6864), .A1(n6810), .B0(n6866), .Y(n6867));
  NAND2X1 g5700(.A(n6854), .B(n6846), .Y(n6868));
  INVX1   g5701(.A(n6868), .Y(n6869));
  NOR2X1  g5702(.A(n6854), .B(n6846), .Y(n6870));
  OAI21X1 g5703(.A0(n6870), .A1(n6869), .B0(n6867), .Y(n6871));
  INVX1   g5704(.A(n6846), .Y(n6872));
  XOR2X1  g5705(.A(n6854), .B(n6872), .Y(n6873));
  OAI21X1 g5706(.A0(n6873), .A1(n6867), .B0(n6871), .Y(n6874));
  AOI22X1 g5707(.A0(n6818), .A1(n5959), .B0(n5910), .B1(n6874), .Y(n6875));
  AOI22X1 g5708(.A0(n6874), .A1(n5911), .B0(n5903), .B1(n6874), .Y(n6879));
  NAND3X1 g5709(.A(n6879), .B(n6875), .C(n6862), .Y(n6880));
  NOR2X1  g5710(.A(n6860), .B(n5902), .Y(n6881));
  AOI21X1 g5711(.A0(n6631), .A1(n6630), .B0(n6860), .Y(n6882));
  NAND4X1 g5712(.A(n5856), .B(n5852), .C(n5850), .D(n6874), .Y(n6883));
  NOR3X1  g5713(.A(n6815), .B(n6753), .C(n6789), .Y(n6884));
  INVX1   g5714(.A(n6854), .Y(n6885));
  XOR2X1  g5715(.A(n6885), .B(n6884), .Y(n6886));
  NAND3X1 g5716(.A(n6791), .B(P2_REG3_REG_18__SCAN_IN), .C(P2_REG3_REG_19__SCAN_IN), .Y(n6887));
  XOR2X1  g5717(.A(n6887), .B(P2_REG3_REG_20__SCAN_IN), .Y(n6888));
  NOR3X1  g5718(.A(n6888), .B(n5890), .C(n5881), .Y(n6889));
  NAND3X1 g5719(.A(n5890), .B(n5889), .C(P2_REG1_REG_20__SCAN_IN), .Y(n6890));
  NAND3X1 g5720(.A(n5886), .B(n5881), .C(P2_REG2_REG_20__SCAN_IN), .Y(n6891));
  NAND3X1 g5721(.A(n5890), .B(n5881), .C(P2_REG0_REG_20__SCAN_IN), .Y(n6892));
  NAND3X1 g5722(.A(n6892), .B(n6891), .C(n6890), .Y(n6893));
  NOR2X1  g5723(.A(n6893), .B(n6889), .Y(n6894));
  OAI22X1 g5724(.A0(n6885), .A1(n5928), .B0(n5965), .B1(n6894), .Y(n6895));
  AOI21X1 g5725(.A0(n6886), .A1(n5924), .B0(n6895), .Y(n6896));
  NAND2X1 g5726(.A(n6896), .B(n6883), .Y(n6897));
  NOR4X1  g5727(.A(n6882), .B(n6881), .C(n6880), .D(n6897), .Y(n6898));
  NAND2X1 g5728(.A(n5862), .B(P2_REG0_REG_19__SCAN_IN), .Y(n6899));
  OAI21X1 g5729(.A0(n6898), .A1(n5862), .B0(n6899), .Y(P2_U3507));
  NOR2X1  g5730(.A(n5867), .B(n5624), .Y(n6901));
  XOR2X1  g5731(.A(n6901), .B(n6894), .Y(n6902));
  INVX1   g5732(.A(n6856), .Y(n6903));
  AOI21X1 g5733(.A0(n8857), .A1(n6774), .B0(n6761), .Y(n6905));
  OAI21X1 g5734(.A0(n6905), .A1(n6762), .B0(n6818), .Y(n6906));
  OAI21X1 g5735(.A0(n6905), .A1(n6762), .B0(n6837), .Y(n6907));
  NAND3X1 g5736(.A(n6907), .B(n6906), .C(n6903), .Y(n6908));
  AOI21X1 g5737(.A0(n6908), .A1(n6868), .B0(n6870), .Y(n6909));
  XOR2X1  g5738(.A(n6909), .B(n6902), .Y(n6910));
  NOR2X1  g5739(.A(n6910), .B(n6128), .Y(n6911));
  NOR2X1  g5740(.A(n6885), .B(n6846), .Y(n6912));
  INVX1   g5741(.A(n6912), .Y(n6913));
  INVX1   g5742(.A(n6894), .Y(n6914));
  OAI22X1 g5743(.A0(n6914), .A1(n6901), .B0(n6854), .B1(n6872), .Y(n6915));
  AOI21X1 g5744(.A0(n6901), .A1(n6914), .B0(n6915), .Y(n6916));
  INVX1   g5745(.A(n6916), .Y(n6917));
  AOI21X1 g5746(.A0(n6913), .A1(n6867), .B0(n6917), .Y(n6918));
  INVX1   g5747(.A(n6918), .Y(n6919));
  NOR2X1  g5748(.A(n6854), .B(n6872), .Y(n6920));
  NOR3X1  g5749(.A(n6914), .B(n5867), .C(n5624), .Y(n6921));
  NOR2X1  g5750(.A(n6901), .B(n6894), .Y(n6922));
  NOR3X1  g5751(.A(n6922), .B(n6921), .C(n6912), .Y(n6923));
  OAI21X1 g5752(.A0(n6920), .A1(n6867), .B0(n6923), .Y(n6924));
  NAND2X1 g5753(.A(n6924), .B(n6919), .Y(n6925));
  OAI22X1 g5754(.A0(n6846), .A1(n6072), .B0(n6071), .B1(n6925), .Y(n6926));
  OAI22X1 g5755(.A0(n6925), .A1(n6097), .B0(n5904), .B1(n6925), .Y(n6931));
  NOR3X1  g5756(.A(n6931), .B(n6926), .C(n6911), .Y(n6932));
  NOR2X1  g5757(.A(n6910), .B(n5902), .Y(n6933));
  AOI21X1 g5758(.A0(n6631), .A1(n6630), .B0(n6910), .Y(n6934));
  NOR2X1  g5759(.A(n6934), .B(n6933), .Y(n6935));
  NAND2X1 g5760(.A(n6935), .B(n6932), .Y(n6936));
  NAND2X1 g5761(.A(n6885), .B(n6884), .Y(n6937));
  XOR2X1  g5762(.A(n6901), .B(n6937), .Y(n6938));
  INVX1   g5763(.A(n6901), .Y(n6939));
  NAND4X1 g5764(.A(P2_REG3_REG_18__SCAN_IN), .B(P2_REG3_REG_20__SCAN_IN), .C(P2_REG3_REG_19__SCAN_IN), .D(n6791), .Y(n6940));
  XOR2X1  g5765(.A(n6940), .B(P2_REG3_REG_21__SCAN_IN), .Y(n6941));
  NOR3X1  g5766(.A(n6941), .B(n5890), .C(n5881), .Y(n6942));
  INVX1   g5767(.A(n6942), .Y(n6943));
  NAND3X1 g5768(.A(n5890), .B(n5889), .C(P2_REG1_REG_21__SCAN_IN), .Y(n6944));
  AOI22X1 g5769(.A0(n5916), .A1(P2_REG2_REG_21__SCAN_IN), .B0(P2_REG0_REG_21__SCAN_IN), .B1(n5920), .Y(n6945));
  NAND3X1 g5770(.A(n6945), .B(n6944), .C(n6943), .Y(n6946));
  INVX1   g5771(.A(n6946), .Y(n6947));
  OAI22X1 g5772(.A0(n6939), .A1(n5928), .B0(n5965), .B1(n6947), .Y(n6948));
  AOI21X1 g5773(.A0(n6938), .A1(n5924), .B0(n6948), .Y(n6949));
  OAI21X1 g5774(.A0(n6925), .A1(n5914), .B0(n6949), .Y(n6950));
  NOR2X1  g5775(.A(n6950), .B(n6936), .Y(n6951));
  NAND2X1 g5776(.A(n5862), .B(P2_REG0_REG_20__SCAN_IN), .Y(n6952));
  OAI21X1 g5777(.A0(n6951), .A1(n5862), .B0(n6952), .Y(P2_U3508));
  NOR2X1  g5778(.A(n5867), .B(n5633), .Y(n6954));
  XOR2X1  g5779(.A(n6954), .B(n6947), .Y(n6955));
  INVX1   g5780(.A(n6921), .Y(n6956));
  INVX1   g5781(.A(n6870), .Y(n6957));
  OAI21X1 g5782(.A0(n6859), .A1(n6869), .B0(n6957), .Y(n6958));
  AOI21X1 g5783(.A0(n6958), .A1(n6956), .B0(n6922), .Y(n6959));
  XOR2X1  g5784(.A(n6959), .B(n6955), .Y(n6960));
  INVX1   g5785(.A(n6960), .Y(n6961));
  NAND2X1 g5786(.A(n6961), .B(n5908), .Y(n6962));
  NOR2X1  g5787(.A(n6915), .B(n6867), .Y(n6963));
  AOI21X1 g5788(.A0(n6854), .A1(n6872), .B0(n6901), .Y(n6964));
  AOI21X1 g5789(.A0(n6901), .A1(n6912), .B0(n6914), .Y(n6965));
  NOR2X1  g5790(.A(n6965), .B(n6964), .Y(n6966));
  NOR2X1  g5791(.A(n6963), .B(n6966), .Y(n6967));
  NOR3X1  g5792(.A(n6946), .B(n5867), .C(n5633), .Y(n6968));
  NOR2X1  g5793(.A(n6954), .B(n6947), .Y(n6969));
  NOR3X1  g5794(.A(n6966), .B(n6969), .C(n6968), .Y(n6970));
  INVX1   g5795(.A(n6970), .Y(n6971));
  OAI22X1 g5796(.A0(n6967), .A1(n6955), .B0(n6963), .B1(n6971), .Y(n6972));
  OAI22X1 g5797(.A0(n6894), .A1(n6072), .B0(n6071), .B1(n6972), .Y(n6973));
  OAI22X1 g5798(.A0(n6972), .A1(n6097), .B0(n5904), .B1(n6972), .Y(n6977));
  NOR2X1  g5799(.A(n6977), .B(n6973), .Y(n6978));
  AOI21X1 g5800(.A0(n6631), .A1(n6630), .B0(n6960), .Y(n6979));
  AOI21X1 g5801(.A0(n6961), .A1(n5901), .B0(n6979), .Y(n6980));
  NAND3X1 g5802(.A(n6980), .B(n6978), .C(n6962), .Y(n6981));
  NAND3X1 g5803(.A(n6939), .B(n6885), .C(n6884), .Y(n6982));
  XOR2X1  g5804(.A(n6954), .B(n6982), .Y(n6983));
  INVX1   g5805(.A(n6954), .Y(n6984));
  INVX1   g5806(.A(P2_REG3_REG_22__SCAN_IN), .Y(n6985));
  INVX1   g5807(.A(P2_REG3_REG_21__SCAN_IN), .Y(n6986));
  NOR2X1  g5808(.A(n6940), .B(n6986), .Y(n6987));
  XOR2X1  g5809(.A(n6987), .B(n6985), .Y(n6988));
  NOR2X1  g5810(.A(n6988), .B(n5894), .Y(n6989));
  INVX1   g5811(.A(P2_REG1_REG_22__SCAN_IN), .Y(n6990));
  NOR3X1  g5812(.A(n5886), .B(n5881), .C(n6990), .Y(n6991));
  NAND3X1 g5813(.A(n5886), .B(n5881), .C(P2_REG2_REG_22__SCAN_IN), .Y(n6992));
  NAND3X1 g5814(.A(n5890), .B(n5881), .C(P2_REG0_REG_22__SCAN_IN), .Y(n6993));
  NAND2X1 g5815(.A(n6993), .B(n6992), .Y(n6994));
  NOR3X1  g5816(.A(n6994), .B(n6991), .C(n6989), .Y(n6995));
  OAI22X1 g5817(.A0(n6984), .A1(n5928), .B0(n5965), .B1(n6995), .Y(n6996));
  AOI21X1 g5818(.A0(n6983), .A1(n5924), .B0(n6996), .Y(n6997));
  OAI21X1 g5819(.A0(n6972), .A1(n5914), .B0(n6997), .Y(n6998));
  NOR2X1  g5820(.A(n6998), .B(n6981), .Y(n6999));
  NAND2X1 g5821(.A(n5862), .B(P2_REG0_REG_21__SCAN_IN), .Y(n7000));
  OAI21X1 g5822(.A0(n6999), .A1(n5862), .B0(n7000), .Y(P2_U3509));
  NOR2X1  g5823(.A(n5867), .B(n5643), .Y(n7002));
  XOR2X1  g5824(.A(n7002), .B(n6995), .Y(n7003));
  INVX1   g5825(.A(n6968), .Y(n7004));
  OAI21X1 g5826(.A0(n6909), .A1(n6921), .B0(n8727), .Y(n7006));
  AOI21X1 g5827(.A0(n7006), .A1(n7004), .B0(n6969), .Y(n7007));
  XOR2X1  g5828(.A(n7007), .B(n7003), .Y(n7008));
  NOR2X1  g5829(.A(n6954), .B(n6946), .Y(n7009));
  INVX1   g5830(.A(n7009), .Y(n7010));
  OAI22X1 g5831(.A0(n6964), .A1(n6965), .B0(n6915), .B1(n6865), .Y(n7011));
  NOR3X1  g5832(.A(n6947), .B(n5867), .C(n5633), .Y(n7012));
  AOI21X1 g5833(.A0(n7011), .A1(n7010), .B0(n7012), .Y(n7013));
  NOR3X1  g5834(.A(n7009), .B(n6915), .C(n6863), .Y(n7014));
  NAND2X1 g5835(.A(n7014), .B(n6810), .Y(n7015));
  NAND2X1 g5836(.A(n7015), .B(n7013), .Y(n7016));
  XOR2X1  g5837(.A(n7016), .B(n7003), .Y(n7017));
  OAI22X1 g5838(.A0(n6947), .A1(n6072), .B0(n6071), .B1(n7017), .Y(n7018));
  OAI22X1 g5839(.A0(n7017), .A1(n6097), .B0(n5904), .B1(n7017), .Y(n7022));
  NOR2X1  g5840(.A(n7022), .B(n7018), .Y(n7023));
  OAI21X1 g5841(.A0(n7008), .A1(n6128), .B0(n7023), .Y(n7024));
  NOR2X1  g5842(.A(n7008), .B(n5902), .Y(n7025));
  AOI21X1 g5843(.A0(n6631), .A1(n6630), .B0(n7008), .Y(n7026));
  NOR3X1  g5844(.A(n6954), .B(n6901), .C(n6937), .Y(n7027));
  INVX1   g5845(.A(n7002), .Y(n7028));
  XOR2X1  g5846(.A(n7028), .B(n7027), .Y(n7029));
  INVX1   g5847(.A(P2_REG3_REG_23__SCAN_IN), .Y(n7030));
  NOR3X1  g5848(.A(n6940), .B(n6985), .C(n6986), .Y(n7031));
  XOR2X1  g5849(.A(n7031), .B(n7030), .Y(n7032));
  INVX1   g5850(.A(n7032), .Y(n7033));
  AOI22X1 g5851(.A0(n5916), .A1(P2_REG2_REG_23__SCAN_IN), .B0(P2_REG0_REG_23__SCAN_IN), .B1(n5920), .Y(n7034));
  INVX1   g5852(.A(n7034), .Y(n7035));
  AOI21X1 g5853(.A0(n5917), .A1(P2_REG1_REG_23__SCAN_IN), .B0(n7035), .Y(n7036));
  INVX1   g5854(.A(n7036), .Y(n7037));
  AOI21X1 g5855(.A0(n7033), .A1(n5919), .B0(n7037), .Y(n7038));
  OAI22X1 g5856(.A0(n7028), .A1(n5928), .B0(n5965), .B1(n7038), .Y(n7039));
  AOI21X1 g5857(.A0(n7029), .A1(n5924), .B0(n7039), .Y(n7040));
  OAI21X1 g5858(.A0(n7017), .A1(n5914), .B0(n7040), .Y(n7041));
  NOR4X1  g5859(.A(n7026), .B(n7025), .C(n7024), .D(n7041), .Y(n7042));
  NAND2X1 g5860(.A(n5862), .B(P2_REG0_REG_22__SCAN_IN), .Y(n7043));
  OAI21X1 g5861(.A0(n7042), .A1(n5862), .B0(n7043), .Y(P2_U3510));
  INVX1   g5862(.A(n6995), .Y(n7045));
  NOR3X1  g5863(.A(n7045), .B(n5867), .C(n5643), .Y(n7046));
  INVX1   g5864(.A(n7046), .Y(n7047));
  NOR2X1  g5865(.A(n5867), .B(n5656), .Y(n7049));
  XOR2X1  g5866(.A(n7049), .B(n7038), .Y(n7050));
  INVX1   g5867(.A(n7050), .Y(n7051));
  NAND3X1 g5868(.A(n7051), .B(n8730), .C(n7047), .Y(n7052));
  INVX1   g5869(.A(n7038), .Y(n7053));
  NOR3X1  g5870(.A(n7053), .B(n5867), .C(n5656), .Y(n7054));
  OAI21X1 g5871(.A0(n3083), .A1(n1149), .B0(n5654), .Y(n7055));
  INVX1   g5872(.A(n5867), .Y(n7056));
  NAND2X1 g5873(.A(n7056), .B(n7055), .Y(n7057));
  AOI22X1 g5874(.A0(n7053), .A1(n7057), .B0(n7028), .B1(n7045), .Y(n7058));
  INVX1   g5875(.A(n7058), .Y(n7059));
  NOR2X1  g5876(.A(n7059), .B(n7054), .Y(n7060));
  OAI21X1 g5877(.A0(n7007), .A1(n7046), .B0(n7060), .Y(n7061));
  AOI21X1 g5878(.A0(n7061), .A1(n7052), .B0(n6128), .Y(n7062));
  NOR3X1  g5879(.A(n6995), .B(n5867), .C(n5643), .Y(n7063));
  OAI21X1 g5880(.A0(n5867), .A1(n5643), .B0(n6995), .Y(n7064));
  AOI21X1 g5881(.A0(n7064), .A1(n7016), .B0(n7063), .Y(n7065));
  XOR2X1  g5882(.A(n7065), .B(n7051), .Y(n7066));
  OAI22X1 g5883(.A0(n6995), .A1(n6072), .B0(n6071), .B1(n7066), .Y(n7067));
  OAI22X1 g5884(.A0(n7066), .A1(n6097), .B0(n5904), .B1(n7066), .Y(n7070));
  NOR3X1  g5885(.A(n7070), .B(n7067), .C(n7062), .Y(n7071));
  AOI21X1 g5886(.A0(n7061), .A1(n7052), .B0(n5902), .Y(n7072));
  AOI22X1 g5887(.A0(n7052), .A1(n7061), .B0(n6631), .B1(n6630), .Y(n7073));
  NOR2X1  g5888(.A(n7073), .B(n7072), .Y(n7074));
  NAND2X1 g5889(.A(n7074), .B(n7071), .Y(n7075));
  OAI21X1 g5890(.A0(n5867), .A1(n5643), .B0(n7027), .Y(n7076));
  XOR2X1  g5891(.A(n7049), .B(n7076), .Y(n7077));
  NOR4X1  g5892(.A(n6985), .B(n6986), .C(n7030), .D(n6940), .Y(n7078));
  XOR2X1  g5893(.A(n7078), .B(P2_REG3_REG_24__SCAN_IN), .Y(n7079));
  NAND3X1 g5894(.A(n5890), .B(n5889), .C(P2_REG1_REG_24__SCAN_IN), .Y(n7080));
  AOI22X1 g5895(.A0(n5916), .A1(P2_REG2_REG_24__SCAN_IN), .B0(P2_REG0_REG_24__SCAN_IN), .B1(n5920), .Y(n7081));
  NAND2X1 g5896(.A(n7081), .B(n7080), .Y(n7082));
  AOI21X1 g5897(.A0(n7079), .A1(n5919), .B0(n7082), .Y(n7083));
  OAI22X1 g5898(.A0(n7057), .A1(n5928), .B0(n5965), .B1(n7083), .Y(n7084));
  AOI21X1 g5899(.A0(n7077), .A1(n5924), .B0(n7084), .Y(n7085));
  OAI21X1 g5900(.A0(n7066), .A1(n5914), .B0(n7085), .Y(n7086));
  NOR2X1  g5901(.A(n7086), .B(n7075), .Y(n7087));
  NAND2X1 g5902(.A(n5862), .B(P2_REG0_REG_23__SCAN_IN), .Y(n7088));
  OAI21X1 g5903(.A0(n7087), .A1(n5862), .B0(n7088), .Y(P2_U3511));
  INVX1   g5904(.A(n7083), .Y(n7090));
  NAND2X1 g5905(.A(n7056), .B(n5664), .Y(n7091));
  XOR2X1  g5906(.A(n7091), .B(n7090), .Y(n7092));
  NAND2X1 g5907(.A(n7047), .B(n6969), .Y(n7094));
  NAND2X1 g5908(.A(n7094), .B(n7058), .Y(n7095));
  NOR3X1  g5909(.A(n7054), .B(n7046), .C(n6968), .Y(n7096));
  XOR2X1  g5910(.A(n8732), .B(n7092), .Y(n7098));
  INVX1   g5911(.A(n7098), .Y(n7099));
  NAND2X1 g5912(.A(n7099), .B(n5908), .Y(n7100));
  NOR3X1  g5913(.A(n7038), .B(n5867), .C(n5656), .Y(n7101));
  INVX1   g5914(.A(n7101), .Y(n7102));
  AOI21X1 g5915(.A0(n7056), .A1(n7055), .B0(n7053), .Y(n7103));
  OAI21X1 g5916(.A0(n7103), .A1(n7065), .B0(n7102), .Y(n7104));
  NAND2X1 g5917(.A(n7092), .B(n7104), .Y(n7107));
  OAI21X1 g5918(.A0(n7104), .A1(n7092), .B0(n7107), .Y(n7108));
  AOI22X1 g5919(.A0(n7053), .A1(n5959), .B0(n5910), .B1(n7108), .Y(n7109));
  AOI22X1 g5920(.A0(n7108), .A1(n5911), .B0(n5903), .B1(n7108), .Y(n7113));
  NAND3X1 g5921(.A(n7113), .B(n7109), .C(n7100), .Y(n7114));
  NOR2X1  g5922(.A(n7098), .B(n5902), .Y(n7115));
  AOI21X1 g5923(.A0(n6631), .A1(n6630), .B0(n7098), .Y(n7116));
  NAND4X1 g5924(.A(n5856), .B(n5852), .C(n5850), .D(n7108), .Y(n7117));
  NOR2X1  g5925(.A(n7049), .B(n7076), .Y(n7118));
  XOR2X1  g5926(.A(n7091), .B(n7118), .Y(n7119));
  NAND2X1 g5927(.A(n7078), .B(P2_REG3_REG_24__SCAN_IN), .Y(n7120));
  XOR2X1  g5928(.A(n7120), .B(P2_REG3_REG_25__SCAN_IN), .Y(n7121));
  INVX1   g5929(.A(n7121), .Y(n7122));
  AOI22X1 g5930(.A0(n5916), .A1(P2_REG2_REG_25__SCAN_IN), .B0(P2_REG0_REG_25__SCAN_IN), .B1(n5920), .Y(n7123));
  INVX1   g5931(.A(n7123), .Y(n7124));
  AOI21X1 g5932(.A0(n5917), .A1(P2_REG1_REG_25__SCAN_IN), .B0(n7124), .Y(n7125));
  INVX1   g5933(.A(n7125), .Y(n7126));
  AOI21X1 g5934(.A0(n7122), .A1(n5919), .B0(n7126), .Y(n7127));
  OAI22X1 g5935(.A0(n7091), .A1(n5928), .B0(n5965), .B1(n7127), .Y(n7128));
  AOI21X1 g5936(.A0(n7119), .A1(n5924), .B0(n7128), .Y(n7129));
  NAND2X1 g5937(.A(n7129), .B(n7117), .Y(n7130));
  NOR4X1  g5938(.A(n7116), .B(n7115), .C(n7114), .D(n7130), .Y(n7131));
  NAND2X1 g5939(.A(n5862), .B(P2_REG0_REG_24__SCAN_IN), .Y(n7132));
  OAI21X1 g5940(.A0(n7131), .A1(n5862), .B0(n7132), .Y(P2_U3512));
  NOR2X1  g5941(.A(n5867), .B(n5673), .Y(n7134));
  XOR2X1  g5942(.A(n7134), .B(n7127), .Y(n7135));
  NOR2X1  g5943(.A(n7091), .B(n7090), .Y(n7136));
  AOI21X1 g5944(.A0(n7056), .A1(n5664), .B0(n7083), .Y(n7138));
  NAND2X1 g5945(.A(n7095), .B(n8764), .Y(n7139));
  INVX1   g5946(.A(n7096), .Y(n7140));
  OAI21X1 g5947(.A0(n7140), .A1(n6959), .B0(n7139), .Y(n7141));
  AOI21X1 g5948(.A0(n7141), .A1(n8762), .B0(n7138), .Y(n7142));
  XOR2X1  g5949(.A(n7142), .B(n7135), .Y(n7143));
  NOR2X1  g5950(.A(n7143), .B(n6128), .Y(n7144));
  INVX1   g5951(.A(n7144), .Y(n7145));
  AOI21X1 g5952(.A0(n7056), .A1(n5664), .B0(n7090), .Y(n7146));
  INVX1   g5953(.A(n7146), .Y(n7147));
  NOR2X1  g5954(.A(n7091), .B(n7083), .Y(n7148));
  AOI21X1 g5955(.A0(n7147), .A1(n7104), .B0(n7148), .Y(n7149));
  NAND2X1 g5956(.A(n7149), .B(n7153), .Y(n7151));
  INVX1   g5957(.A(n7127), .Y(n7152));
  XOR2X1  g5958(.A(n7134), .B(n7152), .Y(n7153));
  OAI21X1 g5959(.A0(n7153), .A1(n7149), .B0(n7151), .Y(n7154));
  AOI22X1 g5960(.A0(n7090), .A1(n5959), .B0(n5910), .B1(n7154), .Y(n7155));
  AOI22X1 g5961(.A0(n7154), .A1(n5911), .B0(n5903), .B1(n7154), .Y(n7159));
  NAND3X1 g5962(.A(n7159), .B(n7155), .C(n7145), .Y(n7160));
  INVX1   g5963(.A(n7143), .Y(n7161));
  OAI21X1 g5964(.A0(n5907), .A1(n5900), .B0(n7161), .Y(n7162));
  OAI21X1 g5965(.A0(n7143), .A1(n5902), .B0(n7162), .Y(n7163));
  NAND4X1 g5966(.A(n5856), .B(n5852), .C(n5850), .D(n7154), .Y(n7164));
  INVX1   g5967(.A(n7091), .Y(n7165));
  NOR3X1  g5968(.A(n7165), .B(n7049), .C(n7076), .Y(n7166));
  INVX1   g5969(.A(n7134), .Y(n7167));
  XOR2X1  g5970(.A(n7167), .B(n7166), .Y(n7168));
  NAND3X1 g5971(.A(n7078), .B(P2_REG3_REG_24__SCAN_IN), .C(P2_REG3_REG_25__SCAN_IN), .Y(n7169));
  XOR2X1  g5972(.A(n7169), .B(P2_REG3_REG_26__SCAN_IN), .Y(n7170));
  INVX1   g5973(.A(n7170), .Y(n7171));
  AOI22X1 g5974(.A0(n5916), .A1(P2_REG2_REG_26__SCAN_IN), .B0(P2_REG0_REG_26__SCAN_IN), .B1(n5920), .Y(n7172));
  INVX1   g5975(.A(n7172), .Y(n7173));
  AOI21X1 g5976(.A0(n5917), .A1(P2_REG1_REG_26__SCAN_IN), .B0(n7173), .Y(n7174));
  INVX1   g5977(.A(n7174), .Y(n7175));
  AOI21X1 g5978(.A0(n7171), .A1(n5919), .B0(n7175), .Y(n7176));
  OAI22X1 g5979(.A0(n7167), .A1(n5928), .B0(n5965), .B1(n7176), .Y(n7177));
  AOI21X1 g5980(.A0(n7168), .A1(n5924), .B0(n7177), .Y(n7178));
  NAND2X1 g5981(.A(n7178), .B(n7164), .Y(n7179));
  NOR3X1  g5982(.A(n7179), .B(n7163), .C(n7160), .Y(n7180));
  NAND2X1 g5983(.A(n5862), .B(P2_REG0_REG_25__SCAN_IN), .Y(n7181));
  OAI21X1 g5984(.A0(n7180), .A1(n5862), .B0(n7181), .Y(P2_U3513));
  INVX1   g5985(.A(n7176), .Y(n7183));
  NOR2X1  g5986(.A(n5867), .B(n5681), .Y(n7184));
  XOR2X1  g5987(.A(n7184), .B(n7183), .Y(n7185));
  NOR3X1  g5988(.A(n7152), .B(n5867), .C(n5673), .Y(n7186));
  OAI21X1 g5989(.A0(n3177), .A1(n1149), .B0(n5671), .Y(n7187));
  AOI21X1 g5990(.A0(n7056), .A1(n7187), .B0(n7127), .Y(n7188));
  OAI21X1 g5991(.A0(n7142), .A1(n7186), .B0(n8758), .Y(n7190));
  XOR2X1  g5992(.A(n7190), .B(n7185), .Y(n7191));
  INVX1   g5993(.A(n7191), .Y(n7192));
  NAND2X1 g5994(.A(n7192), .B(n5908), .Y(n7193));
  OAI21X1 g5995(.A0(n5867), .A1(n5673), .B0(n7127), .Y(n7194));
  OAI21X1 g5996(.A0(n7184), .A1(n7183), .B0(n7194), .Y(n7195));
  NOR3X1  g5997(.A(n7176), .B(n5867), .C(n5681), .Y(n7196));
  NOR2X1  g5998(.A(n7196), .B(n7195), .Y(n7197));
  NOR3X1  g5999(.A(n7127), .B(n5867), .C(n5673), .Y(n7198));
  INVX1   g6000(.A(n7198), .Y(n7199));
  NAND2X1 g6001(.A(n7199), .B(n7149), .Y(n7200));
  NOR2X1  g6002(.A(n7185), .B(n7198), .Y(n7201));
  INVX1   g6003(.A(n7201), .Y(n7202));
  AOI21X1 g6004(.A0(n7056), .A1(n7187), .B0(n7152), .Y(n7203));
  NOR2X1  g6005(.A(n7203), .B(n7149), .Y(n7204));
  NOR2X1  g6006(.A(n7204), .B(n7202), .Y(n7205));
  AOI21X1 g6007(.A0(n7200), .A1(n7197), .B0(n7205), .Y(n7206));
  AOI22X1 g6008(.A0(n7152), .A1(n5959), .B0(n5910), .B1(n7206), .Y(n7207));
  AOI22X1 g6009(.A0(n7206), .A1(n5911), .B0(n5903), .B1(n7206), .Y(n7212));
  NAND3X1 g6010(.A(n7212), .B(n7207), .C(n7193), .Y(n7213));
  NOR2X1  g6011(.A(n7191), .B(n5902), .Y(n7214));
  AOI21X1 g6012(.A0(n6631), .A1(n6630), .B0(n7191), .Y(n7215));
  NAND4X1 g6013(.A(n5856), .B(n5852), .C(n5850), .D(n7206), .Y(n7216));
  NOR4X1  g6014(.A(n7165), .B(n7049), .C(n7076), .D(n7134), .Y(n7217));
  OAI21X1 g6015(.A0(n3264), .A1(n1149), .B0(n5679), .Y(n7218));
  NAND2X1 g6016(.A(n7056), .B(n7218), .Y(n7219));
  XOR2X1  g6017(.A(n7219), .B(n7217), .Y(n7220));
  NAND4X1 g6018(.A(P2_REG3_REG_26__SCAN_IN), .B(P2_REG3_REG_24__SCAN_IN), .C(P2_REG3_REG_25__SCAN_IN), .D(n7078), .Y(n7221));
  XOR2X1  g6019(.A(n7221), .B(P2_REG3_REG_27__SCAN_IN), .Y(n7222));
  INVX1   g6020(.A(n7222), .Y(n7223));
  AOI22X1 g6021(.A0(n5916), .A1(P2_REG2_REG_27__SCAN_IN), .B0(P2_REG0_REG_27__SCAN_IN), .B1(n5920), .Y(n7224));
  INVX1   g6022(.A(n7224), .Y(n7225));
  AOI21X1 g6023(.A0(n5917), .A1(P2_REG1_REG_27__SCAN_IN), .B0(n7225), .Y(n7226));
  INVX1   g6024(.A(n7226), .Y(n7227));
  AOI21X1 g6025(.A0(n7223), .A1(n5919), .B0(n7227), .Y(n7228));
  OAI22X1 g6026(.A0(n7219), .A1(n5928), .B0(n5965), .B1(n7228), .Y(n7229));
  AOI21X1 g6027(.A0(n7220), .A1(n5924), .B0(n7229), .Y(n7230));
  NAND2X1 g6028(.A(n7230), .B(n7216), .Y(n7231));
  NOR4X1  g6029(.A(n7215), .B(n7214), .C(n7213), .D(n7231), .Y(n7232));
  NAND2X1 g6030(.A(n5862), .B(P2_REG0_REG_26__SCAN_IN), .Y(n7233));
  OAI21X1 g6031(.A0(n7232), .A1(n5862), .B0(n7233), .Y(P2_U3514));
  AOI21X1 g6032(.A0(n7056), .A1(n7218), .B0(n7176), .Y(n7235));
  INVX1   g6033(.A(n7235), .Y(n7236));
  INVX1   g6034(.A(n7138), .Y(n7238));
  AOI21X1 g6035(.A0(n8733), .A1(n8756), .B0(n7188), .Y(n7240));
  NAND3X1 g6036(.A(n7176), .B(n7056), .C(n7218), .Y(n7241));
  INVX1   g6037(.A(n7228), .Y(n7242));
  OAI21X1 g6038(.A0(n5694), .A1(n5692), .B0(n7056), .Y(n7243));
  XOR2X1  g6039(.A(n7243), .B(n7242), .Y(n7244));
  NAND2X1 g6040(.A(n8904), .B(n7241), .Y(n7246));
  AOI21X1 g6041(.A0(n7240), .A1(n7236), .B0(n7246), .Y(n7247));
  NAND2X1 g6042(.A(n7244), .B(n7236), .Y(n7248));
  AOI21X1 g6043(.A0(n7190), .A1(n7241), .B0(n7248), .Y(n7249));
  OAI21X1 g6044(.A0(n7249), .A1(n7247), .B0(n5908), .Y(n7250));
  INVX1   g6045(.A(n7196), .Y(n7251));
  AOI21X1 g6046(.A0(n7219), .A1(n7176), .B0(n7203), .Y(n7252));
  OAI21X1 g6047(.A0(n7198), .A1(n7148), .B0(n7252), .Y(n7253));
  NAND3X1 g6048(.A(n7252), .B(n7147), .C(n7104), .Y(n7254));
  NAND3X1 g6049(.A(n7254), .B(n7253), .C(n7251), .Y(n7255));
  XOR2X1  g6050(.A(n7255), .B(n8904), .Y(n7256));
  AOI22X1 g6051(.A0(n7183), .A1(n5959), .B0(n5910), .B1(n7256), .Y(n7257));
  NOR2X1  g6052(.A(n7198), .B(n7148), .Y(n7258));
  NOR2X1  g6053(.A(n7258), .B(n7195), .Y(n7259));
  AOI22X1 g6054(.A0(n7256), .A1(n5911), .B0(n5903), .B1(n7256), .Y(n7265));
  NAND3X1 g6055(.A(n7265), .B(n7257), .C(n7250), .Y(n7266));
  NOR2X1  g6056(.A(n7249), .B(n7247), .Y(n7267));
  NOR2X1  g6057(.A(n7267), .B(n5902), .Y(n7268));
  AOI21X1 g6058(.A0(n6631), .A1(n6630), .B0(n7267), .Y(n7269));
  NAND4X1 g6059(.A(n5856), .B(n5852), .C(n5850), .D(n7256), .Y(n7270));
  NAND2X1 g6060(.A(n7219), .B(n7217), .Y(n7271));
  NOR2X1  g6061(.A(n5867), .B(n5695), .Y(n7272));
  XOR2X1  g6062(.A(n7272), .B(n7271), .Y(n7273));
  INVX1   g6063(.A(P2_REG3_REG_28__SCAN_IN), .Y(n7274));
  INVX1   g6064(.A(P2_REG3_REG_27__SCAN_IN), .Y(n7275));
  NOR2X1  g6065(.A(n7221), .B(n7275), .Y(n7276));
  XOR2X1  g6066(.A(n7276), .B(n7274), .Y(n7277));
  INVX1   g6067(.A(n7277), .Y(n7278));
  AOI22X1 g6068(.A0(n5916), .A1(P2_REG2_REG_28__SCAN_IN), .B0(P2_REG0_REG_28__SCAN_IN), .B1(n5920), .Y(n7279));
  INVX1   g6069(.A(n7279), .Y(n7280));
  AOI21X1 g6070(.A0(n5917), .A1(P2_REG1_REG_28__SCAN_IN), .B0(n7280), .Y(n7281));
  INVX1   g6071(.A(n7281), .Y(n7282));
  AOI21X1 g6072(.A0(n7278), .A1(n5919), .B0(n7282), .Y(n7283));
  OAI22X1 g6073(.A0(n7243), .A1(n5928), .B0(n5965), .B1(n7283), .Y(n7284));
  AOI21X1 g6074(.A0(n7273), .A1(n5924), .B0(n7284), .Y(n7285));
  NAND2X1 g6075(.A(n7285), .B(n7270), .Y(n7286));
  NOR4X1  g6076(.A(n7269), .B(n7268), .C(n7266), .D(n7286), .Y(n7287));
  NAND2X1 g6077(.A(n5862), .B(P2_REG0_REG_27__SCAN_IN), .Y(n7288));
  OAI21X1 g6078(.A0(n7287), .A1(n5862), .B0(n7288), .Y(P2_U3515));
  NOR2X1  g6079(.A(n5867), .B(n5704), .Y(n7290));
  XOR2X1  g6080(.A(n7290), .B(n7283), .Y(n7291));
  INVX1   g6081(.A(n7291), .Y(n7292));
  NOR2X1  g6082(.A(n7272), .B(n7242), .Y(n7293));
  NAND2X1 g6083(.A(n7243), .B(n7228), .Y(n7294));
  NOR2X1  g6084(.A(n7243), .B(n7228), .Y(n7295));
  AOI21X1 g6085(.A0(n7294), .A1(n7259), .B0(n7295), .Y(n7296));
  OAI21X1 g6086(.A0(n7293), .A1(n7251), .B0(n7296), .Y(n7297));
  NAND2X1 g6087(.A(n7252), .B(n7104), .Y(n7298));
  NOR3X1  g6088(.A(n7298), .B(n7293), .C(n7146), .Y(n7299));
  NOR2X1  g6089(.A(n7299), .B(n7297), .Y(n7300));
  XOR2X1  g6090(.A(n7300), .B(n7292), .Y(n7301));
  OAI22X1 g6091(.A0(n7228), .A1(n6072), .B0(n6071), .B1(n7301), .Y(n7302));
  OAI22X1 g6092(.A0(n7301), .A1(n6097), .B0(n5904), .B1(n7301), .Y(n7306));
  NOR2X1  g6093(.A(n7306), .B(n7302), .Y(n7307));
  AOI22X1 g6094(.A0(n7228), .A1(n7272), .B0(n7184), .B1(n7176), .Y(n7308));
  OAI21X1 g6095(.A0(n7242), .A1(n7235), .B0(n7243), .Y(n7309));
  OAI21X1 g6096(.A0(n7228), .A1(n7236), .B0(n7309), .Y(n7310));
  AOI21X1 g6097(.A0(n7308), .A1(n7190), .B0(n7310), .Y(n7311));
  XOR2X1  g6098(.A(n7311), .B(n7291), .Y(n7312));
  AOI21X1 g6099(.A0(n6128), .A1(n6631), .B0(n7312), .Y(n7313));
  AOI21X1 g6100(.A0(n5902), .A1(n6630), .B0(n7312), .Y(n7314));
  NOR2X1  g6101(.A(n7314), .B(n7313), .Y(n7315));
  NAND2X1 g6102(.A(n7315), .B(n7307), .Y(n7316));
  NOR2X1  g6103(.A(n7301), .B(n5914), .Y(n7317));
  NOR2X1  g6104(.A(n7272), .B(n7271), .Y(n7318));
  XOR2X1  g6105(.A(n7290), .B(n7318), .Y(n7319));
  NOR4X1  g6106(.A(n5894), .B(n7274), .C(n7275), .D(n7221), .Y(n7320));
  NAND3X1 g6107(.A(n5890), .B(n5881), .C(P2_REG0_REG_29__SCAN_IN), .Y(n7321));
  INVX1   g6108(.A(n7321), .Y(n7322));
  AOI22X1 g6109(.A0(n5916), .A1(P2_REG2_REG_29__SCAN_IN), .B0(P2_REG1_REG_29__SCAN_IN), .B1(n5917), .Y(n7323));
  INVX1   g6110(.A(n7323), .Y(n7324));
  NOR3X1  g6111(.A(n7324), .B(n7322), .C(n7320), .Y(n7325));
  INVX1   g6112(.A(n7325), .Y(n7326));
  AOI22X1 g6113(.A0(n7290), .A1(n6060), .B0(n5915), .B1(n7326), .Y(n7327));
  OAI21X1 g6114(.A0(n7319), .A1(n5925), .B0(n7327), .Y(n7328));
  NOR3X1  g6115(.A(n7328), .B(n7317), .C(n7316), .Y(n7329));
  NAND2X1 g6116(.A(n5862), .B(P2_REG0_REG_28__SCAN_IN), .Y(n7330));
  OAI21X1 g6117(.A0(n7329), .A1(n5862), .B0(n7330), .Y(P2_U3516));
  OAI21X1 g6118(.A0(n3343), .A1(n3341), .B0(n1156), .Y(n7332));
  AOI21X1 g6119(.A0(n5710), .A1(n7332), .B0(n5867), .Y(n7333));
  XOR2X1  g6120(.A(n7333), .B(n7325), .Y(n7334));
  OAI21X1 g6121(.A0(n3322), .A1(n1149), .B0(n5702), .Y(n7335));
  NAND2X1 g6122(.A(n7056), .B(n7335), .Y(n7336));
  NAND2X1 g6123(.A(n7272), .B(n7242), .Y(n7337));
  OAI21X1 g6124(.A0(n7293), .A1(n7253), .B0(n7337), .Y(n7338));
  AOI21X1 g6125(.A0(n7294), .A1(n7196), .B0(n7338), .Y(n7339));
  NAND4X1 g6126(.A(n7252), .B(n7147), .C(n7104), .D(n7294), .Y(n7340));
  AOI21X1 g6127(.A0(n7340), .A1(n7339), .B0(n7336), .Y(n7341));
  AOI21X1 g6128(.A0(n7300), .A1(n7336), .B0(n7283), .Y(n7342));
  NOR3X1  g6129(.A(n7342), .B(n7341), .C(n7334), .Y(n7343));
  XOR2X1  g6130(.A(n7333), .B(n7326), .Y(n7344));
  OAI21X1 g6131(.A0(n7299), .A1(n7297), .B0(n7290), .Y(n7345));
  INVX1   g6132(.A(n7283), .Y(n7346));
  NAND2X1 g6133(.A(n7340), .B(n7339), .Y(n7347));
  OAI21X1 g6134(.A0(n7347), .A1(n7290), .B0(n7346), .Y(n7348));
  AOI21X1 g6135(.A0(n7348), .A1(n7345), .B0(n7344), .Y(n7349));
  OAI22X1 g6136(.A0(n7343), .A1(n7349), .B0(n5911), .B1(n5910), .Y(n7350));
  AOI21X1 g6137(.A0(n7056), .A1(n7335), .B0(n7283), .Y(n7351));
  INVX1   g6138(.A(n7308), .Y(n7352));
  INVX1   g6139(.A(n7310), .Y(n7353));
  OAI21X1 g6140(.A0(n7352), .A1(n7240), .B0(n7353), .Y(n7354));
  NOR3X1  g6141(.A(n7344), .B(n7354), .C(n7351), .Y(n7355));
  NOR3X1  g6142(.A(n7346), .B(n5867), .C(n5704), .Y(n7356));
  NOR2X1  g6143(.A(n7334), .B(n7356), .Y(n7357));
  NAND2X1 g6144(.A(n7357), .B(n7354), .Y(n7358));
  NOR2X1  g6145(.A(n7334), .B(n8750), .Y(n7360));
  NOR3X1  g6146(.A(n7344), .B(n7336), .C(n7346), .Y(n7361));
  NOR2X1  g6147(.A(n7361), .B(n7360), .Y(n7362));
  NAND2X1 g6148(.A(n7362), .B(n7358), .Y(n7363));
  OAI22X1 g6149(.A0(n7355), .A1(n7363), .B0(n5908), .B1(n5901), .Y(n7364));
  NAND2X1 g6150(.A(n7364), .B(n7350), .Y(n7365));
  NOR3X1  g6151(.A(n7334), .B(n7311), .C(n7356), .Y(n7366));
  NOR4X1  g6152(.A(n7360), .B(n7366), .C(n7355), .D(n7361), .Y(n7367));
  NOR2X1  g6153(.A(n5848), .B(n5850), .Y(n7368));
  INVX1   g6154(.A(n7368), .Y(n7369));
  INVX1   g6155(.A(P2_B_REG_SCAN_IN), .Y(n7370));
  OAI21X1 g6156(.A0(n5869), .A1(n7370), .B0(n5871), .Y(n7371));
  NAND3X1 g6157(.A(n5886), .B(n5881), .C(P2_REG2_REG_30__SCAN_IN), .Y(n7372));
  NAND3X1 g6158(.A(n5890), .B(n5881), .C(P2_REG0_REG_30__SCAN_IN), .Y(n7373));
  NAND2X1 g6159(.A(n7373), .B(n7372), .Y(n7374));
  AOI21X1 g6160(.A0(n5917), .A1(P2_REG1_REG_30__SCAN_IN), .B0(n7374), .Y(n7375));
  NOR3X1  g6161(.A(n7375), .B(n7371), .C(n7369), .Y(n7376));
  AOI21X1 g6162(.A0(n7346), .A1(n5959), .B0(n7376), .Y(n7377));
  OAI21X1 g6163(.A0(n7367), .A1(n6630), .B0(n7377), .Y(n7378));
  NOR2X1  g6164(.A(n7342), .B(n7341), .Y(n7381));
  XOR2X1  g6165(.A(n7381), .B(n7344), .Y(n7382));
  OAI22X1 g6166(.A0(n7367), .A1(n6631), .B0(n5904), .B1(n7382), .Y(n7383));
  NOR3X1  g6167(.A(n7290), .B(n7272), .C(n7271), .Y(n7384));
  NAND2X1 g6168(.A(n5710), .B(n7332), .Y(n7385));
  NAND2X1 g6169(.A(n7056), .B(n7385), .Y(n7386));
  XOR2X1  g6170(.A(n7386), .B(n7384), .Y(n7387));
  AOI22X1 g6171(.A0(n7333), .A1(n6060), .B0(n5924), .B1(n7387), .Y(n7388));
  OAI21X1 g6172(.A0(n7382), .A1(n5914), .B0(n7388), .Y(n7389));
  NOR4X1  g6173(.A(n7383), .B(n7378), .C(n7365), .D(n7389), .Y(n7390));
  NAND2X1 g6174(.A(n5862), .B(P2_REG0_REG_29__SCAN_IN), .Y(n7391));
  OAI21X1 g6175(.A0(n7390), .A1(n5862), .B0(n7391), .Y(P2_U3517));
  NOR4X1  g6176(.A(n7290), .B(n7272), .C(n7271), .D(n7333), .Y(n7393));
  OAI21X1 g6177(.A0(n5720), .A1(n5718), .B0(n7056), .Y(n7394));
  XOR2X1  g6178(.A(n7394), .B(n7393), .Y(n7395));
  NAND3X1 g6179(.A(n5886), .B(n5881), .C(P2_REG2_REG_31__SCAN_IN), .Y(n7396));
  NAND3X1 g6180(.A(n5890), .B(n5881), .C(P2_REG0_REG_31__SCAN_IN), .Y(n7397));
  NAND2X1 g6181(.A(n7397), .B(n7396), .Y(n7398));
  AOI21X1 g6182(.A0(n5917), .A1(P2_REG1_REG_31__SCAN_IN), .B0(n7398), .Y(n7399));
  NOR3X1  g6183(.A(n7399), .B(n7371), .C(n7369), .Y(n7400));
  INVX1   g6184(.A(n7400), .Y(n7401));
  OAI21X1 g6185(.A0(n7394), .A1(n5928), .B0(n7401), .Y(n7402));
  AOI21X1 g6186(.A0(n7395), .A1(n5924), .B0(n7402), .Y(n7403));
  NAND2X1 g6187(.A(n5862), .B(P2_REG0_REG_30__SCAN_IN), .Y(n7404));
  OAI21X1 g6188(.A0(n7403), .A1(n5862), .B0(n7404), .Y(P2_U3518));
  INVX1   g6189(.A(n7393), .Y(n7406));
  NOR2X1  g6190(.A(n5867), .B(n5721), .Y(n7407));
  NOR2X1  g6191(.A(n7407), .B(n7406), .Y(n7408));
  NAND2X1 g6192(.A(n7056), .B(n5728), .Y(n7409));
  XOR2X1  g6193(.A(n7409), .B(n7408), .Y(n7410));
  OAI21X1 g6194(.A0(n7409), .A1(n5928), .B0(n7401), .Y(n7411));
  AOI21X1 g6195(.A0(n7410), .A1(n5924), .B0(n7411), .Y(n7412));
  NAND2X1 g6196(.A(n5862), .B(P2_REG0_REG_31__SCAN_IN), .Y(n7413));
  OAI21X1 g6197(.A0(n7412), .A1(n5862), .B0(n7413), .Y(P2_U3519));
  INVX1   g6198(.A(n5861), .Y(n7415));
  NAND4X1 g6199(.A(n5859), .B(n5837), .C(n5743), .D(n7415), .Y(n7416));
  NAND2X1 g6200(.A(n7416), .B(P2_REG1_REG_0__SCAN_IN), .Y(n7417));
  OAI21X1 g6201(.A0(n7416), .A1(n5932), .B0(n7417), .Y(P2_U3520));
  NAND2X1 g6202(.A(n7416), .B(P2_REG1_REG_1__SCAN_IN), .Y(n7419));
  OAI21X1 g6203(.A0(n7416), .A1(n5978), .B0(n7419), .Y(P2_U3521));
  NAND2X1 g6204(.A(n7416), .B(P2_REG1_REG_2__SCAN_IN), .Y(n7421));
  OAI21X1 g6205(.A0(n7416), .A1(n6019), .B0(n7421), .Y(P2_U3522));
  NAND2X1 g6206(.A(n7416), .B(P2_REG1_REG_3__SCAN_IN), .Y(n7423));
  OAI21X1 g6207(.A0(n7416), .A1(n6068), .B0(n7423), .Y(P2_U3523));
  NAND2X1 g6208(.A(n7416), .B(P2_REG1_REG_4__SCAN_IN), .Y(n7425));
  OAI21X1 g6209(.A0(n7416), .A1(n6125), .B0(n7425), .Y(P2_U3524));
  NAND2X1 g6210(.A(n7416), .B(P2_REG1_REG_5__SCAN_IN), .Y(n7427));
  OAI21X1 g6211(.A0(n7416), .A1(n6176), .B0(n7427), .Y(P2_U3525));
  NAND2X1 g6212(.A(n7416), .B(P2_REG1_REG_6__SCAN_IN), .Y(n7429));
  OAI21X1 g6213(.A0(n7416), .A1(n6227), .B0(n7429), .Y(P2_U3526));
  NAND2X1 g6214(.A(n7416), .B(P2_REG1_REG_7__SCAN_IN), .Y(n7431));
  OAI21X1 g6215(.A0(n7416), .A1(n6279), .B0(n7431), .Y(P2_U3527));
  NAND2X1 g6216(.A(n7416), .B(P2_REG1_REG_8__SCAN_IN), .Y(n7433));
  OAI21X1 g6217(.A0(n7416), .A1(n6331), .B0(n7433), .Y(P2_U3528));
  NAND2X1 g6218(.A(n7416), .B(P2_REG1_REG_9__SCAN_IN), .Y(n7435));
  OAI21X1 g6219(.A0(n7416), .A1(n6378), .B0(n7435), .Y(P2_U3529));
  NAND2X1 g6220(.A(n7416), .B(P2_REG1_REG_10__SCAN_IN), .Y(n7437));
  OAI21X1 g6221(.A0(n7416), .A1(n6434), .B0(n7437), .Y(P2_U3530));
  NAND2X1 g6222(.A(n7416), .B(P2_REG1_REG_11__SCAN_IN), .Y(n7439));
  OAI21X1 g6223(.A0(n7416), .A1(n6498), .B0(n7439), .Y(P2_U3531));
  NAND2X1 g6224(.A(n7416), .B(P2_REG1_REG_12__SCAN_IN), .Y(n7441));
  OAI21X1 g6225(.A0(n7416), .A1(n6550), .B0(n7441), .Y(P2_U3532));
  NAND2X1 g6226(.A(n7416), .B(P2_REG1_REG_13__SCAN_IN), .Y(n7443));
  OAI21X1 g6227(.A0(n7416), .A1(n6601), .B0(n7443), .Y(P2_U3533));
  NAND2X1 g6228(.A(n7416), .B(P2_REG1_REG_14__SCAN_IN), .Y(n7445));
  OAI21X1 g6229(.A0(n7416), .A1(n6650), .B0(n7445), .Y(P2_U3534));
  NAND2X1 g6230(.A(n7416), .B(P2_REG1_REG_15__SCAN_IN), .Y(n7447));
  OAI21X1 g6231(.A0(n7416), .A1(n6694), .B0(n7447), .Y(P2_U3535));
  NAND2X1 g6232(.A(n7416), .B(P2_REG1_REG_16__SCAN_IN), .Y(n7449));
  OAI21X1 g6233(.A0(n7416), .A1(n6744), .B0(n7449), .Y(P2_U3536));
  NAND2X1 g6234(.A(n7416), .B(P2_REG1_REG_17__SCAN_IN), .Y(n7451));
  OAI21X1 g6235(.A0(n7416), .A1(n6803), .B0(n7451), .Y(P2_U3537));
  NAND2X1 g6236(.A(n7416), .B(P2_REG1_REG_18__SCAN_IN), .Y(n7453));
  OAI21X1 g6237(.A0(n7416), .A1(n6850), .B0(n7453), .Y(P2_U3538));
  NAND2X1 g6238(.A(n7416), .B(P2_REG1_REG_19__SCAN_IN), .Y(n7455));
  OAI21X1 g6239(.A0(n7416), .A1(n6898), .B0(n7455), .Y(P2_U3539));
  NAND2X1 g6240(.A(n7416), .B(P2_REG1_REG_20__SCAN_IN), .Y(n7457));
  OAI21X1 g6241(.A0(n7416), .A1(n6951), .B0(n7457), .Y(P2_U3540));
  NAND2X1 g6242(.A(n7416), .B(P2_REG1_REG_21__SCAN_IN), .Y(n7459));
  OAI21X1 g6243(.A0(n7416), .A1(n6999), .B0(n7459), .Y(P2_U3541));
  NAND2X1 g6244(.A(n7416), .B(P2_REG1_REG_22__SCAN_IN), .Y(n7461));
  OAI21X1 g6245(.A0(n7416), .A1(n7042), .B0(n7461), .Y(P2_U3542));
  NAND2X1 g6246(.A(n7416), .B(P2_REG1_REG_23__SCAN_IN), .Y(n7463));
  OAI21X1 g6247(.A0(n7416), .A1(n7087), .B0(n7463), .Y(P2_U3543));
  NAND2X1 g6248(.A(n7416), .B(P2_REG1_REG_24__SCAN_IN), .Y(n7465));
  OAI21X1 g6249(.A0(n7416), .A1(n7131), .B0(n7465), .Y(P2_U3544));
  NAND2X1 g6250(.A(n7416), .B(P2_REG1_REG_25__SCAN_IN), .Y(n7467));
  OAI21X1 g6251(.A0(n7416), .A1(n7180), .B0(n7467), .Y(P2_U3545));
  NAND2X1 g6252(.A(n7416), .B(P2_REG1_REG_26__SCAN_IN), .Y(n7469));
  OAI21X1 g6253(.A0(n7416), .A1(n7232), .B0(n7469), .Y(P2_U3546));
  NAND2X1 g6254(.A(n7416), .B(P2_REG1_REG_27__SCAN_IN), .Y(n7471));
  OAI21X1 g6255(.A0(n7416), .A1(n7287), .B0(n7471), .Y(P2_U3547));
  NAND2X1 g6256(.A(n7416), .B(P2_REG1_REG_28__SCAN_IN), .Y(n7473));
  OAI21X1 g6257(.A0(n7416), .A1(n7329), .B0(n7473), .Y(P2_U3548));
  NAND2X1 g6258(.A(n7416), .B(P2_REG1_REG_29__SCAN_IN), .Y(n7475));
  OAI21X1 g6259(.A0(n7416), .A1(n7390), .B0(n7475), .Y(P2_U3549));
  NAND2X1 g6260(.A(n7416), .B(P2_REG1_REG_30__SCAN_IN), .Y(n7477));
  OAI21X1 g6261(.A0(n7416), .A1(n7403), .B0(n7477), .Y(P2_U3550));
  NAND2X1 g6262(.A(n7416), .B(P2_REG1_REG_31__SCAN_IN), .Y(n7479));
  OAI21X1 g6263(.A0(n7416), .A1(n7412), .B0(n7479), .Y(P2_U3551));
  NOR4X1  g6264(.A(n5853), .B(n5847), .C(n5843), .D(n5855), .Y(n7481));
  INVX1   g6265(.A(n7481), .Y(n7482));
  INVX1   g6266(.A(n5837), .Y(n7483));
  OAI21X1 g6267(.A0(n5856), .A1(n5853), .B0(n7368), .Y(n7484));
  INVX1   g6268(.A(n7484), .Y(n7485));
  NOR4X1  g6269(.A(n7415), .B(n5840), .C(n7483), .D(n7485), .Y(n7486));
  INVX1   g6270(.A(n7486), .Y(n7487));
  AOI21X1 g6271(.A0(n7487), .A1(n7482), .B0(n5750), .Y(n7488));
  INVX1   g6272(.A(n7488), .Y(n7489));
  NOR2X1  g6273(.A(n7489), .B(n5965), .Y(n7490));
  NAND2X1 g6274(.A(n7488), .B(n5913), .Y(n7491));
  OAI21X1 g6275(.A0(n7488), .A1(n5879), .B0(n7491), .Y(n7492));
  AOI21X1 g6276(.A0(n7490), .A1(n5922), .B0(n7492), .Y(n7493));
  NAND3X1 g6277(.A(n5853), .B(n5848), .C(n5850), .Y(n7494));
  NOR2X1  g6278(.A(n7494), .B(n7489), .Y(n7495));
  NOR4X1  g6279(.A(n5742), .B(n5735), .C(P2_U3152), .D(n7482), .Y(n7496));
  AOI22X1 g6280(.A0(n7495), .A1(n5877), .B0(P2_REG3_REG_0__SCAN_IN), .B1(n7496), .Y(n7497));
  NOR3X1  g6281(.A(n7489), .B(n5925), .C(n5856), .Y(n7498));
  NOR4X1  g6282(.A(n5855), .B(n5853), .C(n5848), .D(n7489), .Y(n7499));
  AOI22X1 g6283(.A0(n7498), .A1(n5877), .B0(n8912), .B1(n7499), .Y(n7500));
  NAND3X1 g6284(.A(n7500), .B(n7497), .C(n7493), .Y(P2_U3296));
  NAND2X1 g6285(.A(n7488), .B(n5962), .Y(n7502));
  OAI21X1 g6286(.A0(n7488), .A1(n5949), .B0(n7502), .Y(n7503));
  AOI21X1 g6287(.A0(n7490), .A1(n5995), .B0(n7503), .Y(n7504));
  AOI22X1 g6288(.A0(n7495), .A1(n5939), .B0(P2_REG3_REG_1__SCAN_IN), .B1(n7496), .Y(n7505));
  AOI22X1 g6289(.A0(n7498), .A1(n5964), .B0(n5943), .B1(n7499), .Y(n7506));
  NAND3X1 g6290(.A(n7506), .B(n7505), .C(n7504), .Y(P2_U3295));
  AOI22X1 g6291(.A0(n7496), .A1(P2_REG3_REG_2__SCAN_IN), .B0(n5997), .B1(n7499), .Y(n7508));
  AOI22X1 g6292(.A0(n7495), .A1(n6046), .B0(n6009), .B1(n7498), .Y(n7509));
  NAND2X1 g6293(.A(n7488), .B(n6006), .Y(n7510));
  AOI22X1 g6294(.A0(n7489), .A1(P2_REG2_REG_2__SCAN_IN), .B0(n6028), .B1(n7490), .Y(n7511));
  NAND4X1 g6295(.A(n7510), .B(n7509), .C(n7508), .D(n7511), .Y(P2_U3294));
  NAND2X1 g6296(.A(n7488), .B(n6056), .Y(n7513));
  AOI22X1 g6297(.A0(n7489), .A1(P2_REG2_REG_3__SCAN_IN), .B0(n6065), .B1(n7490), .Y(n7514));
  AOI22X1 g6298(.A0(n7496), .A1(n6026), .B0(n6040), .B1(n7499), .Y(n7515));
  NOR4X1  g6299(.A(n6059), .B(n5925), .C(n5856), .D(n7489), .Y(n7516));
  AOI21X1 g6300(.A0(n7495), .A1(n6033), .B0(n7516), .Y(n7517));
  NAND4X1 g6301(.A(n7515), .B(n7514), .C(n7513), .D(n7517), .Y(P2_U3293));
  NOR3X1  g6302(.A(n6109), .B(n6098), .C(n6096), .Y(n7519));
  INVX1   g6303(.A(n7490), .Y(n7520));
  OAI22X1 g6304(.A0(n7488), .A1(n6087), .B0(n6121), .B1(n7520), .Y(n7521));
  INVX1   g6305(.A(n7496), .Y(n7522));
  INVX1   g6306(.A(n7499), .Y(n7523));
  OAI22X1 g6307(.A0(n7522), .A1(n6062), .B0(n6095), .B1(n7523), .Y(n7524));
  INVX1   g6308(.A(n7495), .Y(n7525));
  NAND4X1 g6309(.A(n6113), .B(n5924), .C(n5855), .D(n7488), .Y(n7526));
  OAI21X1 g6310(.A0(n7525), .A1(n6077), .B0(n7526), .Y(n7527));
  NOR3X1  g6311(.A(n7527), .B(n7524), .C(n7521), .Y(n7528));
  OAI21X1 g6312(.A0(n7489), .A1(n7519), .B0(n7528), .Y(P2_U3292));
  OAI22X1 g6313(.A0(n7488), .A1(n6114), .B0(n6172), .B1(n7520), .Y(n7530));
  OAI22X1 g6314(.A0(n7522), .A1(n6119), .B0(n6153), .B1(n7523), .Y(n7531));
  NAND4X1 g6315(.A(n6162), .B(n5924), .C(n5855), .D(n7488), .Y(n7532));
  OAI21X1 g6316(.A0(n7525), .A1(n6142), .B0(n7532), .Y(n7533));
  NOR3X1  g6317(.A(n7533), .B(n7531), .C(n7530), .Y(n7534));
  OAI21X1 g6318(.A0(n7489), .A1(n6159), .B0(n7534), .Y(P2_U3291));
  OAI22X1 g6319(.A0(n7488), .A1(n6163), .B0(n6223), .B1(n7520), .Y(n7536));
  OAI22X1 g6320(.A0(n7522), .A1(n6168), .B0(n6206), .B1(n7523), .Y(n7537));
  NAND4X1 g6321(.A(n6214), .B(n5924), .C(n5855), .D(n7488), .Y(n7538));
  OAI21X1 g6322(.A0(n7525), .A1(n6215), .B0(n7538), .Y(n7539));
  NOR3X1  g6323(.A(n7539), .B(n7537), .C(n7536), .Y(n7540));
  OAI21X1 g6324(.A0(n7489), .A1(n6211), .B0(n7540), .Y(P2_U3290));
  NOR3X1  g6325(.A(n6262), .B(n6258), .C(n6247), .Y(n7542));
  INVX1   g6326(.A(n6221), .Y(n7543));
  AOI22X1 g6327(.A0(n7496), .A1(n7543), .B0(n6265), .B1(n7498), .Y(n7544));
  OAI21X1 g6328(.A0(n7525), .A1(n6264), .B0(n7544), .Y(n7545));
  AOI22X1 g6329(.A0(n7489), .A1(P2_REG2_REG_7__SCAN_IN), .B0(n6292), .B1(n7490), .Y(n7546));
  OAI21X1 g6330(.A0(n7523), .A1(n6246), .B0(n7546), .Y(n7547));
  NOR2X1  g6331(.A(n7547), .B(n7545), .Y(n7548));
  OAI21X1 g6332(.A0(n7489), .A1(n7542), .B0(n7548), .Y(P2_U3289));
  NOR3X1  g6333(.A(n6312), .B(n6309), .C(n6296), .Y(n7550));
  NOR2X1  g6334(.A(n7523), .B(n6295), .Y(n7551));
  AOI22X1 g6335(.A0(n7489), .A1(P2_REG2_REG_8__SCAN_IN), .B0(n6354), .B1(n7490), .Y(n7552));
  INVX1   g6336(.A(n7494), .Y(n7553));
  NAND3X1 g6337(.A(n7553), .B(n7488), .C(n6289), .Y(n7554));
  INVX1   g6338(.A(n6273), .Y(n7555));
  AOI22X1 g6339(.A0(n7496), .A1(n7555), .B0(n6317), .B1(n7498), .Y(n7556));
  NAND3X1 g6340(.A(n7556), .B(n7554), .C(n7552), .Y(n7557));
  NOR2X1  g6341(.A(n7557), .B(n7551), .Y(n7558));
  OAI21X1 g6342(.A0(n7489), .A1(n7550), .B0(n7558), .Y(P2_U3288));
  NOR3X1  g6343(.A(n6362), .B(n6359), .C(n6349), .Y(n7560));
  AOI22X1 g6344(.A0(n7489), .A1(P2_REG2_REG_9__SCAN_IN), .B0(n6386), .B1(n7490), .Y(n7561));
  NAND3X1 g6345(.A(n7553), .B(n7488), .C(n6338), .Y(n7562));
  INVX1   g6346(.A(n6325), .Y(n7563));
  AOI22X1 g6347(.A0(n7496), .A1(n7563), .B0(n6365), .B1(n7498), .Y(n7564));
  NAND3X1 g6348(.A(n7564), .B(n7562), .C(n7561), .Y(n7565));
  AOI21X1 g6349(.A0(n7499), .A1(n6360), .B0(n7565), .Y(n7566));
  OAI21X1 g6350(.A0(n7489), .A1(n7560), .B0(n7566), .Y(P2_U3287));
  NOR3X1  g6351(.A(n6414), .B(n6410), .C(n6401), .Y(n7568));
  NOR2X1  g6352(.A(n7523), .B(n6400), .Y(n7569));
  AOI22X1 g6353(.A0(n7489), .A1(P2_REG2_REG_10__SCAN_IN), .B0(n6391), .B1(n7495), .Y(n7570));
  NAND3X1 g6354(.A(n7481), .B(n6384), .C(n5743), .Y(n7571));
  AOI22X1 g6355(.A0(n7490), .A1(n6451), .B0(n6417), .B1(n7498), .Y(n7572));
  NAND3X1 g6356(.A(n7572), .B(n7571), .C(n7570), .Y(n7573));
  NOR2X1  g6357(.A(n7573), .B(n7569), .Y(n7574));
  OAI21X1 g6358(.A0(n7489), .A1(n7568), .B0(n7574), .Y(P2_U3286));
  OAI21X1 g6359(.A0(n6483), .A1(n6481), .B0(n7488), .Y(n7576));
  NOR2X1  g6360(.A(n7523), .B(n6470), .Y(n7577));
  AOI22X1 g6361(.A0(n7489), .A1(P2_REG2_REG_11__SCAN_IN), .B0(n6493), .B1(n7490), .Y(n7578));
  NAND3X1 g6362(.A(n7553), .B(n7488), .C(n6443), .Y(n7579));
  INVX1   g6363(.A(n6428), .Y(n7580));
  AOI22X1 g6364(.A0(n7496), .A1(n7580), .B0(n6485), .B1(n7498), .Y(n7581));
  NAND3X1 g6365(.A(n7581), .B(n7579), .C(n7578), .Y(n7582));
  NOR2X1  g6366(.A(n7582), .B(n7577), .Y(n7583));
  NAND2X1 g6367(.A(n7583), .B(n7576), .Y(P2_U3285));
  NOR3X1  g6368(.A(n6535), .B(n6527), .C(n6516), .Y(n7585));
  NOR2X1  g6369(.A(n7523), .B(n6525), .Y(n7586));
  INVX1   g6370(.A(n6537), .Y(n7587));
  NOR4X1  g6371(.A(n7587), .B(n5925), .C(n5856), .D(n7489), .Y(n7588));
  INVX1   g6372(.A(P2_REG2_REG_12__SCAN_IN), .Y(n7589));
  OAI22X1 g6373(.A0(n7488), .A1(n7589), .B0(n6528), .B1(n7525), .Y(n7590));
  OAI22X1 g6374(.A0(n7520), .A1(n6546), .B0(n6490), .B1(n7522), .Y(n7591));
  NOR4X1  g6375(.A(n7590), .B(n7588), .C(n7586), .D(n7591), .Y(n7592));
  OAI21X1 g6376(.A0(n7489), .A1(n7585), .B0(n7592), .Y(P2_U3284));
  NOR3X1  g6377(.A(n6585), .B(n6581), .C(n6573), .Y(n7594));
  NOR2X1  g6378(.A(n7523), .B(n6569), .Y(n7595));
  NAND4X1 g6379(.A(n6587), .B(n5924), .C(n5855), .D(n7488), .Y(n7596));
  AOI22X1 g6380(.A0(n7489), .A1(P2_REG2_REG_13__SCAN_IN), .B0(n6558), .B1(n7495), .Y(n7597));
  INVX1   g6381(.A(n6542), .Y(n7598));
  AOI22X1 g6382(.A0(n7490), .A1(n6660), .B0(n7598), .B1(n7496), .Y(n7599));
  NAND3X1 g6383(.A(n7599), .B(n7597), .C(n7596), .Y(n7600));
  NOR2X1  g6384(.A(n7600), .B(n7595), .Y(n7601));
  OAI21X1 g6385(.A0(n7489), .A1(n7594), .B0(n7601), .Y(P2_U3283));
  NOR3X1  g6386(.A(n6632), .B(n6629), .C(n6628), .Y(n7603));
  NOR2X1  g6387(.A(n7523), .B(n6622), .Y(n7604));
  NOR4X1  g6388(.A(n6637), .B(n5925), .C(n5856), .D(n7489), .Y(n7605));
  INVX1   g6389(.A(P2_REG2_REG_14__SCAN_IN), .Y(n7606));
  OAI22X1 g6390(.A0(n7488), .A1(n7606), .B0(n6634), .B1(n7525), .Y(n7607));
  OAI22X1 g6391(.A0(n7520), .A1(n6646), .B0(n6595), .B1(n7522), .Y(n7608));
  NOR4X1  g6392(.A(n7607), .B(n7605), .C(n7604), .D(n7608), .Y(n7609));
  OAI21X1 g6393(.A0(n7489), .A1(n7603), .B0(n7609), .Y(P2_U3282));
  NOR3X1  g6394(.A(n6677), .B(n6676), .C(n6675), .Y(n7611));
  NOR2X1  g6395(.A(n7523), .B(n6669), .Y(n7612));
  NAND4X1 g6396(.A(n6679), .B(n5924), .C(n5855), .D(n7488), .Y(n7613));
  AOI22X1 g6397(.A0(n7489), .A1(P2_REG2_REG_15__SCAN_IN), .B0(n6657), .B1(n7495), .Y(n7614));
  AOI22X1 g6398(.A0(n7490), .A1(n6689), .B0(n6643), .B1(n7496), .Y(n7615));
  NAND3X1 g6399(.A(n7615), .B(n7614), .C(n7613), .Y(n7616));
  NOR2X1  g6400(.A(n7616), .B(n7612), .Y(n7617));
  OAI21X1 g6401(.A0(n7489), .A1(n7611), .B0(n7617), .Y(P2_U3281));
  NOR3X1  g6402(.A(n6727), .B(n6726), .C(n6725), .Y(n7619));
  NOR2X1  g6403(.A(n7523), .B(n6718), .Y(n7620));
  INVX1   g6404(.A(n6729), .Y(n7621));
  NOR4X1  g6405(.A(n7621), .B(n5925), .C(n5856), .D(n7489), .Y(n7622));
  INVX1   g6406(.A(P2_REG2_REG_16__SCAN_IN), .Y(n7623));
  OAI22X1 g6407(.A0(n7488), .A1(n7623), .B0(n6731), .B1(n7525), .Y(n7624));
  OAI22X1 g6408(.A0(n7520), .A1(n6740), .B0(n6686), .B1(n7522), .Y(n7625));
  NOR4X1  g6409(.A(n7624), .B(n7622), .C(n7620), .D(n7625), .Y(n7626));
  OAI21X1 g6410(.A0(n7489), .A1(n7619), .B0(n7626), .Y(P2_U3280));
  NOR3X1  g6411(.A(n6788), .B(n6784), .C(n6771), .Y(n7628));
  NOR2X1  g6412(.A(n7523), .B(n6766), .Y(n7629));
  NAND4X1 g6413(.A(n6790), .B(n5924), .C(n5855), .D(n7488), .Y(n7630));
  NAND3X1 g6414(.A(n7553), .B(n7488), .C(n6753), .Y(n7631));
  INVX1   g6415(.A(P2_REG2_REG_17__SCAN_IN), .Y(n7632));
  OAI22X1 g6416(.A0(n7488), .A1(n7632), .B0(n6734), .B1(n7522), .Y(n7633));
  AOI21X1 g6417(.A0(n7490), .A1(n6818), .B0(n7633), .Y(n7634));
  NAND3X1 g6418(.A(n7634), .B(n7631), .C(n7630), .Y(n7635));
  NOR2X1  g6419(.A(n7635), .B(n7629), .Y(n7636));
  OAI21X1 g6420(.A0(n7489), .A1(n7628), .B0(n7636), .Y(P2_U3279));
  NOR3X1  g6421(.A(n6833), .B(n6826), .C(n6822), .Y(n7638));
  NOR2X1  g6422(.A(n7523), .B(n6821), .Y(n7639));
  NAND4X1 g6423(.A(n6835), .B(n5924), .C(n5855), .D(n7488), .Y(n7640));
  NAND3X1 g6424(.A(n7553), .B(n7488), .C(n6815), .Y(n7641));
  NAND3X1 g6425(.A(n7488), .B(n6872), .C(n5915), .Y(n7642));
  AOI22X1 g6426(.A0(n7489), .A1(P2_REG2_REG_18__SCAN_IN), .B0(n6792), .B1(n7496), .Y(n7643));
  NAND4X1 g6427(.A(n7642), .B(n7641), .C(n7640), .D(n7643), .Y(n7644));
  NOR2X1  g6428(.A(n7644), .B(n7639), .Y(n7645));
  OAI21X1 g6429(.A0(n7489), .A1(n7638), .B0(n7645), .Y(P2_U3278));
  NOR3X1  g6430(.A(n6882), .B(n6881), .C(n6880), .Y(n7647));
  NAND4X1 g6431(.A(n6886), .B(n5924), .C(n5855), .D(n7488), .Y(n7648));
  NAND3X1 g6432(.A(n7553), .B(n7488), .C(n6854), .Y(n7649));
  NAND3X1 g6433(.A(n7488), .B(n6914), .C(n5915), .Y(n7650));
  INVX1   g6434(.A(n6839), .Y(n7651));
  AOI22X1 g6435(.A0(n7489), .A1(P2_REG2_REG_19__SCAN_IN), .B0(n7651), .B1(n7496), .Y(n7652));
  NAND4X1 g6436(.A(n7650), .B(n7649), .C(n7648), .D(n7652), .Y(n7653));
  AOI21X1 g6437(.A0(n7499), .A1(n6874), .B0(n7653), .Y(n7654));
  OAI21X1 g6438(.A0(n7489), .A1(n7647), .B0(n7654), .Y(P2_U3277));
  NAND2X1 g6439(.A(n7488), .B(n6936), .Y(n7656));
  NAND3X1 g6440(.A(n7499), .B(n6924), .C(n6919), .Y(n7657));
  NAND2X1 g6441(.A(n7498), .B(n6938), .Y(n7658));
  INVX1   g6442(.A(n6888), .Y(n7659));
  AOI22X1 g6443(.A0(n7489), .A1(P2_REG2_REG_20__SCAN_IN), .B0(n7659), .B1(n7496), .Y(n7660));
  OAI21X1 g6444(.A0(n7520), .A1(n6947), .B0(n7660), .Y(n7661));
  AOI21X1 g6445(.A0(n7495), .A1(n6901), .B0(n7661), .Y(n7662));
  NAND4X1 g6446(.A(n7658), .B(n7657), .C(n7656), .D(n7662), .Y(P2_U3276));
  NAND2X1 g6447(.A(n7488), .B(n6981), .Y(n7664));
  INVX1   g6448(.A(n6972), .Y(n7665));
  NAND2X1 g6449(.A(n7499), .B(n7665), .Y(n7666));
  NAND2X1 g6450(.A(n7498), .B(n6983), .Y(n7667));
  INVX1   g6451(.A(n6941), .Y(n7668));
  AOI22X1 g6452(.A0(n7489), .A1(P2_REG2_REG_21__SCAN_IN), .B0(n7668), .B1(n7496), .Y(n7669));
  OAI21X1 g6453(.A0(n7520), .A1(n6995), .B0(n7669), .Y(n7670));
  AOI21X1 g6454(.A0(n7495), .A1(n6954), .B0(n7670), .Y(n7671));
  NAND4X1 g6455(.A(n7667), .B(n7666), .C(n7664), .D(n7671), .Y(P2_U3275));
  NOR3X1  g6456(.A(n7026), .B(n7025), .C(n7024), .Y(n7673));
  NOR2X1  g6457(.A(n7523), .B(n7017), .Y(n7674));
  NAND2X1 g6458(.A(n7498), .B(n7029), .Y(n7675));
  NAND2X1 g6459(.A(n7495), .B(n7002), .Y(n7676));
  NAND3X1 g6460(.A(n7488), .B(n7053), .C(n5915), .Y(n7677));
  INVX1   g6461(.A(n6988), .Y(n7678));
  AOI22X1 g6462(.A0(n7489), .A1(P2_REG2_REG_22__SCAN_IN), .B0(n7678), .B1(n7496), .Y(n7679));
  NAND4X1 g6463(.A(n7677), .B(n7676), .C(n7675), .D(n7679), .Y(n7680));
  NOR2X1  g6464(.A(n7680), .B(n7674), .Y(n7681));
  OAI21X1 g6465(.A0(n7489), .A1(n7673), .B0(n7681), .Y(P2_U3274));
  NAND2X1 g6466(.A(n7488), .B(n7075), .Y(n7683));
  INVX1   g6467(.A(n7066), .Y(n7684));
  NAND2X1 g6468(.A(n7499), .B(n7684), .Y(n7685));
  NAND2X1 g6469(.A(n7498), .B(n7077), .Y(n7686));
  AOI22X1 g6470(.A0(n7489), .A1(P2_REG2_REG_23__SCAN_IN), .B0(n7033), .B1(n7496), .Y(n7687));
  OAI21X1 g6471(.A0(n7520), .A1(n7083), .B0(n7687), .Y(n7688));
  AOI21X1 g6472(.A0(n7495), .A1(n7049), .B0(n7688), .Y(n7689));
  NAND4X1 g6473(.A(n7686), .B(n7685), .C(n7683), .D(n7689), .Y(P2_U3273));
  NOR3X1  g6474(.A(n7116), .B(n7115), .C(n7114), .Y(n7691));
  NAND2X1 g6475(.A(n7498), .B(n7119), .Y(n7692));
  AOI22X1 g6476(.A0(n7489), .A1(P2_REG2_REG_24__SCAN_IN), .B0(n7079), .B1(n7496), .Y(n7693));
  OAI21X1 g6477(.A0(n7520), .A1(n7127), .B0(n7693), .Y(n7694));
  AOI21X1 g6478(.A0(n7495), .A1(n7165), .B0(n7694), .Y(n7695));
  NAND2X1 g6479(.A(n7695), .B(n7692), .Y(n7696));
  AOI21X1 g6480(.A0(n7499), .A1(n7108), .B0(n7696), .Y(n7697));
  OAI21X1 g6481(.A0(n7489), .A1(n7691), .B0(n7697), .Y(P2_U3272));
  OAI21X1 g6482(.A0(n7163), .A1(n7160), .B0(n7488), .Y(n7699));
  NAND2X1 g6483(.A(n7499), .B(n7154), .Y(n7700));
  NAND2X1 g6484(.A(n7498), .B(n7168), .Y(n7701));
  AOI22X1 g6485(.A0(n7489), .A1(P2_REG2_REG_25__SCAN_IN), .B0(n7122), .B1(n7496), .Y(n7702));
  OAI21X1 g6486(.A0(n7520), .A1(n7176), .B0(n7702), .Y(n7703));
  AOI21X1 g6487(.A0(n7495), .A1(n7134), .B0(n7703), .Y(n7704));
  NAND4X1 g6488(.A(n7701), .B(n7700), .C(n7699), .D(n7704), .Y(P2_U3271));
  NOR3X1  g6489(.A(n7215), .B(n7214), .C(n7213), .Y(n7706));
  NAND2X1 g6490(.A(n7498), .B(n7220), .Y(n7707));
  AOI22X1 g6491(.A0(n7489), .A1(P2_REG2_REG_26__SCAN_IN), .B0(n7171), .B1(n7496), .Y(n7708));
  OAI21X1 g6492(.A0(n7520), .A1(n7228), .B0(n7708), .Y(n7709));
  AOI21X1 g6493(.A0(n7495), .A1(n7184), .B0(n7709), .Y(n7710));
  NAND2X1 g6494(.A(n7710), .B(n7707), .Y(n7711));
  AOI21X1 g6495(.A0(n7499), .A1(n7206), .B0(n7711), .Y(n7712));
  OAI21X1 g6496(.A0(n7489), .A1(n7706), .B0(n7712), .Y(P2_U3270));
  NOR3X1  g6497(.A(n7269), .B(n7268), .C(n7266), .Y(n7714));
  NAND2X1 g6498(.A(n7498), .B(n7273), .Y(n7715));
  AOI22X1 g6499(.A0(n7489), .A1(P2_REG2_REG_27__SCAN_IN), .B0(n7223), .B1(n7496), .Y(n7716));
  OAI21X1 g6500(.A0(n7520), .A1(n7283), .B0(n7716), .Y(n7717));
  AOI21X1 g6501(.A0(n7495), .A1(n7272), .B0(n7717), .Y(n7718));
  NAND2X1 g6502(.A(n7718), .B(n7715), .Y(n7719));
  AOI21X1 g6503(.A0(n7499), .A1(n7256), .B0(n7719), .Y(n7720));
  OAI21X1 g6504(.A0(n7489), .A1(n7714), .B0(n7720), .Y(P2_U3269));
  NOR4X1  g6505(.A(n7313), .B(n7306), .C(n7302), .D(n7314), .Y(n7722));
  NOR2X1  g6506(.A(n7523), .B(n7301), .Y(n7723));
  INVX1   g6507(.A(n7498), .Y(n7724));
  AOI22X1 g6508(.A0(n7489), .A1(P2_REG2_REG_28__SCAN_IN), .B0(n7278), .B1(n7496), .Y(n7725));
  OAI21X1 g6509(.A0(n7520), .A1(n7325), .B0(n7725), .Y(n7726));
  AOI21X1 g6510(.A0(n7495), .A1(n7290), .B0(n7726), .Y(n7727));
  OAI21X1 g6511(.A0(n7724), .A1(n7319), .B0(n7727), .Y(n7728));
  NOR2X1  g6512(.A(n7728), .B(n7723), .Y(n7729));
  OAI21X1 g6513(.A0(n7489), .A1(n7722), .B0(n7729), .Y(P2_U3268));
  NOR3X1  g6514(.A(n7383), .B(n7378), .C(n7365), .Y(n7731));
  XOR2X1  g6515(.A(n7381), .B(n7334), .Y(n7732));
  NAND2X1 g6516(.A(n7498), .B(n7387), .Y(n7733));
  NAND2X1 g6517(.A(n7495), .B(n7333), .Y(n7734));
  NOR4X1  g6518(.A(n7221), .B(n7274), .C(n7275), .D(n7522), .Y(n7735));
  AOI21X1 g6519(.A0(n7489), .A1(P2_REG2_REG_29__SCAN_IN), .B0(n7735), .Y(n7736));
  NAND3X1 g6520(.A(n7736), .B(n7734), .C(n7733), .Y(n7737));
  AOI21X1 g6521(.A0(n7499), .A1(n7732), .B0(n7737), .Y(n7738));
  OAI21X1 g6522(.A0(n7489), .A1(n7731), .B0(n7738), .Y(P2_U3267));
  NAND2X1 g6523(.A(n7498), .B(n7395), .Y(n7740));
  NAND2X1 g6524(.A(n7495), .B(n7407), .Y(n7741));
  NAND2X1 g6525(.A(n7488), .B(n7400), .Y(n7742));
  NAND2X1 g6526(.A(n7489), .B(P2_REG2_REG_30__SCAN_IN), .Y(n7743));
  NAND4X1 g6527(.A(n7742), .B(n7741), .C(n7740), .D(n7743), .Y(P2_U3266));
  NAND2X1 g6528(.A(n7498), .B(n7410), .Y(n7745));
  AOI21X1 g6529(.A0(n5727), .A1(n5726), .B0(n5867), .Y(n7746));
  NAND2X1 g6530(.A(n7495), .B(n7746), .Y(n7747));
  NAND2X1 g6531(.A(n7489), .B(P2_REG2_REG_31__SCAN_IN), .Y(n7748));
  NAND4X1 g6532(.A(n7747), .B(n7745), .C(n7742), .D(n7748), .Y(P2_U3265));
  NOR4X1  g6533(.A(n5739), .B(n5737), .C(n5735), .D(n5741), .Y(n7750));
  AOI21X1 g6534(.A0(n5871), .A1(n5869), .B0(n5734), .Y(n7751));
  AOI22X1 g6535(.A0(n5869), .A1(n5871), .B0(n5847), .B1(n5843), .Y(n7752));
  NOR4X1  g6536(.A(n7751), .B(n7750), .C(P2_U3152), .D(n7752), .Y(n7753));
  NOR4X1  g6537(.A(n5742), .B(n5735), .C(P2_U3152), .D(n7753), .Y(n7754));
  NOR2X1  g6538(.A(n5871), .B(n5869), .Y(n7755));
  INVX1   g6539(.A(n7755), .Y(n7756));
  INVX1   g6540(.A(P2_REG2_REG_18__SCAN_IN), .Y(n7757));
  AOI22X1 g6541(.A0(n6701), .A1(n7623), .B0(n7632), .B1(n6750), .Y(n7758));
  NOR2X1  g6542(.A(n6655), .B(P2_REG2_REG_15__SCAN_IN), .Y(n7759));
  INVX1   g6543(.A(P2_REG2_REG_13__SCAN_IN), .Y(n7760));
  NAND2X1 g6544(.A(n6555), .B(n7760), .Y(n7761));
  NOR2X1  g6545(.A(n6440), .B(n6420), .Y(n7762));
  INVX1   g6546(.A(n7762), .Y(n7763));
  AOI22X1 g6547(.A0(n6503), .A1(n7589), .B0(n7760), .B1(n6555), .Y(n7764));
  INVX1   g6548(.A(n7764), .Y(n7765));
  NOR2X1  g6549(.A(n6503), .B(n7589), .Y(n7766));
  AOI21X1 g6550(.A0(n6556), .A1(P2_REG2_REG_13__SCAN_IN), .B0(n7766), .Y(n7767));
  OAI21X1 g6551(.A0(n7765), .A1(n7763), .B0(n7767), .Y(n7768));
  NOR2X1  g6552(.A(n6286), .B(n6266), .Y(n7769));
  AOI22X1 g6553(.A0(n6335), .A1(n6318), .B0(n6366), .B1(n6388), .Y(n7770));
  NAND2X1 g6554(.A(n6336), .B(P2_REG2_REG_9__SCAN_IN), .Y(n7771));
  OAI21X1 g6555(.A0(n6388), .A1(n6366), .B0(n7771), .Y(n7772));
  AOI21X1 g6556(.A0(n7770), .A1(n7769), .B0(n7772), .Y(n7773));
  AOI21X1 g6557(.A0(n6388), .A1(n6366), .B0(n7773), .Y(n7774));
  AOI22X1 g6558(.A0(n6182), .A1(n6163), .B0(n6216), .B1(n6236), .Y(n7775));
  AOI22X1 g6559(.A0(n6074), .A1(n6087), .B0(n6114), .B1(n6130), .Y(n7776));
  OAI22X1 g6560(.A0(n5988), .A1(P2_REG2_REG_2__SCAN_IN), .B0(P2_REG2_REG_3__SCAN_IN), .B1(n6031), .Y(n7777));
  NOR2X1  g6561(.A(n5477), .B(n5879), .Y(n7778));
  INVX1   g6562(.A(n7778), .Y(n7779));
  AOI21X1 g6563(.A0(n5936), .A1(n5949), .B0(n7779), .Y(n7780));
  NOR2X1  g6564(.A(n5936), .B(n5949), .Y(n7781));
  NOR2X1  g6565(.A(n7781), .B(n7780), .Y(n7782));
  NOR2X1  g6566(.A(n6030), .B(n6010), .Y(n7783));
  NOR2X1  g6567(.A(n6031), .B(P2_REG2_REG_3__SCAN_IN), .Y(n7784));
  NOR3X1  g6568(.A(n7784), .B(n5987), .C(n5969), .Y(n7785));
  NOR2X1  g6569(.A(n7785), .B(n7783), .Y(n7786));
  OAI21X1 g6570(.A0(n7782), .A1(n7777), .B0(n7786), .Y(n7787));
  NAND2X1 g6571(.A(n7787), .B(n7776), .Y(n7788));
  INVX1   g6572(.A(n6130), .Y(n7789));
  NOR3X1  g6573(.A(n6074), .B(n6114), .C(n6087), .Y(n7790));
  OAI21X1 g6574(.A0(n6074), .A1(n6087), .B0(n6114), .Y(n7791));
  AOI21X1 g6575(.A0(n7791), .A1(n7789), .B0(n7790), .Y(n7792));
  NAND2X1 g6576(.A(n7792), .B(n7788), .Y(n7793));
  NAND2X1 g6577(.A(n7793), .B(n7775), .Y(n7794));
  NOR3X1  g6578(.A(n6182), .B(n6216), .C(n6163), .Y(n7795));
  OAI21X1 g6579(.A0(n6182), .A1(n6163), .B0(n6216), .Y(n7796));
  AOI21X1 g6580(.A0(n7796), .A1(n6237), .B0(n7795), .Y(n7797));
  NAND2X1 g6581(.A(n7797), .B(n7794), .Y(n7798));
  NOR2X1  g6582(.A(n6287), .B(P2_REG2_REG_8__SCAN_IN), .Y(n7799));
  INVX1   g6583(.A(n7799), .Y(n7800));
  NAND3X1 g6584(.A(n7800), .B(n7798), .C(n7770), .Y(n7801));
  INVX1   g6585(.A(n7801), .Y(n7802));
  NOR2X1  g6586(.A(n7802), .B(n7774), .Y(n7803));
  INVX1   g6587(.A(n7803), .Y(n7804));
  AOI21X1 g6588(.A0(n6440), .A1(n6420), .B0(n7765), .Y(n7805));
  AOI22X1 g6589(.A0(n7804), .A1(n7805), .B0(n7768), .B1(n7761), .Y(n7806));
  AOI21X1 g6590(.A0(n6606), .A1(n7606), .B0(n7806), .Y(n7807));
  AOI21X1 g6591(.A0(n6607), .A1(P2_REG2_REG_14__SCAN_IN), .B0(n7807), .Y(n7808));
  NOR2X1  g6592(.A(n7808), .B(n7759), .Y(n7809));
  AOI21X1 g6593(.A0(n6655), .A1(P2_REG2_REG_15__SCAN_IN), .B0(n7809), .Y(n7810));
  INVX1   g6594(.A(n7810), .Y(n7811));
  NOR2X1  g6595(.A(n6701), .B(n7623), .Y(n7812));
  NAND2X1 g6596(.A(n7812), .B(P2_REG2_REG_17__SCAN_IN), .Y(n7813));
  NOR2X1  g6597(.A(n7812), .B(P2_REG2_REG_17__SCAN_IN), .Y(n7814));
  OAI21X1 g6598(.A0(n7814), .A1(n6750), .B0(n7813), .Y(n7815));
  AOI21X1 g6599(.A0(n7811), .A1(n7758), .B0(n7815), .Y(n7816));
  OAI21X1 g6600(.A0(n6812), .A1(n7757), .B0(n7816), .Y(n7817));
  XOR2X1  g6601(.A(n5855), .B(P2_REG2_REG_19__SCAN_IN), .Y(n7818));
  AOI21X1 g6602(.A0(n6812), .A1(n7757), .B0(n7818), .Y(n7819));
  NAND2X1 g6603(.A(n7819), .B(n7817), .Y(n7820));
  AOI21X1 g6604(.A0(n6812), .A1(n7757), .B0(n7816), .Y(n7821));
  OAI21X1 g6605(.A0(n6812), .A1(n7757), .B0(n7818), .Y(n7822));
  OAI21X1 g6606(.A0(n7822), .A1(n7821), .B0(n7820), .Y(n7823));
  OAI22X1 g6607(.A0(n7756), .A1(n7823), .B0(n5866), .B1(n5855), .Y(n7824));
  INVX1   g6608(.A(P2_REG1_REG_18__SCAN_IN), .Y(n7825));
  INVX1   g6609(.A(P2_REG1_REG_16__SCAN_IN), .Y(n7826));
  INVX1   g6610(.A(P2_REG1_REG_17__SCAN_IN), .Y(n7827));
  AOI22X1 g6611(.A0(n6701), .A1(n7826), .B0(n7827), .B1(n6750), .Y(n7828));
  INVX1   g6612(.A(P2_REG1_REG_15__SCAN_IN), .Y(n7829));
  NOR2X1  g6613(.A(n6606), .B(n6590), .Y(n7830));
  NAND2X1 g6614(.A(n6606), .B(n6590), .Y(n7831));
  NOR2X1  g6615(.A(n6440), .B(n6423), .Y(n7832));
  INVX1   g6616(.A(n7832), .Y(n7833));
  INVX1   g6617(.A(P2_REG1_REG_12__SCAN_IN), .Y(n7834));
  AOI22X1 g6618(.A0(n6503), .A1(n7834), .B0(n6539), .B1(n6555), .Y(n7835));
  INVX1   g6619(.A(n7835), .Y(n7836));
  NOR2X1  g6620(.A(n6503), .B(n7834), .Y(n7837));
  AOI21X1 g6621(.A0(n6556), .A1(P2_REG1_REG_13__SCAN_IN), .B0(n7837), .Y(n7838));
  OAI21X1 g6622(.A0(n7836), .A1(n7833), .B0(n7838), .Y(n7839));
  OAI21X1 g6623(.A0(n6556), .A1(P2_REG1_REG_13__SCAN_IN), .B0(n7839), .Y(n7840));
  NOR2X1  g6624(.A(n6286), .B(n6269), .Y(n7841));
  AOI22X1 g6625(.A0(n6335), .A1(n6321), .B0(n6369), .B1(n6388), .Y(n7842));
  NAND2X1 g6626(.A(n6336), .B(P2_REG1_REG_9__SCAN_IN), .Y(n7843));
  OAI21X1 g6627(.A0(n6388), .A1(n6369), .B0(n7843), .Y(n7844));
  AOI21X1 g6628(.A0(n7842), .A1(n7841), .B0(n7844), .Y(n7845));
  AOI21X1 g6629(.A0(n6388), .A1(n6369), .B0(n7845), .Y(n7846));
  INVX1   g6630(.A(P2_REG1_REG_6__SCAN_IN), .Y(n7847));
  AOI22X1 g6631(.A0(n6182), .A1(n7847), .B0(n6219), .B1(n6236), .Y(n7848));
  AOI22X1 g6632(.A0(n6074), .A1(n6090), .B0(n6117), .B1(n6130), .Y(n7849));
  AOI22X1 g6633(.A0(n5987), .A1(n5968), .B0(n6013), .B1(n6030), .Y(n7850));
  INVX1   g6634(.A(n7850), .Y(n7851));
  NOR2X1  g6635(.A(n5477), .B(n5878), .Y(n7852));
  INVX1   g6636(.A(n7852), .Y(n7853));
  AOI21X1 g6637(.A0(n5936), .A1(n5948), .B0(n7853), .Y(n7854));
  NOR2X1  g6638(.A(n5936), .B(n5948), .Y(n7855));
  NOR2X1  g6639(.A(n7855), .B(n7854), .Y(n7856));
  NOR2X1  g6640(.A(n6030), .B(n6013), .Y(n7857));
  NOR2X1  g6641(.A(n6031), .B(P2_REG1_REG_3__SCAN_IN), .Y(n7858));
  NOR3X1  g6642(.A(n7858), .B(n5987), .C(n5968), .Y(n7859));
  NOR2X1  g6643(.A(n7859), .B(n7857), .Y(n7860));
  OAI21X1 g6644(.A0(n7856), .A1(n7851), .B0(n7860), .Y(n7861));
  NAND2X1 g6645(.A(n7861), .B(n7849), .Y(n7862));
  NOR3X1  g6646(.A(n6074), .B(n6117), .C(n6090), .Y(n7863));
  OAI21X1 g6647(.A0(n6074), .A1(n6090), .B0(n6117), .Y(n7864));
  AOI21X1 g6648(.A0(n7864), .A1(n7789), .B0(n7863), .Y(n7865));
  NAND2X1 g6649(.A(n7865), .B(n7862), .Y(n7866));
  NAND2X1 g6650(.A(n7866), .B(n7848), .Y(n7867));
  NOR3X1  g6651(.A(n6182), .B(n6219), .C(n7847), .Y(n7868));
  OAI21X1 g6652(.A0(n6182), .A1(n7847), .B0(n6219), .Y(n7869));
  AOI21X1 g6653(.A0(n7869), .A1(n6237), .B0(n7868), .Y(n7870));
  NAND2X1 g6654(.A(n7870), .B(n7867), .Y(n7871));
  NOR2X1  g6655(.A(n6287), .B(P2_REG1_REG_8__SCAN_IN), .Y(n7872));
  INVX1   g6656(.A(n7872), .Y(n7873));
  NAND3X1 g6657(.A(n7873), .B(n7871), .C(n7842), .Y(n7874));
  INVX1   g6658(.A(n7874), .Y(n7875));
  NOR2X1  g6659(.A(n7875), .B(n7846), .Y(n7876));
  OAI21X1 g6660(.A0(n6441), .A1(P2_REG1_REG_11__SCAN_IN), .B0(n7835), .Y(n7877));
  OAI21X1 g6661(.A0(n7877), .A1(n7876), .B0(n7840), .Y(n7878));
  AOI21X1 g6662(.A0(n7878), .A1(n7831), .B0(n7830), .Y(n7879));
  AOI21X1 g6663(.A0(n6654), .A1(n7829), .B0(n7879), .Y(n7880));
  AOI21X1 g6664(.A0(n6655), .A1(P2_REG1_REG_15__SCAN_IN), .B0(n7880), .Y(n7881));
  INVX1   g6665(.A(n7881), .Y(n7882));
  NOR3X1  g6666(.A(n6701), .B(n7827), .C(n7826), .Y(n7883));
  OAI21X1 g6667(.A0(n6701), .A1(n7826), .B0(n7827), .Y(n7884));
  AOI21X1 g6668(.A0(n7884), .A1(n6751), .B0(n7883), .Y(n7885));
  INVX1   g6669(.A(n7885), .Y(n7886));
  AOI21X1 g6670(.A0(n7882), .A1(n7828), .B0(n7886), .Y(n7887));
  OAI21X1 g6671(.A0(n6812), .A1(n7825), .B0(n7887), .Y(n7888));
  XOR2X1  g6672(.A(n5855), .B(P2_REG1_REG_19__SCAN_IN), .Y(n7889));
  AOI21X1 g6673(.A0(n6812), .A1(n7825), .B0(n7889), .Y(n7890));
  NAND2X1 g6674(.A(n7890), .B(n7888), .Y(n7891));
  AOI21X1 g6675(.A0(n6812), .A1(n7825), .B0(n7887), .Y(n7892));
  OAI21X1 g6676(.A0(n6812), .A1(n7825), .B0(n7889), .Y(n7893));
  OAI21X1 g6677(.A0(n7893), .A1(n7892), .B0(n7891), .Y(n7894));
  NOR2X1  g6678(.A(n7894), .B(n5864), .Y(n7895));
  OAI21X1 g6679(.A0(n7895), .A1(n7824), .B0(n7754), .Y(n7896));
  NAND2X1 g6680(.A(n7750), .B(P2_STATE_REG_SCAN_IN), .Y(n7897));
  INVX1   g6681(.A(n7897), .Y(P2_U3966));
  NOR2X1  g6682(.A(n5871), .B(n5864), .Y(n7899));
  INVX1   g6683(.A(n7899), .Y(n7900));
  NOR2X1  g6684(.A(n7900), .B(n7894), .Y(n7901));
  OAI21X1 g6685(.A0(n7901), .A1(n7824), .B0(P2_U3966), .Y(n7902));
  NOR4X1  g6686(.A(n7753), .B(n5734), .C(P2_U3152), .D(n7756), .Y(n7903));
  INVX1   g6687(.A(n7903), .Y(n7904));
  NOR2X1  g6688(.A(n7904), .B(n7823), .Y(n7905));
  NOR4X1  g6689(.A(n5864), .B(n5734), .C(P2_U3152), .D(n7753), .Y(n7906));
  INVX1   g6690(.A(n7906), .Y(n7907));
  NOR2X1  g6691(.A(n7907), .B(n7894), .Y(n7908));
  NOR4X1  g6692(.A(n5866), .B(n5734), .C(P2_U3152), .D(n7753), .Y(n7909));
  INVX1   g6693(.A(n7909), .Y(n7910));
  AOI22X1 g6694(.A0(P2_ADDR_REG_19__SCAN_IN), .A1(n7753), .B0(P2_REG3_REG_19__SCAN_IN), .B1(P2_U3152), .Y(n7911));
  OAI21X1 g6695(.A0(n7910), .A1(n5855), .B0(n7911), .Y(n7912));
  NOR3X1  g6696(.A(n7912), .B(n7908), .C(n7905), .Y(n7913));
  NAND3X1 g6697(.A(n7913), .B(n7902), .C(n7896), .Y(P2_U3264));
  XOR2X1  g6698(.A(n6812), .B(P2_REG2_REG_18__SCAN_IN), .Y(n7915));
  XOR2X1  g6699(.A(n7915), .B(n7816), .Y(n7916));
  NAND2X1 g6700(.A(n7916), .B(n7755), .Y(n7917));
  OAI21X1 g6701(.A0(n6812), .A1(n5866), .B0(n7917), .Y(n7918));
  XOR2X1  g6702(.A(n6812), .B(P2_REG1_REG_18__SCAN_IN), .Y(n7919));
  XOR2X1  g6703(.A(n7919), .B(n7887), .Y(n7920));
  INVX1   g6704(.A(n7920), .Y(n7921));
  NOR2X1  g6705(.A(n7921), .B(n5864), .Y(n7922));
  OAI21X1 g6706(.A0(n7922), .A1(n7918), .B0(n7754), .Y(n7923));
  NOR2X1  g6707(.A(n7921), .B(n7900), .Y(n7924));
  OAI21X1 g6708(.A0(n7924), .A1(n7918), .B0(P2_U3966), .Y(n7925));
  NAND2X1 g6709(.A(n7916), .B(n7903), .Y(n7926));
  AOI22X1 g6710(.A0(P2_ADDR_REG_18__SCAN_IN), .A1(n7753), .B0(P2_REG3_REG_18__SCAN_IN), .B1(P2_U3152), .Y(n7927));
  OAI21X1 g6711(.A0(n7910), .A1(n6812), .B0(n7927), .Y(n7928));
  AOI21X1 g6712(.A0(n7920), .A1(n7906), .B0(n7928), .Y(n7929));
  NAND4X1 g6713(.A(n7926), .B(n7925), .C(n7923), .D(n7929), .Y(P2_U3263));
  NOR2X1  g6714(.A(n7812), .B(n7811), .Y(n7931));
  OAI21X1 g6715(.A0(n6750), .A1(n7632), .B0(n7758), .Y(n7932));
  AOI21X1 g6716(.A0(n6701), .A1(n7623), .B0(n7810), .Y(n7933));
  XOR2X1  g6717(.A(n6750), .B(P2_REG2_REG_17__SCAN_IN), .Y(n7934));
  OAI21X1 g6718(.A0(n6701), .A1(n7623), .B0(n7934), .Y(n7935));
  OAI22X1 g6719(.A0(n7933), .A1(n7935), .B0(n7932), .B1(n7931), .Y(n7936));
  OAI22X1 g6720(.A0(n7756), .A1(n7936), .B0(n6750), .B1(n5866), .Y(n7937));
  NOR2X1  g6721(.A(n6701), .B(n7826), .Y(n7938));
  NOR2X1  g6722(.A(n7938), .B(n7882), .Y(n7939));
  OAI21X1 g6723(.A0(n6750), .A1(n7827), .B0(n7828), .Y(n7940));
  NOR2X1  g6724(.A(n6702), .B(P2_REG1_REG_16__SCAN_IN), .Y(n7941));
  XOR2X1  g6725(.A(n6750), .B(n7827), .Y(n7942));
  NOR2X1  g6726(.A(n7942), .B(n7938), .Y(n7943));
  OAI21X1 g6727(.A0(n7881), .A1(n7941), .B0(n7943), .Y(n7944));
  OAI21X1 g6728(.A0(n7940), .A1(n7939), .B0(n7944), .Y(n7945));
  NOR2X1  g6729(.A(n7945), .B(n5864), .Y(n7946));
  OAI21X1 g6730(.A0(n7946), .A1(n7937), .B0(n7754), .Y(n7947));
  NOR2X1  g6731(.A(n7945), .B(n7900), .Y(n7948));
  OAI21X1 g6732(.A0(n7948), .A1(n7937), .B0(P2_U3966), .Y(n7949));
  NOR2X1  g6733(.A(n7936), .B(n7904), .Y(n7950));
  NOR2X1  g6734(.A(n7945), .B(n7907), .Y(n7951));
  AOI22X1 g6735(.A0(P2_ADDR_REG_17__SCAN_IN), .A1(n7753), .B0(P2_REG3_REG_17__SCAN_IN), .B1(P2_U3152), .Y(n7952));
  OAI21X1 g6736(.A0(n7910), .A1(n6750), .B0(n7952), .Y(n7953));
  NOR3X1  g6737(.A(n7953), .B(n7951), .C(n7950), .Y(n7954));
  NAND3X1 g6738(.A(n7954), .B(n7949), .C(n7947), .Y(P2_U3262));
  INVX1   g6739(.A(n7754), .Y(n7956));
  XOR2X1  g6740(.A(n6701), .B(n7623), .Y(n7957));
  NOR2X1  g6741(.A(n7957), .B(n7810), .Y(n7959));
  AOI21X1 g6742(.A0(n7957), .A1(n7810), .B0(n7959), .Y(n7960));
  OAI22X1 g6743(.A0(n7756), .A1(n7960), .B0(n6701), .B1(n5866), .Y(n7961));
  XOR2X1  g6744(.A(n6701), .B(P2_REG1_REG_16__SCAN_IN), .Y(n7962));
  OAI21X1 g6745(.A0(n7938), .A1(n7941), .B0(n7882), .Y(n7963));
  OAI21X1 g6746(.A0(n7962), .A1(n7882), .B0(n7963), .Y(n7964));
  AOI21X1 g6747(.A0(n7964), .A1(n5869), .B0(n7961), .Y(n7965));
  AOI21X1 g6748(.A0(n7964), .A1(n7899), .B0(n7961), .Y(n7966));
  NOR2X1  g6749(.A(n7966), .B(n7897), .Y(n7967));
  AOI22X1 g6750(.A0(P2_ADDR_REG_16__SCAN_IN), .A1(n7753), .B0(P2_REG3_REG_16__SCAN_IN), .B1(P2_U3152), .Y(n7968));
  OAI21X1 g6751(.A0(n7910), .A1(n6701), .B0(n7968), .Y(n7969));
  AOI21X1 g6752(.A0(n7964), .A1(n7906), .B0(n7969), .Y(n7970));
  OAI21X1 g6753(.A0(n7960), .A1(n7904), .B0(n7970), .Y(n7971));
  NOR2X1  g6754(.A(n7971), .B(n7967), .Y(n7972));
  OAI21X1 g6755(.A0(n7965), .A1(n7956), .B0(n7972), .Y(P2_U3261));
  XOR2X1  g6756(.A(n6654), .B(P2_REG2_REG_15__SCAN_IN), .Y(n7974));
  XOR2X1  g6757(.A(n7974), .B(n7808), .Y(n7975));
  NAND2X1 g6758(.A(n7975), .B(n7755), .Y(n7976));
  OAI21X1 g6759(.A0(n6654), .A1(n5866), .B0(n7976), .Y(n7977));
  XOR2X1  g6760(.A(n6654), .B(n7829), .Y(n7978));
  XOR2X1  g6761(.A(n7978), .B(n7879), .Y(n7979));
  NOR2X1  g6762(.A(n7979), .B(n5864), .Y(n7980));
  OAI21X1 g6763(.A0(n7980), .A1(n7977), .B0(n7754), .Y(n7981));
  NOR2X1  g6764(.A(n7979), .B(n7900), .Y(n7982));
  OAI21X1 g6765(.A0(n7982), .A1(n7977), .B0(P2_U3966), .Y(n7983));
  NAND2X1 g6766(.A(n7975), .B(n7903), .Y(n7984));
  NOR2X1  g6767(.A(n7979), .B(n7907), .Y(n7985));
  AOI22X1 g6768(.A0(P2_ADDR_REG_15__SCAN_IN), .A1(n7753), .B0(P2_REG3_REG_15__SCAN_IN), .B1(P2_U3152), .Y(n7986));
  OAI21X1 g6769(.A0(n7910), .A1(n6654), .B0(n7986), .Y(n7987));
  NOR2X1  g6770(.A(n7987), .B(n7985), .Y(n7988));
  NAND4X1 g6771(.A(n7984), .B(n7983), .C(n7981), .D(n7988), .Y(P2_U3260));
  XOR2X1  g6772(.A(n6606), .B(P2_REG2_REG_14__SCAN_IN), .Y(n7990));
  XOR2X1  g6773(.A(n7990), .B(n7806), .Y(n7991));
  NAND2X1 g6774(.A(n7991), .B(n7755), .Y(n7992));
  OAI21X1 g6775(.A0(n6606), .A1(n5866), .B0(n7992), .Y(n7993));
  XOR2X1  g6776(.A(n6606), .B(P2_REG1_REG_14__SCAN_IN), .Y(n7994));
  XOR2X1  g6777(.A(n7994), .B(n7878), .Y(n7995));
  NOR2X1  g6778(.A(n7995), .B(n5864), .Y(n7996));
  OAI21X1 g6779(.A0(n7996), .A1(n7993), .B0(n7754), .Y(n7997));
  NOR2X1  g6780(.A(n7995), .B(n7900), .Y(n7998));
  OAI21X1 g6781(.A0(n7998), .A1(n7993), .B0(P2_U3966), .Y(n7999));
  NAND2X1 g6782(.A(n7991), .B(n7903), .Y(n8000));
  NOR2X1  g6783(.A(n7995), .B(n7907), .Y(n8001));
  AOI22X1 g6784(.A0(P2_ADDR_REG_14__SCAN_IN), .A1(n7753), .B0(P2_REG3_REG_14__SCAN_IN), .B1(P2_U3152), .Y(n8002));
  OAI21X1 g6785(.A0(n7910), .A1(n6606), .B0(n8002), .Y(n8003));
  NOR2X1  g6786(.A(n8003), .B(n8001), .Y(n8004));
  NAND4X1 g6787(.A(n8000), .B(n7999), .C(n7997), .D(n8004), .Y(P2_U3259));
  NAND2X1 g6788(.A(n6440), .B(n6420), .Y(n8006));
  AOI21X1 g6789(.A0(n8006), .A1(n7804), .B0(n7762), .Y(n8007));
  INVX1   g6790(.A(n8007), .Y(n8008));
  AOI21X1 g6791(.A0(n6556), .A1(P2_REG2_REG_13__SCAN_IN), .B0(n7765), .Y(n8009));
  OAI21X1 g6792(.A0(n8008), .A1(n7766), .B0(n8009), .Y(n8010));
  NOR2X1  g6793(.A(n6504), .B(P2_REG2_REG_12__SCAN_IN), .Y(n8011));
  XOR2X1  g6794(.A(n6555), .B(n7760), .Y(n8012));
  NOR2X1  g6795(.A(n8012), .B(n7766), .Y(n8013));
  OAI21X1 g6796(.A0(n8007), .A1(n8011), .B0(n8013), .Y(n8014));
  NAND2X1 g6797(.A(n8014), .B(n8010), .Y(n8015));
  OAI22X1 g6798(.A0(n7756), .A1(n8015), .B0(n6555), .B1(n5866), .Y(n8016));
  INVX1   g6799(.A(n7876), .Y(n8017));
  NOR2X1  g6800(.A(n6441), .B(P2_REG1_REG_11__SCAN_IN), .Y(n8018));
  INVX1   g6801(.A(n8018), .Y(n8019));
  AOI21X1 g6802(.A0(n8019), .A1(n8017), .B0(n7832), .Y(n8020));
  INVX1   g6803(.A(n8020), .Y(n8021));
  AOI21X1 g6804(.A0(n6556), .A1(P2_REG1_REG_13__SCAN_IN), .B0(n7836), .Y(n8022));
  OAI21X1 g6805(.A0(n8021), .A1(n7837), .B0(n8022), .Y(n8023));
  NOR2X1  g6806(.A(n6504), .B(P2_REG1_REG_12__SCAN_IN), .Y(n8024));
  XOR2X1  g6807(.A(n6555), .B(n6539), .Y(n8025));
  NOR2X1  g6808(.A(n8025), .B(n7837), .Y(n8026));
  OAI21X1 g6809(.A0(n8020), .A1(n8024), .B0(n8026), .Y(n8027));
  NAND2X1 g6810(.A(n8027), .B(n8023), .Y(n8028));
  NOR2X1  g6811(.A(n8028), .B(n5864), .Y(n8029));
  OAI21X1 g6812(.A0(n8029), .A1(n8016), .B0(n7754), .Y(n8030));
  NOR2X1  g6813(.A(n8028), .B(n7900), .Y(n8031));
  OAI21X1 g6814(.A0(n8031), .A1(n8016), .B0(P2_U3966), .Y(n8032));
  NOR2X1  g6815(.A(n8015), .B(n7904), .Y(n8033));
  NOR2X1  g6816(.A(n8028), .B(n7907), .Y(n8034));
  AOI22X1 g6817(.A0(P2_ADDR_REG_13__SCAN_IN), .A1(n7753), .B0(P2_REG3_REG_13__SCAN_IN), .B1(P2_U3152), .Y(n8035));
  OAI21X1 g6818(.A0(n7910), .A1(n6555), .B0(n8035), .Y(n8036));
  NOR3X1  g6819(.A(n8036), .B(n8034), .C(n8033), .Y(n8037));
  NAND3X1 g6820(.A(n8037), .B(n8032), .C(n8030), .Y(P2_U3258));
  XOR2X1  g6821(.A(n6503), .B(n7589), .Y(n8039));
  NOR2X1  g6822(.A(n8039), .B(n8007), .Y(n8041));
  AOI21X1 g6823(.A0(n8039), .A1(n8007), .B0(n8041), .Y(n8042));
  OAI22X1 g6824(.A0(n7756), .A1(n8042), .B0(n6503), .B1(n5866), .Y(n8043));
  XOR2X1  g6825(.A(n6503), .B(P2_REG1_REG_12__SCAN_IN), .Y(n8044));
  OAI21X1 g6826(.A0(n7837), .A1(n8024), .B0(n8021), .Y(n8045));
  OAI21X1 g6827(.A0(n8044), .A1(n8021), .B0(n8045), .Y(n8046));
  AOI21X1 g6828(.A0(n8046), .A1(n5869), .B0(n8043), .Y(n8047));
  AOI21X1 g6829(.A0(n8046), .A1(n7899), .B0(n8043), .Y(n8048));
  NOR2X1  g6830(.A(n8048), .B(n7897), .Y(n8049));
  AOI22X1 g6831(.A0(P2_ADDR_REG_12__SCAN_IN), .A1(n7753), .B0(P2_REG3_REG_12__SCAN_IN), .B1(P2_U3152), .Y(n8050));
  OAI21X1 g6832(.A0(n7910), .A1(n6503), .B0(n8050), .Y(n8051));
  AOI21X1 g6833(.A0(n8046), .A1(n7906), .B0(n8051), .Y(n8052));
  OAI21X1 g6834(.A0(n8042), .A1(n7904), .B0(n8052), .Y(n8053));
  NOR2X1  g6835(.A(n8053), .B(n8049), .Y(n8054));
  OAI21X1 g6836(.A0(n8047), .A1(n7956), .B0(n8054), .Y(P2_U3257));
  XOR2X1  g6837(.A(n6440), .B(n6420), .Y(n8056));
  AOI21X1 g6838(.A0(n8006), .A1(n7763), .B0(n7803), .Y(n8057));
  AOI21X1 g6839(.A0(n8056), .A1(n7803), .B0(n8057), .Y(n8058));
  OAI22X1 g6840(.A0(n7756), .A1(n8058), .B0(n6440), .B1(n5866), .Y(n8059));
  XOR2X1  g6841(.A(n6440), .B(n6423), .Y(n8060));
  AOI21X1 g6842(.A0(n8019), .A1(n7833), .B0(n7876), .Y(n8061));
  AOI21X1 g6843(.A0(n8060), .A1(n7876), .B0(n8061), .Y(n8062));
  NOR2X1  g6844(.A(n8062), .B(n5864), .Y(n8063));
  OAI21X1 g6845(.A0(n8063), .A1(n8059), .B0(n7754), .Y(n8064));
  NOR2X1  g6846(.A(n8062), .B(n7900), .Y(n8065));
  OAI21X1 g6847(.A0(n8065), .A1(n8059), .B0(P2_U3966), .Y(n8066));
  AOI22X1 g6848(.A0(P2_ADDR_REG_11__SCAN_IN), .A1(n7753), .B0(P2_REG3_REG_11__SCAN_IN), .B1(P2_U3152), .Y(n8067));
  OAI21X1 g6849(.A0(n7910), .A1(n6440), .B0(n8067), .Y(n8068));
  OAI22X1 g6850(.A0(n8058), .A1(n7904), .B0(n7907), .B1(n8062), .Y(n8069));
  NOR2X1  g6851(.A(n8069), .B(n8068), .Y(n8070));
  NAND3X1 g6852(.A(n8070), .B(n8066), .C(n8064), .Y(P2_U3256));
  NAND2X1 g6853(.A(n6389), .B(P2_REG2_REG_10__SCAN_IN), .Y(n8072));
  AOI21X1 g6854(.A0(n7800), .A1(n7798), .B0(n7769), .Y(n8073));
  NAND2X1 g6855(.A(n8073), .B(n7771), .Y(n8074));
  NAND3X1 g6856(.A(n8074), .B(n8072), .C(n7770), .Y(n8075));
  AOI21X1 g6857(.A0(n6335), .A1(n6318), .B0(n8073), .Y(n8076));
  AOI22X1 g6858(.A0(n6336), .A1(P2_REG2_REG_9__SCAN_IN), .B0(n6366), .B1(n6389), .Y(n8077));
  OAI21X1 g6859(.A0(n6389), .A1(n6366), .B0(n8077), .Y(n8078));
  OAI21X1 g6860(.A0(n8078), .A1(n8076), .B0(n8075), .Y(n8079));
  OAI22X1 g6861(.A0(n7756), .A1(n8079), .B0(n6388), .B1(n5866), .Y(n8080));
  NAND2X1 g6862(.A(n6389), .B(P2_REG1_REG_10__SCAN_IN), .Y(n8081));
  AOI21X1 g6863(.A0(n7873), .A1(n7871), .B0(n7841), .Y(n8082));
  NAND2X1 g6864(.A(n8082), .B(n7843), .Y(n8083));
  NAND3X1 g6865(.A(n8083), .B(n8081), .C(n7842), .Y(n8084));
  AOI21X1 g6866(.A0(n6335), .A1(n6321), .B0(n8082), .Y(n8085));
  AOI22X1 g6867(.A0(n6336), .A1(P2_REG1_REG_9__SCAN_IN), .B0(n6369), .B1(n6389), .Y(n8086));
  OAI21X1 g6868(.A0(n6389), .A1(n6369), .B0(n8086), .Y(n8087));
  OAI21X1 g6869(.A0(n8087), .A1(n8085), .B0(n8084), .Y(n8088));
  NOR2X1  g6870(.A(n8088), .B(n5864), .Y(n8089));
  OAI21X1 g6871(.A0(n8089), .A1(n8080), .B0(n7754), .Y(n8090));
  NOR2X1  g6872(.A(n8088), .B(n7900), .Y(n8091));
  OAI21X1 g6873(.A0(n8091), .A1(n8080), .B0(P2_U3966), .Y(n8092));
  NOR2X1  g6874(.A(n8079), .B(n7904), .Y(n8093));
  NOR2X1  g6875(.A(n8088), .B(n7907), .Y(n8094));
  AOI22X1 g6876(.A0(P2_ADDR_REG_10__SCAN_IN), .A1(n7753), .B0(P2_REG3_REG_10__SCAN_IN), .B1(P2_U3152), .Y(n8095));
  OAI21X1 g6877(.A0(n7910), .A1(n6388), .B0(n8095), .Y(n8096));
  NOR3X1  g6878(.A(n8096), .B(n8094), .C(n8093), .Y(n8097));
  NAND3X1 g6879(.A(n8097), .B(n8092), .C(n8090), .Y(P2_U3255));
  XOR2X1  g6880(.A(n6335), .B(n6318), .Y(n8099));
  NOR2X1  g6881(.A(n8099), .B(n8073), .Y(n8101));
  AOI21X1 g6882(.A0(n8099), .A1(n8073), .B0(n8101), .Y(n8102));
  OAI22X1 g6883(.A0(n7756), .A1(n8102), .B0(n6335), .B1(n5866), .Y(n8103));
  XOR2X1  g6884(.A(n6335), .B(n6321), .Y(n8104));
  NOR2X1  g6885(.A(n8104), .B(n8082), .Y(n8106));
  AOI21X1 g6886(.A0(n8104), .A1(n8082), .B0(n8106), .Y(n8107));
  NOR2X1  g6887(.A(n8107), .B(n5864), .Y(n8108));
  OAI21X1 g6888(.A0(n8108), .A1(n8103), .B0(n7754), .Y(n8109));
  NOR2X1  g6889(.A(n8107), .B(n7900), .Y(n8110));
  OAI21X1 g6890(.A0(n8110), .A1(n8103), .B0(P2_U3966), .Y(n8111));
  AOI22X1 g6891(.A0(P2_ADDR_REG_9__SCAN_IN), .A1(n7753), .B0(P2_REG3_REG_9__SCAN_IN), .B1(P2_U3152), .Y(n8112));
  OAI21X1 g6892(.A0(n7910), .A1(n6335), .B0(n8112), .Y(n8113));
  OAI22X1 g6893(.A0(n8102), .A1(n7904), .B0(n7907), .B1(n8107), .Y(n8114));
  NOR2X1  g6894(.A(n8114), .B(n8113), .Y(n8115));
  NAND3X1 g6895(.A(n8115), .B(n8111), .C(n8109), .Y(P2_U3254));
  XOR2X1  g6896(.A(n6286), .B(P2_REG2_REG_8__SCAN_IN), .Y(n8117));
  NOR2X1  g6897(.A(n8117), .B(n7798), .Y(n8118));
  AOI21X1 g6898(.A0(n8117), .A1(n7798), .B0(n8118), .Y(n8120));
  INVX1   g6899(.A(n8120), .Y(n8121));
  NAND2X1 g6900(.A(n8121), .B(n7903), .Y(n8122));
  AOI22X1 g6901(.A0(P2_ADDR_REG_8__SCAN_IN), .A1(n7753), .B0(P2_REG3_REG_8__SCAN_IN), .B1(P2_U3152), .Y(n8123));
  XOR2X1  g6902(.A(n6286), .B(P2_REG1_REG_8__SCAN_IN), .Y(n8124));
  OAI21X1 g6903(.A0(n7872), .A1(n7841), .B0(n7871), .Y(n8125));
  OAI21X1 g6904(.A0(n8124), .A1(n7871), .B0(n8125), .Y(n8126));
  AOI22X1 g6905(.A0(n7909), .A1(n6287), .B0(n7906), .B1(n8126), .Y(n8127));
  OAI22X1 g6906(.A0(n7756), .A1(n8120), .B0(n6286), .B1(n5866), .Y(n8128));
  AOI21X1 g6907(.A0(n8126), .A1(n7899), .B0(n8128), .Y(n8129));
  NOR2X1  g6908(.A(n8129), .B(n7897), .Y(n8130));
  AOI21X1 g6909(.A0(n8126), .A1(n5869), .B0(n8128), .Y(n8131));
  NOR2X1  g6910(.A(n8131), .B(n7956), .Y(n8132));
  NOR2X1  g6911(.A(n8132), .B(n8130), .Y(n8133));
  NAND4X1 g6912(.A(n8127), .B(n8123), .C(n8122), .D(n8133), .Y(P2_U3253));
  NOR2X1  g6913(.A(n6182), .B(n6163), .Y(n8135));
  INVX1   g6914(.A(n7775), .Y(n8136));
  AOI21X1 g6915(.A0(n6237), .A1(P2_REG2_REG_7__SCAN_IN), .B0(n8136), .Y(n8137));
  OAI21X1 g6916(.A0(n8135), .A1(n7793), .B0(n8137), .Y(n8138));
  AOI22X1 g6917(.A0(n7788), .A1(n7792), .B0(n6182), .B1(n6163), .Y(n8139));
  AOI21X1 g6918(.A0(n6237), .A1(n6216), .B0(n8135), .Y(n8140));
  OAI21X1 g6919(.A0(n6237), .A1(n6216), .B0(n8140), .Y(n8141));
  OAI21X1 g6920(.A0(n8141), .A1(n8139), .B0(n8138), .Y(n8142));
  NOR2X1  g6921(.A(n8142), .B(n7904), .Y(n8143));
  INVX1   g6922(.A(n7753), .Y(n8144));
  OAI22X1 g6923(.A0(n1048), .A1(n8144), .B0(n6271), .B1(P2_STATE_REG_SCAN_IN), .Y(n8145));
  NOR2X1  g6924(.A(n8145), .B(n8143), .Y(n8146));
  NOR2X1  g6925(.A(n6182), .B(n7847), .Y(n8147));
  INVX1   g6926(.A(n7848), .Y(n8148));
  AOI21X1 g6927(.A0(n6237), .A1(P2_REG1_REG_7__SCAN_IN), .B0(n8148), .Y(n8149));
  OAI21X1 g6928(.A0(n8147), .A1(n7866), .B0(n8149), .Y(n8150));
  AOI22X1 g6929(.A0(n7862), .A1(n7865), .B0(n6182), .B1(n7847), .Y(n8151));
  AOI21X1 g6930(.A0(n6237), .A1(n6219), .B0(n8147), .Y(n8152));
  OAI21X1 g6931(.A0(n6237), .A1(n6219), .B0(n8152), .Y(n8153));
  OAI21X1 g6932(.A0(n8153), .A1(n8151), .B0(n8150), .Y(n8154));
  NOR2X1  g6933(.A(n8154), .B(n7900), .Y(n8155));
  OAI22X1 g6934(.A0(n7756), .A1(n8142), .B0(n6236), .B1(n5866), .Y(n8156));
  OAI21X1 g6935(.A0(n8156), .A1(n8155), .B0(P2_U3966), .Y(n8157));
  NOR2X1  g6936(.A(n8154), .B(n5864), .Y(n8158));
  OAI21X1 g6937(.A0(n8158), .A1(n8156), .B0(n7754), .Y(n8159));
  NOR2X1  g6938(.A(n8154), .B(n7907), .Y(n8160));
  AOI21X1 g6939(.A0(n7909), .A1(n6237), .B0(n8160), .Y(n8161));
  NAND4X1 g6940(.A(n8159), .B(n8157), .C(n8146), .D(n8161), .Y(P2_U3252));
  XOR2X1  g6941(.A(n6182), .B(P2_REG2_REG_6__SCAN_IN), .Y(n8163));
  NOR2X1  g6942(.A(n8163), .B(n7793), .Y(n8164));
  AOI21X1 g6943(.A0(n8163), .A1(n7793), .B0(n8164), .Y(n8166));
  OAI22X1 g6944(.A0(n7756), .A1(n8166), .B0(n6182), .B1(n5866), .Y(n8167));
  XOR2X1  g6945(.A(n6182), .B(P2_REG1_REG_6__SCAN_IN), .Y(n8168));
  NOR2X1  g6946(.A(n8168), .B(n7866), .Y(n8169));
  AOI21X1 g6947(.A0(n8168), .A1(n7866), .B0(n8169), .Y(n8171));
  NOR2X1  g6948(.A(n8171), .B(n5864), .Y(n8172));
  OAI21X1 g6949(.A0(n8172), .A1(n8167), .B0(n7754), .Y(n8173));
  NOR2X1  g6950(.A(n8171), .B(n7900), .Y(n8174));
  OAI21X1 g6951(.A0(n8174), .A1(n8167), .B0(P2_U3966), .Y(n8175));
  AOI22X1 g6952(.A0(P2_ADDR_REG_6__SCAN_IN), .A1(n7753), .B0(P2_REG3_REG_6__SCAN_IN), .B1(P2_U3152), .Y(n8176));
  NOR2X1  g6953(.A(n8171), .B(n7907), .Y(n8177));
  OAI22X1 g6954(.A0(n7910), .A1(n6182), .B0(n7904), .B1(n8166), .Y(n8178));
  NOR2X1  g6955(.A(n8178), .B(n8177), .Y(n8179));
  NAND4X1 g6956(.A(n8176), .B(n8175), .C(n8173), .D(n8179), .Y(P2_U3251));
  NOR2X1  g6957(.A(n6074), .B(n6087), .Y(n8181));
  INVX1   g6958(.A(n7780), .Y(n8182));
  NOR2X1  g6959(.A(n8182), .B(n7777), .Y(n8183));
  NOR2X1  g6960(.A(n5987), .B(n5969), .Y(n8184));
  NOR2X1  g6961(.A(n5988), .B(P2_REG2_REG_2__SCAN_IN), .Y(n8185));
  NOR3X1  g6962(.A(n8185), .B(n5936), .C(n5949), .Y(n8186));
  NOR2X1  g6963(.A(n8186), .B(n8184), .Y(n8187));
  NOR2X1  g6964(.A(n8187), .B(n7784), .Y(n8188));
  NOR4X1  g6965(.A(n8183), .B(n8181), .C(n7783), .D(n8188), .Y(n8189));
  OAI21X1 g6966(.A0(n6130), .A1(n6114), .B0(n7776), .Y(n8190));
  NOR3X1  g6967(.A(n8188), .B(n8183), .C(n7783), .Y(n8191));
  AOI21X1 g6968(.A0(n6074), .A1(n6087), .B0(n8191), .Y(n8192));
  AOI21X1 g6969(.A0(n7789), .A1(n6114), .B0(n8181), .Y(n8193));
  OAI21X1 g6970(.A0(n7789), .A1(n6114), .B0(n8193), .Y(n8194));
  OAI22X1 g6971(.A0(n8192), .A1(n8194), .B0(n8190), .B1(n8189), .Y(n8195));
  OAI22X1 g6972(.A0(n7756), .A1(n8195), .B0(n6130), .B1(n5866), .Y(n8196));
  NOR2X1  g6973(.A(n6074), .B(n6090), .Y(n8197));
  INVX1   g6974(.A(n7854), .Y(n8198));
  NOR2X1  g6975(.A(n8198), .B(n7851), .Y(n8199));
  NOR2X1  g6976(.A(n5988), .B(P2_REG1_REG_2__SCAN_IN), .Y(n8200));
  NOR3X1  g6977(.A(n8200), .B(n5936), .C(n5948), .Y(n8201));
  AOI21X1 g6978(.A0(n5988), .A1(P2_REG1_REG_2__SCAN_IN), .B0(n8201), .Y(n8202));
  NOR2X1  g6979(.A(n8202), .B(n7858), .Y(n8203));
  NOR4X1  g6980(.A(n8199), .B(n8197), .C(n7857), .D(n8203), .Y(n8204));
  OAI21X1 g6981(.A0(n6130), .A1(n6117), .B0(n7849), .Y(n8205));
  NOR3X1  g6982(.A(n8203), .B(n8199), .C(n7857), .Y(n8206));
  AOI21X1 g6983(.A0(n6074), .A1(n6090), .B0(n8206), .Y(n8207));
  AOI21X1 g6984(.A0(n7789), .A1(n6117), .B0(n8197), .Y(n8208));
  OAI21X1 g6985(.A0(n7789), .A1(n6117), .B0(n8208), .Y(n8209));
  OAI22X1 g6986(.A0(n8207), .A1(n8209), .B0(n8205), .B1(n8204), .Y(n8210));
  NOR2X1  g6987(.A(n8210), .B(n5864), .Y(n8211));
  OAI21X1 g6988(.A0(n8211), .A1(n8196), .B0(n7754), .Y(n8212));
  NOR2X1  g6989(.A(n8210), .B(n7900), .Y(n8213));
  OAI21X1 g6990(.A0(n8213), .A1(n8196), .B0(P2_U3966), .Y(n8214));
  AOI22X1 g6991(.A0(P2_ADDR_REG_5__SCAN_IN), .A1(n7753), .B0(P2_REG3_REG_5__SCAN_IN), .B1(P2_U3152), .Y(n8215));
  NOR2X1  g6992(.A(n8210), .B(n7907), .Y(n8216));
  OAI22X1 g6993(.A0(n7910), .A1(n6130), .B0(n7904), .B1(n8195), .Y(n8217));
  NOR2X1  g6994(.A(n8217), .B(n8216), .Y(n8218));
  NAND4X1 g6995(.A(n8215), .B(n8214), .C(n8212), .D(n8218), .Y(P2_U3250));
  XOR2X1  g6996(.A(n6074), .B(n6087), .Y(n8220));
  NOR2X1  g6997(.A(n8220), .B(n8191), .Y(n8222));
  AOI21X1 g6998(.A0(n8220), .A1(n8191), .B0(n8222), .Y(n8223));
  OAI22X1 g6999(.A0(n7756), .A1(n8223), .B0(n6074), .B1(n5866), .Y(n8224));
  XOR2X1  g7000(.A(n6074), .B(n6090), .Y(n8225));
  NOR2X1  g7001(.A(n8225), .B(n8206), .Y(n8227));
  AOI21X1 g7002(.A0(n8225), .A1(n8206), .B0(n8227), .Y(n8228));
  NOR2X1  g7003(.A(n8228), .B(n5864), .Y(n8229));
  OAI21X1 g7004(.A0(n8229), .A1(n8224), .B0(n7754), .Y(n8230));
  NOR2X1  g7005(.A(n8228), .B(n7900), .Y(n8231));
  OAI21X1 g7006(.A0(n8231), .A1(n8224), .B0(P2_U3966), .Y(n8232));
  AOI22X1 g7007(.A0(P2_ADDR_REG_4__SCAN_IN), .A1(n7753), .B0(P2_REG3_REG_4__SCAN_IN), .B1(P2_U3152), .Y(n8233));
  NOR2X1  g7008(.A(n8228), .B(n7907), .Y(n8234));
  OAI22X1 g7009(.A0(n7910), .A1(n6074), .B0(n7904), .B1(n8223), .Y(n8235));
  NOR2X1  g7010(.A(n8235), .B(n8234), .Y(n8236));
  NAND4X1 g7011(.A(n8233), .B(n8232), .C(n8230), .D(n8236), .Y(P2_U3249));
  OAI21X1 g7012(.A0(n8182), .A1(n8185), .B0(n8187), .Y(n8238));
  XOR2X1  g7013(.A(n6030), .B(P2_REG2_REG_3__SCAN_IN), .Y(n8239));
  OAI21X1 g7014(.A0(n7783), .A1(n7784), .B0(n8238), .Y(n8240));
  OAI21X1 g7015(.A0(n8239), .A1(n8238), .B0(n8240), .Y(n8241));
  NAND2X1 g7016(.A(n8241), .B(n7903), .Y(n8242));
  AOI22X1 g7017(.A0(n7755), .A1(n8241), .B0(n6031), .B1(n5871), .Y(n8243));
  OAI21X1 g7018(.A0(n8198), .A1(n8200), .B0(n8202), .Y(n8244));
  XOR2X1  g7019(.A(n6030), .B(P2_REG1_REG_3__SCAN_IN), .Y(n8245));
  NOR2X1  g7020(.A(n8245), .B(n8244), .Y(n8246));
  AOI21X1 g7021(.A0(n8245), .A1(n8244), .B0(n8246), .Y(n8248));
  INVX1   g7022(.A(n8248), .Y(n8249));
  NAND2X1 g7023(.A(n8249), .B(n5869), .Y(n8250));
  AOI21X1 g7024(.A0(n8250), .A1(n8243), .B0(n7956), .Y(n8251));
  NOR2X1  g7025(.A(n8144), .B(n1053), .Y(n8252));
  NAND2X1 g7026(.A(n8249), .B(n7899), .Y(n8253));
  AOI21X1 g7027(.A0(n8253), .A1(n8243), .B0(n7897), .Y(n8254));
  NOR2X1  g7028(.A(n6026), .B(P2_STATE_REG_SCAN_IN), .Y(n8255));
  NOR4X1  g7029(.A(n8254), .B(n8252), .C(n8251), .D(n8255), .Y(n8256));
  AOI22X1 g7030(.A0(n7909), .A1(n6031), .B0(n7906), .B1(n8249), .Y(n8257));
  NAND3X1 g7031(.A(n8257), .B(n8256), .C(n8242), .Y(P2_U3248));
  NOR3X1  g7032(.A(n8184), .B(n7782), .C(n8185), .Y(n8259));
  XOR2X1  g7033(.A(n5987), .B(n5969), .Y(n8260));
  NOR3X1  g7034(.A(n8260), .B(n7781), .C(n7780), .Y(n8261));
  NOR2X1  g7035(.A(n8261), .B(n8259), .Y(n8262));
  NAND2X1 g7036(.A(n8262), .B(n7903), .Y(n8263));
  NOR4X1  g7037(.A(n8259), .B(n5871), .C(n5869), .D(n8261), .Y(n8264));
  INVX1   g7038(.A(n7856), .Y(n8265));
  XOR2X1  g7039(.A(n5987), .B(n5968), .Y(n8266));
  NOR3X1  g7040(.A(n8266), .B(n7855), .C(n7854), .Y(n8268));
  AOI21X1 g7041(.A0(n8266), .A1(n8265), .B0(n8268), .Y(n8269));
  INVX1   g7042(.A(n8269), .Y(n8270));
  OAI22X1 g7043(.A0(n5987), .A1(n5866), .B0(n5864), .B1(n8270), .Y(n8271));
  OAI21X1 g7044(.A0(n8271), .A1(n8264), .B0(n7754), .Y(n8272));
  NOR2X1  g7045(.A(n5987), .B(n5866), .Y(n8273));
  NOR2X1  g7046(.A(n8270), .B(n7900), .Y(n8274));
  NOR3X1  g7047(.A(n8274), .B(n8273), .C(n8264), .Y(n8275));
  OAI22X1 g7048(.A0(n7897), .A1(n8275), .B0(n5971), .B1(P2_STATE_REG_SCAN_IN), .Y(n8276));
  AOI21X1 g7049(.A0(n7753), .A1(P2_ADDR_REG_2__SCAN_IN), .B0(n8276), .Y(n8277));
  AOI22X1 g7050(.A0(n7909), .A1(n5988), .B0(n7906), .B1(n8269), .Y(n8278));
  NAND4X1 g7051(.A(n8277), .B(n8272), .C(n8263), .D(n8278), .Y(P2_U3247));
  XOR2X1  g7052(.A(n5936), .B(n5949), .Y(n8280));
  XOR2X1  g7053(.A(n8280), .B(n7779), .Y(n8281));
  INVX1   g7054(.A(n8281), .Y(n8282));
  NAND2X1 g7055(.A(n8282), .B(n7903), .Y(n8283));
  XOR2X1  g7056(.A(n5936), .B(n5948), .Y(n8284));
  XOR2X1  g7057(.A(n8284), .B(n7853), .Y(n8285));
  INVX1   g7058(.A(n8285), .Y(n8286));
  AOI22X1 g7059(.A0(n5937), .A1(n5871), .B0(n5869), .B1(n8286), .Y(n8287));
  OAI21X1 g7060(.A0(n8281), .A1(n7756), .B0(n8287), .Y(n8288));
  NAND2X1 g7061(.A(n8288), .B(n7754), .Y(n8289));
  OAI22X1 g7062(.A0(n7756), .A1(n8281), .B0(n5936), .B1(n5866), .Y(n8290));
  AOI21X1 g7063(.A0(n8286), .A1(n7899), .B0(n8290), .Y(n8291));
  OAI22X1 g7064(.A0(n7897), .A1(n8291), .B0(n5951), .B1(P2_STATE_REG_SCAN_IN), .Y(n8292));
  AOI21X1 g7065(.A0(n7753), .A1(P2_ADDR_REG_1__SCAN_IN), .B0(n8292), .Y(n8293));
  AOI22X1 g7066(.A0(n7909), .A1(n5937), .B0(n7906), .B1(n8286), .Y(n8294));
  NAND4X1 g7067(.A(n8293), .B(n8289), .C(n8283), .D(n8294), .Y(P2_U3246));
  XOR2X1  g7068(.A(n5477), .B(P2_REG2_REG_0__SCAN_IN), .Y(n8296));
  INVX1   g7069(.A(n8296), .Y(n8297));
  NAND2X1 g7070(.A(n8297), .B(n7903), .Y(n8298));
  XOR2X1  g7071(.A(n5477), .B(P2_REG1_REG_0__SCAN_IN), .Y(n8299));
  INVX1   g7072(.A(n8299), .Y(n8300));
  AOI22X1 g7073(.A0(n5875), .A1(n5871), .B0(n5869), .B1(n8300), .Y(n8301));
  OAI21X1 g7074(.A0(n8296), .A1(n7756), .B0(n8301), .Y(n8302));
  NAND2X1 g7075(.A(n8302), .B(n7754), .Y(n8303));
  OAI22X1 g7076(.A0(n7756), .A1(n8296), .B0(n5477), .B1(n5866), .Y(n8304));
  AOI21X1 g7077(.A0(n8300), .A1(n7899), .B0(n8304), .Y(n8305));
  OAI22X1 g7078(.A0(n7897), .A1(n8305), .B0(n5893), .B1(P2_STATE_REG_SCAN_IN), .Y(n8306));
  AOI21X1 g7079(.A0(n7753), .A1(P2_ADDR_REG_0__SCAN_IN), .B0(n8306), .Y(n8307));
  AOI22X1 g7080(.A0(n7909), .A1(n5875), .B0(n7906), .B1(n8300), .Y(n8308));
  NAND4X1 g7081(.A(n8307), .B(n8303), .C(n8298), .D(n8308), .Y(P2_U3245));
  NAND2X1 g7082(.A(n7897), .B(P2_DATAO_REG_0__SCAN_IN), .Y(n8310));
  OAI21X1 g7083(.A0(n7897), .A1(n5897), .B0(n8310), .Y(P2_U3552));
  NAND2X1 g7084(.A(n7897), .B(P2_DATAO_REG_1__SCAN_IN), .Y(n8312));
  OAI21X1 g7085(.A0(n7897), .A1(n5954), .B0(n8312), .Y(P2_U3553));
  NAND2X1 g7086(.A(n7897), .B(P2_DATAO_REG_2__SCAN_IN), .Y(n8314));
  OAI21X1 g7087(.A0(n7897), .A1(n5974), .B0(n8314), .Y(P2_U3554));
  NAND2X1 g7088(.A(n7897), .B(P2_DATAO_REG_3__SCAN_IN), .Y(n8316));
  OAI21X1 g7089(.A0(n7897), .A1(n6015), .B0(n8316), .Y(P2_U3555));
  NAND2X1 g7090(.A(n7897), .B(P2_DATAO_REG_4__SCAN_IN), .Y(n8318));
  OAI21X1 g7091(.A0(n7897), .A1(n6092), .B0(n8318), .Y(P2_U3556));
  NAND2X1 g7092(.A(n7897), .B(P2_DATAO_REG_5__SCAN_IN), .Y(n8320));
  OAI21X1 g7093(.A0(n7897), .A1(n6121), .B0(n8320), .Y(P2_U3557));
  NAND2X1 g7094(.A(n7897), .B(P2_DATAO_REG_6__SCAN_IN), .Y(n8322));
  OAI21X1 g7095(.A0(n7897), .A1(n6172), .B0(n8322), .Y(P2_U3558));
  NAND2X1 g7096(.A(n7897), .B(P2_DATAO_REG_7__SCAN_IN), .Y(n8324));
  OAI21X1 g7097(.A0(n7897), .A1(n6223), .B0(n8324), .Y(P2_U3559));
  NAND2X1 g7098(.A(n7897), .B(P2_DATAO_REG_8__SCAN_IN), .Y(n8326));
  OAI21X1 g7099(.A0(n7897), .A1(n6275), .B0(n8326), .Y(P2_U3560));
  NAND2X1 g7100(.A(n7897), .B(P2_DATAO_REG_9__SCAN_IN), .Y(n8328));
  OAI21X1 g7101(.A0(n7897), .A1(n6327), .B0(n8328), .Y(P2_U3561));
  NAND2X1 g7102(.A(n7897), .B(P2_DATAO_REG_10__SCAN_IN), .Y(n8330));
  OAI21X1 g7103(.A0(n7897), .A1(n6374), .B0(n8330), .Y(P2_U3562));
  NAND2X1 g7104(.A(n7897), .B(P2_DATAO_REG_11__SCAN_IN), .Y(n8332));
  OAI21X1 g7105(.A0(n7897), .A1(n6430), .B0(n8332), .Y(P2_U3563));
  NAND2X1 g7106(.A(n7897), .B(P2_DATAO_REG_12__SCAN_IN), .Y(n8334));
  OAI21X1 g7107(.A0(n7897), .A1(n6494), .B0(n8334), .Y(P2_U3564));
  NAND2X1 g7108(.A(n7897), .B(P2_DATAO_REG_13__SCAN_IN), .Y(n8336));
  OAI21X1 g7109(.A0(n7897), .A1(n6546), .B0(n8336), .Y(P2_U3565));
  NAND2X1 g7110(.A(n7897), .B(P2_DATAO_REG_14__SCAN_IN), .Y(n8338));
  OAI21X1 g7111(.A0(n7897), .A1(n6597), .B0(n8338), .Y(P2_U3566));
  NAND2X1 g7112(.A(n7897), .B(P2_DATAO_REG_15__SCAN_IN), .Y(n8340));
  OAI21X1 g7113(.A0(n7897), .A1(n6646), .B0(n8340), .Y(P2_U3567));
  NAND2X1 g7114(.A(n7897), .B(P2_DATAO_REG_16__SCAN_IN), .Y(n8342));
  OAI21X1 g7115(.A0(n7897), .A1(n6690), .B0(n8342), .Y(P2_U3568));
  NAND2X1 g7116(.A(n7897), .B(P2_DATAO_REG_17__SCAN_IN), .Y(n8344));
  OAI21X1 g7117(.A0(n7897), .A1(n6740), .B0(n8344), .Y(P2_U3569));
  NAND2X1 g7118(.A(n7897), .B(P2_DATAO_REG_18__SCAN_IN), .Y(n8346));
  OAI21X1 g7119(.A0(n7897), .A1(n6799), .B0(n8346), .Y(P2_U3570));
  NAND2X1 g7120(.A(n7897), .B(P2_DATAO_REG_19__SCAN_IN), .Y(n8348));
  OAI21X1 g7121(.A0(n7897), .A1(n6846), .B0(n8348), .Y(P2_U3571));
  NAND2X1 g7122(.A(n7897), .B(P2_DATAO_REG_20__SCAN_IN), .Y(n8350));
  OAI21X1 g7123(.A0(n7897), .A1(n6894), .B0(n8350), .Y(P2_U3572));
  NAND2X1 g7124(.A(n7897), .B(P2_DATAO_REG_21__SCAN_IN), .Y(n8352));
  OAI21X1 g7125(.A0(n7897), .A1(n6947), .B0(n8352), .Y(P2_U3573));
  NAND2X1 g7126(.A(n7897), .B(P2_DATAO_REG_22__SCAN_IN), .Y(n8354));
  OAI21X1 g7127(.A0(n7897), .A1(n6995), .B0(n8354), .Y(P2_U3574));
  NAND2X1 g7128(.A(n7897), .B(P2_DATAO_REG_23__SCAN_IN), .Y(n8356));
  OAI21X1 g7129(.A0(n7897), .A1(n7038), .B0(n8356), .Y(P2_U3575));
  NAND2X1 g7130(.A(n7897), .B(P2_DATAO_REG_24__SCAN_IN), .Y(n8358));
  OAI21X1 g7131(.A0(n7897), .A1(n7083), .B0(n8358), .Y(P2_U3576));
  NAND2X1 g7132(.A(n7897), .B(P2_DATAO_REG_25__SCAN_IN), .Y(n8360));
  OAI21X1 g7133(.A0(n7897), .A1(n7127), .B0(n8360), .Y(P2_U3577));
  NAND2X1 g7134(.A(n7897), .B(P2_DATAO_REG_26__SCAN_IN), .Y(n8362));
  OAI21X1 g7135(.A0(n7897), .A1(n7176), .B0(n8362), .Y(P2_U3578));
  NAND2X1 g7136(.A(n7897), .B(P2_DATAO_REG_27__SCAN_IN), .Y(n8364));
  OAI21X1 g7137(.A0(n7897), .A1(n7228), .B0(n8364), .Y(P2_U3579));
  NAND2X1 g7138(.A(n7897), .B(P2_DATAO_REG_28__SCAN_IN), .Y(n8366));
  OAI21X1 g7139(.A0(n7897), .A1(n7283), .B0(n8366), .Y(P2_U3580));
  NAND2X1 g7140(.A(n7897), .B(P2_DATAO_REG_29__SCAN_IN), .Y(n8368));
  OAI21X1 g7141(.A0(n7897), .A1(n7325), .B0(n8368), .Y(P2_U3581));
  NAND2X1 g7142(.A(n7897), .B(P2_DATAO_REG_30__SCAN_IN), .Y(n8370));
  OAI21X1 g7143(.A0(n7897), .A1(n7375), .B0(n8370), .Y(P2_U3582));
  NAND2X1 g7144(.A(n7897), .B(P2_DATAO_REG_31__SCAN_IN), .Y(n8372));
  OAI21X1 g7145(.A0(n7897), .A1(n7399), .B0(n8372), .Y(P2_U3583));
  NOR4X1  g7146(.A(n5853), .B(n5848), .C(n5850), .D(n5856), .Y(n8374));
  AOI21X1 g7147(.A0(n8374), .A1(n7755), .B0(n5735), .Y(n8375));
  NOR2X1  g7148(.A(n7750), .B(P2_U3152), .Y(n8376));
  OAI21X1 g7149(.A0(n5850), .A1(n5734), .B0(n8376), .Y(n8377));
  OAI21X1 g7150(.A0(n8377), .A1(n8375), .B0(P2_B_REG_SCAN_IN), .Y(n8378));
  INVX1   g7151(.A(n8374), .Y(n8379));
  NOR3X1  g7152(.A(n8379), .B(n7756), .C(n5750), .Y(n8380));
  AOI21X1 g7153(.A0(n5735), .A1(P2_STATE_REG_SCAN_IN), .B0(n8380), .Y(n8381));
  NOR3X1  g7154(.A(n5855), .B(n5853), .C(n5847), .Y(n8382));
  INVX1   g7155(.A(n7399), .Y(n8383));
  NOR3X1  g7156(.A(n5855), .B(n5848), .C(n5843), .Y(n8384));
  AOI21X1 g7157(.A0(n5855), .A1(n5735), .B0(n5848), .Y(n8385));
  OAI21X1 g7158(.A0(n5856), .A1(n5843), .B0(n8385), .Y(n8386));
  AOI21X1 g7159(.A0(n7368), .A1(n5856), .B0(n8386), .Y(n8387));
  INVX1   g7160(.A(n8387), .Y(n8388));
  AOI22X1 g7161(.A0(n8384), .A1(n7746), .B0(n8383), .B1(n8388), .Y(n8389));
  AOI22X1 g7162(.A0(n8384), .A1(n8383), .B0(n7746), .B1(n8388), .Y(n8390));
  INVX1   g7163(.A(n8390), .Y(n8391));
  XOR2X1  g7164(.A(n8391), .B(n8389), .Y(n8392));
  INVX1   g7165(.A(n8384), .Y(n8393));
  OAI22X1 g7166(.A0(n8393), .A1(n7375), .B0(n7394), .B1(n8387), .Y(n8394));
  OAI22X1 g7167(.A0(n7325), .A1(n8393), .B0(n7283), .B1(n5735), .Y(n8395));
  AOI21X1 g7168(.A0(n8388), .A1(n7333), .B0(n8395), .Y(n8396));
  AOI21X1 g7169(.A0(n8388), .A1(n7326), .B0(n5734), .Y(n8397));
  OAI21X1 g7170(.A0(n8393), .A1(n7386), .B0(n8397), .Y(n8398));
  NOR2X1  g7171(.A(n8398), .B(n8396), .Y(n8399));
  INVX1   g7172(.A(n7375), .Y(n8400));
  AOI22X1 g7173(.A0(n8384), .A1(n7407), .B0(n8400), .B1(n8388), .Y(n8401));
  AOI21X1 g7174(.A0(n8401), .A1(n8394), .B0(n8399), .Y(n8402));
  AOI22X1 g7175(.A0(n7346), .A1(n8384), .B0(n7242), .B1(n5734), .Y(n8403));
  OAI21X1 g7176(.A0(n8387), .A1(n7336), .B0(n8403), .Y(n8404));
  NAND3X1 g7177(.A(n8384), .B(n7056), .C(n7335), .Y(n8405));
  AOI21X1 g7178(.A0(n8388), .A1(n7346), .B0(n5734), .Y(n8406));
  NAND3X1 g7179(.A(n8406), .B(n8405), .C(n8404), .Y(n8407));
  NAND2X1 g7180(.A(n8388), .B(n7272), .Y(n8408));
  AOI22X1 g7181(.A0(n7242), .A1(n8384), .B0(n7183), .B1(n5734), .Y(n8409));
  AOI21X1 g7182(.A0(n8388), .A1(n7242), .B0(n5734), .Y(n8410));
  OAI21X1 g7183(.A0(n8393), .A1(n7243), .B0(n8410), .Y(n8411));
  AOI21X1 g7184(.A0(n8409), .A1(n8408), .B0(n8411), .Y(n8412));
  NAND3X1 g7185(.A(n8388), .B(n7056), .C(n7218), .Y(n8413));
  AOI22X1 g7186(.A0(n7183), .A1(n8384), .B0(n7152), .B1(n5734), .Y(n8414));
  AOI21X1 g7187(.A0(n8388), .A1(n7183), .B0(n5734), .Y(n8415));
  OAI21X1 g7188(.A0(n8393), .A1(n7219), .B0(n8415), .Y(n8416));
  AOI21X1 g7189(.A0(n8414), .A1(n8413), .B0(n8416), .Y(n8417));
  AOI21X1 g7190(.A0(n8388), .A1(n7152), .B0(n5734), .Y(n8418));
  INVX1   g7191(.A(n8418), .Y(n8419));
  AOI21X1 g7192(.A0(n8384), .A1(n7134), .B0(n8419), .Y(n8420));
  AOI22X1 g7193(.A0(n7152), .A1(n8384), .B0(n7090), .B1(n5734), .Y(n8421));
  OAI21X1 g7194(.A0(n8387), .A1(n7167), .B0(n8421), .Y(n8422));
  NOR4X1  g7195(.A(n8420), .B(n8417), .C(n8412), .D(n8422), .Y(n8423));
  NAND4X1 g7196(.A(n8407), .B(n8402), .C(n8392), .D(n8423), .Y(n8424));
  OAI21X1 g7197(.A0(n8387), .A1(n7243), .B0(n8409), .Y(n8425));
  INVX1   g7198(.A(n8411), .Y(n8426));
  NOR2X1  g7199(.A(n8426), .B(n8425), .Y(n8427));
  NAND4X1 g7200(.A(n8407), .B(n8402), .C(n8392), .D(n8427), .Y(n8428));
  NAND3X1 g7201(.A(n8416), .B(n8414), .C(n8413), .Y(n8429));
  AOI21X1 g7202(.A0(n8426), .A1(n8425), .B0(n8429), .Y(n8430));
  NAND4X1 g7203(.A(n8407), .B(n8402), .C(n8392), .D(n8430), .Y(n8431));
  NAND3X1 g7204(.A(n8431), .B(n8428), .C(n8424), .Y(n8432));
  NOR4X1  g7205(.A(n5848), .B(n5850), .C(n5735), .D(n5856), .Y(n8433));
  NOR2X1  g7206(.A(n8390), .B(n8389), .Y(n8434));
  AOI21X1 g7207(.A0(n8433), .A1(n8389), .B0(n8434), .Y(n8435));
  OAI21X1 g7208(.A0(n8433), .A1(n8391), .B0(n8435), .Y(n8436));
  NAND2X1 g7209(.A(n8398), .B(n8396), .Y(n8437));
  AOI21X1 g7210(.A0(n8401), .A1(n8394), .B0(n8437), .Y(n8438));
  NOR2X1  g7211(.A(n8401), .B(n8394), .Y(n8439));
  OAI21X1 g7212(.A0(n8439), .A1(n8438), .B0(n8392), .Y(n8440));
  NAND2X1 g7213(.A(n8422), .B(n8420), .Y(n8441));
  AOI21X1 g7214(.A0(n8388), .A1(n7090), .B0(n5734), .Y(n8442));
  OAI21X1 g7215(.A0(n8393), .A1(n7091), .B0(n8442), .Y(n8443));
  NAND3X1 g7216(.A(n8388), .B(n7056), .C(n5664), .Y(n8444));
  AOI22X1 g7217(.A0(n7090), .A1(n8384), .B0(n7053), .B1(n5734), .Y(n8445));
  NAND3X1 g7218(.A(n8445), .B(n8444), .C(n8443), .Y(n8446));
  AOI21X1 g7219(.A0(n8388), .A1(n7053), .B0(n5734), .Y(n8447));
  OAI21X1 g7220(.A0(n8393), .A1(n7057), .B0(n8447), .Y(n8448));
  AOI22X1 g7221(.A0(n7053), .A1(n8384), .B0(n7045), .B1(n5734), .Y(n8449));
  INVX1   g7222(.A(n8449), .Y(n8450));
  AOI21X1 g7223(.A0(n8388), .A1(n7049), .B0(n8450), .Y(n8451));
  NAND2X1 g7224(.A(n8451), .B(n8448), .Y(n8452));
  NAND2X1 g7225(.A(n8384), .B(n7002), .Y(n8453));
  AOI21X1 g7226(.A0(n8388), .A1(n7045), .B0(n5734), .Y(n8454));
  AOI22X1 g7227(.A0(n7045), .A1(n8384), .B0(n6946), .B1(n5734), .Y(n8455));
  OAI21X1 g7228(.A0(n8387), .A1(n7028), .B0(n8455), .Y(n8456));
  AOI21X1 g7229(.A0(n8454), .A1(n8453), .B0(n8456), .Y(n8457));
  AOI22X1 g7230(.A0(n6946), .A1(n8384), .B0(n6914), .B1(n5734), .Y(n8458));
  INVX1   g7231(.A(n8458), .Y(n8459));
  AOI21X1 g7232(.A0(n8388), .A1(n6954), .B0(n8459), .Y(n8460));
  AOI21X1 g7233(.A0(n8388), .A1(n6946), .B0(n5734), .Y(n8461));
  OAI21X1 g7234(.A0(n8393), .A1(n6984), .B0(n8461), .Y(n8462));
  AOI22X1 g7235(.A0(n6914), .A1(n8384), .B0(n6872), .B1(n5734), .Y(n8463));
  OAI21X1 g7236(.A0(n8387), .A1(n6939), .B0(n8463), .Y(n8464));
  INVX1   g7237(.A(n8464), .Y(n8465));
  AOI21X1 g7238(.A0(n8388), .A1(n6914), .B0(n5734), .Y(n8466));
  OAI21X1 g7239(.A0(n8393), .A1(n6939), .B0(n8466), .Y(n8467));
  OAI22X1 g7240(.A0(n8465), .A1(n8467), .B0(n8462), .B1(n8460), .Y(n8468));
  AOI22X1 g7241(.A0(n6872), .A1(n8384), .B0(n6818), .B1(n5734), .Y(n8469));
  OAI21X1 g7242(.A0(n8387), .A1(n6885), .B0(n8469), .Y(n8470));
  INVX1   g7243(.A(n8470), .Y(n8471));
  AOI21X1 g7244(.A0(n8388), .A1(n6872), .B0(n5734), .Y(n8472));
  OAI21X1 g7245(.A0(n8393), .A1(n6885), .B0(n8472), .Y(n8473));
  NAND2X1 g7246(.A(n8473), .B(n8471), .Y(n8474));
  NOR2X1  g7247(.A(n8474), .B(n8468), .Y(n8475));
  INVX1   g7248(.A(n8460), .Y(n8476));
  INVX1   g7249(.A(n8462), .Y(n8477));
  NAND2X1 g7250(.A(n8467), .B(n8465), .Y(n8478));
  AOI21X1 g7251(.A0(n8477), .A1(n8476), .B0(n8478), .Y(n8479));
  NOR2X1  g7252(.A(n8477), .B(n8476), .Y(n8480));
  NOR4X1  g7253(.A(n8479), .B(n8475), .C(n8457), .D(n8480), .Y(n8481));
  OAI22X1 g7254(.A0(n6799), .A1(n8393), .B0(n6740), .B1(n5735), .Y(n8482));
  AOI21X1 g7255(.A0(n8388), .A1(n6815), .B0(n8482), .Y(n8483));
  AOI21X1 g7256(.A0(n8388), .A1(n6818), .B0(n5734), .Y(n8484));
  OAI21X1 g7257(.A0(n8393), .A1(n6837), .B0(n8484), .Y(n8485));
  AOI22X1 g7258(.A0(n6747), .A1(n8384), .B0(n6689), .B1(n5734), .Y(n8486));
  OAI21X1 g7259(.A0(n8387), .A1(n6754), .B0(n8486), .Y(n8487));
  INVX1   g7260(.A(n8487), .Y(n8488));
  AOI21X1 g7261(.A0(n8388), .A1(n6747), .B0(n5734), .Y(n8489));
  OAI21X1 g7262(.A0(n8393), .A1(n6754), .B0(n8489), .Y(n8490));
  AOI22X1 g7263(.A0(n8488), .A1(n8490), .B0(n8485), .B1(n8483), .Y(n8491));
  INVX1   g7264(.A(n8491), .Y(n8492));
  OAI22X1 g7265(.A0(n6690), .A1(n8393), .B0(n6646), .B1(n5735), .Y(n8493));
  AOI21X1 g7266(.A0(n8388), .A1(n6704), .B0(n8493), .Y(n8494));
  AOI21X1 g7267(.A0(n8388), .A1(n6689), .B0(n5734), .Y(n8495));
  OAI21X1 g7268(.A0(n8393), .A1(n6731), .B0(n8495), .Y(n8496));
  NOR3X1  g7269(.A(n8496), .B(n8494), .C(n8492), .Y(n8497));
  NAND2X1 g7270(.A(n8485), .B(n8483), .Y(n8498));
  NOR2X1  g7271(.A(n8485), .B(n8483), .Y(n8499));
  NOR2X1  g7272(.A(n8490), .B(n8488), .Y(n8500));
  AOI21X1 g7273(.A0(n8500), .A1(n8498), .B0(n8499), .Y(n8501));
  OAI21X1 g7274(.A0(n8473), .A1(n8471), .B0(n8501), .Y(n8502));
  NOR3X1  g7275(.A(n8502), .B(n8497), .C(n8468), .Y(n8503));
  AOI21X1 g7276(.A0(n8388), .A1(n6660), .B0(n5734), .Y(n8504));
  OAI21X1 g7277(.A0(n8393), .A1(n6634), .B0(n8504), .Y(n8505));
  OAI22X1 g7278(.A0(n6597), .A1(n8393), .B0(n6546), .B1(n5735), .Y(n8506));
  AOI21X1 g7279(.A0(n8388), .A1(n6609), .B0(n8506), .Y(n8507));
  NAND2X1 g7280(.A(n8507), .B(n8505), .Y(n8508));
  AOI21X1 g7281(.A0(n8388), .A1(n6545), .B0(n5734), .Y(n8509));
  OAI21X1 g7282(.A0(n8393), .A1(n6559), .B0(n8509), .Y(n8510));
  INVX1   g7283(.A(n8510), .Y(n8511));
  AOI22X1 g7284(.A0(n6545), .A1(n8384), .B0(n6493), .B1(n5734), .Y(n8512));
  OAI21X1 g7285(.A0(n8387), .A1(n6559), .B0(n8512), .Y(n8513));
  AOI21X1 g7286(.A0(n8388), .A1(n6493), .B0(n5734), .Y(n8514));
  OAI21X1 g7287(.A0(n8393), .A1(n6528), .B0(n8514), .Y(n8515));
  OAI22X1 g7288(.A0(n6494), .A1(n8393), .B0(n6430), .B1(n5735), .Y(n8516));
  AOI21X1 g7289(.A0(n8388), .A1(n6506), .B0(n8516), .Y(n8517));
  AOI21X1 g7290(.A0(n8388), .A1(n6451), .B0(n5734), .Y(n8518));
  OAI21X1 g7291(.A0(n8393), .A1(n6453), .B0(n8518), .Y(n8519));
  AOI22X1 g7292(.A0(n6451), .A1(n8384), .B0(n6386), .B1(n5734), .Y(n8520));
  OAI21X1 g7293(.A0(n8387), .A1(n6453), .B0(n8520), .Y(n8521));
  INVX1   g7294(.A(n8521), .Y(n8522));
  AOI22X1 g7295(.A0(n8519), .A1(n8522), .B0(n8517), .B1(n8515), .Y(n8523));
  AOI22X1 g7296(.A0(n6354), .A1(n8384), .B0(n6292), .B1(n5734), .Y(n8524));
  OAI21X1 g7297(.A0(n8387), .A1(n6364), .B0(n8524), .Y(n8525));
  OAI21X1 g7298(.A0(n8387), .A1(n6327), .B0(n5735), .Y(n8526));
  AOI21X1 g7299(.A0(n8384), .A1(n6338), .B0(n8526), .Y(n8527));
  AOI22X1 g7300(.A0(n6292), .A1(n8384), .B0(n6234), .B1(n5734), .Y(n8528));
  INVX1   g7301(.A(n8528), .Y(n8529));
  AOI21X1 g7302(.A0(n8388), .A1(n6289), .B0(n8529), .Y(n8530));
  AOI21X1 g7303(.A0(n8388), .A1(n6292), .B0(n5734), .Y(n8531));
  OAI21X1 g7304(.A0(n8393), .A1(n6314), .B0(n8531), .Y(n8532));
  NOR2X1  g7305(.A(n8532), .B(n8530), .Y(n8533));
  AOI21X1 g7306(.A0(n8527), .A1(n8525), .B0(n8533), .Y(n8534));
  OAI22X1 g7307(.A0(n6172), .A1(n8393), .B0(n6121), .B1(n5735), .Y(n8535));
  AOI21X1 g7308(.A0(n8388), .A1(n6185), .B0(n8535), .Y(n8536));
  AOI21X1 g7309(.A0(n8388), .A1(n6231), .B0(n5734), .Y(n8537));
  OAI21X1 g7310(.A0(n8393), .A1(n6215), .B0(n8537), .Y(n8538));
  OAI22X1 g7311(.A0(n6121), .A1(n8393), .B0(n6092), .B1(n5735), .Y(n8539));
  AOI21X1 g7312(.A0(n8388), .A1(n6133), .B0(n8539), .Y(n8540));
  AOI21X1 g7313(.A0(n8388), .A1(n6146), .B0(n5734), .Y(n8541));
  OAI21X1 g7314(.A0(n8393), .A1(n6142), .B0(n8541), .Y(n8542));
  AOI22X1 g7315(.A0(n8540), .A1(n8542), .B0(n8538), .B1(n8536), .Y(n8543));
  AOI22X1 g7316(.A0(n6112), .A1(n8388), .B0(n6028), .B1(n5734), .Y(n8544));
  OAI21X1 g7317(.A0(n8393), .A1(n6092), .B0(n8544), .Y(n8545));
  OAI21X1 g7318(.A0(n8387), .A1(n6092), .B0(n5735), .Y(n8546));
  AOI21X1 g7319(.A0(n8384), .A1(n6112), .B0(n8546), .Y(n8547));
  NAND3X1 g7320(.A(n8547), .B(n8545), .C(n8543), .Y(n8548));
  NAND2X1 g7321(.A(n8538), .B(n8536), .Y(n8549));
  NOR2X1  g7322(.A(n8542), .B(n8540), .Y(n8550));
  OAI22X1 g7323(.A0(n6223), .A1(n8393), .B0(n6172), .B1(n5735), .Y(n8551));
  AOI21X1 g7324(.A0(n8388), .A1(n6239), .B0(n8551), .Y(n8552));
  AOI21X1 g7325(.A0(n8388), .A1(n6234), .B0(n5734), .Y(n8553));
  OAI21X1 g7326(.A0(n8393), .A1(n6264), .B0(n8553), .Y(n8554));
  OAI22X1 g7327(.A0(n8552), .A1(n8554), .B0(n8538), .B1(n8536), .Y(n8555));
  AOI21X1 g7328(.A0(n8550), .A1(n8549), .B0(n8555), .Y(n8556));
  AOI22X1 g7329(.A0(n8384), .A1(n6028), .B0(n6033), .B1(n8388), .Y(n8557));
  OAI21X1 g7330(.A0(n5974), .A1(n5735), .B0(n8557), .Y(n8558));
  OAI21X1 g7331(.A0(n8387), .A1(n6015), .B0(n5735), .Y(n8559));
  AOI21X1 g7332(.A0(n8384), .A1(n6033), .B0(n8559), .Y(n8560));
  NAND2X1 g7333(.A(n8560), .B(n8558), .Y(n8561));
  AOI22X1 g7334(.A0(n6046), .A1(n8388), .B0(n5922), .B1(n5734), .Y(n8562));
  OAI21X1 g7335(.A0(n8393), .A1(n5974), .B0(n8562), .Y(n8563));
  AOI21X1 g7336(.A0(n8384), .A1(n6046), .B0(n5734), .Y(n8564));
  OAI21X1 g7337(.A0(n8387), .A1(n5974), .B0(n8564), .Y(n8565));
  INVX1   g7338(.A(n8565), .Y(n8566));
  NOR2X1  g7339(.A(n8566), .B(n8563), .Y(n8567));
  OAI22X1 g7340(.A0(n8558), .A1(n8560), .B0(n8547), .B1(n8545), .Y(n8568));
  AOI21X1 g7341(.A0(n8567), .A1(n8561), .B0(n8568), .Y(n8569));
  NAND2X1 g7342(.A(n8569), .B(n8543), .Y(n8570));
  NAND4X1 g7343(.A(n8556), .B(n8548), .C(n8534), .D(n8570), .Y(n8571));
  NAND3X1 g7344(.A(n8554), .B(n8552), .C(n8534), .Y(n8572));
  NAND2X1 g7345(.A(n8532), .B(n8530), .Y(n8573));
  AOI21X1 g7346(.A0(n8527), .A1(n8525), .B0(n8573), .Y(n8574));
  AOI21X1 g7347(.A0(n8388), .A1(n6386), .B0(n5734), .Y(n8575));
  OAI21X1 g7348(.A0(n8393), .A1(n6419), .B0(n8575), .Y(n8576));
  INVX1   g7349(.A(n8576), .Y(n8577));
  AOI22X1 g7350(.A0(n6386), .A1(n8384), .B0(n6354), .B1(n5734), .Y(n8578));
  OAI21X1 g7351(.A0(n8387), .A1(n6419), .B0(n8578), .Y(n8579));
  OAI22X1 g7352(.A0(n8577), .A1(n8579), .B0(n8527), .B1(n8525), .Y(n8580));
  NOR2X1  g7353(.A(n8580), .B(n8574), .Y(n8581));
  NAND4X1 g7354(.A(n8572), .B(n8571), .C(n8523), .D(n8581), .Y(n8582));
  AOI22X1 g7355(.A0(n8563), .A1(n8566), .B0(n8560), .B1(n8558), .Y(n8583));
  NAND4X1 g7356(.A(n8556), .B(n8548), .C(n8534), .D(n8583), .Y(n8584));
  AOI21X1 g7357(.A0(n8384), .A1(n5939), .B0(n5734), .Y(n8585));
  OAI21X1 g7358(.A0(n8387), .A1(n5954), .B0(n8585), .Y(n8586));
  OAI22X1 g7359(.A0(n5967), .A1(n8387), .B0(n5897), .B1(n5735), .Y(n8587));
  AOI21X1 g7360(.A0(n8384), .A1(n5922), .B0(n8587), .Y(n8588));
  OAI22X1 g7361(.A0(n8393), .A1(n5897), .B0(n5923), .B1(n8387), .Y(n8589));
  AOI21X1 g7362(.A0(n8384), .A1(n5877), .B0(n5734), .Y(n8590));
  OAI21X1 g7363(.A0(n8387), .A1(n5897), .B0(n8590), .Y(n8591));
  NOR2X1  g7364(.A(n5848), .B(n5734), .Y(n8592));
  OAI21X1 g7365(.A0(n5855), .A1(n5843), .B0(n8592), .Y(n8593));
  NAND2X1 g7366(.A(n8593), .B(n8591), .Y(n8594));
  NOR2X1  g7367(.A(n8593), .B(n8591), .Y(n8595));
  AOI21X1 g7368(.A0(n8594), .A1(n8589), .B0(n8595), .Y(n8596));
  OAI21X1 g7369(.A0(n8588), .A1(n8586), .B0(n8596), .Y(n8597));
  NAND2X1 g7370(.A(n8588), .B(n8586), .Y(n8598));
  AOI21X1 g7371(.A0(n8598), .A1(n8597), .B0(n8584), .Y(n8599));
  NOR2X1  g7372(.A(n8599), .B(n8582), .Y(n8600));
  NAND3X1 g7373(.A(n8579), .B(n8577), .C(n8523), .Y(n8601));
  NAND2X1 g7374(.A(n8517), .B(n8515), .Y(n8602));
  NOR2X1  g7375(.A(n8522), .B(n8519), .Y(n8603));
  NAND2X1 g7376(.A(n8603), .B(n8602), .Y(n8604));
  NOR2X1  g7377(.A(n8517), .B(n8515), .Y(n8605));
  AOI21X1 g7378(.A0(n8513), .A1(n8511), .B0(n8605), .Y(n8606));
  NAND3X1 g7379(.A(n8606), .B(n8604), .C(n8601), .Y(n8607));
  OAI22X1 g7380(.A0(n8600), .A1(n8607), .B0(n8513), .B1(n8511), .Y(n8608));
  OAI21X1 g7381(.A0(n8507), .A1(n8505), .B0(n8608), .Y(n8609));
  AOI22X1 g7382(.A0(n6645), .A1(n8384), .B0(n6660), .B1(n5734), .Y(n8610));
  OAI21X1 g7383(.A0(n8387), .A1(n6678), .B0(n8610), .Y(n8611));
  INVX1   g7384(.A(n8611), .Y(n8612));
  AOI21X1 g7385(.A0(n8388), .A1(n6645), .B0(n5734), .Y(n8613));
  OAI21X1 g7386(.A0(n8393), .A1(n6678), .B0(n8613), .Y(n8614));
  NOR2X1  g7387(.A(n8614), .B(n8612), .Y(n8615));
  AOI21X1 g7388(.A0(n8609), .A1(n8508), .B0(n8615), .Y(n8616));
  AOI22X1 g7389(.A0(n8612), .A1(n8614), .B0(n8496), .B1(n8494), .Y(n8617));
  NAND2X1 g7390(.A(n8617), .B(n8491), .Y(n8618));
  OAI21X1 g7391(.A0(n8618), .A1(n8616), .B0(n8503), .Y(n8619));
  NAND4X1 g7392(.A(n8481), .B(n8452), .C(n8446), .D(n8619), .Y(n8620));
  NAND3X1 g7393(.A(n8384), .B(n7056), .C(n5664), .Y(n8621));
  NAND2X1 g7394(.A(n8445), .B(n8444), .Y(n8622));
  NAND3X1 g7395(.A(n8622), .B(n8442), .C(n8621), .Y(n8623));
  NAND3X1 g7396(.A(n8456), .B(n8454), .C(n8453), .Y(n8624));
  OAI21X1 g7397(.A0(n8451), .A1(n8448), .B0(n8624), .Y(n8625));
  NAND3X1 g7398(.A(n8625), .B(n8452), .C(n8446), .Y(n8626));
  NAND4X1 g7399(.A(n8623), .B(n8620), .C(n8441), .D(n8626), .Y(n8627));
  NOR3X1  g7400(.A(n8627), .B(n8417), .C(n8412), .Y(n8628));
  NAND4X1 g7401(.A(n8407), .B(n8402), .C(n8392), .D(n8628), .Y(n8629));
  AOI21X1 g7402(.A0(n8406), .A1(n8405), .B0(n8404), .Y(n8630));
  NAND3X1 g7403(.A(n8630), .B(n8402), .C(n8392), .Y(n8631));
  NAND4X1 g7404(.A(n8629), .B(n8440), .C(n8436), .D(n8631), .Y(n8632));
  OAI22X1 g7405(.A0(n8432), .A1(n8632), .B0(n8382), .B1(n5900), .Y(n8633));
  NOR2X1  g7406(.A(n5848), .B(n5843), .Y(n8634));
  AOI21X1 g7407(.A0(n5857), .A1(n5843), .B0(n8634), .Y(n8635));
  NOR4X1  g7408(.A(n8632), .B(n8432), .C(n5853), .D(n8635), .Y(n8636));
  NAND2X1 g7409(.A(n8383), .B(n8400), .Y(n8639));
  AOI22X1 g7410(.A0(n7325), .A1(n7333), .B0(n7407), .B1(n8639), .Y(n8640));
  NAND2X1 g7411(.A(n8383), .B(n7409), .Y(n8642));
  NAND4X1 g7412(.A(n8642), .B(n8640), .C(n7336), .D(n7346), .Y(n8645));
  NAND2X1 g7413(.A(n8639), .B(n7407), .Y(n8647));
  NAND4X1 g7414(.A(n8642), .B(n7326), .C(n7386), .D(n8647), .Y(n8648));
  NOR4X1  g7415(.A(n7399), .B(n7407), .C(n7375), .D(n7409), .Y(n8649));
  OAI21X1 g7416(.A0(n8383), .A1(n7409), .B0(n5843), .Y(n8650));
  NOR2X1  g7417(.A(n8650), .B(n8649), .Y(n8651));
  NAND3X1 g7418(.A(n8651), .B(n8648), .C(n8645), .Y(n8652));
  OAI22X1 g7419(.A0(n7346), .A1(n7336), .B0(n7243), .B1(n7242), .Y(n8655));
  AOI21X1 g7420(.A0(n8383), .A1(n7409), .B0(n8655), .Y(n8656));
  NAND4X1 g7421(.A(n8656), .B(n8640), .C(n7219), .D(n7183), .Y(n8659));
  NAND4X1 g7422(.A(n7242), .B(n8640), .C(n7243), .D(n8656), .Y(n8660));
  OAI21X1 g7423(.A0(n5867), .A1(n5643), .B0(n7045), .Y(n8671));
  OAI22X1 g7424(.A0(n6846), .A1(n6854), .B0(n6815), .B1(n6799), .Y(n8672));
  NAND2X1 g7425(.A(n6753), .B(n6740), .Y(n8673));
  NOR2X1  g7426(.A(n8673), .B(n8672), .Y(n8674));
  NAND2X1 g7427(.A(n6815), .B(n6799), .Y(n8679));
  OAI21X1 g7428(.A0(n8679), .A1(n6870), .B0(n6868), .Y(n8681));
  NOR3X1  g7429(.A(n8681), .B(n6921), .C(n8674), .Y(n8682));
  NOR2X1  g7430(.A(n6657), .B(n6646), .Y(n8683));
  AOI22X1 g7431(.A0(n6374), .A1(n6391), .B0(n6239), .B1(n6223), .Y(n8684));
  AOI22X1 g7432(.A0(n6327), .A1(n6338), .B0(n6289), .B1(n6275), .Y(n8685));
  NAND2X1 g7433(.A(n8685), .B(n8684), .Y(n8686));
  OAI22X1 g7434(.A0(n6231), .A1(n6215), .B0(n6142), .B1(n6146), .Y(n8687));
  NOR2X1  g7435(.A(n6077), .B(n6065), .Y(n8688));
  NOR3X1  g7436(.A(n8688), .B(n8687), .C(n8686), .Y(n8689));
  NAND3X1 g7437(.A(n6028), .B(n8689), .C(n6034), .Y(n8691));
  AOI22X1 g7438(.A0(n6146), .A1(n6142), .B0(n6077), .B1(n6065), .Y(n8692));
  AOI22X1 g7439(.A0(n6234), .A1(n6264), .B0(n6215), .B1(n6231), .Y(n8693));
  OAI21X1 g7440(.A0(n8692), .A1(n8687), .B0(n8693), .Y(n8694));
  NAND3X1 g7441(.A(n8694), .B(n8685), .C(n8684), .Y(n8695));
  OAI22X1 g7442(.A0(n6327), .A1(n6338), .B0(n6289), .B1(n6275), .Y(n8697));
  AOI22X1 g7443(.A0(n6374), .A1(n6391), .B0(n6338), .B1(n6327), .Y(n8698));
  OAI22X1 g7444(.A0(n6430), .A1(n6443), .B0(n6391), .B1(n6374), .Y(n8699));
  AOI21X1 g7445(.A0(n8698), .A1(n8697), .B0(n8699), .Y(n8700));
  NAND4X1 g7446(.A(n6611), .B(n8695), .C(n8691), .D(n8700), .Y(n8701));
  NAND3X1 g7447(.A(n6033), .B(n6027), .C(n6025), .Y(n8702));
  NOR3X1  g7448(.A(n5896), .B(n5892), .C(n5923), .Y(n8704));
  OAI21X1 g7449(.A0(n5954), .A1(n5939), .B0(n8704), .Y(n8705));
  AOI22X1 g7450(.A0(n5974), .A1(n6046), .B0(n5939), .B1(n5954), .Y(n8706));
  NAND4X1 g7451(.A(n8705), .B(n8702), .C(n8689), .D(n8706), .Y(n8707));
  NAND4X1 g7452(.A(n8702), .B(n8689), .C(n5990), .D(n5995), .Y(n8710));
  NAND2X1 g7453(.A(n8710), .B(n8707), .Y(n8711));
  OAI22X1 g7454(.A0(n6545), .A1(n6559), .B0(n6528), .B1(n6493), .Y(n8713));
  AOI21X1 g7455(.A0(n6450), .A1(n6611), .B0(n8713), .Y(n8714));
  OAI21X1 g7456(.A0(n8711), .A1(n8701), .B0(n8714), .Y(n8715));
  AOI22X1 g7457(.A0(n6660), .A1(n6634), .B0(n6559), .B1(n6545), .Y(n8716));
  AOI21X1 g7458(.A0(n8716), .A1(n8715), .B0(n6778), .Y(n8718));
  OAI22X1 g7459(.A0(n8718), .A1(n8683), .B0(n6731), .B1(n6689), .Y(n8720));
  OAI22X1 g7460(.A0(n6740), .A1(n6753), .B0(n6704), .B1(n6690), .Y(n8721));
  NOR2X1  g7461(.A(n8721), .B(n8672), .Y(n8722));
  AOI22X1 g7462(.A0(n8722), .A1(n8720), .B0(n6954), .B1(n6947), .Y(n8725));
  NAND2X1 g7463(.A(n8725), .B(n8682), .Y(n8726));
  OAI21X1 g7464(.A0(n5867), .A1(n5624), .B0(n6914), .Y(n8727));
  AOI21X1 g7465(.A0(n6947), .A1(n6954), .B0(n8727), .Y(n8728));
  AOI21X1 g7466(.A0(n6946), .A1(n6984), .B0(n8728), .Y(n8729));
  NAND3X1 g7467(.A(n8729), .B(n8726), .C(n8671), .Y(n8730));
  AOI22X1 g7468(.A0(n7038), .A1(n7049), .B0(n7002), .B1(n6995), .Y(n8731));
  AOI22X1 g7469(.A0(n8730), .A1(n8731), .B0(n7053), .B1(n7057), .Y(n8732));
  AOI21X1 g7470(.A0(n8732), .A1(n7238), .B0(n7136), .Y(n8733));
  AOI21X1 g7471(.A0(n8733), .A1(n7152), .B0(n7167), .Y(n8734));
  OAI22X1 g7472(.A0(n7152), .A1(n8733), .B0(n7183), .B1(n7219), .Y(n8735));
  NOR2X1  g7473(.A(n8735), .B(n8734), .Y(n8736));
  NAND3X1 g7474(.A(n8736), .B(n8656), .C(n8640), .Y(n8737));
  NAND3X1 g7475(.A(n8737), .B(n8660), .C(n8659), .Y(n8738));
  NOR2X1  g7476(.A(n8738), .B(n8652), .Y(n8739));
  NOR3X1  g7477(.A(n5856), .B(n5847), .C(n5843), .Y(n8740));
  OAI21X1 g7478(.A0(n5867), .A1(n5712), .B0(n7326), .Y(n8747));
  OAI21X1 g7479(.A0(n5867), .A1(n5704), .B0(n7346), .Y(n8750));
  NOR2X1  g7480(.A(n7228), .B(n7272), .Y(n8752));
  NAND3X1 g7481(.A(n7127), .B(n7056), .C(n7187), .Y(n8756));
  OAI21X1 g7482(.A0(n5867), .A1(n5673), .B0(n7152), .Y(n8758));
  NAND3X1 g7483(.A(n7083), .B(n7056), .C(n5664), .Y(n8762));
  NAND3X1 g7484(.A(n7038), .B(n7056), .C(n7055), .Y(n8764));
  OAI21X1 g7485(.A0(n5867), .A1(n5656), .B0(n7053), .Y(n8766));
  OAI21X1 g7486(.A0(n5867), .A1(n5633), .B0(n6946), .Y(n8774));
  NOR2X1  g7487(.A(n6028), .B(n6034), .Y(n8782));
  OAI22X1 g7488(.A0(n6065), .A1(n6077), .B0(n5967), .B1(n5922), .Y(n8786));
  NOR3X1  g7489(.A(n5958), .B(n5922), .C(n5923), .Y(n8789));
  NAND2X1 g7490(.A(n5939), .B(n5877), .Y(n8790));
  OAI22X1 g7491(.A0(n8790), .A1(n5958), .B0(n5990), .B1(n5995), .Y(n8792));
  NOR4X1  g7492(.A(n8789), .B(n8786), .C(n8782), .D(n8792), .Y(n8793));
  NAND2X1 g7493(.A(n5995), .B(n5990), .Y(n8795));
  NOR3X1  g7494(.A(n8795), .B(n8688), .C(n8782), .Y(n8796));
  NAND2X1 g7495(.A(n6028), .B(n6034), .Y(n8797));
  NOR2X1  g7496(.A(n8797), .B(n8688), .Y(n8798));
  NAND2X1 g7497(.A(n6231), .B(n6215), .Y(n8804));
  NAND3X1 g7498(.A(n8692), .B(n8804), .C(n6305), .Y(n8808));
  NOR4X1  g7499(.A(n8798), .B(n8796), .C(n8793), .D(n8808), .Y(n8809));
  NAND3X1 g7500(.A(n6189), .B(n8804), .C(n6305), .Y(n8811));
  NOR2X1  g7501(.A(n6231), .B(n6215), .Y(n8812));
  NAND2X1 g7502(.A(n8812), .B(n6305), .Y(n8813));
  NOR3X1  g7503(.A(n6341), .B(n6403), .C(n6448), .Y(n8823));
  NAND3X1 g7504(.A(n8823), .B(n8813), .C(n8811), .Y(n8824));
  NAND3X1 g7505(.A(n6292), .B(n6447), .C(n6314), .Y(n8827));
  NOR2X1  g7506(.A(n8827), .B(n6403), .Y(n8828));
  OAI21X1 g7507(.A0(n6546), .A1(n6558), .B0(n6454), .Y(n8834));
  OAI21X1 g7508(.A0(n6494), .A1(n6506), .B0(n6508), .Y(n8838));
  NOR3X1  g7509(.A(n8838), .B(n8834), .C(n8828), .Y(n8839));
  OAI21X1 g7510(.A0(n8824), .A1(n8809), .B0(n8839), .Y(n8840));
  NAND2X1 g7511(.A(n6494), .B(n6506), .Y(n8842));
  NOR2X1  g7512(.A(n8842), .B(n6565), .Y(n8843));
  NAND2X1 g7513(.A(n6646), .B(n6657), .Y(n8848));
  NOR3X1  g7514(.A(n6778), .B(n6564), .C(n8843), .Y(n8852));
  NAND2X1 g7515(.A(n6690), .B(n6704), .Y(n8854));
  NOR3X1  g7516(.A(n6451), .B(n6565), .C(n6453), .Y(n8855));
  OAI21X1 g7517(.A0(n6494), .A1(n6506), .B0(n8855), .Y(n8856));
  NAND4X1 g7518(.A(n8854), .B(n8852), .C(n8840), .D(n8856), .Y(n8857));
  NAND2X1 g7519(.A(n8683), .B(n8854), .Y(n8861));
  NAND4X1 g7520(.A(n6660), .B(n8848), .C(n6634), .D(n8854), .Y(n8862));
  NAND2X1 g7521(.A(n6689), .B(n6731), .Y(n8864));
  NAND3X1 g7522(.A(n8864), .B(n8862), .C(n8861), .Y(n8865));
  AOI21X1 g7523(.A0(n6747), .A1(n6754), .B0(n8865), .Y(n8866));
  OAI22X1 g7524(.A0(n6747), .A1(n6754), .B0(n6837), .B1(n6818), .Y(n8869));
  AOI21X1 g7525(.A0(n8866), .A1(n8857), .B0(n8869), .Y(n8870));
  AOI22X1 g7526(.A0(n6894), .A1(n6901), .B0(n6854), .B1(n6846), .Y(n8876));
  OAI21X1 g7527(.A0(n8672), .A1(n8870), .B0(n8876), .Y(n8877));
  NAND3X1 g7528(.A(n8877), .B(n8727), .C(n8774), .Y(n8878));
  NAND3X1 g7529(.A(n8878), .B(n7004), .C(n7047), .Y(n8879));
  NAND3X1 g7530(.A(n8879), .B(n8671), .C(n8766), .Y(n8880));
  NAND3X1 g7531(.A(n8880), .B(n8764), .C(n8762), .Y(n8881));
  NAND3X1 g7532(.A(n8881), .B(n7238), .C(n8758), .Y(n8882));
  NAND3X1 g7533(.A(n8882), .B(n8756), .C(n7241), .Y(n8883));
  OAI21X1 g7534(.A0(n7176), .A1(n7184), .B0(n8883), .Y(n8884));
  AOI22X1 g7535(.A0(n7283), .A1(n7290), .B0(n7272), .B1(n7228), .Y(n8885));
  OAI21X1 g7536(.A0(n8884), .A1(n8752), .B0(n8885), .Y(n8886));
  NAND3X1 g7537(.A(n8886), .B(n8750), .C(n8747), .Y(n8887));
  NAND2X1 g7538(.A(n7325), .B(n7333), .Y(n8888));
  NAND4X1 g7539(.A(n8887), .B(n8642), .C(n7394), .D(n8888), .Y(n8889));
  NAND2X1 g7540(.A(n7399), .B(n7746), .Y(n8890));
  OAI22X1 g7541(.A0(n8639), .A1(n8740), .B0(n7375), .B1(n5847), .Y(n8891));
  INVX1   g7542(.A(n8891), .Y(n8892));
  AOI21X1 g7543(.A0(n8383), .A1(n7409), .B0(n8892), .Y(n8893));
  NAND3X1 g7544(.A(n8893), .B(n8888), .C(n8887), .Y(n8894));
  NAND2X1 g7545(.A(n8893), .B(n7394), .Y(n8895));
  NAND4X1 g7546(.A(n8894), .B(n8890), .C(n8889), .D(n8895), .Y(n8896));
  OAI21X1 g7547(.A0(n8896), .A1(n5843), .B0(n5901), .Y(n8897));
  NOR2X1  g7548(.A(n8897), .B(n8739), .Y(n8898));
  AOI21X1 g7549(.A0(n5924), .A1(n5855), .B0(n5908), .Y(n8899));
  XOR2X1  g7550(.A(n7394), .B(n7375), .Y(n8900));
  XOR2X1  g7551(.A(n7746), .B(n7399), .Y(n8901));
  XOR2X1  g7552(.A(n7243), .B(n7228), .Y(n8904));
  XOR2X1  g7553(.A(n6954), .B(n6946), .Y(n8908));
  XOR2X1  g7554(.A(n6901), .B(n6914), .Y(n8909));
  OAI22X1 g7555(.A0(n6080), .A1(n6082), .B0(n5993), .B1(n5991), .Y(n8911));
  XOR2X1  g7556(.A(n5897), .B(n5923), .Y(n8912));
  NOR4X1  g7557(.A(n8911), .B(n6093), .C(n5940), .D(n8912), .Y(n8913));
  NAND4X1 g7558(.A(n6134), .B(n8913), .C(n6186), .D(n6244), .Y(n8916));
  NOR2X1  g7559(.A(n6355), .B(n6293), .Y(n8918));
  NAND3X1 g7560(.A(n8918), .B(n6396), .C(n6444), .Y(n8919));
  NAND4X1 g7561(.A(n6610), .B(n6574), .C(n6507), .D(n6658), .Y(n8923));
  NOR4X1  g7562(.A(n8919), .B(n8916), .C(n6716), .D(n8923), .Y(n8924));
  NAND3X1 g7563(.A(n8924), .B(n6772), .C(n6816), .Y(n8925));
  NOR4X1  g7564(.A(n8909), .B(n8908), .C(n6873), .D(n8925), .Y(n8926));
  NAND4X1 g7565(.A(n7003), .B(n7050), .C(n7092), .D(n8926), .Y(n8927));
  NOR4X1  g7566(.A(n7185), .B(n8904), .C(n7153), .D(n8927), .Y(n8928));
  NAND4X1 g7567(.A(n7291), .B(n7334), .C(n8901), .D(n8928), .Y(n8929));
  NOR2X1  g7568(.A(n8929), .B(n8900), .Y(n8930));
  NOR2X1  g7569(.A(n5855), .B(n5847), .Y(n8931));
  NAND2X1 g7570(.A(n8931), .B(n5853), .Y(n8932));
  OAI21X1 g7571(.A0(n8930), .A1(n8932), .B0(n8378), .Y(n8933));
  AOI21X1 g7572(.A0(n8930), .A1(n5927), .B0(n8933), .Y(n8934));
  OAI21X1 g7573(.A0(n8899), .A1(n8896), .B0(n8934), .Y(n8935));
  NOR3X1  g7574(.A(n8935), .B(n8898), .C(n8636), .Y(n8936));
  AOI22X1 g7575(.A0(n8633), .A1(n8936), .B0(n8381), .B1(n8378), .Y(P2_U3244));
  NOR4X1  g7576(.A(n5853), .B(n5847), .C(n5843), .D(n5856), .Y(n8938));
  NOR2X1  g7577(.A(n8938), .B(n6597), .Y(n8939));
  INVX1   g7578(.A(n8939), .Y(n8940));
  NOR2X1  g7579(.A(n5852), .B(n5848), .Y(n8941));
  NOR3X1  g7580(.A(n8941), .B(n8931), .C(n5926), .Y(n8942));
  XOR2X1  g7581(.A(n8942), .B(n6609), .Y(n8943));
  NOR2X1  g7582(.A(n8943), .B(n8940), .Y(n8944));
  INVX1   g7583(.A(n8944), .Y(n8945));
  NAND2X1 g7584(.A(n8943), .B(n8940), .Y(n8946));
  INVX1   g7585(.A(n8946), .Y(n8947));
  XOR2X1  g7586(.A(n8942), .B(n6558), .Y(n8948));
  AOI21X1 g7587(.A0(n6544), .A1(n6538), .B0(n8938), .Y(n8949));
  INVX1   g7588(.A(n8949), .Y(n8950));
  XOR2X1  g7589(.A(n8942), .B(n6443), .Y(n8951));
  NOR3X1  g7590(.A(n8951), .B(n8938), .C(n6430), .Y(n8952));
  INVX1   g7591(.A(n8938), .Y(n8953));
  NAND2X1 g7592(.A(n8953), .B(n6493), .Y(n8954));
  XOR2X1  g7593(.A(n8942), .B(n6506), .Y(n8955));
  AOI22X1 g7594(.A0(n8954), .A1(n8955), .B0(n8950), .B1(n8948), .Y(n8956));
  NAND2X1 g7595(.A(n8956), .B(n8952), .Y(n8957));
  INVX1   g7596(.A(n8948), .Y(n8958));
  NOR2X1  g7597(.A(n8955), .B(n8954), .Y(n8959));
  AOI21X1 g7598(.A0(n8949), .A1(n8958), .B0(n8959), .Y(n8960));
  AOI22X1 g7599(.A0(n8957), .A1(n8960), .B0(n8950), .B1(n8948), .Y(n8961));
  AOI21X1 g7600(.A0(n6385), .A1(n6383), .B0(n8938), .Y(n8962));
  INVX1   g7601(.A(n8962), .Y(n8963));
  XOR2X1  g7602(.A(n8942), .B(n6391), .Y(n8964));
  INVX1   g7603(.A(n8964), .Y(n8965));
  NOR2X1  g7604(.A(n8938), .B(n6327), .Y(n8966));
  INVX1   g7605(.A(n8966), .Y(n8967));
  OAI21X1 g7606(.A0(n6274), .A1(n6268), .B0(n8953), .Y(n8968));
  XOR2X1  g7607(.A(n8942), .B(n6289), .Y(n8969));
  NOR2X1  g7608(.A(n8969), .B(n8968), .Y(n8970));
  NAND2X1 g7609(.A(n8969), .B(n8968), .Y(n8971));
  OAI21X1 g7610(.A0(n6171), .A1(n6165), .B0(n8953), .Y(n8972));
  XOR2X1  g7611(.A(n8942), .B(n6185), .Y(n8973));
  NOR2X1  g7612(.A(n8938), .B(n6223), .Y(n8974));
  INVX1   g7613(.A(n8974), .Y(n8975));
  XOR2X1  g7614(.A(n8942), .B(n6239), .Y(n8976));
  AOI22X1 g7615(.A0(n8975), .A1(n8976), .B0(n8973), .B1(n8972), .Y(n8977));
  OAI21X1 g7616(.A0(n6120), .A1(n6116), .B0(n8953), .Y(n8978));
  XOR2X1  g7617(.A(n8942), .B(n6133), .Y(n8979));
  NOR2X1  g7618(.A(n8979), .B(n8978), .Y(n8980));
  AOI21X1 g7619(.A0(n6064), .A1(n6061), .B0(n8938), .Y(n8981));
  AOI21X1 g7620(.A0(n5985), .A1(n5984), .B0(n8938), .Y(n8982));
  XOR2X1  g7621(.A(n8942), .B(n5990), .Y(n8983));
  OAI21X1 g7622(.A0(n6014), .A1(n6012), .B0(n8953), .Y(n8984));
  INVX1   g7623(.A(n8984), .Y(n8985));
  XOR2X1  g7624(.A(n8942), .B(n6033), .Y(n8986));
  INVX1   g7625(.A(n8986), .Y(n8987));
  OAI22X1 g7626(.A0(n8985), .A1(n8987), .B0(n8983), .B1(n8982), .Y(n8988));
  OAI21X1 g7627(.A0(n5953), .A1(n5950), .B0(n8953), .Y(n8989));
  XOR2X1  g7628(.A(n8942), .B(n5939), .Y(n8990));
  NOR2X1  g7629(.A(n8990), .B(n8989), .Y(n8991));
  NAND2X1 g7630(.A(n8990), .B(n8989), .Y(n8992));
  NOR2X1  g7631(.A(n8941), .B(n5926), .Y(n8993));
  OAI21X1 g7632(.A0(n5855), .A1(n5847), .B0(n8993), .Y(n8994));
  AOI21X1 g7633(.A0(n5946), .A1(n5945), .B0(n8938), .Y(n8995));
  OAI21X1 g7634(.A0(n8994), .A1(n5877), .B0(n8995), .Y(n8996));
  OAI21X1 g7635(.A0(n8942), .A1(n5877), .B0(n8996), .Y(n8997));
  AOI21X1 g7636(.A0(n8997), .A1(n8992), .B0(n8991), .Y(n8998));
  XOR2X1  g7637(.A(n8942), .B(n6046), .Y(n8999));
  NOR3X1  g7638(.A(n8999), .B(n8938), .C(n5974), .Y(n9000));
  NAND2X1 g7639(.A(n8983), .B(n8982), .Y(n9001));
  AOI21X1 g7640(.A0(n9001), .A1(n8984), .B0(n8986), .Y(n9002));
  AOI21X1 g7641(.A0(n9000), .A1(n8985), .B0(n9002), .Y(n9003));
  OAI21X1 g7642(.A0(n8998), .A1(n8988), .B0(n9003), .Y(n9004));
  NAND2X1 g7643(.A(n9004), .B(n8981), .Y(n9005));
  XOR2X1  g7644(.A(n8942), .B(n6112), .Y(n9006));
  INVX1   g7645(.A(n9006), .Y(n9007));
  OAI21X1 g7646(.A0(n9004), .A1(n8981), .B0(n9007), .Y(n9008));
  AOI22X1 g7647(.A0(n9005), .A1(n9008), .B0(n8979), .B1(n8978), .Y(n9009));
  OAI21X1 g7648(.A0(n9009), .A1(n8980), .B0(n8977), .Y(n9010));
  NOR2X1  g7649(.A(n8973), .B(n8972), .Y(n9011));
  INVX1   g7650(.A(n9011), .Y(n9012));
  AOI21X1 g7651(.A0(n9012), .A1(n8975), .B0(n8976), .Y(n9013));
  AOI21X1 g7652(.A0(n9011), .A1(n8974), .B0(n9013), .Y(n9014));
  NAND2X1 g7653(.A(n9014), .B(n9010), .Y(n9015));
  AOI21X1 g7654(.A0(n9015), .A1(n8971), .B0(n8970), .Y(n9016));
  NOR2X1  g7655(.A(n9016), .B(n8967), .Y(n9017));
  XOR2X1  g7656(.A(n8942), .B(n6338), .Y(n9018));
  AOI21X1 g7657(.A0(n9016), .A1(n8967), .B0(n9018), .Y(n9019));
  OAI22X1 g7658(.A0(n9017), .A1(n9019), .B0(n8965), .B1(n8962), .Y(n9020));
  OAI21X1 g7659(.A0(n8964), .A1(n8963), .B0(n9020), .Y(n9021));
  OAI21X1 g7660(.A0(n8938), .A1(n6430), .B0(n8951), .Y(n9022));
  NAND2X1 g7661(.A(n9022), .B(n8956), .Y(n9023));
  INVX1   g7662(.A(n9023), .Y(n9024));
  AOI21X1 g7663(.A0(n9024), .A1(n9021), .B0(n8961), .Y(n9025));
  OAI21X1 g7664(.A0(n9025), .A1(n8947), .B0(n8945), .Y(n9026));
  XOR2X1  g7665(.A(n8942), .B(n6657), .Y(n9027));
  NOR2X1  g7666(.A(n8938), .B(n6646), .Y(n9028));
  XOR2X1  g7667(.A(n9028), .B(n9027), .Y(n9029));
  XOR2X1  g7668(.A(n9029), .B(n9026), .Y(n9030));
  NOR3X1  g7669(.A(n5861), .B(n5840), .C(n7483), .Y(n9031));
  INVX1   g7670(.A(n9031), .Y(n9032));
  NAND2X1 g7671(.A(n8931), .B(n5843), .Y(n9033));
  NAND2X1 g7672(.A(n5847), .B(n5850), .Y(n9034));
  AOI22X1 g7673(.A0(n5903), .A1(n5848), .B0(n5855), .B1(n5924), .Y(n9035));
  NAND4X1 g7674(.A(n9034), .B(n9033), .C(n6097), .D(n9035), .Y(n9036));
  INVX1   g7675(.A(n9036), .Y(n9037));
  NOR3X1  g7676(.A(n9037), .B(n9032), .C(n5750), .Y(n9038));
  INVX1   g7677(.A(n9038), .Y(n9039));
  NOR4X1  g7678(.A(n5742), .B(n5735), .C(P2_U3152), .D(n7494), .Y(n9040));
  NOR2X1  g7679(.A(n9037), .B(n9031), .Y(n9041));
  NOR4X1  g7680(.A(n7750), .B(n7485), .C(n5735), .D(n9041), .Y(n9042));
  NOR2X1  g7681(.A(n9042), .B(P2_U3152), .Y(n9043));
  AOI21X1 g7682(.A0(n9040), .A1(n9032), .B0(n9043), .Y(n9044));
  INVX1   g7683(.A(n9044), .Y(n9045));
  NOR2X1  g7684(.A(n8379), .B(n5750), .Y(n9046));
  INVX1   g7685(.A(n9046), .Y(n9047));
  NOR4X1  g7686(.A(n5861), .B(n5840), .C(n7483), .D(n5866), .Y(n9048));
  NOR4X1  g7687(.A(n5861), .B(n5840), .C(n7483), .D(n5871), .Y(n9049));
  INVX1   g7688(.A(n9049), .Y(n9050));
  OAI22X1 g7689(.A0(n9031), .A1(n6642), .B0(n6597), .B1(n9050), .Y(n9051));
  AOI21X1 g7690(.A0(n9048), .A1(n6689), .B0(n9051), .Y(n9052));
  AOI22X1 g7691(.A0(n9031), .A1(n9040), .B0(n7481), .B1(n5743), .Y(n9053));
  AOI22X1 g7692(.A0(n6657), .A1(n9145), .B0(P2_REG3_REG_15__SCAN_IN), .B1(P2_U3152), .Y(n9055));
  OAI21X1 g7693(.A0(n9052), .A1(n9047), .B0(n9055), .Y(n9056));
  AOI21X1 g7694(.A0(n9045), .A1(n6643), .B0(n9056), .Y(n9057));
  OAI21X1 g7695(.A0(n9039), .A1(n9030), .B0(n9057), .Y(P2_U3243));
  XOR2X1  g7696(.A(n8942), .B(n7134), .Y(n9059));
  INVX1   g7697(.A(n9059), .Y(n9060));
  NOR2X1  g7698(.A(n8938), .B(n7127), .Y(n9061));
  NOR2X1  g7699(.A(n9061), .B(n9060), .Y(n9062));
  NAND2X1 g7700(.A(n8953), .B(n7090), .Y(n9063));
  XOR2X1  g7701(.A(n8994), .B(n7091), .Y(n9064));
  NOR2X1  g7702(.A(n9064), .B(n9063), .Y(n9065));
  NAND2X1 g7703(.A(n9064), .B(n9063), .Y(n9066));
  NOR2X1  g7704(.A(n8938), .B(n7038), .Y(n9067));
  INVX1   g7705(.A(n9067), .Y(n9068));
  XOR2X1  g7706(.A(n8942), .B(n7049), .Y(n9069));
  NOR2X1  g7707(.A(n9069), .B(n9068), .Y(n9070));
  INVX1   g7708(.A(n9070), .Y(n9071));
  NAND2X1 g7709(.A(n9069), .B(n9068), .Y(n9072));
  INVX1   g7710(.A(n9072), .Y(n9073));
  XOR2X1  g7711(.A(n8942), .B(n7002), .Y(n9074));
  NOR3X1  g7712(.A(n9074), .B(n8938), .C(n6995), .Y(n9075));
  NOR2X1  g7713(.A(n8938), .B(n6995), .Y(n9076));
  INVX1   g7714(.A(n9074), .Y(n9077));
  NOR2X1  g7715(.A(n9077), .B(n9076), .Y(n9078));
  INVX1   g7716(.A(n9078), .Y(n9079));
  XOR2X1  g7717(.A(n8942), .B(n6954), .Y(n9080));
  INVX1   g7718(.A(n9080), .Y(n9081));
  NOR2X1  g7719(.A(n8938), .B(n6947), .Y(n9082));
  NOR2X1  g7720(.A(n8938), .B(n6846), .Y(n9083));
  INVX1   g7721(.A(n9083), .Y(n9084));
  XOR2X1  g7722(.A(n8942), .B(n6854), .Y(n9085));
  NOR2X1  g7723(.A(n9085), .B(n9084), .Y(n9086));
  INVX1   g7724(.A(n9086), .Y(n9087));
  INVX1   g7725(.A(n9082), .Y(n9088));
  OAI21X1 g7726(.A0(n6893), .A1(n6889), .B0(n8953), .Y(n9089));
  XOR2X1  g7727(.A(n8942), .B(n6901), .Y(n9090));
  AOI22X1 g7728(.A0(n9089), .A1(n9090), .B0(n9088), .B1(n9080), .Y(n9091));
  INVX1   g7729(.A(n9091), .Y(n9092));
  NOR2X1  g7730(.A(n9090), .B(n9089), .Y(n9093));
  AOI21X1 g7731(.A0(n9082), .A1(n9081), .B0(n9093), .Y(n9094));
  OAI21X1 g7732(.A0(n9092), .A1(n9087), .B0(n9094), .Y(n9095));
  OAI21X1 g7733(.A0(n9082), .A1(n9081), .B0(n9095), .Y(n9096));
  XOR2X1  g7734(.A(n8942), .B(n6815), .Y(n9097));
  NOR3X1  g7735(.A(n9097), .B(n8938), .C(n6799), .Y(n9098));
  NOR2X1  g7736(.A(n8938), .B(n6799), .Y(n9099));
  INVX1   g7737(.A(n9097), .Y(n9100));
  NOR2X1  g7738(.A(n9100), .B(n9099), .Y(n9101));
  INVX1   g7739(.A(n9101), .Y(n9102));
  NAND2X1 g7740(.A(n8953), .B(n6689), .Y(n9103));
  XOR2X1  g7741(.A(n8942), .B(n6704), .Y(n9104));
  NOR2X1  g7742(.A(n6737), .B(n6735), .Y(n9105));
  AOI21X1 g7743(.A0(n6738), .A1(n9105), .B0(n8938), .Y(n9106));
  INVX1   g7744(.A(n9106), .Y(n9107));
  XOR2X1  g7745(.A(n8942), .B(n6753), .Y(n9108));
  AOI22X1 g7746(.A0(n9107), .A1(n9108), .B0(n9104), .B1(n9103), .Y(n9109));
  INVX1   g7747(.A(n9109), .Y(n9110));
  NOR3X1  g7748(.A(n9027), .B(n8938), .C(n6646), .Y(n9111));
  INVX1   g7749(.A(n9027), .Y(n9112));
  NOR2X1  g7750(.A(n9028), .B(n9112), .Y(n9113));
  INVX1   g7751(.A(n9113), .Y(n9114));
  AOI21X1 g7752(.A0(n9114), .A1(n9026), .B0(n9111), .Y(n9115));
  NOR2X1  g7753(.A(n9104), .B(n9103), .Y(n9116));
  INVX1   g7754(.A(n9116), .Y(n9117));
  AOI21X1 g7755(.A0(n9117), .A1(n9107), .B0(n9108), .Y(n9118));
  AOI21X1 g7756(.A0(n9116), .A1(n9106), .B0(n9118), .Y(n9119));
  OAI21X1 g7757(.A0(n9115), .A1(n9110), .B0(n9119), .Y(n9120));
  AOI21X1 g7758(.A0(n9120), .A1(n9102), .B0(n9098), .Y(n9121));
  AOI21X1 g7759(.A0(n9085), .A1(n9084), .B0(n9092), .Y(n9122));
  INVX1   g7760(.A(n9122), .Y(n9123));
  OAI21X1 g7761(.A0(n9123), .A1(n9121), .B0(n9096), .Y(n9124));
  AOI21X1 g7762(.A0(n9124), .A1(n9079), .B0(n9075), .Y(n9125));
  OAI21X1 g7763(.A0(n9125), .A1(n9073), .B0(n9071), .Y(n9126));
  AOI21X1 g7764(.A0(n9126), .A1(n9066), .B0(n9065), .Y(n9127));
  NOR2X1  g7765(.A(n9127), .B(n9062), .Y(n9128));
  NOR2X1  g7766(.A(n8938), .B(n7176), .Y(n9129));
  INVX1   g7767(.A(n9129), .Y(n9130));
  XOR2X1  g7768(.A(n8942), .B(n7184), .Y(n9131));
  INVX1   g7769(.A(n9131), .Y(n9132));
  AOI22X1 g7770(.A0(n9130), .A1(n9132), .B0(n9061), .B1(n9060), .Y(n9133));
  OAI21X1 g7771(.A0(n9132), .A1(n9130), .B0(n9133), .Y(n9134));
  NOR2X1  g7772(.A(n9134), .B(n9128), .Y(n9135));
  INVX1   g7773(.A(n9065), .Y(n9136));
  NAND2X1 g7774(.A(n9061), .B(n9060), .Y(n9137));
  NAND2X1 g7775(.A(n9137), .B(n9136), .Y(n9138));
  AOI21X1 g7776(.A0(n9126), .A1(n9066), .B0(n9138), .Y(n9139));
  OAI22X1 g7777(.A0(n9129), .A1(n9132), .B0(n9061), .B1(n9060), .Y(n9140));
  INVX1   g7778(.A(n9140), .Y(n9141));
  OAI21X1 g7779(.A0(n9131), .A1(n9130), .B0(n9141), .Y(n9142));
  OAI21X1 g7780(.A0(n9142), .A1(n9139), .B0(n9038), .Y(n9143));
  NAND4X1 g7781(.A(n7415), .B(n5841), .C(n5837), .D(n7553), .Y(n9144));
  AOI21X1 g7782(.A0(n9144), .A1(n7482), .B0(n5750), .Y(n9145));
  OAI21X1 g7783(.A0(n9031), .A1(n7494), .B0(n9042), .Y(n9146));
  INVX1   g7784(.A(n9048), .Y(n9148));
  AOI22X1 g7785(.A0(n9032), .A1(n7171), .B0(n7152), .B1(n9049), .Y(n9149));
  OAI21X1 g7786(.A0(n9148), .A1(n7228), .B0(n9149), .Y(n9150));
  AOI22X1 g7787(.A0(n9046), .A1(n9150), .B0(P2_REG3_REG_26__SCAN_IN), .B1(P2_U3152), .Y(n9151));
  OAI21X1 g7788(.A0(n9044), .A1(n7170), .B0(n9151), .Y(n9152));
  AOI21X1 g7789(.A0(n9145), .A1(n7184), .B0(n9152), .Y(n9153));
  OAI21X1 g7790(.A0(n9143), .A1(n9135), .B0(n9153), .Y(P2_U3242));
  NOR2X1  g7791(.A(n9009), .B(n8980), .Y(n9155));
  XOR2X1  g7792(.A(n8973), .B(n8972), .Y(n9156));
  NOR2X1  g7793(.A(n9156), .B(n9155), .Y(n9158));
  AOI21X1 g7794(.A0(n9156), .A1(n9155), .B0(n9158), .Y(n9159));
  NOR2X1  g7795(.A(n9148), .B(n6223), .Y(n9160));
  OAI22X1 g7796(.A0(n9031), .A1(n6168), .B0(n6121), .B1(n9050), .Y(n9161));
  OAI21X1 g7797(.A0(n9161), .A1(n9160), .B0(n9046), .Y(n9162));
  AOI22X1 g7798(.A0(n6185), .A1(n9145), .B0(P2_REG3_REG_6__SCAN_IN), .B1(P2_U3152), .Y(n9163));
  NAND2X1 g7799(.A(n9163), .B(n9162), .Y(n9164));
  AOI21X1 g7800(.A0(n9045), .A1(n6169), .B0(n9164), .Y(n9165));
  OAI21X1 g7801(.A0(n9159), .A1(n9039), .B0(n9165), .Y(P2_U3241));
  XOR2X1  g7802(.A(n9097), .B(n9099), .Y(n9167));
  XOR2X1  g7803(.A(n9167), .B(n9120), .Y(n9168));
  AOI22X1 g7804(.A0(n9032), .A1(n6792), .B0(n6747), .B1(n9049), .Y(n9169));
  OAI21X1 g7805(.A0(n9148), .A1(n6846), .B0(n9169), .Y(n9170));
  AOI22X1 g7806(.A0(n9046), .A1(n9170), .B0(P2_REG3_REG_18__SCAN_IN), .B1(P2_U3152), .Y(n9171));
  OAI21X1 g7807(.A0(n9044), .A1(n6793), .B0(n9171), .Y(n9172));
  AOI21X1 g7808(.A0(n9145), .A1(n6815), .B0(n9172), .Y(n9173));
  OAI21X1 g7809(.A0(n9168), .A1(n9039), .B0(n9173), .Y(P2_U3240));
  NAND2X1 g7810(.A(n9045), .B(P2_REG3_REG_2__SCAN_IN), .Y(n9175));
  NOR2X1  g7811(.A(n9148), .B(n6015), .Y(n9176));
  OAI22X1 g7812(.A0(n9031), .A1(n5971), .B0(n5954), .B1(n9050), .Y(n9177));
  OAI21X1 g7813(.A0(n9177), .A1(n9176), .B0(n9046), .Y(n9178));
  NAND2X1 g7814(.A(n9145), .B(n6046), .Y(n9179));
  XOR2X1  g7815(.A(n8983), .B(n8982), .Y(n9180));
  NAND2X1 g7816(.A(n9180), .B(n8998), .Y(n9181));
  OAI21X1 g7817(.A0(n9180), .A1(n8998), .B0(n9181), .Y(n9183));
  AOI22X1 g7818(.A0(n9038), .A1(n9183), .B0(P2_REG3_REG_2__SCAN_IN), .B1(P2_U3152), .Y(n9184));
  NAND4X1 g7819(.A(n9179), .B(n9178), .C(n9175), .D(n9184), .Y(P2_U3239));
  NOR2X1  g7820(.A(n8938), .B(n6430), .Y(n9186));
  XOR2X1  g7821(.A(n8951), .B(n9186), .Y(n9187));
  NOR2X1  g7822(.A(n9187), .B(n9021), .Y(n9188));
  AOI21X1 g7823(.A0(n9187), .A1(n9021), .B0(n9188), .Y(n9190));
  OAI22X1 g7824(.A0(n9031), .A1(n6428), .B0(n6374), .B1(n9050), .Y(n9191));
  AOI21X1 g7825(.A0(n9048), .A1(n6493), .B0(n9191), .Y(n9192));
  AOI22X1 g7826(.A0(n6443), .A1(n9145), .B0(P2_REG3_REG_11__SCAN_IN), .B1(P2_U3152), .Y(n9193));
  OAI21X1 g7827(.A0(n9192), .A1(n9047), .B0(n9193), .Y(n9194));
  AOI21X1 g7828(.A0(n9045), .A1(n7580), .B0(n9194), .Y(n9195));
  OAI21X1 g7829(.A0(n9190), .A1(n9039), .B0(n9195), .Y(P2_U3238));
  XOR2X1  g7830(.A(n9074), .B(n9076), .Y(n9197));
  XOR2X1  g7831(.A(n9197), .B(n9124), .Y(n9198));
  AOI22X1 g7832(.A0(n9032), .A1(n7678), .B0(n7053), .B1(n9048), .Y(n9199));
  OAI21X1 g7833(.A0(n9050), .A1(n6947), .B0(n9199), .Y(n9200));
  AOI22X1 g7834(.A0(n9046), .A1(n9200), .B0(P2_REG3_REG_22__SCAN_IN), .B1(P2_U3152), .Y(n9201));
  OAI21X1 g7835(.A0(n9044), .A1(n6988), .B0(n9201), .Y(n9202));
  AOI21X1 g7836(.A0(n9145), .A1(n7002), .B0(n9202), .Y(n9203));
  OAI21X1 g7837(.A0(n9198), .A1(n9039), .B0(n9203), .Y(P2_U3237));
  INVX1   g7838(.A(n8959), .Y(n9205));
  AOI21X1 g7839(.A0(n9022), .A1(n9021), .B0(n8952), .Y(n9206));
  OAI21X1 g7840(.A0(n8950), .A1(n8948), .B0(n8956), .Y(n9207));
  AOI21X1 g7841(.A0(n9206), .A1(n9205), .B0(n9207), .Y(n9208));
  AOI21X1 g7842(.A0(n8955), .A1(n8954), .B0(n9206), .Y(n9209));
  AOI21X1 g7843(.A0(n8950), .A1(n8958), .B0(n8959), .Y(n9210));
  OAI21X1 g7844(.A0(n8950), .A1(n8958), .B0(n9210), .Y(n9211));
  OAI21X1 g7845(.A0(n9211), .A1(n9209), .B0(n9038), .Y(n9212));
  OAI22X1 g7846(.A0(n9031), .A1(n6542), .B0(n6494), .B1(n9050), .Y(n9213));
  AOI21X1 g7847(.A0(n9048), .A1(n6660), .B0(n9213), .Y(n9214));
  AOI22X1 g7848(.A0(n6558), .A1(n9145), .B0(P2_REG3_REG_13__SCAN_IN), .B1(P2_U3152), .Y(n9215));
  OAI21X1 g7849(.A0(n9214), .A1(n9047), .B0(n9215), .Y(n9216));
  AOI21X1 g7850(.A0(n9045), .A1(n7598), .B0(n9216), .Y(n9217));
  OAI21X1 g7851(.A0(n9212), .A1(n9208), .B0(n9217), .Y(P2_U3236));
  XOR2X1  g7852(.A(n9090), .B(n9089), .Y(n9219));
  AOI21X1 g7853(.A0(n9085), .A1(n9084), .B0(n9121), .Y(n9220));
  NOR2X1  g7854(.A(n9220), .B(n9086), .Y(n9221));
  NOR2X1  g7855(.A(n9219), .B(n9221), .Y(n9223));
  AOI21X1 g7856(.A0(n9221), .A1(n9219), .B0(n9223), .Y(n9224));
  AOI22X1 g7857(.A0(n9032), .A1(n7659), .B0(n6872), .B1(n9049), .Y(n9225));
  OAI21X1 g7858(.A0(n9148), .A1(n6947), .B0(n9225), .Y(n9226));
  AOI22X1 g7859(.A0(n9046), .A1(n9226), .B0(P2_REG3_REG_20__SCAN_IN), .B1(P2_U3152), .Y(n9227));
  OAI21X1 g7860(.A0(n9044), .A1(n6888), .B0(n9227), .Y(n9228));
  AOI21X1 g7861(.A0(n9145), .A1(n6901), .B0(n9228), .Y(n9229));
  OAI21X1 g7862(.A0(n9224), .A1(n9039), .B0(n9229), .Y(P2_U3235));
  AOI21X1 g7863(.A0(n8379), .A1(n7494), .B0(n5750), .Y(n9231));
  AOI21X1 g7864(.A0(n9231), .A1(n9032), .B0(n9043), .Y(n9232));
  XOR2X1  g7865(.A(n8942), .B(n5923), .Y(n9233));
  XOR2X1  g7866(.A(n8995), .B(n8942), .Y(n9234));
  XOR2X1  g7867(.A(n9234), .B(n9233), .Y(n9235));
  NOR3X1  g7868(.A(n8379), .B(n5954), .C(n5750), .Y(n9236));
  AOI22X1 g7869(.A0(n9048), .A1(n9236), .B0(P2_REG3_REG_0__SCAN_IN), .B1(P2_U3152), .Y(n9237));
  OAI21X1 g7870(.A0(n9235), .A1(n9039), .B0(n9237), .Y(n9238));
  AOI21X1 g7871(.A0(n9145), .A1(n5877), .B0(n9238), .Y(n9239));
  OAI21X1 g7872(.A0(n9232), .A1(n5893), .B0(n9239), .Y(P2_U3234));
  XOR2X1  g7873(.A(n9018), .B(n8967), .Y(n9241));
  XOR2X1  g7874(.A(n9241), .B(n9016), .Y(n9242));
  OAI22X1 g7875(.A0(n9031), .A1(n6325), .B0(n6275), .B1(n9050), .Y(n9243));
  AOI21X1 g7876(.A0(n9048), .A1(n6386), .B0(n9243), .Y(n9244));
  AOI22X1 g7877(.A0(n6338), .A1(n9145), .B0(P2_REG3_REG_9__SCAN_IN), .B1(P2_U3152), .Y(n9245));
  OAI21X1 g7878(.A0(n9244), .A1(n9047), .B0(n9245), .Y(n9246));
  AOI21X1 g7879(.A0(n9045), .A1(n7563), .B0(n9246), .Y(n9247));
  OAI21X1 g7880(.A0(n9242), .A1(n9039), .B0(n9247), .Y(P2_U3233));
  NAND2X1 g7881(.A(n9045), .B(n6063), .Y(n9249));
  NOR2X1  g7882(.A(n9148), .B(n6121), .Y(n9250));
  OAI22X1 g7883(.A0(n9031), .A1(n6062), .B0(n6015), .B1(n9050), .Y(n9251));
  OAI21X1 g7884(.A0(n9251), .A1(n9250), .B0(n9046), .Y(n9252));
  XOR2X1  g7885(.A(n9007), .B(n8981), .Y(n9253));
  XOR2X1  g7886(.A(n9253), .B(n9004), .Y(n9254));
  NAND4X1 g7887(.A(n9036), .B(n9031), .C(n5743), .D(n9254), .Y(n9255));
  AOI22X1 g7888(.A0(n6112), .A1(n9145), .B0(P2_REG3_REG_4__SCAN_IN), .B1(P2_U3152), .Y(n9256));
  NAND4X1 g7889(.A(n9255), .B(n9252), .C(n9249), .D(n9256), .Y(P2_U3232));
  NOR2X1  g7890(.A(n9125), .B(n9073), .Y(n9258));
  NOR2X1  g7891(.A(n9258), .B(n9070), .Y(n9259));
  XOR2X1  g7892(.A(n9064), .B(n9063), .Y(n9260));
  AOI21X1 g7893(.A0(n9066), .A1(n9136), .B0(n9259), .Y(n9261));
  AOI21X1 g7894(.A0(n9260), .A1(n9259), .B0(n9261), .Y(n9262));
  NAND3X1 g7895(.A(n9146), .B(n7079), .C(P2_STATE_REG_SCAN_IN), .Y(n9263));
  AOI22X1 g7896(.A0(n9032), .A1(n7079), .B0(n7152), .B1(n9048), .Y(n9264));
  OAI21X1 g7897(.A0(n9050), .A1(n7038), .B0(n9264), .Y(n9265));
  AOI22X1 g7898(.A0(n9046), .A1(n9265), .B0(P2_REG3_REG_24__SCAN_IN), .B1(P2_U3152), .Y(n9266));
  NAND2X1 g7899(.A(n9266), .B(n9263), .Y(n9267));
  AOI21X1 g7900(.A0(n9145), .A1(n7165), .B0(n9267), .Y(n9268));
  OAI21X1 g7901(.A0(n9262), .A1(n9039), .B0(n9268), .Y(P2_U3231));
  OAI21X1 g7902(.A0(n9108), .A1(n9107), .B0(n9109), .Y(n9270));
  AOI21X1 g7903(.A0(n9117), .A1(n9115), .B0(n9270), .Y(n9271));
  AOI21X1 g7904(.A0(n9104), .A1(n9103), .B0(n9115), .Y(n9272));
  INVX1   g7905(.A(n9108), .Y(n9273));
  AOI21X1 g7906(.A0(n9273), .A1(n9107), .B0(n9116), .Y(n9274));
  OAI21X1 g7907(.A0(n9273), .A1(n9107), .B0(n9274), .Y(n9275));
  OAI21X1 g7908(.A0(n9275), .A1(n9272), .B0(n9038), .Y(n9276));
  OAI22X1 g7909(.A0(n9031), .A1(n6734), .B0(n6690), .B1(n9050), .Y(n9277));
  AOI21X1 g7910(.A0(n9048), .A1(n6818), .B0(n9277), .Y(n9278));
  OAI22X1 g7911(.A0(n9047), .A1(n9278), .B0(n6732), .B1(P2_STATE_REG_SCAN_IN), .Y(n9279));
  OAI22X1 g7912(.A0(n9044), .A1(n6734), .B0(n6754), .B1(n9053), .Y(n9280));
  NOR2X1  g7913(.A(n9280), .B(n9279), .Y(n9281));
  OAI21X1 g7914(.A0(n9276), .A1(n9271), .B0(n9281), .Y(P2_U3230));
  NAND2X1 g7915(.A(n9008), .B(n9005), .Y(n9283));
  XOR2X1  g7916(.A(n8979), .B(n8978), .Y(n9284));
  XOR2X1  g7917(.A(n9284), .B(n9283), .Y(n9285));
  NAND2X1 g7918(.A(n9285), .B(n9038), .Y(n9286));
  NAND2X1 g7919(.A(n9048), .B(n6231), .Y(n9287));
  AOI22X1 g7920(.A0(n9032), .A1(n6144), .B0(n6065), .B1(n9049), .Y(n9288));
  AOI21X1 g7921(.A0(n9288), .A1(n9287), .B0(n9047), .Y(n9289));
  AOI22X1 g7922(.A0(n6133), .A1(n9145), .B0(P2_REG3_REG_5__SCAN_IN), .B1(P2_U3152), .Y(n9290));
  OAI21X1 g7923(.A0(n9044), .A1(n6119), .B0(n9290), .Y(n9291));
  NOR2X1  g7924(.A(n9291), .B(n9289), .Y(n9292));
  NAND2X1 g7925(.A(n9292), .B(n9286), .Y(P2_U3229));
  XOR2X1  g7926(.A(n9104), .B(n9103), .Y(n9294));
  NOR2X1  g7927(.A(n9294), .B(n9115), .Y(n9296));
  AOI21X1 g7928(.A0(n9294), .A1(n9115), .B0(n9296), .Y(n9297));
  OAI22X1 g7929(.A0(n9031), .A1(n6686), .B0(n6646), .B1(n9050), .Y(n9298));
  AOI21X1 g7930(.A0(n9048), .A1(n6747), .B0(n9298), .Y(n9299));
  AOI22X1 g7931(.A0(n6704), .A1(n9145), .B0(P2_REG3_REG_16__SCAN_IN), .B1(P2_U3152), .Y(n9300));
  OAI21X1 g7932(.A0(n9299), .A1(n9047), .B0(n9300), .Y(n9301));
  AOI21X1 g7933(.A0(n9045), .A1(n6687), .B0(n9301), .Y(n9302));
  OAI21X1 g7934(.A0(n9297), .A1(n9039), .B0(n9302), .Y(P2_U3228));
  XOR2X1  g7935(.A(n9061), .B(n9060), .Y(n9304));
  NOR2X1  g7936(.A(n9304), .B(n9127), .Y(n9306));
  AOI21X1 g7937(.A0(n9304), .A1(n9127), .B0(n9306), .Y(n9307));
  AOI22X1 g7938(.A0(n9032), .A1(n7122), .B0(n7183), .B1(n9048), .Y(n9308));
  OAI21X1 g7939(.A0(n9050), .A1(n7083), .B0(n9308), .Y(n9309));
  AOI22X1 g7940(.A0(n9046), .A1(n9309), .B0(P2_REG3_REG_25__SCAN_IN), .B1(P2_U3152), .Y(n9310));
  OAI21X1 g7941(.A0(n9044), .A1(n7121), .B0(n9310), .Y(n9311));
  AOI21X1 g7942(.A0(n9145), .A1(n7134), .B0(n9311), .Y(n9312));
  OAI21X1 g7943(.A0(n9307), .A1(n9039), .B0(n9312), .Y(P2_U3227));
  XOR2X1  g7944(.A(n8955), .B(n8954), .Y(n9314));
  NOR2X1  g7945(.A(n9314), .B(n9206), .Y(n9316));
  AOI21X1 g7946(.A0(n9314), .A1(n9206), .B0(n9316), .Y(n9317));
  OAI22X1 g7947(.A0(n9031), .A1(n6490), .B0(n6430), .B1(n9050), .Y(n9318));
  AOI21X1 g7948(.A0(n9048), .A1(n6545), .B0(n9318), .Y(n9319));
  AOI22X1 g7949(.A0(n6506), .A1(n9145), .B0(P2_REG3_REG_12__SCAN_IN), .B1(P2_U3152), .Y(n9320));
  OAI21X1 g7950(.A0(n9319), .A1(n9047), .B0(n9320), .Y(n9321));
  AOI21X1 g7951(.A0(n9045), .A1(n6491), .B0(n9321), .Y(n9322));
  OAI21X1 g7952(.A0(n9317), .A1(n9039), .B0(n9322), .Y(P2_U3226));
  NOR3X1  g7953(.A(n9220), .B(n9093), .C(n9086), .Y(n9324));
  OAI21X1 g7954(.A0(n9088), .A1(n9080), .B0(n9091), .Y(n9325));
  NOR2X1  g7955(.A(n9325), .B(n9324), .Y(n9326));
  AOI21X1 g7956(.A0(n9090), .A1(n9089), .B0(n9221), .Y(n9327));
  AOI21X1 g7957(.A0(n9088), .A1(n9081), .B0(n9093), .Y(n9328));
  OAI21X1 g7958(.A0(n9088), .A1(n9081), .B0(n9328), .Y(n9329));
  OAI21X1 g7959(.A0(n9329), .A1(n9327), .B0(n9038), .Y(n9330));
  AOI22X1 g7960(.A0(n9032), .A1(n7668), .B0(n6914), .B1(n9049), .Y(n9331));
  OAI21X1 g7961(.A0(n9148), .A1(n6995), .B0(n9331), .Y(n9332));
  AOI22X1 g7962(.A0(n9046), .A1(n9332), .B0(P2_REG3_REG_21__SCAN_IN), .B1(P2_U3152), .Y(n9333));
  OAI21X1 g7963(.A0(n9044), .A1(n6941), .B0(n9333), .Y(n9334));
  AOI21X1 g7964(.A0(n9145), .A1(n6954), .B0(n9334), .Y(n9335));
  OAI21X1 g7965(.A0(n9330), .A1(n9326), .B0(n9335), .Y(P2_U3225));
  NAND2X1 g7966(.A(n9045), .B(P2_REG3_REG_1__SCAN_IN), .Y(n9337));
  NOR2X1  g7967(.A(n9148), .B(n5974), .Y(n9338));
  OAI22X1 g7968(.A0(n9031), .A1(n5951), .B0(n5897), .B1(n9050), .Y(n9339));
  OAI21X1 g7969(.A0(n9339), .A1(n9338), .B0(n9046), .Y(n9340));
  NAND2X1 g7970(.A(n9145), .B(n5939), .Y(n9341));
  XOR2X1  g7971(.A(n8990), .B(n8989), .Y(n9342));
  XOR2X1  g7972(.A(n9342), .B(n8997), .Y(n9343));
  AOI22X1 g7973(.A0(n9038), .A1(n9343), .B0(P2_REG3_REG_1__SCAN_IN), .B1(P2_U3152), .Y(n9344));
  NAND4X1 g7974(.A(n9341), .B(n9340), .C(n9337), .D(n9344), .Y(P2_U3224));
  XOR2X1  g7975(.A(n8969), .B(n8968), .Y(n9346));
  XOR2X1  g7976(.A(n9346), .B(n9015), .Y(n9347));
  NAND2X1 g7977(.A(n9347), .B(n9038), .Y(n9348));
  OAI22X1 g7978(.A0(n9031), .A1(n6273), .B0(n6223), .B1(n9050), .Y(n9349));
  AOI21X1 g7979(.A0(n9048), .A1(n6354), .B0(n9349), .Y(n9350));
  AOI22X1 g7980(.A0(n6289), .A1(n9145), .B0(P2_REG3_REG_8__SCAN_IN), .B1(P2_U3152), .Y(n9351));
  OAI21X1 g7981(.A0(n9350), .A1(n9047), .B0(n9351), .Y(n9352));
  AOI21X1 g7982(.A0(n9045), .A1(n7555), .B0(n9352), .Y(n9353));
  NAND2X1 g7983(.A(n9353), .B(n9348), .Y(P2_U3223));
  XOR2X1  g7984(.A(n8994), .B(n7243), .Y(n9355));
  OAI21X1 g7985(.A0(n8938), .A1(n7228), .B0(n9355), .Y(n9356));
  INVX1   g7986(.A(n9356), .Y(n9357));
  NAND2X1 g7987(.A(n9141), .B(n9066), .Y(n9358));
  NOR2X1  g7988(.A(n9358), .B(n9357), .Y(n9359));
  NOR2X1  g7989(.A(n8938), .B(n7283), .Y(n9360));
  XOR2X1  g7990(.A(n9360), .B(n8994), .Y(n9361));
  XOR2X1  g7991(.A(n9361), .B(n7290), .Y(n9362));
  NOR3X1  g7992(.A(n9355), .B(n8938), .C(n7228), .Y(n9363));
  INVX1   g7993(.A(n9363), .Y(n9364));
  NOR2X1  g7994(.A(n9131), .B(n9130), .Y(n9365));
  AOI21X1 g7995(.A0(n9137), .A1(n9136), .B0(n9140), .Y(n9366));
  OAI21X1 g7996(.A0(n9366), .A1(n9365), .B0(n9356), .Y(n9367));
  NAND3X1 g7997(.A(n9367), .B(n9364), .C(n9362), .Y(n9368));
  AOI21X1 g7998(.A0(n9359), .A1(n9126), .B0(n9368), .Y(n9369));
  NOR3X1  g7999(.A(n9366), .B(n9363), .C(n9365), .Y(n9370));
  OAI21X1 g8000(.A0(n9358), .A1(n9259), .B0(n9370), .Y(n9371));
  NOR2X1  g8001(.A(n9362), .B(n9357), .Y(n9372));
  AOI21X1 g8002(.A0(n9372), .A1(n9371), .B0(n9369), .Y(n9373));
  AOI22X1 g8003(.A0(n9032), .A1(n7278), .B0(n7326), .B1(n9048), .Y(n9374));
  OAI21X1 g8004(.A0(n9050), .A1(n7228), .B0(n9374), .Y(n9375));
  AOI22X1 g8005(.A0(n9046), .A1(n9375), .B0(P2_REG3_REG_28__SCAN_IN), .B1(P2_U3152), .Y(n9376));
  OAI21X1 g8006(.A0(n9044), .A1(n7277), .B0(n9376), .Y(n9377));
  AOI21X1 g8007(.A0(n9145), .A1(n7290), .B0(n9377), .Y(n9378));
  OAI21X1 g8008(.A0(n9373), .A1(n9039), .B0(n9378), .Y(P2_U3222));
  XOR2X1  g8009(.A(n9085), .B(n9084), .Y(n9380));
  NOR2X1  g8010(.A(n9380), .B(n9121), .Y(n9382));
  AOI21X1 g8011(.A0(n9380), .A1(n9121), .B0(n9382), .Y(n9383));
  AOI22X1 g8012(.A0(n9032), .A1(n7651), .B0(n6818), .B1(n9049), .Y(n9384));
  OAI21X1 g8013(.A0(n9148), .A1(n6894), .B0(n9384), .Y(n9385));
  AOI22X1 g8014(.A0(n9046), .A1(n9385), .B0(P2_REG3_REG_19__SCAN_IN), .B1(P2_U3152), .Y(n9386));
  OAI21X1 g8015(.A0(n9044), .A1(n6839), .B0(n9386), .Y(n9387));
  AOI21X1 g8016(.A0(n9145), .A1(n6854), .B0(n9387), .Y(n9388));
  OAI21X1 g8017(.A0(n9383), .A1(n9039), .B0(n9388), .Y(P2_U3221));
  NAND2X1 g8018(.A(n9048), .B(n6065), .Y(n9390));
  AOI22X1 g8019(.A0(n9032), .A1(n6026), .B0(n5995), .B1(n9049), .Y(n9391));
  AOI21X1 g8020(.A0(n9391), .A1(n9390), .B0(n9047), .Y(n9392));
  NOR2X1  g8021(.A(n9053), .B(n6034), .Y(n9393));
  NAND2X1 g8022(.A(n9001), .B(n8998), .Y(n9394));
  AOI21X1 g8023(.A0(n8987), .A1(n8985), .B0(n8988), .Y(n9395));
  NOR2X1  g8024(.A(n8983), .B(n8982), .Y(n9396));
  OAI21X1 g8025(.A0(n8986), .A1(n8985), .B0(n9001), .Y(n9397));
  AOI21X1 g8026(.A0(n8986), .A1(n8985), .B0(n9397), .Y(n9398));
  OAI21X1 g8027(.A0(n8998), .A1(n9396), .B0(n9398), .Y(n9399));
  NAND4X1 g8028(.A(n9036), .B(n9031), .C(n5743), .D(n9399), .Y(n9400));
  AOI21X1 g8029(.A0(n9395), .A1(n9394), .B0(n9400), .Y(n9401));
  NOR4X1  g8030(.A(n9393), .B(n9392), .C(n8255), .D(n9401), .Y(n9402));
  OAI21X1 g8031(.A0(n9044), .A1(P2_REG3_REG_3__SCAN_IN), .B0(n9402), .Y(P2_U3220));
  NOR2X1  g8032(.A(n9019), .B(n9017), .Y(n9404));
  XOR2X1  g8033(.A(n8964), .B(n8963), .Y(n9405));
  XOR2X1  g8034(.A(n9405), .B(n9404), .Y(n9406));
  OAI22X1 g8035(.A0(n9031), .A1(n6372), .B0(n6327), .B1(n9050), .Y(n9407));
  AOI21X1 g8036(.A0(n9048), .A1(n6451), .B0(n9407), .Y(n9408));
  AOI22X1 g8037(.A0(n6391), .A1(n9145), .B0(P2_REG3_REG_10__SCAN_IN), .B1(P2_U3152), .Y(n9409));
  OAI21X1 g8038(.A0(n9408), .A1(n9047), .B0(n9409), .Y(n9410));
  AOI21X1 g8039(.A0(n9045), .A1(n6384), .B0(n9410), .Y(n9411));
  OAI21X1 g8040(.A0(n9406), .A1(n9039), .B0(n9411), .Y(P2_U3219));
  XOR2X1  g8041(.A(n9069), .B(n9068), .Y(n9413));
  XOR2X1  g8042(.A(n9413), .B(n9125), .Y(n9414));
  AOI22X1 g8043(.A0(n9032), .A1(n7033), .B0(n7090), .B1(n9048), .Y(n9415));
  OAI21X1 g8044(.A0(n9050), .A1(n6995), .B0(n9415), .Y(n9416));
  AOI22X1 g8045(.A0(n9046), .A1(n9416), .B0(P2_REG3_REG_23__SCAN_IN), .B1(P2_U3152), .Y(n9417));
  OAI21X1 g8046(.A0(n9044), .A1(n7032), .B0(n9417), .Y(n9418));
  AOI21X1 g8047(.A0(n9145), .A1(n7049), .B0(n9418), .Y(n9419));
  OAI21X1 g8048(.A0(n9414), .A1(n9039), .B0(n9419), .Y(P2_U3218));
  XOR2X1  g8049(.A(n8943), .B(n8940), .Y(n9421));
  XOR2X1  g8050(.A(n9421), .B(n9025), .Y(n9422));
  NOR2X1  g8051(.A(n9044), .B(n6595), .Y(n9423));
  OAI22X1 g8052(.A0(n9031), .A1(n6595), .B0(n6546), .B1(n9050), .Y(n9424));
  AOI21X1 g8053(.A0(n9048), .A1(n6645), .B0(n9424), .Y(n9425));
  AOI22X1 g8054(.A0(n6609), .A1(n9145), .B0(P2_REG3_REG_14__SCAN_IN), .B1(P2_U3152), .Y(n9426));
  OAI21X1 g8055(.A0(n9425), .A1(n9047), .B0(n9426), .Y(n9427));
  NOR2X1  g8056(.A(n9427), .B(n9423), .Y(n9428));
  OAI21X1 g8057(.A0(n9422), .A1(n9039), .B0(n9428), .Y(P2_U3217));
  NOR2X1  g8058(.A(n9366), .B(n9365), .Y(n9430));
  OAI21X1 g8059(.A0(n9358), .A1(n9259), .B0(n9430), .Y(n9431));
  NOR2X1  g8060(.A(n8938), .B(n7228), .Y(n9432));
  XOR2X1  g8061(.A(n9432), .B(n9355), .Y(n9433));
  XOR2X1  g8062(.A(n9433), .B(n9431), .Y(n9434));
  NOR2X1  g8063(.A(n9148), .B(n7283), .Y(n9435));
  OAI22X1 g8064(.A0(n9031), .A1(n7222), .B0(n7176), .B1(n9050), .Y(n9436));
  OAI21X1 g8065(.A0(n9436), .A1(n9435), .B0(n9046), .Y(n9437));
  NAND2X1 g8066(.A(P2_REG3_REG_27__SCAN_IN), .B(P2_U3152), .Y(n9438));
  NAND3X1 g8067(.A(n9146), .B(n7223), .C(P2_STATE_REG_SCAN_IN), .Y(n9439));
  NAND3X1 g8068(.A(n9439), .B(n9438), .C(n9437), .Y(n9440));
  AOI21X1 g8069(.A0(n9145), .A1(n7272), .B0(n9440), .Y(n9441));
  OAI21X1 g8070(.A0(n9434), .A1(n9039), .B0(n9441), .Y(P2_U3216));
  NOR3X1  g8071(.A(n9011), .B(n9009), .C(n8980), .Y(n9443));
  OAI21X1 g8072(.A0(n8976), .A1(n8975), .B0(n8977), .Y(n9444));
  INVX1   g8073(.A(n8972), .Y(n9445));
  INVX1   g8074(.A(n8973), .Y(n9446));
  OAI22X1 g8075(.A0(n8980), .A1(n9009), .B0(n9446), .B1(n9445), .Y(n9447));
  OAI22X1 g8076(.A0(n8974), .A1(n8976), .B0(n8973), .B1(n8972), .Y(n9448));
  AOI21X1 g8077(.A0(n8976), .A1(n8974), .B0(n9448), .Y(n9449));
  AOI21X1 g8078(.A0(n9449), .A1(n9447), .B0(n9039), .Y(n9450));
  OAI21X1 g8079(.A0(n9444), .A1(n9443), .B0(n9450), .Y(n9451));
  OAI22X1 g8080(.A0(n9031), .A1(n6221), .B0(n6172), .B1(n9050), .Y(n9452));
  AOI21X1 g8081(.A0(n9048), .A1(n6292), .B0(n9452), .Y(n9453));
  AOI22X1 g8082(.A0(n6239), .A1(n9145), .B0(P2_REG3_REG_7__SCAN_IN), .B1(P2_U3152), .Y(n9454));
  OAI21X1 g8083(.A0(n9453), .A1(n9047), .B0(n9454), .Y(n9455));
  AOI21X1 g8084(.A0(n9045), .A1(n7543), .B0(n9455), .Y(n9456));
  NAND2X1 g8085(.A(n9456), .B(n9451), .Y(P2_U3215));
  NOR2X1  g8086(.A(n5742), .B(n5735), .Y(n9458));
  NAND2X1 g8087(.A(n7752), .B(n9458), .Y(n9459));
  NOR2X1  g8088(.A(n7751), .B(P2_U3152), .Y(n9460));
  NAND2X1 g8089(.A(n9460), .B(n9459), .Y(P2_U3151));
endmodule


