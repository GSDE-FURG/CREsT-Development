//Converted to Combinational , Module name: s420 , Timestamp: 2018-12-03T15:51:01.631077 
module s420 ( X, Clear, C_16, C_15, C_14, C_13, C_12, C_11, C_10, C_9, C_8, C_7, C_6, C_5, C_4, C_3, C_2, C_0, Y_4, Y_3, Y_2, Y_1, Y_8, Y_7, Y_6, Y_5, Y_12, Y_11, Y_10, Y_9, Y_16, Y_15, Y_14, Y_13, W, Z, n43, n48, n53, n58, n63, n68, n73, n78, n83, n88, n93, n98, n103, n108, n113, n118 );
input C_1, X, Clear, C_16, C_15, C_14, C_13, C_12, C_11, C_10, C_9, C_8, C_7, C_6, C_5, C_4, C_3, C_2, C_0, Y_4, Y_3, Y_2, Y_1, Y_8, Y_7, Y_6, Y_5, Y_12, Y_11, Y_10, Y_9, Y_16, Y_15, Y_14, Y_13;
output W, Z, n43, n48, n53, n58, n63, n68, n73, n78, n83, n88, n93, n98, n103, n108, n113, n118;
wire n69, n70, n72, n73_1, n74, n75, n76, n77, n78_1, n79, n80, n81, n82, n83_1, n84, n85, n86, n87, n88_1, n89, n90, n91, n92, n93_1, n94, n95, n96, n97, n98_1, n99, n100, n101, n102, n103_1, n104, n105, n106, n107, n108_1, n109, n110, n111, n112, n113_1, n114, n115, n116, n117, n119, n120, n121, n122, n123, n124, n126, n127, n129, n132, n133, n134, n135, n136, n138, n139, n140, n144, n145, n146, n147, n148, n149, n151, n152, n153, n157, n158, n159, n160, n161, n163, n164, n165;
INVX1    g00(.A(Y_16), .Y(n69));
NAND3X1  g01(.A(Y_13), .B(Y_14), .C(Y_15), .Y(n70));
NOR2X1   g02(.A(n70), .B(n69), .Y(W));
INVX1    g03(.A(C_14), .Y(n72));
INVX1    g04(.A(Y_14), .Y(n73_1));
INVX1    g05(.A(Y_8), .Y(n74));
INVX1    g06(.A(Y_7), .Y(n75));
INVX1    g07(.A(Y_9), .Y(n76));
INVX1    g08(.A(X), .Y(n77));
OR4X1    g09(.A(Y_2), .B(Y_3), .C(n77), .D(Y_1), .Y(n78_1));
NOR4X1   g10(.A(Y_5), .B(Y_6), .C(Y_4), .D(n78_1), .Y(n79));
NAND4X1  g11(.A(n76), .B(n75), .C(n74), .D(n79), .Y(n80));
OR4X1    g12(.A(Y_10), .B(Y_11), .C(Y_12), .D(n80), .Y(n81));
OR4X1    g13(.A(Y_13), .B(n73_1), .C(n72), .D(n81), .Y(n82));
NAND2X1  g14(.A(Y_13), .B(C_13), .Y(n83_1));
NOR2X1   g15(.A(n83_1), .B(n81), .Y(n84));
NAND2X1  g16(.A(Y_12), .B(C_12), .Y(n85));
NOR4X1   g17(.A(n80), .B(Y_10), .C(Y_11), .D(n85), .Y(n86));
NAND2X1  g18(.A(Y_11), .B(C_11), .Y(n87));
NOR3X1   g19(.A(n87), .B(n80), .C(Y_10), .Y(n88_1));
NAND2X1  g20(.A(Y_10), .B(C_10), .Y(n89));
OR2X1    g21(.A(n89), .B(n80), .Y(n90));
AND2X1   g22(.A(Y_9), .B(C_9), .Y(n91));
NAND4X1  g23(.A(n79), .B(n75), .C(n74), .D(n91), .Y(n92));
NAND4X1  g24(.A(n75), .B(Y_8), .C(C_8), .D(n79), .Y(n93_1));
AND2X1   g25(.A(Y_7), .B(C_7), .Y(n94));
AND2X1   g26(.A(n94), .B(n79), .Y(n95));
NAND2X1  g27(.A(Y_6), .B(C_6), .Y(n96));
NOR4X1   g28(.A(n78_1), .B(Y_5), .C(Y_4), .D(n96), .Y(n97));
NAND2X1  g29(.A(Y_5), .B(C_5), .Y(n98_1));
NOR3X1   g30(.A(n98_1), .B(n78_1), .C(Y_4), .Y(n99));
NAND2X1  g31(.A(Y_4), .B(C_4), .Y(n100));
OR2X1    g32(.A(n100), .B(n78_1), .Y(n101));
INVX1    g33(.A(Y_2), .Y(n102));
INVX1    g34(.A(Y_1), .Y(n103_1));
AND2X1   g35(.A(Y_3), .B(C_3), .Y(n104));
NAND4X1  g36(.A(n103_1), .B(n102), .C(X), .D(n104), .Y(n105));
NAND4X1  g37(.A(Y_2), .B(C_2), .C(X), .D(n103_1), .Y(n106));
AND2X1   g38(.A(Y_1), .B(C_1), .Y(n107));
OAI21X1  g39(.A0(n107), .A1(C_0), .B0(X), .Y(n108_1));
NAND4X1  g40(.A(n106), .B(n105), .C(n101), .D(n108_1), .Y(n109));
NOR4X1   g41(.A(n99), .B(n97), .C(n95), .D(n109), .Y(n110));
NAND4X1  g42(.A(n93_1), .B(n92), .C(n90), .D(n110), .Y(n111));
NOR4X1   g43(.A(n88_1), .B(n86), .C(n84), .D(n111), .Y(n112));
NOR3X1   g44(.A(n81), .B(Y_13), .C(Y_14), .Y(n113_1));
AND2X1   g45(.A(Y_15), .B(C_15), .Y(n114));
NAND2X1  g46(.A(Y_16), .B(C_16), .Y(n115));
NOR2X1   g47(.A(n115), .B(Y_15), .Y(n116));
OAI21X1  g48(.A0(n116), .A1(n114), .B0(n113_1), .Y(n117));
NAND3X1  g49(.A(n117), .B(n112), .C(n82), .Y(Z));
INVX1    g50(.A(Clear), .Y(n119));
NAND4X1  g51(.A(Y_2), .B(n119), .C(X), .D(Y_1), .Y(n120));
INVX1    g52(.A(Y_4), .Y(n121));
NAND2X1  g53(.A(Y_3), .B(n121), .Y(n122));
NAND3X1  g54(.A(Y_1), .B(Y_2), .C(Y_3), .Y(n123));
NAND4X1  g55(.A(Y_4), .B(n119), .C(X), .D(n123), .Y(n124));
OAI21X1  g56(.A0(n122), .A1(n120), .B0(n124), .Y(n43));
NAND2X1  g57(.A(n119), .B(X), .Y(n126));
OAI21X1  g58(.A0(n103_1), .A1(n102), .B0(Y_3), .Y(n127));
OAI22X1  g59(.A0(n120), .A1(Y_3), .B0(n126), .B1(n127), .Y(n48));
NOR3X1   g60(.A(n103_1), .B(Clear), .C(n77), .Y(n129));
NOR3X1   g61(.A(Y_1), .B(Clear), .C(n77), .Y(n58));
MX2X1    g62(.A(n129), .B(n58), .S0(Y_2), .Y(n53));
NOR3X1   g63(.A(n123), .B(n121), .C(Clear), .Y(n132));
AND2X1   g64(.A(n132), .B(Y_5), .Y(n133));
NAND4X1  g65(.A(Y_6), .B(Y_7), .C(n74), .D(n133), .Y(n134));
NAND3X1  g66(.A(Y_5), .B(Y_6), .C(Y_7), .Y(n135));
NAND3X1  g67(.A(n135), .B(n132), .C(Y_8), .Y(n136));
NAND2X1  g68(.A(n136), .B(n134), .Y(n63));
NAND2X1  g69(.A(Y_5), .B(Y_6), .Y(n138));
NAND3X1  g70(.A(n138), .B(n132), .C(Y_7), .Y(n139));
NAND4X1  g71(.A(Y_5), .B(Y_6), .C(n75), .D(n132), .Y(n140));
NAND2X1  g72(.A(n140), .B(n139), .Y(n68));
NOR4X1   g73(.A(Y_5), .B(n121), .C(Clear), .D(n123), .Y(n78));
MX2X1    g74(.A(n133), .B(n78), .S0(Y_6), .Y(n73));
INVX1    g75(.A(Y_12), .Y(n144));
NOR4X1   g76(.A(n76), .B(n74), .C(Clear), .D(n135), .Y(n145));
NAND4X1  g77(.A(Y_10), .B(Y_11), .C(n144), .D(n145), .Y(n146));
NOR3X1   g78(.A(n135), .B(n74), .C(Clear), .Y(n147));
NAND3X1  g79(.A(Y_9), .B(Y_10), .C(Y_11), .Y(n148));
NAND3X1  g80(.A(n148), .B(n147), .C(Y_12), .Y(n149));
NAND2X1  g81(.A(n149), .B(n146), .Y(n83));
NAND2X1  g82(.A(n145), .B(Y_10), .Y(n151));
NAND2X1  g83(.A(Y_9), .B(Y_10), .Y(n152));
NAND3X1  g84(.A(n152), .B(n147), .C(Y_11), .Y(n153));
OAI21X1  g85(.A0(n151), .A1(Y_11), .B0(n153), .Y(n88));
NOR4X1   g86(.A(Y_9), .B(n74), .C(Clear), .D(n135), .Y(n98));
MX2X1    g87(.A(n145), .B(n98), .S0(Y_10), .Y(n93));
INVX1    g88(.A(Y_13), .Y(n157));
NOR4X1   g89(.A(n157), .B(n144), .C(Clear), .D(n148), .Y(n158));
NAND4X1  g90(.A(Y_14), .B(Y_15), .C(n69), .D(n158), .Y(n159));
NOR3X1   g91(.A(n148), .B(n144), .C(Clear), .Y(n160));
NAND3X1  g92(.A(n160), .B(n70), .C(Y_16), .Y(n161));
NAND2X1  g93(.A(n161), .B(n159), .Y(n103));
NAND2X1  g94(.A(n158), .B(Y_14), .Y(n163));
NAND2X1  g95(.A(Y_13), .B(Y_14), .Y(n164));
NAND3X1  g96(.A(n160), .B(n164), .C(Y_15), .Y(n165));
OAI21X1  g97(.A0(n163), .A1(Y_15), .B0(n165), .Y(n108));
NOR4X1   g98(.A(Y_13), .B(n144), .C(Clear), .D(n148), .Y(n118));
MX2X1    g99(.A(n158), .B(n118), .S0(Y_14), .Y(n113));
endmodule
