// Benchmark "b14_C" written by ABC on Wed Aug 05 14:40:44 2020

module b14_C ( 
    WR_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_,
    DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_,
    DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_,
    DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_,
    DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_,
    DATAI_1_, DATAI_0_, RD_REG_SCAN_IN, STATE_REG_SCAN_IN,
    REG3_REG_7__SCAN_IN, REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN,
    REG3_REG_23__SCAN_IN, REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN,
    REG3_REG_19__SCAN_IN, REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN,
    REG3_REG_1__SCAN_IN, REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN,
    REG3_REG_25__SCAN_IN, REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN,
    REG3_REG_17__SCAN_IN, REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN,
    REG3_REG_9__SCAN_IN, REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN,
    REG3_REG_13__SCAN_IN, IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN,
    IR_REG_2__SCAN_IN, IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN,
    IR_REG_5__SCAN_IN, IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN,
    IR_REG_8__SCAN_IN, IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN,
    IR_REG_11__SCAN_IN, IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN,
    IR_REG_14__SCAN_IN, IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN,
    IR_REG_17__SCAN_IN, IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN,
    IR_REG_20__SCAN_IN, IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN,
    IR_REG_23__SCAN_IN, IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN,
    IR_REG_26__SCAN_IN, IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN,
    IR_REG_29__SCAN_IN, IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN,
    D_REG_0__SCAN_IN, D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
    D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN,
    D_REG_8__SCAN_IN, D_REG_9__SCAN_IN, D_REG_10__SCAN_IN,
    D_REG_11__SCAN_IN, D_REG_12__SCAN_IN, D_REG_13__SCAN_IN,
    D_REG_14__SCAN_IN, D_REG_15__SCAN_IN, D_REG_16__SCAN_IN,
    D_REG_17__SCAN_IN, D_REG_18__SCAN_IN, D_REG_19__SCAN_IN,
    D_REG_20__SCAN_IN, D_REG_21__SCAN_IN, D_REG_22__SCAN_IN,
    D_REG_23__SCAN_IN, D_REG_24__SCAN_IN, D_REG_25__SCAN_IN,
    D_REG_26__SCAN_IN, D_REG_27__SCAN_IN, D_REG_28__SCAN_IN,
    D_REG_29__SCAN_IN, D_REG_30__SCAN_IN, D_REG_31__SCAN_IN,
    REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN,
    REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN,
    REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN,
    REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN,
    REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN,
    REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN,
    REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN,
    REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN,
    REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN,
    REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN,
    REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN,
    REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN,
    REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN,
    REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN,
    REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN,
    REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN,
    REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN,
    REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN,
    REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN,
    REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN,
    REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN,
    REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN,
    REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN,
    REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN,
    REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN,
    REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN,
    REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN,
    REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN,
    REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN,
    REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN,
    REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN,
    REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN,
    ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN,
    ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN,
    ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN,
    ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN,
    ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN,
    ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN,
    ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN,
    DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN,
    DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN,
    DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN,
    DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN,
    DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN,
    DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN,
    DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN,
    DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN,
    DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN,
    DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN,
    DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN, REG3_REG_15__SCAN_IN,
    REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN,
    REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN,
    U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
    U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
    U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
    U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
    U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
    U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
    U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
    U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
    U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
    U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
    U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
    U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
    U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
    U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
    U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
    U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
    U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
    U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
    U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
    U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
    U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
    U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
    U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
    U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
    U3211, U3210, U3149, U3148, U4043  );
  input  WR_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
    DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
    DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
    DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
    DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
    DATAI_2_, DATAI_1_, DATAI_0_, RD_REG_SCAN_IN, STATE_REG_SCAN_IN,
    REG3_REG_7__SCAN_IN, REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN,
    REG3_REG_23__SCAN_IN, REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN,
    REG3_REG_19__SCAN_IN, REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN,
    REG3_REG_1__SCAN_IN, REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN,
    REG3_REG_25__SCAN_IN, REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN,
    REG3_REG_17__SCAN_IN, REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN,
    REG3_REG_9__SCAN_IN, REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN,
    REG3_REG_13__SCAN_IN, IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN,
    IR_REG_2__SCAN_IN, IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN,
    IR_REG_5__SCAN_IN, IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN,
    IR_REG_8__SCAN_IN, IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN,
    IR_REG_11__SCAN_IN, IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN,
    IR_REG_14__SCAN_IN, IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN,
    IR_REG_17__SCAN_IN, IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN,
    IR_REG_20__SCAN_IN, IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN,
    IR_REG_23__SCAN_IN, IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN,
    IR_REG_26__SCAN_IN, IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN,
    IR_REG_29__SCAN_IN, IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN,
    D_REG_0__SCAN_IN, D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
    D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN,
    D_REG_8__SCAN_IN, D_REG_9__SCAN_IN, D_REG_10__SCAN_IN,
    D_REG_11__SCAN_IN, D_REG_12__SCAN_IN, D_REG_13__SCAN_IN,
    D_REG_14__SCAN_IN, D_REG_15__SCAN_IN, D_REG_16__SCAN_IN,
    D_REG_17__SCAN_IN, D_REG_18__SCAN_IN, D_REG_19__SCAN_IN,
    D_REG_20__SCAN_IN, D_REG_21__SCAN_IN, D_REG_22__SCAN_IN,
    D_REG_23__SCAN_IN, D_REG_24__SCAN_IN, D_REG_25__SCAN_IN,
    D_REG_26__SCAN_IN, D_REG_27__SCAN_IN, D_REG_28__SCAN_IN,
    D_REG_29__SCAN_IN, D_REG_30__SCAN_IN, D_REG_31__SCAN_IN,
    REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN,
    REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN,
    REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN,
    REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN,
    REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN,
    REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN,
    REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN,
    REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN,
    REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN,
    REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN,
    REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN,
    REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN,
    REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN,
    REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN,
    REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN,
    REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN,
    REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN,
    REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN,
    REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN,
    REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN,
    REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN,
    REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN,
    REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN,
    REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN,
    REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN,
    REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN,
    REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN,
    REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN,
    REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN,
    REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN,
    REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN,
    REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN,
    ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN,
    ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN,
    ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN,
    ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN,
    ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN,
    ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN,
    ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN,
    DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN,
    DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN,
    DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN,
    DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN,
    DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN,
    DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN,
    DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN,
    DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN,
    DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN,
    DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN,
    DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN, REG3_REG_15__SCAN_IN,
    REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN,
    REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
    U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
    U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
    U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
    U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
    U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
    U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
    U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
    U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
    U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
    U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
    U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
    U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
    U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
    U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
    U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
    U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
    U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
    U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
    U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
    U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
    U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
    U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
    U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
    U3211, U3210, U3149, U3148, U4043;
  wire n576, n577, n579, n580, n582, n583, n585, n586, n587, n589, n590,
    n591, n593, n594, n595, n597, n598, n599, n600, n601, n602, n603, n605,
    n606, n607, n609, n610, n611, n612, n613, n615, n616, n618, n619, n620,
    n621, n622, n623, n624, n625, n626, n628, n629, n631, n632, n633, n634,
    n635, n636, n637, n639, n640, n642, n643, n644, n645, n646, n647, n648,
    n649, n651, n652, n653, n655, n656, n657, n658, n659, n661, n662, n663,
    n664, n665, n667, n668, n669, n670, n671, n673, n674, n675, n676, n677,
    n679, n680, n681, n682, n683, n685, n686, n687, n688, n690, n691, n692,
    n693, n694, n695, n697, n698, n699, n701, n702, n703, n704, n705, n707,
    n708, n709, n710, n711, n712, n713, n715, n716, n717, n718, n719, n720,
    n722, n723, n724, n726, n727, n728, n729, n730, n732, n733, n734, n735,
    n736, n737, n738, n740, n741, n742, n743, n744, n745, n746, n748, n749,
    n750, n752, n753, n754, n756, n757, n758, n759, n760, n761, n762, n763,
    n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
    n776, n777, n778, n779, n780, n781, n782, n784, n785, n786, n787, n789,
    n791, n793, n795, n797, n799, n801, n803, n805, n807, n809, n811, n813,
    n815, n817, n819, n821, n823, n825, n827, n829, n831, n833, n835, n837,
    n839, n841, n843, n845, n847, n849, n850, n851, n852, n853, n854, n855,
    n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
    n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
    n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
    n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
    n904, n905, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
    n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
    n929, n930, n931, n932, n933, n934, n936, n937, n938, n939, n940, n941,
    n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
    n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
    n966, n967, n968, n970, n971, n972, n973, n974, n975, n976, n977, n978,
    n979, n980, n981, n982, n983, n984, n985, n986, n987, n989, n990, n991,
    n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
    n1003, n1004, n1005, n1006, n1008, n1009, n1010, n1011, n1012, n1013,
    n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
    n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
    n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
    n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
    n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1064,
    n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
    n1075, n1076, n1077, n1078, n1079, n1080, n1082, n1083, n1084, n1085,
    n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
    n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
    n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1116,
    n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
    n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
    n1137, n1138, n1139, n1140, n1141, n1142, n1144, n1145, n1146, n1147,
    n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
    n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
    n1168, n1169, n1170, n1171, n1172, n1174, n1175, n1176, n1177, n1178,
    n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
    n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
    n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
    n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
    n1219, n1220, n1221, n1222, n1224, n1225, n1226, n1227, n1228, n1229,
    n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
    n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
    n1250, n1251, n1252, n1253, n1255, n1256, n1257, n1258, n1259, n1260,
    n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
    n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1280, n1281,
    n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
    n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
    n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
    n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
    n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
    n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
    n1342, n1343, n1344, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
    n1353, n1354, n1355, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
    n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
    n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
    n1384, n1385, n1386, n1387, n1388, n1390, n1391, n1392, n1393, n1394,
    n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
    n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1414, n1415,
    n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
    n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
    n1436, n1437, n1438, n1439, n1441, n1442, n1443, n1444, n1445, n1446,
    n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
    n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
    n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
    n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
    n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1497,
    n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
    n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
    n1518, n1519, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
    n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
    n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
    n1549, n1550, n1551, n1552, n1554, n1555, n1556, n1557, n1558, n1559,
    n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1570,
    n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
    n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
    n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
    n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
    n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
    n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
    n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
    n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1652,
    n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
    n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
    n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
    n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
    n1695, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
    n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
    n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
    n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
    n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1744, n1745, n1746,
    n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
    n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
    n1767, n1768, n1769, n1770, n1772, n1773, n1774, n1775, n1776, n1777,
    n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
    n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1797, n1798,
    n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
    n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1818, n1819,
    n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
    n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
    n1841, n1842, n1843, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
    n1852, n1853, n1854, n1855, n1856, n1857, n1859, n1860, n1861, n1862,
    n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
    n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
    n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1892, n1893,
    n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1903, n1904,
    n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
    n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
    n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1933, n1934, n1935,
    n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
    n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
    n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
    n1966, n1967, n1968, n1969, n1970, n1972, n1973, n1974, n1975, n1976,
    n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
    n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
    n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
    n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2016, n2017,
    n2018, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2029,
    n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
    n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
    n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
    n2060, n2061, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
    n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
    n2081, n2082, n2083, n2084, n2086, n2087, n2088, n2089, n2090, n2091,
    n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
    n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2110, n2111, n2112,
    n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
    n2123, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
    n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
    n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2154, n2155,
    n2156, n2157, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
    n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2177, n2178,
    n2179, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
    n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
    n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2211, n2212,
    n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
    n2223, n2224, n2225, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
    n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
    n2244, n2245, n2246, n2247, n2248, n2254, n2255, n2256, n2257, n2258,
    n2259, n2263, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
    n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2283,
    n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
    n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
    n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
    n2314, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
    n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2338, n2339,
    n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
    n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
    n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2372, n2373,
    n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
    n2384, n2385, n2386, n2388, n2389, n2390, n2392, n2393, n2394, n2395,
    n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
    n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2416,
    n2417, n2420, n2421, n2422, n2423, n2424, n2425, n2427, n2428, n2429,
    n2430, n2431, n2432, n2433, n2434, n2435, n2437, n2438, n2439, n2440,
    n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2451,
    n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2460, n2461, n2462,
    n2464, n2466, n2468, n2470, n2472, n2474, n2476, n2478, n2480, n2482,
    n2484, n2486, n2488, n2490, n2492, n2494, n2496, n2498, n2500, n2502,
    n2504, n2506, n2508, n2510, n2512, n2514, n2516, n2518, n2520, n2522,
    n2524, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
    n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2544, n2545,
    n2546, n2547, n2548, n2549, n2551, n2552, n2553, n2554, n2556, n2557,
    n2558, n2559, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
    n2569, n2570, n2572, n2573, n2574, n2575, n2576, n2578, n2579, n2580,
    n2581, n2583, n2584, n2585, n2586, n2587, n2589, n2590, n2591, n2592,
    n2593, n2594, n2595, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
    n2605, n2606, n2607, n2608, n2609, n2611, n2612, n2613, n2614, n2615,
    n2616, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2626, n2627,
    n2628, n2629, n2630, n2631, n2633, n2634, n2635, n2636, n2637, n2638,
    n2639, n2640, n2642, n2643, n2644, n2645, n2646, n2647, n2649, n2650,
    n2651, n2652, n2653, n2654, n2656, n2657, n2658, n2659, n2660, n2661,
    n2662, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2673,
    n2674, n2675, n2676, n2677, n2678, n2680, n2681, n2682, n2683, n2684,
    n2685, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2695, n2696,
    n2697, n2698, n2699, n2700, n2702, n2703, n2704, n2705, n2706, n2707,
    n2708, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2718, n2719,
    n2720, n2721, n2722, n2723, n2724, n2726, n2727, n2728, n2729, n2730,
    n2731, n2732, n2733, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
    n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2752, n2753,
    n2754, n2755, n2756, n2757, n2758, n2759, n2761, n2762, n2763, n2764,
    n2766, n2767, n2768, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
    n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
    n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
    n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
    n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
    n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
    n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
    n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2845, n2846, n2847,
    n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
    n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
    n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
    n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
    n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
    n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
    n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
    n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
    n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
    n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2947, n2948, n2949,
    n2950, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
    n2961, n2962, n2963, n2965, n2966, n2968, n2969, n2970, n2971, n2972,
    n2973, n2974, n2975, n2976, n2977, n2979, n2980, n2981, n2982, n2983,
    n2984, n2985, n2986, n2987, n2988, n2989, n2991, n2992, n2993, n2994,
    n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3005,
    n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
    n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026,
    n3027, n3028, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
    n3038, n3039, n3040, n3041, n3043, n3044, n3045, n3046, n3047, n3048,
    n3049, n3050, n3051, n3052, n3053, n3054, n3056, n3057, n3058, n3059,
    n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3068, n3069, n3070,
    n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3080, n3081,
    n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
    n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
    n3103, n3104, n3105, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
    n3114, n3115, n3116, n3117, n3118, n3120, n3122, n3123, n3124, n3125,
    n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3136, n3137,
    n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
    n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
    n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
    n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3178,
    n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
    n3189, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
    n3200, n3201, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
    n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3220, n3221,
    n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3231, n3233,
    n3235, n3237, n3239, n3241, n3243, n3245, n3247, n3249, n3251, n3253,
    n3255, n3257, n3259, n3261, n3263, n3265, n3267, n3269, n3271, n3273,
    n3275, n3277, n3279, n3281, n3283, n3285, n3287, n3289, n3291, n3293,
    n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
    n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
    n3315, n3316, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
    n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
    n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
    n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
    n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
    n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
    n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
    n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
    n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
    n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
    n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
    n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
    n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3444, n3445, n3446,
    n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
    n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
    n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
    n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
    n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
    n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
    n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
    n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
    n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
    n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
    n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
    n3557, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
    n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
    n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
    n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
    n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
    n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
    n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
    n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
    n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
    n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
    n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
    n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3679,
    n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
    n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
    n3700, n3701, n3702, n3703, n3704, n3705, n3707, n3708, n3709, n3710,
    n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
    n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
    n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
    n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
    n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
    n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
    n3771, n3772, n3773, n3774, n3776, n3777, n3781, n3782, n3783, n3784,
    n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
    n3795, n3796, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
    n3806, n3807, n3808, n3811, n3812, n3814, n3815, n3816, n3817, n3820,
    n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3833, n3834,
    n3835, n3836, n3837, n3838, n3839, n3840, n3842, n3844, n3845, n3846,
    n3847, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3857, n3858,
    n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3867, n3868, n3869,
    n3870, n3872, n3873, n3874, n3876, n3878, n3881, n3882, n3883, n3884,
    n3885, n3888, n3889, n3890, n3891, n3894, n3895, n3896, n3897, n3899,
    n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
    n3910, n3911, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
    n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
    n3931, n3932, n3933, n3934, n3935, n3937, n3938, n3939, n3940, n3941,
    n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
    n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
    n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
    n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
    n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
    n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
    n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
    n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
    n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
    n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
    n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
    n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
    n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
    n4072, n4073, n4074, n4075, n4077, n4078, n4079, n4080, n4081, n4082,
    n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
    n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
    n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
    n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
    n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
    n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
    n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
    n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
    n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
    n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
    n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
    n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
    n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
    n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4224,
    n4225, n4229, n4230, n4231, n4233, n4234, n4235, n4236, n4238, n4239,
    n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4248, n4249, n4250,
    n4251, n4252, n4253, n4254, n4256, n4257, n4258, n4260, n4261, n4262,
    n4263, n4264, n4265, n4266, n4268, n4269, n4270, n4271, n4272, n4273,
    n4274, n4275, n4276, n4277, n4278, n4279, n4281, n4282, n4283, n4284,
    n4285, n4286, n4287, n4288, n4290, n4291, n4292, n4293, n4294, n4295,
    n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4306,
    n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
    n4317, n4318, n4319, n4320, n4322, n4323, n4324, n4325, n4326, n4327,
    n4328, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4339,
    n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4349, n4350,
    n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4360, n4361,
    n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
    n4372, n4373, n4374, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
    n4383, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
    n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
    n4405, n4407, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416,
    n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
    n4428, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
    n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4449, n4450,
    n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
    n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
    n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4479, n4480, n4481,
    n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4490, n4491, n4492,
    n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4502, n4503,
    n4504, n4505, n4506, n4507, n4508, n4510, n4511, n4512, n4513, n4514,
    n4515, n4516, n4517, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
    n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4536, n4537,
    n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547;
  INVX1   g0000(.A(IR_REG_0__SCAN_IN), .Y(n576));
  NAND2X1 g0001(.A(IR_REG_31__SCAN_IN), .B(STATE_REG_SCAN_IN), .Y(n577));
  INVX1   g0002(.A(STATE_REG_SCAN_IN), .Y(U3149));
  NOR2X1  g0003(.A(IR_REG_31__SCAN_IN), .B(U3149), .Y(n579));
  AOI22X1 g0004(.A0(IR_REG_0__SCAN_IN), .A1(n579), .B0(U3149), .B1(DATAI_0_), .Y(n580));
  OAI21X1 g0005(.A0(n577), .A1(n576), .B0(n580), .Y(U3352));
  XOR2X1  g0006(.A(IR_REG_1__SCAN_IN), .B(n576), .Y(n582));
  AOI22X1 g0007(.A0(IR_REG_1__SCAN_IN), .A1(n579), .B0(U3149), .B1(DATAI_1_), .Y(n583));
  OAI21X1 g0008(.A0(n582), .A1(n577), .B0(n583), .Y(U3351));
  NOR2X1  g0009(.A(IR_REG_1__SCAN_IN), .B(IR_REG_0__SCAN_IN), .Y(n585));
  XOR2X1  g0010(.A(n585), .B(IR_REG_2__SCAN_IN), .Y(n586));
  AOI22X1 g0011(.A0(IR_REG_2__SCAN_IN), .A1(n579), .B0(U3149), .B1(DATAI_2_), .Y(n587));
  OAI21X1 g0012(.A0(n586), .A1(n577), .B0(n587), .Y(U3350));
  NOR3X1  g0013(.A(IR_REG_2__SCAN_IN), .B(IR_REG_1__SCAN_IN), .C(IR_REG_0__SCAN_IN), .Y(n589));
  XOR2X1  g0014(.A(n589), .B(IR_REG_3__SCAN_IN), .Y(n590));
  AOI22X1 g0015(.A0(IR_REG_3__SCAN_IN), .A1(n579), .B0(U3149), .B1(DATAI_3_), .Y(n591));
  OAI21X1 g0016(.A0(n590), .A1(n577), .B0(n591), .Y(U3349));
  NOR4X1  g0017(.A(IR_REG_2__SCAN_IN), .B(IR_REG_1__SCAN_IN), .C(IR_REG_0__SCAN_IN), .D(IR_REG_3__SCAN_IN), .Y(n593));
  XOR2X1  g0018(.A(n593), .B(IR_REG_4__SCAN_IN), .Y(n594));
  AOI22X1 g0019(.A0(IR_REG_4__SCAN_IN), .A1(n579), .B0(U3149), .B1(DATAI_4_), .Y(n595));
  OAI21X1 g0020(.A0(n594), .A1(n577), .B0(n595), .Y(U3348));
  INVX1   g0021(.A(IR_REG_4__SCAN_IN), .Y(n597));
  NAND2X1 g0022(.A(n593), .B(n597), .Y(n598));
  NAND2X1 g0023(.A(n598), .B(IR_REG_5__SCAN_IN), .Y(n599));
  NOR3X1  g0024(.A(IR_REG_5__SCAN_IN), .B(IR_REG_4__SCAN_IN), .C(IR_REG_3__SCAN_IN), .Y(n600));
  NAND2X1 g0025(.A(n600), .B(n589), .Y(n601));
  NAND2X1 g0026(.A(n601), .B(n599), .Y(n602));
  AOI22X1 g0027(.A0(IR_REG_5__SCAN_IN), .A1(n579), .B0(U3149), .B1(DATAI_5_), .Y(n603));
  OAI21X1 g0028(.A0(n602), .A1(n577), .B0(n603), .Y(U3347));
  INVX1   g0029(.A(IR_REG_6__SCAN_IN), .Y(n605));
  XOR2X1  g0030(.A(n601), .B(n605), .Y(n606));
  AOI22X1 g0031(.A0(IR_REG_6__SCAN_IN), .A1(n579), .B0(U3149), .B1(DATAI_6_), .Y(n607));
  OAI21X1 g0032(.A0(n606), .A1(n577), .B0(n607), .Y(U3346));
  NAND3X1 g0033(.A(n600), .B(n589), .C(n605), .Y(n609));
  NOR3X1  g0034(.A(n601), .B(IR_REG_7__SCAN_IN), .C(IR_REG_6__SCAN_IN), .Y(n610));
  AOI21X1 g0035(.A0(n609), .A1(IR_REG_7__SCAN_IN), .B0(n610), .Y(n611));
  NAND3X1 g0036(.A(n611), .B(IR_REG_31__SCAN_IN), .C(STATE_REG_SCAN_IN), .Y(n612));
  AOI22X1 g0037(.A0(IR_REG_7__SCAN_IN), .A1(n579), .B0(U3149), .B1(DATAI_7_), .Y(n613));
  NAND2X1 g0038(.A(n613), .B(n612), .Y(U3345));
  XOR2X1  g0039(.A(n610), .B(IR_REG_8__SCAN_IN), .Y(n615));
  AOI22X1 g0040(.A0(IR_REG_8__SCAN_IN), .A1(n579), .B0(U3149), .B1(DATAI_8_), .Y(n616));
  OAI21X1 g0041(.A0(n615), .A1(n577), .B0(n616), .Y(U3344));
  INVX1   g0042(.A(IR_REG_8__SCAN_IN), .Y(n618));
  NOR2X1  g0043(.A(IR_REG_7__SCAN_IN), .B(IR_REG_6__SCAN_IN), .Y(n619));
  NAND4X1 g0044(.A(n600), .B(n589), .C(n618), .D(n619), .Y(n620));
  INVX1   g0045(.A(IR_REG_9__SCAN_IN), .Y(n621));
  NAND3X1 g0046(.A(n619), .B(n621), .C(n618), .Y(n622));
  NOR2X1  g0047(.A(n622), .B(n601), .Y(n623));
  AOI21X1 g0048(.A0(n620), .A1(IR_REG_9__SCAN_IN), .B0(n623), .Y(n624));
  NAND3X1 g0049(.A(n624), .B(IR_REG_31__SCAN_IN), .C(STATE_REG_SCAN_IN), .Y(n625));
  AOI22X1 g0050(.A0(IR_REG_9__SCAN_IN), .A1(n579), .B0(U3149), .B1(DATAI_9_), .Y(n626));
  NAND2X1 g0051(.A(n626), .B(n625), .Y(U3343));
  XOR2X1  g0052(.A(n623), .B(IR_REG_10__SCAN_IN), .Y(n628));
  AOI22X1 g0053(.A0(IR_REG_10__SCAN_IN), .A1(n579), .B0(U3149), .B1(DATAI_10_), .Y(n629));
  OAI21X1 g0054(.A0(n628), .A1(n577), .B0(n629), .Y(U3342));
  INVX1   g0055(.A(IR_REG_10__SCAN_IN), .Y(n631));
  INVX1   g0056(.A(IR_REG_11__SCAN_IN), .Y(n632));
  AOI21X1 g0057(.A0(n623), .A1(n631), .B0(n632), .Y(n633));
  NOR4X1  g0058(.A(n601), .B(IR_REG_11__SCAN_IN), .C(IR_REG_10__SCAN_IN), .D(n622), .Y(n634));
  NOR2X1  g0059(.A(n634), .B(n633), .Y(n635));
  NAND3X1 g0060(.A(n635), .B(IR_REG_31__SCAN_IN), .C(STATE_REG_SCAN_IN), .Y(n636));
  AOI22X1 g0061(.A0(IR_REG_11__SCAN_IN), .A1(n579), .B0(U3149), .B1(DATAI_11_), .Y(n637));
  NAND2X1 g0062(.A(n637), .B(n636), .Y(U3341));
  XOR2X1  g0063(.A(n634), .B(IR_REG_12__SCAN_IN), .Y(n639));
  AOI22X1 g0064(.A0(IR_REG_12__SCAN_IN), .A1(n579), .B0(U3149), .B1(DATAI_12_), .Y(n640));
  OAI21X1 g0065(.A0(n639), .A1(n577), .B0(n640), .Y(U3340));
  INVX1   g0066(.A(IR_REG_13__SCAN_IN), .Y(n642));
  NAND2X1 g0067(.A(n632), .B(n631), .Y(n643));
  NOR4X1  g0068(.A(n622), .B(n601), .C(IR_REG_12__SCAN_IN), .D(n643), .Y(n644));
  NOR4X1  g0069(.A(IR_REG_9__SCAN_IN), .B(IR_REG_8__SCAN_IN), .C(IR_REG_7__SCAN_IN), .D(IR_REG_12__SCAN_IN), .Y(n645));
  NOR4X1  g0070(.A(IR_REG_11__SCAN_IN), .B(IR_REG_10__SCAN_IN), .C(IR_REG_6__SCAN_IN), .D(IR_REG_13__SCAN_IN), .Y(n646));
  NAND4X1 g0071(.A(n645), .B(n600), .C(n589), .D(n646), .Y(n647));
  OAI21X1 g0072(.A0(n644), .A1(n642), .B0(n647), .Y(n648));
  AOI22X1 g0073(.A0(IR_REG_13__SCAN_IN), .A1(n579), .B0(U3149), .B1(DATAI_13_), .Y(n649));
  OAI21X1 g0074(.A0(n648), .A1(n577), .B0(n649), .Y(U3339));
  INVX1   g0075(.A(IR_REG_14__SCAN_IN), .Y(n651));
  XOR2X1  g0076(.A(n647), .B(n651), .Y(n652));
  AOI22X1 g0077(.A0(IR_REG_14__SCAN_IN), .A1(n579), .B0(U3149), .B1(DATAI_14_), .Y(n653));
  OAI21X1 g0078(.A0(n652), .A1(n577), .B0(n653), .Y(U3338));
  OAI21X1 g0079(.A0(n647), .A1(IR_REG_14__SCAN_IN), .B0(IR_REG_15__SCAN_IN), .Y(n655));
  INVX1   g0080(.A(IR_REG_15__SCAN_IN), .Y(n656));
  NAND2X1 g0081(.A(n656), .B(n651), .Y(n657));
  OAI21X1 g0082(.A0(n657), .A1(n647), .B0(n655), .Y(n658));
  AOI22X1 g0083(.A0(IR_REG_15__SCAN_IN), .A1(n579), .B0(U3149), .B1(DATAI_15_), .Y(n659));
  OAI21X1 g0084(.A0(n658), .A1(n577), .B0(n659), .Y(U3337));
  INVX1   g0085(.A(IR_REG_16__SCAN_IN), .Y(n661));
  NOR2X1  g0086(.A(n657), .B(n647), .Y(n662));
  XOR2X1  g0087(.A(n662), .B(n661), .Y(n663));
  NAND3X1 g0088(.A(n663), .B(IR_REG_31__SCAN_IN), .C(STATE_REG_SCAN_IN), .Y(n664));
  AOI22X1 g0089(.A0(IR_REG_16__SCAN_IN), .A1(n579), .B0(U3149), .B1(DATAI_16_), .Y(n665));
  NAND2X1 g0090(.A(n665), .B(n664), .Y(U3336));
  INVX1   g0091(.A(IR_REG_17__SCAN_IN), .Y(n667));
  NOR3X1  g0092(.A(n657), .B(n647), .C(IR_REG_16__SCAN_IN), .Y(n668));
  NAND4X1 g0093(.A(n661), .B(n656), .C(n651), .D(n667), .Y(n669));
  OAI22X1 g0094(.A0(n668), .A1(n667), .B0(n647), .B1(n669), .Y(n670));
  AOI22X1 g0095(.A0(IR_REG_17__SCAN_IN), .A1(n579), .B0(U3149), .B1(DATAI_17_), .Y(n671));
  OAI21X1 g0096(.A0(n670), .A1(n577), .B0(n671), .Y(U3335));
  INVX1   g0097(.A(IR_REG_18__SCAN_IN), .Y(n673));
  NOR2X1  g0098(.A(n669), .B(n647), .Y(n674));
  XOR2X1  g0099(.A(n674), .B(n673), .Y(n675));
  NAND3X1 g0100(.A(n675), .B(IR_REG_31__SCAN_IN), .C(STATE_REG_SCAN_IN), .Y(n676));
  AOI22X1 g0101(.A0(IR_REG_18__SCAN_IN), .A1(n579), .B0(U3149), .B1(DATAI_18_), .Y(n677));
  NAND2X1 g0102(.A(n677), .B(n676), .Y(U3334));
  INVX1   g0103(.A(IR_REG_19__SCAN_IN), .Y(n679));
  NOR3X1  g0104(.A(n669), .B(n647), .C(IR_REG_18__SCAN_IN), .Y(n680));
  NAND3X1 g0105(.A(n674), .B(n679), .C(n673), .Y(n681));
  OAI21X1 g0106(.A0(n680), .A1(n679), .B0(n681), .Y(n682));
  AOI22X1 g0107(.A0(IR_REG_19__SCAN_IN), .A1(n579), .B0(U3149), .B1(DATAI_19_), .Y(n683));
  OAI21X1 g0108(.A0(n682), .A1(n577), .B0(n683), .Y(U3333));
  NAND2X1 g0109(.A(n679), .B(n673), .Y(n685));
  NOR3X1  g0110(.A(n685), .B(n669), .C(n647), .Y(n686));
  XOR2X1  g0111(.A(n686), .B(IR_REG_20__SCAN_IN), .Y(n687));
  AOI22X1 g0112(.A0(IR_REG_20__SCAN_IN), .A1(n579), .B0(U3149), .B1(DATAI_20_), .Y(n688));
  OAI21X1 g0113(.A0(n687), .A1(n577), .B0(n688), .Y(U3332));
  INVX1   g0114(.A(IR_REG_21__SCAN_IN), .Y(n690));
  NOR4X1  g0115(.A(n669), .B(n647), .C(IR_REG_20__SCAN_IN), .D(n685), .Y(n691));
  INVX1   g0116(.A(IR_REG_20__SCAN_IN), .Y(n692));
  NAND2X1 g0117(.A(n690), .B(n692), .Y(n693));
  OAI22X1 g0118(.A0(n691), .A1(n690), .B0(n681), .B1(n693), .Y(n694));
  AOI22X1 g0119(.A0(IR_REG_21__SCAN_IN), .A1(n579), .B0(U3149), .B1(DATAI_21_), .Y(n695));
  OAI21X1 g0120(.A0(n694), .A1(n577), .B0(n695), .Y(U3331));
  NOR4X1  g0121(.A(n685), .B(n669), .C(n647), .D(n693), .Y(n697));
  XOR2X1  g0122(.A(n697), .B(IR_REG_22__SCAN_IN), .Y(n698));
  AOI22X1 g0123(.A0(IR_REG_22__SCAN_IN), .A1(n579), .B0(U3149), .B1(DATAI_22_), .Y(n699));
  OAI21X1 g0124(.A0(n698), .A1(n577), .B0(n699), .Y(U3330));
  INVX1   g0125(.A(IR_REG_22__SCAN_IN), .Y(n701));
  NAND2X1 g0126(.A(n697), .B(n701), .Y(n702));
  XOR2X1  g0127(.A(n702), .B(IR_REG_23__SCAN_IN), .Y(n703));
  INVX1   g0128(.A(n703), .Y(n704));
  AOI22X1 g0129(.A0(IR_REG_23__SCAN_IN), .A1(n579), .B0(U3149), .B1(DATAI_23_), .Y(n705));
  OAI21X1 g0130(.A0(n704), .A1(n577), .B0(n705), .Y(U3329));
  INVX1   g0131(.A(IR_REG_23__SCAN_IN), .Y(n707));
  NOR4X1  g0132(.A(IR_REG_16__SCAN_IN), .B(IR_REG_15__SCAN_IN), .C(IR_REG_14__SCAN_IN), .D(IR_REG_17__SCAN_IN), .Y(n708));
  NOR4X1  g0133(.A(IR_REG_20__SCAN_IN), .B(IR_REG_19__SCAN_IN), .C(IR_REG_18__SCAN_IN), .D(IR_REG_21__SCAN_IN), .Y(n709));
  NAND4X1 g0134(.A(n708), .B(n707), .C(n701), .D(n709), .Y(n710));
  NOR2X1  g0135(.A(n710), .B(n647), .Y(n711));
  XOR2X1  g0136(.A(n711), .B(IR_REG_24__SCAN_IN), .Y(n712));
  AOI22X1 g0137(.A0(IR_REG_24__SCAN_IN), .A1(n579), .B0(U3149), .B1(DATAI_24_), .Y(n713));
  OAI21X1 g0138(.A0(n712), .A1(n577), .B0(n713), .Y(U3328));
  INVX1   g0139(.A(IR_REG_25__SCAN_IN), .Y(n715));
  NOR3X1  g0140(.A(n710), .B(n647), .C(IR_REG_24__SCAN_IN), .Y(n716));
  INVX1   g0141(.A(IR_REG_24__SCAN_IN), .Y(n717));
  NAND3X1 g0142(.A(n711), .B(n715), .C(n717), .Y(n718));
  OAI21X1 g0143(.A0(n716), .A1(n715), .B0(n718), .Y(n719));
  AOI22X1 g0144(.A0(IR_REG_25__SCAN_IN), .A1(n579), .B0(U3149), .B1(DATAI_25_), .Y(n720));
  OAI21X1 g0145(.A0(n719), .A1(n577), .B0(n720), .Y(U3327));
  NOR4X1  g0146(.A(n647), .B(IR_REG_25__SCAN_IN), .C(IR_REG_24__SCAN_IN), .D(n710), .Y(n722));
  XOR2X1  g0147(.A(n722), .B(IR_REG_26__SCAN_IN), .Y(n723));
  AOI22X1 g0148(.A0(IR_REG_26__SCAN_IN), .A1(n579), .B0(U3149), .B1(DATAI_26_), .Y(n724));
  OAI21X1 g0149(.A0(n723), .A1(n577), .B0(n724), .Y(U3326));
  INVX1   g0150(.A(IR_REG_27__SCAN_IN), .Y(n726));
  INVX1   g0151(.A(IR_REG_26__SCAN_IN), .Y(n727));
  NAND2X1 g0152(.A(n722), .B(n727), .Y(n728));
  XOR2X1  g0153(.A(n728), .B(n726), .Y(n729));
  AOI22X1 g0154(.A0(IR_REG_27__SCAN_IN), .A1(n579), .B0(U3149), .B1(DATAI_27_), .Y(n730));
  OAI21X1 g0155(.A0(n729), .A1(n577), .B0(n730), .Y(U3325));
  INVX1   g0156(.A(IR_REG_28__SCAN_IN), .Y(n732));
  NAND4X1 g0157(.A(n727), .B(n715), .C(n717), .D(n726), .Y(n733));
  NOR3X1  g0158(.A(n733), .B(n710), .C(n647), .Y(n734));
  NOR4X1  g0159(.A(n710), .B(n647), .C(IR_REG_28__SCAN_IN), .D(n733), .Y(n735));
  INVX1   g0160(.A(n735), .Y(n736));
  OAI21X1 g0161(.A0(n734), .A1(n732), .B0(n736), .Y(n737));
  AOI22X1 g0162(.A0(IR_REG_28__SCAN_IN), .A1(n579), .B0(U3149), .B1(DATAI_28_), .Y(n738));
  OAI21X1 g0163(.A0(n737), .A1(n577), .B0(n738), .Y(U3324));
  INVX1   g0164(.A(IR_REG_29__SCAN_IN), .Y(n740));
  NOR2X1  g0165(.A(n733), .B(n647), .Y(n741));
  NAND2X1 g0166(.A(n740), .B(n732), .Y(n742));
  NOR2X1  g0167(.A(n742), .B(n710), .Y(n743));
  NAND2X1 g0168(.A(n743), .B(n741), .Y(n744));
  OAI21X1 g0169(.A0(n735), .A1(n740), .B0(n744), .Y(n745));
  AOI22X1 g0170(.A0(IR_REG_29__SCAN_IN), .A1(n579), .B0(U3149), .B1(DATAI_29_), .Y(n746));
  OAI21X1 g0171(.A0(n745), .A1(n577), .B0(n746), .Y(U3323));
  NOR4X1  g0172(.A(n733), .B(n710), .C(n647), .D(n742), .Y(n748));
  XOR2X1  g0173(.A(n748), .B(IR_REG_30__SCAN_IN), .Y(n749));
  AOI22X1 g0174(.A0(IR_REG_30__SCAN_IN), .A1(n579), .B0(U3149), .B1(DATAI_30_), .Y(n750));
  OAI21X1 g0175(.A0(n749), .A1(n577), .B0(n750), .Y(U3322));
  INVX1   g0176(.A(IR_REG_30__SCAN_IN), .Y(n752));
  NAND4X1 g0177(.A(IR_REG_31__SCAN_IN), .B(n752), .C(STATE_REG_SCAN_IN), .D(n748), .Y(n753));
  NAND2X1 g0178(.A(U3149), .B(DATAI_31_), .Y(n754));
  NAND2X1 g0179(.A(n754), .B(n753), .Y(U3321));
  NOR2X1  g0180(.A(IR_REG_31__SCAN_IN), .B(n707), .Y(n756));
  AOI21X1 g0181(.A0(n703), .A1(IR_REG_31__SCAN_IN), .B0(n756), .Y(n757));
  INVX1   g0182(.A(n757), .Y(n758));
  INVX1   g0183(.A(IR_REG_31__SCAN_IN), .Y(n759));
  NOR2X1  g0184(.A(n716), .B(n715), .Y(n760));
  NOR3X1  g0185(.A(n722), .B(n760), .C(n759), .Y(n761));
  AOI21X1 g0186(.A0(n759), .A1(IR_REG_25__SCAN_IN), .B0(n761), .Y(n762));
  NOR2X1  g0187(.A(n712), .B(n759), .Y(n763));
  AOI21X1 g0188(.A0(n759), .A1(IR_REG_24__SCAN_IN), .B0(n763), .Y(n764));
  NOR2X1  g0189(.A(n723), .B(n759), .Y(n765));
  AOI21X1 g0190(.A0(n759), .A1(IR_REG_26__SCAN_IN), .B0(n765), .Y(n766));
  NOR3X1  g0191(.A(n766), .B(n764), .C(n762), .Y(n767));
  NOR3X1  g0192(.A(n767), .B(n758), .C(U3149), .Y(n768));
  INVX1   g0193(.A(n768), .Y(n769));
  NAND2X1 g0194(.A(n759), .B(IR_REG_26__SCAN_IN), .Y(n770));
  OAI21X1 g0195(.A0(n723), .A1(n759), .B0(n770), .Y(n771));
  NAND4X1 g0196(.A(n764), .B(n762), .C(B_REG_SCAN_IN), .D(n771), .Y(n772));
  INVX1   g0197(.A(B_REG_SCAN_IN), .Y(n773));
  NAND2X1 g0198(.A(n759), .B(IR_REG_24__SCAN_IN), .Y(n774));
  OAI21X1 g0199(.A0(n712), .A1(n759), .B0(n774), .Y(n775));
  AOI21X1 g0200(.A0(n775), .A1(n773), .B0(n766), .Y(n776));
  NAND2X1 g0201(.A(n776), .B(n772), .Y(n777));
  INVX1   g0202(.A(n777), .Y(n778));
  NOR2X1  g0203(.A(n778), .B(n769), .Y(n779));
  INVX1   g0204(.A(n779), .Y(n780));
  AOI21X1 g0205(.A0(n771), .A1(n762), .B0(n775), .Y(n781));
  OAI21X1 g0206(.A0(n778), .A1(n769), .B0(D_REG_0__SCAN_IN), .Y(n782));
  OAI21X1 g0207(.A0(n781), .A1(n780), .B0(n782), .Y(U3458));
  NAND2X1 g0208(.A(n759), .B(IR_REG_25__SCAN_IN), .Y(n784));
  OAI21X1 g0209(.A0(n719), .A1(n759), .B0(n784), .Y(n785));
  NOR2X1  g0210(.A(n771), .B(n785), .Y(n786));
  OAI21X1 g0211(.A0(n778), .A1(n769), .B0(D_REG_1__SCAN_IN), .Y(n787));
  OAI21X1 g0212(.A0(n786), .A1(n780), .B0(n787), .Y(U3459));
  INVX1   g0213(.A(D_REG_2__SCAN_IN), .Y(n789));
  AOI21X1 g0214(.A0(n777), .A1(n768), .B0(n789), .Y(U3320));
  INVX1   g0215(.A(D_REG_3__SCAN_IN), .Y(n791));
  AOI21X1 g0216(.A0(n777), .A1(n768), .B0(n791), .Y(U3319));
  INVX1   g0217(.A(D_REG_4__SCAN_IN), .Y(n793));
  AOI21X1 g0218(.A0(n777), .A1(n768), .B0(n793), .Y(U3318));
  INVX1   g0219(.A(D_REG_5__SCAN_IN), .Y(n795));
  AOI21X1 g0220(.A0(n777), .A1(n768), .B0(n795), .Y(U3317));
  INVX1   g0221(.A(D_REG_6__SCAN_IN), .Y(n797));
  AOI21X1 g0222(.A0(n777), .A1(n768), .B0(n797), .Y(U3316));
  INVX1   g0223(.A(D_REG_7__SCAN_IN), .Y(n799));
  AOI21X1 g0224(.A0(n777), .A1(n768), .B0(n799), .Y(U3315));
  INVX1   g0225(.A(D_REG_8__SCAN_IN), .Y(n801));
  AOI21X1 g0226(.A0(n777), .A1(n768), .B0(n801), .Y(U3314));
  INVX1   g0227(.A(D_REG_9__SCAN_IN), .Y(n803));
  AOI21X1 g0228(.A0(n777), .A1(n768), .B0(n803), .Y(U3313));
  INVX1   g0229(.A(D_REG_10__SCAN_IN), .Y(n805));
  AOI21X1 g0230(.A0(n777), .A1(n768), .B0(n805), .Y(U3312));
  INVX1   g0231(.A(D_REG_11__SCAN_IN), .Y(n807));
  AOI21X1 g0232(.A0(n777), .A1(n768), .B0(n807), .Y(U3311));
  INVX1   g0233(.A(D_REG_12__SCAN_IN), .Y(n809));
  AOI21X1 g0234(.A0(n777), .A1(n768), .B0(n809), .Y(U3310));
  INVX1   g0235(.A(D_REG_13__SCAN_IN), .Y(n811));
  AOI21X1 g0236(.A0(n777), .A1(n768), .B0(n811), .Y(U3309));
  INVX1   g0237(.A(D_REG_14__SCAN_IN), .Y(n813));
  AOI21X1 g0238(.A0(n777), .A1(n768), .B0(n813), .Y(U3308));
  INVX1   g0239(.A(D_REG_15__SCAN_IN), .Y(n815));
  AOI21X1 g0240(.A0(n777), .A1(n768), .B0(n815), .Y(U3307));
  INVX1   g0241(.A(D_REG_16__SCAN_IN), .Y(n817));
  AOI21X1 g0242(.A0(n777), .A1(n768), .B0(n817), .Y(U3306));
  INVX1   g0243(.A(D_REG_17__SCAN_IN), .Y(n819));
  AOI21X1 g0244(.A0(n777), .A1(n768), .B0(n819), .Y(U3305));
  INVX1   g0245(.A(D_REG_18__SCAN_IN), .Y(n821));
  AOI21X1 g0246(.A0(n777), .A1(n768), .B0(n821), .Y(U3304));
  INVX1   g0247(.A(D_REG_19__SCAN_IN), .Y(n823));
  AOI21X1 g0248(.A0(n777), .A1(n768), .B0(n823), .Y(U3303));
  INVX1   g0249(.A(D_REG_20__SCAN_IN), .Y(n825));
  AOI21X1 g0250(.A0(n777), .A1(n768), .B0(n825), .Y(U3302));
  INVX1   g0251(.A(D_REG_21__SCAN_IN), .Y(n827));
  AOI21X1 g0252(.A0(n777), .A1(n768), .B0(n827), .Y(U3301));
  INVX1   g0253(.A(D_REG_22__SCAN_IN), .Y(n829));
  AOI21X1 g0254(.A0(n777), .A1(n768), .B0(n829), .Y(U3300));
  INVX1   g0255(.A(D_REG_23__SCAN_IN), .Y(n831));
  AOI21X1 g0256(.A0(n777), .A1(n768), .B0(n831), .Y(U3299));
  INVX1   g0257(.A(D_REG_24__SCAN_IN), .Y(n833));
  AOI21X1 g0258(.A0(n777), .A1(n768), .B0(n833), .Y(U3298));
  INVX1   g0259(.A(D_REG_25__SCAN_IN), .Y(n835));
  AOI21X1 g0260(.A0(n777), .A1(n768), .B0(n835), .Y(U3297));
  INVX1   g0261(.A(D_REG_26__SCAN_IN), .Y(n837));
  AOI21X1 g0262(.A0(n777), .A1(n768), .B0(n837), .Y(U3296));
  INVX1   g0263(.A(D_REG_27__SCAN_IN), .Y(n839));
  AOI21X1 g0264(.A0(n777), .A1(n768), .B0(n839), .Y(U3295));
  INVX1   g0265(.A(D_REG_28__SCAN_IN), .Y(n841));
  AOI21X1 g0266(.A0(n777), .A1(n768), .B0(n841), .Y(U3294));
  INVX1   g0267(.A(D_REG_29__SCAN_IN), .Y(n843));
  AOI21X1 g0268(.A0(n777), .A1(n768), .B0(n843), .Y(U3293));
  INVX1   g0269(.A(D_REG_30__SCAN_IN), .Y(n845));
  AOI21X1 g0270(.A0(n777), .A1(n768), .B0(n845), .Y(U3292));
  INVX1   g0271(.A(D_REG_31__SCAN_IN), .Y(n847));
  AOI21X1 g0272(.A0(n777), .A1(n768), .B0(n847), .Y(U3291));
  OAI21X1 g0273(.A0(D_REG_7__SCAN_IN), .A1(D_REG_3__SCAN_IN), .B0(n778), .Y(n849));
  OAI21X1 g0274(.A0(D_REG_9__SCAN_IN), .A1(D_REG_8__SCAN_IN), .B0(n778), .Y(n850));
  OAI21X1 g0275(.A0(D_REG_10__SCAN_IN), .A1(D_REG_5__SCAN_IN), .B0(n778), .Y(n851));
  OAI21X1 g0276(.A0(D_REG_6__SCAN_IN), .A1(D_REG_4__SCAN_IN), .B0(n778), .Y(n852));
  NAND4X1 g0277(.A(n851), .B(n850), .C(n849), .D(n852), .Y(n853));
  OAI21X1 g0278(.A0(D_REG_28__SCAN_IN), .A1(D_REG_27__SCAN_IN), .B0(n778), .Y(n854));
  OAI21X1 g0279(.A0(D_REG_26__SCAN_IN), .A1(D_REG_25__SCAN_IN), .B0(n778), .Y(n855));
  OAI21X1 g0280(.A0(D_REG_31__SCAN_IN), .A1(D_REG_30__SCAN_IN), .B0(n778), .Y(n856));
  OAI21X1 g0281(.A0(D_REG_29__SCAN_IN), .A1(D_REG_2__SCAN_IN), .B0(n778), .Y(n857));
  NAND4X1 g0282(.A(n856), .B(n855), .C(n854), .D(n857), .Y(n858));
  OAI21X1 g0283(.A0(D_REG_21__SCAN_IN), .A1(D_REG_20__SCAN_IN), .B0(n778), .Y(n859));
  OAI21X1 g0284(.A0(D_REG_19__SCAN_IN), .A1(D_REG_18__SCAN_IN), .B0(n778), .Y(n860));
  OAI21X1 g0285(.A0(D_REG_23__SCAN_IN), .A1(D_REG_22__SCAN_IN), .B0(n778), .Y(n861));
  AOI21X1 g0286(.A0(n813), .A1(n809), .B0(n777), .Y(n862));
  AOI21X1 g0287(.A0(n811), .A1(n807), .B0(n777), .Y(n863));
  AOI21X1 g0288(.A0(n833), .A1(n817), .B0(n777), .Y(n864));
  AOI21X1 g0289(.A0(n819), .A1(n815), .B0(n777), .Y(n865));
  NOR4X1  g0290(.A(n864), .B(n863), .C(n862), .D(n865), .Y(n866));
  NAND4X1 g0291(.A(n861), .B(n860), .C(n859), .D(n866), .Y(n867));
  NOR3X1  g0292(.A(n867), .B(n858), .C(n853), .Y(n868));
  AOI21X1 g0293(.A0(n776), .A1(n772), .B0(n786), .Y(n869));
  AOI21X1 g0294(.A0(n778), .A1(D_REG_1__SCAN_IN), .B0(n869), .Y(n870));
  NOR2X1  g0295(.A(n691), .B(n690), .Y(n871));
  NOR3X1  g0296(.A(n697), .B(n871), .C(n759), .Y(n872));
  AOI21X1 g0297(.A0(n759), .A1(IR_REG_21__SCAN_IN), .B0(n872), .Y(n873));
  NOR2X1  g0298(.A(IR_REG_31__SCAN_IN), .B(n701), .Y(n874));
  INVX1   g0299(.A(n874), .Y(n875));
  OAI21X1 g0300(.A0(n698), .A1(n759), .B0(n875), .Y(n876));
  NOR2X1  g0301(.A(n687), .B(n759), .Y(n877));
  AOI21X1 g0302(.A0(n759), .A1(IR_REG_20__SCAN_IN), .B0(n877), .Y(n878));
  NOR2X1  g0303(.A(n680), .B(n679), .Y(n879));
  NOR3X1  g0304(.A(n686), .B(n879), .C(n759), .Y(n880));
  AOI21X1 g0305(.A0(n759), .A1(IR_REG_19__SCAN_IN), .B0(n880), .Y(n881));
  AOI22X1 g0306(.A0(n878), .A1(n881), .B0(n876), .B1(n873), .Y(n882));
  NAND2X1 g0307(.A(n759), .B(IR_REG_21__SCAN_IN), .Y(n883));
  OAI21X1 g0308(.A0(n694), .A1(n759), .B0(n883), .Y(n884));
  XOR2X1  g0309(.A(n697), .B(n701), .Y(n885));
  AOI21X1 g0310(.A0(n885), .A1(IR_REG_31__SCAN_IN), .B0(n874), .Y(n886));
  NAND2X1 g0311(.A(n886), .B(n884), .Y(n887));
  NAND2X1 g0312(.A(n759), .B(IR_REG_20__SCAN_IN), .Y(n888));
  OAI21X1 g0313(.A0(n687), .A1(n759), .B0(n888), .Y(n889));
  NAND2X1 g0314(.A(n889), .B(n873), .Y(n890));
  NAND3X1 g0315(.A(n890), .B(n887), .C(n882), .Y(n891));
  AOI22X1 g0316(.A0(n772), .A1(n776), .B0(n766), .B1(n764), .Y(n892));
  AOI21X1 g0317(.A0(n778), .A1(D_REG_0__SCAN_IN), .B0(n892), .Y(n893));
  INVX1   g0318(.A(n893), .Y(n894));
  NOR2X1  g0319(.A(n894), .B(n769), .Y(n895));
  NAND4X1 g0320(.A(n891), .B(n870), .C(n868), .D(n895), .Y(n896));
  INVX1   g0321(.A(DATAI_0_), .Y(n897));
  NAND2X1 g0322(.A(n759), .B(IR_REG_27__SCAN_IN), .Y(n898));
  OAI21X1 g0323(.A0(n729), .A1(n759), .B0(n898), .Y(n899));
  NOR2X1  g0324(.A(n737), .B(n759), .Y(n900));
  NOR2X1  g0325(.A(IR_REG_31__SCAN_IN), .B(n732), .Y(n901));
  NOR3X1  g0326(.A(n901), .B(n900), .C(n899), .Y(n902));
  NAND2X1 g0327(.A(IR_REG_31__SCAN_IN), .B(IR_REG_0__SCAN_IN), .Y(n903));
  INVX1   g0328(.A(n903), .Y(n904));
  NOR2X1  g0329(.A(IR_REG_31__SCAN_IN), .B(n576), .Y(n905));
  INVX1   g0330(.A(n576), .Y(n907));
  NAND2X1 g0331(.A(n907), .B(n902), .Y(n908));
  OAI21X1 g0332(.A0(n902), .A1(n897), .B0(n908), .Y(n909));
  INVX1   g0333(.A(REG2_REG_0__SCAN_IN), .Y(n910));
  NOR2X1  g0334(.A(IR_REG_31__SCAN_IN), .B(n752), .Y(n911));
  INVX1   g0335(.A(n911), .Y(n912));
  OAI21X1 g0336(.A0(n749), .A1(n759), .B0(n912), .Y(n913));
  NOR2X1  g0337(.A(n735), .B(n740), .Y(n914));
  NOR3X1  g0338(.A(n748), .B(n914), .C(n759), .Y(n915));
  NOR2X1  g0339(.A(IR_REG_31__SCAN_IN), .B(n740), .Y(n916));
  NOR3X1  g0340(.A(n916), .B(n915), .C(n913), .Y(n917));
  NAND2X1 g0341(.A(n917), .B(REG0_REG_0__SCAN_IN), .Y(n918));
  NOR2X1  g0342(.A(n916), .B(n915), .Y(n919));
  NAND2X1 g0343(.A(n919), .B(n913), .Y(n920));
  OAI21X1 g0344(.A0(n920), .A1(n910), .B0(n918), .Y(n921));
  INVX1   g0345(.A(REG3_REG_0__SCAN_IN), .Y(n922));
  INVX1   g0346(.A(REG1_REG_0__SCAN_IN), .Y(n923));
  XOR2X1  g0347(.A(n748), .B(n752), .Y(n924));
  AOI21X1 g0348(.A0(n924), .A1(IR_REG_31__SCAN_IN), .B0(n911), .Y(n925));
  OAI21X1 g0349(.A0(n916), .A1(n915), .B0(n925), .Y(n926));
  OAI21X1 g0350(.A0(n916), .A1(n915), .B0(n913), .Y(n927));
  OAI22X1 g0351(.A0(n926), .A1(n923), .B0(n922), .B1(n927), .Y(n928));
  NOR2X1  g0352(.A(n928), .B(n921), .Y(n929));
  XOR2X1  g0353(.A(n929), .B(n909), .Y(n930));
  NOR3X1  g0354(.A(n881), .B(n889), .C(n886), .Y(n931));
  INVX1   g0355(.A(n931), .Y(n932));
  NOR2X1  g0356(.A(n932), .B(n930), .Y(n933));
  INVX1   g0357(.A(n933), .Y(n934));
  NOR3X1  g0358(.A(n881), .B(n878), .C(n873), .Y(n936));
  NAND2X1 g0359(.A(n759), .B(IR_REG_19__SCAN_IN), .Y(n937));
  OAI21X1 g0360(.A0(n682), .A1(n759), .B0(n937), .Y(n938));
  NOR3X1  g0361(.A(n938), .B(n878), .C(n886), .Y(n939));
  OAI21X1 g0362(.A0(n939), .A1(n936), .B0(n3791), .Y(n940));
  NOR3X1  g0363(.A(n881), .B(n878), .C(n886), .Y(n941));
  NAND3X1 g0364(.A(n881), .B(n889), .C(n884), .Y(n942));
  INVX1   g0365(.A(n942), .Y(n943));
  OAI21X1 g0366(.A0(n943), .A1(n941), .B0(n3791), .Y(n944));
  NOR4X1  g0367(.A(n889), .B(n876), .C(n873), .D(n938), .Y(n945));
  NOR4X1  g0368(.A(n889), .B(n886), .C(n884), .D(n938), .Y(n946));
  OAI21X1 g0369(.A0(n946), .A1(n945), .B0(n3791), .Y(n947));
  NAND4X1 g0370(.A(n944), .B(n940), .C(n934), .D(n947), .Y(n948));
  NOR3X1  g0371(.A(n881), .B(n889), .C(n876), .Y(n949));
  INVX1   g0372(.A(n949), .Y(n950));
  NOR4X1  g0373(.A(n900), .B(n886), .C(n873), .D(n901), .Y(n951));
  NOR3X1  g0374(.A(n916), .B(n915), .C(n925), .Y(n952));
  AOI22X1 g0375(.A0(n917), .A1(REG0_REG_1__SCAN_IN), .B0(REG2_REG_1__SCAN_IN), .B1(n952), .Y(n953));
  NOR2X1  g0376(.A(n919), .B(n913), .Y(n954));
  NOR2X1  g0377(.A(n919), .B(n925), .Y(n955));
  AOI22X1 g0378(.A0(n954), .A1(REG1_REG_1__SCAN_IN), .B0(REG3_REG_1__SCAN_IN), .B1(n955), .Y(n956));
  NAND2X1 g0379(.A(n956), .B(n953), .Y(n957));
  NOR2X1  g0380(.A(n902), .B(n897), .Y(n958));
  AOI21X1 g0381(.A0(n907), .A1(n902), .B0(n958), .Y(n959));
  NOR3X1  g0382(.A(n889), .B(n876), .C(n884), .Y(n960));
  INVX1   g0383(.A(n960), .Y(n961));
  NOR3X1  g0384(.A(n878), .B(n876), .C(n884), .Y(n962));
  INVX1   g0385(.A(n962), .Y(n963));
  AOI21X1 g0386(.A0(n963), .A1(n961), .B0(n959), .Y(n964));
  AOI21X1 g0387(.A0(n957), .A1(n951), .B0(n964), .Y(n965));
  OAI21X1 g0388(.A0(n950), .A1(n930), .B0(n965), .Y(n966));
  NOR2X1  g0389(.A(n966), .B(n948), .Y(n967));
  NAND2X1 g0390(.A(n896), .B(REG0_REG_0__SCAN_IN), .Y(n968));
  OAI21X1 g0391(.A0(n967), .A1(n896), .B0(n968), .Y(U3467));
  INVX1   g0392(.A(DATAI_1_), .Y(n970));
  NAND2X1 g0393(.A(n759), .B(IR_REG_1__SCAN_IN), .Y(n971));
  OAI21X1 g0394(.A0(n582), .A1(n759), .B0(n971), .Y(n972));
  NAND2X1 g0395(.A(n972), .B(n902), .Y(n973));
  OAI21X1 g0396(.A0(n902), .A1(n970), .B0(n973), .Y(n974));
  XOR2X1  g0397(.A(n974), .B(n957), .Y(n975));
  NOR2X1  g0398(.A(n929), .B(n959), .Y(n976));
  INVX1   g0399(.A(n976), .Y(n977));
  XOR2X1  g0400(.A(n977), .B(n975), .Y(n978));
  INVX1   g0401(.A(n978), .Y(n979));
  OAI21X1 g0402(.A0(n946), .A1(n939), .B0(n979), .Y(n980));
  AOI22X1 g0403(.A0(n917), .A1(REG0_REG_0__SCAN_IN), .B0(REG2_REG_0__SCAN_IN), .B1(n952), .Y(n981));
  INVX1   g0404(.A(n916), .Y(n982));
  OAI21X1 g0405(.A0(n745), .A1(n759), .B0(n982), .Y(n983));
  NAND3X1 g0406(.A(n983), .B(n925), .C(REG1_REG_0__SCAN_IN), .Y(n984));
  NAND3X1 g0407(.A(n983), .B(n913), .C(REG3_REG_0__SCAN_IN), .Y(n985));
  NAND3X1 g0408(.A(n985), .B(n984), .C(n981), .Y(n986));
  NOR2X1  g0409(.A(n986), .B(n959), .Y(n987));
  XOR2X1  g0410(.A(n975), .B(n987), .Y(n989));
  AOI22X1 g0411(.A0(n979), .A1(n945), .B0(n936), .B1(n989), .Y(n990));
  NOR2X1  g0412(.A(n901), .B(n900), .Y(n991));
  NOR3X1  g0413(.A(n991), .B(n886), .C(n873), .Y(n992));
  AOI22X1 g0414(.A0(n989), .A1(n943), .B0(n986), .B1(n992), .Y(n993));
  OAI21X1 g0415(.A0(n941), .A1(n931), .B0(n989), .Y(n994));
  NAND4X1 g0416(.A(n993), .B(n990), .C(n980), .D(n994), .Y(n995));
  NOR2X1  g0417(.A(n978), .B(n950), .Y(n996));
  NOR2X1  g0418(.A(n902), .B(n970), .Y(n997));
  AOI21X1 g0419(.A0(n972), .A1(n902), .B0(n997), .Y(n998));
  XOR2X1  g0420(.A(n998), .B(n909), .Y(n999));
  AOI22X1 g0421(.A0(n917), .A1(REG0_REG_2__SCAN_IN), .B0(REG2_REG_2__SCAN_IN), .B1(n952), .Y(n1000));
  AOI22X1 g0422(.A0(n954), .A1(REG1_REG_2__SCAN_IN), .B0(REG3_REG_2__SCAN_IN), .B1(n955), .Y(n1001));
  NAND2X1 g0423(.A(n1001), .B(n1000), .Y(n1002));
  AOI22X1 g0424(.A0(n974), .A1(n962), .B0(n951), .B1(n1002), .Y(n1003));
  OAI21X1 g0425(.A0(n999), .A1(n961), .B0(n1003), .Y(n1004));
  NOR3X1  g0426(.A(n1004), .B(n996), .C(n995), .Y(n1005));
  NAND2X1 g0427(.A(n896), .B(REG0_REG_1__SCAN_IN), .Y(n1006));
  OAI21X1 g0428(.A0(n1005), .A1(n896), .B0(n1006), .Y(U3469));
  INVX1   g0429(.A(DATAI_2_), .Y(n1008));
  NAND2X1 g0430(.A(n759), .B(IR_REG_2__SCAN_IN), .Y(n1009));
  OAI21X1 g0431(.A0(n586), .A1(n759), .B0(n1009), .Y(n1010));
  NAND2X1 g0432(.A(n1010), .B(n902), .Y(n1011));
  OAI21X1 g0433(.A0(n902), .A1(n1008), .B0(n1011), .Y(n1012));
  XOR2X1  g0434(.A(n1012), .B(n1002), .Y(n1013));
  INVX1   g0435(.A(REG2_REG_1__SCAN_IN), .Y(n1014));
  NAND2X1 g0436(.A(n917), .B(REG0_REG_1__SCAN_IN), .Y(n1015));
  OAI21X1 g0437(.A0(n920), .A1(n1014), .B0(n1015), .Y(n1016));
  INVX1   g0438(.A(REG3_REG_1__SCAN_IN), .Y(n1017));
  INVX1   g0439(.A(REG1_REG_1__SCAN_IN), .Y(n1018));
  OAI22X1 g0440(.A0(n926), .A1(n1018), .B0(n1017), .B1(n927), .Y(n1019));
  NOR2X1  g0441(.A(n1019), .B(n1016), .Y(n1020));
  AOI21X1 g0442(.A0(n998), .A1(n1020), .B0(n977), .Y(n1021));
  INVX1   g0443(.A(n1021), .Y(n1022));
  OAI21X1 g0444(.A0(n998), .A1(n1020), .B0(n1022), .Y(n1023));
  NOR2X1  g0445(.A(n998), .B(n1020), .Y(n1024));
  NOR2X1  g0446(.A(n902), .B(n1008), .Y(n1025));
  AOI21X1 g0447(.A0(n1010), .A1(n902), .B0(n1025), .Y(n1026));
  NOR2X1  g0448(.A(n1026), .B(n1002), .Y(n1027));
  INVX1   g0449(.A(REG2_REG_2__SCAN_IN), .Y(n1028));
  NAND2X1 g0450(.A(n917), .B(REG0_REG_2__SCAN_IN), .Y(n1029));
  OAI21X1 g0451(.A0(n920), .A1(n1028), .B0(n1029), .Y(n1030));
  INVX1   g0452(.A(REG1_REG_2__SCAN_IN), .Y(n1031));
  INVX1   g0453(.A(REG3_REG_2__SCAN_IN), .Y(n1032));
  OAI22X1 g0454(.A0(n926), .A1(n1031), .B0(n1032), .B1(n927), .Y(n1033));
  NOR2X1  g0455(.A(n1033), .B(n1030), .Y(n1034));
  NOR2X1  g0456(.A(n1012), .B(n1034), .Y(n1035));
  NOR4X1  g0457(.A(n1027), .B(n1021), .C(n1024), .D(n1035), .Y(n1036));
  AOI21X1 g0458(.A0(n1023), .A1(n1013), .B0(n1036), .Y(n1037));
  AOI22X1 g0459(.A0(n992), .A1(n957), .B0(n945), .B1(n1037), .Y(n1038));
  OAI21X1 g0460(.A0(n946), .A1(n939), .B0(n1037), .Y(n1039));
  XOR2X1  g0461(.A(n1026), .B(n1002), .Y(n1040));
  INVX1   g0462(.A(n987), .Y(n1041));
  OAI21X1 g0463(.A0(n957), .A1(n1041), .B0(n998), .Y(n1042));
  OAI21X1 g0464(.A0(n1020), .A1(n987), .B0(n1042), .Y(n1043));
  XOR2X1  g0465(.A(n1043), .B(n1040), .Y(n1044));
  OAI21X1 g0466(.A0(n943), .A1(n941), .B0(n1044), .Y(n1045));
  OAI21X1 g0467(.A0(n936), .A1(n931), .B0(n1044), .Y(n1046));
  NAND4X1 g0468(.A(n1045), .B(n1039), .C(n1038), .D(n1046), .Y(n1047));
  NAND2X1 g0469(.A(n1037), .B(n949), .Y(n1048));
  NAND2X1 g0470(.A(n998), .B(n959), .Y(n1049));
  XOR2X1  g0471(.A(n1049), .B(n1012), .Y(n1050));
  INVX1   g0472(.A(n951), .Y(n1051));
  INVX1   g0473(.A(REG2_REG_3__SCAN_IN), .Y(n1052));
  NAND2X1 g0474(.A(n917), .B(REG0_REG_3__SCAN_IN), .Y(n1053));
  OAI21X1 g0475(.A0(n920), .A1(n1052), .B0(n1053), .Y(n1054));
  INVX1   g0476(.A(REG1_REG_3__SCAN_IN), .Y(n1055));
  OAI22X1 g0477(.A0(n926), .A1(n1055), .B0(REG3_REG_3__SCAN_IN), .B1(n927), .Y(n1056));
  NOR2X1  g0478(.A(n1056), .B(n1054), .Y(n1057));
  OAI22X1 g0479(.A0(n1026), .A1(n963), .B0(n1051), .B1(n1057), .Y(n1058));
  AOI21X1 g0480(.A0(n1050), .A1(n960), .B0(n1058), .Y(n1059));
  NAND2X1 g0481(.A(n1059), .B(n1048), .Y(n1060));
  NOR2X1  g0482(.A(n1060), .B(n1047), .Y(n1061));
  NAND2X1 g0483(.A(n896), .B(REG0_REG_2__SCAN_IN), .Y(n1062));
  OAI21X1 g0484(.A0(n1061), .A1(n896), .B0(n1062), .Y(U3471));
  NOR2X1  g0485(.A(n1012), .B(n1002), .Y(n1064));
  NOR2X1  g0486(.A(n1026), .B(n1034), .Y(n1065));
  INVX1   g0487(.A(n1064), .Y(n1066));
  AOI21X1 g0488(.A0(n1066), .A1(n1024), .B0(n1065), .Y(n1067));
  OAI21X1 g0489(.A0(n1022), .A1(n1064), .B0(n1067), .Y(n1068));
  INVX1   g0490(.A(DATAI_3_), .Y(n1069));
  NAND2X1 g0491(.A(n759), .B(IR_REG_3__SCAN_IN), .Y(n1070));
  OAI21X1 g0492(.A0(n590), .A1(n759), .B0(n1070), .Y(n1071));
  NAND2X1 g0493(.A(n1071), .B(n902), .Y(n1072));
  OAI21X1 g0494(.A0(n902), .A1(n1069), .B0(n1072), .Y(n1073));
  XOR2X1  g0495(.A(n1073), .B(n1057), .Y(n1074));
  NOR2X1  g0496(.A(n1074), .B(n1068), .Y(n1075));
  AOI22X1 g0497(.A0(n917), .A1(REG0_REG_3__SCAN_IN), .B0(REG2_REG_3__SCAN_IN), .B1(n952), .Y(n1076));
  INVX1   g0498(.A(REG3_REG_3__SCAN_IN), .Y(n1077));
  AOI22X1 g0499(.A0(n954), .A1(REG1_REG_3__SCAN_IN), .B0(n1077), .B1(n955), .Y(n1078));
  NAND2X1 g0500(.A(n1078), .B(n1076), .Y(n1079));
  XOR2X1  g0501(.A(n1073), .B(n1079), .Y(n1080));
  AOI21X1 g0502(.A0(n1074), .A1(n1068), .B0(n1075), .Y(n1082));
  INVX1   g0503(.A(n1082), .Y(n1083));
  AOI22X1 g0504(.A0(n1002), .A1(n992), .B0(n945), .B1(n1083), .Y(n1084));
  OAI21X1 g0505(.A0(n946), .A1(n939), .B0(n1083), .Y(n1085));
  INVX1   g0506(.A(n941), .Y(n1086));
  NOR2X1  g0507(.A(n1074), .B(n1027), .Y(n1087));
  OAI21X1 g0508(.A0(n1043), .A1(n1035), .B0(n1087), .Y(n1088));
  INVX1   g0509(.A(n1043), .Y(n1089));
  NOR2X1  g0510(.A(n902), .B(n1069), .Y(n1090));
  AOI21X1 g0511(.A0(n1071), .A1(n902), .B0(n1090), .Y(n1091));
  NOR2X1  g0512(.A(n1091), .B(n1079), .Y(n1092));
  NOR2X1  g0513(.A(n1073), .B(n1057), .Y(n1093));
  NOR3X1  g0514(.A(n1093), .B(n1092), .C(n1035), .Y(n1094));
  OAI21X1 g0515(.A0(n1089), .A1(n1027), .B0(n1094), .Y(n1095));
  AOI22X1 g0516(.A0(n1088), .A1(n1095), .B0(n942), .B1(n1086), .Y(n1096));
  NAND3X1 g0517(.A(n938), .B(n889), .C(n884), .Y(n1097));
  AOI22X1 g0518(.A0(n1088), .A1(n1095), .B0(n1097), .B1(n932), .Y(n1098));
  NOR2X1  g0519(.A(n1098), .B(n1096), .Y(n1099));
  NAND3X1 g0520(.A(n1099), .B(n1085), .C(n1084), .Y(n1100));
  NOR3X1  g0521(.A(n1012), .B(n974), .C(n909), .Y(n1101));
  XOR2X1  g0522(.A(n1091), .B(n1101), .Y(n1102));
  INVX1   g0523(.A(REG2_REG_4__SCAN_IN), .Y(n1103));
  NAND2X1 g0524(.A(n917), .B(REG0_REG_4__SCAN_IN), .Y(n1104));
  OAI21X1 g0525(.A0(n920), .A1(n1103), .B0(n1104), .Y(n1105));
  INVX1   g0526(.A(REG1_REG_4__SCAN_IN), .Y(n1106));
  XOR2X1  g0527(.A(REG3_REG_4__SCAN_IN), .B(n1077), .Y(n1107));
  OAI22X1 g0528(.A0(n927), .A1(n1107), .B0(n926), .B1(n1106), .Y(n1108));
  NOR2X1  g0529(.A(n1108), .B(n1105), .Y(n1109));
  OAI22X1 g0530(.A0(n1091), .A1(n963), .B0(n1051), .B1(n1109), .Y(n1110));
  AOI21X1 g0531(.A0(n1102), .A1(n960), .B0(n1110), .Y(n1111));
  OAI21X1 g0532(.A0(n1082), .A1(n950), .B0(n1111), .Y(n1112));
  NOR2X1  g0533(.A(n1112), .B(n1100), .Y(n1113));
  NAND2X1 g0534(.A(n896), .B(REG0_REG_3__SCAN_IN), .Y(n1114));
  OAI21X1 g0535(.A0(n1113), .A1(n896), .B0(n1114), .Y(U3473));
  INVX1   g0536(.A(n945), .Y(n1116));
  INVX1   g0537(.A(n992), .Y(n1117));
  NOR2X1  g0538(.A(n1091), .B(n1057), .Y(n1118));
  AOI22X1 g0539(.A0(n917), .A1(REG0_REG_4__SCAN_IN), .B0(REG2_REG_4__SCAN_IN), .B1(n952), .Y(n1119));
  INVX1   g0540(.A(n1107), .Y(n1120));
  AOI22X1 g0541(.A0(n955), .A1(n1120), .B0(n954), .B1(REG1_REG_4__SCAN_IN), .Y(n1121));
  NAND2X1 g0542(.A(n1121), .B(n1119), .Y(n1122));
  NAND2X1 g0543(.A(n759), .B(IR_REG_4__SCAN_IN), .Y(n1123));
  OAI21X1 g0544(.A0(n594), .A1(n759), .B0(n1123), .Y(n1124));
  INVX1   g0545(.A(DATAI_4_), .Y(n1125));
  NOR2X1  g0546(.A(n902), .B(n1125), .Y(n1126));
  AOI21X1 g0547(.A0(n1124), .A1(n902), .B0(n1126), .Y(n1127));
  XOR2X1  g0548(.A(n1127), .B(n1122), .Y(n1128));
  NOR2X1  g0549(.A(n1073), .B(n1079), .Y(n1129));
  NOR2X1  g0550(.A(n1129), .B(n1067), .Y(n1130));
  NOR3X1  g0551(.A(n1129), .B(n1022), .C(n1064), .Y(n1131));
  NOR4X1  g0552(.A(n1130), .B(n1128), .C(n1118), .D(n1131), .Y(n1132));
  NOR3X1  g0553(.A(n1131), .B(n1130), .C(n1118), .Y(n1133));
  NAND2X1 g0554(.A(n1124), .B(n902), .Y(n1134));
  OAI21X1 g0555(.A0(n902), .A1(n1125), .B0(n1134), .Y(n1135));
  XOR2X1  g0556(.A(n1135), .B(n1122), .Y(n1136));
  NOR2X1  g0557(.A(n1136), .B(n1133), .Y(n1137));
  NOR2X1  g0558(.A(n1137), .B(n1132), .Y(n1138));
  OAI22X1 g0559(.A0(n1057), .A1(n1117), .B0(n1116), .B1(n1138), .Y(n1139));
  INVX1   g0560(.A(n939), .Y(n1140));
  INVX1   g0561(.A(n946), .Y(n1141));
  AOI21X1 g0562(.A0(n1141), .A1(n1140), .B0(n1138), .Y(n1142));
  AOI22X1 g0563(.A0(n1057), .A1(n1073), .B0(n1012), .B1(n1034), .Y(n1144));
  NAND2X1 g0564(.A(n1144), .B(n1043), .Y(n1145));
  INVX1   g0565(.A(n1035), .Y(n1146));
  AOI21X1 g0566(.A0(n1057), .A1(n1146), .B0(n1073), .Y(n1147));
  AOI21X1 g0567(.A0(n1079), .A1(n1035), .B0(n1147), .Y(n1148));
  NAND2X1 g0568(.A(n1148), .B(n1145), .Y(n1149));
  XOR2X1  g0569(.A(n1149), .B(n1136), .Y(n1150));
  INVX1   g0570(.A(n1150), .Y(n1151));
  OAI21X1 g0571(.A0(n943), .A1(n941), .B0(n1151), .Y(n1152));
  OAI21X1 g0572(.A0(n936), .A1(n931), .B0(n1151), .Y(n1153));
  NAND2X1 g0573(.A(n1153), .B(n1152), .Y(n1154));
  NOR4X1  g0574(.A(n1012), .B(n974), .C(n909), .D(n1073), .Y(n1155));
  NOR4X1  g0575(.A(n1073), .B(n1049), .C(n1012), .D(n1135), .Y(n1156));
  INVX1   g0576(.A(n1156), .Y(n1157));
  OAI21X1 g0577(.A0(n1127), .A1(n1155), .B0(n1157), .Y(n1158));
  NOR2X1  g0578(.A(n1158), .B(n961), .Y(n1159));
  INVX1   g0579(.A(REG2_REG_5__SCAN_IN), .Y(n1160));
  NAND2X1 g0580(.A(n917), .B(REG0_REG_5__SCAN_IN), .Y(n1161));
  OAI21X1 g0581(.A0(n920), .A1(n1160), .B0(n1161), .Y(n1162));
  INVX1   g0582(.A(REG1_REG_5__SCAN_IN), .Y(n1163));
  NAND2X1 g0583(.A(REG3_REG_4__SCAN_IN), .B(REG3_REG_3__SCAN_IN), .Y(n1164));
  XOR2X1  g0584(.A(n1164), .B(REG3_REG_5__SCAN_IN), .Y(n1165));
  OAI22X1 g0585(.A0(n927), .A1(n1165), .B0(n926), .B1(n1163), .Y(n1166));
  NOR2X1  g0586(.A(n1166), .B(n1162), .Y(n1167));
  OAI22X1 g0587(.A0(n1127), .A1(n963), .B0(n1051), .B1(n1167), .Y(n1168));
  NOR2X1  g0588(.A(n1168), .B(n1159), .Y(n1169));
  OAI21X1 g0589(.A0(n1138), .A1(n950), .B0(n1169), .Y(n1170));
  NOR4X1  g0590(.A(n1154), .B(n1142), .C(n1139), .D(n1170), .Y(n1171));
  NAND2X1 g0591(.A(n896), .B(REG0_REG_4__SCAN_IN), .Y(n1172));
  OAI21X1 g0592(.A0(n1171), .A1(n896), .B0(n1172), .Y(U3475));
  INVX1   g0593(.A(DATAI_5_), .Y(n1174));
  NAND2X1 g0594(.A(n759), .B(IR_REG_5__SCAN_IN), .Y(n1175));
  OAI21X1 g0595(.A0(n602), .A1(n759), .B0(n1175), .Y(n1176));
  NAND2X1 g0596(.A(n1176), .B(n902), .Y(n1177));
  OAI21X1 g0597(.A0(n902), .A1(n1174), .B0(n1177), .Y(n1178));
  XOR2X1  g0598(.A(n1178), .B(n1167), .Y(n1179));
  NAND2X1 g0599(.A(n1135), .B(n1109), .Y(n1180));
  NOR2X1  g0600(.A(n1135), .B(n1109), .Y(n1181));
  AOI21X1 g0601(.A0(n1149), .A1(n1180), .B0(n1181), .Y(n1182));
  XOR2X1  g0602(.A(n1182), .B(n1179), .Y(n1183));
  NOR2X1  g0603(.A(n1183), .B(n942), .Y(n1184));
  NOR2X1  g0604(.A(n1127), .B(n1109), .Y(n1185));
  NOR4X1  g0605(.A(n1131), .B(n1130), .C(n1118), .D(n1185), .Y(n1186));
  NOR2X1  g0606(.A(n902), .B(n1174), .Y(n1187));
  AOI21X1 g0607(.A0(n1176), .A1(n902), .B0(n1187), .Y(n1188));
  NOR2X1  g0608(.A(n1188), .B(n1167), .Y(n1189));
  AOI22X1 g0609(.A0(n1167), .A1(n1188), .B0(n1127), .B1(n1109), .Y(n1190));
  INVX1   g0610(.A(n1190), .Y(n1191));
  NOR3X1  g0611(.A(n1191), .B(n1189), .C(n1186), .Y(n1192));
  AOI22X1 g0612(.A0(n917), .A1(REG0_REG_5__SCAN_IN), .B0(REG2_REG_5__SCAN_IN), .B1(n952), .Y(n1193));
  INVX1   g0613(.A(n1165), .Y(n1194));
  AOI22X1 g0614(.A0(n955), .A1(n1194), .B0(n954), .B1(REG1_REG_5__SCAN_IN), .Y(n1195));
  NAND2X1 g0615(.A(n1195), .B(n1193), .Y(n1196));
  NOR2X1  g0616(.A(n1188), .B(n1196), .Y(n1197));
  NOR2X1  g0617(.A(n1178), .B(n1167), .Y(n1198));
  AOI21X1 g0618(.A0(n1127), .A1(n1109), .B0(n1133), .Y(n1199));
  NOR4X1  g0619(.A(n1198), .B(n1197), .C(n1185), .D(n1199), .Y(n1200));
  NOR2X1  g0620(.A(n1200), .B(n1192), .Y(n1201));
  AOI22X1 g0621(.A0(n1122), .A1(n992), .B0(n945), .B1(n1201), .Y(n1202));
  INVX1   g0622(.A(n1202), .Y(n1203));
  OAI21X1 g0623(.A0(n946), .A1(n939), .B0(n1201), .Y(n1204));
  INVX1   g0624(.A(n1204), .Y(n1205));
  INVX1   g0625(.A(n1183), .Y(n1206));
  OAI21X1 g0626(.A0(n941), .A1(n931), .B0(n1206), .Y(n1207));
  OAI21X1 g0627(.A0(n1183), .A1(n1097), .B0(n1207), .Y(n1208));
  NOR4X1  g0628(.A(n1205), .B(n1203), .C(n1184), .D(n1208), .Y(n1209));
  INVX1   g0629(.A(n1209), .Y(n1210));
  NOR3X1  g0630(.A(n1200), .B(n1192), .C(n950), .Y(n1211));
  XOR2X1  g0631(.A(n1178), .B(n1156), .Y(n1212));
  AOI22X1 g0632(.A0(n917), .A1(REG0_REG_6__SCAN_IN), .B0(REG2_REG_6__SCAN_IN), .B1(n952), .Y(n1213));
  NAND3X1 g0633(.A(REG3_REG_4__SCAN_IN), .B(REG3_REG_5__SCAN_IN), .C(REG3_REG_3__SCAN_IN), .Y(n1214));
  XOR2X1  g0634(.A(n1214), .B(REG3_REG_6__SCAN_IN), .Y(n1215));
  INVX1   g0635(.A(n1215), .Y(n1216));
  AOI22X1 g0636(.A0(n955), .A1(n1216), .B0(n954), .B1(REG1_REG_6__SCAN_IN), .Y(n1217));
  NAND2X1 g0637(.A(n1217), .B(n1213), .Y(n1218));
  AOI22X1 g0638(.A0(n1178), .A1(n962), .B0(n951), .B1(n1218), .Y(n1219));
  OAI21X1 g0639(.A0(n1212), .A1(n961), .B0(n1219), .Y(n1220));
  NOR3X1  g0640(.A(n1220), .B(n1211), .C(n1210), .Y(n1221));
  NAND2X1 g0641(.A(n896), .B(REG0_REG_5__SCAN_IN), .Y(n1222));
  OAI21X1 g0642(.A0(n1221), .A1(n896), .B0(n1222), .Y(U3477));
  OAI21X1 g0643(.A0(n1178), .A1(n1167), .B0(n1182), .Y(n1224));
  NAND2X1 g0644(.A(n759), .B(IR_REG_6__SCAN_IN), .Y(n1225));
  OAI21X1 g0645(.A0(n606), .A1(n759), .B0(n1225), .Y(n1226));
  INVX1   g0646(.A(DATAI_6_), .Y(n1227));
  NOR2X1  g0647(.A(n902), .B(n1227), .Y(n1228));
  AOI21X1 g0648(.A0(n1226), .A1(n902), .B0(n1228), .Y(n1229));
  XOR2X1  g0649(.A(n1229), .B(n1218), .Y(n1230));
  NOR2X1  g0650(.A(n1230), .B(n1197), .Y(n1231));
  NAND2X1 g0651(.A(n1231), .B(n1224), .Y(n1232));
  NOR2X1  g0652(.A(n1182), .B(n1197), .Y(n1233));
  AOI22X1 g0653(.A0(n1218), .A1(n1229), .B0(n1188), .B1(n1196), .Y(n1234));
  OAI21X1 g0654(.A0(n1229), .A1(n1218), .B0(n1234), .Y(n1235));
  OAI21X1 g0655(.A0(n1235), .A1(n1233), .B0(n1232), .Y(n1236));
  INVX1   g0656(.A(n1236), .Y(n1237));
  NOR2X1  g0657(.A(n1237), .B(n942), .Y(n1238));
  NAND3X1 g0658(.A(n1178), .B(n1135), .C(n1122), .Y(n1239));
  AOI21X1 g0659(.A0(n1135), .A1(n1122), .B0(n1178), .Y(n1240));
  OAI21X1 g0660(.A0(n1240), .A1(n1167), .B0(n1239), .Y(n1241));
  NAND2X1 g0661(.A(n1073), .B(n1079), .Y(n1242));
  OAI21X1 g0662(.A0(n1073), .A1(n1079), .B0(n1065), .Y(n1243));
  AOI21X1 g0663(.A0(n1243), .A1(n1242), .B0(n1191), .Y(n1244));
  NOR2X1  g0664(.A(n1244), .B(n1241), .Y(n1245));
  INVX1   g0665(.A(n1129), .Y(n1246));
  NAND4X1 g0666(.A(n1246), .B(n1021), .C(n1066), .D(n1190), .Y(n1247));
  NAND4X1 g0667(.A(n1246), .B(n1066), .C(n1024), .D(n1190), .Y(n1248));
  NAND3X1 g0668(.A(n1248), .B(n1247), .C(n1245), .Y(n1249));
  NOR2X1  g0669(.A(n1249), .B(n1230), .Y(n1250));
  NAND2X1 g0670(.A(n1226), .B(n902), .Y(n1251));
  OAI21X1 g0671(.A0(n902), .A1(n1227), .B0(n1251), .Y(n1252));
  XOR2X1  g0672(.A(n1252), .B(n1218), .Y(n1253));
  AOI21X1 g0673(.A0(n1230), .A1(n1249), .B0(n1250), .Y(n1255));
  INVX1   g0674(.A(n1255), .Y(n1256));
  AOI22X1 g0675(.A0(n1196), .A1(n992), .B0(n945), .B1(n1256), .Y(n1257));
  OAI21X1 g0676(.A0(n946), .A1(n939), .B0(n1256), .Y(n1258));
  NAND2X1 g0677(.A(n1258), .B(n1257), .Y(n1259));
  NOR2X1  g0678(.A(n1237), .B(n1097), .Y(n1260));
  OAI21X1 g0679(.A0(n941), .A1(n931), .B0(n1236), .Y(n1261));
  INVX1   g0680(.A(n1261), .Y(n1262));
  NOR4X1  g0681(.A(n1260), .B(n1259), .C(n1238), .D(n1262), .Y(n1263));
  INVX1   g0682(.A(n1263), .Y(n1264));
  NOR2X1  g0683(.A(n1255), .B(n950), .Y(n1265));
  OAI21X1 g0684(.A0(n1178), .A1(n1157), .B0(n1252), .Y(n1266));
  NAND2X1 g0685(.A(n1229), .B(n1188), .Y(n1267));
  OAI21X1 g0686(.A0(n1267), .A1(n1157), .B0(n1266), .Y(n1268));
  AOI22X1 g0687(.A0(n917), .A1(REG0_REG_7__SCAN_IN), .B0(REG2_REG_7__SCAN_IN), .B1(n952), .Y(n1269));
  NAND4X1 g0688(.A(REG3_REG_4__SCAN_IN), .B(REG3_REG_5__SCAN_IN), .C(REG3_REG_3__SCAN_IN), .D(REG3_REG_6__SCAN_IN), .Y(n1270));
  XOR2X1  g0689(.A(n1270), .B(REG3_REG_7__SCAN_IN), .Y(n1271));
  INVX1   g0690(.A(n1271), .Y(n1272));
  AOI22X1 g0691(.A0(n955), .A1(n1272), .B0(n954), .B1(REG1_REG_7__SCAN_IN), .Y(n1273));
  NAND2X1 g0692(.A(n1273), .B(n1269), .Y(n1274));
  AOI22X1 g0693(.A0(n1252), .A1(n962), .B0(n951), .B1(n1274), .Y(n1275));
  OAI21X1 g0694(.A0(n1268), .A1(n961), .B0(n1275), .Y(n1276));
  NOR3X1  g0695(.A(n1276), .B(n1265), .C(n1264), .Y(n1277));
  NAND2X1 g0696(.A(n896), .B(REG0_REG_6__SCAN_IN), .Y(n1278));
  OAI21X1 g0697(.A0(n1277), .A1(n896), .B0(n1278), .Y(U3479));
  INVX1   g0698(.A(REG2_REG_6__SCAN_IN), .Y(n1280));
  NAND2X1 g0699(.A(n917), .B(REG0_REG_6__SCAN_IN), .Y(n1281));
  OAI21X1 g0700(.A0(n920), .A1(n1280), .B0(n1281), .Y(n1282));
  INVX1   g0701(.A(REG1_REG_6__SCAN_IN), .Y(n1283));
  OAI22X1 g0702(.A0(n927), .A1(n1215), .B0(n926), .B1(n1283), .Y(n1284));
  NOR2X1  g0703(.A(n1284), .B(n1282), .Y(n1285));
  NOR2X1  g0704(.A(n1229), .B(n1285), .Y(n1286));
  INVX1   g0705(.A(DATAI_7_), .Y(n1287));
  INVX1   g0706(.A(IR_REG_7__SCAN_IN), .Y(n1288));
  NAND2X1 g0707(.A(n611), .B(IR_REG_31__SCAN_IN), .Y(n1289));
  OAI21X1 g0708(.A0(IR_REG_31__SCAN_IN), .A1(n1288), .B0(n1289), .Y(n1290));
  NAND2X1 g0709(.A(n1290), .B(n902), .Y(n1291));
  OAI21X1 g0710(.A0(n902), .A1(n1287), .B0(n1291), .Y(n1292));
  INVX1   g0711(.A(REG2_REG_7__SCAN_IN), .Y(n1293));
  NAND2X1 g0712(.A(n917), .B(REG0_REG_7__SCAN_IN), .Y(n1294));
  OAI21X1 g0713(.A0(n920), .A1(n1293), .B0(n1294), .Y(n1295));
  INVX1   g0714(.A(REG1_REG_7__SCAN_IN), .Y(n1296));
  OAI22X1 g0715(.A0(n927), .A1(n1271), .B0(n926), .B1(n1296), .Y(n1297));
  NOR2X1  g0716(.A(n1297), .B(n1295), .Y(n1298));
  NOR2X1  g0717(.A(n902), .B(n1287), .Y(n1299));
  AOI21X1 g0718(.A0(n1290), .A1(n902), .B0(n1299), .Y(n1300));
  AOI22X1 g0719(.A0(n1298), .A1(n1300), .B0(n1229), .B1(n1285), .Y(n1301));
  INVX1   g0720(.A(n1301), .Y(n1302));
  AOI21X1 g0721(.A0(n1292), .A1(n1274), .B0(n1302), .Y(n1303));
  OAI21X1 g0722(.A0(n1286), .A1(n1249), .B0(n1303), .Y(n1304));
  INVX1   g0723(.A(n1249), .Y(n1305));
  AOI21X1 g0724(.A0(n1229), .A1(n1285), .B0(n1305), .Y(n1306));
  NOR2X1  g0725(.A(n1300), .B(n1274), .Y(n1307));
  NOR2X1  g0726(.A(n1292), .B(n1298), .Y(n1308));
  NOR3X1  g0727(.A(n1308), .B(n1307), .C(n1286), .Y(n1309));
  INVX1   g0728(.A(n1309), .Y(n1310));
  OAI21X1 g0729(.A0(n1310), .A1(n1306), .B0(n1304), .Y(n1311));
  INVX1   g0730(.A(n1311), .Y(n1312));
  AOI22X1 g0731(.A0(n1218), .A1(n992), .B0(n945), .B1(n1312), .Y(n1313));
  OAI21X1 g0732(.A0(n946), .A1(n939), .B0(n1312), .Y(n1314));
  XOR2X1  g0733(.A(n1292), .B(n1298), .Y(n1315));
  NOR2X1  g0734(.A(n1229), .B(n1218), .Y(n1316));
  OAI21X1 g0735(.A0(n1188), .A1(n1196), .B0(n1181), .Y(n1317));
  AOI21X1 g0736(.A0(n1317), .A1(n1234), .B0(n1316), .Y(n1318));
  OAI22X1 g0737(.A0(n1218), .A1(n1229), .B0(n1127), .B1(n1122), .Y(n1319));
  NOR2X1  g0738(.A(n1319), .B(n1197), .Y(n1320));
  AOI21X1 g0739(.A0(n1320), .A1(n1149), .B0(n1318), .Y(n1321));
  XOR2X1  g0740(.A(n1321), .B(n1315), .Y(n1322));
  INVX1   g0741(.A(n1322), .Y(n1323));
  OAI21X1 g0742(.A0(n943), .A1(n941), .B0(n1323), .Y(n1324));
  OAI21X1 g0743(.A0(n936), .A1(n931), .B0(n1323), .Y(n1325));
  NAND4X1 g0744(.A(n1324), .B(n1314), .C(n1313), .D(n1325), .Y(n1326));
  NOR2X1  g0745(.A(n1311), .B(n950), .Y(n1327));
  NOR3X1  g0746(.A(n1252), .B(n1178), .C(n1157), .Y(n1328));
  XOR2X1  g0747(.A(n1292), .B(n1328), .Y(n1329));
  INVX1   g0748(.A(REG2_REG_8__SCAN_IN), .Y(n1330));
  NAND2X1 g0749(.A(n917), .B(REG0_REG_8__SCAN_IN), .Y(n1331));
  OAI21X1 g0750(.A0(n920), .A1(n1330), .B0(n1331), .Y(n1332));
  INVX1   g0751(.A(REG1_REG_8__SCAN_IN), .Y(n1333));
  INVX1   g0752(.A(REG3_REG_8__SCAN_IN), .Y(n1334));
  INVX1   g0753(.A(REG3_REG_7__SCAN_IN), .Y(n1335));
  NOR2X1  g0754(.A(n1270), .B(n1335), .Y(n1336));
  XOR2X1  g0755(.A(n1336), .B(n1334), .Y(n1337));
  OAI22X1 g0756(.A0(n927), .A1(n1337), .B0(n926), .B1(n1333), .Y(n1338));
  NOR2X1  g0757(.A(n1338), .B(n1332), .Y(n1339));
  INVX1   g0758(.A(n1339), .Y(n1340));
  AOI22X1 g0759(.A0(n1292), .A1(n962), .B0(n951), .B1(n1340), .Y(n1341));
  OAI21X1 g0760(.A0(n1329), .A1(n961), .B0(n1341), .Y(n1342));
  NOR3X1  g0761(.A(n1342), .B(n1327), .C(n1326), .Y(n1343));
  NAND2X1 g0762(.A(n896), .B(REG0_REG_7__SCAN_IN), .Y(n1344));
  OAI21X1 g0763(.A0(n1343), .A1(n896), .B0(n1344), .Y(U3481));
  NAND3X1 g0764(.A(n1292), .B(n1252), .C(n1218), .Y(n1346));
  AOI21X1 g0765(.A0(n1252), .A1(n1218), .B0(n1292), .Y(n1347));
  OAI21X1 g0766(.A0(n1347), .A1(n1298), .B0(n1346), .Y(n1348));
  AOI21X1 g0767(.A0(n1301), .A1(n1249), .B0(n1348), .Y(n1349));
  INVX1   g0768(.A(DATAI_8_), .Y(n1350));
  NAND2X1 g0769(.A(n759), .B(IR_REG_8__SCAN_IN), .Y(n1351));
  OAI21X1 g0770(.A0(n615), .A1(n759), .B0(n1351), .Y(n1352));
  NAND2X1 g0771(.A(n1352), .B(n902), .Y(n1353));
  OAI21X1 g0772(.A0(n902), .A1(n1350), .B0(n1353), .Y(n1354));
  XOR2X1  g0773(.A(n1354), .B(n1339), .Y(n1355));
  NOR2X1  g0774(.A(n902), .B(n1350), .Y(n1357));
  AOI21X1 g0775(.A0(n1352), .A1(n902), .B0(n1357), .Y(n1358));
  XOR2X1  g0776(.A(n1358), .B(n1339), .Y(n1359));
  NOR2X1  g0777(.A(n1359), .B(n1349), .Y(n1360));
  AOI21X1 g0778(.A0(n1359), .A1(n1349), .B0(n1360), .Y(n1361));
  OAI22X1 g0779(.A0(n1298), .A1(n1117), .B0(n1116), .B1(n1361), .Y(n1362));
  AOI21X1 g0780(.A0(n1141), .A1(n1140), .B0(n1361), .Y(n1363));
  OAI21X1 g0781(.A0(n1292), .A1(n1298), .B0(n1321), .Y(n1364));
  NOR2X1  g0782(.A(n1355), .B(n1307), .Y(n1365));
  NAND2X1 g0783(.A(n1365), .B(n1364), .Y(n1366));
  NOR2X1  g0784(.A(n1359), .B(n1308), .Y(n1367));
  OAI21X1 g0785(.A0(n1321), .A1(n1307), .B0(n1367), .Y(n1368));
  NAND2X1 g0786(.A(n1368), .B(n1366), .Y(n1369));
  OAI21X1 g0787(.A0(n943), .A1(n941), .B0(n1369), .Y(n1370));
  OAI21X1 g0788(.A0(n936), .A1(n931), .B0(n1369), .Y(n1371));
  NAND2X1 g0789(.A(n1371), .B(n1370), .Y(n1372));
  NAND4X1 g0790(.A(n1229), .B(n1188), .C(n1156), .D(n1300), .Y(n1373));
  XOR2X1  g0791(.A(n1354), .B(n1373), .Y(n1374));
  INVX1   g0792(.A(REG2_REG_9__SCAN_IN), .Y(n1375));
  NAND2X1 g0793(.A(n917), .B(REG0_REG_9__SCAN_IN), .Y(n1376));
  OAI21X1 g0794(.A0(n920), .A1(n1375), .B0(n1376), .Y(n1377));
  INVX1   g0795(.A(REG1_REG_9__SCAN_IN), .Y(n1378));
  INVX1   g0796(.A(REG3_REG_9__SCAN_IN), .Y(n1379));
  NOR3X1  g0797(.A(n1270), .B(n1334), .C(n1335), .Y(n1380));
  XOR2X1  g0798(.A(n1380), .B(n1379), .Y(n1381));
  OAI22X1 g0799(.A0(n927), .A1(n1381), .B0(n926), .B1(n1378), .Y(n1382));
  NOR2X1  g0800(.A(n1382), .B(n1377), .Y(n1383));
  OAI22X1 g0801(.A0(n1358), .A1(n963), .B0(n1051), .B1(n1383), .Y(n1384));
  AOI21X1 g0802(.A0(n1374), .A1(n960), .B0(n1384), .Y(n1385));
  OAI21X1 g0803(.A0(n1361), .A1(n950), .B0(n1385), .Y(n1386));
  NOR4X1  g0804(.A(n1372), .B(n1363), .C(n1362), .D(n1386), .Y(n1387));
  NAND2X1 g0805(.A(n896), .B(REG0_REG_8__SCAN_IN), .Y(n1388));
  OAI21X1 g0806(.A0(n1387), .A1(n896), .B0(n1388), .Y(U3483));
  AOI22X1 g0807(.A0(n917), .A1(REG0_REG_9__SCAN_IN), .B0(REG2_REG_9__SCAN_IN), .B1(n952), .Y(n1390));
  INVX1   g0808(.A(n1382), .Y(n1391));
  NAND2X1 g0809(.A(n1391), .B(n1390), .Y(n1392));
  NAND2X1 g0810(.A(n624), .B(IR_REG_31__SCAN_IN), .Y(n1393));
  OAI21X1 g0811(.A0(IR_REG_31__SCAN_IN), .A1(n621), .B0(n1393), .Y(n1394));
  INVX1   g0812(.A(DATAI_9_), .Y(n1395));
  NOR2X1  g0813(.A(n902), .B(n1395), .Y(n1396));
  AOI21X1 g0814(.A0(n1394), .A1(n902), .B0(n1396), .Y(n1397));
  XOR2X1  g0815(.A(n1397), .B(n1392), .Y(n1398));
  NOR3X1  g0816(.A(n1358), .B(n1338), .C(n1332), .Y(n1399));
  NOR4X1  g0817(.A(n1319), .B(n1307), .C(n1197), .D(n1399), .Y(n1400));
  AOI22X1 g0818(.A0(n1339), .A1(n1354), .B0(n1292), .B1(n1298), .Y(n1401));
  NAND2X1 g0819(.A(n1401), .B(n1318), .Y(n1402));
  NAND2X1 g0820(.A(n1340), .B(n1308), .Y(n1403));
  OAI21X1 g0821(.A0(n1340), .A1(n1308), .B0(n1358), .Y(n1404));
  NAND3X1 g0822(.A(n1404), .B(n1403), .C(n1402), .Y(n1405));
  AOI21X1 g0823(.A0(n1400), .A1(n1149), .B0(n1405), .Y(n1406));
  XOR2X1  g0824(.A(n1406), .B(n1398), .Y(n1407));
  INVX1   g0825(.A(n1407), .Y(n1408));
  AOI22X1 g0826(.A0(n1340), .A1(n992), .B0(n943), .B1(n1408), .Y(n1409));
  INVX1   g0827(.A(n1409), .Y(n1410));
  OAI21X1 g0828(.A0(n941), .A1(n931), .B0(n1408), .Y(n1411));
  OAI21X1 g0829(.A0(n1407), .A1(n1097), .B0(n1411), .Y(n1412));
  NOR3X1  g0830(.A(n1354), .B(n1338), .C(n1332), .Y(n1414));
  OAI21X1 g0831(.A0(n1338), .A1(n1332), .B0(n1354), .Y(n1415));
  OAI21X1 g0832(.A0(n1414), .A1(n1349), .B0(n1415), .Y(n1416));
  INVX1   g0833(.A(n1416), .Y(n1417));
  XOR2X1  g0834(.A(n1397), .B(n1383), .Y(n1418));
  NOR2X1  g0835(.A(n1418), .B(n1417), .Y(n1419));
  AOI21X1 g0836(.A0(n1417), .A1(n1418), .B0(n1419), .Y(n1420));
  INVX1   g0837(.A(n1420), .Y(n1421));
  OAI21X1 g0838(.A0(n945), .A1(n939), .B0(n1421), .Y(n1422));
  OAI21X1 g0839(.A0(n1420), .A1(n1141), .B0(n1422), .Y(n1423));
  NOR4X1  g0840(.A(n1292), .B(n1267), .C(n1157), .D(n1354), .Y(n1424));
  XOR2X1  g0841(.A(n1424), .B(n1397), .Y(n1425));
  INVX1   g0842(.A(REG2_REG_10__SCAN_IN), .Y(n1426));
  NAND2X1 g0843(.A(n917), .B(REG0_REG_10__SCAN_IN), .Y(n1427));
  OAI21X1 g0844(.A0(n920), .A1(n1426), .B0(n1427), .Y(n1428));
  INVX1   g0845(.A(REG1_REG_10__SCAN_IN), .Y(n1429));
  INVX1   g0846(.A(REG3_REG_10__SCAN_IN), .Y(n1430));
  NOR4X1  g0847(.A(n1379), .B(n1334), .C(n1335), .D(n1270), .Y(n1431));
  XOR2X1  g0848(.A(n1431), .B(n1430), .Y(n1432));
  OAI22X1 g0849(.A0(n927), .A1(n1432), .B0(n926), .B1(n1429), .Y(n1433));
  NOR2X1  g0850(.A(n1433), .B(n1428), .Y(n1434));
  OAI22X1 g0851(.A0(n1397), .A1(n963), .B0(n1051), .B1(n1434), .Y(n1435));
  AOI21X1 g0852(.A0(n1425), .A1(n960), .B0(n1435), .Y(n1436));
  OAI21X1 g0853(.A0(n1420), .A1(n950), .B0(n1436), .Y(n1437));
  NOR4X1  g0854(.A(n1423), .B(n1412), .C(n1410), .D(n1437), .Y(n1438));
  NAND2X1 g0855(.A(n896), .B(REG0_REG_9__SCAN_IN), .Y(n1439));
  OAI21X1 g0856(.A0(n1438), .A1(n896), .B0(n1439), .Y(U3485));
  AOI22X1 g0857(.A0(n917), .A1(REG0_REG_10__SCAN_IN), .B0(REG2_REG_10__SCAN_IN), .B1(n952), .Y(n1441));
  INVX1   g0858(.A(n1432), .Y(n1442));
  AOI22X1 g0859(.A0(n955), .A1(n1442), .B0(n954), .B1(REG1_REG_10__SCAN_IN), .Y(n1443));
  NAND2X1 g0860(.A(n1443), .B(n1441), .Y(n1444));
  NAND2X1 g0861(.A(n759), .B(IR_REG_10__SCAN_IN), .Y(n1445));
  OAI21X1 g0862(.A0(n628), .A1(n759), .B0(n1445), .Y(n1446));
  INVX1   g0863(.A(DATAI_10_), .Y(n1447));
  NOR2X1  g0864(.A(n902), .B(n1447), .Y(n1448));
  AOI21X1 g0865(.A0(n1446), .A1(n902), .B0(n1448), .Y(n1449));
  XOR2X1  g0866(.A(n1449), .B(n1444), .Y(n1450));
  INVX1   g0867(.A(n1397), .Y(n1451));
  NOR2X1  g0868(.A(n1451), .B(n1383), .Y(n1452));
  NOR2X1  g0869(.A(n1397), .B(n1392), .Y(n1453));
  NOR2X1  g0870(.A(n1406), .B(n1453), .Y(n1454));
  NOR2X1  g0871(.A(n1454), .B(n1452), .Y(n1455));
  XOR2X1  g0872(.A(n1455), .B(n1450), .Y(n1456));
  INVX1   g0873(.A(n1456), .Y(n1457));
  OAI21X1 g0874(.A0(n941), .A1(n931), .B0(n1457), .Y(n1458));
  OAI21X1 g0875(.A0(n1456), .A1(n1097), .B0(n1458), .Y(n1459));
  NAND2X1 g0876(.A(n1451), .B(n1392), .Y(n1460));
  INVX1   g0877(.A(n1449), .Y(n1461));
  NAND2X1 g0878(.A(n1449), .B(n1434), .Y(n1462));
  OAI21X1 g0879(.A0(n1451), .A1(n1392), .B0(n1462), .Y(n1463));
  AOI21X1 g0880(.A0(n1461), .A1(n1444), .B0(n1463), .Y(n1464));
  INVX1   g0881(.A(n1464), .Y(n1465));
  AOI21X1 g0882(.A0(n1460), .A1(n1417), .B0(n1465), .Y(n1466));
  NAND2X1 g0883(.A(n1397), .B(n1383), .Y(n1467));
  OAI21X1 g0884(.A0(n1397), .A1(n1383), .B0(n1450), .Y(n1468));
  AOI21X1 g0885(.A0(n1467), .A1(n1416), .B0(n1468), .Y(n1469));
  NOR3X1  g0886(.A(n1469), .B(n1466), .C(n1140), .Y(n1470));
  AOI22X1 g0887(.A0(n1392), .A1(n992), .B0(n943), .B1(n1457), .Y(n1471));
  INVX1   g0888(.A(n1471), .Y(n1472));
  NOR2X1  g0889(.A(n1469), .B(n1466), .Y(n1473));
  OAI21X1 g0890(.A0(n946), .A1(n945), .B0(n1473), .Y(n1474));
  INVX1   g0891(.A(n1474), .Y(n1475));
  NOR4X1  g0892(.A(n1472), .B(n1470), .C(n1459), .D(n1475), .Y(n1476));
  INVX1   g0893(.A(n1476), .Y(n1477));
  NAND2X1 g0894(.A(n1473), .B(n949), .Y(n1478));
  NAND4X1 g0895(.A(n1358), .B(n1300), .C(n1328), .D(n1397), .Y(n1479));
  XOR2X1  g0896(.A(n1461), .B(n1479), .Y(n1480));
  INVX1   g0897(.A(REG2_REG_11__SCAN_IN), .Y(n1481));
  NAND2X1 g0898(.A(n917), .B(REG0_REG_11__SCAN_IN), .Y(n1482));
  OAI21X1 g0899(.A0(n920), .A1(n1481), .B0(n1482), .Y(n1483));
  INVX1   g0900(.A(REG1_REG_11__SCAN_IN), .Y(n1484));
  INVX1   g0901(.A(REG3_REG_11__SCAN_IN), .Y(n1485));
  NAND2X1 g0902(.A(REG3_REG_9__SCAN_IN), .B(REG3_REG_8__SCAN_IN), .Y(n1486));
  NOR4X1  g0903(.A(n1270), .B(n1430), .C(n1335), .D(n1486), .Y(n1487));
  XOR2X1  g0904(.A(n1487), .B(n1485), .Y(n1488));
  OAI22X1 g0905(.A0(n927), .A1(n1488), .B0(n926), .B1(n1484), .Y(n1489));
  NOR2X1  g0906(.A(n1489), .B(n1483), .Y(n1490));
  OAI22X1 g0907(.A0(n1449), .A1(n963), .B0(n1051), .B1(n1490), .Y(n1491));
  AOI21X1 g0908(.A0(n1480), .A1(n960), .B0(n1491), .Y(n1492));
  NAND2X1 g0909(.A(n1492), .B(n1478), .Y(n1493));
  NOR2X1  g0910(.A(n1493), .B(n1477), .Y(n1494));
  NAND2X1 g0911(.A(n896), .B(REG0_REG_10__SCAN_IN), .Y(n1495));
  OAI21X1 g0912(.A0(n1494), .A1(n896), .B0(n1495), .Y(U3487));
  OAI21X1 g0913(.A0(n1461), .A1(n1434), .B0(n1455), .Y(n1497));
  NOR2X1  g0914(.A(n1449), .B(n1444), .Y(n1498));
  AOI22X1 g0915(.A0(n917), .A1(REG0_REG_11__SCAN_IN), .B0(REG2_REG_11__SCAN_IN), .B1(n952), .Y(n1499));
  INVX1   g0916(.A(n1488), .Y(n1500));
  AOI22X1 g0917(.A0(n955), .A1(n1500), .B0(n954), .B1(REG1_REG_11__SCAN_IN), .Y(n1501));
  NAND2X1 g0918(.A(n1501), .B(n1499), .Y(n1502));
  NAND2X1 g0919(.A(n635), .B(IR_REG_31__SCAN_IN), .Y(n1503));
  OAI21X1 g0920(.A0(IR_REG_31__SCAN_IN), .A1(n632), .B0(n1503), .Y(n1504));
  INVX1   g0921(.A(DATAI_11_), .Y(n1505));
  NOR2X1  g0922(.A(n902), .B(n1505), .Y(n1506));
  AOI21X1 g0923(.A0(n1504), .A1(n902), .B0(n1506), .Y(n1507));
  XOR2X1  g0924(.A(n1507), .B(n1502), .Y(n1508));
  NOR2X1  g0925(.A(n1508), .B(n1498), .Y(n1509));
  INVX1   g0926(.A(n1498), .Y(n1510));
  OAI21X1 g0927(.A0(n1454), .A1(n1452), .B0(n1510), .Y(n1511));
  NOR2X1  g0928(.A(n1461), .B(n1434), .Y(n1512));
  NOR2X1  g0929(.A(n1507), .B(n1502), .Y(n1513));
  INVX1   g0930(.A(n1507), .Y(n1514));
  NOR2X1  g0931(.A(n1514), .B(n1490), .Y(n1515));
  NOR3X1  g0932(.A(n1515), .B(n1513), .C(n1512), .Y(n1516));
  AOI22X1 g0933(.A0(n1511), .A1(n1516), .B0(n1509), .B1(n1497), .Y(n1517));
  INVX1   g0934(.A(n1517), .Y(n1518));
  NAND2X1 g0935(.A(n1518), .B(n943), .Y(n1519));
  NOR3X1  g0936(.A(n1463), .B(n1414), .C(n1302), .Y(n1521));
  NAND2X1 g0937(.A(n1358), .B(n1339), .Y(n1522));
  NAND4X1 g0938(.A(n1467), .B(n1522), .C(n1348), .D(n1462), .Y(n1523));
  AOI22X1 g0939(.A0(n1444), .A1(n1461), .B0(n1451), .B1(n1392), .Y(n1524));
  OAI21X1 g0940(.A0(n1463), .A1(n1415), .B0(n1524), .Y(n1525));
  NAND2X1 g0941(.A(n1525), .B(n1462), .Y(n1526));
  NAND2X1 g0942(.A(n1526), .B(n1523), .Y(n1527));
  AOI21X1 g0943(.A0(n1521), .A1(n1249), .B0(n1527), .Y(n1528));
  XOR2X1  g0944(.A(n1507), .B(n1490), .Y(n1529));
  NOR2X1  g0945(.A(n1529), .B(n1528), .Y(n1530));
  AOI21X1 g0946(.A0(n1528), .A1(n1529), .B0(n1530), .Y(n1531));
  INVX1   g0947(.A(n1531), .Y(n1532));
  AOI22X1 g0948(.A0(n1444), .A1(n992), .B0(n945), .B1(n1532), .Y(n1533));
  OAI21X1 g0949(.A0(n946), .A1(n939), .B0(n1532), .Y(n1534));
  NAND3X1 g0950(.A(n1534), .B(n1533), .C(n1519), .Y(n1535));
  NOR2X1  g0951(.A(n1517), .B(n1097), .Y(n1536));
  AOI21X1 g0952(.A0(n1086), .A1(n932), .B0(n1517), .Y(n1537));
  NAND3X1 g0953(.A(n1449), .B(n1424), .C(n1397), .Y(n1538));
  XOR2X1  g0954(.A(n1538), .B(n1514), .Y(n1539));
  INVX1   g0955(.A(REG2_REG_12__SCAN_IN), .Y(n1540));
  NAND2X1 g0956(.A(n917), .B(REG0_REG_12__SCAN_IN), .Y(n1541));
  OAI21X1 g0957(.A0(n920), .A1(n1540), .B0(n1541), .Y(n1542));
  INVX1   g0958(.A(REG1_REG_12__SCAN_IN), .Y(n1543));
  NAND3X1 g0959(.A(n1431), .B(REG3_REG_11__SCAN_IN), .C(REG3_REG_10__SCAN_IN), .Y(n1544));
  XOR2X1  g0960(.A(n1544), .B(REG3_REG_12__SCAN_IN), .Y(n1545));
  OAI22X1 g0961(.A0(n927), .A1(n1545), .B0(n926), .B1(n1543), .Y(n1546));
  NOR2X1  g0962(.A(n1546), .B(n1542), .Y(n1547));
  OAI22X1 g0963(.A0(n1507), .A1(n963), .B0(n1051), .B1(n1547), .Y(n1548));
  AOI21X1 g0964(.A0(n1539), .A1(n960), .B0(n1548), .Y(n1549));
  OAI21X1 g0965(.A0(n1531), .A1(n950), .B0(n1549), .Y(n1550));
  NOR4X1  g0966(.A(n1537), .B(n1536), .C(n1535), .D(n1550), .Y(n1551));
  NAND2X1 g0967(.A(n896), .B(REG0_REG_11__SCAN_IN), .Y(n1552));
  OAI21X1 g0968(.A0(n1551), .A1(n896), .B0(n1552), .Y(U3489));
  NOR2X1  g0969(.A(n1514), .B(n1502), .Y(n1554));
  NAND2X1 g0970(.A(n1514), .B(n1502), .Y(n1555));
  OAI21X1 g0971(.A0(n1554), .A1(n1528), .B0(n1555), .Y(n1556));
  INVX1   g0972(.A(DATAI_12_), .Y(n1557));
  NAND2X1 g0973(.A(n759), .B(IR_REG_12__SCAN_IN), .Y(n1558));
  OAI21X1 g0974(.A0(n639), .A1(n759), .B0(n1558), .Y(n1559));
  NAND2X1 g0975(.A(n1559), .B(n902), .Y(n1560));
  OAI21X1 g0976(.A0(n902), .A1(n1557), .B0(n1560), .Y(n1561));
  XOR2X1  g0977(.A(n1561), .B(n1547), .Y(n1562));
  NOR2X1  g0978(.A(n1556), .B(n1562), .Y(n1563));
  AOI22X1 g0979(.A0(n917), .A1(REG0_REG_12__SCAN_IN), .B0(REG2_REG_12__SCAN_IN), .B1(n952), .Y(n1564));
  INVX1   g0980(.A(n1545), .Y(n1565));
  AOI22X1 g0981(.A0(n955), .A1(n1565), .B0(n954), .B1(REG1_REG_12__SCAN_IN), .Y(n1566));
  NAND2X1 g0982(.A(n1566), .B(n1564), .Y(n1567));
  XOR2X1  g0983(.A(n1561), .B(n1567), .Y(n1568));
  AOI21X1 g0984(.A0(n1562), .A1(n1556), .B0(n1563), .Y(n1570));
  AOI21X1 g0985(.A0(n1141), .A1(n1140), .B0(n1570), .Y(n1571));
  INVX1   g0986(.A(n1513), .Y(n1572));
  OAI22X1 g0987(.A0(n1502), .A1(n1507), .B0(n1449), .B1(n1444), .Y(n1573));
  NOR3X1  g0988(.A(n1573), .B(n1406), .C(n1453), .Y(n1574));
  AOI22X1 g0989(.A0(n1502), .A1(n1507), .B0(n1449), .B1(n1444), .Y(n1575));
  NAND3X1 g0990(.A(n1572), .B(n1510), .C(n1452), .Y(n1576));
  NAND2X1 g0991(.A(n1576), .B(n1575), .Y(n1577));
  AOI21X1 g0992(.A0(n1577), .A1(n1572), .B0(n1574), .Y(n1578));
  XOR2X1  g0993(.A(n1578), .B(n1562), .Y(n1579));
  OAI22X1 g0994(.A0(n1570), .A1(n1116), .B0(n1097), .B1(n1579), .Y(n1580));
  INVX1   g0995(.A(n1579), .Y(n1581));
  AOI22X1 g0996(.A0(n1502), .A1(n992), .B0(n943), .B1(n1581), .Y(n1582));
  OAI21X1 g0997(.A0(n941), .A1(n931), .B0(n1581), .Y(n1583));
  NAND2X1 g0998(.A(n1583), .B(n1582), .Y(n1584));
  NAND4X1 g0999(.A(n1449), .B(n1424), .C(n1397), .D(n1507), .Y(n1585));
  XOR2X1  g1000(.A(n1561), .B(n1585), .Y(n1586));
  NOR2X1  g1001(.A(n902), .B(n1557), .Y(n1587));
  AOI21X1 g1002(.A0(n1559), .A1(n902), .B0(n1587), .Y(n1588));
  AOI22X1 g1003(.A0(n917), .A1(REG0_REG_13__SCAN_IN), .B0(REG2_REG_13__SCAN_IN), .B1(n952), .Y(n1589));
  NAND4X1 g1004(.A(REG3_REG_11__SCAN_IN), .B(REG3_REG_12__SCAN_IN), .C(REG3_REG_10__SCAN_IN), .D(n1431), .Y(n1590));
  XOR2X1  g1005(.A(n1590), .B(REG3_REG_13__SCAN_IN), .Y(n1591));
  INVX1   g1006(.A(n1591), .Y(n1592));
  AOI22X1 g1007(.A0(n955), .A1(n1592), .B0(n954), .B1(REG1_REG_13__SCAN_IN), .Y(n1593));
  NAND2X1 g1008(.A(n1593), .B(n1589), .Y(n1594));
  INVX1   g1009(.A(n1594), .Y(n1595));
  OAI22X1 g1010(.A0(n1588), .A1(n963), .B0(n1051), .B1(n1595), .Y(n1596));
  AOI21X1 g1011(.A0(n1586), .A1(n960), .B0(n1596), .Y(n1597));
  OAI21X1 g1012(.A0(n1570), .A1(n950), .B0(n1597), .Y(n1598));
  NOR4X1  g1013(.A(n1584), .B(n1580), .C(n1571), .D(n1598), .Y(n1599));
  NAND2X1 g1014(.A(n896), .B(REG0_REG_12__SCAN_IN), .Y(n1600));
  OAI21X1 g1015(.A0(n1599), .A1(n896), .B0(n1600), .Y(U3491));
  NAND2X1 g1016(.A(n759), .B(IR_REG_13__SCAN_IN), .Y(n1602));
  OAI21X1 g1017(.A0(n648), .A1(n759), .B0(n1602), .Y(n1603));
  INVX1   g1018(.A(DATAI_13_), .Y(n1604));
  NOR2X1  g1019(.A(n902), .B(n1604), .Y(n1605));
  AOI21X1 g1020(.A0(n1603), .A1(n902), .B0(n1605), .Y(n1606));
  XOR2X1  g1021(.A(n1606), .B(n1594), .Y(n1607));
  INVX1   g1022(.A(n1406), .Y(n1608));
  NOR2X1  g1023(.A(n1588), .B(n1567), .Y(n1609));
  NOR3X1  g1024(.A(n1573), .B(n1609), .C(n1453), .Y(n1610));
  AOI22X1 g1025(.A0(n1588), .A1(n1567), .B0(n1572), .B1(n1577), .Y(n1611));
  NOR2X1  g1026(.A(n1611), .B(n1609), .Y(n1612));
  AOI21X1 g1027(.A0(n1610), .A1(n1608), .B0(n1612), .Y(n1613));
  XOR2X1  g1028(.A(n1613), .B(n1607), .Y(n1614));
  INVX1   g1029(.A(n1614), .Y(n1615));
  OAI21X1 g1030(.A0(n941), .A1(n931), .B0(n1615), .Y(n1616));
  OAI21X1 g1031(.A0(n1614), .A1(n1097), .B0(n1616), .Y(n1617));
  NOR2X1  g1032(.A(n1588), .B(n1547), .Y(n1618));
  NAND2X1 g1033(.A(n1603), .B(n902), .Y(n1619));
  OAI21X1 g1034(.A0(n902), .A1(n1604), .B0(n1619), .Y(n1620));
  AOI22X1 g1035(.A0(n1595), .A1(n1606), .B0(n1588), .B1(n1547), .Y(n1621));
  INVX1   g1036(.A(n1621), .Y(n1622));
  AOI21X1 g1037(.A0(n1620), .A1(n1594), .B0(n1622), .Y(n1623));
  OAI21X1 g1038(.A0(n1618), .A1(n1556), .B0(n1623), .Y(n1624));
  INVX1   g1039(.A(n1556), .Y(n1625));
  AOI21X1 g1040(.A0(n1588), .A1(n1547), .B0(n1625), .Y(n1626));
  OAI21X1 g1041(.A0(n1588), .A1(n1547), .B0(n1607), .Y(n1627));
  OAI21X1 g1042(.A0(n1627), .A1(n1626), .B0(n1624), .Y(n1628));
  AOI22X1 g1043(.A0(n1567), .A1(n992), .B0(n943), .B1(n1615), .Y(n1629));
  OAI21X1 g1044(.A0(n1628), .A1(n1140), .B0(n1629), .Y(n1630));
  INVX1   g1045(.A(n1628), .Y(n1631));
  OAI21X1 g1046(.A0(n946), .A1(n945), .B0(n1631), .Y(n1632));
  INVX1   g1047(.A(n1632), .Y(n1633));
  NOR3X1  g1048(.A(n1561), .B(n1538), .C(n1514), .Y(n1634));
  XOR2X1  g1049(.A(n1634), .B(n1606), .Y(n1635));
  AOI22X1 g1050(.A0(n917), .A1(REG0_REG_14__SCAN_IN), .B0(REG2_REG_14__SCAN_IN), .B1(n952), .Y(n1636));
  INVX1   g1051(.A(n1636), .Y(n1637));
  INVX1   g1052(.A(REG1_REG_14__SCAN_IN), .Y(n1638));
  INVX1   g1053(.A(REG3_REG_14__SCAN_IN), .Y(n1639));
  INVX1   g1054(.A(REG3_REG_12__SCAN_IN), .Y(n1640));
  INVX1   g1055(.A(REG3_REG_13__SCAN_IN), .Y(n1641));
  NOR3X1  g1056(.A(n1544), .B(n1641), .C(n1640), .Y(n1642));
  XOR2X1  g1057(.A(n1642), .B(n1639), .Y(n1643));
  OAI22X1 g1058(.A0(n927), .A1(n1643), .B0(n926), .B1(n1638), .Y(n1644));
  NOR2X1  g1059(.A(n1644), .B(n1637), .Y(n1645));
  OAI22X1 g1060(.A0(n1606), .A1(n963), .B0(n1051), .B1(n1645), .Y(n1646));
  AOI21X1 g1061(.A0(n1635), .A1(n960), .B0(n1646), .Y(n1647));
  OAI21X1 g1062(.A0(n1628), .A1(n950), .B0(n1647), .Y(n1648));
  NOR4X1  g1063(.A(n1633), .B(n1630), .C(n1617), .D(n1648), .Y(n1649));
  NAND2X1 g1064(.A(n896), .B(REG0_REG_13__SCAN_IN), .Y(n1650));
  OAI21X1 g1065(.A0(n1649), .A1(n896), .B0(n1650), .Y(U3493));
  NAND3X1 g1066(.A(n1621), .B(n1514), .C(n1502), .Y(n1652));
  AOI22X1 g1067(.A0(n1594), .A1(n1620), .B0(n1561), .B1(n1567), .Y(n1653));
  AOI22X1 g1068(.A0(n1652), .A1(n1653), .B0(n1606), .B1(n1595), .Y(n1654));
  NOR3X1  g1069(.A(n1622), .B(n1554), .C(n1528), .Y(n1655));
  NOR2X1  g1070(.A(n1655), .B(n1654), .Y(n1656));
  INVX1   g1071(.A(DATAI_14_), .Y(n1657));
  NOR2X1  g1072(.A(IR_REG_31__SCAN_IN), .B(n651), .Y(n1658));
  INVX1   g1073(.A(n1658), .Y(n1659));
  OAI21X1 g1074(.A0(n652), .A1(n759), .B0(n1659), .Y(n1660));
  NAND2X1 g1075(.A(n1660), .B(n902), .Y(n1661));
  OAI21X1 g1076(.A0(n902), .A1(n1657), .B0(n1661), .Y(n1662));
  XOR2X1  g1077(.A(n3794), .B(n1656), .Y(n1665));
  AOI21X1 g1078(.A0(n1141), .A1(n1140), .B0(n1665), .Y(n1666));
  NOR2X1  g1079(.A(n1606), .B(n1594), .Y(n1667));
  INVX1   g1080(.A(n1667), .Y(n1668));
  NAND2X1 g1081(.A(n1610), .B(n1668), .Y(n1669));
  AOI21X1 g1082(.A0(n1593), .A1(n1589), .B0(n1620), .Y(n1670));
  AOI21X1 g1083(.A0(n1612), .A1(n1668), .B0(n1670), .Y(n1671));
  OAI21X1 g1084(.A0(n1669), .A1(n1406), .B0(n1671), .Y(n1672));
  XOR2X1  g1085(.A(n1672), .B(n3794), .Y(n1673));
  OAI22X1 g1086(.A0(n1665), .A1(n1116), .B0(n1097), .B1(n1673), .Y(n1674));
  INVX1   g1087(.A(n1673), .Y(n1675));
  AOI22X1 g1088(.A0(n1594), .A1(n992), .B0(n943), .B1(n1675), .Y(n1676));
  OAI21X1 g1089(.A0(n941), .A1(n931), .B0(n1675), .Y(n1677));
  NAND2X1 g1090(.A(n1677), .B(n1676), .Y(n1678));
  NOR4X1  g1091(.A(n1561), .B(n1538), .C(n1514), .D(n1620), .Y(n1679));
  NOR2X1  g1092(.A(n902), .B(n1657), .Y(n1680));
  AOI21X1 g1093(.A0(n1660), .A1(n902), .B0(n1680), .Y(n1681));
  XOR2X1  g1094(.A(n1681), .B(n1679), .Y(n1682));
  AOI22X1 g1095(.A0(n917), .A1(REG0_REG_15__SCAN_IN), .B0(REG2_REG_15__SCAN_IN), .B1(n952), .Y(n1683));
  INVX1   g1096(.A(REG1_REG_15__SCAN_IN), .Y(n1684));
  NAND2X1 g1097(.A(n1642), .B(REG3_REG_14__SCAN_IN), .Y(n1685));
  XOR2X1  g1098(.A(n1685), .B(REG3_REG_15__SCAN_IN), .Y(n1686));
  OAI22X1 g1099(.A0(n927), .A1(n1686), .B0(n926), .B1(n1684), .Y(n1687));
  INVX1   g1100(.A(n1687), .Y(n1688));
  NAND2X1 g1101(.A(n1688), .B(n1683), .Y(n1689));
  INVX1   g1102(.A(n1689), .Y(n1690));
  OAI22X1 g1103(.A0(n1681), .A1(n963), .B0(n1051), .B1(n1690), .Y(n1691));
  AOI21X1 g1104(.A0(n1682), .A1(n960), .B0(n1691), .Y(n1692));
  OAI21X1 g1105(.A0(n1665), .A1(n950), .B0(n1692), .Y(n1693));
  NOR4X1  g1106(.A(n1678), .B(n1674), .C(n1666), .D(n1693), .Y(n1694));
  NAND2X1 g1107(.A(n896), .B(REG0_REG_14__SCAN_IN), .Y(n1695));
  OAI21X1 g1108(.A0(n1694), .A1(n896), .B0(n1695), .Y(U3495));
  NOR2X1  g1109(.A(IR_REG_31__SCAN_IN), .B(n656), .Y(n1697));
  INVX1   g1110(.A(n1697), .Y(n1698));
  OAI21X1 g1111(.A0(n658), .A1(n759), .B0(n1698), .Y(n1699));
  INVX1   g1112(.A(DATAI_15_), .Y(n1700));
  NOR2X1  g1113(.A(n902), .B(n1700), .Y(n1701));
  AOI21X1 g1114(.A0(n1699), .A1(n902), .B0(n1701), .Y(n1702));
  XOR2X1  g1115(.A(n1702), .B(n1689), .Y(n1703));
  NOR3X1  g1116(.A(n1681), .B(n1644), .C(n1637), .Y(n1704));
  INVX1   g1117(.A(n1704), .Y(n1705));
  NOR2X1  g1118(.A(n1662), .B(n1645), .Y(n1706));
  AOI21X1 g1119(.A0(n1672), .A1(n1705), .B0(n1706), .Y(n1707));
  XOR2X1  g1120(.A(n1707), .B(n1703), .Y(n1708));
  NOR2X1  g1121(.A(n1708), .B(n942), .Y(n1709));
  INVX1   g1122(.A(n1645), .Y(n1710));
  AOI21X1 g1123(.A0(n1662), .A1(n1710), .B0(n1654), .Y(n1711));
  NOR3X1  g1124(.A(n1662), .B(n1644), .C(n1637), .Y(n1712));
  NOR2X1  g1125(.A(n1712), .B(n1711), .Y(n1713));
  NOR4X1  g1126(.A(n1622), .B(n1554), .C(n1528), .D(n1712), .Y(n1714));
  NOR2X1  g1127(.A(n1714), .B(n1713), .Y(n1715));
  XOR2X1  g1128(.A(n1715), .B(n1703), .Y(n1716));
  AOI22X1 g1129(.A0(n1710), .A1(n992), .B0(n945), .B1(n1716), .Y(n1717));
  OAI21X1 g1130(.A0(n946), .A1(n939), .B0(n1716), .Y(n1718));
  NAND2X1 g1131(.A(n1718), .B(n1717), .Y(n1719));
  NOR2X1  g1132(.A(n1708), .B(n1097), .Y(n1720));
  AOI21X1 g1133(.A0(n1086), .A1(n932), .B0(n1708), .Y(n1721));
  NOR4X1  g1134(.A(n1720), .B(n1719), .C(n1709), .D(n1721), .Y(n1722));
  INVX1   g1135(.A(n1722), .Y(n1723));
  NAND2X1 g1136(.A(n1716), .B(n949), .Y(n1724));
  NAND2X1 g1137(.A(n1681), .B(n1606), .Y(n1725));
  NOR4X1  g1138(.A(n1561), .B(n1538), .C(n1514), .D(n1725), .Y(n1726));
  XOR2X1  g1139(.A(n1726), .B(n1702), .Y(n1727));
  AOI22X1 g1140(.A0(n917), .A1(REG0_REG_16__SCAN_IN), .B0(REG2_REG_16__SCAN_IN), .B1(n952), .Y(n1728));
  INVX1   g1141(.A(REG1_REG_16__SCAN_IN), .Y(n1729));
  INVX1   g1142(.A(REG3_REG_16__SCAN_IN), .Y(n1730));
  NAND2X1 g1143(.A(REG3_REG_15__SCAN_IN), .B(REG3_REG_14__SCAN_IN), .Y(n1731));
  NOR4X1  g1144(.A(n1544), .B(n1641), .C(n1640), .D(n1731), .Y(n1732));
  XOR2X1  g1145(.A(n1732), .B(n1730), .Y(n1733));
  OAI22X1 g1146(.A0(n927), .A1(n1733), .B0(n926), .B1(n1729), .Y(n1734));
  INVX1   g1147(.A(n1734), .Y(n1735));
  NAND2X1 g1148(.A(n1735), .B(n1728), .Y(n1736));
  INVX1   g1149(.A(n1736), .Y(n1737));
  OAI22X1 g1150(.A0(n1702), .A1(n963), .B0(n1051), .B1(n1737), .Y(n1738));
  AOI21X1 g1151(.A0(n1727), .A1(n960), .B0(n1738), .Y(n1739));
  NAND2X1 g1152(.A(n1739), .B(n1724), .Y(n1740));
  NOR2X1  g1153(.A(n1740), .B(n1723), .Y(n1741));
  NAND2X1 g1154(.A(n896), .B(REG0_REG_15__SCAN_IN), .Y(n1742));
  OAI21X1 g1155(.A0(n1741), .A1(n896), .B0(n1742), .Y(U3497));
  INVX1   g1156(.A(n1702), .Y(n1744));
  OAI21X1 g1157(.A0(n1744), .A1(n1690), .B0(n1707), .Y(n1745));
  NOR2X1  g1158(.A(IR_REG_31__SCAN_IN), .B(n661), .Y(n1746));
  AOI21X1 g1159(.A0(n663), .A1(IR_REG_31__SCAN_IN), .B0(n1746), .Y(n1747));
  INVX1   g1160(.A(n1747), .Y(n1748));
  INVX1   g1161(.A(DATAI_16_), .Y(n1749));
  NOR2X1  g1162(.A(n902), .B(n1749), .Y(n1750));
  AOI21X1 g1163(.A0(n1748), .A1(n902), .B0(n1750), .Y(n1751));
  XOR2X1  g1164(.A(n1751), .B(n1736), .Y(n1752));
  AOI21X1 g1165(.A0(n1744), .A1(n1690), .B0(n1752), .Y(n1753));
  NAND2X1 g1166(.A(n1744), .B(n1690), .Y(n1754));
  INVX1   g1167(.A(n1707), .Y(n1755));
  AOI22X1 g1168(.A0(n1736), .A1(n1751), .B0(n1702), .B1(n1689), .Y(n1756));
  OAI21X1 g1169(.A0(n1751), .A1(n1736), .B0(n1756), .Y(n1757));
  AOI21X1 g1170(.A0(n1755), .A1(n1754), .B0(n1757), .Y(n1758));
  AOI21X1 g1171(.A0(n1753), .A1(n1745), .B0(n1758), .Y(n1759));
  NOR2X1  g1172(.A(n1759), .B(n942), .Y(n1760));
  NOR3X1  g1173(.A(n1712), .B(n1622), .C(n1554), .Y(n1761));
  NOR2X1  g1174(.A(n1744), .B(n1689), .Y(n1762));
  INVX1   g1175(.A(n1762), .Y(n1763));
  NAND2X1 g1176(.A(n1763), .B(n1761), .Y(n1764));
  AOI21X1 g1177(.A0(n1688), .A1(n1683), .B0(n1702), .Y(n1765));
  AOI21X1 g1178(.A0(n1763), .A1(n1713), .B0(n1765), .Y(n1766));
  OAI21X1 g1179(.A0(n1764), .A1(n1528), .B0(n1766), .Y(n1767));
  NOR2X1  g1180(.A(n1767), .B(n1752), .Y(n1768));
  INVX1   g1181(.A(n1751), .Y(n1769));
  XOR2X1  g1182(.A(n1769), .B(n1736), .Y(n1770));
  AOI21X1 g1183(.A0(n1752), .A1(n1767), .B0(n1768), .Y(n1772));
  INVX1   g1184(.A(n1772), .Y(n1773));
  AOI22X1 g1185(.A0(n1689), .A1(n992), .B0(n945), .B1(n1773), .Y(n1774));
  OAI21X1 g1186(.A0(n946), .A1(n939), .B0(n1773), .Y(n1775));
  NAND2X1 g1187(.A(n1775), .B(n1774), .Y(n1776));
  NOR2X1  g1188(.A(n1759), .B(n1097), .Y(n1777));
  AOI21X1 g1189(.A0(n1086), .A1(n932), .B0(n1759), .Y(n1778));
  NOR4X1  g1190(.A(n1777), .B(n1776), .C(n1760), .D(n1778), .Y(n1779));
  INVX1   g1191(.A(n1779), .Y(n1780));
  NAND2X1 g1192(.A(n1726), .B(n1702), .Y(n1781));
  XOR2X1  g1193(.A(n1769), .B(n1781), .Y(n1782));
  AOI22X1 g1194(.A0(n917), .A1(REG0_REG_17__SCAN_IN), .B0(REG2_REG_17__SCAN_IN), .B1(n952), .Y(n1783));
  INVX1   g1195(.A(REG1_REG_17__SCAN_IN), .Y(n1784));
  NAND2X1 g1196(.A(n1732), .B(REG3_REG_16__SCAN_IN), .Y(n1785));
  XOR2X1  g1197(.A(n1785), .B(REG3_REG_17__SCAN_IN), .Y(n1786));
  OAI22X1 g1198(.A0(n927), .A1(n1786), .B0(n926), .B1(n1784), .Y(n1787));
  INVX1   g1199(.A(n1787), .Y(n1788));
  NAND2X1 g1200(.A(n1788), .B(n1783), .Y(n1789));
  INVX1   g1201(.A(n1789), .Y(n1790));
  OAI22X1 g1202(.A0(n1751), .A1(n963), .B0(n1051), .B1(n1790), .Y(n1791));
  AOI21X1 g1203(.A0(n1782), .A1(n960), .B0(n1791), .Y(n1792));
  OAI21X1 g1204(.A0(n1772), .A1(n950), .B0(n1792), .Y(n1793));
  NOR2X1  g1205(.A(n1793), .B(n1780), .Y(n1794));
  NAND2X1 g1206(.A(n896), .B(REG0_REG_16__SCAN_IN), .Y(n1795));
  OAI21X1 g1207(.A0(n1794), .A1(n896), .B0(n1795), .Y(U3499));
  NAND2X1 g1208(.A(n1769), .B(n1736), .Y(n1797));
  INVX1   g1209(.A(n1797), .Y(n1798));
  NOR2X1  g1210(.A(n1798), .B(n1767), .Y(n1799));
  NOR2X1  g1211(.A(n670), .B(n759), .Y(n1800));
  NOR2X1  g1212(.A(IR_REG_31__SCAN_IN), .B(n667), .Y(n1801));
  NOR2X1  g1213(.A(n1801), .B(n1800), .Y(n1802));
  INVX1   g1214(.A(n1802), .Y(n1803));
  INVX1   g1215(.A(DATAI_17_), .Y(n1804));
  NOR2X1  g1216(.A(n902), .B(n1804), .Y(n1805));
  AOI21X1 g1217(.A0(n1803), .A1(n902), .B0(n1805), .Y(n1806));
  AOI22X1 g1218(.A0(n1790), .A1(n1806), .B0(n1751), .B1(n1737), .Y(n1807));
  OAI21X1 g1219(.A0(n1806), .A1(n1790), .B0(n1807), .Y(n1808));
  OAI21X1 g1220(.A0(n1769), .A1(n1736), .B0(n1767), .Y(n1809));
  XOR2X1  g1221(.A(n1806), .B(n1789), .Y(n1810));
  NAND3X1 g1222(.A(n1810), .B(n1809), .C(n1797), .Y(n1811));
  OAI21X1 g1223(.A0(n1808), .A1(n1799), .B0(n1811), .Y(n1812));
  INVX1   g1224(.A(n1812), .Y(n1813));
  AOI22X1 g1225(.A0(n1736), .A1(n992), .B0(n945), .B1(n1813), .Y(n1814));
  OAI21X1 g1226(.A0(n946), .A1(n939), .B0(n1813), .Y(n1815));
  NAND2X1 g1227(.A(n1769), .B(n1737), .Y(n1816));
  NAND3X1 g1228(.A(n1816), .B(n1754), .C(n1706), .Y(n1818));
  AOI21X1 g1229(.A0(n1818), .A1(n1756), .B0(n3825), .Y(n1819));
  NOR3X1  g1230(.A(n3825), .B(n3826), .C(n1704), .Y(n1821));
  AOI21X1 g1231(.A0(n1821), .A1(n1672), .B0(n1819), .Y(n1822));
  XOR2X1  g1232(.A(n1822), .B(n1810), .Y(n1823));
  INVX1   g1233(.A(n1823), .Y(n1824));
  OAI21X1 g1234(.A0(n943), .A1(n941), .B0(n1824), .Y(n1825));
  OAI21X1 g1235(.A0(n936), .A1(n931), .B0(n1824), .Y(n1826));
  NAND4X1 g1236(.A(n1825), .B(n1815), .C(n1814), .D(n1826), .Y(n1827));
  INVX1   g1237(.A(n1806), .Y(n1828));
  NAND3X1 g1238(.A(n1751), .B(n1726), .C(n1702), .Y(n1829));
  XOR2X1  g1239(.A(n1829), .B(n1828), .Y(n1830));
  AOI22X1 g1240(.A0(n917), .A1(REG0_REG_18__SCAN_IN), .B0(REG2_REG_18__SCAN_IN), .B1(n952), .Y(n1831));
  INVX1   g1241(.A(REG1_REG_18__SCAN_IN), .Y(n1832));
  NAND3X1 g1242(.A(n1732), .B(REG3_REG_17__SCAN_IN), .C(REG3_REG_16__SCAN_IN), .Y(n1833));
  XOR2X1  g1243(.A(n1833), .B(REG3_REG_18__SCAN_IN), .Y(n1834));
  OAI22X1 g1244(.A0(n927), .A1(n1834), .B0(n926), .B1(n1832), .Y(n1835));
  INVX1   g1245(.A(n1835), .Y(n1836));
  NAND2X1 g1246(.A(n1836), .B(n1831), .Y(n1837));
  INVX1   g1247(.A(n1837), .Y(n1838));
  OAI22X1 g1248(.A0(n1806), .A1(n963), .B0(n1051), .B1(n1838), .Y(n1839));
  AOI21X1 g1249(.A0(n1830), .A1(n960), .B0(n1839), .Y(n1840));
  OAI21X1 g1250(.A0(n1812), .A1(n950), .B0(n1840), .Y(n1841));
  NOR2X1  g1251(.A(n1841), .B(n1827), .Y(n1842));
  NAND2X1 g1252(.A(n896), .B(REG0_REG_17__SCAN_IN), .Y(n1843));
  OAI21X1 g1253(.A0(n1842), .A1(n896), .B0(n1843), .Y(U3501));
  AOI21X1 g1254(.A0(n1806), .A1(n1797), .B0(n1790), .Y(n1845));
  AOI21X1 g1255(.A0(n1828), .A1(n1798), .B0(n1845), .Y(n1846));
  INVX1   g1256(.A(n1846), .Y(n1847));
  AOI21X1 g1257(.A0(n1807), .A1(n1767), .B0(n1847), .Y(n1848));
  NOR2X1  g1258(.A(IR_REG_31__SCAN_IN), .B(n673), .Y(n1849));
  AOI21X1 g1259(.A0(n675), .A1(IR_REG_31__SCAN_IN), .B0(n1849), .Y(n1850));
  INVX1   g1260(.A(n1850), .Y(n1851));
  INVX1   g1261(.A(DATAI_18_), .Y(n1852));
  NOR2X1  g1262(.A(n902), .B(n1852), .Y(n1853));
  AOI21X1 g1263(.A0(n1851), .A1(n902), .B0(n1853), .Y(n1854));
  XOR2X1  g1264(.A(n1854), .B(n1837), .Y(n1855));
  INVX1   g1265(.A(n1855), .Y(n1856));
  INVX1   g1266(.A(n1854), .Y(n1857));
  NOR2X1  g1267(.A(n1856), .B(n1848), .Y(n1859));
  AOI21X1 g1268(.A0(n1856), .A1(n1848), .B0(n1859), .Y(n1860));
  AOI21X1 g1269(.A0(n1141), .A1(n1140), .B0(n1860), .Y(n1861));
  NOR2X1  g1270(.A(n1806), .B(n1789), .Y(n1862));
  NOR4X1  g1271(.A(n3825), .B(n3826), .C(n1704), .D(n1862), .Y(n1863));
  INVX1   g1272(.A(n1862), .Y(n1864));
  NOR2X1  g1273(.A(n1828), .B(n1790), .Y(n1865));
  AOI21X1 g1274(.A0(n1819), .A1(n1864), .B0(n1865), .Y(n1866));
  INVX1   g1275(.A(n1866), .Y(n1867));
  AOI21X1 g1276(.A0(n1863), .A1(n1672), .B0(n1867), .Y(n1868));
  XOR2X1  g1277(.A(n1868), .B(n1855), .Y(n1869));
  OAI22X1 g1278(.A0(n1860), .A1(n1116), .B0(n1097), .B1(n1869), .Y(n1870));
  INVX1   g1279(.A(n1869), .Y(n1871));
  AOI22X1 g1280(.A0(n1789), .A1(n992), .B0(n943), .B1(n1871), .Y(n1872));
  OAI21X1 g1281(.A0(n941), .A1(n931), .B0(n1871), .Y(n1873));
  NAND2X1 g1282(.A(n1873), .B(n1872), .Y(n1874));
  NAND4X1 g1283(.A(n1751), .B(n1726), .C(n1702), .D(n1806), .Y(n1875));
  XOR2X1  g1284(.A(n1857), .B(n1875), .Y(n1876));
  AOI22X1 g1285(.A0(n917), .A1(REG0_REG_19__SCAN_IN), .B0(REG2_REG_19__SCAN_IN), .B1(n952), .Y(n1877));
  INVX1   g1286(.A(REG3_REG_19__SCAN_IN), .Y(n1878));
  INVX1   g1287(.A(REG3_REG_18__SCAN_IN), .Y(n1879));
  NOR2X1  g1288(.A(n1833), .B(n1879), .Y(n1880));
  XOR2X1  g1289(.A(n1880), .B(n1878), .Y(n1881));
  INVX1   g1290(.A(n1881), .Y(n1882));
  AOI22X1 g1291(.A0(n955), .A1(n1882), .B0(n954), .B1(REG1_REG_19__SCAN_IN), .Y(n1883));
  NAND2X1 g1292(.A(n1883), .B(n1877), .Y(n1884));
  INVX1   g1293(.A(n1884), .Y(n1885));
  OAI22X1 g1294(.A0(n1854), .A1(n963), .B0(n1051), .B1(n1885), .Y(n1886));
  AOI21X1 g1295(.A0(n1876), .A1(n960), .B0(n1886), .Y(n1887));
  OAI21X1 g1296(.A0(n1860), .A1(n950), .B0(n1887), .Y(n1888));
  NOR4X1  g1297(.A(n1874), .B(n1870), .C(n1861), .D(n1888), .Y(n1889));
  NAND2X1 g1298(.A(n896), .B(REG0_REG_18__SCAN_IN), .Y(n1890));
  OAI21X1 g1299(.A0(n1889), .A1(n896), .B0(n1890), .Y(U3503));
  NOR2X1  g1300(.A(n1857), .B(n1837), .Y(n1892));
  NAND2X1 g1301(.A(n1857), .B(n1837), .Y(n1893));
  OAI21X1 g1302(.A0(n1892), .A1(n1848), .B0(n1893), .Y(n1894));
  INVX1   g1303(.A(DATAI_19_), .Y(n1895));
  NOR2X1  g1304(.A(n902), .B(n1895), .Y(n1896));
  AOI21X1 g1305(.A0(n902), .A1(n938), .B0(n1896), .Y(n1897));
  XOR2X1  g1306(.A(n1897), .B(n1884), .Y(n1898));
  NOR2X1  g1307(.A(n1894), .B(n1898), .Y(n1899));
  INVX1   g1308(.A(n1897), .Y(n1900));
  XOR2X1  g1309(.A(n1900), .B(n1884), .Y(n1901));
  AOI21X1 g1310(.A0(n1898), .A1(n1894), .B0(n1899), .Y(n1903));
  INVX1   g1311(.A(n1903), .Y(n1904));
  OAI21X1 g1312(.A0(n946), .A1(n939), .B0(n1904), .Y(n1905));
  NOR2X1  g1313(.A(n1854), .B(n1837), .Y(n1906));
  NOR2X1  g1314(.A(n1857), .B(n1838), .Y(n1907));
  INVX1   g1315(.A(n1907), .Y(n1908));
  OAI21X1 g1316(.A0(n1868), .A1(n1906), .B0(n1908), .Y(n1909));
  INVX1   g1317(.A(n1909), .Y(n1910));
  XOR2X1  g1318(.A(n1910), .B(n1898), .Y(n1911));
  INVX1   g1319(.A(n1911), .Y(n1912));
  AOI22X1 g1320(.A0(n1904), .A1(n945), .B0(n936), .B1(n1912), .Y(n1913));
  AOI22X1 g1321(.A0(n1837), .A1(n992), .B0(n943), .B1(n1912), .Y(n1914));
  OAI21X1 g1322(.A0(n941), .A1(n931), .B0(n1912), .Y(n1915));
  NAND4X1 g1323(.A(n1914), .B(n1913), .C(n1905), .D(n1915), .Y(n1916));
  NOR2X1  g1324(.A(n1857), .B(n1828), .Y(n1917));
  NAND4X1 g1325(.A(n1751), .B(n1726), .C(n1702), .D(n1917), .Y(n1918));
  XOR2X1  g1326(.A(n1918), .B(n1900), .Y(n1919));
  NOR3X1  g1327(.A(n1833), .B(n1879), .C(n1878), .Y(n1920));
  XOR2X1  g1328(.A(n1920), .B(REG3_REG_20__SCAN_IN), .Y(n1921));
  NAND2X1 g1329(.A(n1921), .B(n955), .Y(n1922));
  NAND3X1 g1330(.A(n983), .B(n925), .C(REG1_REG_20__SCAN_IN), .Y(n1923));
  AOI22X1 g1331(.A0(n917), .A1(REG0_REG_20__SCAN_IN), .B0(REG2_REG_20__SCAN_IN), .B1(n952), .Y(n1924));
  NAND3X1 g1332(.A(n1924), .B(n1923), .C(n1922), .Y(n1925));
  INVX1   g1333(.A(n1925), .Y(n1926));
  OAI22X1 g1334(.A0(n1897), .A1(n963), .B0(n1051), .B1(n1926), .Y(n1927));
  AOI21X1 g1335(.A0(n1919), .A1(n960), .B0(n1927), .Y(n1928));
  OAI21X1 g1336(.A0(n1903), .A1(n950), .B0(n1928), .Y(n1929));
  NOR2X1  g1337(.A(n1929), .B(n1916), .Y(n1930));
  NAND2X1 g1338(.A(n896), .B(REG0_REG_19__SCAN_IN), .Y(n1931));
  OAI21X1 g1339(.A0(n1930), .A1(n896), .B0(n1931), .Y(U3505));
  AOI21X1 g1340(.A0(n1883), .A1(n1877), .B0(n1897), .Y(n1933));
  INVX1   g1341(.A(DATAI_20_), .Y(n1934));
  NOR2X1  g1342(.A(n902), .B(n1934), .Y(n1935));
  OAI22X1 g1343(.A0(n1925), .A1(n1935), .B0(n1900), .B1(n1884), .Y(n1936));
  AOI21X1 g1344(.A0(n1935), .A1(n1925), .B0(n1936), .Y(n1937));
  OAI21X1 g1345(.A0(n1933), .A1(n1894), .B0(n1937), .Y(n1938));
  INVX1   g1346(.A(n1933), .Y(n1939));
  OAI21X1 g1347(.A0(n1900), .A1(n1884), .B0(n1894), .Y(n1940));
  INVX1   g1348(.A(n1935), .Y(n1941));
  XOR2X1  g1349(.A(n1941), .B(n1925), .Y(n1942));
  NAND3X1 g1350(.A(n1942), .B(n1940), .C(n1939), .Y(n1943));
  NAND2X1 g1351(.A(n1943), .B(n1938), .Y(n1944));
  INVX1   g1352(.A(n1944), .Y(n1945));
  AOI22X1 g1353(.A0(n1884), .A1(n992), .B0(n945), .B1(n1945), .Y(n1946));
  OAI21X1 g1354(.A0(n946), .A1(n939), .B0(n1945), .Y(n1947));
  NOR2X1  g1355(.A(n1897), .B(n1884), .Y(n1948));
  AOI21X1 g1356(.A0(n1883), .A1(n1877), .B0(n1900), .Y(n1949));
  INVX1   g1357(.A(n1949), .Y(n1950));
  OAI21X1 g1358(.A0(n1910), .A1(n1948), .B0(n1950), .Y(n1951));
  XOR2X1  g1359(.A(n1951), .B(n1942), .Y(n1952));
  OAI21X1 g1360(.A0(n943), .A1(n941), .B0(n1952), .Y(n1953));
  OAI21X1 g1361(.A0(n936), .A1(n931), .B0(n1952), .Y(n1954));
  NAND4X1 g1362(.A(n1953), .B(n1947), .C(n1946), .D(n1954), .Y(n1955));
  NOR2X1  g1363(.A(n1918), .B(n1900), .Y(n1956));
  XOR2X1  g1364(.A(n1941), .B(n1956), .Y(n1957));
  INVX1   g1365(.A(REG3_REG_20__SCAN_IN), .Y(n1958));
  NOR4X1  g1366(.A(n1879), .B(n1958), .C(n1878), .D(n1833), .Y(n1959));
  XOR2X1  g1367(.A(n1959), .B(REG3_REG_21__SCAN_IN), .Y(n1960));
  NAND2X1 g1368(.A(n1960), .B(n955), .Y(n1961));
  NAND3X1 g1369(.A(n983), .B(n925), .C(REG1_REG_21__SCAN_IN), .Y(n1962));
  AOI22X1 g1370(.A0(n917), .A1(REG0_REG_21__SCAN_IN), .B0(REG2_REG_21__SCAN_IN), .B1(n952), .Y(n1963));
  NAND3X1 g1371(.A(n1963), .B(n1962), .C(n1961), .Y(n1964));
  INVX1   g1372(.A(n1964), .Y(n1965));
  OAI22X1 g1373(.A0(n1941), .A1(n963), .B0(n1051), .B1(n1965), .Y(n1966));
  AOI21X1 g1374(.A0(n1957), .A1(n960), .B0(n1966), .Y(n1967));
  OAI21X1 g1375(.A0(n1944), .A1(n950), .B0(n1967), .Y(n1968));
  NOR2X1  g1376(.A(n1968), .B(n1955), .Y(n1969));
  NAND2X1 g1377(.A(n896), .B(REG0_REG_20__SCAN_IN), .Y(n1970));
  OAI21X1 g1378(.A0(n1969), .A1(n896), .B0(n1970), .Y(U3506));
  INVX1   g1379(.A(DATAI_21_), .Y(n1972));
  NOR2X1  g1380(.A(n902), .B(n1972), .Y(n1973));
  INVX1   g1381(.A(n1973), .Y(n1974));
  XOR2X1  g1382(.A(n1974), .B(n1964), .Y(n1975));
  INVX1   g1383(.A(n1936), .Y(n1976));
  AOI21X1 g1384(.A0(n1935), .A1(n1933), .B0(n1925), .Y(n1977));
  AOI21X1 g1385(.A0(n1941), .A1(n1939), .B0(n1977), .Y(n1978));
  AOI21X1 g1386(.A0(n1976), .A1(n1894), .B0(n1978), .Y(n1979));
  NAND2X1 g1387(.A(n1976), .B(n1894), .Y(n1980));
  NOR2X1  g1388(.A(n1974), .B(n1964), .Y(n1981));
  NOR2X1  g1389(.A(n1973), .B(n1965), .Y(n1982));
  NOR3X1  g1390(.A(n1978), .B(n1982), .C(n1981), .Y(n1983));
  NAND2X1 g1391(.A(n1983), .B(n1980), .Y(n1984));
  OAI21X1 g1392(.A0(n1979), .A1(n1975), .B0(n1984), .Y(n1985));
  AOI21X1 g1393(.A0(n1141), .A1(n1140), .B0(n1985), .Y(n1986));
  NOR2X1  g1394(.A(n1941), .B(n1925), .Y(n1987));
  INVX1   g1395(.A(n1987), .Y(n1988));
  NOR2X1  g1396(.A(n1935), .B(n1926), .Y(n1989));
  AOI21X1 g1397(.A0(n1988), .A1(n1949), .B0(n1989), .Y(n1990));
  INVX1   g1398(.A(n1990), .Y(n1991));
  NOR2X1  g1399(.A(n1987), .B(n1948), .Y(n1992));
  AOI21X1 g1400(.A0(n1992), .A1(n1909), .B0(n1991), .Y(n1993));
  XOR2X1  g1401(.A(n1993), .B(n1975), .Y(n1994));
  OAI22X1 g1402(.A0(n1985), .A1(n1116), .B0(n1097), .B1(n1994), .Y(n1995));
  NOR2X1  g1403(.A(n1995), .B(n1986), .Y(n1996));
  INVX1   g1404(.A(n1994), .Y(n1997));
  AOI22X1 g1405(.A0(n1925), .A1(n992), .B0(n943), .B1(n1997), .Y(n1998));
  OAI21X1 g1406(.A0(n941), .A1(n931), .B0(n1997), .Y(n1999));
  NAND3X1 g1407(.A(n1999), .B(n1998), .C(n1996), .Y(n2000));
  NOR3X1  g1408(.A(n1935), .B(n1918), .C(n1900), .Y(n2001));
  XOR2X1  g1409(.A(n2001), .B(n1974), .Y(n2002));
  INVX1   g1410(.A(REG3_REG_22__SCAN_IN), .Y(n2003));
  NAND2X1 g1411(.A(n1959), .B(REG3_REG_21__SCAN_IN), .Y(n2004));
  XOR2X1  g1412(.A(n2004), .B(n2003), .Y(n2005));
  NAND3X1 g1413(.A(n983), .B(n925), .C(REG1_REG_22__SCAN_IN), .Y(n2006));
  AOI22X1 g1414(.A0(n917), .A1(REG0_REG_22__SCAN_IN), .B0(REG2_REG_22__SCAN_IN), .B1(n952), .Y(n2007));
  NAND2X1 g1415(.A(n2007), .B(n2006), .Y(n2008));
  AOI21X1 g1416(.A0(n2005), .A1(n955), .B0(n2008), .Y(n2009));
  OAI22X1 g1417(.A0(n1974), .A1(n963), .B0(n1051), .B1(n2009), .Y(n2010));
  AOI21X1 g1418(.A0(n2002), .A1(n960), .B0(n2010), .Y(n2011));
  OAI21X1 g1419(.A0(n1985), .A1(n950), .B0(n2011), .Y(n2012));
  NOR2X1  g1420(.A(n2012), .B(n2000), .Y(n2013));
  NAND2X1 g1421(.A(n896), .B(REG0_REG_21__SCAN_IN), .Y(n2014));
  OAI21X1 g1422(.A0(n2013), .A1(n896), .B0(n2014), .Y(U3507));
  INVX1   g1423(.A(DATAI_22_), .Y(n2016));
  NOR2X1  g1424(.A(n902), .B(n2016), .Y(n2017));
  XOR2X1  g1425(.A(n2017), .B(n2009), .Y(n2018));
  OAI21X1 g1426(.A0(n1993), .A1(n1981), .B0(n3876), .Y(n2020));
  INVX1   g1427(.A(n2020), .Y(n2021));
  XOR2X1  g1428(.A(n2021), .B(n2018), .Y(n2022));
  NOR2X1  g1429(.A(n2022), .B(n942), .Y(n2023));
  INVX1   g1430(.A(n1981), .Y(n2024));
  NAND3X1 g1431(.A(n1992), .B(n2024), .C(n1909), .Y(n2025));
  NOR2X1  g1432(.A(n1990), .B(n1981), .Y(n2026));
  NOR2X1  g1433(.A(n2026), .B(n1982), .Y(n2027));
  XOR2X1  g1434(.A(n2020), .B(n2018), .Y(n2029));
  NAND2X1 g1435(.A(n2029), .B(n941), .Y(n2030));
  NOR2X1  g1436(.A(n1973), .B(n1964), .Y(n2031));
  NOR3X1  g1437(.A(n2031), .B(n1936), .C(n1892), .Y(n2032));
  INVX1   g1438(.A(n2032), .Y(n2033));
  NOR3X1  g1439(.A(n2031), .B(n1936), .C(n1893), .Y(n2034));
  NOR2X1  g1440(.A(n1974), .B(n1965), .Y(n2035));
  NOR3X1  g1441(.A(n2035), .B(n2034), .C(n1978), .Y(n2036));
  OAI22X1 g1442(.A0(n2033), .A1(n1846), .B0(n2031), .B1(n2036), .Y(n2037));
  NAND2X1 g1443(.A(n2032), .B(n1807), .Y(n2038));
  INVX1   g1444(.A(n2038), .Y(n2039));
  AOI21X1 g1445(.A0(n2039), .A1(n1767), .B0(n2037), .Y(n2040));
  XOR2X1  g1446(.A(n2040), .B(n2018), .Y(n2041));
  AOI22X1 g1447(.A0(n1964), .A1(n992), .B0(n945), .B1(n2041), .Y(n2042));
  OAI21X1 g1448(.A0(n946), .A1(n939), .B0(n2041), .Y(n2043));
  NAND3X1 g1449(.A(n2043), .B(n2042), .C(n2030), .Y(n2044));
  AOI21X1 g1450(.A0(n1097), .A1(n932), .B0(n2022), .Y(n2045));
  NOR4X1  g1451(.A(n1935), .B(n1918), .C(n1900), .D(n1973), .Y(n2046));
  INVX1   g1452(.A(n2017), .Y(n2047));
  XOR2X1  g1453(.A(n2047), .B(n2046), .Y(n2048));
  NAND2X1 g1454(.A(n2048), .B(n960), .Y(n2049));
  INVX1   g1455(.A(REG3_REG_23__SCAN_IN), .Y(n2050));
  NAND3X1 g1456(.A(n1959), .B(REG3_REG_22__SCAN_IN), .C(REG3_REG_21__SCAN_IN), .Y(n2051));
  XOR2X1  g1457(.A(n2051), .B(n2050), .Y(n2052));
  NAND3X1 g1458(.A(n983), .B(n925), .C(REG1_REG_23__SCAN_IN), .Y(n2053));
  AOI22X1 g1459(.A0(n917), .A1(REG0_REG_23__SCAN_IN), .B0(REG2_REG_23__SCAN_IN), .B1(n952), .Y(n2054));
  NAND2X1 g1460(.A(n2054), .B(n2053), .Y(n2055));
  AOI21X1 g1461(.A0(n2052), .A1(n955), .B0(n2055), .Y(n2056));
  OAI22X1 g1462(.A0(n2047), .A1(n963), .B0(n1051), .B1(n2056), .Y(n2057));
  AOI21X1 g1463(.A0(n2041), .A1(n949), .B0(n2057), .Y(n2058));
  NAND2X1 g1464(.A(n2058), .B(n2049), .Y(n2059));
  NOR4X1  g1465(.A(n2045), .B(n2044), .C(n2023), .D(n2059), .Y(n2060));
  NAND2X1 g1466(.A(n896), .B(REG0_REG_22__SCAN_IN), .Y(n2061));
  OAI21X1 g1467(.A0(n2060), .A1(n896), .B0(n2061), .Y(U3508));
  NOR2X1  g1468(.A(n2017), .B(n2009), .Y(n2063));
  INVX1   g1469(.A(n2063), .Y(n2064));
  INVX1   g1470(.A(DATAI_23_), .Y(n2065));
  NOR2X1  g1471(.A(n902), .B(n2065), .Y(n2066));
  XOR2X1  g1472(.A(n2066), .B(n2056), .Y(n2067));
  AOI21X1 g1473(.A0(n2017), .A1(n2009), .B0(n2067), .Y(n2068));
  INVX1   g1474(.A(n2068), .Y(n2069));
  AOI21X1 g1475(.A0(n2021), .A1(n2064), .B0(n2069), .Y(n2070));
  INVX1   g1476(.A(n2056), .Y(n2071));
  INVX1   g1477(.A(n2066), .Y(n2072));
  NOR2X1  g1478(.A(n2072), .B(n2071), .Y(n2073));
  AOI21X1 g1479(.A0(n2072), .A1(n2071), .B0(n2063), .Y(n2074));
  INVX1   g1480(.A(n2074), .Y(n2075));
  INVX1   g1481(.A(n2009), .Y(n2076));
  NOR2X1  g1482(.A(n2047), .B(n2076), .Y(n2077));
  NOR2X1  g1483(.A(n2021), .B(n2077), .Y(n2078));
  NOR3X1  g1484(.A(n2078), .B(n2075), .C(n2073), .Y(n2079));
  OAI21X1 g1485(.A0(n2079), .A1(n2070), .B0(n931), .Y(n2080));
  NOR2X1  g1486(.A(n2075), .B(n2073), .Y(n2081));
  NAND3X1 g1487(.A(n2081), .B(n2027), .C(n2025), .Y(n2082));
  NAND2X1 g1488(.A(n2068), .B(n2020), .Y(n2083));
  INVX1   g1489(.A(n2067), .Y(n2084));
  NAND3X1 g1490(.A(n2092), .B(n2083), .C(n2082), .Y(n2086));
  NAND2X1 g1491(.A(n2086), .B(n941), .Y(n2087));
  INVX1   g1492(.A(n1993), .Y(n2088));
  NAND3X1 g1493(.A(n2068), .B(n2088), .C(n2024), .Y(n2089));
  NOR4X1  g1494(.A(n2073), .B(n2026), .C(n1982), .D(n2075), .Y(n2090));
  NOR3X1  g1495(.A(n2073), .B(n2047), .C(n2076), .Y(n2091));
  AOI22X1 g1496(.A0(n2074), .A1(n2091), .B0(n2084), .B1(n2063), .Y(n2092));
  OAI21X1 g1497(.A0(n2069), .A1(n3876), .B0(n2092), .Y(n2093));
  AOI21X1 g1498(.A0(n2090), .A1(n2025), .B0(n2093), .Y(n2094));
  AOI21X1 g1499(.A0(n2094), .A1(n2089), .B0(n1097), .Y(n2095));
  AOI21X1 g1500(.A0(n2094), .A1(n2089), .B0(n942), .Y(n2096));
  NOR2X1  g1501(.A(n2017), .B(n2076), .Y(n2097));
  NOR2X1  g1502(.A(n2097), .B(n2038), .Y(n2098));
  NAND2X1 g1503(.A(n2017), .B(n2076), .Y(n2099));
  OAI21X1 g1504(.A0(n2017), .A1(n2076), .B0(n2037), .Y(n2100));
  NAND2X1 g1505(.A(n2100), .B(n2099), .Y(n2101));
  AOI21X1 g1506(.A0(n2098), .A1(n1767), .B0(n2101), .Y(n2102));
  XOR2X1  g1507(.A(n2102), .B(n2084), .Y(n2103));
  OAI22X1 g1508(.A0(n2009), .A1(n1117), .B0(n1116), .B1(n2103), .Y(n2104));
  AOI21X1 g1509(.A0(n1141), .A1(n1140), .B0(n2103), .Y(n2105));
  NOR4X1  g1510(.A(n2104), .B(n2096), .C(n2095), .D(n2105), .Y(n2106));
  NAND3X1 g1511(.A(n2106), .B(n2087), .C(n2080), .Y(n2107));
  OAI21X1 g1512(.A0(n2097), .A1(n2040), .B0(n2099), .Y(n2108));
  NAND3X1 g1513(.A(n2047), .B(n2001), .C(n1974), .Y(n2110));
  XOR2X1  g1514(.A(n2110), .B(n2066), .Y(n2111));
  INVX1   g1515(.A(REG3_REG_24__SCAN_IN), .Y(n2112));
  NAND4X1 g1516(.A(REG3_REG_22__SCAN_IN), .B(REG3_REG_21__SCAN_IN), .C(REG3_REG_23__SCAN_IN), .D(n1959), .Y(n2113));
  XOR2X1  g1517(.A(n2113), .B(n2112), .Y(n2114));
  NAND3X1 g1518(.A(n983), .B(n925), .C(REG1_REG_24__SCAN_IN), .Y(n2115));
  AOI22X1 g1519(.A0(n917), .A1(REG0_REG_24__SCAN_IN), .B0(REG2_REG_24__SCAN_IN), .B1(n952), .Y(n2116));
  NAND2X1 g1520(.A(n2116), .B(n2115), .Y(n2117));
  AOI21X1 g1521(.A0(n2114), .A1(n955), .B0(n2117), .Y(n2118));
  OAI22X1 g1522(.A0(n2072), .A1(n963), .B0(n1051), .B1(n2118), .Y(n2119));
  AOI21X1 g1523(.A0(n2111), .A1(n960), .B0(n2119), .Y(n2120));
  OAI21X1 g1524(.A0(n2103), .A1(n950), .B0(n2120), .Y(n2121));
  NOR2X1  g1525(.A(n2121), .B(n2107), .Y(n2122));
  NAND2X1 g1526(.A(n896), .B(REG0_REG_23__SCAN_IN), .Y(n2123));
  OAI21X1 g1527(.A0(n2122), .A1(n896), .B0(n2123), .Y(U3509));
  INVX1   g1528(.A(DATAI_24_), .Y(n2125));
  NOR2X1  g1529(.A(n902), .B(n2125), .Y(n2126));
  XOR2X1  g1530(.A(n2126), .B(n2118), .Y(n2127));
  AOI22X1 g1531(.A0(n2056), .A1(n2066), .B0(n2017), .B1(n2009), .Y(n2128));
  INVX1   g1532(.A(n2128), .Y(n2129));
  NOR2X1  g1533(.A(n2129), .B(n1981), .Y(n2130));
  NAND3X1 g1534(.A(n2128), .B(n1974), .C(n1964), .Y(n2131));
  AOI21X1 g1535(.A0(n2131), .A1(n2074), .B0(n2073), .Y(n2132));
  AOI21X1 g1536(.A0(n2130), .A1(n1991), .B0(n2132), .Y(n2133));
  INVX1   g1537(.A(n2133), .Y(n2134));
  NOR4X1  g1538(.A(n1981), .B(n1987), .C(n1948), .D(n2129), .Y(n2135));
  AOI21X1 g1539(.A0(n2135), .A1(n1909), .B0(n2134), .Y(n2136));
  XOR2X1  g1540(.A(n2136), .B(n2127), .Y(n2137));
  NOR2X1  g1541(.A(n2137), .B(n942), .Y(n2138));
  NOR2X1  g1542(.A(n2072), .B(n2056), .Y(n2139));
  INVX1   g1543(.A(n2139), .Y(n2140));
  NOR2X1  g1544(.A(n2066), .B(n2071), .Y(n2141));
  OAI21X1 g1545(.A0(n2141), .A1(n2102), .B0(n2140), .Y(n2142));
  NOR2X1  g1546(.A(n2142), .B(n2127), .Y(n2143));
  AOI21X1 g1547(.A0(n2127), .A1(n2142), .B0(n2143), .Y(n2145));
  OAI22X1 g1548(.A0(n2056), .A1(n1117), .B0(n1116), .B1(n2145), .Y(n2146));
  AOI21X1 g1549(.A0(n1141), .A1(n1140), .B0(n2145), .Y(n2147));
  NOR3X1  g1550(.A(n2147), .B(n2146), .C(n2138), .Y(n2148));
  NOR2X1  g1551(.A(n2137), .B(n1097), .Y(n2149));
  AOI21X1 g1552(.A0(n1086), .A1(n932), .B0(n2137), .Y(n2150));
  NOR2X1  g1553(.A(n2150), .B(n2149), .Y(n2151));
  NAND2X1 g1554(.A(n2151), .B(n2148), .Y(n2152));
  INVX1   g1555(.A(n2141), .Y(n2154));
  AOI21X1 g1556(.A0(n2154), .A1(n2108), .B0(n2139), .Y(n2155));
  INVX1   g1557(.A(n2126), .Y(n2156));
  XOR2X1  g1558(.A(n2156), .B(n2118), .Y(n2157));
  NAND4X1 g1559(.A(n2047), .B(n2001), .C(n1974), .D(n2072), .Y(n2160));
  XOR2X1  g1560(.A(n2126), .B(n2160), .Y(n2161));
  INVX1   g1561(.A(REG3_REG_25__SCAN_IN), .Y(n2162));
  NOR2X1  g1562(.A(n2113), .B(n2112), .Y(n2163));
  XOR2X1  g1563(.A(n2163), .B(n2162), .Y(n2164));
  INVX1   g1564(.A(n2164), .Y(n2165));
  AOI22X1 g1565(.A0(n917), .A1(REG0_REG_25__SCAN_IN), .B0(REG2_REG_25__SCAN_IN), .B1(n952), .Y(n2166));
  INVX1   g1566(.A(n2166), .Y(n2167));
  AOI21X1 g1567(.A0(n954), .A1(REG1_REG_25__SCAN_IN), .B0(n2167), .Y(n2168));
  INVX1   g1568(.A(n2168), .Y(n2169));
  AOI21X1 g1569(.A0(n2165), .A1(n955), .B0(n2169), .Y(n2170));
  OAI22X1 g1570(.A0(n2156), .A1(n963), .B0(n1051), .B1(n2170), .Y(n2171));
  AOI21X1 g1571(.A0(n2161), .A1(n960), .B0(n2171), .Y(n2172));
  OAI21X1 g1572(.A0(n2145), .A1(n950), .B0(n2172), .Y(n2173));
  NOR2X1  g1573(.A(n2173), .B(n2152), .Y(n2174));
  NAND2X1 g1574(.A(n896), .B(REG0_REG_24__SCAN_IN), .Y(n2175));
  OAI21X1 g1575(.A0(n2174), .A1(n896), .B0(n2175), .Y(U3510));
  INVX1   g1576(.A(DATAI_25_), .Y(n2177));
  NOR2X1  g1577(.A(n902), .B(n2177), .Y(n2178));
  XOR2X1  g1578(.A(n2178), .B(n2170), .Y(n2179));
  INVX1   g1579(.A(n2118), .Y(n2181));
  NOR2X1  g1580(.A(n2126), .B(n2181), .Y(n2182));
  INVX1   g1581(.A(n2182), .Y(n2183));
  NOR2X1  g1582(.A(n2156), .B(n2118), .Y(n2184));
  AOI21X1 g1583(.A0(n2183), .A1(n2142), .B0(n2184), .Y(n2185));
  INVX1   g1584(.A(n2178), .Y(n2186));
  XOR2X1  g1585(.A(n2186), .B(n2170), .Y(n2187));
  NOR2X1  g1586(.A(n2187), .B(n2185), .Y(n2188));
  AOI21X1 g1587(.A0(n2185), .A1(n2187), .B0(n2188), .Y(n2189));
  INVX1   g1588(.A(n2189), .Y(n2190));
  OAI21X1 g1589(.A0(n946), .A1(n939), .B0(n2190), .Y(n2191));
  NOR2X1  g1590(.A(n2156), .B(n2181), .Y(n2192));
  NOR2X1  g1591(.A(n2126), .B(n2118), .Y(n2193));
  INVX1   g1592(.A(n2193), .Y(n2194));
  OAI21X1 g1593(.A0(n2133), .A1(n2192), .B0(n2194), .Y(n2195));
  INVX1   g1594(.A(n2192), .Y(n2196));
  NAND2X1 g1595(.A(n2135), .B(n2196), .Y(n2197));
  INVX1   g1596(.A(n2197), .Y(n2198));
  AOI21X1 g1597(.A0(n2198), .A1(n1909), .B0(n2195), .Y(n2199));
  XOR2X1  g1598(.A(n2199), .B(n2179), .Y(n2200));
  INVX1   g1599(.A(n2200), .Y(n2201));
  AOI22X1 g1600(.A0(n2190), .A1(n945), .B0(n936), .B1(n2201), .Y(n2202));
  AOI22X1 g1601(.A0(n2181), .A1(n992), .B0(n943), .B1(n2201), .Y(n2203));
  OAI21X1 g1602(.A0(n941), .A1(n931), .B0(n2201), .Y(n2204));
  NAND4X1 g1603(.A(n2203), .B(n2202), .C(n2191), .D(n2204), .Y(n2205));
  INVX1   g1604(.A(n2184), .Y(n2206));
  OAI21X1 g1605(.A0(n2155), .A1(n2182), .B0(n2206), .Y(n2207));
  NOR2X1  g1606(.A(n2189), .B(n950), .Y(n2211));
  NOR3X1  g1607(.A(n2126), .B(n2110), .C(n2066), .Y(n2212));
  XOR2X1  g1608(.A(n2212), .B(n2186), .Y(n2213));
  NAND2X1 g1609(.A(n2213), .B(n960), .Y(n2214));
  INVX1   g1610(.A(REG3_REG_26__SCAN_IN), .Y(n2215));
  NOR3X1  g1611(.A(n2113), .B(n2112), .C(n2162), .Y(n2216));
  XOR2X1  g1612(.A(n2216), .B(n2215), .Y(n2217));
  AOI22X1 g1613(.A0(n917), .A1(REG0_REG_26__SCAN_IN), .B0(REG2_REG_26__SCAN_IN), .B1(n952), .Y(n2218));
  INVX1   g1614(.A(n2218), .Y(n2219));
  AOI21X1 g1615(.A0(n954), .A1(REG1_REG_26__SCAN_IN), .B0(n2219), .Y(n2220));
  OAI21X1 g1616(.A0(n2217), .A1(n927), .B0(n2220), .Y(n2221));
  AOI22X1 g1617(.A0(n2178), .A1(n962), .B0(n951), .B1(n2221), .Y(n2222));
  NAND2X1 g1618(.A(n2222), .B(n2214), .Y(n2223));
  NOR3X1  g1619(.A(n2223), .B(n2211), .C(n2205), .Y(n2224));
  NAND2X1 g1620(.A(n896), .B(REG0_REG_25__SCAN_IN), .Y(n2225));
  OAI21X1 g1621(.A0(n2224), .A1(n896), .B0(n2225), .Y(U3511));
  OAI21X1 g1622(.A0(n2186), .A1(n2170), .B0(n2185), .Y(n2227));
  INVX1   g1623(.A(DATAI_26_), .Y(n2228));
  NOR2X1  g1624(.A(n902), .B(n2228), .Y(n2229));
  INVX1   g1625(.A(n2170), .Y(n2230));
  OAI22X1 g1626(.A0(n2221), .A1(n2229), .B0(n2178), .B1(n2230), .Y(n2231));
  AOI21X1 g1627(.A0(n2229), .A1(n2221), .B0(n2231), .Y(n2232));
  INVX1   g1628(.A(n2229), .Y(n2233));
  XOR2X1  g1629(.A(n2233), .B(n2221), .Y(n2234));
  OAI21X1 g1630(.A0(n2186), .A1(n2170), .B0(n2234), .Y(n2235));
  NOR2X1  g1631(.A(n2178), .B(n2230), .Y(n2236));
  NOR2X1  g1632(.A(n2236), .B(n2185), .Y(n2237));
  NOR2X1  g1633(.A(n2237), .B(n2235), .Y(n2238));
  AOI21X1 g1634(.A0(n2232), .A1(n2227), .B0(n2238), .Y(n2239));
  NAND2X1 g1635(.A(n2239), .B(n945), .Y(n2240));
  OAI21X1 g1636(.A0(n946), .A1(n939), .B0(n2239), .Y(n2241));
  NOR2X1  g1637(.A(n2186), .B(n2230), .Y(n2242));
  NOR2X1  g1638(.A(n2178), .B(n2170), .Y(n2243));
  INVX1   g1639(.A(n2243), .Y(n2244));
  OAI21X1 g1640(.A0(n2199), .A1(n2242), .B0(n2244), .Y(n2245));
  INVX1   g1641(.A(n2245), .Y(n2246));
  XOR2X1  g1642(.A(n2246), .B(n2234), .Y(n2247));
  NOR2X1  g1643(.A(n2247), .B(n1086), .Y(n2248));
  OAI22X1 g1644(.A0(n2170), .A1(n1117), .B0(n942), .B1(n2247), .Y(n2254));
  AOI21X1 g1645(.A0(n1097), .A1(n932), .B0(n2247), .Y(n2255));
  NOR3X1  g1646(.A(n2255), .B(n2254), .C(n2248), .Y(n2256));
  NAND3X1 g1647(.A(n2256), .B(n2241), .C(n2240), .Y(n2257));
  NOR2X1  g1648(.A(n2186), .B(n2170), .Y(n2258));
  NOR2X1  g1649(.A(n2229), .B(n2221), .Y(n2259));
  OAI21X1 g1650(.A0(n2207), .A1(n2258), .B0(n2232), .Y(n2263));
  OAI21X1 g1651(.A0(n2237), .A1(n2235), .B0(n2263), .Y(n2265));
  NOR4X1  g1652(.A(n2126), .B(n2110), .C(n2066), .D(n2178), .Y(n2266));
  XOR2X1  g1653(.A(n2233), .B(n2266), .Y(n2267));
  INVX1   g1654(.A(REG3_REG_27__SCAN_IN), .Y(n2268));
  NOR4X1  g1655(.A(n2215), .B(n2112), .C(n2162), .D(n2113), .Y(n2269));
  XOR2X1  g1656(.A(n2269), .B(n2268), .Y(n2270));
  INVX1   g1657(.A(n2270), .Y(n2271));
  AOI22X1 g1658(.A0(n917), .A1(REG0_REG_27__SCAN_IN), .B0(REG2_REG_27__SCAN_IN), .B1(n952), .Y(n2272));
  INVX1   g1659(.A(n2272), .Y(n2273));
  AOI21X1 g1660(.A0(n954), .A1(REG1_REG_27__SCAN_IN), .B0(n2273), .Y(n2274));
  INVX1   g1661(.A(n2274), .Y(n2275));
  AOI21X1 g1662(.A0(n2271), .A1(n955), .B0(n2275), .Y(n2276));
  OAI22X1 g1663(.A0(n2233), .A1(n963), .B0(n1051), .B1(n2276), .Y(n2277));
  AOI21X1 g1664(.A0(n2267), .A1(n960), .B0(n2277), .Y(n2278));
  OAI21X1 g1665(.A0(n2265), .A1(n950), .B0(n2278), .Y(n2279));
  NOR2X1  g1666(.A(n2279), .B(n2257), .Y(n2280));
  NAND2X1 g1667(.A(n896), .B(REG0_REG_26__SCAN_IN), .Y(n2281));
  OAI21X1 g1668(.A0(n2280), .A1(n896), .B0(n2281), .Y(U3512));
  INVX1   g1669(.A(n2221), .Y(n2283));
  NOR2X1  g1670(.A(n2229), .B(n2283), .Y(n2284));
  INVX1   g1671(.A(n2284), .Y(n2285));
  INVX1   g1672(.A(DATAI_27_), .Y(n2286));
  NOR2X1  g1673(.A(n902), .B(n2286), .Y(n2287));
  XOR2X1  g1674(.A(n2287), .B(n2276), .Y(n2288));
  XOR2X1  g1675(.A(n2288), .B(n2285), .Y(n2289));
  INVX1   g1676(.A(n2289), .Y(n2290));
  NOR2X1  g1677(.A(n2233), .B(n2221), .Y(n2291));
  NOR2X1  g1678(.A(n2288), .B(n2291), .Y(n2292));
  AOI21X1 g1679(.A0(n2292), .A1(n2245), .B0(n2290), .Y(n2293));
  INVX1   g1680(.A(n2288), .Y(n2294));
  NOR3X1  g1681(.A(n2294), .B(n2246), .C(n2291), .Y(n2295));
  NOR3X1  g1682(.A(n2295), .B(n2293), .C(n1086), .Y(n2296));
  INVX1   g1683(.A(n2292), .Y(n2297));
  NOR2X1  g1684(.A(n2246), .B(n2291), .Y(n2298));
  OAI22X1 g1685(.A0(n2297), .A1(n2246), .B0(n2289), .B1(n2298), .Y(n2299));
  NAND2X1 g1686(.A(n2140), .B(n2102), .Y(n2300));
  NOR3X1  g1687(.A(n2231), .B(n2182), .C(n2141), .Y(n2301));
  AOI21X1 g1688(.A0(n2229), .A1(n2221), .B0(n2258), .Y(n2302));
  OAI22X1 g1689(.A0(n2259), .A1(n2302), .B0(n2231), .B1(n2206), .Y(n2303));
  AOI21X1 g1690(.A0(n2301), .A1(n2300), .B0(n2303), .Y(n2304));
  XOR2X1  g1691(.A(n2304), .B(n2288), .Y(n2305));
  AOI22X1 g1692(.A0(n2221), .A1(n992), .B0(n945), .B1(n2305), .Y(n2306));
  OAI21X1 g1693(.A0(n946), .A1(n939), .B0(n2305), .Y(n2307));
  NAND2X1 g1694(.A(n2307), .B(n2306), .Y(n2308));
  AOI21X1 g1695(.A0(n2299), .A1(n943), .B0(n2308), .Y(n2309));
  NAND2X1 g1696(.A(n2299), .B(n936), .Y(n2310));
  AOI21X1 g1697(.A0(n2246), .A1(n2285), .B0(n2297), .Y(n2311));
  NOR3X1  g1698(.A(n2298), .B(n2294), .C(n2284), .Y(n2312));
  OAI21X1 g1699(.A0(n2312), .A1(n2311), .B0(n931), .Y(n2313));
  NAND3X1 g1700(.A(n2313), .B(n2310), .C(n2309), .Y(n2314));
  XOR2X1  g1701(.A(n2304), .B(n2294), .Y(n2320));
  NAND3X1 g1702(.A(n2233), .B(n2212), .C(n2186), .Y(n2321));
  XOR2X1  g1703(.A(n2321), .B(n2287), .Y(n2322));
  INVX1   g1704(.A(n2287), .Y(n2323));
  NAND2X1 g1705(.A(n2269), .B(REG3_REG_27__SCAN_IN), .Y(n2324));
  XOR2X1  g1706(.A(n2324), .B(REG3_REG_28__SCAN_IN), .Y(n2325));
  INVX1   g1707(.A(n2325), .Y(n2326));
  AOI22X1 g1708(.A0(n917), .A1(REG0_REG_28__SCAN_IN), .B0(REG2_REG_28__SCAN_IN), .B1(n952), .Y(n2327));
  INVX1   g1709(.A(n2327), .Y(n2328));
  AOI21X1 g1710(.A0(n954), .A1(REG1_REG_28__SCAN_IN), .B0(n2328), .Y(n2329));
  INVX1   g1711(.A(n2329), .Y(n2330));
  AOI21X1 g1712(.A0(n2326), .A1(n955), .B0(n2330), .Y(n2331));
  OAI22X1 g1713(.A0(n2323), .A1(n963), .B0(n1051), .B1(n2331), .Y(n2332));
  AOI21X1 g1714(.A0(n2322), .A1(n960), .B0(n2332), .Y(n2333));
  OAI21X1 g1715(.A0(n2320), .A1(n950), .B0(n2333), .Y(n2334));
  NOR3X1  g1716(.A(n2334), .B(n2314), .C(n2296), .Y(n2335));
  NAND2X1 g1717(.A(n896), .B(REG0_REG_27__SCAN_IN), .Y(n2336));
  OAI21X1 g1718(.A0(n2335), .A1(n896), .B0(n2336), .Y(U3513));
  INVX1   g1719(.A(DATAI_28_), .Y(n2338));
  NOR2X1  g1720(.A(n902), .B(n2338), .Y(n2339));
  XOR2X1  g1721(.A(n2339), .B(n2331), .Y(n2340));
  INVX1   g1722(.A(n2340), .Y(n2341));
  INVX1   g1723(.A(n2276), .Y(n2342));
  AOI21X1 g1724(.A0(n2276), .A1(n2285), .B0(n2287), .Y(n2343));
  AOI21X1 g1725(.A0(n2342), .A1(n2284), .B0(n2343), .Y(n2344));
  AOI21X1 g1726(.A0(n2287), .A1(n2276), .B0(n2291), .Y(n2345));
  NAND2X1 g1727(.A(n2345), .B(n2245), .Y(n2346));
  NAND2X1 g1728(.A(n2346), .B(n2344), .Y(n2347));
  XOR2X1  g1729(.A(n2347), .B(n2341), .Y(n2348));
  NOR2X1  g1730(.A(n2348), .B(n1086), .Y(n2349));
  NOR2X1  g1731(.A(n2287), .B(n2342), .Y(n2353));
  NOR4X1  g1732(.A(n2231), .B(n2182), .C(n2141), .D(n2353), .Y(n2354));
  NOR3X1  g1733(.A(n2353), .B(n2231), .C(n2206), .Y(n2355));
  NOR2X1  g1734(.A(n2323), .B(n2276), .Y(n2356));
  NOR3X1  g1735(.A(n2353), .B(n2302), .C(n2259), .Y(n2357));
  NOR3X1  g1736(.A(n2357), .B(n2356), .C(n2355), .Y(n2358));
  INVX1   g1737(.A(n2358), .Y(n2359));
  AOI21X1 g1738(.A0(n2354), .A1(n2300), .B0(n2359), .Y(n2360));
  XOR2X1  g1739(.A(n2360), .B(n2341), .Y(n2361));
  OAI22X1 g1740(.A0(n2276), .A1(n1117), .B0(n1116), .B1(n2361), .Y(n2362));
  AOI21X1 g1741(.A0(n1141), .A1(n1140), .B0(n2361), .Y(n2363));
  NOR2X1  g1742(.A(n2363), .B(n2362), .Y(n2364));
  OAI21X1 g1743(.A0(n2348), .A1(n942), .B0(n2364), .Y(n2365));
  INVX1   g1744(.A(n2348), .Y(n2366));
  OAI21X1 g1745(.A0(n936), .A1(n931), .B0(n2366), .Y(n2367));
  INVX1   g1746(.A(n2367), .Y(n2368));
  INVX1   g1747(.A(n2356), .Y(n2369));
  OAI21X1 g1748(.A0(n2353), .A1(n2304), .B0(n2369), .Y(n2370));
  NAND4X1 g1749(.A(n2233), .B(n2212), .C(n2186), .D(n2323), .Y(n2372));
  XOR2X1  g1750(.A(n2339), .B(n2372), .Y(n2373));
  INVX1   g1751(.A(n2339), .Y(n2374));
  NAND3X1 g1752(.A(n2269), .B(REG3_REG_28__SCAN_IN), .C(REG3_REG_27__SCAN_IN), .Y(n2375));
  INVX1   g1753(.A(n2375), .Y(n2376));
  AOI22X1 g1754(.A0(n952), .A1(REG2_REG_29__SCAN_IN), .B0(REG1_REG_29__SCAN_IN), .B1(n954), .Y(n2377));
  INVX1   g1755(.A(n2377), .Y(n2378));
  AOI21X1 g1756(.A0(n917), .A1(REG0_REG_29__SCAN_IN), .B0(n2378), .Y(n2379));
  INVX1   g1757(.A(n2379), .Y(n2380));
  AOI21X1 g1758(.A0(n2376), .A1(n955), .B0(n2380), .Y(n2381));
  OAI22X1 g1759(.A0(n2374), .A1(n963), .B0(n1051), .B1(n2381), .Y(n2382));
  AOI21X1 g1760(.A0(n2373), .A1(n960), .B0(n2382), .Y(n2383));
  OAI21X1 g1761(.A0(n2361), .A1(n950), .B0(n2383), .Y(n2384));
  NOR4X1  g1762(.A(n2368), .B(n2365), .C(n2349), .D(n2384), .Y(n2385));
  NAND2X1 g1763(.A(n896), .B(REG0_REG_28__SCAN_IN), .Y(n2386));
  OAI21X1 g1764(.A0(n2385), .A1(n896), .B0(n2386), .Y(U3514));
  INVX1   g1765(.A(DATAI_29_), .Y(n2388));
  NOR2X1  g1766(.A(n902), .B(n2388), .Y(n2389));
  XOR2X1  g1767(.A(n2389), .B(n2381), .Y(n2390));
  NAND2X1 g1768(.A(n2370), .B(n2339), .Y(n2392));
  INVX1   g1769(.A(n2331), .Y(n2393));
  OAI21X1 g1770(.A0(n2370), .A1(n2339), .B0(n2393), .Y(n2394));
  NAND2X1 g1771(.A(n2394), .B(n2392), .Y(n2395));
  XOR2X1  g1772(.A(n2395), .B(n3804), .Y(n2396));
  NOR2X1  g1773(.A(n2360), .B(n2374), .Y(n2397));
  AOI21X1 g1774(.A0(n2360), .A1(n2374), .B0(n2331), .Y(n2398));
  NOR2X1  g1775(.A(n2398), .B(n2397), .Y(n2399));
  XOR2X1  g1776(.A(n2399), .B(n3804), .Y(n2400));
  NOR2X1  g1777(.A(n886), .B(n873), .Y(n2401));
  INVX1   g1778(.A(n2401), .Y(n2402));
  AOI21X1 g1779(.A0(n991), .A1(n773), .B0(n902), .Y(n2403));
  AOI22X1 g1780(.A0(n917), .A1(REG0_REG_30__SCAN_IN), .B0(REG2_REG_30__SCAN_IN), .B1(n952), .Y(n2404));
  INVX1   g1781(.A(n2404), .Y(n2405));
  AOI21X1 g1782(.A0(n954), .A1(REG1_REG_30__SCAN_IN), .B0(n2405), .Y(n2406));
  NOR3X1  g1783(.A(n2406), .B(n2403), .C(n2402), .Y(n2407));
  AOI21X1 g1784(.A0(n2393), .A1(n992), .B0(n2407), .Y(n2408));
  OAI21X1 g1785(.A0(n2400), .A1(n1141), .B0(n2408), .Y(n2409));
  AOI21X1 g1786(.A0(n1116), .A1(n1140), .B0(n2400), .Y(n2410));
  NOR2X1  g1787(.A(n2410), .B(n2409), .Y(n2411));
  AOI21X1 g1788(.A0(n2339), .A1(n2331), .B0(n2390), .Y(n2412));
  NAND2X1 g1789(.A(n2412), .B(n2347), .Y(n2413));
  NOR2X1  g1790(.A(n2339), .B(n2331), .Y(n2414));
  NOR3X1  g1791(.A(n3804), .B(n2374), .C(n2393), .Y(n2416));
  NOR3X1  g1792(.A(n2390), .B(n2339), .C(n2331), .Y(n2417));
  INVX1   g1793(.A(n2389), .Y(n2420));
  NOR3X1  g1794(.A(n2339), .B(n2321), .C(n2287), .Y(n2421));
  XOR2X1  g1795(.A(n2421), .B(n2389), .Y(n2422));
  OAI22X1 g1796(.A0(n2420), .A1(n963), .B0(n961), .B1(n2422), .Y(n2423));
  AOI21X1 g1797(.A0(n2430), .A1(n931), .B0(n2423), .Y(n2424));
  NOR2X1  g1798(.A(n2417), .B(n2416), .Y(n2425));
  OAI21X1 g1799(.A0(n2276), .A1(n2285), .B0(n2390), .Y(n2427));
  NOR3X1  g1800(.A(n2427), .B(n2343), .C(n2414), .Y(n2428));
  NAND2X1 g1801(.A(n2428), .B(n2346), .Y(n2429));
  NAND3X1 g1802(.A(n2429), .B(n2413), .C(n2425), .Y(n2430));
  NAND2X1 g1803(.A(n2430), .B(n941), .Y(n2431));
  OAI21X1 g1804(.A0(n943), .A1(n936), .B0(n2430), .Y(n2432));
  NAND4X1 g1805(.A(n2431), .B(n2424), .C(n2411), .D(n2432), .Y(n2433));
  AOI21X1 g1806(.A0(n2396), .A1(n949), .B0(n2433), .Y(n2434));
  NAND2X1 g1807(.A(n896), .B(REG0_REG_29__SCAN_IN), .Y(n2435));
  OAI21X1 g1808(.A0(n2434), .A1(n896), .B0(n2435), .Y(U3515));
  NOR4X1  g1809(.A(n2339), .B(n2321), .C(n2287), .D(n2389), .Y(n2437));
  INVX1   g1810(.A(DATAI_30_), .Y(n2438));
  NOR2X1  g1811(.A(n902), .B(n2438), .Y(n2439));
  INVX1   g1812(.A(n2439), .Y(n2440));
  XOR2X1  g1813(.A(n2440), .B(n2437), .Y(n2441));
  AOI22X1 g1814(.A0(n917), .A1(REG0_REG_31__SCAN_IN), .B0(REG2_REG_31__SCAN_IN), .B1(n952), .Y(n2442));
  INVX1   g1815(.A(n2442), .Y(n2443));
  AOI21X1 g1816(.A0(n954), .A1(REG1_REG_31__SCAN_IN), .B0(n2443), .Y(n2444));
  NOR3X1  g1817(.A(n2444), .B(n2403), .C(n2402), .Y(n2445));
  INVX1   g1818(.A(n2445), .Y(n2446));
  OAI21X1 g1819(.A0(n2440), .A1(n963), .B0(n2446), .Y(n2447));
  AOI21X1 g1820(.A0(n2441), .A1(n960), .B0(n2447), .Y(n2448));
  NAND2X1 g1821(.A(n896), .B(REG0_REG_30__SCAN_IN), .Y(n2449));
  OAI21X1 g1822(.A0(n2448), .A1(n896), .B0(n2449), .Y(U3516));
  INVX1   g1823(.A(DATAI_31_), .Y(n2451));
  NOR2X1  g1824(.A(n902), .B(n2451), .Y(n2452));
  NAND3X1 g1825(.A(n2440), .B(n2421), .C(n2420), .Y(n2453));
  XOR2X1  g1826(.A(n2453), .B(n2452), .Y(n2454));
  INVX1   g1827(.A(n2452), .Y(n2455));
  OAI21X1 g1828(.A0(n2455), .A1(n963), .B0(n2446), .Y(n2456));
  AOI21X1 g1829(.A0(n2454), .A1(n960), .B0(n2456), .Y(n2457));
  NAND2X1 g1830(.A(n896), .B(REG0_REG_31__SCAN_IN), .Y(n2458));
  OAI21X1 g1831(.A0(n2457), .A1(n896), .B0(n2458), .Y(U3517));
  NOR2X1  g1832(.A(n893), .B(n769), .Y(n2460));
  NAND4X1 g1833(.A(n891), .B(n870), .C(n868), .D(n2460), .Y(n2461));
  NAND2X1 g1834(.A(n2461), .B(REG1_REG_0__SCAN_IN), .Y(n2462));
  OAI21X1 g1835(.A0(n2461), .A1(n967), .B0(n2462), .Y(U3518));
  NAND2X1 g1836(.A(n2461), .B(REG1_REG_1__SCAN_IN), .Y(n2464));
  OAI21X1 g1837(.A0(n2461), .A1(n1005), .B0(n2464), .Y(U3519));
  NAND2X1 g1838(.A(n2461), .B(REG1_REG_2__SCAN_IN), .Y(n2466));
  OAI21X1 g1839(.A0(n2461), .A1(n1061), .B0(n2466), .Y(U3520));
  NAND2X1 g1840(.A(n2461), .B(REG1_REG_3__SCAN_IN), .Y(n2468));
  OAI21X1 g1841(.A0(n2461), .A1(n1113), .B0(n2468), .Y(U3521));
  NAND2X1 g1842(.A(n2461), .B(REG1_REG_4__SCAN_IN), .Y(n2470));
  OAI21X1 g1843(.A0(n2461), .A1(n1171), .B0(n2470), .Y(U3522));
  NAND2X1 g1844(.A(n2461), .B(REG1_REG_5__SCAN_IN), .Y(n2472));
  OAI21X1 g1845(.A0(n2461), .A1(n1221), .B0(n2472), .Y(U3523));
  NAND2X1 g1846(.A(n2461), .B(REG1_REG_6__SCAN_IN), .Y(n2474));
  OAI21X1 g1847(.A0(n2461), .A1(n1277), .B0(n2474), .Y(U3524));
  NAND2X1 g1848(.A(n2461), .B(REG1_REG_7__SCAN_IN), .Y(n2476));
  OAI21X1 g1849(.A0(n2461), .A1(n1343), .B0(n2476), .Y(U3525));
  NAND2X1 g1850(.A(n2461), .B(REG1_REG_8__SCAN_IN), .Y(n2478));
  OAI21X1 g1851(.A0(n2461), .A1(n1387), .B0(n2478), .Y(U3526));
  NAND2X1 g1852(.A(n2461), .B(REG1_REG_9__SCAN_IN), .Y(n2480));
  OAI21X1 g1853(.A0(n2461), .A1(n1438), .B0(n2480), .Y(U3527));
  NAND2X1 g1854(.A(n2461), .B(REG1_REG_10__SCAN_IN), .Y(n2482));
  OAI21X1 g1855(.A0(n2461), .A1(n1494), .B0(n2482), .Y(U3528));
  NAND2X1 g1856(.A(n2461), .B(REG1_REG_11__SCAN_IN), .Y(n2484));
  OAI21X1 g1857(.A0(n2461), .A1(n1551), .B0(n2484), .Y(U3529));
  NAND2X1 g1858(.A(n2461), .B(REG1_REG_12__SCAN_IN), .Y(n2486));
  OAI21X1 g1859(.A0(n2461), .A1(n1599), .B0(n2486), .Y(U3530));
  NAND2X1 g1860(.A(n2461), .B(REG1_REG_13__SCAN_IN), .Y(n2488));
  OAI21X1 g1861(.A0(n2461), .A1(n1649), .B0(n2488), .Y(U3531));
  NAND2X1 g1862(.A(n2461), .B(REG1_REG_14__SCAN_IN), .Y(n2490));
  OAI21X1 g1863(.A0(n2461), .A1(n1694), .B0(n2490), .Y(U3532));
  NAND2X1 g1864(.A(n2461), .B(REG1_REG_15__SCAN_IN), .Y(n2492));
  OAI21X1 g1865(.A0(n2461), .A1(n1741), .B0(n2492), .Y(U3533));
  NAND2X1 g1866(.A(n2461), .B(REG1_REG_16__SCAN_IN), .Y(n2494));
  OAI21X1 g1867(.A0(n2461), .A1(n1794), .B0(n2494), .Y(U3534));
  NAND2X1 g1868(.A(n2461), .B(REG1_REG_17__SCAN_IN), .Y(n2496));
  OAI21X1 g1869(.A0(n2461), .A1(n1842), .B0(n2496), .Y(U3535));
  NAND2X1 g1870(.A(n2461), .B(REG1_REG_18__SCAN_IN), .Y(n2498));
  OAI21X1 g1871(.A0(n2461), .A1(n1889), .B0(n2498), .Y(U3536));
  NAND2X1 g1872(.A(n2461), .B(REG1_REG_19__SCAN_IN), .Y(n2500));
  OAI21X1 g1873(.A0(n2461), .A1(n1930), .B0(n2500), .Y(U3537));
  NAND2X1 g1874(.A(n2461), .B(REG1_REG_20__SCAN_IN), .Y(n2502));
  OAI21X1 g1875(.A0(n2461), .A1(n1969), .B0(n2502), .Y(U3538));
  NAND2X1 g1876(.A(n2461), .B(REG1_REG_21__SCAN_IN), .Y(n2504));
  OAI21X1 g1877(.A0(n2461), .A1(n2013), .B0(n2504), .Y(U3539));
  NAND2X1 g1878(.A(n2461), .B(REG1_REG_22__SCAN_IN), .Y(n2506));
  OAI21X1 g1879(.A0(n2461), .A1(n2060), .B0(n2506), .Y(U3540));
  NAND2X1 g1880(.A(n2461), .B(REG1_REG_23__SCAN_IN), .Y(n2508));
  OAI21X1 g1881(.A0(n2461), .A1(n2122), .B0(n2508), .Y(U3541));
  NAND2X1 g1882(.A(n2461), .B(REG1_REG_24__SCAN_IN), .Y(n2510));
  OAI21X1 g1883(.A0(n2461), .A1(n2174), .B0(n2510), .Y(U3542));
  NAND2X1 g1884(.A(n2461), .B(REG1_REG_25__SCAN_IN), .Y(n2512));
  OAI21X1 g1885(.A0(n2461), .A1(n2224), .B0(n2512), .Y(U3543));
  NAND2X1 g1886(.A(n2461), .B(REG1_REG_26__SCAN_IN), .Y(n2514));
  OAI21X1 g1887(.A0(n2461), .A1(n2280), .B0(n2514), .Y(U3544));
  NAND2X1 g1888(.A(n2461), .B(REG1_REG_27__SCAN_IN), .Y(n2516));
  OAI21X1 g1889(.A0(n2461), .A1(n2335), .B0(n2516), .Y(U3545));
  NAND2X1 g1890(.A(n2461), .B(REG1_REG_28__SCAN_IN), .Y(n2518));
  OAI21X1 g1891(.A0(n2461), .A1(n2385), .B0(n2518), .Y(U3546));
  NAND2X1 g1892(.A(n2461), .B(REG1_REG_29__SCAN_IN), .Y(n2520));
  OAI21X1 g1893(.A0(n2461), .A1(n2434), .B0(n2520), .Y(U3547));
  NAND2X1 g1894(.A(n2461), .B(REG1_REG_30__SCAN_IN), .Y(n2522));
  OAI21X1 g1895(.A0(n2461), .A1(n2448), .B0(n2522), .Y(U3548));
  NAND2X1 g1896(.A(n2461), .B(REG1_REG_31__SCAN_IN), .Y(n2524));
  OAI21X1 g1897(.A0(n2461), .A1(n2457), .B0(n2524), .Y(U3549));
  NOR4X1  g1898(.A(n889), .B(n876), .C(n884), .D(n881), .Y(n2526));
  INVX1   g1899(.A(n868), .Y(n2527));
  AOI21X1 g1900(.A0(n881), .A1(n878), .B0(n2402), .Y(n2528));
  NOR4X1  g1901(.A(n894), .B(n870), .C(n2527), .D(n2528), .Y(n2529));
  OAI21X1 g1902(.A0(n2529), .A1(n2526), .B0(n768), .Y(n2530));
  NOR2X1  g1903(.A(n2530), .B(n1051), .Y(n2531));
  NAND2X1 g1904(.A(n2531), .B(n957), .Y(n2532));
  INVX1   g1905(.A(n2530), .Y(n2533));
  NOR2X1  g1906(.A(n2533), .B(n910), .Y(n2534));
  AOI21X1 g1907(.A0(n2533), .A1(n948), .B0(n2534), .Y(n2535));
  NOR2X1  g1908(.A(n2530), .B(n963), .Y(n2536));
  NOR4X1  g1909(.A(n881), .B(n889), .C(n873), .D(n2530), .Y(n2537));
  AOI22X1 g1910(.A0(n2536), .A1(n909), .B0(n3791), .B1(n2537), .Y(n2538));
  NOR3X1  g1911(.A(n2530), .B(n961), .C(n938), .Y(n2539));
  INVX1   g1912(.A(n2526), .Y(n2540));
  NOR4X1  g1913(.A(n767), .B(n758), .C(U3149), .D(n2540), .Y(n2541));
  AOI22X1 g1914(.A0(n2539), .A1(n909), .B0(REG3_REG_0__SCAN_IN), .B1(n2541), .Y(n2542));
  NAND4X1 g1915(.A(n2538), .B(n2535), .C(n2532), .D(n2542), .Y(U3290));
  NAND2X1 g1916(.A(n2531), .B(n1002), .Y(n2544));
  NOR2X1  g1917(.A(n2533), .B(n1014), .Y(n2545));
  AOI21X1 g1918(.A0(n2533), .A1(n995), .B0(n2545), .Y(n2546));
  AOI22X1 g1919(.A0(n2536), .A1(n974), .B0(n979), .B1(n2537), .Y(n2547));
  NOR4X1  g1920(.A(n999), .B(n961), .C(n938), .D(n2530), .Y(n2548));
  AOI21X1 g1921(.A0(n2541), .A1(REG3_REG_1__SCAN_IN), .B0(n2548), .Y(n2549));
  NAND4X1 g1922(.A(n2547), .B(n2546), .C(n2544), .D(n2549), .Y(U3289));
  AOI22X1 g1923(.A0(n2537), .A1(n1037), .B0(REG3_REG_2__SCAN_IN), .B1(n2541), .Y(n2551));
  AOI22X1 g1924(.A0(n2536), .A1(n1012), .B0(n1050), .B1(n2539), .Y(n2552));
  NAND2X1 g1925(.A(n2533), .B(n1047), .Y(n2553));
  AOI22X1 g1926(.A0(n2530), .A1(REG2_REG_2__SCAN_IN), .B0(n1079), .B1(n2531), .Y(n2554));
  NAND4X1 g1927(.A(n2553), .B(n2552), .C(n2551), .D(n2554), .Y(U3288));
  NAND2X1 g1928(.A(n2533), .B(n1100), .Y(n2556));
  AOI22X1 g1929(.A0(n2530), .A1(REG2_REG_3__SCAN_IN), .B0(n1122), .B1(n2531), .Y(n2557));
  AOI22X1 g1930(.A0(n2537), .A1(n1083), .B0(n1077), .B1(n2541), .Y(n2558));
  AOI22X1 g1931(.A0(n2536), .A1(n1073), .B0(n1102), .B1(n2539), .Y(n2559));
  NAND4X1 g1932(.A(n2558), .B(n2557), .C(n2556), .D(n2559), .Y(U3287));
  NOR3X1  g1933(.A(n1154), .B(n1142), .C(n1139), .Y(n2561));
  INVX1   g1934(.A(n2531), .Y(n2562));
  OAI22X1 g1935(.A0(n2533), .A1(n1103), .B0(n1167), .B1(n2562), .Y(n2563));
  INVX1   g1936(.A(n2537), .Y(n2564));
  INVX1   g1937(.A(n2541), .Y(n2565));
  OAI22X1 g1938(.A0(n2564), .A1(n1138), .B0(n1107), .B1(n2565), .Y(n2566));
  INVX1   g1939(.A(n2536), .Y(n2567));
  INVX1   g1940(.A(n2539), .Y(n2568));
  OAI22X1 g1941(.A0(n2567), .A1(n1127), .B0(n1158), .B1(n2568), .Y(n2569));
  NOR3X1  g1942(.A(n2569), .B(n2566), .C(n2563), .Y(n2570));
  OAI21X1 g1943(.A0(n2530), .A1(n2561), .B0(n2570), .Y(U3286));
  OAI22X1 g1944(.A0(n2533), .A1(n1160), .B0(n1285), .B1(n2562), .Y(n2572));
  NOR3X1  g1945(.A(n2564), .B(n1200), .C(n1192), .Y(n2573));
  NOR3X1  g1946(.A(n2540), .B(n1165), .C(n769), .Y(n2574));
  OAI22X1 g1947(.A0(n2567), .A1(n1188), .B0(n1212), .B1(n2568), .Y(n2575));
  NOR4X1  g1948(.A(n2574), .B(n2573), .C(n2572), .D(n2575), .Y(n2576));
  OAI21X1 g1949(.A0(n2530), .A1(n1209), .B0(n2576), .Y(U3285));
  OAI22X1 g1950(.A0(n2533), .A1(n1280), .B0(n1298), .B1(n2562), .Y(n2578));
  OAI22X1 g1951(.A0(n2564), .A1(n1255), .B0(n1215), .B1(n2565), .Y(n2579));
  OAI22X1 g1952(.A0(n2567), .A1(n1229), .B0(n1268), .B1(n2568), .Y(n2580));
  NOR3X1  g1953(.A(n2580), .B(n2579), .C(n2578), .Y(n2581));
  OAI21X1 g1954(.A0(n2530), .A1(n1263), .B0(n2581), .Y(U3284));
  NAND2X1 g1955(.A(n2533), .B(n1326), .Y(n2583));
  OAI22X1 g1956(.A0(n2533), .A1(n1293), .B0(n1339), .B1(n2562), .Y(n2584));
  OAI22X1 g1957(.A0(n2564), .A1(n1311), .B0(n1271), .B1(n2565), .Y(n2585));
  OAI22X1 g1958(.A0(n2567), .A1(n1300), .B0(n1329), .B1(n2568), .Y(n2586));
  NOR3X1  g1959(.A(n2586), .B(n2585), .C(n2584), .Y(n2587));
  NAND2X1 g1960(.A(n2587), .B(n2583), .Y(U3283));
  NOR3X1  g1961(.A(n1372), .B(n1363), .C(n1362), .Y(n2589));
  INVX1   g1962(.A(n1337), .Y(n2590));
  AOI22X1 g1963(.A0(n2539), .A1(n1374), .B0(n2590), .B1(n2541), .Y(n2591));
  OAI21X1 g1964(.A0(n2567), .A1(n1358), .B0(n2591), .Y(n2592));
  AOI22X1 g1965(.A0(n2530), .A1(REG2_REG_8__SCAN_IN), .B0(n1392), .B1(n2531), .Y(n2593));
  OAI21X1 g1966(.A0(n2564), .A1(n1361), .B0(n2593), .Y(n2594));
  NOR2X1  g1967(.A(n2594), .B(n2592), .Y(n2595));
  OAI21X1 g1968(.A0(n2530), .A1(n2589), .B0(n2595), .Y(U3282));
  NOR3X1  g1969(.A(n1423), .B(n1412), .C(n1410), .Y(n2597));
  AOI22X1 g1970(.A0(n2530), .A1(REG2_REG_9__SCAN_IN), .B0(n1444), .B1(n2531), .Y(n2598));
  NAND2X1 g1971(.A(n2536), .B(n1451), .Y(n2599));
  INVX1   g1972(.A(n1381), .Y(n2600));
  AOI22X1 g1973(.A0(n2539), .A1(n1425), .B0(n2600), .B1(n2541), .Y(n2601));
  NAND3X1 g1974(.A(n2601), .B(n2599), .C(n2598), .Y(n2602));
  AOI21X1 g1975(.A0(n2537), .A1(n1421), .B0(n2602), .Y(n2603));
  OAI21X1 g1976(.A0(n2530), .A1(n2597), .B0(n2603), .Y(U3281));
  AOI22X1 g1977(.A0(n2530), .A1(REG2_REG_10__SCAN_IN), .B0(n1502), .B1(n2531), .Y(n2605));
  NAND2X1 g1978(.A(n2536), .B(n1461), .Y(n2606));
  AOI22X1 g1979(.A0(n2539), .A1(n1480), .B0(n1442), .B1(n2541), .Y(n2607));
  NAND3X1 g1980(.A(n2607), .B(n2606), .C(n2605), .Y(n2608));
  AOI21X1 g1981(.A0(n2537), .A1(n1473), .B0(n2608), .Y(n2609));
  OAI21X1 g1982(.A0(n2530), .A1(n1476), .B0(n2609), .Y(U3280));
  NOR3X1  g1983(.A(n1537), .B(n1536), .C(n1535), .Y(n2611));
  AOI22X1 g1984(.A0(n2539), .A1(n1539), .B0(n1500), .B1(n2541), .Y(n2612));
  OAI21X1 g1985(.A0(n2567), .A1(n1507), .B0(n2612), .Y(n2613));
  AOI22X1 g1986(.A0(n2530), .A1(REG2_REG_11__SCAN_IN), .B0(n1567), .B1(n2531), .Y(n2614));
  OAI21X1 g1987(.A0(n2564), .A1(n1531), .B0(n2614), .Y(n2615));
  NOR2X1  g1988(.A(n2615), .B(n2613), .Y(n2616));
  OAI21X1 g1989(.A0(n2530), .A1(n2611), .B0(n2616), .Y(U3279));
  NOR3X1  g1990(.A(n1584), .B(n1580), .C(n1571), .Y(n2618));
  NOR2X1  g1991(.A(n2564), .B(n1570), .Y(n2619));
  AOI22X1 g1992(.A0(n2530), .A1(REG2_REG_12__SCAN_IN), .B0(n1594), .B1(n2531), .Y(n2620));
  NAND2X1 g1993(.A(n2536), .B(n1561), .Y(n2621));
  AOI22X1 g1994(.A0(n2539), .A1(n1586), .B0(n1565), .B1(n2541), .Y(n2622));
  NAND3X1 g1995(.A(n2622), .B(n2621), .C(n2620), .Y(n2623));
  NOR2X1  g1996(.A(n2623), .B(n2619), .Y(n2624));
  OAI21X1 g1997(.A0(n2530), .A1(n2618), .B0(n2624), .Y(U3278));
  NOR3X1  g1998(.A(n1633), .B(n1630), .C(n1617), .Y(n2626));
  AOI22X1 g1999(.A0(n2530), .A1(REG2_REG_13__SCAN_IN), .B0(n1620), .B1(n2536), .Y(n2627));
  NAND3X1 g2000(.A(n2526), .B(n1592), .C(n768), .Y(n2628));
  AOI22X1 g2001(.A0(n2531), .A1(n1710), .B0(n1635), .B1(n2539), .Y(n2629));
  NAND3X1 g2002(.A(n2629), .B(n2628), .C(n2627), .Y(n2630));
  AOI21X1 g2003(.A0(n2537), .A1(n1631), .B0(n2630), .Y(n2631));
  OAI21X1 g2004(.A0(n2530), .A1(n2626), .B0(n2631), .Y(U3277));
  NOR3X1  g2005(.A(n1678), .B(n1674), .C(n1666), .Y(n2633));
  NOR2X1  g2006(.A(n2564), .B(n1665), .Y(n2634));
  NAND2X1 g2007(.A(n2539), .B(n1682), .Y(n2635));
  AOI22X1 g2008(.A0(n2530), .A1(REG2_REG_14__SCAN_IN), .B0(n1689), .B1(n2531), .Y(n2636));
  INVX1   g2009(.A(n1643), .Y(n2637));
  AOI22X1 g2010(.A0(n2536), .A1(n1662), .B0(n2637), .B1(n2541), .Y(n2638));
  NAND3X1 g2011(.A(n2638), .B(n2636), .C(n2635), .Y(n2639));
  NOR2X1  g2012(.A(n2639), .B(n2634), .Y(n2640));
  OAI21X1 g2013(.A0(n2530), .A1(n2633), .B0(n2640), .Y(U3276));
  NAND2X1 g2014(.A(n2539), .B(n1727), .Y(n2642));
  AOI22X1 g2015(.A0(n2530), .A1(REG2_REG_15__SCAN_IN), .B0(n1744), .B1(n2536), .Y(n2643));
  INVX1   g2016(.A(n1686), .Y(n2644));
  AOI22X1 g2017(.A0(n2531), .A1(n1736), .B0(n2644), .B1(n2541), .Y(n2645));
  NAND3X1 g2018(.A(n2645), .B(n2643), .C(n2642), .Y(n2646));
  AOI21X1 g2019(.A0(n2537), .A1(n1716), .B0(n2646), .Y(n2647));
  OAI21X1 g2020(.A0(n2530), .A1(n1722), .B0(n2647), .Y(U3275));
  NAND2X1 g2021(.A(n2539), .B(n1782), .Y(n2649));
  AOI22X1 g2022(.A0(n2530), .A1(REG2_REG_16__SCAN_IN), .B0(n1769), .B1(n2536), .Y(n2650));
  INVX1   g2023(.A(n1733), .Y(n2651));
  AOI22X1 g2024(.A0(n2531), .A1(n1789), .B0(n2651), .B1(n2541), .Y(n2652));
  NAND3X1 g2025(.A(n2652), .B(n2650), .C(n2649), .Y(n2653));
  AOI21X1 g2026(.A0(n2537), .A1(n1773), .B0(n2653), .Y(n2654));
  OAI21X1 g2027(.A0(n2530), .A1(n1779), .B0(n2654), .Y(U3274));
  NAND2X1 g2028(.A(n2533), .B(n1827), .Y(n2656));
  NAND2X1 g2029(.A(n2539), .B(n1830), .Y(n2657));
  AOI22X1 g2030(.A0(n2530), .A1(REG2_REG_17__SCAN_IN), .B0(n1828), .B1(n2536), .Y(n2658));
  INVX1   g2031(.A(n1786), .Y(n2659));
  AOI22X1 g2032(.A0(n2531), .A1(n1837), .B0(n2659), .B1(n2541), .Y(n2660));
  NAND3X1 g2033(.A(n2660), .B(n2658), .C(n2657), .Y(n2661));
  AOI21X1 g2034(.A0(n2537), .A1(n1813), .B0(n2661), .Y(n2662));
  NAND2X1 g2035(.A(n2662), .B(n2656), .Y(U3273));
  NOR3X1  g2036(.A(n1874), .B(n1870), .C(n1861), .Y(n2664));
  NOR2X1  g2037(.A(n2564), .B(n1860), .Y(n2665));
  NAND2X1 g2038(.A(n2539), .B(n1876), .Y(n2666));
  AOI22X1 g2039(.A0(n2530), .A1(REG2_REG_18__SCAN_IN), .B0(n1857), .B1(n2536), .Y(n2667));
  INVX1   g2040(.A(n1834), .Y(n2668));
  AOI22X1 g2041(.A0(n2531), .A1(n1884), .B0(n2668), .B1(n2541), .Y(n2669));
  NAND3X1 g2042(.A(n2669), .B(n2667), .C(n2666), .Y(n2670));
  NOR2X1  g2043(.A(n2670), .B(n2665), .Y(n2671));
  OAI21X1 g2044(.A0(n2530), .A1(n2664), .B0(n2671), .Y(U3272));
  NAND2X1 g2045(.A(n2533), .B(n1916), .Y(n2673));
  NAND2X1 g2046(.A(n2539), .B(n1919), .Y(n2674));
  AOI22X1 g2047(.A0(n2530), .A1(REG2_REG_19__SCAN_IN), .B0(n1900), .B1(n2536), .Y(n2675));
  AOI22X1 g2048(.A0(n2531), .A1(n1925), .B0(n1882), .B1(n2541), .Y(n2676));
  NAND3X1 g2049(.A(n2676), .B(n2675), .C(n2674), .Y(n2677));
  AOI21X1 g2050(.A0(n2537), .A1(n1904), .B0(n2677), .Y(n2678));
  NAND2X1 g2051(.A(n2678), .B(n2673), .Y(U3271));
  NAND2X1 g2052(.A(n2533), .B(n1955), .Y(n2680));
  NAND2X1 g2053(.A(n2539), .B(n1957), .Y(n2681));
  AOI22X1 g2054(.A0(n2530), .A1(REG2_REG_20__SCAN_IN), .B0(n1935), .B1(n2536), .Y(n2682));
  AOI22X1 g2055(.A0(n2531), .A1(n1964), .B0(n1921), .B1(n2541), .Y(n2683));
  NAND3X1 g2056(.A(n2683), .B(n2682), .C(n2681), .Y(n2684));
  AOI21X1 g2057(.A0(n2537), .A1(n1945), .B0(n2684), .Y(n2685));
  NAND2X1 g2058(.A(n2685), .B(n2680), .Y(U3270));
  NAND2X1 g2059(.A(n2533), .B(n2000), .Y(n2687));
  NOR2X1  g2060(.A(n2564), .B(n1985), .Y(n2688));
  NAND2X1 g2061(.A(n2539), .B(n2002), .Y(n2689));
  AOI22X1 g2062(.A0(n2530), .A1(REG2_REG_21__SCAN_IN), .B0(n1973), .B1(n2536), .Y(n2690));
  AOI22X1 g2063(.A0(n2531), .A1(n2076), .B0(n1960), .B1(n2541), .Y(n2691));
  NAND3X1 g2064(.A(n2691), .B(n2690), .C(n2689), .Y(n2692));
  NOR2X1  g2065(.A(n2692), .B(n2688), .Y(n2693));
  NAND2X1 g2066(.A(n2693), .B(n2687), .Y(U3269));
  NOR3X1  g2067(.A(n2045), .B(n2044), .C(n2023), .Y(n2695));
  NAND2X1 g2068(.A(n2539), .B(n2048), .Y(n2696));
  AOI22X1 g2069(.A0(n2530), .A1(REG2_REG_22__SCAN_IN), .B0(n2017), .B1(n2536), .Y(n2697));
  AOI22X1 g2070(.A0(n2531), .A1(n2071), .B0(n2005), .B1(n2541), .Y(n2698));
  NAND3X1 g2071(.A(n2698), .B(n2697), .C(n2696), .Y(n2699));
  AOI21X1 g2072(.A0(n2537), .A1(n2041), .B0(n2699), .Y(n2700));
  OAI21X1 g2073(.A0(n2530), .A1(n2695), .B0(n2700), .Y(U3268));
  NAND2X1 g2074(.A(n2533), .B(n2107), .Y(n2702));
  NOR2X1  g2075(.A(n2564), .B(n2103), .Y(n2703));
  NAND2X1 g2076(.A(n2539), .B(n2111), .Y(n2704));
  AOI22X1 g2077(.A0(n2530), .A1(REG2_REG_23__SCAN_IN), .B0(n2066), .B1(n2536), .Y(n2705));
  AOI22X1 g2078(.A0(n2531), .A1(n2181), .B0(n2052), .B1(n2541), .Y(n2706));
  NAND3X1 g2079(.A(n2706), .B(n2705), .C(n2704), .Y(n2707));
  NOR2X1  g2080(.A(n2707), .B(n2703), .Y(n2708));
  NAND2X1 g2081(.A(n2708), .B(n2702), .Y(U3267));
  NAND2X1 g2082(.A(n2533), .B(n2152), .Y(n2710));
  NOR2X1  g2083(.A(n2564), .B(n2145), .Y(n2711));
  NAND2X1 g2084(.A(n2539), .B(n2161), .Y(n2712));
  AOI22X1 g2085(.A0(n2530), .A1(REG2_REG_24__SCAN_IN), .B0(n2126), .B1(n2536), .Y(n2713));
  AOI22X1 g2086(.A0(n2531), .A1(n2230), .B0(n2114), .B1(n2541), .Y(n2714));
  NAND3X1 g2087(.A(n2714), .B(n2713), .C(n2712), .Y(n2715));
  NOR2X1  g2088(.A(n2715), .B(n2711), .Y(n2716));
  NAND2X1 g2089(.A(n2716), .B(n2710), .Y(U3266));
  NAND2X1 g2090(.A(n2533), .B(n2205), .Y(n2718));
  NOR2X1  g2091(.A(n2564), .B(n2189), .Y(n2719));
  NAND2X1 g2092(.A(n2539), .B(n2213), .Y(n2720));
  AOI22X1 g2093(.A0(n2530), .A1(REG2_REG_25__SCAN_IN), .B0(n2178), .B1(n2536), .Y(n2721));
  AOI22X1 g2094(.A0(n2531), .A1(n2221), .B0(n2165), .B1(n2541), .Y(n2722));
  NAND3X1 g2095(.A(n2722), .B(n2721), .C(n2720), .Y(n2723));
  NOR2X1  g2096(.A(n2723), .B(n2719), .Y(n2724));
  NAND2X1 g2097(.A(n2724), .B(n2718), .Y(U3265));
  NAND2X1 g2098(.A(n2533), .B(n2257), .Y(n2726));
  NOR2X1  g2099(.A(n2564), .B(n2265), .Y(n2727));
  NAND2X1 g2100(.A(n2539), .B(n2267), .Y(n2728));
  AOI22X1 g2101(.A0(n2530), .A1(REG2_REG_26__SCAN_IN), .B0(n2229), .B1(n2536), .Y(n2729));
  INVX1   g2102(.A(n2217), .Y(n2730));
  AOI22X1 g2103(.A0(n2531), .A1(n2342), .B0(n2730), .B1(n2541), .Y(n2731));
  NAND3X1 g2104(.A(n2731), .B(n2729), .C(n2728), .Y(n2732));
  NOR2X1  g2105(.A(n2732), .B(n2727), .Y(n2733));
  NAND2X1 g2106(.A(n2733), .B(n2726), .Y(U3264));
  OAI21X1 g2107(.A0(n2314), .A1(n2296), .B0(n2533), .Y(n2735));
  NOR2X1  g2108(.A(n2564), .B(n2320), .Y(n2736));
  NAND2X1 g2109(.A(n2539), .B(n2322), .Y(n2737));
  AOI22X1 g2110(.A0(n2530), .A1(REG2_REG_27__SCAN_IN), .B0(n2287), .B1(n2536), .Y(n2738));
  AOI22X1 g2111(.A0(n2531), .A1(n2393), .B0(n2271), .B1(n2541), .Y(n2739));
  NAND3X1 g2112(.A(n2739), .B(n2738), .C(n2737), .Y(n2740));
  NOR2X1  g2113(.A(n2740), .B(n2736), .Y(n2741));
  NAND2X1 g2114(.A(n2741), .B(n2735), .Y(U3263));
  NOR3X1  g2115(.A(n2368), .B(n2365), .C(n2349), .Y(n2743));
  NOR2X1  g2116(.A(n2564), .B(n2361), .Y(n2744));
  NAND2X1 g2117(.A(n2539), .B(n2373), .Y(n2745));
  AOI22X1 g2118(.A0(n2530), .A1(REG2_REG_28__SCAN_IN), .B0(n2339), .B1(n2536), .Y(n2746));
  INVX1   g2119(.A(n2381), .Y(n2747));
  AOI22X1 g2120(.A0(n2531), .A1(n2747), .B0(n2326), .B1(n2541), .Y(n2748));
  NAND3X1 g2121(.A(n2748), .B(n2746), .C(n2745), .Y(n2749));
  NOR2X1  g2122(.A(n2749), .B(n2744), .Y(n2750));
  OAI21X1 g2123(.A0(n2530), .A1(n2743), .B0(n2750), .Y(U3262));
  NAND2X1 g2124(.A(n2537), .B(n2396), .Y(n2752));
  AOI22X1 g2125(.A0(n2430), .A1(n931), .B0(n941), .B1(n2430), .Y(n2753));
  NAND3X1 g2126(.A(n2753), .B(n2432), .C(n2411), .Y(n2754));
  NAND2X1 g2127(.A(n2530), .B(REG2_REG_29__SCAN_IN), .Y(n2755));
  OAI21X1 g2128(.A0(n2565), .A1(n2375), .B0(n2755), .Y(n2756));
  AOI21X1 g2129(.A0(n2536), .A1(n2389), .B0(n2756), .Y(n2757));
  OAI21X1 g2130(.A0(n2568), .A1(n2422), .B0(n2757), .Y(n2758));
  AOI21X1 g2131(.A0(n2754), .A1(n2533), .B0(n2758), .Y(n2759));
  NAND2X1 g2132(.A(n2759), .B(n2752), .Y(U3354));
  NAND2X1 g2133(.A(n2539), .B(n2441), .Y(n2761));
  NAND2X1 g2134(.A(n2536), .B(n2439), .Y(n2762));
  NAND2X1 g2135(.A(n2533), .B(n2445), .Y(n2763));
  NAND2X1 g2136(.A(n2530), .B(REG2_REG_30__SCAN_IN), .Y(n2764));
  NAND4X1 g2137(.A(n2763), .B(n2762), .C(n2761), .D(n2764), .Y(U3261));
  NAND2X1 g2138(.A(n2539), .B(n2454), .Y(n2766));
  NAND2X1 g2139(.A(n2536), .B(n2452), .Y(n2767));
  NAND2X1 g2140(.A(n2530), .B(REG2_REG_31__SCAN_IN), .Y(n2768));
  NAND4X1 g2141(.A(n2767), .B(n2766), .C(n2763), .D(n2768), .Y(U3260));
  NOR2X1  g2142(.A(n1802), .B(n1784), .Y(n2770));
  NOR3X1  g2143(.A(n1801), .B(n1800), .C(REG1_REG_17__SCAN_IN), .Y(n2771));
  INVX1   g2144(.A(n2771), .Y(n2772));
  NOR2X1  g2145(.A(n1747), .B(n1729), .Y(n2773));
  INVX1   g2146(.A(n2773), .Y(n2774));
  NOR2X1  g2147(.A(n1748), .B(REG1_REG_16__SCAN_IN), .Y(n2775));
  INVX1   g2148(.A(n1603), .Y(n2776));
  INVX1   g2149(.A(n1559), .Y(n2777));
  NOR2X1  g2150(.A(n2777), .B(n1543), .Y(n2778));
  INVX1   g2151(.A(n1504), .Y(n2779));
  NOR2X1  g2152(.A(n2779), .B(n1484), .Y(n2780));
  INVX1   g2153(.A(n2780), .Y(n2781));
  INVX1   g2154(.A(n1394), .Y(n2782));
  NOR2X1  g2155(.A(n2782), .B(n1378), .Y(n2783));
  NOR2X1  g2156(.A(n1394), .B(REG1_REG_9__SCAN_IN), .Y(n2784));
  INVX1   g2157(.A(n2784), .Y(n2785));
  INVX1   g2158(.A(n1352), .Y(n2786));
  INVX1   g2159(.A(n1290), .Y(n2787));
  NOR2X1  g2160(.A(n2787), .B(n1296), .Y(n2788));
  INVX1   g2161(.A(n1226), .Y(n2789));
  NOR2X1  g2162(.A(n2789), .B(n1283), .Y(n2790));
  INVX1   g2163(.A(n2790), .Y(n2791));
  INVX1   g2164(.A(n1124), .Y(n2792));
  NOR2X1  g2165(.A(n2792), .B(n1106), .Y(n2793));
  NOR2X1  g2166(.A(n1124), .B(REG1_REG_4__SCAN_IN), .Y(n2794));
  INVX1   g2167(.A(n2794), .Y(n2795));
  INVX1   g2168(.A(n1010), .Y(n2796));
  NOR2X1  g2169(.A(n2796), .B(n1031), .Y(n2797));
  NAND2X1 g2170(.A(n2796), .B(n1031), .Y(n2798));
  OAI21X1 g2171(.A0(n905), .A1(n904), .B0(REG1_REG_0__SCAN_IN), .Y(n2799));
  NAND2X1 g2172(.A(n759), .B(IR_REG_0__SCAN_IN), .Y(n2800));
  AOI21X1 g2173(.A0(n2800), .A1(n903), .B0(n923), .Y(n2801));
  OAI21X1 g2174(.A0(n2801), .A1(REG1_REG_1__SCAN_IN), .B0(n972), .Y(n2802));
  OAI21X1 g2175(.A0(n2799), .A1(n1018), .B0(n2802), .Y(n2803));
  AOI21X1 g2176(.A0(n2803), .A1(n2798), .B0(n2797), .Y(n2804));
  NAND2X1 g2177(.A(n2804), .B(n1055), .Y(n2805));
  NAND2X1 g2178(.A(n2805), .B(n1071), .Y(n2806));
  OAI21X1 g2179(.A0(n2804), .A1(n1055), .B0(n2806), .Y(n2807));
  AOI21X1 g2180(.A0(n2807), .A1(n2795), .B0(n2793), .Y(n2808));
  NOR2X1  g2181(.A(n2808), .B(n1163), .Y(n2809));
  INVX1   g2182(.A(n1176), .Y(n2810));
  AOI21X1 g2183(.A0(n2808), .A1(n1163), .B0(n2810), .Y(n2811));
  OAI22X1 g2184(.A0(n2809), .A1(n2811), .B0(n1226), .B1(REG1_REG_6__SCAN_IN), .Y(n2812));
  AOI22X1 g2185(.A0(n2791), .A1(n2812), .B0(n2787), .B1(n1296), .Y(n2813));
  OAI21X1 g2186(.A0(n2813), .A1(n2788), .B0(REG1_REG_8__SCAN_IN), .Y(n2814));
  NOR3X1  g2187(.A(n2813), .B(n2788), .C(REG1_REG_8__SCAN_IN), .Y(n2815));
  OAI21X1 g2188(.A0(n2815), .A1(n2786), .B0(n2814), .Y(n2816));
  AOI21X1 g2189(.A0(n2816), .A1(n2785), .B0(n2783), .Y(n2817));
  NOR2X1  g2190(.A(n2817), .B(n1429), .Y(n2818));
  INVX1   g2191(.A(n1446), .Y(n2819));
  AOI21X1 g2192(.A0(n2817), .A1(n1429), .B0(n2819), .Y(n2820));
  OAI22X1 g2193(.A0(n2818), .A1(n2820), .B0(n1504), .B1(REG1_REG_11__SCAN_IN), .Y(n2821));
  AOI22X1 g2194(.A0(n2781), .A1(n2821), .B0(n2777), .B1(n1543), .Y(n2822));
  OAI21X1 g2195(.A0(n2822), .A1(n2778), .B0(REG1_REG_13__SCAN_IN), .Y(n2823));
  NOR3X1  g2196(.A(n2822), .B(n2778), .C(REG1_REG_13__SCAN_IN), .Y(n2824));
  OAI21X1 g2197(.A0(n2824), .A1(n2776), .B0(n2823), .Y(n2825));
  NAND2X1 g2198(.A(n2825), .B(REG1_REG_14__SCAN_IN), .Y(n2826));
  OAI21X1 g2199(.A0(n2825), .A1(REG1_REG_14__SCAN_IN), .B0(n1660), .Y(n2827));
  AOI21X1 g2200(.A0(n2827), .A1(n2826), .B0(n1684), .Y(n2828));
  NAND3X1 g2201(.A(n2827), .B(n2826), .C(n1684), .Y(n2829));
  AOI21X1 g2202(.A0(n2829), .A1(n1699), .B0(n2828), .Y(n2830));
  OAI21X1 g2203(.A0(n2830), .A1(n2775), .B0(n2774), .Y(n2831));
  AOI21X1 g2204(.A0(n2831), .A1(n2772), .B0(n2770), .Y(n2832));
  OAI21X1 g2205(.A0(n1850), .A1(n1832), .B0(n2832), .Y(n2833));
  NOR2X1  g2206(.A(n1851), .B(REG1_REG_18__SCAN_IN), .Y(n2834));
  XOR2X1  g2207(.A(n881), .B(REG1_REG_19__SCAN_IN), .Y(n2835));
  NOR2X1  g2208(.A(n2835), .B(n2834), .Y(n2836));
  NAND2X1 g2209(.A(n2836), .B(n2833), .Y(n2837));
  INVX1   g2210(.A(n2835), .Y(n2838));
  AOI21X1 g2211(.A0(n1851), .A1(REG1_REG_18__SCAN_IN), .B0(n2838), .Y(n2839));
  OAI21X1 g2212(.A0(n2834), .A1(n2832), .B0(n2839), .Y(n2840));
  NAND3X1 g2213(.A(n771), .B(n775), .C(n785), .Y(n2841));
  NOR2X1  g2214(.A(n2841), .B(n758), .Y(n2842));
  AOI21X1 g2215(.A0(n2402), .A1(n2841), .B0(n758), .Y(n2843));
  OAI21X1 g2216(.A0(n2843), .A1(n902), .B0(STATE_REG_SCAN_IN), .Y(U3148));
  NOR2X1  g2217(.A(U3148), .B(n2842), .Y(n2845));
  NOR2X1  g2218(.A(n2845), .B(n769), .Y(n2846));
  NOR4X1  g2219(.A(n889), .B(n876), .C(n884), .D(n938), .Y(n2847));
  NOR2X1  g2220(.A(n889), .B(n886), .Y(n2848));
  NAND2X1 g2221(.A(n2848), .B(n881), .Y(n2849));
  NAND3X1 g2222(.A(n963), .B(n2849), .C(n932), .Y(n2850));
  OAI21X1 g2223(.A0(n878), .A1(n886), .B0(n873), .Y(n2851));
  NOR4X1  g2224(.A(n2850), .B(n2847), .C(n2526), .D(n2851), .Y(n2852));
  NOR2X1  g2225(.A(n2852), .B(n899), .Y(n2853));
  NAND4X1 g2226(.A(n2846), .B(n2840), .C(n2837), .D(n2853), .Y(n2854));
  NOR4X1  g2227(.A(n899), .B(n757), .C(U3149), .D(n2845), .Y(n2855));
  NAND3X1 g2228(.A(n2855), .B(n2840), .C(n2837), .Y(n2856));
  INVX1   g2229(.A(n2846), .Y(n2857));
  INVX1   g2230(.A(REG2_REG_17__SCAN_IN), .Y(n2858));
  NOR2X1  g2231(.A(n1802), .B(n2858), .Y(n2859));
  INVX1   g2232(.A(n2859), .Y(n2860));
  NOR3X1  g2233(.A(n1801), .B(n1800), .C(REG2_REG_17__SCAN_IN), .Y(n2861));
  INVX1   g2234(.A(REG2_REG_16__SCAN_IN), .Y(n2862));
  NOR2X1  g2235(.A(n1747), .B(n2862), .Y(n2863));
  NOR2X1  g2236(.A(n1748), .B(REG2_REG_16__SCAN_IN), .Y(n2864));
  INVX1   g2237(.A(n2864), .Y(n2865));
  INVX1   g2238(.A(REG2_REG_15__SCAN_IN), .Y(n2866));
  INVX1   g2239(.A(n1699), .Y(n2867));
  NOR2X1  g2240(.A(n2867), .B(n2866), .Y(n2868));
  INVX1   g2241(.A(n2868), .Y(n2869));
  NOR2X1  g2242(.A(n1699), .B(REG2_REG_15__SCAN_IN), .Y(n2870));
  INVX1   g2243(.A(REG2_REG_14__SCAN_IN), .Y(n2871));
  INVX1   g2244(.A(n1660), .Y(n2872));
  NOR2X1  g2245(.A(n2872), .B(n2871), .Y(n2873));
  NOR2X1  g2246(.A(n1660), .B(REG2_REG_14__SCAN_IN), .Y(n2874));
  INVX1   g2247(.A(n2874), .Y(n2875));
  INVX1   g2248(.A(REG2_REG_13__SCAN_IN), .Y(n2876));
  NOR2X1  g2249(.A(n2776), .B(n2876), .Y(n2877));
  INVX1   g2250(.A(n2877), .Y(n2878));
  NOR2X1  g2251(.A(n1603), .B(REG2_REG_13__SCAN_IN), .Y(n2879));
  NOR2X1  g2252(.A(n2777), .B(n1540), .Y(n2880));
  NOR2X1  g2253(.A(n1559), .B(REG2_REG_12__SCAN_IN), .Y(n2881));
  INVX1   g2254(.A(n2881), .Y(n2882));
  NOR2X1  g2255(.A(n2779), .B(n1481), .Y(n2883));
  INVX1   g2256(.A(n2883), .Y(n2884));
  NOR2X1  g2257(.A(n1504), .B(REG2_REG_11__SCAN_IN), .Y(n2885));
  NOR2X1  g2258(.A(n2819), .B(n1426), .Y(n2886));
  NOR2X1  g2259(.A(n1446), .B(REG2_REG_10__SCAN_IN), .Y(n2887));
  INVX1   g2260(.A(n2887), .Y(n2888));
  NOR2X1  g2261(.A(n2782), .B(n1375), .Y(n2889));
  INVX1   g2262(.A(n2889), .Y(n2890));
  NOR2X1  g2263(.A(n1394), .B(REG2_REG_9__SCAN_IN), .Y(n2891));
  NOR2X1  g2264(.A(n2786), .B(n1330), .Y(n2892));
  NOR2X1  g2265(.A(n1352), .B(REG2_REG_8__SCAN_IN), .Y(n2893));
  INVX1   g2266(.A(n2893), .Y(n2894));
  NOR2X1  g2267(.A(n2787), .B(n1293), .Y(n2895));
  INVX1   g2268(.A(n2895), .Y(n2896));
  NOR2X1  g2269(.A(n1290), .B(REG2_REG_7__SCAN_IN), .Y(n2897));
  NOR2X1  g2270(.A(n2789), .B(n1280), .Y(n2898));
  NOR2X1  g2271(.A(n1226), .B(REG2_REG_6__SCAN_IN), .Y(n2899));
  INVX1   g2272(.A(n2899), .Y(n2900));
  INVX1   g2273(.A(n1071), .Y(n2901));
  NOR2X1  g2274(.A(n582), .B(n759), .Y(n2902));
  AOI21X1 g2275(.A0(n759), .A1(IR_REG_1__SCAN_IN), .B0(n2902), .Y(n2903));
  OAI21X1 g2276(.A0(n905), .A1(n904), .B0(REG2_REG_0__SCAN_IN), .Y(n2904));
  AOI21X1 g2277(.A0(n2800), .A1(n903), .B0(n910), .Y(n2905));
  OAI21X1 g2278(.A0(n2905), .A1(n972), .B0(REG2_REG_1__SCAN_IN), .Y(n2906));
  OAI21X1 g2279(.A0(n2904), .A1(n2903), .B0(n2906), .Y(n2907));
  OAI21X1 g2280(.A0(n1010), .A1(REG2_REG_2__SCAN_IN), .B0(n2907), .Y(n2908));
  OAI21X1 g2281(.A0(n2796), .A1(n1028), .B0(n2908), .Y(n2909));
  OAI21X1 g2282(.A0(n1071), .A1(REG2_REG_3__SCAN_IN), .B0(n2909), .Y(n2910));
  OAI21X1 g2283(.A0(n2901), .A1(n1052), .B0(n2910), .Y(n2911));
  OAI21X1 g2284(.A0(n1124), .A1(REG2_REG_4__SCAN_IN), .B0(n2911), .Y(n2912));
  OAI21X1 g2285(.A0(n2792), .A1(n1103), .B0(n2912), .Y(n2913));
  OAI21X1 g2286(.A0(n1176), .A1(REG2_REG_5__SCAN_IN), .B0(n2913), .Y(n2914));
  OAI21X1 g2287(.A0(n2810), .A1(n1160), .B0(n2914), .Y(n2915));
  AOI21X1 g2288(.A0(n2915), .A1(n2900), .B0(n2898), .Y(n2916));
  OAI21X1 g2289(.A0(n2916), .A1(n2897), .B0(n2896), .Y(n2917));
  AOI21X1 g2290(.A0(n2917), .A1(n2894), .B0(n2892), .Y(n2918));
  OAI21X1 g2291(.A0(n2918), .A1(n2891), .B0(n2890), .Y(n2919));
  AOI21X1 g2292(.A0(n2919), .A1(n2888), .B0(n2886), .Y(n2920));
  OAI21X1 g2293(.A0(n2920), .A1(n2885), .B0(n2884), .Y(n2921));
  AOI21X1 g2294(.A0(n2921), .A1(n2882), .B0(n2880), .Y(n2922));
  OAI21X1 g2295(.A0(n2922), .A1(n2879), .B0(n2878), .Y(n2923));
  AOI21X1 g2296(.A0(n2923), .A1(n2875), .B0(n2873), .Y(n2924));
  OAI21X1 g2297(.A0(n2924), .A1(n2870), .B0(n2869), .Y(n2925));
  AOI21X1 g2298(.A0(n2925), .A1(n2865), .B0(n2863), .Y(n2926));
  OAI21X1 g2299(.A0(n2926), .A1(n2861), .B0(n2860), .Y(n2927));
  AOI21X1 g2300(.A0(n1851), .A1(REG2_REG_18__SCAN_IN), .B0(n2927), .Y(n2928));
  NOR2X1  g2301(.A(n1851), .B(REG2_REG_18__SCAN_IN), .Y(n2929));
  XOR2X1  g2302(.A(n881), .B(REG2_REG_19__SCAN_IN), .Y(n2930));
  NOR3X1  g2303(.A(n2930), .B(n2929), .C(n2928), .Y(n2931));
  INVX1   g2304(.A(n2929), .Y(n2932));
  INVX1   g2305(.A(REG2_REG_18__SCAN_IN), .Y(n2933));
  OAI21X1 g2306(.A0(n1850), .A1(n2933), .B0(n2930), .Y(n2934));
  AOI21X1 g2307(.A0(n2932), .A1(n2927), .B0(n2934), .Y(n2935));
  OAI21X1 g2308(.A0(n901), .A1(n900), .B0(n899), .Y(n2936));
  NOR2X1  g2309(.A(n2936), .B(n2852), .Y(n2937));
  NOR4X1  g2310(.A(n2935), .B(n2931), .C(n2857), .D(n2936), .Y(n2939));
  NOR4X1  g2311(.A(n2845), .B(n757), .C(U3149), .D(n2936), .Y(n2940));
  INVX1   g2312(.A(n2940), .Y(n2941));
  NOR3X1  g2313(.A(n2941), .B(n2935), .C(n2931), .Y(n2942));
  INVX1   g2314(.A(n991), .Y(n2943));
  NOR4X1  g2315(.A(n2943), .B(n757), .C(U3149), .D(n2845), .Y(n2944));
  NAND2X1 g2316(.A(n2944), .B(n938), .Y(n2945));
  NAND3X1 g2317(.A(n991), .B(n2846), .C(n938), .Y(n2947));
  AOI22X1 g2318(.A0(ADDR_REG_19__SCAN_IN), .A1(n2845), .B0(REG3_REG_19__SCAN_IN), .B1(U3149), .Y(n2948));
  NAND3X1 g2319(.A(n2948), .B(n2947), .C(n2945), .Y(n2949));
  NOR3X1  g2320(.A(n2949), .B(n2942), .C(n2939), .Y(n2950));
  NAND3X1 g2321(.A(n2950), .B(n2856), .C(n2854), .Y(U3259));
  XOR2X1  g2322(.A(n1850), .B(REG1_REG_18__SCAN_IN), .Y(n2952));
  XOR2X1  g2323(.A(n2952), .B(n2832), .Y(n2953));
  NAND3X1 g2324(.A(n2953), .B(n2853), .C(n2846), .Y(n2954));
  NAND2X1 g2325(.A(n2953), .B(n2855), .Y(n2955));
  XOR2X1  g2326(.A(n1850), .B(n2933), .Y(n2956));
  XOR2X1  g2327(.A(n2956), .B(n2927), .Y(n2957));
  NAND3X1 g2328(.A(n2957), .B(n2937), .C(n2846), .Y(n2958));
  NAND2X1 g2329(.A(n2944), .B(n1851), .Y(n2959));
  NAND3X1 g2330(.A(n991), .B(n2846), .C(n1851), .Y(n2960));
  AOI22X1 g2331(.A0(REG3_REG_18__SCAN_IN), .A1(U3149), .B0(ADDR_REG_18__SCAN_IN), .B1(n2845), .Y(n2961));
  NAND3X1 g2332(.A(n2961), .B(n2960), .C(n2959), .Y(n2962));
  AOI21X1 g2333(.A0(n2957), .A1(n2940), .B0(n2962), .Y(n2963));
  NAND4X1 g2334(.A(n2958), .B(n2955), .C(n2954), .D(n2963), .Y(U3258));
  XOR2X1  g2335(.A(n1802), .B(n1784), .Y(n2965));
  XOR2X1  g2336(.A(n2965), .B(n2831), .Y(n2966));
  XOR2X1  g2337(.A(n1802), .B(n2858), .Y(n2968));
  XOR2X1  g2338(.A(n2968), .B(n2926), .Y(n2969));
  OAI22X1 g2339(.A0(n2943), .A1(n1802), .B0(n2936), .B1(n2969), .Y(n2970));
  AOI21X1 g2340(.A0(n2966), .A1(n2853), .B0(n2970), .Y(n2971));
  NAND2X1 g2341(.A(n2845), .B(ADDR_REG_17__SCAN_IN), .Y(n2972));
  NAND2X1 g2342(.A(REG3_REG_17__SCAN_IN), .B(U3149), .Y(n2973));
  NAND2X1 g2343(.A(n2973), .B(n2972), .Y(n2974));
  AOI21X1 g2344(.A0(n2944), .A1(n1803), .B0(n2974), .Y(n2975));
  OAI21X1 g2345(.A0(n2969), .A1(n2941), .B0(n2975), .Y(n2976));
  AOI21X1 g2346(.A0(n2966), .A1(n2855), .B0(n2976), .Y(n2977));
  OAI21X1 g2347(.A0(n2971), .A1(n2857), .B0(n2977), .Y(U3257));
  XOR2X1  g2348(.A(n1747), .B(REG1_REG_16__SCAN_IN), .Y(n2979));
  XOR2X1  g2349(.A(n2979), .B(n2830), .Y(n2980));
  XOR2X1  g2350(.A(n1747), .B(REG2_REG_16__SCAN_IN), .Y(n2981));
  XOR2X1  g2351(.A(n2981), .B(n2925), .Y(n2982));
  OAI22X1 g2352(.A0(n2943), .A1(n1747), .B0(n2936), .B1(n2982), .Y(n2983));
  AOI21X1 g2353(.A0(n2980), .A1(n2853), .B0(n2983), .Y(n2984));
  NAND2X1 g2354(.A(n2845), .B(ADDR_REG_16__SCAN_IN), .Y(n2985));
  OAI21X1 g2355(.A0(n1730), .A1(STATE_REG_SCAN_IN), .B0(n2985), .Y(n2986));
  AOI21X1 g2356(.A0(n2944), .A1(n1748), .B0(n2986), .Y(n2987));
  OAI21X1 g2357(.A0(n2982), .A1(n2941), .B0(n2987), .Y(n2988));
  AOI21X1 g2358(.A0(n2980), .A1(n2855), .B0(n2988), .Y(n2989));
  OAI21X1 g2359(.A0(n2984), .A1(n2857), .B0(n2989), .Y(U3256));
  NAND2X1 g2360(.A(n2827), .B(n2826), .Y(n2991));
  XOR2X1  g2361(.A(n2991), .B(n1684), .Y(n2992));
  XOR2X1  g2362(.A(n2992), .B(n2867), .Y(n2993));
  XOR2X1  g2363(.A(n1699), .B(REG2_REG_15__SCAN_IN), .Y(n2994));
  XOR2X1  g2364(.A(n2994), .B(n2924), .Y(n2995));
  OAI22X1 g2365(.A0(n2943), .A1(n2867), .B0(n2936), .B1(n2995), .Y(n2996));
  AOI21X1 g2366(.A0(n2993), .A1(n2853), .B0(n2996), .Y(n2997));
  NAND2X1 g2367(.A(n2845), .B(ADDR_REG_15__SCAN_IN), .Y(n2998));
  NAND2X1 g2368(.A(REG3_REG_15__SCAN_IN), .B(U3149), .Y(n2999));
  NAND2X1 g2369(.A(n2999), .B(n2998), .Y(n3000));
  AOI21X1 g2370(.A0(n2944), .A1(n1699), .B0(n3000), .Y(n3001));
  OAI21X1 g2371(.A0(n2995), .A1(n2941), .B0(n3001), .Y(n3002));
  AOI21X1 g2372(.A0(n2993), .A1(n2855), .B0(n3002), .Y(n3003));
  OAI21X1 g2373(.A0(n2997), .A1(n2857), .B0(n3003), .Y(U3255));
  XOR2X1  g2374(.A(n2825), .B(REG1_REG_14__SCAN_IN), .Y(n3005));
  XOR2X1  g2375(.A(n3005), .B(n1660), .Y(n3006));
  XOR2X1  g2376(.A(n1660), .B(n2871), .Y(n3007));
  XOR2X1  g2377(.A(n3007), .B(n2923), .Y(n3008));
  OAI22X1 g2378(.A0(n2943), .A1(n2872), .B0(n2936), .B1(n3008), .Y(n3009));
  AOI21X1 g2379(.A0(n3006), .A1(n2853), .B0(n3009), .Y(n3010));
  NAND2X1 g2380(.A(n2845), .B(ADDR_REG_14__SCAN_IN), .Y(n3011));
  OAI21X1 g2381(.A0(n1639), .A1(STATE_REG_SCAN_IN), .B0(n3011), .Y(n3012));
  AOI21X1 g2382(.A0(n2944), .A1(n1660), .B0(n3012), .Y(n3013));
  OAI21X1 g2383(.A0(n3008), .A1(n2941), .B0(n3013), .Y(n3014));
  AOI21X1 g2384(.A0(n3006), .A1(n2855), .B0(n3014), .Y(n3015));
  OAI21X1 g2385(.A0(n3010), .A1(n2857), .B0(n3015), .Y(U3254));
  NOR2X1  g2386(.A(n2822), .B(n2778), .Y(n3017));
  XOR2X1  g2387(.A(n3017), .B(REG1_REG_13__SCAN_IN), .Y(n3018));
  XOR2X1  g2388(.A(n3018), .B(n2776), .Y(n3019));
  XOR2X1  g2389(.A(n1603), .B(REG2_REG_13__SCAN_IN), .Y(n3020));
  XOR2X1  g2390(.A(n3020), .B(n2922), .Y(n3021));
  OAI22X1 g2391(.A0(n2943), .A1(n2776), .B0(n2936), .B1(n3021), .Y(n3022));
  AOI21X1 g2392(.A0(n3019), .A1(n2853), .B0(n3022), .Y(n3023));
  NAND2X1 g2393(.A(n2845), .B(ADDR_REG_13__SCAN_IN), .Y(n3024));
  OAI21X1 g2394(.A0(n1641), .A1(STATE_REG_SCAN_IN), .B0(n3024), .Y(n3025));
  AOI21X1 g2395(.A0(n2944), .A1(n1603), .B0(n3025), .Y(n3026));
  OAI21X1 g2396(.A0(n3021), .A1(n2941), .B0(n3026), .Y(n3027));
  AOI21X1 g2397(.A0(n3019), .A1(n2855), .B0(n3027), .Y(n3028));
  OAI21X1 g2398(.A0(n3023), .A1(n2857), .B0(n3028), .Y(U3253));
  NAND2X1 g2399(.A(n2821), .B(n2781), .Y(n3030));
  XOR2X1  g2400(.A(n1559), .B(REG1_REG_12__SCAN_IN), .Y(n3031));
  XOR2X1  g2401(.A(n3031), .B(n3030), .Y(n3032));
  XOR2X1  g2402(.A(n1559), .B(n1540), .Y(n3033));
  XOR2X1  g2403(.A(n3033), .B(n2921), .Y(n3034));
  OAI22X1 g2404(.A0(n2943), .A1(n2777), .B0(n2936), .B1(n3034), .Y(n3035));
  AOI21X1 g2405(.A0(n3032), .A1(n2853), .B0(n3035), .Y(n3036));
  NAND2X1 g2406(.A(n2845), .B(ADDR_REG_12__SCAN_IN), .Y(n3037));
  OAI21X1 g2407(.A0(n1640), .A1(STATE_REG_SCAN_IN), .B0(n3037), .Y(n3038));
  AOI21X1 g2408(.A0(n2944), .A1(n1559), .B0(n3038), .Y(n3039));
  OAI21X1 g2409(.A0(n3034), .A1(n2941), .B0(n3039), .Y(n3040));
  AOI21X1 g2410(.A0(n3032), .A1(n2855), .B0(n3040), .Y(n3041));
  OAI21X1 g2411(.A0(n3036), .A1(n2857), .B0(n3041), .Y(U3252));
  NOR2X1  g2412(.A(n2820), .B(n2818), .Y(n3043));
  XOR2X1  g2413(.A(n1504), .B(n1484), .Y(n3044));
  XOR2X1  g2414(.A(n3044), .B(n3043), .Y(n3045));
  XOR2X1  g2415(.A(n1504), .B(REG2_REG_11__SCAN_IN), .Y(n3046));
  XOR2X1  g2416(.A(n3046), .B(n2920), .Y(n3047));
  OAI22X1 g2417(.A0(n2943), .A1(n2779), .B0(n2936), .B1(n3047), .Y(n3048));
  AOI21X1 g2418(.A0(n3045), .A1(n2853), .B0(n3048), .Y(n3049));
  NAND2X1 g2419(.A(n2845), .B(ADDR_REG_11__SCAN_IN), .Y(n3050));
  OAI21X1 g2420(.A0(n1485), .A1(STATE_REG_SCAN_IN), .B0(n3050), .Y(n3051));
  AOI21X1 g2421(.A0(n2944), .A1(n1504), .B0(n3051), .Y(n3052));
  OAI21X1 g2422(.A0(n3047), .A1(n2941), .B0(n3052), .Y(n3053));
  AOI21X1 g2423(.A0(n3045), .A1(n2855), .B0(n3053), .Y(n3054));
  OAI21X1 g2424(.A0(n3049), .A1(n2857), .B0(n3054), .Y(U3251));
  XOR2X1  g2425(.A(n2817), .B(n1429), .Y(n3056));
  XOR2X1  g2426(.A(n3056), .B(n1446), .Y(n3057));
  XOR2X1  g2427(.A(n1446), .B(n1426), .Y(n3058));
  XOR2X1  g2428(.A(n3058), .B(n2919), .Y(n3059));
  OAI22X1 g2429(.A0(n2943), .A1(n2819), .B0(n2936), .B1(n3059), .Y(n3060));
  AOI21X1 g2430(.A0(n3057), .A1(n2853), .B0(n3060), .Y(n3061));
  NAND2X1 g2431(.A(n2845), .B(ADDR_REG_10__SCAN_IN), .Y(n3062));
  OAI21X1 g2432(.A0(n1430), .A1(STATE_REG_SCAN_IN), .B0(n3062), .Y(n3063));
  AOI21X1 g2433(.A0(n2944), .A1(n1446), .B0(n3063), .Y(n3064));
  OAI21X1 g2434(.A0(n3059), .A1(n2941), .B0(n3064), .Y(n3065));
  AOI21X1 g2435(.A0(n3057), .A1(n2855), .B0(n3065), .Y(n3066));
  OAI21X1 g2436(.A0(n3061), .A1(n2857), .B0(n3066), .Y(U3250));
  XOR2X1  g2437(.A(n1394), .B(REG1_REG_9__SCAN_IN), .Y(n3068));
  XOR2X1  g2438(.A(n3068), .B(n2816), .Y(n3069));
  XOR2X1  g2439(.A(n1394), .B(REG2_REG_9__SCAN_IN), .Y(n3070));
  XOR2X1  g2440(.A(n3070), .B(n2918), .Y(n3071));
  OAI22X1 g2441(.A0(n2943), .A1(n2782), .B0(n2936), .B1(n3071), .Y(n3072));
  AOI21X1 g2442(.A0(n3069), .A1(n2853), .B0(n3072), .Y(n3073));
  NAND2X1 g2443(.A(n2845), .B(ADDR_REG_9__SCAN_IN), .Y(n3074));
  OAI21X1 g2444(.A0(n1379), .A1(STATE_REG_SCAN_IN), .B0(n3074), .Y(n3075));
  AOI21X1 g2445(.A0(n2944), .A1(n1394), .B0(n3075), .Y(n3076));
  OAI21X1 g2446(.A0(n3071), .A1(n2941), .B0(n3076), .Y(n3077));
  AOI21X1 g2447(.A0(n3069), .A1(n2855), .B0(n3077), .Y(n3078));
  OAI21X1 g2448(.A0(n3073), .A1(n2857), .B0(n3078), .Y(U3249));
  NOR2X1  g2449(.A(n2813), .B(n2788), .Y(n3080));
  XOR2X1  g2450(.A(n3080), .B(n1333), .Y(n3081));
  XOR2X1  g2451(.A(n3081), .B(n1352), .Y(n3082));
  XOR2X1  g2452(.A(n1352), .B(n1330), .Y(n3083));
  XOR2X1  g2453(.A(n3083), .B(n2917), .Y(n3084));
  OAI22X1 g2454(.A0(n2943), .A1(n2786), .B0(n2936), .B1(n3084), .Y(n3085));
  AOI21X1 g2455(.A0(n3082), .A1(n2853), .B0(n3085), .Y(n3086));
  NAND2X1 g2456(.A(n2845), .B(ADDR_REG_8__SCAN_IN), .Y(n3087));
  OAI21X1 g2457(.A0(n1334), .A1(STATE_REG_SCAN_IN), .B0(n3087), .Y(n3088));
  AOI21X1 g2458(.A0(n2944), .A1(n1352), .B0(n3088), .Y(n3089));
  OAI21X1 g2459(.A0(n3084), .A1(n2941), .B0(n3089), .Y(n3090));
  AOI21X1 g2460(.A0(n3082), .A1(n2855), .B0(n3090), .Y(n3091));
  OAI21X1 g2461(.A0(n3086), .A1(n2857), .B0(n3091), .Y(U3248));
  INVX1   g2462(.A(n2812), .Y(n3093));
  NOR2X1  g2463(.A(n3093), .B(n2790), .Y(n3094));
  XOR2X1  g2464(.A(n1290), .B(n1296), .Y(n3095));
  XOR2X1  g2465(.A(n3095), .B(n3094), .Y(n3096));
  NAND2X1 g2466(.A(n3096), .B(n2853), .Y(n3097));
  XOR2X1  g2467(.A(n1290), .B(n1293), .Y(n3098));
  XOR2X1  g2468(.A(n3098), .B(n2916), .Y(n3099));
  AOI22X1 g2469(.A0(n991), .A1(n1290), .B0(n2937), .B1(n3099), .Y(n3100));
  NAND2X1 g2470(.A(n3100), .B(n3097), .Y(n3101));
  NAND2X1 g2471(.A(n3101), .B(n2846), .Y(n3102));
  NAND2X1 g2472(.A(n3099), .B(n2940), .Y(n3103));
  AOI22X1 g2473(.A0(ADDR_REG_7__SCAN_IN), .A1(n2845), .B0(REG3_REG_7__SCAN_IN), .B1(U3149), .Y(n3104));
  AOI22X1 g2474(.A0(n2944), .A1(n1290), .B0(n2855), .B1(n3096), .Y(n3105));
  NAND4X1 g2475(.A(n3104), .B(n3103), .C(n3102), .D(n3105), .Y(U3247));
  NOR2X1  g2476(.A(n2811), .B(n2809), .Y(n3107));
  XOR2X1  g2477(.A(n1226), .B(n1283), .Y(n3108));
  XOR2X1  g2478(.A(n3108), .B(n3107), .Y(n3109));
  XOR2X1  g2479(.A(n1226), .B(n1280), .Y(n3110));
  XOR2X1  g2480(.A(n3110), .B(n2915), .Y(n3111));
  INVX1   g2481(.A(n3111), .Y(n3112));
  AOI22X1 g2482(.A0(n3109), .A1(n2853), .B0(n2937), .B1(n3112), .Y(n3113));
  OAI21X1 g2483(.A0(n2943), .A1(n2789), .B0(n3113), .Y(n3114));
  NAND2X1 g2484(.A(n3114), .B(n2846), .Y(n3115));
  NAND2X1 g2485(.A(n3112), .B(n2940), .Y(n3116));
  AOI22X1 g2486(.A0(REG3_REG_6__SCAN_IN), .A1(U3149), .B0(ADDR_REG_6__SCAN_IN), .B1(n2845), .Y(n3117));
  AOI22X1 g2487(.A0(n2944), .A1(n1226), .B0(n2855), .B1(n3109), .Y(n3118));
  NAND4X1 g2488(.A(n3117), .B(n3116), .C(n3115), .D(n3118), .Y(U3246));
  NOR3X1  g2489(.A(n2852), .B(n2810), .C(n2943), .Y(n3120));
  XOR2X1  g2490(.A(n2808), .B(n1163), .Y(n3122));
  XOR2X1  g2491(.A(n3122), .B(n2810), .Y(n3123));
  XOR2X1  g2492(.A(n1176), .B(n1160), .Y(n3124));
  XOR2X1  g2493(.A(n3124), .B(n2913), .Y(n3125));
  OAI22X1 g2494(.A0(n3123), .A1(n899), .B0(n2936), .B1(n3125), .Y(n3126));
  NOR2X1  g2495(.A(n3126), .B(n3120), .Y(n3127));
  AOI22X1 g2496(.A0(ADDR_REG_5__SCAN_IN), .A1(n2845), .B0(REG3_REG_5__SCAN_IN), .B1(U3149), .Y(n3128));
  OAI21X1 g2497(.A0(n3125), .A1(n2941), .B0(n3128), .Y(n3129));
  INVX1   g2498(.A(n2855), .Y(n3130));
  INVX1   g2499(.A(n2944), .Y(n3131));
  OAI22X1 g2500(.A0(n3131), .A1(n2810), .B0(n3130), .B1(n3123), .Y(n3132));
  NOR2X1  g2501(.A(n3132), .B(n3129), .Y(n3133));
  OAI21X1 g2502(.A0(n3127), .A1(n2857), .B0(n3133), .Y(U3245));
  NOR3X1  g2503(.A(n2841), .B(n758), .C(U3149), .Y(U4043));
  INVX1   g2504(.A(U4043), .Y(n3136));
  NAND2X1 g2505(.A(n886), .B(n873), .Y(n3137));
  NOR2X1  g2506(.A(n881), .B(n884), .Y(n3138));
  AOI21X1 g2507(.A0(n889), .A1(n884), .B0(n3138), .Y(n3139));
  AOI21X1 g2508(.A0(n3139), .A1(n3137), .B0(n767), .Y(n3140));
  NAND2X1 g2509(.A(n938), .B(n873), .Y(n3141));
  NOR3X1  g2510(.A(n938), .B(n889), .C(n886), .Y(n3142));
  AOI21X1 g2511(.A0(n938), .A1(n884), .B0(n878), .Y(n3143));
  NOR3X1  g2512(.A(n3143), .B(n3142), .C(n936), .Y(n3144));
  AOI21X1 g2513(.A0(n3144), .A1(n3141), .B0(n767), .Y(n3145));
  NAND3X1 g2514(.A(n878), .B(n884), .C(n2841), .Y(n3146));
  OAI22X1 g2515(.A0(n959), .A1(n3146), .B0(n576), .B1(n2841), .Y(n3147));
  AOI21X1 g2516(.A0(n3145), .A1(n986), .B0(n3147), .Y(n3148));
  XOR2X1  g2517(.A(n3148), .B(n3140), .Y(n3149));
  NOR2X1  g2518(.A(n876), .B(n884), .Y(n3150));
  OAI21X1 g2519(.A0(n878), .A1(n873), .B0(n3141), .Y(n3151));
  OAI21X1 g2520(.A0(n3151), .A1(n3150), .B0(n2841), .Y(n3152));
  NAND4X1 g2521(.A(n942), .B(n1097), .C(n890), .D(n2849), .Y(n3153));
  AOI21X1 g2522(.A0(n3141), .A1(n3137), .B0(n767), .Y(n3154));
  AOI21X1 g2523(.A0(n3153), .A1(n2841), .B0(n3154), .Y(n3155));
  NOR3X1  g2524(.A(n889), .B(n873), .C(n767), .Y(n3156));
  AOI22X1 g2525(.A0(n986), .A1(n3156), .B0(n767), .B1(REG1_REG_0__SCAN_IN), .Y(n3157));
  OAI21X1 g2526(.A0(n3155), .A1(n959), .B0(n3157), .Y(n3158));
  XOR2X1  g2527(.A(n3158), .B(n3152), .Y(n3159));
  XOR2X1  g2528(.A(n3159), .B(n3149), .Y(n3160));
  NOR2X1  g2529(.A(n991), .B(n899), .Y(n3161));
  NAND3X1 g2530(.A(n2800), .B(n903), .C(REG2_REG_0__SCAN_IN), .Y(n3162));
  AOI21X1 g2531(.A0(n899), .A1(n910), .B0(n991), .Y(n3163));
  OAI22X1 g2532(.A0(n3162), .A1(n2936), .B0(n576), .B1(n3163), .Y(n3164));
  AOI21X1 g2533(.A0(n3161), .A1(n3160), .B0(n3164), .Y(n3165));
  XOR2X1  g2534(.A(n1124), .B(n1106), .Y(n3166));
  XOR2X1  g2535(.A(n3166), .B(n2807), .Y(n3167));
  XOR2X1  g2536(.A(n1124), .B(n1103), .Y(n3168));
  XOR2X1  g2537(.A(n3168), .B(n2911), .Y(n3169));
  OAI22X1 g2538(.A0(n3167), .A1(n899), .B0(n2936), .B1(n3169), .Y(n3170));
  AOI21X1 g2539(.A0(n991), .A1(n1124), .B0(n3170), .Y(n3171));
  NOR2X1  g2540(.A(n3171), .B(n2857), .Y(n3172));
  AOI22X1 g2541(.A0(ADDR_REG_4__SCAN_IN), .A1(n2845), .B0(REG3_REG_4__SCAN_IN), .B1(U3149), .Y(n3173));
  OAI21X1 g2542(.A0(n3169), .A1(n2941), .B0(n3173), .Y(n3174));
  OAI22X1 g2543(.A0(n3131), .A1(n2792), .B0(n3130), .B1(n3167), .Y(n3175));
  NOR3X1  g2544(.A(n3175), .B(n3174), .C(n3172), .Y(n3176));
  OAI21X1 g2545(.A0(n3165), .A1(n3136), .B0(n3176), .Y(U3244));
  XOR2X1  g2546(.A(n2804), .B(n1055), .Y(n3178));
  XOR2X1  g2547(.A(n3178), .B(n2901), .Y(n3179));
  INVX1   g2548(.A(n3179), .Y(n3180));
  XOR2X1  g2549(.A(n1071), .B(n1052), .Y(n3181));
  XOR2X1  g2550(.A(n3181), .B(n2909), .Y(n3182));
  INVX1   g2551(.A(n3182), .Y(n3183));
  AOI22X1 g2552(.A0(n3180), .A1(n2853), .B0(n2937), .B1(n3183), .Y(n3184));
  OAI21X1 g2553(.A0(n2943), .A1(n2901), .B0(n3184), .Y(n3185));
  NAND2X1 g2554(.A(n3185), .B(n2846), .Y(n3186));
  NAND2X1 g2555(.A(n3183), .B(n2940), .Y(n3187));
  AOI22X1 g2556(.A0(ADDR_REG_3__SCAN_IN), .A1(n2845), .B0(REG3_REG_3__SCAN_IN), .B1(U3149), .Y(n3188));
  AOI22X1 g2557(.A0(n2944), .A1(n1071), .B0(n2855), .B1(n3180), .Y(n3189));
  NAND4X1 g2558(.A(n3188), .B(n3187), .C(n3186), .D(n3189), .Y(U3243));
  XOR2X1  g2559(.A(n1010), .B(n1031), .Y(n3191));
  XOR2X1  g2560(.A(n3191), .B(n2803), .Y(n3192));
  XOR2X1  g2561(.A(n1010), .B(n1028), .Y(n3193));
  XOR2X1  g2562(.A(n3193), .B(n2907), .Y(n3194));
  OAI22X1 g2563(.A0(n3192), .A1(n899), .B0(n2936), .B1(n3194), .Y(n3195));
  AOI21X1 g2564(.A0(n991), .A1(n1010), .B0(n3195), .Y(n3196));
  NOR2X1  g2565(.A(n3196), .B(n2857), .Y(n3197));
  AOI22X1 g2566(.A0(REG3_REG_2__SCAN_IN), .A1(U3149), .B0(ADDR_REG_2__SCAN_IN), .B1(n2845), .Y(n3198));
  OAI21X1 g2567(.A0(n3194), .A1(n2941), .B0(n3198), .Y(n3199));
  OAI22X1 g2568(.A0(n3131), .A1(n2796), .B0(n3130), .B1(n3192), .Y(n3200));
  NOR3X1  g2569(.A(n3200), .B(n3199), .C(n3197), .Y(n3201));
  OAI21X1 g2570(.A0(n3165), .A1(n3136), .B0(n3201), .Y(U3242));
  XOR2X1  g2571(.A(n2799), .B(n972), .Y(n3203));
  NOR2X1  g2572(.A(n2799), .B(n1018), .Y(n3204));
  NOR3X1  g2573(.A(n2801), .B(n972), .C(n1018), .Y(n3205));
  AOI21X1 g2574(.A0(n3204), .A1(n972), .B0(n3205), .Y(n3206));
  OAI21X1 g2575(.A0(n3203), .A1(REG1_REG_1__SCAN_IN), .B0(n3206), .Y(n3207));
  XOR2X1  g2576(.A(n2905), .B(n1014), .Y(n3208));
  NOR3X1  g2577(.A(n2904), .B(n2903), .C(n1014), .Y(n3209));
  NOR3X1  g2578(.A(n2905), .B(n2903), .C(REG2_REG_1__SCAN_IN), .Y(n3210));
  NOR2X1  g2579(.A(n3210), .B(n3209), .Y(n3211));
  OAI21X1 g2580(.A0(n3208), .A1(n972), .B0(n3211), .Y(n3212));
  AOI22X1 g2581(.A0(n3207), .A1(n2853), .B0(n2937), .B1(n3212), .Y(n3213));
  OAI21X1 g2582(.A0(n2943), .A1(n2903), .B0(n3213), .Y(n3214));
  NAND2X1 g2583(.A(n3214), .B(n2846), .Y(n3215));
  NAND2X1 g2584(.A(n3212), .B(n2940), .Y(n3216));
  AOI22X1 g2585(.A0(ADDR_REG_1__SCAN_IN), .A1(n2845), .B0(REG3_REG_1__SCAN_IN), .B1(U3149), .Y(n3217));
  AOI22X1 g2586(.A0(n2944), .A1(n972), .B0(n2855), .B1(n3207), .Y(n3218));
  NAND4X1 g2587(.A(n3217), .B(n3216), .C(n3215), .D(n3218), .Y(U3241));
  XOR2X1  g2588(.A(n576), .B(REG1_REG_0__SCAN_IN), .Y(n3220));
  INVX1   g2589(.A(n3220), .Y(n3221));
  XOR2X1  g2590(.A(n576), .B(REG2_REG_0__SCAN_IN), .Y(n3222));
  INVX1   g2591(.A(n3222), .Y(n3223));
  AOI22X1 g2592(.A0(n3221), .A1(n2853), .B0(n2937), .B1(n3223), .Y(n3224));
  OAI21X1 g2593(.A0(n2943), .A1(n576), .B0(n3224), .Y(n3225));
  NAND2X1 g2594(.A(n3225), .B(n2846), .Y(n3226));
  NAND2X1 g2595(.A(n3223), .B(n2940), .Y(n3227));
  AOI22X1 g2596(.A0(ADDR_REG_0__SCAN_IN), .A1(n2845), .B0(REG3_REG_0__SCAN_IN), .B1(U3149), .Y(n3228));
  AOI22X1 g2597(.A0(n2944), .A1(n907), .B0(n2855), .B1(n3221), .Y(n3229));
  NAND4X1 g2598(.A(n3228), .B(n3227), .C(n3226), .D(n3229), .Y(U3240));
  NAND2X1 g2599(.A(n3136), .B(DATAO_REG_0__SCAN_IN), .Y(n3231));
  OAI21X1 g2600(.A0(n3136), .A1(n929), .B0(n3231), .Y(U3550));
  NAND2X1 g2601(.A(n3136), .B(DATAO_REG_1__SCAN_IN), .Y(n3233));
  OAI21X1 g2602(.A0(n3136), .A1(n1020), .B0(n3233), .Y(U3551));
  NAND2X1 g2603(.A(n3136), .B(DATAO_REG_2__SCAN_IN), .Y(n3235));
  OAI21X1 g2604(.A0(n3136), .A1(n1034), .B0(n3235), .Y(U3552));
  NAND2X1 g2605(.A(n3136), .B(DATAO_REG_3__SCAN_IN), .Y(n3237));
  OAI21X1 g2606(.A0(n3136), .A1(n1057), .B0(n3237), .Y(U3553));
  NAND2X1 g2607(.A(n3136), .B(DATAO_REG_4__SCAN_IN), .Y(n3239));
  OAI21X1 g2608(.A0(n3136), .A1(n1109), .B0(n3239), .Y(U3554));
  NAND2X1 g2609(.A(n3136), .B(DATAO_REG_5__SCAN_IN), .Y(n3241));
  OAI21X1 g2610(.A0(n3136), .A1(n1167), .B0(n3241), .Y(U3555));
  NAND2X1 g2611(.A(n3136), .B(DATAO_REG_6__SCAN_IN), .Y(n3243));
  OAI21X1 g2612(.A0(n3136), .A1(n1285), .B0(n3243), .Y(U3556));
  NAND2X1 g2613(.A(n3136), .B(DATAO_REG_7__SCAN_IN), .Y(n3245));
  OAI21X1 g2614(.A0(n3136), .A1(n1298), .B0(n3245), .Y(U3557));
  NAND2X1 g2615(.A(n3136), .B(DATAO_REG_8__SCAN_IN), .Y(n3247));
  OAI21X1 g2616(.A0(n3136), .A1(n1339), .B0(n3247), .Y(U3558));
  NAND2X1 g2617(.A(n3136), .B(DATAO_REG_9__SCAN_IN), .Y(n3249));
  OAI21X1 g2618(.A0(n3136), .A1(n1383), .B0(n3249), .Y(U3559));
  NAND2X1 g2619(.A(n3136), .B(DATAO_REG_10__SCAN_IN), .Y(n3251));
  OAI21X1 g2620(.A0(n3136), .A1(n1434), .B0(n3251), .Y(U3560));
  NAND2X1 g2621(.A(n3136), .B(DATAO_REG_11__SCAN_IN), .Y(n3253));
  OAI21X1 g2622(.A0(n3136), .A1(n1490), .B0(n3253), .Y(U3561));
  NAND2X1 g2623(.A(n3136), .B(DATAO_REG_12__SCAN_IN), .Y(n3255));
  OAI21X1 g2624(.A0(n3136), .A1(n1547), .B0(n3255), .Y(U3562));
  NAND2X1 g2625(.A(n3136), .B(DATAO_REG_13__SCAN_IN), .Y(n3257));
  OAI21X1 g2626(.A0(n3136), .A1(n1595), .B0(n3257), .Y(U3563));
  NAND2X1 g2627(.A(n3136), .B(DATAO_REG_14__SCAN_IN), .Y(n3259));
  OAI21X1 g2628(.A0(n3136), .A1(n1645), .B0(n3259), .Y(U3564));
  NAND2X1 g2629(.A(n3136), .B(DATAO_REG_15__SCAN_IN), .Y(n3261));
  OAI21X1 g2630(.A0(n3136), .A1(n1690), .B0(n3261), .Y(U3565));
  NAND2X1 g2631(.A(n3136), .B(DATAO_REG_16__SCAN_IN), .Y(n3263));
  OAI21X1 g2632(.A0(n3136), .A1(n1737), .B0(n3263), .Y(U3566));
  NAND2X1 g2633(.A(n3136), .B(DATAO_REG_17__SCAN_IN), .Y(n3265));
  OAI21X1 g2634(.A0(n3136), .A1(n1790), .B0(n3265), .Y(U3567));
  NAND2X1 g2635(.A(n3136), .B(DATAO_REG_18__SCAN_IN), .Y(n3267));
  OAI21X1 g2636(.A0(n3136), .A1(n1838), .B0(n3267), .Y(U3568));
  NAND2X1 g2637(.A(n3136), .B(DATAO_REG_19__SCAN_IN), .Y(n3269));
  OAI21X1 g2638(.A0(n3136), .A1(n1885), .B0(n3269), .Y(U3569));
  NAND2X1 g2639(.A(n3136), .B(DATAO_REG_20__SCAN_IN), .Y(n3271));
  OAI21X1 g2640(.A0(n3136), .A1(n1926), .B0(n3271), .Y(U3570));
  NAND2X1 g2641(.A(n3136), .B(DATAO_REG_21__SCAN_IN), .Y(n3273));
  OAI21X1 g2642(.A0(n3136), .A1(n1965), .B0(n3273), .Y(U3571));
  NAND2X1 g2643(.A(n3136), .B(DATAO_REG_22__SCAN_IN), .Y(n3275));
  OAI21X1 g2644(.A0(n3136), .A1(n2009), .B0(n3275), .Y(U3572));
  NAND2X1 g2645(.A(n3136), .B(DATAO_REG_23__SCAN_IN), .Y(n3277));
  OAI21X1 g2646(.A0(n3136), .A1(n2056), .B0(n3277), .Y(U3573));
  NAND2X1 g2647(.A(n3136), .B(DATAO_REG_24__SCAN_IN), .Y(n3279));
  OAI21X1 g2648(.A0(n3136), .A1(n2118), .B0(n3279), .Y(U3574));
  NAND2X1 g2649(.A(n3136), .B(DATAO_REG_25__SCAN_IN), .Y(n3281));
  OAI21X1 g2650(.A0(n3136), .A1(n2170), .B0(n3281), .Y(U3575));
  NAND2X1 g2651(.A(n3136), .B(DATAO_REG_26__SCAN_IN), .Y(n3283));
  OAI21X1 g2652(.A0(n3136), .A1(n2283), .B0(n3283), .Y(U3576));
  NAND2X1 g2653(.A(n3136), .B(DATAO_REG_27__SCAN_IN), .Y(n3285));
  OAI21X1 g2654(.A0(n3136), .A1(n2276), .B0(n3285), .Y(U3577));
  NAND2X1 g2655(.A(n3136), .B(DATAO_REG_28__SCAN_IN), .Y(n3287));
  OAI21X1 g2656(.A0(n3136), .A1(n2331), .B0(n3287), .Y(U3578));
  NAND2X1 g2657(.A(n3136), .B(DATAO_REG_29__SCAN_IN), .Y(n3289));
  OAI21X1 g2658(.A0(n3136), .A1(n2381), .B0(n3289), .Y(U3579));
  NAND2X1 g2659(.A(n3136), .B(DATAO_REG_30__SCAN_IN), .Y(n3291));
  OAI21X1 g2660(.A0(n3136), .A1(n2406), .B0(n3291), .Y(U3580));
  NAND2X1 g2661(.A(n3136), .B(DATAO_REG_31__SCAN_IN), .Y(n3293));
  OAI21X1 g2662(.A0(n3136), .A1(n2444), .B0(n3293), .Y(U3581));
  NOR2X1  g2663(.A(n2287), .B(n2276), .Y(n3295));
  NAND4X1 g2664(.A(n955), .B(REG3_REG_28__SCAN_IN), .C(REG3_REG_27__SCAN_IN), .D(n2269), .Y(n3296));
  AOI21X1 g2665(.A0(n2379), .A1(n3296), .B0(n2389), .Y(n3297));
  NOR2X1  g2666(.A(n2439), .B(n2406), .Y(n3298));
  INVX1   g2667(.A(n2444), .Y(n3299));
  NOR2X1  g2668(.A(n2455), .B(n3299), .Y(n3300));
  NOR4X1  g2669(.A(n3298), .B(n3297), .C(n3295), .D(n3300), .Y(n3301));
  INVX1   g2670(.A(n3301), .Y(n3302));
  NOR2X1  g2671(.A(n3302), .B(n2414), .Y(n3303));
  INVX1   g2672(.A(n3303), .Y(n3304));
  NAND3X1 g2673(.A(n2196), .B(n2072), .C(n2071), .Y(n3305));
  NOR2X1  g2674(.A(n2243), .B(n2193), .Y(n3306));
  NAND3X1 g2675(.A(n3306), .B(n3305), .C(n2285), .Y(n3307));
  INVX1   g2676(.A(n1865), .Y(n3308));
  OAI22X1 g2677(.A0(n3308), .A1(n1906), .B0(n1769), .B1(n1737), .Y(n3309));
  AOI22X1 g2678(.A0(n1884), .A1(n1897), .B0(n1854), .B1(n1837), .Y(n3310));
  INVX1   g2679(.A(n3310), .Y(n3311));
  NOR4X1  g2680(.A(n3309), .B(n1982), .C(n1989), .D(n3311), .Y(n3312));
  AOI21X1 g2681(.A0(n1702), .A1(n1689), .B0(n1706), .Y(n3313));
  AOI22X1 g2682(.A0(n1594), .A1(n1606), .B0(n1588), .B1(n1567), .Y(n3314));
  NAND3X1 g2683(.A(n3314), .B(n3313), .C(n3312), .Y(n3315));
  AOI22X1 g2684(.A0(n1392), .A1(n1397), .B0(n1358), .B1(n1340), .Y(n3316));
  NOR3X1  g2685(.A(n1609), .B(n1514), .C(n1490), .Y(n3318));
  NOR4X1  g2686(.A(n3829), .B(n1512), .C(n1308), .D(n3318), .Y(n3319));
  INVX1   g2687(.A(n3319), .Y(n3320));
  AOI21X1 g2688(.A0(n1229), .A1(n1218), .B0(n3320), .Y(n3321));
  AOI21X1 g2689(.A0(n938), .A1(n886), .B0(n884), .Y(n3322));
  INVX1   g2690(.A(n3322), .Y(n3323));
  AOI21X1 g2691(.A0(n3323), .A1(n909), .B0(n929), .Y(n3324));
  NOR3X1  g2692(.A(n1316), .B(n1178), .C(n1167), .Y(n3325));
  AOI22X1 g2693(.A0(n998), .A1(n957), .B0(n959), .B1(n3322), .Y(n3326));
  INVX1   g2694(.A(n3326), .Y(n3327));
  NOR3X1  g2695(.A(n3327), .B(n3325), .C(n3324), .Y(n3328));
  NOR3X1  g2696(.A(n1181), .B(n1093), .C(n1035), .Y(n3329));
  NAND4X1 g2697(.A(n3328), .B(n3321), .C(n2064), .D(n3329), .Y(n3330));
  NOR4X1  g2698(.A(n3315), .B(n3307), .C(n3304), .D(n3330), .Y(n3331));
  INVX1   g2699(.A(n3307), .Y(n3332));
  NOR3X1  g2700(.A(n2192), .B(n2073), .C(n2064), .Y(n3333));
  NOR2X1  g2701(.A(n3333), .B(n3315), .Y(n3334));
  NAND3X1 g2702(.A(n3334), .B(n3332), .C(n1513), .Y(n3335));
  NOR2X1  g2703(.A(n3335), .B(n3304), .Y(n3336));
  NOR4X1  g2704(.A(n3318), .B(n3315), .C(n1510), .D(n3333), .Y(n3337));
  NAND3X1 g2705(.A(n3337), .B(n3332), .C(n3303), .Y(n3338));
  INVX1   g2706(.A(n3338), .Y(n3339));
  NOR3X1  g2707(.A(n3339), .B(n3336), .C(n3331), .Y(n3340));
  INVX1   g2708(.A(n2414), .Y(n3341));
  NOR4X1  g2709(.A(n3298), .B(n3297), .C(n2323), .D(n3300), .Y(n3342));
  NAND3X1 g2710(.A(n3342), .B(n3341), .C(n2276), .Y(n3343));
  NOR4X1  g2711(.A(n3298), .B(n3297), .C(n2374), .D(n3300), .Y(n3344));
  NAND2X1 g2712(.A(n3344), .B(n2331), .Y(n3345));
  NOR2X1  g2713(.A(n3298), .B(n2420), .Y(n3346));
  AOI22X1 g2714(.A0(n2439), .A1(n2406), .B0(n2381), .B1(n3346), .Y(n3347));
  NOR2X1  g2715(.A(n3347), .B(n3300), .Y(n3348));
  AOI21X1 g2716(.A0(n2455), .A1(n3299), .B0(n3348), .Y(n3349));
  NAND3X1 g2717(.A(n3349), .B(n3345), .C(n3343), .Y(n3350));
  AOI21X1 g2718(.A0(n2285), .A1(n2242), .B0(n2291), .Y(n3351));
  NAND2X1 g2719(.A(n3321), .B(n1197), .Y(n3352));
  NOR4X1  g2720(.A(n3333), .B(n3315), .C(n3307), .D(n3352), .Y(n3353));
  NAND2X1 g2721(.A(n3353), .B(n3303), .Y(n3354));
  OAI21X1 g2722(.A0(n3351), .A1(n3304), .B0(n3354), .Y(n3355));
  NOR2X1  g2723(.A(n3355), .B(n3350), .Y(n3356));
  NOR4X1  g2724(.A(n3307), .B(n1982), .C(n1989), .D(n3333), .Y(n3357));
  NOR4X1  g2725(.A(n3302), .B(n2414), .C(n1864), .D(n3311), .Y(n3358));
  NAND4X1 g2726(.A(n3341), .B(n1950), .C(n1906), .D(n3301), .Y(n3359));
  INVX1   g2727(.A(n3359), .Y(n3360));
  OAI21X1 g2728(.A0(n3360), .A1(n3358), .B0(n3357), .Y(n3361));
  NAND3X1 g2729(.A(n3361), .B(n3356), .C(n3340), .Y(n3362));
  NOR2X1  g2730(.A(n3333), .B(n3307), .Y(n3363));
  NOR4X1  g2731(.A(n3315), .B(n1229), .C(n1218), .D(n3320), .Y(n3364));
  NAND4X1 g2732(.A(n3363), .B(n3301), .C(n3341), .D(n3364), .Y(n3365));
  NAND3X1 g2733(.A(n3312), .B(n3301), .C(n3826), .Y(n3366));
  NOR2X1  g2734(.A(n3366), .B(n2414), .Y(n3367));
  NAND2X1 g2735(.A(n3367), .B(n3363), .Y(n3368));
  NAND2X1 g2736(.A(n3313), .B(n3312), .Y(n3369));
  NOR4X1  g2737(.A(n3302), .B(n2414), .C(n1668), .D(n3369), .Y(n3370));
  NOR4X1  g2738(.A(n2414), .B(n1897), .C(n1884), .D(n3302), .Y(n3371));
  AOI22X1 g2739(.A0(n3370), .A1(n3363), .B0(n3357), .B1(n3371), .Y(n3372));
  NOR4X1  g2740(.A(n2073), .B(n2077), .C(n1981), .D(n2192), .Y(n3373));
  NOR3X1  g2741(.A(n3373), .B(n3302), .C(n2414), .Y(n3374));
  NAND2X1 g2742(.A(n3374), .B(n3363), .Y(n3375));
  INVX1   g2743(.A(n1027), .Y(n3376));
  NOR4X1  g2744(.A(n1181), .B(n1093), .C(n3376), .D(n2414), .Y(n3377));
  INVX1   g2745(.A(n3321), .Y(n3378));
  NOR4X1  g2746(.A(n3325), .B(n3378), .C(n3315), .D(n3333), .Y(n3379));
  NAND4X1 g2747(.A(n3377), .B(n3332), .C(n3301), .D(n3379), .Y(n3380));
  NAND2X1 g2748(.A(n3380), .B(n3375), .Y(n3381));
  INVX1   g2749(.A(n3363), .Y(n3382));
  OAI21X1 g2750(.A0(n1135), .A1(n1109), .B0(n1092), .Y(n3383));
  NOR3X1  g2751(.A(n3383), .B(n3302), .C(n2414), .Y(n3384));
  NAND3X1 g2752(.A(n3384), .B(n3379), .C(n3332), .Y(n3385));
  AOI21X1 g2753(.A0(n1702), .A1(n1689), .B0(n1705), .Y(n3386));
  NAND4X1 g2754(.A(n3312), .B(n3301), .C(n3341), .D(n3386), .Y(n3387));
  OAI21X1 g2755(.A0(n3387), .A1(n3382), .B0(n3385), .Y(n3388));
  NOR2X1  g2756(.A(n3388), .B(n3381), .Y(n3389));
  NAND4X1 g2757(.A(n3372), .B(n3368), .C(n3365), .D(n3389), .Y(n3390));
  NOR3X1  g2758(.A(n3318), .B(n2284), .C(n1512), .Y(n3391));
  NAND4X1 g2759(.A(n3334), .B(n3306), .C(n3305), .D(n3391), .Y(n3392));
  INVX1   g2760(.A(n3392), .Y(n3393));
  NOR4X1  g2761(.A(n2414), .B(n1397), .C(n1392), .D(n3302), .Y(n3394));
  NAND2X1 g2762(.A(n3394), .B(n3393), .Y(n3395));
  OAI21X1 g2763(.A0(n1906), .A1(n3308), .B0(n3825), .Y(n3396));
  NOR4X1  g2764(.A(n3311), .B(n3302), .C(n2414), .D(n3396), .Y(n3397));
  NAND2X1 g2765(.A(n3397), .B(n3357), .Y(n3398));
  NOR3X1  g2766(.A(n1670), .B(n1588), .C(n1567), .Y(n3399));
  NAND4X1 g2767(.A(n3313), .B(n3312), .C(n3301), .D(n3399), .Y(n3400));
  NOR2X1  g2768(.A(n3400), .B(n2414), .Y(n3401));
  NOR4X1  g2769(.A(n2414), .B(n1982), .C(n1988), .D(n3302), .Y(n3402));
  OAI21X1 g2770(.A0(n3402), .A1(n3401), .B0(n3363), .Y(n3403));
  NAND4X1 g2771(.A(n3301), .B(n3341), .C(n1307), .D(n3316), .Y(n3404));
  NOR2X1  g2772(.A(n3404), .B(n3392), .Y(n3405));
  NAND2X1 g2773(.A(n3379), .B(n3332), .Y(n3406));
  NOR4X1  g2774(.A(n3302), .B(n2414), .C(n1180), .D(n3406), .Y(n3407));
  NOR2X1  g2775(.A(n998), .B(n957), .Y(n3408));
  NAND4X1 g2776(.A(n3301), .B(n3341), .C(n3408), .D(n3329), .Y(n3409));
  NOR4X1  g2777(.A(n1452), .B(n1358), .C(n1340), .D(n2414), .Y(n3410));
  NAND2X1 g2778(.A(n3410), .B(n3301), .Y(n3411));
  OAI22X1 g2779(.A0(n3409), .A1(n3406), .B0(n3392), .B1(n3411), .Y(n3412));
  NOR3X1  g2780(.A(n3412), .B(n3407), .C(n3405), .Y(n3413));
  NAND4X1 g2781(.A(n3403), .B(n3398), .C(n3395), .D(n3413), .Y(n3414));
  NOR3X1  g2782(.A(n3414), .B(n3390), .C(n3362), .Y(n3415));
  INVX1   g2783(.A(n3415), .Y(n3416));
  NAND2X1 g2784(.A(n3416), .B(n2402), .Y(n3417));
  NOR3X1  g2785(.A(n889), .B(n886), .C(n757), .Y(n3418));
  INVX1   g2786(.A(n3418), .Y(n3419));
  INVX1   g2787(.A(n2848), .Y(n3420));
  AOI22X1 g2788(.A0(n1002), .A1(n757), .B0(n3420), .B1(n1073), .Y(n3421));
  OAI21X1 g2789(.A0(n3419), .A1(n1057), .B0(n3421), .Y(n3422));
  NOR2X1  g2790(.A(n3299), .B(n2406), .Y(n3423));
  AOI21X1 g2791(.A0(n1078), .A1(n1076), .B0(n878), .Y(n3424));
  NOR2X1  g2792(.A(n3419), .B(n1091), .Y(n3425));
  OAI21X1 g2793(.A0(n1057), .A1(n876), .B0(n758), .Y(n3426));
  NOR3X1  g2794(.A(n3426), .B(n3425), .C(n3424), .Y(n3427));
  NAND2X1 g2795(.A(n3427), .B(n3422), .Y(n3428));
  AOI22X1 g2796(.A0(n1079), .A1(n757), .B0(n3420), .B1(n1135), .Y(n3429));
  OAI21X1 g2797(.A0(n3419), .A1(n1109), .B0(n3429), .Y(n3430));
  AOI21X1 g2798(.A0(n1121), .A1(n1119), .B0(n878), .Y(n3431));
  NOR2X1  g2799(.A(n3419), .B(n1127), .Y(n3432));
  OAI21X1 g2800(.A0(n1109), .A1(n876), .B0(n758), .Y(n3433));
  NOR3X1  g2801(.A(n3433), .B(n3432), .C(n3431), .Y(n3434));
  OAI21X1 g2802(.A0(n1019), .A1(n1016), .B0(n3418), .Y(n3435));
  AOI22X1 g2803(.A0(n3420), .A1(n974), .B0(n986), .B1(n757), .Y(n3436));
  NAND2X1 g2804(.A(n3436), .B(n3435), .Y(n3437));
  AOI21X1 g2805(.A0(n956), .A1(n953), .B0(n878), .Y(n3438));
  NOR2X1  g2806(.A(n3419), .B(n998), .Y(n3439));
  OAI21X1 g2807(.A0(n1020), .A1(n876), .B0(n758), .Y(n3440));
  NOR3X1  g2808(.A(n3440), .B(n3439), .C(n3438), .Y(n3441));
  AOI22X1 g2809(.A0(n3437), .A1(n3441), .B0(n3434), .B1(n3430), .Y(n3442));
  AOI21X1 g2810(.A0(n986), .A1(n886), .B0(n757), .Y(n3444));
  OAI21X1 g2811(.A0(n3419), .A1(n959), .B0(n3444), .Y(n3445));
  AOI21X1 g2812(.A0(n986), .A1(n889), .B0(n3445), .Y(n3446));
  OAI22X1 g2813(.A0(n2848), .A1(n959), .B0(n929), .B1(n3419), .Y(n3447));
  NAND3X1 g2814(.A(n3447), .B(n3446), .C(n3441), .Y(n3448));
  AOI22X1 g2815(.A0(n3420), .A1(n909), .B0(n986), .B1(n3418), .Y(n3449));
  AOI21X1 g2816(.A0(n3436), .A1(n3435), .B0(n3449), .Y(n3450));
  AOI22X1 g2817(.A0(n957), .A1(n757), .B0(n3420), .B1(n1012), .Y(n3451));
  OAI21X1 g2818(.A0(n3419), .A1(n1034), .B0(n3451), .Y(n3452));
  AOI21X1 g2819(.A0(n1001), .A1(n1000), .B0(n878), .Y(n3453));
  NOR2X1  g2820(.A(n3419), .B(n1026), .Y(n3454));
  OAI21X1 g2821(.A0(n1034), .A1(n876), .B0(n758), .Y(n3455));
  NOR3X1  g2822(.A(n3455), .B(n3454), .C(n3453), .Y(n3456));
  AOI22X1 g2823(.A0(n3452), .A1(n3456), .B0(n3450), .B1(n3446), .Y(n3457));
  NAND4X1 g2824(.A(n3448), .B(n3442), .C(n3428), .D(n3457), .Y(n3458));
  NAND2X1 g2825(.A(n3434), .B(n3430), .Y(n3459));
  OAI22X1 g2826(.A0(n1020), .A1(n758), .B0(n2848), .B1(n1026), .Y(n3460));
  AOI21X1 g2827(.A0(n3418), .A1(n1002), .B0(n3460), .Y(n3461));
  OAI21X1 g2828(.A0(n1033), .A1(n1030), .B0(n889), .Y(n3462));
  NAND2X1 g2829(.A(n3418), .B(n1012), .Y(n3463));
  AOI21X1 g2830(.A0(n1002), .A1(n886), .B0(n757), .Y(n3464));
  NAND3X1 g2831(.A(n3464), .B(n3463), .C(n3462), .Y(n3465));
  NAND4X1 g2832(.A(n3461), .B(n3459), .C(n3428), .D(n3465), .Y(n3466));
  NOR2X1  g2833(.A(n3427), .B(n3422), .Y(n3467));
  NAND2X1 g2834(.A(n3467), .B(n3459), .Y(n3468));
  AOI21X1 g2835(.A0(n1195), .A1(n1193), .B0(n878), .Y(n3469));
  NOR2X1  g2836(.A(n3419), .B(n1188), .Y(n3470));
  OAI21X1 g2837(.A0(n1167), .A1(n876), .B0(n758), .Y(n3471));
  NOR3X1  g2838(.A(n3471), .B(n3470), .C(n3469), .Y(n3472));
  AOI22X1 g2839(.A0(n1122), .A1(n757), .B0(n3420), .B1(n1178), .Y(n3473));
  OAI21X1 g2840(.A0(n3419), .A1(n1167), .B0(n3473), .Y(n3474));
  OAI22X1 g2841(.A0(n3472), .A1(n3474), .B0(n3434), .B1(n3430), .Y(n3475));
  AOI21X1 g2842(.A0(n1273), .A1(n1269), .B0(n878), .Y(n3476));
  NOR2X1  g2843(.A(n3419), .B(n1300), .Y(n3477));
  OAI21X1 g2844(.A0(n1298), .A1(n876), .B0(n758), .Y(n3478));
  NOR3X1  g2845(.A(n3478), .B(n3477), .C(n3476), .Y(n3479));
  AOI22X1 g2846(.A0(n1218), .A1(n757), .B0(n3420), .B1(n1292), .Y(n3480));
  OAI21X1 g2847(.A0(n3419), .A1(n1298), .B0(n3480), .Y(n3481));
  AOI21X1 g2848(.A0(n1217), .A1(n1213), .B0(n878), .Y(n3482));
  NOR2X1  g2849(.A(n3419), .B(n1229), .Y(n3483));
  OAI21X1 g2850(.A0(n1285), .A1(n876), .B0(n758), .Y(n3484));
  NOR3X1  g2851(.A(n3484), .B(n3483), .C(n3482), .Y(n3485));
  AOI22X1 g2852(.A0(n1196), .A1(n757), .B0(n3420), .B1(n1252), .Y(n3486));
  OAI21X1 g2853(.A0(n3419), .A1(n1285), .B0(n3486), .Y(n3487));
  OAI22X1 g2854(.A0(n3485), .A1(n3487), .B0(n3481), .B1(n3479), .Y(n3488));
  NOR2X1  g2855(.A(n3488), .B(n3475), .Y(n3489));
  NAND4X1 g2856(.A(n3468), .B(n3466), .C(n3458), .D(n3489), .Y(n3490));
  AOI21X1 g2857(.A0(n1274), .A1(n886), .B0(n757), .Y(n3491));
  OAI21X1 g2858(.A0(n3419), .A1(n1300), .B0(n3491), .Y(n3492));
  OAI22X1 g2859(.A0(n1285), .A1(n758), .B0(n2848), .B1(n1300), .Y(n3493));
  AOI21X1 g2860(.A0(n3418), .A1(n1274), .B0(n3493), .Y(n3494));
  OAI21X1 g2861(.A0(n3492), .A1(n3476), .B0(n3494), .Y(n3495));
  AOI21X1 g2862(.A0(n1218), .A1(n886), .B0(n757), .Y(n3496));
  OAI21X1 g2863(.A0(n3419), .A1(n1229), .B0(n3496), .Y(n3497));
  OAI22X1 g2864(.A0(n1167), .A1(n758), .B0(n2848), .B1(n1229), .Y(n3498));
  AOI21X1 g2865(.A0(n3418), .A1(n1218), .B0(n3498), .Y(n3499));
  OAI21X1 g2866(.A0(n3497), .A1(n3482), .B0(n3499), .Y(n3500));
  NAND4X1 g2867(.A(n3495), .B(n3474), .C(n3472), .D(n3500), .Y(n3501));
  NAND3X1 g2868(.A(n3487), .B(n3485), .C(n3495), .Y(n3502));
  OAI22X1 g2869(.A0(n1383), .A1(n758), .B0(n2848), .B1(n1449), .Y(n3503));
  AOI21X1 g2870(.A0(n3418), .A1(n1444), .B0(n3503), .Y(n3504));
  AOI21X1 g2871(.A0(n1443), .A1(n1441), .B0(n878), .Y(n3505));
  AOI21X1 g2872(.A0(n1444), .A1(n886), .B0(n757), .Y(n3506));
  OAI21X1 g2873(.A0(n3419), .A1(n1449), .B0(n3506), .Y(n3507));
  NOR3X1  g2874(.A(n3507), .B(n3505), .C(n3504), .Y(n3508));
  AOI21X1 g2875(.A0(n1391), .A1(n1390), .B0(n3419), .Y(n3509));
  OAI22X1 g2876(.A0(n1339), .A1(n758), .B0(n2848), .B1(n1397), .Y(n3510));
  NOR2X1  g2877(.A(n3510), .B(n3509), .Y(n3511));
  AOI21X1 g2878(.A0(n1391), .A1(n1390), .B0(n878), .Y(n3512));
  NOR2X1  g2879(.A(n3419), .B(n1397), .Y(n3513));
  OAI21X1 g2880(.A0(n1383), .A1(n876), .B0(n758), .Y(n3514));
  NOR4X1  g2881(.A(n3513), .B(n3512), .C(n3511), .D(n3514), .Y(n3515));
  AOI22X1 g2882(.A0(n1274), .A1(n757), .B0(n3420), .B1(n1354), .Y(n3516));
  OAI21X1 g2883(.A0(n3419), .A1(n1339), .B0(n3516), .Y(n3517));
  NOR2X1  g2884(.A(n1339), .B(n878), .Y(n3518));
  NOR2X1  g2885(.A(n3419), .B(n1358), .Y(n3519));
  OAI21X1 g2886(.A0(n1339), .A1(n876), .B0(n758), .Y(n3520));
  NOR3X1  g2887(.A(n3520), .B(n3519), .C(n3518), .Y(n3521));
  NAND2X1 g2888(.A(n3521), .B(n3517), .Y(n3522));
  NAND2X1 g2889(.A(n3481), .B(n3479), .Y(n3523));
  NAND2X1 g2890(.A(n3523), .B(n3522), .Y(n3524));
  NOR3X1  g2891(.A(n3524), .B(n3515), .C(n3508), .Y(n3525));
  NAND4X1 g2892(.A(n3502), .B(n3501), .C(n3490), .D(n3525), .Y(n3526));
  NOR4X1  g2893(.A(n3517), .B(n3515), .C(n3508), .D(n3521), .Y(n3527));
  NOR3X1  g2894(.A(n3514), .B(n3513), .C(n3512), .Y(n3528));
  NOR4X1  g2895(.A(n3510), .B(n3509), .C(n3508), .D(n3528), .Y(n3529));
  AOI21X1 g2896(.A0(n1593), .A1(n1589), .B0(n878), .Y(n3530));
  AOI21X1 g2897(.A0(n1594), .A1(n886), .B0(n757), .Y(n3531));
  OAI21X1 g2898(.A0(n3419), .A1(n1606), .B0(n3531), .Y(n3532));
  OAI22X1 g2899(.A0(n1547), .A1(n758), .B0(n2848), .B1(n1606), .Y(n3533));
  AOI21X1 g2900(.A0(n3418), .A1(n1594), .B0(n3533), .Y(n3534));
  OAI21X1 g2901(.A0(n3532), .A1(n3530), .B0(n3534), .Y(n3535));
  AOI21X1 g2902(.A0(n1566), .A1(n1564), .B0(n878), .Y(n3536));
  AOI21X1 g2903(.A0(n1567), .A1(n886), .B0(n757), .Y(n3537));
  OAI21X1 g2904(.A0(n3419), .A1(n1588), .B0(n3537), .Y(n3538));
  OAI22X1 g2905(.A0(n1490), .A1(n758), .B0(n2848), .B1(n1588), .Y(n3539));
  AOI21X1 g2906(.A0(n3418), .A1(n1567), .B0(n3539), .Y(n3540));
  OAI21X1 g2907(.A0(n3538), .A1(n3536), .B0(n3540), .Y(n3541));
  AOI21X1 g2908(.A0(n1501), .A1(n1499), .B0(n878), .Y(n3542));
  AOI21X1 g2909(.A0(n1502), .A1(n886), .B0(n757), .Y(n3543));
  OAI21X1 g2910(.A0(n3419), .A1(n1507), .B0(n3543), .Y(n3544));
  OAI22X1 g2911(.A0(n1434), .A1(n758), .B0(n2848), .B1(n1507), .Y(n3545));
  AOI21X1 g2912(.A0(n3418), .A1(n1502), .B0(n3545), .Y(n3546));
  OAI21X1 g2913(.A0(n3544), .A1(n3542), .B0(n3546), .Y(n3547));
  OAI21X1 g2914(.A0(n3507), .A1(n3505), .B0(n3504), .Y(n3548));
  NAND4X1 g2915(.A(n3547), .B(n3541), .C(n3535), .D(n3548), .Y(n3549));
  NOR3X1  g2916(.A(n3549), .B(n3529), .C(n3527), .Y(n3550));
  NOR3X1  g2917(.A(n3546), .B(n3544), .C(n3542), .Y(n3551));
  NAND3X1 g2918(.A(n3551), .B(n3541), .C(n3535), .Y(n3552));
  NOR3X1  g2919(.A(n3540), .B(n3538), .C(n3536), .Y(n3553));
  NAND2X1 g2920(.A(n3553), .B(n3535), .Y(n3554));
  NOR2X1  g2921(.A(n3532), .B(n3530), .Y(n3555));
  AOI22X1 g2922(.A0(n1567), .A1(n757), .B0(n3420), .B1(n1620), .Y(n3556));
  OAI21X1 g2923(.A0(n3419), .A1(n1595), .B0(n3556), .Y(n3557));
  NOR2X1  g2924(.A(n1645), .B(n878), .Y(n3559));
  NOR2X1  g2925(.A(n3419), .B(n1681), .Y(n3560));
  OAI21X1 g2926(.A0(n1645), .A1(n876), .B0(n758), .Y(n3561));
  NOR3X1  g2927(.A(n3561), .B(n3560), .C(n3559), .Y(n3562));
  AOI22X1 g2928(.A0(n1594), .A1(n757), .B0(n3420), .B1(n1662), .Y(n3563));
  OAI21X1 g2929(.A0(n3419), .A1(n1645), .B0(n3563), .Y(n3564));
  AOI22X1 g2930(.A0(n3562), .A1(n3564), .B0(n3557), .B1(n3555), .Y(n3565));
  NAND3X1 g2931(.A(n3565), .B(n3554), .C(n3552), .Y(n3566));
  AOI21X1 g2932(.A0(n3550), .A1(n3526), .B0(n3566), .Y(n3567));
  AOI22X1 g2933(.A0(n1710), .A1(n757), .B0(n3420), .B1(n1744), .Y(n3568));
  OAI21X1 g2934(.A0(n3419), .A1(n1690), .B0(n3568), .Y(n3569));
  AOI21X1 g2935(.A0(n1688), .A1(n1683), .B0(n878), .Y(n3570));
  NOR2X1  g2936(.A(n3419), .B(n1702), .Y(n3571));
  AOI21X1 g2937(.A0(n1688), .A1(n1683), .B0(n876), .Y(n3572));
  NOR4X1  g2938(.A(n3571), .B(n3570), .C(n757), .D(n3572), .Y(n3573));
  OAI22X1 g2939(.A0(n3569), .A1(n3573), .B0(n3564), .B1(n3562), .Y(n3574));
  AOI21X1 g2940(.A0(n1735), .A1(n1728), .B0(n878), .Y(n3575));
  NOR2X1  g2941(.A(n3419), .B(n1751), .Y(n3576));
  OAI21X1 g2942(.A0(n1737), .A1(n876), .B0(n758), .Y(n3577));
  OAI22X1 g2943(.A0(n1690), .A1(n758), .B0(n2848), .B1(n1751), .Y(n3578));
  AOI21X1 g2944(.A0(n3418), .A1(n1736), .B0(n3578), .Y(n3579));
  NOR4X1  g2945(.A(n3577), .B(n3576), .C(n3575), .D(n3579), .Y(n3580));
  AOI21X1 g2946(.A0(n3573), .A1(n3569), .B0(n3580), .Y(n3581));
  OAI21X1 g2947(.A0(n3574), .A1(n3567), .B0(n3581), .Y(n3582));
  NOR3X1  g2948(.A(n3577), .B(n3576), .C(n3575), .Y(n3583));
  AOI21X1 g2949(.A0(n1735), .A1(n1728), .B0(n3419), .Y(n3584));
  NOR3X1  g2950(.A(n3578), .B(n3584), .C(n3583), .Y(n3585));
  OAI22X1 g2951(.A0(n1737), .A1(n758), .B0(n2848), .B1(n1806), .Y(n3586));
  AOI21X1 g2952(.A0(n3418), .A1(n1789), .B0(n3586), .Y(n3587));
  AOI21X1 g2953(.A0(n1788), .A1(n1783), .B0(n878), .Y(n3588));
  INVX1   g2954(.A(n3588), .Y(n3589));
  NAND2X1 g2955(.A(n3418), .B(n1828), .Y(n3590));
  AOI21X1 g2956(.A0(n1789), .A1(n886), .B0(n757), .Y(n3591));
  NAND3X1 g2957(.A(n3591), .B(n3590), .C(n3589), .Y(n3592));
  AOI21X1 g2958(.A0(n3592), .A1(n3587), .B0(n3585), .Y(n3593));
  NOR2X1  g2959(.A(n3592), .B(n3587), .Y(n3594));
  AOI21X1 g2960(.A0(n1836), .A1(n1831), .B0(n878), .Y(n3595));
  NOR2X1  g2961(.A(n3419), .B(n1854), .Y(n3596));
  AOI21X1 g2962(.A0(n1836), .A1(n1831), .B0(n876), .Y(n3597));
  NOR4X1  g2963(.A(n3596), .B(n3595), .C(n757), .D(n3597), .Y(n3598));
  AOI22X1 g2964(.A0(n1789), .A1(n757), .B0(n3420), .B1(n1857), .Y(n3599));
  OAI21X1 g2965(.A0(n3419), .A1(n1838), .B0(n3599), .Y(n3600));
  AOI21X1 g2966(.A0(n3600), .A1(n3598), .B0(n3594), .Y(n3601));
  INVX1   g2967(.A(n3601), .Y(n3602));
  AOI21X1 g2968(.A0(n3593), .A1(n3582), .B0(n3602), .Y(n3603));
  AOI22X1 g2969(.A0(n1900), .A1(n3420), .B0(n1884), .B1(n3418), .Y(n3604));
  OAI21X1 g2970(.A0(n1838), .A1(n758), .B0(n3604), .Y(n3605));
  AOI21X1 g2971(.A0(n1883), .A1(n1877), .B0(n878), .Y(n3606));
  NOR2X1  g2972(.A(n3419), .B(n1897), .Y(n3607));
  AOI21X1 g2973(.A0(n1883), .A1(n1877), .B0(n876), .Y(n3608));
  NOR4X1  g2974(.A(n3607), .B(n3606), .C(n757), .D(n3608), .Y(n3609));
  OAI22X1 g2975(.A0(n3605), .A1(n3609), .B0(n3600), .B1(n3598), .Y(n3610));
  NOR2X1  g2976(.A(n1926), .B(n878), .Y(n3611));
  AOI21X1 g2977(.A0(n3418), .A1(n1935), .B0(n757), .Y(n3612));
  OAI21X1 g2978(.A0(n1926), .A1(n876), .B0(n3612), .Y(n3613));
  NOR2X1  g2979(.A(n3613), .B(n3611), .Y(n3614));
  AOI22X1 g2980(.A0(n1884), .A1(n757), .B0(n3420), .B1(n1935), .Y(n3615));
  OAI21X1 g2981(.A0(n3419), .A1(n1926), .B0(n3615), .Y(n3616));
  AOI22X1 g2982(.A0(n3614), .A1(n3616), .B0(n3609), .B1(n3605), .Y(n3617));
  OAI21X1 g2983(.A0(n3610), .A1(n3603), .B0(n3617), .Y(n3618));
  NOR2X1  g2984(.A(n3616), .B(n3614), .Y(n3619));
  AOI22X1 g2985(.A0(n1973), .A1(n3420), .B0(n1964), .B1(n3418), .Y(n3620));
  OAI21X1 g2986(.A0(n1926), .A1(n758), .B0(n3620), .Y(n3621));
  NOR2X1  g2987(.A(n1965), .B(n878), .Y(n3622));
  AOI21X1 g2988(.A0(n3418), .A1(n1973), .B0(n757), .Y(n3623));
  OAI21X1 g2989(.A0(n1965), .A1(n876), .B0(n3623), .Y(n3624));
  NOR2X1  g2990(.A(n3624), .B(n3622), .Y(n3625));
  NOR2X1  g2991(.A(n3625), .B(n3621), .Y(n3626));
  NOR2X1  g2992(.A(n3626), .B(n3619), .Y(n3627));
  NOR2X1  g2993(.A(n2009), .B(n878), .Y(n3628));
  AOI21X1 g2994(.A0(n3418), .A1(n2017), .B0(n757), .Y(n3629));
  OAI21X1 g2995(.A0(n2009), .A1(n876), .B0(n3629), .Y(n3630));
  NOR2X1  g2996(.A(n3630), .B(n3628), .Y(n3631));
  AOI22X1 g2997(.A0(n1964), .A1(n757), .B0(n3420), .B1(n2017), .Y(n3632));
  OAI21X1 g2998(.A0(n3419), .A1(n2009), .B0(n3632), .Y(n3633));
  AOI22X1 g2999(.A0(n3631), .A1(n3633), .B0(n3625), .B1(n3621), .Y(n3634));
  INVX1   g3000(.A(n3634), .Y(n3635));
  AOI21X1 g3001(.A0(n3627), .A1(n3618), .B0(n3635), .Y(n3636));
  AOI22X1 g3002(.A0(n2076), .A1(n757), .B0(n3420), .B1(n2066), .Y(n3637));
  OAI21X1 g3003(.A0(n3419), .A1(n2056), .B0(n3637), .Y(n3638));
  NOR2X1  g3004(.A(n2056), .B(n878), .Y(n3639));
  AOI21X1 g3005(.A0(n3418), .A1(n2066), .B0(n757), .Y(n3640));
  OAI21X1 g3006(.A0(n2056), .A1(n876), .B0(n3640), .Y(n3641));
  NOR2X1  g3007(.A(n3641), .B(n3639), .Y(n3642));
  OAI22X1 g3008(.A0(n3638), .A1(n3642), .B0(n3633), .B1(n3631), .Y(n3643));
  NOR2X1  g3009(.A(n2118), .B(n878), .Y(n3644));
  AOI21X1 g3010(.A0(n3418), .A1(n2126), .B0(n757), .Y(n3645));
  OAI21X1 g3011(.A0(n2118), .A1(n876), .B0(n3645), .Y(n3646));
  NOR2X1  g3012(.A(n3646), .B(n3644), .Y(n3647));
  AOI22X1 g3013(.A0(n2071), .A1(n757), .B0(n3420), .B1(n2126), .Y(n3648));
  OAI21X1 g3014(.A0(n3419), .A1(n2118), .B0(n3648), .Y(n3649));
  AOI22X1 g3015(.A0(n3647), .A1(n3649), .B0(n3642), .B1(n3638), .Y(n3650));
  OAI21X1 g3016(.A0(n3643), .A1(n3636), .B0(n3650), .Y(n3651));
  NOR2X1  g3017(.A(n3649), .B(n3647), .Y(n3652));
  AOI22X1 g3018(.A0(n2181), .A1(n757), .B0(n3420), .B1(n2178), .Y(n3653));
  OAI21X1 g3019(.A0(n3419), .A1(n2170), .B0(n3653), .Y(n3654));
  NAND2X1 g3020(.A(n2230), .B(n889), .Y(n3655));
  OAI21X1 g3021(.A0(n3419), .A1(n2186), .B0(n758), .Y(n3656));
  AOI21X1 g3022(.A0(n2230), .A1(n886), .B0(n3656), .Y(n3657));
  AOI21X1 g3023(.A0(n3657), .A1(n3655), .B0(n3654), .Y(n3658));
  NOR2X1  g3024(.A(n3658), .B(n3652), .Y(n3659));
  NAND3X1 g3025(.A(n3657), .B(n3655), .C(n3654), .Y(n3660));
  NOR2X1  g3026(.A(n2283), .B(n878), .Y(n3661));
  AOI21X1 g3027(.A0(n3418), .A1(n2229), .B0(n757), .Y(n3662));
  OAI21X1 g3028(.A0(n2283), .A1(n876), .B0(n3662), .Y(n3663));
  NOR2X1  g3029(.A(n3663), .B(n3661), .Y(n3664));
  AOI22X1 g3030(.A0(n2230), .A1(n757), .B0(n3420), .B1(n2229), .Y(n3665));
  OAI21X1 g3031(.A0(n3419), .A1(n2283), .B0(n3665), .Y(n3666));
  NAND2X1 g3032(.A(n3666), .B(n3664), .Y(n3667));
  NAND2X1 g3033(.A(n3667), .B(n3660), .Y(n3668));
  AOI21X1 g3034(.A0(n3659), .A1(n3651), .B0(n3668), .Y(n3669));
  AOI22X1 g3035(.A0(n2221), .A1(n757), .B0(n3420), .B1(n2287), .Y(n3670));
  OAI21X1 g3036(.A0(n3419), .A1(n2276), .B0(n3670), .Y(n3671));
  NOR2X1  g3037(.A(n2276), .B(n878), .Y(n3672));
  AOI21X1 g3038(.A0(n3418), .A1(n2287), .B0(n757), .Y(n3673));
  OAI21X1 g3039(.A0(n2276), .A1(n876), .B0(n3673), .Y(n3674));
  NOR2X1  g3040(.A(n3674), .B(n3672), .Y(n3675));
  OAI22X1 g3041(.A0(n3671), .A1(n3675), .B0(n3666), .B1(n3664), .Y(n3676));
  AOI21X1 g3042(.A0(n3418), .A1(n2339), .B0(n757), .Y(n3679));
  OAI21X1 g3043(.A0(n2331), .A1(n876), .B0(n3679), .Y(n3680));
  AOI21X1 g3044(.A0(n2393), .A1(n889), .B0(n3680), .Y(n3681));
  AOI22X1 g3045(.A0(n2342), .A1(n757), .B0(n3420), .B1(n2339), .Y(n3682));
  OAI21X1 g3046(.A0(n3419), .A1(n2331), .B0(n3682), .Y(n3683));
  AOI22X1 g3047(.A0(n3681), .A1(n3683), .B0(n3675), .B1(n3671), .Y(n3684));
  OAI21X1 g3048(.A0(n3676), .A1(n3669), .B0(n3684), .Y(n3685));
  AOI22X1 g3049(.A0(n2389), .A1(n3420), .B0(n2747), .B1(n3418), .Y(n3686));
  OAI21X1 g3050(.A0(n2331), .A1(n758), .B0(n3686), .Y(n3687));
  AOI21X1 g3051(.A0(n2379), .A1(n3296), .B0(n878), .Y(n3688));
  AOI21X1 g3052(.A0(n2379), .A1(n3296), .B0(n876), .Y(n3689));
  OAI21X1 g3053(.A0(n3419), .A1(n2420), .B0(n758), .Y(n3690));
  NOR3X1  g3054(.A(n3690), .B(n3689), .C(n3688), .Y(n3691));
  OAI22X1 g3055(.A0(n3687), .A1(n3691), .B0(n3683), .B1(n3681), .Y(n3692));
  INVX1   g3056(.A(n3692), .Y(n3693));
  INVX1   g3057(.A(n2406), .Y(n3694));
  NAND3X1 g3058(.A(n3299), .B(n3694), .C(n889), .Y(n3695));
  AOI22X1 g3059(.A0(n2439), .A1(n3418), .B0(n3694), .B1(n886), .Y(n3696));
  NAND2X1 g3060(.A(n3696), .B(n3695), .Y(n3697));
  INVX1   g3061(.A(n3697), .Y(n3698));
  AOI22X1 g3062(.A0(n2439), .A1(n3420), .B0(n3694), .B1(n3418), .Y(n3699));
  INVX1   g3063(.A(n3699), .Y(n3700));
  AOI22X1 g3064(.A0(n3698), .A1(n3700), .B0(n3691), .B1(n3687), .Y(n3701));
  INVX1   g3065(.A(n3701), .Y(n3702));
  AOI21X1 g3066(.A0(n3693), .A1(n3685), .B0(n3702), .Y(n3703));
  AOI22X1 g3067(.A0(n2452), .A1(n3420), .B0(n3299), .B1(n3418), .Y(n3704));
  INVX1   g3068(.A(n3704), .Y(n3705));
  OAI22X1 g3069(.A0(n2455), .A1(n3419), .B0(n2444), .B1(n876), .Y(n3707));
  AOI21X1 g3070(.A0(n3299), .A1(n889), .B0(n3707), .Y(n3708));
  XOR2X1  g3071(.A(n3708), .B(n3705), .Y(n3709));
  OAI21X1 g3072(.A0(n3700), .A1(n3698), .B0(n3709), .Y(n3710));
  NOR3X1  g3073(.A(n3704), .B(n3420), .C(n758), .Y(n3711));
  OAI21X1 g3074(.A0(n3420), .A1(n758), .B0(n3704), .Y(n3712));
  NOR2X1  g3075(.A(n3712), .B(n3708), .Y(n3713));
  AOI21X1 g3076(.A0(n3711), .A1(n3708), .B0(n3713), .Y(n3714));
  OAI21X1 g3077(.A0(n3710), .A1(n3703), .B0(n3714), .Y(n3715));
  OAI21X1 g3078(.A0(n3715), .A1(n2402), .B0(n3417), .Y(n3716));
  OAI22X1 g3079(.A0(n1034), .A1(n758), .B0(n2848), .B1(n1091), .Y(n3717));
  AOI21X1 g3080(.A0(n3418), .A1(n1079), .B0(n3717), .Y(n3718));
  NOR4X1  g3081(.A(n3425), .B(n3424), .C(n3718), .D(n3426), .Y(n3719));
  OAI22X1 g3082(.A0(n1057), .A1(n758), .B0(n2848), .B1(n1127), .Y(n3720));
  AOI21X1 g3083(.A0(n3418), .A1(n1122), .B0(n3720), .Y(n3721));
  OAI21X1 g3084(.A0(n1108), .A1(n1105), .B0(n889), .Y(n3722));
  NAND2X1 g3085(.A(n3418), .B(n1135), .Y(n3723));
  AOI21X1 g3086(.A0(n1122), .A1(n886), .B0(n757), .Y(n3724));
  NAND3X1 g3087(.A(n3724), .B(n3723), .C(n3722), .Y(n3725));
  AOI21X1 g3088(.A0(n956), .A1(n953), .B0(n3419), .Y(n3726));
  OAI22X1 g3089(.A0(n2848), .A1(n998), .B0(n929), .B1(n758), .Y(n3727));
  NOR2X1  g3090(.A(n3727), .B(n3726), .Y(n3728));
  OAI21X1 g3091(.A0(n1019), .A1(n1016), .B0(n889), .Y(n3729));
  NAND2X1 g3092(.A(n3418), .B(n974), .Y(n3730));
  AOI21X1 g3093(.A0(n957), .A1(n886), .B0(n757), .Y(n3731));
  NAND3X1 g3094(.A(n3731), .B(n3730), .C(n3729), .Y(n3732));
  OAI22X1 g3095(.A0(n3728), .A1(n3732), .B0(n3725), .B1(n3721), .Y(n3733));
  NAND2X1 g3096(.A(n986), .B(n889), .Y(n3734));
  NAND2X1 g3097(.A(n3418), .B(n909), .Y(n3735));
  NAND3X1 g3098(.A(n3444), .B(n3735), .C(n3734), .Y(n3736));
  NOR3X1  g3099(.A(n3449), .B(n3736), .C(n3732), .Y(n3737));
  OAI21X1 g3100(.A0(n3727), .A1(n3726), .B0(n3447), .Y(n3738));
  OAI22X1 g3101(.A0(n3461), .A1(n3465), .B0(n3738), .B1(n3736), .Y(n3739));
  NOR4X1  g3102(.A(n3737), .B(n3733), .C(n3719), .D(n3739), .Y(n3740));
  NOR2X1  g3103(.A(n3725), .B(n3721), .Y(n3741));
  NOR4X1  g3104(.A(n3452), .B(n3741), .C(n3719), .D(n3456), .Y(n3742));
  NOR3X1  g3105(.A(n3741), .B(n3427), .C(n3422), .Y(n3743));
  NAND2X1 g3106(.A(n3725), .B(n3721), .Y(n3744));
  AOI21X1 g3107(.A0(n1196), .A1(n886), .B0(n757), .Y(n3745));
  OAI21X1 g3108(.A0(n3419), .A1(n1188), .B0(n3745), .Y(n3746));
  OAI22X1 g3109(.A0(n1109), .A1(n758), .B0(n2848), .B1(n1188), .Y(n3747));
  AOI21X1 g3110(.A0(n3418), .A1(n1196), .B0(n3747), .Y(n3748));
  OAI21X1 g3111(.A0(n3746), .A1(n3469), .B0(n3748), .Y(n3749));
  NAND4X1 g3112(.A(n3495), .B(n3749), .C(n3744), .D(n3500), .Y(n3750));
  NOR4X1  g3113(.A(n3743), .B(n3742), .C(n3740), .D(n3750), .Y(n3751));
  NOR2X1  g3114(.A(n3515), .B(n3508), .Y(n3752));
  AOI22X1 g3115(.A0(n3517), .A1(n3521), .B0(n3481), .B1(n3479), .Y(n3753));
  NAND4X1 g3116(.A(n3752), .B(n3502), .C(n3501), .D(n3753), .Y(n3754));
  OAI21X1 g3117(.A0(n3754), .A1(n3751), .B0(n3550), .Y(n3755));
  NOR2X1  g3118(.A(n3557), .B(n3555), .Y(n3756));
  NOR4X1  g3119(.A(n3544), .B(n3542), .C(n3756), .D(n3546), .Y(n3757));
  NAND2X1 g3120(.A(n3565), .B(n3554), .Y(n3758));
  AOI21X1 g3121(.A0(n3757), .A1(n3541), .B0(n3758), .Y(n3759));
  AOI21X1 g3122(.A0(n3759), .A1(n3755), .B0(n3574), .Y(n3760));
  INVX1   g3123(.A(n3581), .Y(n3761));
  OAI21X1 g3124(.A0(n3761), .A1(n3760), .B0(n3593), .Y(n3762));
  AOI21X1 g3125(.A0(n3601), .A1(n3762), .B0(n3610), .Y(n3763));
  INVX1   g3126(.A(n3617), .Y(n3764));
  OAI21X1 g3127(.A0(n3764), .A1(n3763), .B0(n3627), .Y(n3765));
  AOI21X1 g3128(.A0(n3634), .A1(n3765), .B0(n3643), .Y(n3766));
  INVX1   g3129(.A(n3650), .Y(n3767));
  OAI21X1 g3130(.A0(n3767), .A1(n3766), .B0(n3659), .Y(n3768));
  NAND3X1 g3131(.A(n3667), .B(n3660), .C(n3768), .Y(n3769));
  INVX1   g3132(.A(n3676), .Y(n3770));
  INVX1   g3133(.A(n3684), .Y(n3771));
  AOI21X1 g3134(.A0(n3770), .A1(n3769), .B0(n3771), .Y(n3772));
  OAI21X1 g3135(.A0(n3692), .A1(n3772), .B0(n3701), .Y(n3773));
  INVX1   g3136(.A(n3710), .Y(n3774));
  AOI21X1 g3137(.A0(n3774), .A1(n3773), .B0(n3713), .Y(n3776));
  NAND3X1 g3138(.A(n889), .B(n876), .C(n884), .Y(n3777));
  XOR2X1  g3139(.A(n1973), .B(n1964), .Y(n3781));
  XOR2X1  g3140(.A(n1935), .B(n1925), .Y(n3782));
  XOR2X1  g3141(.A(n2440), .B(n2406), .Y(n3783));
  XOR2X1  g3142(.A(n2455), .B(n2444), .Y(n3784));
  NOR4X1  g3143(.A(n3783), .B(n3782), .C(n3781), .D(n3784), .Y(n3785));
  NOR4X1  g3144(.A(n1529), .B(n1418), .C(n1359), .D(n1856), .Y(n3786));
  XOR2X1  g3145(.A(n1449), .B(n1434), .Y(n3787));
  NOR4X1  g3146(.A(n1901), .B(n1568), .C(n1136), .D(n3787), .Y(n3788));
  NAND4X1 g3147(.A(n3786), .B(n3785), .C(n2067), .D(n3788), .Y(n3789));
  XOR2X1  g3148(.A(n1292), .B(n1274), .Y(n3790));
  XOR2X1  g3149(.A(n929), .B(n959), .Y(n3791));
  NOR4X1  g3150(.A(n3790), .B(n1770), .C(n1253), .D(n3791), .Y(n3792));
  XOR2X1  g3151(.A(n1620), .B(n1594), .Y(n3793));
  XOR2X1  g3152(.A(n1681), .B(n1645), .Y(n3794));
  XOR2X1  g3153(.A(n1744), .B(n1689), .Y(n3795));
  NOR4X1  g3154(.A(n3794), .B(n3793), .C(n975), .D(n3795), .Y(n3796));
  XOR2X1  g3155(.A(n1178), .B(n1196), .Y(n3798));
  XOR2X1  g3156(.A(n1828), .B(n1789), .Y(n3799));
  NOR4X1  g3157(.A(n3798), .B(n1080), .C(n1013), .D(n3799), .Y(n3800));
  NAND4X1 g3158(.A(n2018), .B(n3796), .C(n3792), .D(n3800), .Y(n3801));
  NOR4X1  g3159(.A(n3789), .B(n2187), .C(n2157), .D(n3801), .Y(n3802));
  XOR2X1  g3160(.A(n2229), .B(n2221), .Y(n3803));
  XOR2X1  g3161(.A(n2420), .B(n2381), .Y(n3804));
  NOR2X1  g3162(.A(n3804), .B(n3803), .Y(n3805));
  NAND4X1 g3163(.A(n3802), .B(n2288), .C(n2340), .D(n3805), .Y(n3806));
  OAI22X1 g3164(.A0(n3777), .A1(n3776), .B0(n890), .B1(n3806), .Y(n3807));
  AOI21X1 g3165(.A0(n3716), .A1(n878), .B0(n3807), .Y(n3808));
  NOR2X1  g3166(.A(n1864), .B(n3311), .Y(n3811));
  OAI22X1 g3167(.A0(n2076), .A1(n2047), .B0(n1974), .B1(n1964), .Y(n3812));
  NAND2X1 g3168(.A(n1857), .B(n1838), .Y(n3814));
  NOR2X1  g3169(.A(n3814), .B(n1949), .Y(n3815));
  OAI22X1 g3170(.A0(n1925), .A1(n1941), .B0(n1897), .B1(n1884), .Y(n3816));
  NOR4X1  g3171(.A(n3815), .B(n3812), .C(n3811), .D(n3816), .Y(n3817));
  NAND2X1 g3172(.A(n1513), .B(n3314), .Y(n3820));
  OAI22X1 g3173(.A0(n1710), .A1(n1681), .B0(n1606), .B1(n1594), .Y(n3824));
  NOR2X1  g3174(.A(n1751), .B(n1736), .Y(n3825));
  NOR2X1  g3175(.A(n1702), .B(n1689), .Y(n3826));
  NOR4X1  g3176(.A(n3825), .B(n3824), .C(n3399), .D(n3826), .Y(n3827));
  NAND3X1 g3177(.A(n3827), .B(n3820), .C(n3817), .Y(n3828));
  OAI22X1 g3178(.A0(n1383), .A1(n1451), .B0(n1354), .B1(n1339), .Y(n3829));
  AOI22X1 g3179(.A0(n1434), .A1(n1461), .B0(n1451), .B1(n1383), .Y(n3830));
  NAND2X1 g3180(.A(n3830), .B(n3829), .Y(n3831));
  NAND2X1 g3181(.A(n1401), .B(n3830), .Y(n3833));
  AOI22X1 g3182(.A0(n1285), .A1(n1252), .B0(n1178), .B1(n1167), .Y(n3834));
  INVX1   g3183(.A(n3834), .Y(n3835));
  NOR2X1  g3184(.A(n1127), .B(n1122), .Y(n3836));
  NAND2X1 g3185(.A(n1091), .B(n1079), .Y(n3837));
  NOR4X1  g3186(.A(n3836), .B(n3835), .C(n3833), .D(n3837), .Y(n3838));
  NAND4X1 g3187(.A(n3827), .B(n3820), .C(n3817), .D(n3838), .Y(n3839));
  INVX1   g3188(.A(n3839), .Y(n3840));
  NOR4X1  g3189(.A(n3836), .B(n3835), .C(n3833), .D(n1092), .Y(n3842));
  NAND2X1 g3190(.A(n1035), .B(n3842), .Y(n3844));
  NOR2X1  g3191(.A(n3844), .B(n3828), .Y(n3845));
  NOR2X1  g3192(.A(n3845), .B(n3840), .Y(n3846));
  OAI21X1 g3193(.A0(n3831), .A1(n3828), .B0(n3846), .Y(n3847));
  INVX1   g3194(.A(n1512), .Y(n3849));
  NOR2X1  g3195(.A(n974), .B(n1020), .Y(n3850));
  NOR3X1  g3196(.A(n3850), .B(n986), .C(n959), .Y(n3851));
  OAI22X1 g3197(.A0(n1002), .A1(n1026), .B0(n998), .B1(n957), .Y(n3852));
  NOR2X1  g3198(.A(n3852), .B(n3851), .Y(n3853));
  NAND2X1 g3199(.A(n3853), .B(n3842), .Y(n3854));
  AOI21X1 g3200(.A0(n3854), .A1(n3849), .B0(n3828), .Y(n3855));
  INVX1   g3201(.A(n1515), .Y(n3857));
  AOI22X1 g3202(.A0(n1196), .A1(n1188), .B0(n1127), .B1(n1122), .Y(n3858));
  AOI22X1 g3203(.A0(n1274), .A1(n1300), .B0(n1229), .B1(n1218), .Y(n3859));
  OAI21X1 g3204(.A0(n3858), .A1(n3835), .B0(n3859), .Y(n3860));
  NAND3X1 g3205(.A(n3860), .B(n1401), .C(n3830), .Y(n3861));
  AOI21X1 g3206(.A0(n3861), .A1(n3857), .B0(n3828), .Y(n3862));
  NOR2X1  g3207(.A(n1769), .B(n1737), .Y(n3863));
  NOR4X1  g3208(.A(n3825), .B(n1645), .C(n1662), .D(n3826), .Y(n3864));
  OAI21X1 g3209(.A0(n3864), .A1(n3863), .B0(n3817), .Y(n3865));
  OAI21X1 g3210(.A0(n1865), .A1(n3311), .B0(n3817), .Y(n3867));
  INVX1   g3211(.A(n3314), .Y(n3868));
  NAND4X1 g3212(.A(n3820), .B(n3868), .C(n3817), .D(n3827), .Y(n3869));
  INVX1   g3213(.A(n3817), .Y(n3870));
  NOR2X1  g3214(.A(n1744), .B(n1690), .Y(n3872));
  NAND2X1 g3215(.A(n3872), .B(n1816), .Y(n3873));
  NOR2X1  g3216(.A(n3873), .B(n3870), .Y(n3874));
  NAND2X1 g3217(.A(n1974), .B(n1964), .Y(n3876));
  OAI21X1 g3218(.A0(n3876), .A1(n2077), .B0(n2074), .Y(n3878));
  NAND2X1 g3219(.A(n1941), .B(n1925), .Y(n3881));
  OAI21X1 g3220(.A0(n3881), .A1(n3812), .B0(n2194), .Y(n3882));
  NOR3X1  g3221(.A(n3882), .B(n3878), .C(n3874), .Y(n3883));
  NAND4X1 g3222(.A(n3869), .B(n3867), .C(n3865), .D(n3883), .Y(n3884));
  NOR4X1  g3223(.A(n3862), .B(n3855), .C(n3847), .D(n3884), .Y(n3885));
  AOI21X1 g3224(.A0(n2073), .A1(n2194), .B0(n2192), .Y(n3888));
  INVX1   g3225(.A(n3888), .Y(n3889));
  NOR2X1  g3226(.A(n3889), .B(n3885), .Y(n3890));
  NOR2X1  g3227(.A(n3890), .B(n2186), .Y(n3891));
  NOR2X1  g3228(.A(n2323), .B(n2342), .Y(n3894));
  AOI21X1 g3229(.A0(n3299), .A1(n3694), .B0(n2440), .Y(n3895));
  NOR3X1  g3230(.A(n3423), .B(n2452), .C(n2444), .Y(n3896));
  NOR3X1  g3231(.A(n3896), .B(n3895), .C(n2389), .Y(n3897));
  NOR3X1  g3232(.A(n3896), .B(n3895), .C(n2381), .Y(n3899));
  NOR2X1  g3233(.A(n3899), .B(n3897), .Y(n3900));
  NOR3X1  g3234(.A(n3900), .B(n3894), .C(n2339), .Y(n3901));
  NOR2X1  g3235(.A(n3901), .B(n2393), .Y(n3902));
  OAI22X1 g3236(.A0(n2221), .A1(n2233), .B0(n2186), .B1(n2230), .Y(n3903));
  NOR4X1  g3237(.A(n3902), .B(n3900), .C(n3894), .D(n3903), .Y(n3904));
  OAI21X1 g3238(.A0(n3890), .A1(n2230), .B0(n3904), .Y(n3905));
  NOR2X1  g3239(.A(n3905), .B(n3891), .Y(n3906));
  NOR3X1  g3240(.A(n3900), .B(n3894), .C(n2331), .Y(n3907));
  NOR2X1  g3241(.A(n3907), .B(n3901), .Y(n3908));
  AOI22X1 g3242(.A0(n2342), .A1(n2323), .B0(n2233), .B1(n2221), .Y(n3909));
  NOR3X1  g3243(.A(n3900), .B(n2331), .C(n2339), .Y(n3910));
  NOR4X1  g3244(.A(n3895), .B(n2381), .C(n2389), .D(n3896), .Y(n3911));
  NOR4X1  g3245(.A(n2444), .B(n2439), .C(n2406), .D(n2455), .Y(n3913));
  NOR4X1  g3246(.A(n3300), .B(n3911), .C(n3910), .D(n3913), .Y(n3914));
  OAI21X1 g3247(.A0(n3909), .A1(n3908), .B0(n3914), .Y(n3915));
  OAI21X1 g3248(.A0(n3915), .A1(n3906), .B0(n936), .Y(n3916));
  NOR2X1  g3249(.A(n3915), .B(n3906), .Y(n3917));
  NOR4X1  g3250(.A(n878), .B(n876), .C(n873), .D(n938), .Y(n3918));
  NAND2X1 g3251(.A(n3918), .B(n3917), .Y(n3919));
  NOR3X1  g3252(.A(n881), .B(n889), .C(n873), .Y(n3920));
  NOR3X1  g3253(.A(n881), .B(n878), .C(n884), .Y(n3921));
  AOI22X1 g3254(.A0(n3806), .A1(n3921), .B0(n3415), .B1(n3920), .Y(n3922));
  NAND3X1 g3255(.A(n3922), .B(n3919), .C(n3916), .Y(n3923));
  AOI21X1 g3256(.A0(n3776), .A1(n2526), .B0(n3923), .Y(n3924));
  OAI21X1 g3257(.A0(n3808), .A1(n938), .B0(n3924), .Y(n3925));
  NOR3X1  g3258(.A(n3419), .B(n3416), .C(n881), .Y(n3926));
  AOI21X1 g3259(.A0(n3925), .A1(n758), .B0(n3926), .Y(n3927));
  NOR3X1  g3260(.A(n938), .B(n889), .C(n873), .Y(n3928));
  INVX1   g3261(.A(n3928), .Y(n3929));
  NOR3X1  g3262(.A(n2936), .B(n3929), .C(n886), .Y(n3930));
  NOR2X1  g3263(.A(n886), .B(n757), .Y(n3931));
  NOR3X1  g3264(.A(n3931), .B(n2842), .C(U3149), .Y(n3932));
  OAI21X1 g3265(.A0(n3930), .A1(n758), .B0(n3932), .Y(n3933));
  NOR4X1  g3266(.A(n3929), .B(n886), .C(n769), .D(n2936), .Y(n3934));
  AOI22X1 g3267(.A0(n3933), .A1(B_REG_SCAN_IN), .B0(n3715), .B1(n3934), .Y(n3935));
  OAI21X1 g3268(.A0(n3927), .A1(U3149), .B0(n3935), .Y(U3239));
  AOI22X1 g3269(.A0(n3145), .A1(n1710), .B0(n1662), .B1(n3156), .Y(n3937));
  OAI22X1 g3270(.A0(n3146), .A1(n1645), .B0(n1681), .B1(n3155), .Y(n3938));
  XOR2X1  g3271(.A(n3938), .B(n3152), .Y(n3939));
  NOR2X1  g3272(.A(n3939), .B(n3937), .Y(n3940));
  NAND2X1 g3273(.A(n3939), .B(n3937), .Y(n3941));
  AOI22X1 g3274(.A0(n3145), .A1(n1392), .B0(n1451), .B1(n3156), .Y(n3942));
  OAI21X1 g3275(.A0(n3138), .A1(n3150), .B0(n2841), .Y(n3943));
  OAI21X1 g3276(.A0(n3144), .A1(n767), .B0(n3943), .Y(n3944));
  AOI22X1 g3277(.A0(n3156), .A1(n1122), .B0(n1135), .B1(n3944), .Y(n3945));
  XOR2X1  g3278(.A(n3945), .B(n3152), .Y(n3946));
  INVX1   g3279(.A(n3946), .Y(n3947));
  AOI22X1 g3280(.A0(n3145), .A1(n1122), .B0(n1135), .B1(n3156), .Y(n3948));
  AOI22X1 g3281(.A0(n3145), .A1(n1002), .B0(n1012), .B1(n3156), .Y(n3949));
  AOI22X1 g3282(.A0(n3156), .A1(n1002), .B0(n1012), .B1(n3944), .Y(n3950));
  XOR2X1  g3283(.A(n3950), .B(n3140), .Y(n3951));
  AOI22X1 g3284(.A0(n3145), .A1(n1079), .B0(n1073), .B1(n3156), .Y(n3952));
  AOI22X1 g3285(.A0(n3156), .A1(n1079), .B0(n1073), .B1(n3944), .Y(n3953));
  XOR2X1  g3286(.A(n3953), .B(n3140), .Y(n3954));
  AOI22X1 g3287(.A0(n3952), .A1(n3954), .B0(n3951), .B1(n3949), .Y(n3955));
  AOI22X1 g3288(.A0(n3156), .A1(n957), .B0(n974), .B1(n3944), .Y(n3956));
  XOR2X1  g3289(.A(n3956), .B(n3152), .Y(n3957));
  OAI21X1 g3290(.A0(n3153), .A1(n3138), .B0(n2841), .Y(n3958));
  OAI22X1 g3291(.A0(n3958), .A1(n1020), .B0(n998), .B1(n3146), .Y(n3959));
  NOR2X1  g3292(.A(n3959), .B(n3957), .Y(n3960));
  NOR3X1  g3293(.A(n3960), .B(n3148), .C(n3152), .Y(n3961));
  AOI22X1 g3294(.A0(n909), .A1(n3156), .B0(n907), .B1(n767), .Y(n3962));
  OAI21X1 g3295(.A0(n3958), .A1(n929), .B0(n3962), .Y(n3963));
  XOR2X1  g3296(.A(n3158), .B(n3140), .Y(n3964));
  OAI21X1 g3297(.A0(n3963), .A1(n3140), .B0(n3964), .Y(n3965));
  NAND2X1 g3298(.A(n3959), .B(n3957), .Y(n3966));
  OAI21X1 g3299(.A0(n3965), .A1(n3960), .B0(n3966), .Y(n3967));
  OAI21X1 g3300(.A0(n3967), .A1(n3961), .B0(n3955), .Y(n3968));
  INVX1   g3301(.A(n3952), .Y(n3969));
  NOR2X1  g3302(.A(n3951), .B(n3949), .Y(n3970));
  OAI22X1 g3303(.A0(n3958), .A1(n1034), .B0(n1026), .B1(n3146), .Y(n3971));
  XOR2X1  g3304(.A(n3950), .B(n3152), .Y(n3972));
  NAND2X1 g3305(.A(n3972), .B(n3971), .Y(n3973));
  AOI21X1 g3306(.A0(n3973), .A1(n3952), .B0(n3954), .Y(n3974));
  AOI21X1 g3307(.A0(n3970), .A1(n3969), .B0(n3974), .Y(n3975));
  AOI22X1 g3308(.A0(n3968), .A1(n3975), .B0(n3948), .B1(n3947), .Y(n3976));
  NOR2X1  g3309(.A(n3948), .B(n3947), .Y(n3977));
  AOI22X1 g3310(.A0(n3156), .A1(n1340), .B0(n1354), .B1(n3944), .Y(n3978));
  XOR2X1  g3311(.A(n3978), .B(n3152), .Y(n3979));
  AOI22X1 g3312(.A0(n3145), .A1(n1340), .B0(n1354), .B1(n3156), .Y(n3980));
  INVX1   g3313(.A(n3980), .Y(n3981));
  NOR2X1  g3314(.A(n3981), .B(n3979), .Y(n3982));
  AOI22X1 g3315(.A0(n3145), .A1(n1218), .B0(n1252), .B1(n3156), .Y(n3983));
  AOI22X1 g3316(.A0(n3156), .A1(n1218), .B0(n1252), .B1(n3944), .Y(n3984));
  XOR2X1  g3317(.A(n3984), .B(n3140), .Y(n3985));
  AOI22X1 g3318(.A0(n3145), .A1(n1274), .B0(n1292), .B1(n3156), .Y(n3986));
  AOI22X1 g3319(.A0(n3156), .A1(n1274), .B0(n1292), .B1(n3944), .Y(n3987));
  XOR2X1  g3320(.A(n3987), .B(n3140), .Y(n3988));
  AOI22X1 g3321(.A0(n3986), .A1(n3988), .B0(n3985), .B1(n3983), .Y(n3989));
  AOI22X1 g3322(.A0(n3145), .A1(n1196), .B0(n1178), .B1(n3156), .Y(n3990));
  AOI22X1 g3323(.A0(n3156), .A1(n1196), .B0(n1178), .B1(n3944), .Y(n3991));
  XOR2X1  g3324(.A(n3991), .B(n3140), .Y(n3992));
  NAND2X1 g3325(.A(n3992), .B(n3990), .Y(n3993));
  NAND2X1 g3326(.A(n3993), .B(n3989), .Y(n3994));
  NOR2X1  g3327(.A(n3994), .B(n3982), .Y(n3995));
  OAI21X1 g3328(.A0(n3977), .A1(n3976), .B0(n3995), .Y(n3996));
  INVX1   g3329(.A(n3986), .Y(n3997));
  XOR2X1  g3330(.A(n3987), .B(n3152), .Y(n3998));
  NOR2X1  g3331(.A(n3985), .B(n3983), .Y(n3999));
  OAI21X1 g3332(.A0(n3999), .A1(n3997), .B0(n3998), .Y(n4000));
  NOR2X1  g3333(.A(n3992), .B(n3990), .Y(n4001));
  AOI22X1 g3334(.A0(n3999), .A1(n3997), .B0(n3989), .B1(n4001), .Y(n4002));
  AOI21X1 g3335(.A0(n4002), .A1(n4000), .B0(n3982), .Y(n4003));
  AOI21X1 g3336(.A0(n3981), .A1(n3979), .B0(n4003), .Y(n4004));
  AOI21X1 g3337(.A0(n4004), .A1(n3996), .B0(n3942), .Y(n4005));
  AOI22X1 g3338(.A0(n3156), .A1(n1392), .B0(n1451), .B1(n3944), .Y(n4006));
  XOR2X1  g3339(.A(n4006), .B(n3140), .Y(n4007));
  NOR2X1  g3340(.A(n4007), .B(n3942), .Y(n4008));
  AOI21X1 g3341(.A0(n4004), .A1(n3996), .B0(n4007), .Y(n4009));
  NOR3X1  g3342(.A(n4009), .B(n4008), .C(n4005), .Y(n4010));
  AOI22X1 g3343(.A0(n3156), .A1(n1567), .B0(n1561), .B1(n3944), .Y(n4011));
  XOR2X1  g3344(.A(n4011), .B(n3140), .Y(n4012));
  AOI22X1 g3345(.A0(n3145), .A1(n1567), .B0(n1561), .B1(n3156), .Y(n4013));
  AOI22X1 g3346(.A0(n3156), .A1(n1594), .B0(n1620), .B1(n3944), .Y(n4014));
  XOR2X1  g3347(.A(n4014), .B(n3140), .Y(n4015));
  AOI22X1 g3348(.A0(n3145), .A1(n1594), .B0(n1620), .B1(n3156), .Y(n4016));
  AOI22X1 g3349(.A0(n4015), .A1(n4016), .B0(n4013), .B1(n4012), .Y(n4017));
  AOI22X1 g3350(.A0(n3156), .A1(n1502), .B0(n1514), .B1(n3944), .Y(n4018));
  XOR2X1  g3351(.A(n4018), .B(n3140), .Y(n4019));
  INVX1   g3352(.A(n4019), .Y(n4020));
  AOI22X1 g3353(.A0(n3145), .A1(n1502), .B0(n1514), .B1(n3156), .Y(n4021));
  INVX1   g3354(.A(n4021), .Y(n4022));
  NOR2X1  g3355(.A(n4022), .B(n4020), .Y(n4023));
  INVX1   g3356(.A(n4023), .Y(n4024));
  AOI22X1 g3357(.A0(n3145), .A1(n1444), .B0(n1461), .B1(n3156), .Y(n4025));
  OAI22X1 g3358(.A0(n3146), .A1(n1434), .B0(n1449), .B1(n3155), .Y(n4026));
  XOR2X1  g3359(.A(n4026), .B(n3152), .Y(n4027));
  NAND2X1 g3360(.A(n4027), .B(n4025), .Y(n4028));
  NAND3X1 g3361(.A(n4028), .B(n4024), .C(n4017), .Y(n4029));
  INVX1   g3362(.A(n4015), .Y(n4030));
  INVX1   g3363(.A(n4016), .Y(n4031));
  NOR2X1  g3364(.A(n4031), .B(n4030), .Y(n4032));
  INVX1   g3365(.A(n4032), .Y(n4033));
  INVX1   g3366(.A(n4017), .Y(n4034));
  NOR4X1  g3367(.A(n4025), .B(n4023), .C(n4034), .D(n4027), .Y(n4035));
  NAND2X1 g3368(.A(n4022), .B(n4020), .Y(n4036));
  INVX1   g3369(.A(n4012), .Y(n4037));
  INVX1   g3370(.A(n4013), .Y(n4038));
  AOI22X1 g3371(.A0(n4030), .A1(n4031), .B0(n4038), .B1(n4037), .Y(n4039));
  OAI21X1 g3372(.A0(n4036), .A1(n4034), .B0(n4039), .Y(n4040));
  AOI21X1 g3373(.A0(n4040), .A1(n4033), .B0(n4035), .Y(n4041));
  OAI21X1 g3374(.A0(n4029), .A1(n4010), .B0(n4041), .Y(n4042));
  AOI21X1 g3375(.A0(n4042), .A1(n3941), .B0(n3940), .Y(n4043));
  AOI22X1 g3376(.A0(n3156), .A1(n1689), .B0(n1744), .B1(n3944), .Y(n4044));
  XOR2X1  g3377(.A(n4044), .B(n3140), .Y(n4045));
  AOI22X1 g3378(.A0(n3145), .A1(n1689), .B0(n1744), .B1(n3156), .Y(n4046));
  XOR2X1  g3379(.A(n4046), .B(n4045), .Y(n4047));
  XOR2X1  g3380(.A(n4047), .B(n4043), .Y(n4048));
  NOR3X1  g3381(.A(n893), .B(n870), .C(n2527), .Y(n4049));
  NOR4X1  g3382(.A(n2847), .B(n946), .C(n945), .D(n3918), .Y(n4050));
  OAI21X1 g3383(.A0(n3920), .A1(n936), .B0(n886), .Y(n4051));
  AOI21X1 g3384(.A0(n881), .A1(n878), .B0(n886), .Y(n4052));
  NAND2X1 g3385(.A(n4052), .B(n873), .Y(n4053));
  NAND3X1 g3386(.A(n4053), .B(n4051), .C(n4050), .Y(n4054));
  NAND3X1 g3387(.A(n4054), .B(n4049), .C(n768), .Y(n4055));
  INVX1   g3388(.A(n4049), .Y(n4056));
  NOR4X1  g3389(.A(n767), .B(n758), .C(U3149), .D(n963), .Y(n4057));
  INVX1   g3390(.A(n2528), .Y(n4058));
  NAND3X1 g3391(.A(n4058), .B(n2841), .C(n757), .Y(n4059));
  AOI21X1 g3392(.A0(n4054), .A1(n4056), .B0(n4059), .Y(n4060));
  NOR2X1  g3393(.A(n4060), .B(U3149), .Y(n4061));
  AOI21X1 g3394(.A0(n4057), .A1(n4056), .B0(n4061), .Y(n4062));
  INVX1   g3395(.A(n4062), .Y(n4063));
  NOR3X1  g3396(.A(n3929), .B(n886), .C(n769), .Y(n4064));
  INVX1   g3397(.A(n4064), .Y(n4065));
  NOR4X1  g3398(.A(n893), .B(n870), .C(n2527), .D(n2943), .Y(n4066));
  NOR4X1  g3399(.A(n893), .B(n870), .C(n2527), .D(n991), .Y(n4067));
  INVX1   g3400(.A(n4067), .Y(n4068));
  OAI22X1 g3401(.A0(n4049), .A1(n1686), .B0(n1645), .B1(n4068), .Y(n4069));
  AOI21X1 g3402(.A0(n4066), .A1(n1736), .B0(n4069), .Y(n4070));
  AOI22X1 g3403(.A0(n4049), .A1(n4057), .B0(n2526), .B1(n768), .Y(n4071));
  INVX1   g3404(.A(n4071), .Y(n4072));
  AOI22X1 g3405(.A0(n1744), .A1(n4072), .B0(REG3_REG_15__SCAN_IN), .B1(U3149), .Y(n4073));
  OAI21X1 g3406(.A0(n4070), .A1(n4065), .B0(n4073), .Y(n4074));
  AOI21X1 g3407(.A0(n4063), .A1(n2644), .B0(n4074), .Y(n4075));
  OAI21X1 g3408(.A0(n4055), .A1(n4048), .B0(n4075), .Y(U3238));
  OAI22X1 g3409(.A0(n3146), .A1(n2170), .B0(n2186), .B1(n3155), .Y(n4077));
  XOR2X1  g3410(.A(n4077), .B(n3152), .Y(n4078));
  INVX1   g3411(.A(n4078), .Y(n4079));
  AOI22X1 g3412(.A0(n3145), .A1(n2230), .B0(n2178), .B1(n3156), .Y(n4080));
  INVX1   g3413(.A(n4080), .Y(n4081));
  NOR2X1  g3414(.A(n4081), .B(n4079), .Y(n4082));
  INVX1   g3415(.A(n4082), .Y(n4083));
  AOI22X1 g3416(.A0(n3145), .A1(n2181), .B0(n2126), .B1(n3156), .Y(n4084));
  OAI22X1 g3417(.A0(n3146), .A1(n2118), .B0(n2156), .B1(n3155), .Y(n4085));
  XOR2X1  g3418(.A(n4085), .B(n3152), .Y(n4086));
  NOR2X1  g3419(.A(n4086), .B(n4084), .Y(n4087));
  INVX1   g3420(.A(n4087), .Y(n4088));
  NAND2X1 g3421(.A(n4086), .B(n4084), .Y(n4089));
  INVX1   g3422(.A(n4089), .Y(n4090));
  AOI22X1 g3423(.A0(n3145), .A1(n2071), .B0(n2066), .B1(n3156), .Y(n4091));
  OAI22X1 g3424(.A0(n3146), .A1(n2056), .B0(n2072), .B1(n3155), .Y(n4092));
  XOR2X1  g3425(.A(n4092), .B(n3152), .Y(n4093));
  NOR2X1  g3426(.A(n4093), .B(n4091), .Y(n4094));
  NAND2X1 g3427(.A(n4093), .B(n4091), .Y(n4095));
  AOI22X1 g3428(.A0(n3145), .A1(n2076), .B0(n2017), .B1(n3156), .Y(n4096));
  OAI22X1 g3429(.A0(n3146), .A1(n2009), .B0(n2047), .B1(n3155), .Y(n4097));
  XOR2X1  g3430(.A(n4097), .B(n3152), .Y(n4098));
  NOR2X1  g3431(.A(n4098), .B(n4096), .Y(n4099));
  INVX1   g3432(.A(n4099), .Y(n4100));
  NAND2X1 g3433(.A(n4098), .B(n4096), .Y(n4101));
  INVX1   g3434(.A(n4101), .Y(n4102));
  AOI22X1 g3435(.A0(n3156), .A1(n1964), .B0(n1973), .B1(n3944), .Y(n4103));
  XOR2X1  g3436(.A(n4103), .B(n3140), .Y(n4104));
  INVX1   g3437(.A(n4104), .Y(n4105));
  AOI22X1 g3438(.A0(n3145), .A1(n1964), .B0(n1973), .B1(n3156), .Y(n4106));
  INVX1   g3439(.A(n4106), .Y(n4107));
  NOR2X1  g3440(.A(n4107), .B(n4105), .Y(n4108));
  INVX1   g3441(.A(n4108), .Y(n4109));
  AOI22X1 g3442(.A0(n3145), .A1(n1884), .B0(n1900), .B1(n3156), .Y(n4110));
  AOI22X1 g3443(.A0(n3156), .A1(n1884), .B0(n1900), .B1(n3944), .Y(n4111));
  XOR2X1  g3444(.A(n4111), .B(n3140), .Y(n4112));
  NOR2X1  g3445(.A(n4112), .B(n4110), .Y(n4113));
  INVX1   g3446(.A(n4113), .Y(n4114));
  AOI22X1 g3447(.A0(n3145), .A1(n1925), .B0(n1935), .B1(n3156), .Y(n4115));
  AOI22X1 g3448(.A0(n3156), .A1(n1925), .B0(n1935), .B1(n3944), .Y(n4116));
  XOR2X1  g3449(.A(n4116), .B(n3140), .Y(n4117));
  AOI22X1 g3450(.A0(n4115), .A1(n4117), .B0(n4106), .B1(n4104), .Y(n4118));
  INVX1   g3451(.A(n4118), .Y(n4119));
  NOR2X1  g3452(.A(n4117), .B(n4115), .Y(n4120));
  AOI21X1 g3453(.A0(n4107), .A1(n4105), .B0(n4120), .Y(n4121));
  OAI21X1 g3454(.A0(n4119), .A1(n4114), .B0(n4121), .Y(n4122));
  AOI22X1 g3455(.A0(n3145), .A1(n1837), .B0(n1857), .B1(n3156), .Y(n4123));
  AOI22X1 g3456(.A0(n3156), .A1(n1837), .B0(n1857), .B1(n3944), .Y(n4124));
  XOR2X1  g3457(.A(n4124), .B(n3140), .Y(n4125));
  NOR2X1  g3458(.A(n4125), .B(n4123), .Y(n4126));
  INVX1   g3459(.A(n4126), .Y(n4127));
  NAND2X1 g3460(.A(n4125), .B(n4123), .Y(n4128));
  INVX1   g3461(.A(n4128), .Y(n4129));
  AOI22X1 g3462(.A0(n3145), .A1(n1736), .B0(n1769), .B1(n3156), .Y(n4130));
  AOI22X1 g3463(.A0(n3156), .A1(n1736), .B0(n1769), .B1(n3944), .Y(n4131));
  XOR2X1  g3464(.A(n4131), .B(n3140), .Y(n4132));
  AOI22X1 g3465(.A0(n3145), .A1(n1789), .B0(n1828), .B1(n3156), .Y(n4133));
  AOI22X1 g3466(.A0(n3156), .A1(n1789), .B0(n1828), .B1(n3944), .Y(n4134));
  XOR2X1  g3467(.A(n4134), .B(n3140), .Y(n4135));
  AOI22X1 g3468(.A0(n4133), .A1(n4135), .B0(n4132), .B1(n4130), .Y(n4136));
  NOR2X1  g3469(.A(n4046), .B(n4045), .Y(n4137));
  INVX1   g3470(.A(n4137), .Y(n4138));
  NAND2X1 g3471(.A(n4046), .B(n4045), .Y(n4139));
  INVX1   g3472(.A(n4139), .Y(n4140));
  OAI21X1 g3473(.A0(n4140), .A1(n4043), .B0(n4138), .Y(n4141));
  INVX1   g3474(.A(n4133), .Y(n4142));
  NOR2X1  g3475(.A(n4132), .B(n4130), .Y(n4143));
  INVX1   g3476(.A(n4143), .Y(n4144));
  AOI21X1 g3477(.A0(n4144), .A1(n4133), .B0(n4135), .Y(n4145));
  AOI21X1 g3478(.A0(n4143), .A1(n4142), .B0(n4145), .Y(n4146));
  INVX1   g3479(.A(n4146), .Y(n4147));
  AOI21X1 g3480(.A0(n4141), .A1(n4136), .B0(n4147), .Y(n4148));
  OAI21X1 g3481(.A0(n4148), .A1(n4129), .B0(n4127), .Y(n4149));
  AOI21X1 g3482(.A0(n4112), .A1(n4110), .B0(n4119), .Y(n4150));
  AOI22X1 g3483(.A0(n4149), .A1(n4150), .B0(n4122), .B1(n4109), .Y(n4151));
  OAI21X1 g3484(.A0(n4151), .A1(n4102), .B0(n4100), .Y(n4152));
  AOI21X1 g3485(.A0(n4152), .A1(n4095), .B0(n4094), .Y(n4153));
  OAI21X1 g3486(.A0(n4153), .A1(n4090), .B0(n4088), .Y(n4154));
  AOI22X1 g3487(.A0(n3145), .A1(n2221), .B0(n2229), .B1(n3156), .Y(n4155));
  OAI22X1 g3488(.A0(n3146), .A1(n2283), .B0(n2233), .B1(n3155), .Y(n4156));
  XOR2X1  g3489(.A(n4156), .B(n3152), .Y(n4157));
  INVX1   g3490(.A(n4157), .Y(n4158));
  NOR2X1  g3491(.A(n4080), .B(n4078), .Y(n4159));
  AOI21X1 g3492(.A0(n4158), .A1(n4155), .B0(n4159), .Y(n4160));
  OAI21X1 g3493(.A0(n4158), .A1(n4155), .B0(n4160), .Y(n4161));
  AOI21X1 g3494(.A0(n4154), .A1(n4083), .B0(n4161), .Y(n4162));
  INVX1   g3495(.A(n4055), .Y(n4163));
  INVX1   g3496(.A(n4094), .Y(n4164));
  INVX1   g3497(.A(n4095), .Y(n4165));
  NAND2X1 g3498(.A(n4122), .B(n4109), .Y(n4166));
  INVX1   g3499(.A(n4136), .Y(n4167));
  INVX1   g3500(.A(n3940), .Y(n4168));
  INVX1   g3501(.A(n3941), .Y(n4169));
  INVX1   g3502(.A(n3942), .Y(n4170));
  INVX1   g3503(.A(n3948), .Y(n4171));
  XOR2X1  g3504(.A(n3953), .B(n3152), .Y(n4172));
  OAI22X1 g3505(.A0(n3969), .A1(n4172), .B0(n3972), .B1(n3971), .Y(n4173));
  XOR2X1  g3506(.A(n3956), .B(n3140), .Y(n4174));
  AOI22X1 g3507(.A0(n3145), .A1(n957), .B0(n974), .B1(n3156), .Y(n4175));
  NAND2X1 g3508(.A(n4175), .B(n4174), .Y(n4176));
  NOR2X1  g3509(.A(n3148), .B(n3152), .Y(n4177));
  NAND2X1 g3510(.A(n4177), .B(n4176), .Y(n4178));
  AOI21X1 g3511(.A0(n3148), .A1(n3152), .B0(n3159), .Y(n4179));
  NOR2X1  g3512(.A(n4175), .B(n4174), .Y(n4180));
  AOI21X1 g3513(.A0(n4179), .A1(n4176), .B0(n4180), .Y(n4181));
  AOI21X1 g3514(.A0(n4181), .A1(n4178), .B0(n4173), .Y(n4182));
  OAI21X1 g3515(.A0(n3970), .A1(n3969), .B0(n4172), .Y(n4183));
  OAI21X1 g3516(.A0(n3973), .A1(n3952), .B0(n4183), .Y(n4184));
  OAI22X1 g3517(.A0(n4182), .A1(n4184), .B0(n4171), .B1(n3946), .Y(n4185));
  INVX1   g3518(.A(n3977), .Y(n4186));
  INVX1   g3519(.A(n3983), .Y(n4187));
  XOR2X1  g3520(.A(n3984), .B(n3152), .Y(n4188));
  OAI22X1 g3521(.A0(n3997), .A1(n3998), .B0(n4188), .B1(n4187), .Y(n4189));
  AOI21X1 g3522(.A0(n3992), .A1(n3990), .B0(n4189), .Y(n4190));
  OAI21X1 g3523(.A0(n3981), .A1(n3979), .B0(n4190), .Y(n4191));
  AOI21X1 g3524(.A0(n4186), .A1(n4185), .B0(n4191), .Y(n4192));
  NAND2X1 g3525(.A(n4188), .B(n4187), .Y(n4193));
  AOI21X1 g3526(.A0(n4193), .A1(n3986), .B0(n3988), .Y(n4194));
  NAND2X1 g3527(.A(n4001), .B(n3989), .Y(n4195));
  OAI21X1 g3528(.A0(n4193), .A1(n3986), .B0(n4195), .Y(n4196));
  NOR2X1  g3529(.A(n4196), .B(n4194), .Y(n4197));
  NAND2X1 g3530(.A(n3981), .B(n3979), .Y(n4198));
  OAI21X1 g3531(.A0(n4197), .A1(n3982), .B0(n4198), .Y(n4199));
  OAI21X1 g3532(.A0(n4199), .A1(n4192), .B0(n4170), .Y(n4200));
  INVX1   g3533(.A(n4008), .Y(n4201));
  INVX1   g3534(.A(n4007), .Y(n4202));
  OAI21X1 g3535(.A0(n4199), .A1(n4192), .B0(n4202), .Y(n4203));
  NAND3X1 g3536(.A(n4203), .B(n4201), .C(n4200), .Y(n4204));
  INVX1   g3537(.A(n4029), .Y(n4205));
  INVX1   g3538(.A(n4041), .Y(n4206));
  AOI21X1 g3539(.A0(n4205), .A1(n4204), .B0(n4206), .Y(n4207));
  OAI21X1 g3540(.A0(n4207), .A1(n4169), .B0(n4168), .Y(n4208));
  AOI21X1 g3541(.A0(n4139), .A1(n4208), .B0(n4137), .Y(n4209));
  OAI21X1 g3542(.A0(n4209), .A1(n4167), .B0(n4146), .Y(n4210));
  AOI21X1 g3543(.A0(n4210), .A1(n4128), .B0(n4126), .Y(n4211));
  INVX1   g3544(.A(n4150), .Y(n4212));
  OAI21X1 g3545(.A0(n4212), .A1(n4211), .B0(n4166), .Y(n4213));
  AOI21X1 g3546(.A0(n4213), .A1(n4101), .B0(n4099), .Y(n4214));
  OAI21X1 g3547(.A0(n4214), .A1(n4165), .B0(n4164), .Y(n4215));
  OAI21X1 g3548(.A0(n4080), .A1(n4078), .B0(n4088), .Y(n4216));
  AOI21X1 g3549(.A0(n4215), .A1(n4089), .B0(n4216), .Y(n4217));
  AOI22X1 g3550(.A0(n4155), .A1(n4157), .B0(n4080), .B1(n4078), .Y(n4218));
  OAI21X1 g3551(.A0(n4157), .A1(n4155), .B0(n4218), .Y(n4219));
  OAI21X1 g3552(.A0(n4219), .A1(n4217), .B0(n4163), .Y(n4220));
  OAI21X1 g3553(.A0(n4049), .A1(n963), .B0(n4060), .Y(n4221));
  OAI22X1 g3554(.A0(n4049), .A1(n2217), .B0(n2170), .B1(n4068), .Y(n4224));
  AOI21X1 g3555(.A0(n4066), .A1(n2342), .B0(n4224), .Y(n4225));
  AOI22X1 g3556(.A0(n2229), .A1(n4072), .B0(REG3_REG_26__SCAN_IN), .B1(U3149), .Y(n4229));
  OAI21X1 g3557(.A0(n4225), .A1(n4065), .B0(n4229), .Y(n4230));
  AOI21X1 g3558(.A0(n4063), .A1(n2730), .B0(n4230), .Y(n4231));
  OAI21X1 g3559(.A0(n4220), .A1(n4162), .B0(n4231), .Y(U3237));
  XOR2X1  g3560(.A(n4188), .B(n4187), .Y(n4233));
  NOR2X1  g3561(.A(n3977), .B(n3976), .Y(n4234));
  INVX1   g3562(.A(n4234), .Y(n4235));
  AOI21X1 g3563(.A0(n3993), .A1(n4235), .B0(n4001), .Y(n4236));
  NOR2X1  g3564(.A(n4233), .B(n4236), .Y(n4238));
  AOI21X1 g3565(.A0(n4236), .A1(n4233), .B0(n4238), .Y(n4239));
  INVX1   g3566(.A(n4066), .Y(n4240));
  NOR2X1  g3567(.A(n4240), .B(n1298), .Y(n4241));
  OAI22X1 g3568(.A0(n4049), .A1(n1215), .B0(n1167), .B1(n4068), .Y(n4242));
  OAI21X1 g3569(.A0(n4242), .A1(n4241), .B0(n4064), .Y(n4243));
  AOI22X1 g3570(.A0(n1252), .A1(n4072), .B0(REG3_REG_6__SCAN_IN), .B1(U3149), .Y(n4244));
  NAND2X1 g3571(.A(n4244), .B(n4243), .Y(n4245));
  AOI21X1 g3572(.A0(n4063), .A1(n1216), .B0(n4245), .Y(n4246));
  OAI21X1 g3573(.A0(n4239), .A1(n4055), .B0(n4246), .Y(U3236));
  XOR2X1  g3574(.A(n4125), .B(n4123), .Y(n4248));
  XOR2X1  g3575(.A(n4248), .B(n4148), .Y(n4249));
  OAI22X1 g3576(.A0(n4049), .A1(n1834), .B0(n1790), .B1(n4068), .Y(n4250));
  AOI21X1 g3577(.A0(n4066), .A1(n1884), .B0(n4250), .Y(n4251));
  AOI22X1 g3578(.A0(n1857), .A1(n4072), .B0(REG3_REG_18__SCAN_IN), .B1(U3149), .Y(n4252));
  OAI21X1 g3579(.A0(n4251), .A1(n4065), .B0(n4252), .Y(n4253));
  AOI21X1 g3580(.A0(n4063), .A1(n2668), .B0(n4253), .Y(n4254));
  OAI21X1 g3581(.A0(n4249), .A1(n4055), .B0(n4254), .Y(U3235));
  NOR2X1  g3582(.A(n3967), .B(n3961), .Y(n4256));
  XOR2X1  g3583(.A(n3972), .B(n3971), .Y(n4257));
  NAND3X1 g3584(.A(n4257), .B(n4181), .C(n4178), .Y(n4258));
  OAI21X1 g3585(.A0(n4257), .A1(n4256), .B0(n4258), .Y(n4260));
  NAND4X1 g3586(.A(n4054), .B(n4049), .C(n768), .D(n4260), .Y(n4261));
  NAND2X1 g3587(.A(n4063), .B(REG3_REG_2__SCAN_IN), .Y(n4262));
  AOI22X1 g3588(.A0(n4056), .A1(REG3_REG_2__SCAN_IN), .B0(n957), .B1(n4067), .Y(n4263));
  OAI21X1 g3589(.A0(n4240), .A1(n1057), .B0(n4263), .Y(n4264));
  OAI22X1 g3590(.A0(n1026), .A1(n4071), .B0(n1032), .B1(STATE_REG_SCAN_IN), .Y(n4265));
  AOI21X1 g3591(.A0(n4264), .A1(n4064), .B0(n4265), .Y(n4266));
  NAND3X1 g3592(.A(n4266), .B(n4262), .C(n4261), .Y(U3234));
  NOR2X1  g3593(.A(n4027), .B(n4025), .Y(n4268));
  AOI21X1 g3594(.A0(n4027), .A1(n4025), .B0(n4010), .Y(n4269));
  XOR2X1  g3595(.A(n4022), .B(n4019), .Y(n4270));
  NOR3X1  g3596(.A(n4270), .B(n4269), .C(n4268), .Y(n4271));
  AOI21X1 g3597(.A0(n4028), .A1(n4204), .B0(n4268), .Y(n4272));
  AOI21X1 g3598(.A0(n4036), .A1(n4024), .B0(n4272), .Y(n4273));
  OAI21X1 g3599(.A0(n4273), .A1(n4271), .B0(n4163), .Y(n4274));
  NAND2X1 g3600(.A(n4063), .B(n1500), .Y(n4275));
  AOI22X1 g3601(.A0(n4056), .A1(n1500), .B0(n1444), .B1(n4067), .Y(n4276));
  OAI21X1 g3602(.A0(n4240), .A1(n1547), .B0(n4276), .Y(n4277));
  OAI22X1 g3603(.A0(n1507), .A1(n4071), .B0(n1485), .B1(STATE_REG_SCAN_IN), .Y(n4278));
  AOI21X1 g3604(.A0(n4277), .A1(n4064), .B0(n4278), .Y(n4279));
  NAND3X1 g3605(.A(n4279), .B(n4275), .C(n4274), .Y(U3233));
  XOR2X1  g3606(.A(n4098), .B(n4096), .Y(n4281));
  XOR2X1  g3607(.A(n4281), .B(n4151), .Y(n4282));
  INVX1   g3608(.A(n2005), .Y(n4283));
  OAI22X1 g3609(.A0(n4049), .A1(n4283), .B0(n1965), .B1(n4068), .Y(n4284));
  AOI21X1 g3610(.A0(n4066), .A1(n2071), .B0(n4284), .Y(n4285));
  AOI22X1 g3611(.A0(n2017), .A1(n4072), .B0(REG3_REG_22__SCAN_IN), .B1(U3149), .Y(n4286));
  OAI21X1 g3612(.A0(n4285), .A1(n4065), .B0(n4286), .Y(n4287));
  AOI21X1 g3613(.A0(n4063), .A1(n2005), .B0(n4287), .Y(n4288));
  OAI21X1 g3614(.A0(n4282), .A1(n4055), .B0(n4288), .Y(U3232));
  NAND2X1 g3615(.A(n4038), .B(n4037), .Y(n4290));
  OAI21X1 g3616(.A0(n4272), .A1(n4023), .B0(n4036), .Y(n4291));
  INVX1   g3617(.A(n4291), .Y(n4292));
  OAI21X1 g3618(.A0(n4016), .A1(n4015), .B0(n4017), .Y(n4293));
  AOI21X1 g3619(.A0(n4292), .A1(n4290), .B0(n4293), .Y(n4294));
  AOI21X1 g3620(.A0(n4013), .A1(n4012), .B0(n4292), .Y(n4295));
  AOI22X1 g3621(.A0(n4030), .A1(n4016), .B0(n4038), .B1(n4037), .Y(n4296));
  OAI21X1 g3622(.A0(n4016), .A1(n4030), .B0(n4296), .Y(n4297));
  OAI21X1 g3623(.A0(n4297), .A1(n4295), .B0(n4163), .Y(n4298));
  NOR2X1  g3624(.A(n4240), .B(n1645), .Y(n4299));
  OAI22X1 g3625(.A0(n4049), .A1(n1591), .B0(n1547), .B1(n4068), .Y(n4300));
  OAI21X1 g3626(.A0(n4300), .A1(n4299), .B0(n4064), .Y(n4301));
  AOI22X1 g3627(.A0(n1620), .A1(n4072), .B0(REG3_REG_13__SCAN_IN), .B1(U3149), .Y(n4302));
  NAND2X1 g3628(.A(n4302), .B(n4301), .Y(n4303));
  AOI21X1 g3629(.A0(n4063), .A1(n1592), .B0(n4303), .Y(n4304));
  OAI21X1 g3630(.A0(n4298), .A1(n4294), .B0(n4304), .Y(U3231));
  INVX1   g3631(.A(n4115), .Y(n4306));
  XOR2X1  g3632(.A(n4117), .B(n4306), .Y(n4307));
  NAND2X1 g3633(.A(n4112), .B(n4110), .Y(n4308));
  AOI21X1 g3634(.A0(n4308), .A1(n4149), .B0(n4113), .Y(n4309));
  INVX1   g3635(.A(n4309), .Y(n4310));
  INVX1   g3636(.A(n4117), .Y(n4311));
  NOR2X1  g3637(.A(n4311), .B(n4306), .Y(n4312));
  OAI21X1 g3638(.A0(n4120), .A1(n4312), .B0(n4310), .Y(n4313));
  OAI21X1 g3639(.A0(n4310), .A1(n4307), .B0(n4313), .Y(n4314));
  NAND2X1 g3640(.A(n4314), .B(n4163), .Y(n4315));
  NAND3X1 g3641(.A(n4221), .B(n1921), .C(STATE_REG_SCAN_IN), .Y(n4316));
  AOI22X1 g3642(.A0(n4056), .A1(n1921), .B0(n1884), .B1(n4067), .Y(n4317));
  OAI21X1 g3643(.A0(n4240), .A1(n1965), .B0(n4317), .Y(n4318));
  OAI22X1 g3644(.A0(n1941), .A1(n4071), .B0(n1958), .B1(STATE_REG_SCAN_IN), .Y(n4319));
  AOI21X1 g3645(.A0(n4318), .A1(n4064), .B0(n4319), .Y(n4320));
  NAND3X1 g3646(.A(n4320), .B(n4316), .C(n4315), .Y(U3230));
  OAI21X1 g3647(.A0(n4064), .A1(n4057), .B0(n4056), .Y(n4322));
  OAI21X1 g3648(.A0(n4060), .A1(U3149), .B0(n4322), .Y(n4323));
  NAND2X1 g3649(.A(n4323), .B(REG3_REG_0__SCAN_IN), .Y(n4324));
  NAND4X1 g3650(.A(n4049), .B(n3160), .C(n768), .D(n4054), .Y(n4325));
  NAND3X1 g3651(.A(n4066), .B(n4064), .C(n957), .Y(n4326));
  OAI21X1 g3652(.A0(n922), .A1(STATE_REG_SCAN_IN), .B0(n4326), .Y(n4327));
  AOI21X1 g3653(.A0(n4072), .A1(n909), .B0(n4327), .Y(n4328));
  NAND3X1 g3654(.A(n4328), .B(n4325), .C(n4324), .Y(U3229));
  NAND2X1 g3655(.A(n4004), .B(n3996), .Y(n4330));
  XOR2X1  g3656(.A(n4007), .B(n4170), .Y(n4331));
  XOR2X1  g3657(.A(n4331), .B(n4330), .Y(n4332));
  OAI22X1 g3658(.A0(n4049), .A1(n1381), .B0(n1339), .B1(n4068), .Y(n4333));
  AOI21X1 g3659(.A0(n4066), .A1(n1444), .B0(n4333), .Y(n4334));
  AOI22X1 g3660(.A0(n1451), .A1(n4072), .B0(REG3_REG_9__SCAN_IN), .B1(U3149), .Y(n4335));
  OAI21X1 g3661(.A0(n4334), .A1(n4065), .B0(n4335), .Y(n4336));
  AOI21X1 g3662(.A0(n4063), .A1(n2600), .B0(n4336), .Y(n4337));
  OAI21X1 g3663(.A0(n4332), .A1(n4055), .B0(n4337), .Y(U3228));
  NOR2X1  g3664(.A(n4184), .B(n4182), .Y(n4339));
  XOR2X1  g3665(.A(n4171), .B(n3946), .Y(n4340));
  XOR2X1  g3666(.A(n4340), .B(n4339), .Y(n4341));
  NOR2X1  g3667(.A(n4240), .B(n1167), .Y(n4342));
  OAI22X1 g3668(.A0(n4049), .A1(n1107), .B0(n1057), .B1(n4068), .Y(n4343));
  OAI21X1 g3669(.A0(n4343), .A1(n4342), .B0(n4064), .Y(n4344));
  AOI22X1 g3670(.A0(n1135), .A1(n4072), .B0(REG3_REG_4__SCAN_IN), .B1(U3149), .Y(n4345));
  NAND2X1 g3671(.A(n4345), .B(n4344), .Y(n4346));
  AOI21X1 g3672(.A0(n4063), .A1(n1120), .B0(n4346), .Y(n4347));
  OAI21X1 g3673(.A0(n4341), .A1(n4055), .B0(n4347), .Y(U3227));
  INVX1   g3674(.A(n4084), .Y(n4349));
  XOR2X1  g3675(.A(n4086), .B(n4349), .Y(n4350));
  NOR2X1  g3676(.A(n4350), .B(n4215), .Y(n4351));
  AOI21X1 g3677(.A0(n4089), .A1(n4088), .B0(n4153), .Y(n4352));
  OAI21X1 g3678(.A0(n4352), .A1(n4351), .B0(n4163), .Y(n4353));
  NAND3X1 g3679(.A(n4221), .B(n2114), .C(STATE_REG_SCAN_IN), .Y(n4354));
  AOI22X1 g3680(.A0(n4056), .A1(n2114), .B0(n2071), .B1(n4067), .Y(n4355));
  OAI21X1 g3681(.A0(n4240), .A1(n2170), .B0(n4355), .Y(n4356));
  OAI22X1 g3682(.A0(n2156), .A1(n4071), .B0(n2112), .B1(STATE_REG_SCAN_IN), .Y(n4357));
  AOI21X1 g3683(.A0(n4356), .A1(n4064), .B0(n4357), .Y(n4358));
  NAND3X1 g3684(.A(n4358), .B(n4354), .C(n4353), .Y(U3226));
  OAI21X1 g3685(.A0(n4135), .A1(n4133), .B0(n4136), .Y(n4360));
  AOI21X1 g3686(.A0(n4144), .A1(n4209), .B0(n4360), .Y(n4361));
  INVX1   g3687(.A(n4130), .Y(n4362));
  INVX1   g3688(.A(n4132), .Y(n4363));
  NOR2X1  g3689(.A(n4363), .B(n4362), .Y(n4364));
  OAI22X1 g3690(.A0(n4142), .A1(n4135), .B0(n4132), .B1(n4130), .Y(n4365));
  AOI21X1 g3691(.A0(n4135), .A1(n4142), .B0(n4365), .Y(n4366));
  OAI21X1 g3692(.A0(n4209), .A1(n4364), .B0(n4366), .Y(n4367));
  NAND2X1 g3693(.A(n4367), .B(n4163), .Y(n4368));
  NOR2X1  g3694(.A(n4240), .B(n1838), .Y(n4369));
  OAI22X1 g3695(.A0(n4049), .A1(n1786), .B0(n1737), .B1(n4068), .Y(n4370));
  OAI21X1 g3696(.A0(n4370), .A1(n4369), .B0(n4064), .Y(n4371));
  AOI22X1 g3697(.A0(n1828), .A1(n4072), .B0(REG3_REG_17__SCAN_IN), .B1(U3149), .Y(n4372));
  NAND2X1 g3698(.A(n4372), .B(n4371), .Y(n4373));
  AOI21X1 g3699(.A0(n4063), .A1(n2659), .B0(n4373), .Y(n4374));
  OAI21X1 g3700(.A0(n4368), .A1(n4361), .B0(n4374), .Y(U3225));
  XOR2X1  g3701(.A(n3992), .B(n3990), .Y(n4376));
  XOR2X1  g3702(.A(n4376), .B(n4234), .Y(n4377));
  NAND2X1 g3703(.A(n4066), .B(n1218), .Y(n4378));
  AOI22X1 g3704(.A0(n4056), .A1(n1194), .B0(n1122), .B1(n4067), .Y(n4379));
  AOI21X1 g3705(.A0(n4379), .A1(n4378), .B0(n4065), .Y(n4380));
  AOI22X1 g3706(.A0(n1178), .A1(n4072), .B0(REG3_REG_5__SCAN_IN), .B1(U3149), .Y(n4381));
  OAI21X1 g3707(.A0(n4062), .A1(n1165), .B0(n4381), .Y(n4382));
  NOR2X1  g3708(.A(n4382), .B(n4380), .Y(n4383));
  OAI21X1 g3709(.A0(n4377), .A1(n4055), .B0(n4383), .Y(U3224));
  XOR2X1  g3710(.A(n4132), .B(n4362), .Y(n4385));
  OAI21X1 g3711(.A0(n4143), .A1(n4364), .B0(n4141), .Y(n4386));
  OAI21X1 g3712(.A0(n4385), .A1(n4141), .B0(n4386), .Y(n4387));
  NAND2X1 g3713(.A(n4387), .B(n4163), .Y(n4388));
  NAND2X1 g3714(.A(n4063), .B(n2651), .Y(n4389));
  AOI22X1 g3715(.A0(n4056), .A1(n2651), .B0(n1689), .B1(n4067), .Y(n4390));
  OAI21X1 g3716(.A0(n4240), .A1(n1790), .B0(n4390), .Y(n4391));
  OAI22X1 g3717(.A0(n1751), .A1(n4071), .B0(n1730), .B1(STATE_REG_SCAN_IN), .Y(n4392));
  AOI21X1 g3718(.A0(n4391), .A1(n4064), .B0(n4392), .Y(n4393));
  NAND3X1 g3719(.A(n4393), .B(n4389), .C(n4388), .Y(U3223));
  XOR2X1  g3720(.A(n4081), .B(n4078), .Y(n4395));
  NOR2X1  g3721(.A(n4395), .B(n4154), .Y(n4396));
  AOI21X1 g3722(.A0(n4215), .A1(n4089), .B0(n4087), .Y(n4397));
  XOR2X1  g3723(.A(n4080), .B(n4078), .Y(n4398));
  NOR2X1  g3724(.A(n4398), .B(n4397), .Y(n4399));
  OAI21X1 g3725(.A0(n4399), .A1(n4396), .B0(n4163), .Y(n4400));
  NAND3X1 g3726(.A(n4221), .B(n2165), .C(STATE_REG_SCAN_IN), .Y(n4401));
  AOI22X1 g3727(.A0(n4056), .A1(n2165), .B0(n2181), .B1(n4067), .Y(n4402));
  OAI21X1 g3728(.A0(n4240), .A1(n2283), .B0(n4402), .Y(n4403));
  OAI22X1 g3729(.A0(n2186), .A1(n4071), .B0(n2162), .B1(STATE_REG_SCAN_IN), .Y(n4404));
  AOI21X1 g3730(.A0(n4403), .A1(n4064), .B0(n4404), .Y(n4405));
  NAND3X1 g3731(.A(n4405), .B(n4401), .C(n4400), .Y(U3222));
  XOR2X1  g3732(.A(n4038), .B(n4012), .Y(n4407));
  NAND2X1 g3733(.A(n4407), .B(n4291), .Y(n4409));
  OAI21X1 g3734(.A0(n4407), .A1(n4291), .B0(n4409), .Y(n4410));
  NAND2X1 g3735(.A(n4410), .B(n4163), .Y(n4411));
  NAND2X1 g3736(.A(n4063), .B(n1565), .Y(n4412));
  AOI22X1 g3737(.A0(n4056), .A1(n1565), .B0(n1502), .B1(n4067), .Y(n4413));
  OAI21X1 g3738(.A0(n4240), .A1(n1595), .B0(n4413), .Y(n4414));
  OAI22X1 g3739(.A0(n1588), .A1(n4071), .B0(n1640), .B1(STATE_REG_SCAN_IN), .Y(n4415));
  AOI21X1 g3740(.A0(n4414), .A1(n4064), .B0(n4415), .Y(n4416));
  NAND3X1 g3741(.A(n4416), .B(n4412), .C(n4411), .Y(U3221));
  AOI21X1 g3742(.A0(n4107), .A1(n4105), .B0(n4119), .Y(n4418));
  OAI21X1 g3743(.A0(n4310), .A1(n4120), .B0(n4418), .Y(n4419));
  OAI22X1 g3744(.A0(n4115), .A1(n4117), .B0(n4107), .B1(n4104), .Y(n4420));
  AOI21X1 g3745(.A0(n4107), .A1(n4104), .B0(n4420), .Y(n4421));
  OAI21X1 g3746(.A0(n4309), .A1(n4312), .B0(n4421), .Y(n4422));
  NAND3X1 g3747(.A(n4422), .B(n4419), .C(n4163), .Y(n4423));
  NAND3X1 g3748(.A(n4221), .B(n1960), .C(STATE_REG_SCAN_IN), .Y(n4424));
  AOI22X1 g3749(.A0(n4056), .A1(n1960), .B0(n1925), .B1(n4067), .Y(n4425));
  OAI21X1 g3750(.A0(n4240), .A1(n2009), .B0(n4425), .Y(n4426));
  NAND2X1 g3751(.A(n4426), .B(n4064), .Y(n4427));
  AOI22X1 g3752(.A0(n1973), .A1(n4072), .B0(REG3_REG_21__SCAN_IN), .B1(U3149), .Y(n4428));
  NAND4X1 g3753(.A(n4427), .B(n4424), .C(n4423), .D(n4428), .Y(U3220));
  NOR2X1  g3754(.A(n4179), .B(n4177), .Y(n4430));
  XOR2X1  g3755(.A(n4175), .B(n3957), .Y(n4431));
  XOR2X1  g3756(.A(n4431), .B(n4430), .Y(n4432));
  NAND4X1 g3757(.A(n4054), .B(n4049), .C(n768), .D(n4432), .Y(n4433));
  NAND2X1 g3758(.A(n4063), .B(REG3_REG_1__SCAN_IN), .Y(n4434));
  AOI22X1 g3759(.A0(n4056), .A1(REG3_REG_1__SCAN_IN), .B0(n986), .B1(n4067), .Y(n4435));
  OAI21X1 g3760(.A0(n4240), .A1(n1034), .B0(n4435), .Y(n4436));
  OAI22X1 g3761(.A0(n998), .A1(n4071), .B0(n1017), .B1(STATE_REG_SCAN_IN), .Y(n4437));
  AOI21X1 g3762(.A0(n4436), .A1(n4064), .B0(n4437), .Y(n4438));
  NAND3X1 g3763(.A(n4438), .B(n4434), .C(n4433), .Y(U3219));
  OAI21X1 g3764(.A0(n3994), .A1(n4234), .B0(n4197), .Y(n4440));
  XOR2X1  g3765(.A(n3980), .B(n3979), .Y(n4441));
  XOR2X1  g3766(.A(n4441), .B(n4440), .Y(n4442));
  OAI22X1 g3767(.A0(n4049), .A1(n1337), .B0(n1298), .B1(n4068), .Y(n4443));
  AOI21X1 g3768(.A0(n4066), .A1(n1392), .B0(n4443), .Y(n4444));
  AOI22X1 g3769(.A0(n1354), .A1(n4072), .B0(REG3_REG_8__SCAN_IN), .B1(U3149), .Y(n4445));
  OAI21X1 g3770(.A0(n4444), .A1(n4065), .B0(n4445), .Y(n4446));
  AOI21X1 g3771(.A0(n4063), .A1(n2590), .B0(n4446), .Y(n4447));
  OAI21X1 g3772(.A0(n4442), .A1(n4055), .B0(n4447), .Y(U3218));
  AOI22X1 g3773(.A0(n3145), .A1(n2342), .B0(n2287), .B1(n3156), .Y(n4449));
  OAI22X1 g3774(.A0(n3146), .A1(n2276), .B0(n2323), .B1(n3155), .Y(n4450));
  XOR2X1  g3775(.A(n4450), .B(n3152), .Y(n4451));
  NAND2X1 g3776(.A(n4451), .B(n4449), .Y(n4452));
  NAND2X1 g3777(.A(n4218), .B(n4087), .Y(n4453));
  NOR2X1  g3778(.A(n4157), .B(n4155), .Y(n4454));
  NOR2X1  g3779(.A(n4454), .B(n4159), .Y(n4455));
  AOI22X1 g3780(.A0(n4453), .A1(n4455), .B0(n4157), .B1(n4155), .Y(n4456));
  INVX1   g3781(.A(n4456), .Y(n4457));
  NAND2X1 g3782(.A(n4218), .B(n4089), .Y(n4458));
  OAI21X1 g3783(.A0(n4458), .A1(n4153), .B0(n4457), .Y(n4459));
  OAI22X1 g3784(.A0(n3958), .A1(n2331), .B0(n2374), .B1(n3146), .Y(n4460));
  XOR2X1  g3785(.A(n4460), .B(n3152), .Y(n4461));
  OAI22X1 g3786(.A0(n3146), .A1(n2331), .B0(n2374), .B1(n3155), .Y(n4462));
  XOR2X1  g3787(.A(n4462), .B(n4461), .Y(n4463));
  INVX1   g3788(.A(n4463), .Y(n4464));
  OAI21X1 g3789(.A0(n4451), .A1(n4449), .B0(n4464), .Y(n4465));
  AOI21X1 g3790(.A0(n4459), .A1(n4452), .B0(n4465), .Y(n4466));
  NAND3X1 g3791(.A(n4218), .B(n4215), .C(n4089), .Y(n4467));
  NOR2X1  g3792(.A(n4451), .B(n4449), .Y(n4468));
  NOR2X1  g3793(.A(n4468), .B(n4456), .Y(n4469));
  NAND2X1 g3794(.A(n4463), .B(n4452), .Y(n4470));
  AOI21X1 g3795(.A0(n4469), .A1(n4467), .B0(n4470), .Y(n4471));
  OAI21X1 g3796(.A0(n4471), .A1(n4466), .B0(n4163), .Y(n4472));
  NAND3X1 g3797(.A(n4221), .B(n2326), .C(STATE_REG_SCAN_IN), .Y(n4473));
  NOR2X1  g3798(.A(n4240), .B(n2381), .Y(n4474));
  OAI22X1 g3799(.A0(n4049), .A1(n2325), .B0(n2276), .B1(n4068), .Y(n4475));
  OAI21X1 g3800(.A0(n4475), .A1(n4474), .B0(n4064), .Y(n4476));
  AOI22X1 g3801(.A0(n2339), .A1(n4072), .B0(REG3_REG_28__SCAN_IN), .B1(U3149), .Y(n4477));
  NAND4X1 g3802(.A(n4476), .B(n4473), .C(n4472), .D(n4477), .Y(U3217));
  INVX1   g3803(.A(n4110), .Y(n4479));
  XOR2X1  g3804(.A(n4112), .B(n4479), .Y(n4480));
  NOR2X1  g3805(.A(n4480), .B(n4149), .Y(n4481));
  AOI21X1 g3806(.A0(n4308), .A1(n4114), .B0(n4211), .Y(n4482));
  OAI21X1 g3807(.A0(n4482), .A1(n4481), .B0(n4163), .Y(n4483));
  NAND2X1 g3808(.A(n4063), .B(n1882), .Y(n4484));
  AOI22X1 g3809(.A0(n4056), .A1(n1882), .B0(n1837), .B1(n4067), .Y(n4485));
  OAI21X1 g3810(.A0(n4240), .A1(n1926), .B0(n4485), .Y(n4486));
  OAI22X1 g3811(.A0(n1897), .A1(n4071), .B0(n1878), .B1(STATE_REG_SCAN_IN), .Y(n4487));
  AOI21X1 g3812(.A0(n4486), .A1(n4064), .B0(n4487), .Y(n4488));
  NAND3X1 g3813(.A(n4488), .B(n4484), .C(n4483), .Y(U3216));
  OAI21X1 g3814(.A0(n3954), .A1(n3952), .B0(n3955), .Y(n4490));
  AOI21X1 g3815(.A0(n3973), .A1(n4256), .B0(n4490), .Y(n4491));
  AOI22X1 g3816(.A0(n4178), .A1(n4181), .B0(n3951), .B1(n3949), .Y(n4492));
  AOI22X1 g3817(.A0(n3952), .A1(n4172), .B0(n3972), .B1(n3971), .Y(n4493));
  OAI21X1 g3818(.A0(n4172), .A1(n3952), .B0(n4493), .Y(n4494));
  OAI21X1 g3819(.A0(n4494), .A1(n4492), .B0(n4163), .Y(n4495));
  OAI22X1 g3820(.A0(n4049), .A1(REG3_REG_3__SCAN_IN), .B0(n1034), .B1(n4068), .Y(n4496));
  AOI21X1 g3821(.A0(n4066), .A1(n1122), .B0(n4496), .Y(n4497));
  AOI22X1 g3822(.A0(n1073), .A1(n4072), .B0(REG3_REG_3__SCAN_IN), .B1(U3149), .Y(n4498));
  OAI21X1 g3823(.A0(n4497), .A1(n4065), .B0(n4498), .Y(n4499));
  AOI21X1 g3824(.A0(n4063), .A1(n1077), .B0(n4499), .Y(n4500));
  OAI21X1 g3825(.A0(n4495), .A1(n4491), .B0(n4500), .Y(U3215));
  XOR2X1  g3826(.A(n4027), .B(n4025), .Y(n4502));
  XOR2X1  g3827(.A(n4502), .B(n4010), .Y(n4503));
  OAI22X1 g3828(.A0(n4049), .A1(n1432), .B0(n1383), .B1(n4068), .Y(n4504));
  AOI21X1 g3829(.A0(n4066), .A1(n1502), .B0(n4504), .Y(n4505));
  AOI22X1 g3830(.A0(n1461), .A1(n4072), .B0(REG3_REG_10__SCAN_IN), .B1(U3149), .Y(n4506));
  OAI21X1 g3831(.A0(n4505), .A1(n4065), .B0(n4506), .Y(n4507));
  AOI21X1 g3832(.A0(n4063), .A1(n1442), .B0(n4507), .Y(n4508));
  OAI21X1 g3833(.A0(n4503), .A1(n4055), .B0(n4508), .Y(U3214));
  XOR2X1  g3834(.A(n4093), .B(n4091), .Y(n4510));
  XOR2X1  g3835(.A(n4510), .B(n4214), .Y(n4511));
  INVX1   g3836(.A(n2052), .Y(n4512));
  OAI22X1 g3837(.A0(n4049), .A1(n4512), .B0(n2009), .B1(n4068), .Y(n4513));
  AOI21X1 g3838(.A0(n4066), .A1(n2181), .B0(n4513), .Y(n4514));
  AOI22X1 g3839(.A0(n2066), .A1(n4072), .B0(REG3_REG_23__SCAN_IN), .B1(U3149), .Y(n4515));
  OAI21X1 g3840(.A0(n4514), .A1(n4065), .B0(n4515), .Y(n4516));
  AOI21X1 g3841(.A0(n4063), .A1(n2052), .B0(n4516), .Y(n4517));
  OAI21X1 g3842(.A0(n4511), .A1(n4055), .B0(n4517), .Y(U3213));
  XOR2X1  g3843(.A(n3939), .B(n3937), .Y(n4519));
  XOR2X1  g3844(.A(n4519), .B(n4207), .Y(n4520));
  OAI22X1 g3845(.A0(n4049), .A1(n1643), .B0(n1595), .B1(n4068), .Y(n4521));
  AOI21X1 g3846(.A0(n4066), .A1(n1689), .B0(n4521), .Y(n4522));
  AOI22X1 g3847(.A0(n1662), .A1(n4072), .B0(REG3_REG_14__SCAN_IN), .B1(U3149), .Y(n4523));
  OAI21X1 g3848(.A0(n4522), .A1(n4065), .B0(n4523), .Y(n4524));
  AOI21X1 g3849(.A0(n4063), .A1(n2637), .B0(n4524), .Y(n4525));
  OAI21X1 g3850(.A0(n4520), .A1(n4055), .B0(n4525), .Y(U3212));
  INVX1   g3851(.A(n4449), .Y(n4527));
  XOR2X1  g3852(.A(n4451), .B(n4527), .Y(n4528));
  XOR2X1  g3853(.A(n4528), .B(n4459), .Y(n4529));
  OAI22X1 g3854(.A0(n4049), .A1(n2270), .B0(n2283), .B1(n4068), .Y(n4530));
  AOI21X1 g3855(.A0(n4066), .A1(n2393), .B0(n4530), .Y(n4531));
  AOI22X1 g3856(.A0(n2287), .A1(n4072), .B0(REG3_REG_27__SCAN_IN), .B1(U3149), .Y(n4532));
  OAI21X1 g3857(.A0(n4531), .A1(n4065), .B0(n4532), .Y(n4533));
  AOI21X1 g3858(.A0(n4063), .A1(n2271), .B0(n4533), .Y(n4534));
  OAI21X1 g3859(.A0(n4529), .A1(n4055), .B0(n4534), .Y(U3211));
  OAI21X1 g3860(.A0(n3988), .A1(n3986), .B0(n3989), .Y(n4536));
  AOI21X1 g3861(.A0(n4236), .A1(n4193), .B0(n4536), .Y(n4537));
  NOR2X1  g3862(.A(n4188), .B(n4187), .Y(n4538));
  OAI22X1 g3863(.A0(n3997), .A1(n3988), .B0(n3985), .B1(n3983), .Y(n4539));
  AOI21X1 g3864(.A0(n3988), .A1(n3997), .B0(n4539), .Y(n4540));
  OAI21X1 g3865(.A0(n4236), .A1(n4538), .B0(n4540), .Y(n4541));
  NAND2X1 g3866(.A(n4541), .B(n4163), .Y(n4542));
  OAI22X1 g3867(.A0(n4049), .A1(n1271), .B0(n1285), .B1(n4068), .Y(n4543));
  AOI21X1 g3868(.A0(n4066), .A1(n1340), .B0(n4543), .Y(n4544));
  AOI22X1 g3869(.A0(n1292), .A1(n4072), .B0(REG3_REG_7__SCAN_IN), .B1(U3149), .Y(n4545));
  OAI21X1 g3870(.A0(n4544), .A1(n4065), .B0(n4545), .Y(n4546));
  AOI21X1 g3871(.A0(n4063), .A1(n1272), .B0(n4546), .Y(n4547));
  OAI21X1 g3872(.A0(n4542), .A1(n4537), .B0(n4547), .Y(U3210));
endmodule


