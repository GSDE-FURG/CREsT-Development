//Converted to Combinational (Partial output: n466) , Module name: s9234_n466 , Timestamp: 2018-12-03T15:51:03.421391 
module s9234_n466 ( g1, g2, g6, g28, g693, g698, g197, g687, g688, g684, g685, g269, g677, g689, g683, g702, g699, g41, g676, g662, g471, g211, g210, g207, g682, g678, g282, g283, g478, g279, g658, g206, g204, g205, g679, g266, g680, g554, g297, g561, g512, g449, g541, g414, g278, g276, g277, g48, g208, g209, g681, g280, g281, g10, g18, g14, g24, n466 );
input g1, g2, g6, g28, g693, g698, g197, g687, g688, g684, g685, g269, g677, g689, g683, g702, g699, g41, g676, g662, g471, g211, g210, g207, g682, g678, g282, g283, g478, g279, g658, g206, g204, g205, g679, g266, g680, g554, g297, g561, g512, g449, g541, g414, g278, g276, g277, g48, g208, g209, g681, g280, g281, g10, g18, g14, g24;
output n466;
wire n1363, n1207, n1354, n1362, n1361, n775, n166, n1186_1, n1185, n1188, n1206, n1353, n1178, n770, n1187, n821, n1359, n1360, n769, n758, n757, n843, n976_1, n974, n809, n943, n1184, n1205, n1197, n1198, n1201_1, n1352, n1208, n941_1, n1357, n1356, n765, n762, n725, n727, n761_1, n975, n972, n973, n792, n1182, n1183, n1203, n1204, n1196_1, n1191_1, n1193, n1194, n1180, n1009, n1200, n1345, n1348, n1351, n940, n920, n1073, n1355, n724, n726_1, n760, n970, n964, n971_1, n963, n1181_1, n1008, n1202, n1195, n1179, n1190, n1192, n802, n1189, n1005, n1006_1, n1199, n1343, n1344, n1347, n1346, n1349, n1350, n939, n911_1, n871_1, n922, n869, n716_1, n723, n968, n969, n960, n961_1, n962, n965, n966_1, n967, n795, n789, n798, n826_1, n813, n805, n906_1, n910, n870, n904, n905, n872, n719, n722, n866_1, n867, n868, n717, n718, n720, n721_1;
NAND4X1  g0655(.A(n1362), .B(n1354), .C(n1207), .D(n1363), .Y(n466));
AOI22X1  g0654(.A0(n1186_1), .A1(n166), .B0(n775), .B1(n1361), .Y(n1363));
NAND3X1  g0498(.A(n1206), .B(n1188), .C(n1185), .Y(n1207));
AOI21X1  g0645(.A0(n1178), .A1(g693), .B0(n1353), .Y(n1354));
AOI22X1  g0653(.A0(n821), .A1(n1187), .B0(n770), .B1(n1361), .Y(n1362));
NAND2X1  g0652(.A(n1360), .B(n1359), .Y(n1361));
NOR4X1   g0067(.A(n757), .B(g698), .C(n758), .D(n769), .Y(n775));
OAI22X1  g0268(.A0(n974), .A1(n976_1), .B0(g197), .B1(n843), .Y(n166));
NOR4X1   g0477(.A(n769), .B(g688), .C(g687), .D(n809), .Y(n1186_1));
NOR3X1   g0476(.A(n1184), .B(n1178), .C(n943), .Y(n1185));
NOR4X1   g0479(.A(n1186_1), .B(n775), .C(n770), .D(n1187), .Y(n1188));
NOR4X1   g0497(.A(n1201_1), .B(n1198), .C(n1197), .D(n1205), .Y(n1206));
OAI21X1  g0644(.A0(n1208), .A1(n843), .B0(n1352), .Y(n1353));
NOR4X1   g0469(.A(n769), .B(g685), .C(g684), .D(n941_1), .Y(n1178));
NOR4X1   g0062(.A(g687), .B(g698), .C(n758), .D(n769), .Y(n770));
NOR4X1   g0478(.A(n769), .B(g688), .C(n757), .D(n809), .Y(n1187));
OAI22X1  g0649(.A0(n1356), .A1(n1357), .B0(g269), .B1(n843), .Y(n821));
NAND2X1  g0650(.A(n765), .B(g693), .Y(n1359));
NAND2X1  g0651(.A(g677), .B(g693), .Y(n1360));
OR4X1    g0061(.A(n761_1), .B(n727), .C(n725), .D(n762), .Y(n769));
INVX1    g0050(.A(g689), .Y(n758));
INVX1    g0049(.A(g687), .Y(n757));
INVX1    g0135(.A(g693), .Y(n843));
NAND2X1  g0267(.A(n975), .B(g197), .Y(n976_1));
AND2X1   g0265(.A(n973), .B(n972), .Y(n974));
OR2X1    g0101(.A(g698), .B(g689), .Y(n809));
NOR4X1   g0234(.A(n769), .B(g685), .C(n792), .D(n941_1), .Y(n943));
NAND2X1  g0475(.A(n1183), .B(n1182), .Y(n1184));
NAND2X1  g0496(.A(n1204), .B(n1203), .Y(n1205));
OR4X1    g0488(.A(n1194), .B(n1193), .C(n1191_1), .D(n1196_1), .Y(n1197));
NOR4X1   g0489(.A(n1009), .B(g683), .C(n792), .D(n1180), .Y(n1198));
NOR3X1   g0492(.A(n1200), .B(n1180), .C(n1009), .Y(n1201_1));
NOR3X1   g0643(.A(n1351), .B(n1348), .C(n1345), .Y(n1352));
INVX1    g0499(.A(n943), .Y(n1208));
INVX1    g0232(.A(n940), .Y(n941_1));
NAND2X1  g0648(.A(n920), .B(g269), .Y(n1357));
AND2X1   g0647(.A(n1355), .B(n1073), .Y(n1356));
INVX1    g0057(.A(g677), .Y(n765));
NAND2X1  g0054(.A(g699), .B(g702), .Y(n762));
INVX1    g0017(.A(g41), .Y(n725));
OAI21X1  g0019(.A0(n726_1), .A1(n724), .B0(g676), .Y(n727));
NAND2X1  g0053(.A(n760), .B(g662), .Y(n761_1));
OR4X1    g0266(.A(g210), .B(g211), .C(g471), .D(n970), .Y(n975));
AND2X1   g0263(.A(n971_1), .B(n964), .Y(n972));
XOR2X1   g0264(.A(n963), .B(g207), .Y(n973));
INVX1    g0084(.A(g684), .Y(n792));
NAND4X1  g0473(.A(n1008), .B(n765), .C(g682), .D(n1181_1), .Y(n1182));
NAND4X1  g0474(.A(n1008), .B(g677), .C(g682), .D(n1181_1), .Y(n1183));
OR2X1    g0494(.A(n1202), .B(g677), .Y(n1203));
OR2X1    g0495(.A(n1202), .B(n765), .Y(n1204));
NOR4X1   g0487(.A(n1179), .B(n762), .C(n725), .D(n1195), .Y(n1196_1));
NOR4X1   g0482(.A(n1179), .B(n762), .C(n725), .D(n1190), .Y(n1191_1));
NOR4X1   g0484(.A(n1189), .B(n1180), .C(n802), .D(n1192), .Y(n1193));
NOR4X1   g0485(.A(n1189), .B(n1180), .C(g678), .D(n1192), .Y(n1194));
OR4X1    g0471(.A(n1006_1), .B(n725), .C(n1005), .D(n1179), .Y(n1180));
INVX1    g0300(.A(n1008), .Y(n1009));
INVX1    g0491(.A(n1199), .Y(n1200));
NAND2X1  g0636(.A(n1344), .B(n1343), .Y(n1345));
OAI22X1  g0639(.A0(n1182), .A1(n1346), .B0(n1347), .B1(n1204), .Y(n1348));
OAI22X1  g0642(.A0(n1183), .A1(n1350), .B0(n1349), .B1(n1203), .Y(n1351));
NOR3X1   g0231(.A(g688), .B(n939), .C(n758), .Y(n940));
OR4X1    g0212(.A(g478), .B(g283), .C(g282), .D(n911_1), .Y(n920));
AND2X1   g0364(.A(n922), .B(n871_1), .Y(n1073));
XOR2X1   g0646(.A(n869), .B(g279), .Y(n1355));
AND2X1   g0016(.A(n723), .B(n716_1), .Y(n724));
OAI21X1  g0018(.A0(n723), .A1(n716_1), .B0(n725), .Y(n726_1));
INVX1    g0052(.A(g658), .Y(n760));
NOR2X1   g0261(.A(n969), .B(n968), .Y(n970));
OR4X1    g0255(.A(n962), .B(n961_1), .C(n960), .D(n963), .Y(n964));
NAND4X1  g0262(.A(n967), .B(n966_1), .C(n965), .D(n970), .Y(n971_1));
NAND3X1  g0254(.A(g205), .B(g204), .C(g206), .Y(n963));
NOR3X1   g0472(.A(n1180), .B(n795), .C(n792), .Y(n1181_1));
NOR4X1   g0299(.A(n939), .B(n789), .C(n758), .D(g688), .Y(n1008));
NAND4X1  g0493(.A(n1008), .B(n826_1), .C(n798), .D(n1181_1), .Y(n1202));
OR4X1    g0486(.A(n813), .B(g679), .C(g678), .D(n1189), .Y(n1195));
OAI21X1  g0470(.A0(g266), .A1(g662), .B0(n760), .Y(n1179));
OR4X1    g0481(.A(g680), .B(n805), .C(n802), .D(n1189), .Y(n1190));
OR2X1    g0483(.A(g680), .B(g679), .Y(n1192));
INVX1    g0094(.A(g678), .Y(n802));
NAND3X1  g0480(.A(g688), .B(g698), .C(g689), .Y(n1189));
INVX1    g0296(.A(g702), .Y(n1005));
INVX1    g0297(.A(g699), .Y(n1006_1));
NOR4X1   g0490(.A(n826_1), .B(n792), .C(g682), .D(n795), .Y(n1199));
NAND2X1  g0634(.A(n1201_1), .B(g554), .Y(n1343));
AOI22X1  g0635(.A0(n1191_1), .A1(g561), .B0(g297), .B1(n1198), .Y(n1344));
INVX1    g0638(.A(g512), .Y(n1347));
INVX1    g0637(.A(g449), .Y(n1346));
INVX1    g0640(.A(g541), .Y(n1349));
INVX1    g0641(.A(g414), .Y(n1350));
INVX1    g0230(.A(g698), .Y(n939));
NOR2X1   g0203(.A(n910), .B(n906_1), .Y(n911_1));
INVX1    g0163(.A(n870), .Y(n871_1));
NAND4X1  g0214(.A(n872), .B(n905), .C(n904), .D(n911_1), .Y(n922));
NAND3X1  g0161(.A(g277), .B(g276), .C(g278), .Y(n869));
INVX1    g0008(.A(g48), .Y(n716_1));
XOR2X1   g0015(.A(n722), .B(n719), .Y(n723));
NOR4X1   g0259(.A(n962), .B(g208), .C(n960), .D(n963), .Y(n968));
XOR2X1   g0260(.A(g209), .B(n961_1), .Y(n969));
INVX1    g0251(.A(g207), .Y(n960));
INVX1    g0252(.A(g208), .Y(n961_1));
INVX1    g0253(.A(g209), .Y(n962));
INVX1    g0256(.A(g471), .Y(n965));
INVX1    g0257(.A(g211), .Y(n966_1));
INVX1    g0258(.A(g210), .Y(n967));
INVX1    g0087(.A(g683), .Y(n795));
INVX1    g0081(.A(g685), .Y(n789));
INVX1    g0090(.A(g682), .Y(n798));
INVX1    g0118(.A(g681), .Y(n826_1));
INVX1    g0105(.A(g680), .Y(n813));
INVX1    g0097(.A(g679), .Y(n805));
XOR2X1   g0198(.A(g280), .B(n866_1), .Y(n906_1));
NOR4X1   g0202(.A(g280), .B(n867), .C(n866_1), .D(n869), .Y(n910));
NOR4X1   g0162(.A(n868), .B(n867), .C(n866_1), .D(n869), .Y(n870));
INVX1    g0196(.A(g282), .Y(n904));
INVX1    g0197(.A(g283), .Y(n905));
INVX1    g0164(.A(g478), .Y(n872));
XOR2X1   g0011(.A(n718), .B(n717), .Y(n719));
XOR2X1   g0014(.A(n721_1), .B(n720), .Y(n722));
INVX1    g0158(.A(g281), .Y(n866_1));
INVX1    g0159(.A(g279), .Y(n867));
INVX1    g0160(.A(g280), .Y(n868));
XOR2X1   g0009(.A(g1), .B(g2), .Y(n717));
XOR2X1   g0010(.A(g10), .B(g6), .Y(n718));
XOR2X1   g0012(.A(g14), .B(g18), .Y(n720));
XOR2X1   g0013(.A(g28), .B(g24), .Y(n721_1));

endmodule
