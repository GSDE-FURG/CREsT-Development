//Converted to Combinational (Partial output: n4425) , Module name: s38417_n4425 , Timestamp: 2018-12-03T15:51:13.866436 
module s38417_n4425 ( g1421, g1211, g1224, g1309, g1345, g1414, g1416, g1418, g1415, g1315, g1312, g1352, g1346, g1326, g1417, g1419, g1378, g1339, g1358, g1372, g1365, g1332, g1394, g1319, g1388, g1412, g1411, g1413, g1391, g1390, g1392, g1400, g1399, g1401, g1403, g1402, g1404, g1409, g1408, g1410, g1406, g1405, g1407, g1397, g1396, g1398, g1385, g1384, g1386, g1393, g1395, g1387, g1389, n4425 );
input g1421, g1211, g1224, g1309, g1345, g1414, g1416, g1418, g1415, g1315, g1312, g1352, g1346, g1326, g1417, g1419, g1378, g1339, g1358, g1372, g1365, g1332, g1394, g1319, g1388, g1412, g1411, g1413, g1391, g1390, g1392, g1400, g1399, g1401, g1403, g1402, g1404, g1409, g1408, g1410, g1406, g1405, g1407, g1397, g1396, g1398, g1385, g1384, g1386, g1393, g1395, g1387, g1389;
output n4425;
wire n7254, n7351, n7212, n7350_1, n7344, n7348, n7349, n7215_1, n7298_1, n7343, n7314, n7324, n7334, n7347, n7296, n7338, n7342, n7313, n7301, n7305, n7309, n7319, n7323, n7328, n7333, n7346, n7345_1, n7284, n7337, n7223, n7341, n7236, n7312_1, n7300, n7247, n7304, n7243, n7308, n7227, n7318, n7322, n7327, n7219, n7332, n7335_1, n7336, n7339, n7340_1, n7310, n7311, n7297, n7299, n7302_1, n7303, n7306, n7307_1, n7317, n7320, n7321_1, n7325_1, n7326, n7331, n7316_1, n7315, n7330_1, n7329;
MX2X1    g2308(.A(n7351), .B(g1421), .S0(n7254), .Y(n4425));
NAND4X1  g2210(.A(g1309), .B(g1224), .C(g1211), .D(n7212), .Y(n7254));
NOR4X1   g2307(.A(n7349), .B(n7348), .C(n7344), .D(n7350_1), .Y(n7351));
INVX1    g2168(.A(g1345), .Y(n7212));
OAI22X1  g2306(.A0(g1416), .A1(n7298_1), .B0(n7215_1), .B1(g1414), .Y(n7350_1));
NOR4X1   g2300(.A(n7334), .B(n7324), .C(n7314), .D(n7343), .Y(n7344));
OAI21X1  g2304(.A0(g1418), .A1(n7296), .B0(n7347), .Y(n7348));
NOR2X1   g2305(.A(g1415), .B(n7296), .Y(n7349));
INVX1    g2171(.A(g1315), .Y(n7215_1));
INVX1    g2254(.A(g1312), .Y(n7298_1));
OR2X1    g2299(.A(n7342), .B(n7338), .Y(n7343));
OR4X1    g2270(.A(n7309), .B(n7305), .C(n7301), .D(n7313), .Y(n7314));
NAND2X1  g2280(.A(n7323), .B(n7319), .Y(n7324));
NAND2X1  g2290(.A(n7333), .B(n7328), .Y(n7334));
AOI22X1  g2303(.A0(n7345_1), .A1(g1312), .B0(g1315), .B1(n7346), .Y(n7347));
INVX1    g2252(.A(g1309), .Y(n7296));
XOR2X1   g2294(.A(n7337), .B(n7284), .Y(n7338));
XOR2X1   g2298(.A(n7341), .B(n7223), .Y(n7342));
XOR2X1   g2269(.A(n7312_1), .B(n7236), .Y(n7313));
XOR2X1   g2257(.A(n7300), .B(g1352), .Y(n7301));
XOR2X1   g2261(.A(n7304), .B(n7247), .Y(n7305));
XOR2X1   g2265(.A(n7308), .B(n7243), .Y(n7309));
XOR2X1   g2275(.A(n7318), .B(n7227), .Y(n7319));
XOR2X1   g2279(.A(n7322), .B(g1346), .Y(n7323));
XOR2X1   g2284(.A(n7327), .B(g1326), .Y(n7328));
XOR2X1   g2289(.A(n7332), .B(n7219), .Y(n7333));
INVX1    g2302(.A(g1417), .Y(n7346));
INVX1    g2301(.A(g1419), .Y(n7345_1));
INVX1    g2240(.A(g1378), .Y(n7284));
NOR2X1   g2293(.A(n7336), .B(n7335_1), .Y(n7337));
INVX1    g2179(.A(g1339), .Y(n7223));
NOR2X1   g2297(.A(n7340_1), .B(n7339), .Y(n7341));
INVX1    g2192(.A(g1358), .Y(n7236));
NOR2X1   g2268(.A(n7311), .B(n7310), .Y(n7312_1));
OR2X1    g2256(.A(n7299), .B(n7297), .Y(n7300));
INVX1    g2203(.A(g1372), .Y(n7247));
NOR2X1   g2260(.A(n7303), .B(n7302_1), .Y(n7304));
INVX1    g2199(.A(g1365), .Y(n7243));
NOR2X1   g2264(.A(n7307_1), .B(n7306), .Y(n7308));
INVX1    g2183(.A(g1332), .Y(n7227));
OAI21X1  g2274(.A0(g1394), .A1(n7296), .B0(n7317), .Y(n7318));
NOR2X1   g2278(.A(n7321_1), .B(n7320), .Y(n7322));
NOR2X1   g2283(.A(n7326), .B(n7325_1), .Y(n7327));
INVX1    g2175(.A(g1319), .Y(n7219));
OAI21X1  g2288(.A0(g1388), .A1(n7296), .B0(n7331), .Y(n7332));
NOR2X1   g2291(.A(g1412), .B(n7296), .Y(n7335_1));
OAI22X1  g2292(.A0(g1413), .A1(n7298_1), .B0(n7215_1), .B1(g1411), .Y(n7336));
NOR2X1   g2295(.A(g1391), .B(n7296), .Y(n7339));
OAI22X1  g2296(.A0(g1392), .A1(n7298_1), .B0(n7215_1), .B1(g1390), .Y(n7340_1));
NOR2X1   g2266(.A(g1400), .B(n7296), .Y(n7310));
OAI22X1  g2267(.A0(g1401), .A1(n7298_1), .B0(n7215_1), .B1(g1399), .Y(n7311));
NOR2X1   g2253(.A(g1403), .B(n7296), .Y(n7297));
OAI22X1  g2255(.A0(g1404), .A1(n7298_1), .B0(n7215_1), .B1(g1402), .Y(n7299));
NOR2X1   g2258(.A(g1409), .B(n7296), .Y(n7302_1));
OAI22X1  g2259(.A0(g1410), .A1(n7298_1), .B0(n7215_1), .B1(g1408), .Y(n7303));
NOR2X1   g2262(.A(g1406), .B(n7296), .Y(n7306));
OAI22X1  g2263(.A0(g1407), .A1(n7298_1), .B0(n7215_1), .B1(g1405), .Y(n7307_1));
AOI22X1  g2273(.A0(n7315), .A1(g1312), .B0(g1315), .B1(n7316_1), .Y(n7317));
NOR2X1   g2276(.A(g1397), .B(n7296), .Y(n7320));
OAI22X1  g2277(.A0(g1398), .A1(n7298_1), .B0(n7215_1), .B1(g1396), .Y(n7321_1));
NOR2X1   g2281(.A(g1385), .B(n7296), .Y(n7325_1));
OAI22X1  g2282(.A0(g1386), .A1(n7298_1), .B0(n7215_1), .B1(g1384), .Y(n7326));
AOI22X1  g2287(.A0(n7329), .A1(g1312), .B0(g1315), .B1(n7330_1), .Y(n7331));
INVX1    g2272(.A(g1393), .Y(n7316_1));
INVX1    g2271(.A(g1395), .Y(n7315));
INVX1    g2286(.A(g1387), .Y(n7330_1));
INVX1    g2285(.A(g1389), .Y(n7329));

endmodule
