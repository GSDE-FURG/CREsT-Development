//Converted to Combinational (Partial output: n161) , Module name: s9234_n161 , Timestamp: 2018-12-03T15:51:03.367424 
module s9234_n161 ( g1, g2, g6, g10, g24, g28, g102, g89, g94, g98, g658, g690, g123, g114, g260, g686, g662, g685, g650, g681, g646, g680, g642, g678, g606, g679, g139, g128, g131, g135, g684, g41, g571, g683, g654, g682, g254, g248, g236, g242, g688, g702, g699, g676, g297, g212, g283, g282, g689, g698, g218, g224, g288, g289, g287, g567, g598, g634, g478, g48, g687, g286, g284, g691, g697, g692, g694, g693, g695, g696, g278, g276, g277, g281, g279, g280, g292, g290, g285, g291, g18, g14, n161 );
input g1, g2, g6, g10, g24, g28, g102, g89, g94, g98, g658, g690, g123, g114, g260, g686, g662, g685, g650, g681, g646, g680, g642, g678, g606, g679, g139, g128, g131, g135, g684, g41, g571, g683, g654, g682, g254, g248, g236, g242, g688, g702, g699, g676, g297, g212, g283, g282, g689, g698, g218, g224, g288, g289, g287, g567, g598, g634, g478, g48, g687, g286, g284, g691, g697, g692, g694, g693, g695, g696, g278, g276, g277, g281, g279, g280, g292, g290, g285, g291, g18, g14;
output n161;
wire n788, n958, n787, n957, n830, n937, n786_1, n780, n784, n956_1, n944, n948, n953, n801_1, n829, n936_1, n785, n783, n955, n954, n767, n942, n943, n947, n949, n950, n952, n951_1, n791_1, n794, n800, n797, n825, n819, n822, n824, n865, n932, n935, n781_1, n782, n941_1, n792, n938, n769, n945, n946_1, n790, n789, n793, n799, n798, n796_1, n795, n820, n818, n823, n804, n815, n821_1, n864, n926_1, n931_1, n933, n934, n940, n762, n727, n761_1, n725, n816_1, n811_1, n817, n807, n803, n802, n814, n863, n842, n851_1, n905, n915, n918, n921_1, n927, n928, n930, n904, n924, n758, n939, n724, n726_1, n760, n810, n763, n806_1, n805, n813, n812, n862, n852, n853, n854, n841_1, n833, n837, n839, n850, n844, n846_1, n848, n871_1, n909, n914, n917, n919, n920, n870, n929, n922, n912, n923, n716_1, n723, n757, n808, n809, n855, n856_1, n861_1, n496, n916, n831_1, n836_1, n834, n835, n838, n849, n843, n845, n847, n908, n889, n903, n913, n916_1, n911_1, n869, n866_1, n867, n868, n872, n907, n719, n722, n860, n857, n858, n859, n887, n888, n901_1, n902, n906_1, n910, n717, n718, n720, n721_1, n886_1, n900, n874, n879, n885, n881_1, n891_1, n894, n899, n896_1, n873, n876_1, n878, n882, n883, n884, n880, n890, n892, n893, n897, n898, n895, n875, n877;
MX2X1    g0250(.A(n787), .B(n958), .S0(n788), .Y(n161));
NOR4X1   g0080(.A(g98), .B(g94), .C(g89), .D(g102), .Y(n788));
OAI21X1  g0249(.A0(n937), .A1(n830), .B0(n957), .Y(n958));
OAI21X1  g0079(.A0(n784), .A1(n780), .B0(n786_1), .Y(n787));
NOR4X1   g0248(.A(n953), .B(n948), .C(n944), .D(n956_1), .Y(n957));
AND2X1   g0122(.A(n829), .B(n801_1), .Y(n830));
MX2X1    g0228(.A(g690), .B(n936_1), .S0(g658), .Y(n937));
NAND3X1  g0078(.A(n784), .B(n785), .C(n780), .Y(n786_1));
INVX1    g0072(.A(g123), .Y(n780));
INVX1    g0076(.A(n783), .Y(n784));
MX2X1    g0247(.A(n954), .B(n955), .S0(g658), .Y(n956_1));
NOR3X1   g0235(.A(n943), .B(n942), .C(n767), .Y(n944));
NOR4X1   g0239(.A(n943), .B(n942), .C(n767), .D(n947), .Y(n948));
AOI22X1  g0244(.A0(n951_1), .A1(n952), .B0(n950), .B1(n949), .Y(n953));
OAI22X1  g0093(.A0(n797), .A1(n800), .B0(n794), .B1(n791_1), .Y(n801_1));
NAND4X1  g0121(.A(n824), .B(n822), .C(n819), .D(n825), .Y(n829));
NAND3X1  g0227(.A(n935), .B(n932), .C(n865), .Y(n936_1));
OR2X1    g0077(.A(g98), .B(g94), .Y(n785));
NAND3X1  g0075(.A(n782), .B(g114), .C(n781_1), .Y(n783));
INVX1    g0246(.A(g260), .Y(n955));
INVX1    g0245(.A(g686), .Y(n954));
AND2X1   g0059(.A(g658), .B(g662), .Y(n767));
NOR4X1   g0233(.A(n938), .B(g685), .C(n792), .D(n941_1), .Y(n942));
NOR4X1   g0234(.A(n769), .B(g685), .C(n792), .D(n941_1), .Y(n943));
AND2X1   g0238(.A(n946_1), .B(n945), .Y(n947));
MX2X1    g0240(.A(g681), .B(g650), .S0(g658), .Y(n949));
MX2X1    g0241(.A(g680), .B(g646), .S0(g658), .Y(n950));
MX2X1    g0243(.A(g678), .B(g642), .S0(g658), .Y(n952));
MX2X1    g0242(.A(g679), .B(g606), .S0(g658), .Y(n951_1));
MX2X1    g0083(.A(n789), .B(n790), .S0(g658), .Y(n791_1));
MX2X1    g0086(.A(n792), .B(n793), .S0(g658), .Y(n794));
MX2X1    g0092(.A(n798), .B(n799), .S0(g658), .Y(n800));
MX2X1    g0089(.A(n795), .B(n796_1), .S0(g658), .Y(n797));
OAI21X1  g0117(.A0(n823), .A1(n818), .B0(n820), .Y(n825));
OAI21X1  g0111(.A0(n818), .A1(n815), .B0(n804), .Y(n819));
OAI21X1  g0114(.A0(n821_1), .A1(n815), .B0(n820), .Y(n822));
OAI21X1  g0116(.A0(n823), .A1(n821_1), .B0(n804), .Y(n824));
INVX1    g0157(.A(n864), .Y(n865));
NAND2X1  g0223(.A(n931_1), .B(n926_1), .Y(n932));
NAND2X1  g0226(.A(n934), .B(n933), .Y(n935));
INVX1    g0073(.A(g139), .Y(n781_1));
NOR3X1   g0074(.A(g135), .B(g131), .C(g128), .Y(n782));
INVX1    g0232(.A(n940), .Y(n941_1));
INVX1    g0084(.A(g684), .Y(n792));
OR4X1    g0229(.A(n761_1), .B(n727), .C(g41), .D(n762), .Y(n938));
OR4X1    g0061(.A(n761_1), .B(n727), .C(n725), .D(n762), .Y(n769));
MX2X1    g0236(.A(g683), .B(g571), .S0(g658), .Y(n945));
MX2X1    g0237(.A(g682), .B(g654), .S0(g658), .Y(n946_1));
INVX1    g0082(.A(g254), .Y(n790));
INVX1    g0081(.A(g685), .Y(n789));
INVX1    g0085(.A(g248), .Y(n793));
INVX1    g0091(.A(g236), .Y(n799));
INVX1    g0090(.A(g682), .Y(n798));
INVX1    g0088(.A(g242), .Y(n796_1));
INVX1    g0087(.A(g683), .Y(n795));
INVX1    g0112(.A(n804), .Y(n820));
NOR3X1   g0110(.A(n817), .B(n811_1), .C(n816_1), .Y(n818));
NOR3X1   g0115(.A(n817), .B(n811_1), .C(n807), .Y(n823));
MX2X1    g0096(.A(n802), .B(n803), .S0(g658), .Y(n804));
NOR3X1   g0107(.A(n814), .B(n811_1), .C(n807), .Y(n815));
NOR3X1   g0113(.A(n814), .B(n811_1), .C(n816_1), .Y(n821_1));
AOI21X1  g0156(.A0(n851_1), .A1(n842), .B0(n863), .Y(n864));
OR4X1    g0217(.A(n921_1), .B(n918), .C(n915), .D(n905), .Y(n926_1));
NOR3X1   g0222(.A(n930), .B(n928), .C(n927), .Y(n931_1));
OR4X1    g0224(.A(n927), .B(n924), .C(n904), .D(n928), .Y(n933));
NOR4X1   g0225(.A(n921_1), .B(n918), .C(n915), .D(n930), .Y(n934));
NOR3X1   g0231(.A(g688), .B(n939), .C(n758), .Y(n940));
NAND2X1  g0054(.A(g699), .B(g702), .Y(n762));
OAI21X1  g0019(.A0(n726_1), .A1(n724), .B0(g676), .Y(n727));
NAND2X1  g0053(.A(n760), .B(g662), .Y(n761_1));
INVX1    g0017(.A(g41), .Y(n725));
INVX1    g0108(.A(n807), .Y(n816_1));
AOI22X1  g0103(.A0(n767), .A1(g297), .B0(n763), .B1(n810), .Y(n811_1));
INVX1    g0109(.A(n814), .Y(n817));
MX2X1    g0099(.A(n805), .B(n806_1), .S0(g658), .Y(n807));
INVX1    g0095(.A(g212), .Y(n803));
INVX1    g0094(.A(g678), .Y(n802));
MX2X1    g0106(.A(n812), .B(n813), .S0(n760), .Y(n814));
NOR4X1   g0155(.A(n854), .B(n853), .C(n852), .D(n862), .Y(n863));
NOR4X1   g0134(.A(n839), .B(n837), .C(n833), .D(n841_1), .Y(n842));
NOR4X1   g0143(.A(n848), .B(n846_1), .C(n844), .D(n850), .Y(n851_1));
INVX1    g0197(.A(g283), .Y(n905));
AOI21X1  g0207(.A0(n914), .A1(n909), .B0(n871_1), .Y(n915));
NOR2X1   g0210(.A(n917), .B(n871_1), .Y(n918));
NAND2X1  g0213(.A(n920), .B(n919), .Y(n921_1));
AOI21X1  g0218(.A0(n914), .A1(n909), .B0(n870), .Y(n927));
NOR2X1   g0219(.A(n917), .B(n870), .Y(n928));
AND2X1   g0221(.A(n929), .B(n917), .Y(n930));
INVX1    g0196(.A(g282), .Y(n904));
OAI21X1  g0216(.A0(n923), .A1(n912), .B0(n922), .Y(n924));
INVX1    g0050(.A(g689), .Y(n758));
INVX1    g0230(.A(g698), .Y(n939));
AND2X1   g0016(.A(n723), .B(n716_1), .Y(n724));
OAI21X1  g0018(.A0(n723), .A1(n716_1), .B0(n725), .Y(n726_1));
INVX1    g0052(.A(g658), .Y(n760));
NOR3X1   g0102(.A(n809), .B(n808), .C(n757), .Y(n810));
NOR4X1   g0055(.A(n761_1), .B(n727), .C(g41), .D(n762), .Y(n763));
INVX1    g0098(.A(g218), .Y(n806_1));
INVX1    g0097(.A(g679), .Y(n805));
INVX1    g0105(.A(g680), .Y(n813));
INVX1    g0104(.A(g224), .Y(n812));
NAND3X1  g0154(.A(n861_1), .B(n856_1), .C(n855), .Y(n862));
XOR2X1   g0144(.A(g288), .B(g682), .Y(n852));
XOR2X1   g0145(.A(g683), .B(g289), .Y(n853));
XOR2X1   g0146(.A(g287), .B(g681), .Y(n854));
NOR4X1   g0133(.A(g634), .B(g598), .C(g567), .D(n496), .Y(n841_1));
NOR4X1   g0125(.A(g634), .B(g598), .C(n831_1), .D(n916), .Y(n833));
NOR4X1   g0129(.A(n835), .B(n834), .C(n831_1), .D(n836_1), .Y(n837));
NOR4X1   g0131(.A(g634), .B(n834), .C(g567), .D(n838), .Y(n839));
NOR4X1   g0142(.A(n836_1), .B(g598), .C(g567), .D(n849), .Y(n850));
NOR4X1   g0136(.A(g634), .B(n834), .C(n831_1), .D(n843), .Y(n844));
NOR4X1   g0138(.A(g598), .B(n845), .C(n831_1), .D(n836_1), .Y(n846_1));
NOR4X1   g0140(.A(n836_1), .B(n834), .C(g567), .D(n847), .Y(n848));
INVX1    g0163(.A(n870), .Y(n871_1));
OAI21X1  g0201(.A0(n903), .A1(n889), .B0(n908), .Y(n909));
INVX1    g0206(.A(n913), .Y(n914));
OAI21X1  g0209(.A0(n903), .A1(n889), .B0(n916_1), .Y(n917));
NAND3X1  g0211(.A(n870), .B(g283), .C(n904), .Y(n919));
OR4X1    g0212(.A(g478), .B(g283), .C(g282), .D(n911_1), .Y(n920));
NOR4X1   g0162(.A(n868), .B(n867), .C(n866_1), .D(n869), .Y(n870));
NOR3X1   g0220(.A(n871_1), .B(g283), .C(n904), .Y(n929));
NAND4X1  g0214(.A(n872), .B(n905), .C(n904), .D(n911_1), .Y(n922));
XOR2X1   g0204(.A(n911_1), .B(n872), .Y(n912));
NAND3X1  g0215(.A(n907), .B(n905), .C(g282), .Y(n923));
INVX1    g0008(.A(g48), .Y(n716_1));
XOR2X1   g0015(.A(n722), .B(n719), .Y(n723));
INVX1    g0049(.A(g687), .Y(n757));
INVX1    g0100(.A(g688), .Y(n808));
OR2X1    g0101(.A(g698), .B(g689), .Y(n809));
XOR2X1   g0147(.A(g286), .B(n813), .Y(n855));
XOR2X1   g0148(.A(g284), .B(n802), .Y(n856_1));
NOR4X1   g0153(.A(n859), .B(n858), .C(n857), .D(n860), .Y(n861_1));
INVX1    g0132(.A(g690), .Y(n496));
INVX1    g0124(.A(g691), .Y(n916));
INVX1    g0123(.A(g567), .Y(n831_1));
INVX1    g0128(.A(g634), .Y(n836_1));
INVX1    g0126(.A(g598), .Y(n834));
INVX1    g0127(.A(g697), .Y(n835));
INVX1    g0130(.A(g692), .Y(n838));
INVX1    g0141(.A(g694), .Y(n849));
INVX1    g0135(.A(g693), .Y(n843));
INVX1    g0137(.A(g695), .Y(n845));
INVX1    g0139(.A(g696), .Y(n847));
NOR3X1   g0200(.A(n907), .B(n905), .C(n904), .Y(n908));
AOI21X1  g0181(.A0(n888), .A1(n887), .B0(n872), .Y(n889));
NOR3X1   g0195(.A(n902), .B(n901_1), .C(g478), .Y(n903));
NOR4X1   g0205(.A(n906_1), .B(n905), .C(n904), .D(n912), .Y(n913));
NOR3X1   g0208(.A(n907), .B(g283), .C(n904), .Y(n916_1));
NOR2X1   g0203(.A(n910), .B(n906_1), .Y(n911_1));
NAND3X1  g0161(.A(g277), .B(g276), .C(g278), .Y(n869));
INVX1    g0158(.A(g281), .Y(n866_1));
INVX1    g0159(.A(g279), .Y(n867));
INVX1    g0160(.A(g280), .Y(n868));
INVX1    g0164(.A(g478), .Y(n872));
INVX1    g0199(.A(n906_1), .Y(n907));
XOR2X1   g0011(.A(n718), .B(n717), .Y(n719));
XOR2X1   g0014(.A(n721_1), .B(n720), .Y(n722));
XOR2X1   g0152(.A(g686), .B(g292), .Y(n860));
XOR2X1   g0149(.A(g290), .B(g684), .Y(n857));
XOR2X1   g0150(.A(g679), .B(g285), .Y(n858));
XOR2X1   g0151(.A(g685), .B(g291), .Y(n859));
NAND2X1  g0179(.A(n886_1), .B(n867), .Y(n887));
NAND2X1  g0180(.A(n886_1), .B(g279), .Y(n888));
NOR2X1   g0193(.A(n900), .B(g279), .Y(n901_1));
NOR2X1   g0194(.A(n900), .B(n867), .Y(n902));
XOR2X1   g0198(.A(g280), .B(n866_1), .Y(n906_1));
NOR4X1   g0202(.A(g280), .B(n867), .C(n866_1), .D(n869), .Y(n910));
XOR2X1   g0009(.A(g1), .B(g2), .Y(n717));
XOR2X1   g0010(.A(g10), .B(g6), .Y(n718));
XOR2X1   g0012(.A(g14), .B(g18), .Y(n720));
XOR2X1   g0013(.A(g28), .B(g24), .Y(n721_1));
AOI22X1  g0178(.A0(n881_1), .A1(n885), .B0(n879), .B1(n874), .Y(n886_1));
OAI22X1  g0192(.A0(n896_1), .A1(n899), .B0(n894), .B1(n891_1), .Y(n900));
OAI21X1  g0166(.A0(n835), .A1(g276), .B0(n873), .Y(n874));
AOI21X1  g0171(.A0(n878), .A1(n876_1), .B0(g278), .Y(n879));
AOI21X1  g0177(.A0(n884), .A1(n883), .B0(n882), .Y(n885));
OAI21X1  g0173(.A0(n843), .A1(g276), .B0(n880), .Y(n881_1));
AND2X1   g0183(.A(n873), .B(n890), .Y(n891_1));
OAI21X1  g0186(.A0(n893), .A1(n892), .B0(n882), .Y(n894));
OAI21X1  g0191(.A0(n898), .A1(n897), .B0(g278), .Y(n899));
AND2X1   g0188(.A(n880), .B(n895), .Y(n896_1));
AOI21X1  g0165(.A0(g696), .A1(g276), .B0(g277), .Y(n873));
NAND2X1  g0168(.A(n875), .B(g695), .Y(n876_1));
AOI21X1  g0170(.A0(g694), .A1(g276), .B0(n877), .Y(n878));
INVX1    g0174(.A(g278), .Y(n882));
NAND2X1  g0175(.A(g691), .B(n875), .Y(n883));
AOI21X1  g0176(.A0(g690), .A1(g276), .B0(n877), .Y(n884));
AOI21X1  g0172(.A0(g692), .A1(g276), .B0(g277), .Y(n880));
NAND2X1  g0182(.A(g697), .B(n875), .Y(n890));
NOR2X1   g0184(.A(g276), .B(n845), .Y(n892));
OAI21X1  g0185(.A0(n849), .A1(n875), .B0(g277), .Y(n893));
NOR2X1   g0189(.A(n916), .B(g276), .Y(n897));
OAI21X1  g0190(.A0(n496), .A1(n875), .B0(g277), .Y(n898));
NAND2X1  g0187(.A(g693), .B(n875), .Y(n895));
INVX1    g0167(.A(g276), .Y(n875));
INVX1    g0169(.A(g277), .Y(n877));

endmodule
