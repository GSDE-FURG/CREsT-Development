//Converted to Combinational , Module name: s510 , Timestamp: 2018-12-03T15:51:01.852024 
module s510 ( john, cnt13, cnt21, cnt284, pcnt6, cnt261, cnt44, pcnt12, pcnt17, cnt591, cnt45, cnt567, pcnt27, cnt283, cnt272, cnt10, cnt511, pcnt241, cnt509, st_5, st_4, st_3, st_2, st_1, st_0, csm, pclr, cclr, vsync, cblank, csync, n53, n58, n63, n68, n73, n78 );
input john, cnt13, cnt21, cnt284, pcnt6, cnt261, cnt44, pcnt12, pcnt17, cnt591, cnt45, cnt567, pcnt27, cnt283, cnt272, cnt10, cnt511, pcnt241, cnt509, st_5, st_4, st_3, st_2, st_1, st_0;
output csm, pclr, cclr, vsync, cblank, csync, n53, n58, n63, n68, n73, n78;
wire pc, n44, n45, n47, n48, n49, n50, n51, n52, n53_1, n54, n55, n56, n58_1, n59, n60, n61, n62, n64, n65, n66, n67, n68_1, n69, n70, n71, n73_1, n74, n75, n76, n77, n79, n80, n81, n82, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n95, n96, n97, n98, n99, n100, n101, n103, n104, n105, n106, n107, n109, n110, n111, n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187;
NOR2X1   g000(.A(st_0), .B(st_1), .Y(n44));
NAND3X1  g001(.A(st_2), .B(st_3), .C(st_5), .Y(n45));
NOR2X1   g002(.A(n45), .B(n44), .Y(csm));
INVX1    g003(.A(st_4), .Y(n47));
INVX1    g004(.A(st_2), .Y(n48));
NAND3X1  g005(.A(st_0), .B(n48), .C(n47), .Y(n49));
INVX1    g006(.A(st_5), .Y(n50));
AND2X1   g007(.A(st_1), .B(st_3), .Y(n51));
NAND2X1  g008(.A(n51), .B(n50), .Y(n52));
INVX1    g009(.A(st_3), .Y(n53_1));
AND2X1   g010(.A(st_0), .B(st_4), .Y(n54));
AND2X1   g011(.A(st_1), .B(st_2), .Y(n55));
NAND3X1  g012(.A(n55), .B(n54), .C(n53_1), .Y(n56));
OAI21X1  g013(.A0(n52), .A1(n49), .B0(n56), .Y(pclr));
NOR4X1   g014(.A(st_2), .B(st_3), .C(st_5), .D(st_1), .Y(n58_1));
AND2X1   g015(.A(n58_1), .B(n47), .Y(n59));
OR2X1    g016(.A(n51), .B(st_5), .Y(n60));
NAND3X1  g017(.A(n54), .B(n51), .C(st_2), .Y(n61));
OAI21X1  g018(.A0(n60), .A1(n49), .B0(n61), .Y(n62));
OR2X1    g019(.A(n62), .B(n59), .Y(pc));
OR2X1    g020(.A(st_3), .B(st_5), .Y(n64));
NAND3X1  g021(.A(n64), .B(st_0), .C(st_1), .Y(n65));
INVX1    g022(.A(st_1), .Y(n66));
NAND3X1  g023(.A(st_0), .B(n66), .C(n50), .Y(n67));
OAI21X1  g024(.A0(n48), .A1(st_4), .B0(st_0), .Y(n68_1));
OR2X1    g025(.A(st_0), .B(st_1), .Y(n69));
NOR4X1   g026(.A(n48), .B(st_3), .C(n50), .D(n69), .Y(n70));
NOR2X1   g027(.A(n70), .B(n59), .Y(n71));
NAND4X1  g028(.A(n68_1), .B(n67), .C(n65), .D(n71), .Y(cclr));
NAND2X1  g029(.A(n55), .B(n47), .Y(n73_1));
AOI21X1  g030(.A0(st_0), .A1(st_1), .B0(st_3), .Y(n74));
NAND3X1  g031(.A(n66), .B(st_2), .C(n50), .Y(n75));
OR2X1    g032(.A(st_4), .B(st_5), .Y(n76));
OAI21X1  g033(.A0(n76), .A1(n44), .B0(n48), .Y(n77));
NAND4X1  g034(.A(n75), .B(n74), .C(n73_1), .D(n77), .Y(vsync));
INVX1    g035(.A(st_0), .Y(n79));
AOI21X1  g036(.A0(st_3), .A1(st_4), .B0(st_5), .Y(n80));
OR4X1    g037(.A(n79), .B(n66), .C(st_2), .D(n80), .Y(n81));
NAND4X1  g038(.A(st_2), .B(st_3), .C(n47), .D(n79), .Y(n82));
NAND3X1  g039(.A(n82), .B(n81), .C(n45), .Y(cblank));
XOR2X1   g040(.A(st_1), .B(st_2), .Y(n84));
AOI22X1  g041(.A0(n64), .A1(st_1), .B0(n47), .B1(n84), .Y(n85));
OR2X1    g042(.A(n85), .B(st_0), .Y(n86));
NAND4X1  g043(.A(st_0), .B(n47), .C(n50), .D(n55), .Y(n87));
NOR2X1   g044(.A(st_4), .B(st_5), .Y(n88));
NOR3X1   g045(.A(n48), .B(n53_1), .C(st_4), .Y(n89));
NOR2X1   g046(.A(st_0), .B(n53_1), .Y(n90));
AOI21X1  g047(.A0(n90), .A1(n88), .B0(n89), .Y(n91));
NOR3X1   g048(.A(n88), .B(n79), .C(st_2), .Y(n92));
AOI21X1  g049(.A0(n54), .A1(n66), .B0(n92), .Y(n93));
NAND4X1  g050(.A(n91), .B(n87), .C(n86), .D(n93), .Y(csync));
NOR3X1   g051(.A(st_0), .B(n66), .C(n50), .Y(n95));
NOR4X1   g052(.A(st_1), .B(st_2), .C(st_4), .D(n79), .Y(n96));
OAI21X1  g053(.A0(n96), .A1(n95), .B0(n53_1), .Y(n97));
NOR2X1   g054(.A(st_0), .B(st_2), .Y(n98));
AOI21X1  g055(.A0(n79), .A1(st_1), .B0(n53_1), .Y(n99));
OAI21X1  g056(.A0(n99), .A1(n98), .B0(st_5), .Y(n100));
NAND3X1  g057(.A(n60), .B(st_0), .C(st_2), .Y(n101));
NAND3X1  g058(.A(n101), .B(n100), .C(n97), .Y(n53));
NAND4X1  g059(.A(st_0), .B(n47), .C(n50), .D(n84), .Y(n103));
OAI21X1  g060(.A0(n58_1), .A1(st_4), .B0(n79), .Y(n104));
NAND4X1  g061(.A(st_2), .B(st_3), .C(st_5), .D(st_1), .Y(n105));
NOR4X1   g062(.A(st_1), .B(st_2), .C(st_5), .D(n79), .Y(n106));
NAND2X1  g063(.A(n106), .B(st_3), .Y(n107));
NAND4X1  g064(.A(n105), .B(n104), .C(n103), .D(n107), .Y(n58));
NAND2X1  g065(.A(st_0), .B(st_4), .Y(n109));
NOR2X1   g066(.A(n109), .B(st_3), .Y(n110));
OAI21X1  g067(.A0(n89), .A1(n110), .B0(n66), .Y(n111));
NOR3X1   g068(.A(n79), .B(st_2), .C(st_4), .Y(n112));
AND2X1   g069(.A(st_0), .B(st_5), .Y(n113));
OAI21X1  g070(.A0(n113), .A1(n112), .B0(st_1), .Y(n114));
NOR3X1   g071(.A(n88), .B(st_2), .C(n53_1), .Y(n115));
AOI21X1  g072(.A0(n90), .A1(n50), .B0(n115), .Y(n116));
NAND3X1  g073(.A(n116), .B(n114), .C(n111), .Y(n63));
NOR3X1   g074(.A(n79), .B(n66), .C(st_2), .Y(n118));
NAND2X1  g075(.A(st_3), .B(n47), .Y(n119));
NAND3X1  g076(.A(st_2), .B(st_3), .C(n47), .Y(n120));
NAND3X1  g077(.A(n66), .B(st_2), .C(st_3), .Y(n121));
NAND2X1  g078(.A(n121), .B(n120), .Y(n122));
AOI21X1  g079(.A0(n119), .A1(n118), .B0(n122), .Y(n123));
NAND2X1  g080(.A(n50), .B(cnt13), .Y(n124));
NAND3X1  g081(.A(n124), .B(n55), .C(n79), .Y(n125));
AOI22X1  g082(.A0(n106), .A1(n47), .B0(n84), .B1(n113), .Y(n126));
OR2X1    g083(.A(n64), .B(n79), .Y(n127));
INVX1    g084(.A(cnt284), .Y(n128));
NOR2X1   g085(.A(pcnt17), .B(n128), .Y(n129));
OAI22X1  g086(.A0(n127), .A1(n129), .B0(n109), .B1(st_3), .Y(n130));
OAI22X1  g087(.A0(n48), .A1(n47), .B0(cnt284), .B1(n75), .Y(n131));
AOI22X1  g088(.A0(n130), .A1(st_1), .B0(n79), .B1(n131), .Y(n132));
NAND4X1  g089(.A(n126), .B(n125), .C(n123), .D(n132), .Y(n68));
NOR3X1   g090(.A(n109), .B(n48), .C(st_3), .Y(n134));
NAND3X1  g091(.A(n54), .B(n66), .C(st_3), .Y(n135));
NAND3X1  g092(.A(n76), .B(n79), .C(st_1), .Y(n136));
NAND2X1  g093(.A(n136), .B(n135), .Y(n137));
OR4X1    g094(.A(n79), .B(st_2), .C(n50), .D(n51), .Y(n138));
OAI21X1  g095(.A0(n120), .A1(n79), .B0(n138), .Y(n139));
NAND3X1  g096(.A(n55), .B(n79), .C(st_3), .Y(n140));
INVX1    g097(.A(cnt511), .Y(n141));
NOR2X1   g098(.A(pcnt241), .B(n141), .Y(n142));
NAND2X1  g099(.A(st_1), .B(st_2), .Y(n143));
OR4X1    g100(.A(st_0), .B(st_3), .C(cnt13), .D(n143), .Y(n144));
OAI21X1  g101(.A0(n142), .A1(n140), .B0(n144), .Y(n145));
OR4X1    g102(.A(n139), .B(n137), .C(n134), .D(n145), .Y(n146));
NAND2X1  g103(.A(n58_1), .B(n47), .Y(n147));
NAND3X1  g104(.A(st_2), .B(n53_1), .C(st_5), .Y(n148));
AOI21X1  g105(.A0(n148), .A1(n147), .B0(st_0), .Y(n149));
INVX1    g106(.A(pcnt12), .Y(n150));
NAND4X1  g107(.A(st_1), .B(n48), .C(n53_1), .D(n79), .Y(n151));
AOI21X1  g108(.A0(n150), .A1(cnt44), .B0(n151), .Y(n152));
AOI21X1  g109(.A0(pcnt17), .A1(cnt284), .B0(st_3), .Y(n153));
NAND4X1  g110(.A(n55), .B(st_0), .C(n50), .D(n153), .Y(n154));
INVX1    g111(.A(cnt567), .Y(n155));
NOR2X1   g112(.A(pcnt27), .B(n155), .Y(n156));
NAND2X1  g113(.A(n98), .B(n51), .Y(n157));
OAI21X1  g114(.A0(n157), .A1(n156), .B0(n154), .Y(n158));
OR4X1    g115(.A(n152), .B(n149), .C(n146), .D(n158), .Y(n73));
INVX1    g116(.A(cnt10), .Y(n160));
NOR4X1   g117(.A(st_0), .B(n53_1), .C(n160), .D(n143), .Y(n161));
OR2X1    g118(.A(st_0), .B(cnt21), .Y(n162));
NAND4X1  g119(.A(n66), .B(st_2), .C(st_3), .D(n162), .Y(n163));
NAND3X1  g120(.A(n98), .B(n53_1), .C(cnt21), .Y(n164));
NAND4X1  g121(.A(st_2), .B(n53_1), .C(cnt45), .D(n44), .Y(n165));
NAND3X1  g122(.A(n98), .B(n51), .C(cnt283), .Y(n166));
NAND4X1  g123(.A(n165), .B(n164), .C(n163), .D(n166), .Y(n167));
OAI21X1  g124(.A0(n167), .A1(n161), .B0(st_4), .Y(n168));
NOR4X1   g125(.A(st_0), .B(n53_1), .C(n141), .D(n143), .Y(n169));
NAND2X1  g126(.A(pcnt6), .B(cnt284), .Y(n170));
OR4X1    g127(.A(n69), .B(n48), .C(st_3), .D(n170), .Y(n171));
OAI21X1  g128(.A0(n157), .A1(n155), .B0(n171), .Y(n172));
OAI21X1  g129(.A0(n172), .A1(n169), .B0(n88), .Y(n173));
AOI22X1  g130(.A0(st_5), .A1(cnt10), .B0(john), .B1(st_4), .Y(n174));
NOR4X1   g131(.A(n143), .B(st_0), .C(st_3), .D(n174), .Y(n175));
NOR4X1   g132(.A(n79), .B(st_1), .C(cnt261), .D(n148), .Y(n176));
MX2X1    g133(.A(cnt591), .B(cnt272), .S0(st_2), .Y(n177));
NOR4X1   g134(.A(n53_1), .B(st_4), .C(st_5), .D(n69), .Y(n178));
AND2X1   g135(.A(n178), .B(n177), .Y(n179));
NOR4X1   g136(.A(n64), .B(n79), .C(st_4), .D(n84), .Y(n180));
NOR4X1   g137(.A(n179), .B(n176), .C(n175), .D(n180), .Y(n181));
NAND4X1  g138(.A(st_1), .B(n48), .C(st_5), .D(n79), .Y(n182));
OAI21X1  g139(.A0(n151), .A1(st_4), .B0(n182), .Y(n183));
NAND2X1  g140(.A(st_5), .B(cnt509), .Y(n184));
NAND3X1  g141(.A(n66), .B(n48), .C(cnt45), .Y(n185));
OAI22X1  g142(.A0(n184), .A1(n121), .B0(n80), .B1(n185), .Y(n186));
AOI22X1  g143(.A0(n183), .A1(cnt44), .B0(n79), .B1(n186), .Y(n187));
NAND4X1  g144(.A(n181), .B(n173), .C(n168), .D(n187), .Y(n78));
endmodule
