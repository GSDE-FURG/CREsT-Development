//Converted to Combinational , Module name: s38417 , Timestamp: 2018-12-03T15:51:11.524459 
module s38417 ( g51, g563, g1249, g1943, g2637, g3212, g3213, g3214, g3215, g3216, g3217, g3218, g3219, g3220, g3221, g3222, g3223, g3224, g3225, g3226, g3227, g3228, g3229, g3230, g3231, g3232, g3233, g3234, g2814, g2817, g2933, g2950, g2883, g2888, g2896, g2892, g2903, g2900, g2908, g2912, g2917, g2924, g2920, g2984, g2985, g2930, g2929, g2879, g2934, g2935, g2938, g2941, g2944, g2947, g2953, g2956, g2959, g2962, g2963, g2966, g2969, g2972, g2975, g2978, g2981, g2874, g1506, g1501, g1496, g1491, g1486, g1481, g1476, g1471, g2877, g2861, g813, g2864, g809, g2867, g805, g2870, g801, g2818, g797, g2821, g793, g2824, g789, g2827, g785, g2830, g2873, g2833, g125, g2836, g121, g2839, g117, g2842, g113, g2845, g109, g2848, g105, g2851, g101, g2854, g97, g2858, g2857, g2200, g2195, g2190, g2185, g2180, g2175, g2170, g2165, g2878, g3129, g3117, g3109, g3210, g3211, g3084, g3085, g3086, g3087, g3091, g3092, g3093, g3094, g3095, g3096, g3097, g3098, g3099, g3100, g3101, g3102, g3103, g3104, g3105, g3106, g3107, g3108, g3155, g3158, g3161, g3164, g3167, g3170, g3173, g3176, g3179, g3182, g3185, g3088, g3191, g3194, g3197, g3198, g3201, g3204, g3207, g3188, g3133, g3132, g3128, g3127, g3126, g3125, g3124, g3123, g3120, g3114, g3113, g3112, g3110, g3111, g3139, g3136, g3134, g3135, g3151, g3142, g3147, g185, g138, g135, g165, g130, g131, g129, g133, g134, g132, g142, g143, g141, g145, g146, g144, g151, g152, g154, g155, g153, g157, g158, g156, g160, g161, g159, g163, g164, g162, g169, g170, g168, g172, g173, g171, g175, g176, g174, g178, g179, g177, g186, g189, g192, g231, g234, g237, g195, g198, g201, g240, g243, g246, g204, g207, g210, g249, g252, g255, g213, g258, g261, g264, g222, g225, g228, g267, g270, g273, g92, g88, g83, g74, g70, g65, g61, g52, g180, g182, g181, g276, g405, g401, g354, g343, g346, g369, g358, g361, g384, g373, g376, g398, g388, g391, g408, g411, g414, g417, g420, g423, g427, g428, g426, g429, g432, g435, g438, g441, g444, g448, g449, g447, g403, g404, g402, g450, g451, g452, g453, g454, g279, g280, g299, g305, g304, g303, g302, g301, g300, g342, g349, g350, g351, g352, g353, g357, g364, g365, g366, g367, g368, g372, g379, g380, g381, g382, g383, g387, g394, g395, g396, g397, g324, g325, g331, g337, g545, g551, g550, g554, g557, g510, g513, g523, g524, g564, g569, g570, g571, g572, g573, g574, g565, g566, g567, g568, g489, g474, g481, g485, g486, g487, g488, g455, g458, g461, g477, g478, g479, g480, g484, g464, g465, g468, g471, g528, g535, g542, g543, g544, g548, g549, g499, g558, g559, g576, g577, g575, g579, g580, g578, g582, g583, g581, g585, g586, g584, g587, g590, g593, g596, g599, g602, g614, g617, g620, g605, g608, g611, g490, g493, g496, g506, g507, g508, g509, g514, g515, g516, g517, g518, g519, g520, g525, g529, g530, g531, g532, g533, g534, g536, g537, g538, g541, g623, g626, g629, g630, g659, g640, g633, g653, g646, g660, g672, g666, g679, g686, g692, g699, g700, g698, g702, g703, g701, g705, g706, g704, g708, g709, g707, g711, g712, g710, g714, g715, g713, g717, g718, g716, g720, g721, g719, g723, g724, g722, g726, g727, g725, g729, g730, g728, g732, g733, g731, g735, g736, g734, g738, g739, g737, g826, g823, g853, g818, g819, g817, g821, g822, g820, g830, g831, g829, g833, g834, g832, g836, g837, g835, g839, g840, g838, g842, g843, g841, g845, g846, g844, g848, g849, g847, g851, g852, g850, g857, g858, g856, g860, g861, g859, g863, g864, g862, g866, g867, g865, g873, g876, g879, g918, g921, g924, g882, g885, g888, g927, g930, g933, g891, g894, g897, g936, g939, g942, g900, g903, g906, g945, g948, g951, g909, g912, g915, g954, g957, g960, g780, g776, g771, g767, g762, g758, g753, g749, g744, g740, g868, g870, g869, g963, g1092, g1088, g996, g1041, g1030, g1033, g1056, g1045, g1048, g1071, g1060, g1063, g1085, g1075, g1078, g1095, g1098, g1101, g1104, g1107, g1110, g1114, g1115, g1113, g1116, g1119, g1122, g1125, g1128, g1131, g1135, g1136, g1134, g999, g1000, g1001, g1002, g1003, g1004, g1005, g1006, g1007, g1009, g1010, g1008, g1090, g1091, g1089, g1137, g1138, g1139, g1140, g1141, g966, g967, g968, g969, g970, g971, g972, g973, g974, g975, g976, g977, g978, g986, g992, g995, g984, g983, g982, g981, g991, g990, g989, g988, g987, g985, g1029, g1036, g1037, g1038, g1039, g1040, g1044, g1051, g1052, g1053, g1054, g1055, g1059, g1066, g1067, g1068, g1069, g1070, g1074, g1081, g1082, g1083, g1084, g1011, g1012, g1018, g1024, g1231, g1237, g1236, g1240, g1243, g1196, g1199, g1209, g1210, g1250, g1255, g1256, g1257, g1258, g1259, g1260, g1251, g1252, g1253, g1254, g1176, g1161, g1168, g1172, g1173, g1174, g1175, g1142, g1145, g1148, g1164, g1165, g1166, g1167, g1171, g1151, g1152, g1155, g1158, g1214, g1221, g1228, g1229, g1230, g1234, g1235, g1186, g1244, g1245, g1262, g1263, g1261, g1265, g1266, g1264, g1268, g1269, g1267, g1271, g1272, g1270, g1273, g1276, g1279, g1282, g1285, g1288, g1300, g1303, g1306, g1291, g1294, g1297, g1177, g1180, g1183, g1192, g1193, g1194, g1195, g1200, g1201, g1202, g1203, g1204, g1205, g1206, g1211, g1215, g1216, g1217, g1218, g1219, g1220, g1222, g1223, g1224, g1227, g1309, g1312, g1315, g1316, g1345, g1326, g1319, g1339, g1332, g1346, g1358, g1352, g1365, g1372, g1378, g1385, g1386, g1384, g1388, g1389, g1387, g1391, g1392, g1390, g1394, g1395, g1393, g1397, g1398, g1396, g1400, g1401, g1399, g1403, g1404, g1402, g1406, g1407, g1405, g1409, g1410, g1408, g1412, g1413, g1411, g1415, g1416, g1414, g1418, g1419, g1417, g1421, g1422, g1420, g1424, g1425, g1423, g1520, g1517, g1547, g1512, g1513, g1511, g1515, g1516, g1514, g1524, g1525, g1523, g1527, g1528, g1526, g1530, g1531, g1529, g1533, g1534, g1532, g1536, g1537, g1535, g1539, g1540, g1538, g1542, g1543, g1541, g1545, g1546, g1544, g1551, g1552, g1550, g1554, g1555, g1553, g1557, g1558, g1556, g1560, g1561, g1559, g1567, g1570, g1573, g1612, g1615, g1618, g1576, g1579, g1582, g1621, g1624, g1627, g1585, g1588, g1591, g1630, g1633, g1636, g1594, g1597, g1600, g1639, g1642, g1645, g1603, g1606, g1609, g1648, g1651, g1654, g1466, g1462, g1457, g1453, g1448, g1444, g1439, g1435, g1430, g1426, g1562, g1564, g1563, g1657, g1786, g1782, g1690, g1735, g1724, g1727, g1750, g1739, g1742, g1765, g1754, g1757, g1779, g1769, g1772, g1789, g1792, g1795, g1798, g1801, g1804, g1808, g1809, g1807, g1810, g1813, g1816, g1819, g1822, g1825, g1829, g1830, g1828, g1693, g1694, g1695, g1696, g1697, g1698, g1699, g1700, g1701, g1703, g1704, g1702, g1784, g1785, g1783, g1831, g1832, g1833, g1834, g1835, g1660, g1661, g1662, g1663, g1664, g1665, g1666, g1667, g1668, g1669, g1670, g1671, g1672, g1680, g1686, g1689, g1678, g1677, g1676, g1675, g1685, g1684, g1683, g1682, g1681, g1679, g1723, g1730, g1731, g1732, g1733, g1734, g1738, g1745, g1746, g1747, g1748, g1749, g1753, g1760, g1761, g1762, g1763, g1764, g1768, g1775, g1776, g1777, g1778, g1705, g1706, g1712, g1718, g1925, g1931, g1930, g1934, g1937, g1890, g1893, g1903, g1904, g1944, g1949, g1950, g1951, g1952, g1953, g1954, g1945, g1946, g1947, g1948, g1870, g1855, g1862, g1866, g1867, g1868, g1869, g1836, g1839, g1842, g1858, g1859, g1860, g1861, g1865, g1845, g1846, g1849, g1852, g1908, g1915, g1922, g1923, g1924, g1928, g1929, g1880, g1938, g1939, g1956, g1957, g1955, g1959, g1960, g1958, g1962, g1963, g1961, g1965, g1966, g1964, g1967, g1970, g1973, g1976, g1979, g1982, g1994, g1997, g2000, g1985, g1988, g1991, g1871, g1874, g1877, g1886, g1887, g1888, g1889, g1894, g1895, g1896, g1897, g1898, g1899, g1900, g1905, g1909, g1910, g1911, g1912, g1913, g1914, g1916, g1917, g1918, g1921, g2003, g2006, g2009, g2010, g2039, g2020, g2013, g2033, g2026, g2040, g2052, g2046, g2059, g2066, g2072, g2079, g2080, g2078, g2082, g2083, g2081, g2085, g2086, g2084, g2088, g2089, g2087, g2091, g2092, g2090, g2094, g2095, g2093, g2097, g2098, g2096, g2100, g2101, g2099, g2103, g2104, g2102, g2106, g2107, g2105, g2109, g2110, g2108, g2112, g2113, g2111, g2115, g2116, g2114, g2118, g2119, g2117, g2214, g2211, g2241, g2206, g2207, g2205, g2209, g2210, g2208, g2218, g2219, g2217, g2221, g2222, g2220, g2224, g2225, g2223, g2227, g2228, g2226, g2230, g2231, g2229, g2233, g2234, g2232, g2236, g2237, g2235, g2239, g2240, g2238, g2245, g2246, g2244, g2248, g2249, g2247, g2251, g2252, g2250, g2254, g2255, g2253, g2261, g2264, g2267, g2306, g2309, g2312, g2270, g2273, g2276, g2315, g2318, g2321, g2279, g2282, g2285, g2324, g2327, g2330, g2288, g2291, g2294, g2333, g2336, g2339, g2297, g2300, g2303, g2342, g2345, g2348, g2160, g2156, g2151, g2147, g2142, g2138, g2133, g2129, g2124, g2120, g2256, g2258, g2257, g2351, g2480, g2476, g2384, g2429, g2418, g2421, g2444, g2433, g2436, g2459, g2448, g2451, g2473, g2463, g2466, g2483, g2486, g2489, g2492, g2495, g2498, g2502, g2503, g2501, g2504, g2507, g2510, g2513, g2516, g2519, g2523, g2524, g2522, g2387, g2388, g2389, g2390, g2391, g2392, g2393, g2394, g2395, g2397, g2398, g2396, g2478, g2479, g2477, g2525, g2526, g2527, g2528, g2529, g2354, g2355, g2356, g2357, g2358, g2359, g2360, g2361, g2362, g2363, g2364, g2365, g2366, g2374, g2380, g2383, g2372, g2371, g2370, g2369, g2379, g2378, g2377, g2376, g2375, g2373, g2417, g2424, g2425, g2426, g2427, g2428, g2432, g2439, g2440, g2441, g2442, g2443, g2447, g2454, g2455, g2456, g2457, g2458, g2462, g2469, g2470, g2471, g2472, g2399, g2400, g2406, g2412, g2619, g2625, g2624, g2628, g2631, g2584, g2587, g2597, g2598, g2638, g2643, g2644, g2645, g2646, g2647, g2648, g2639, g2640, g2641, g2642, g2564, g2549, g2556, g2560, g2561, g2562, g2563, g2530, g2533, g2536, g2552, g2553, g2554, g2555, g2559, g2539, g2540, g2543, g2546, g2602, g2609, g2616, g2617, g2618, g2622, g2623, g2574, g2632, g2633, g2650, g2651, g2649, g2653, g2654, g2652, g2656, g2657, g2655, g2659, g2660, g2658, g2661, g2664, g2667, g2670, g2673, g2676, g2688, g2691, g2694, g2679, g2682, g2685, g2565, g2568, g2571, g2580, g2581, g2582, g2583, g2588, g2589, g2590, g2591, g2592, g2593, g2594, g2599, g2603, g2604, g2605, g2606, g2607, g2608, g2610, g2611, g2612, g2615, g2697, g2700, g2703, g2704, g2733, g2714, g2707, g2727, g2720, g2734, g2746, g2740, g2753, g2760, g2766, g2773, g2774, g2772, g2776, g2777, g2775, g2779, g2780, g2778, g2782, g2783, g2781, g2785, g2786, g2784, g2788, g2789, g2787, g2791, g2792, g2790, g2794, g2795, g2793, g2797, g2798, g2796, g2800, g2801, g2799, g2803, g2804, g2802, g2806, g2807, g2805, g2809, g2810, g2808, g2812, g2813, g2811, g3054, g3079, g3080, g3043, g3044, g3045, g3046, g3047, g3048, g3049, g3050, g3051, g3052, g3053, g3055, g3056, g3057, g3058, g3059, g3060, g3061, g3062, g3063, g3064, g3065, g3066, g3067, g3068, g3069, g3070, g3071, g3072, g3073, g3074, g3075, g3076, g3077, g3078, g2997, g2993, g2998, g3006, g3002, g3013, g3010, g3024, g3018, g3028, g3036, g3032, g3040, g2986, g2987, g3083, g2992, g2990, g2991, g3993, g4088, g4090, g4200, g4321, g4323, g4450, g4590, g5388, g5437, g5472, g5511, g5549, g5555, g5595, g5612, g5629, g5637, g5648, g5657, g5686, g5695, g5738, g5747, g5796, g6225, g6231, g6313, g6368, g6442, g6447, g6485, g6518, g6573, g6642, g6677, g6712, g6750, g6782, g6837, g6895, g6911, g6944, g6979, g7014, g7052, g7084, g7161, g7194, g7229, g7264, g7302, g7334, g7357, g7390, g7425, g7487, g7519, g7909, g7956, g7961, g8007, g8012, g8021, g8023, g8030, g8082, g8087, g8096, g8106, g8167, g8175, g8249, g8251, g8258, g8259, g8260, g8261, g8262, g8263, g8264, g8265, g8266, g8267, g8268, g8269, g8270, g8271, g8272, g8273, g8274, g8275, g16297, g16355, g16399, g16437, g16496, g24734, g25420, g25435, g25442, g25489, g26104, g26135, g26149, g27380, n269, n274, n279, n284, n289, n294, n299, n304, n309, n314, n319, n324, n329, n334, n339, n344, n349, n354, n358, n363, n368, n373, n378, n383, n388, n393, n398, n403, n408, n413, n418, n423, n428, n433, n438, n443, n448, n453, n458, n463, n468, n473, n478, n483, n488, n493, n498, n503, n507, n512, n516, n521, n525, n530, n534, n539, n543, n548, n552, n557, n561, n566, n570, n575, n579, n584, n588, n593, n597, n602, n606, n611, n615, n620, n624, n629, n633, n638, n642, n647, n651, n656, n660, n665, n670, n675, n680, n685, n690, n695, n700, n705, n710, n714, n718, n723, n728, n733, n738, n743, n748, n753, n758, n763, n768, n773, n778, n783, n788, n793, n798, n803, n808, n813, n818, n823, n828, n833, n838, n843, n848, n853, n858, n863, n868, n873, n878, n883, n888, n893, n898, n903, n908, n913, n918, n923, n928, n933, n938, n943, n948, n953, n958, n963, n968, n973, n978, n983, n988, n993, n998, n1003, n1008, n1013, n1018, n1023, n1028, n1033, n1038, n1043, n1048, n1053, n1057, n1061, n1066, n1071, n1076, n1081, n1086, n1091, n1096, n1101, n1106, n1111, n1116, n1121, n1126, n1131, n1136, n1141, n1146, n1151, n1156, n1161, n1166, n1171, n1176, n1181, n1186, n1191, n1196, n1201, n1206, n1211, n1216, n1221, n1226, n1231, n1236, n1241, n1246, n1251, n1256, n1261, n1266, n1271, n1276, n1281, n1286, n1291, n1296, n1301, n1306, n1311, n1316, n1321, n1326, n1331, n1336, n1341, n1346, n1351, n1356, n1361, n1366, n1371, n1376, n1381, n1386, n1391, n1396, n1401, n1406, n1411, n1416, n1421, n1426, n1431, n1436, n1441, n1446, n1451, n1456, n1461, n1466, n1471, n1476, n1480, n1484, n1489, n1493, n1497, n1502, n1507, n1512, n1517, n1522, n1527, n1532, n1537, n1542, n1547, n1552, n1557, n1562, n1567, n1572, n1577, n1582, n1587, n1592, n1597, n1602, n1607, n1612, n1617, n1622, n1627, n1632, n1637, n1642, n1647, n1652, n1657, n1662, n1667, n1672, n1677, n1682, n1687, n1692, n1697, n1702, n1707, n1712, n1717, n1722, n1727, n1732, n1736, n1741, n1745, n1750, n1754, n1759, n1763, n1768, n1772, n1777, n1781, n1786, n1790, n1795, n1799, n1804, n1808, n1813, n1818, n1823, n1828, n1833, n1838, n1843, n1848, n1853, n1858, n1863, n1868, n1873, n1878, n1882, n1887, n1891, n1896, n1900, n1905, n1909, n1914, n1918, n1923, n1927, n1932, n1936, n1941, n1945, n1950, n1954, n1959, n1963, n1968, n1972, n1977, n1981, n1986, n1990, n1994, n1999, n2003, n2007, n2012, n2017, n2022, n2027, n2031, n2035, n2040, n2044, n2049, n2053, n2058, n2062, n2067, n2071, n2076, n2080, n2085, n2089, n2094, n2098, n2102, n2107, n2112, n2117, n2122, n2127, n2132, n2137, n2142, n2147, n2152, n2157, n2162, n2167, n2172, n2177, n2182, n2186, n2190, n2195, n2199, n2204, n2209, n2213, n2218, n2222, n2227, n2232, n2237, n2242, n2247, n2252, n2257, n2262, n2267, n2272, n2277, n2282, n2287, n2292, n2297, n2302, n2307, n2312, n2317, n2322, n2327, n2332, n2337, n2342, n2347, n2352, n2357, n2362, n2367, n2372, n2377, n2382, n2387, n2392, n2397, n2402, n2407, n2412, n2416, n2421, n2426, n2431, n2436, n2441, n2446, n2451, n2456, n2461, n2466, n2471, n2475, n2479, n2484, n2489, n2494, n2499, n2504, n2509, n2514, n2519, n2524, n2529, n2534, n2539, n2544, n2549, n2554, n2559, n2564, n2569, n2574, n2579, n2584, n2589, n2594, n2599, n2604, n2609, n2614, n2619, n2624, n2629, n2634, n2639, n2644, n2649, n2654, n2659, n2664, n2669, n2674, n2679, n2684, n2689, n2694, n2699, n2704, n2709, n2714, n2719, n2724, n2729, n2734, n2739, n2744, n2749, n2754, n2758, n2762, n2767, n2772, n2777, n2782, n2787, n2792, n2797, n2802, n2807, n2812, n2817, n2822, n2827, n2832, n2837, n2842, n2847, n2852, n2857, n2862, n2867, n2872, n2877, n2882, n2887, n2892, n2897, n2902, n2907, n2912, n2917, n2922, n2927, n2932, n2937, n2942, n2947, n2952, n2957, n2962, n2967, n2972, n2977, n2982, n2987, n2992, n2997, n3002, n3007, n3012, n3017, n3022, n3027, n3032, n3037, n3042, n3047, n3052, n3057, n3062, n3067, n3072, n3077, n3082, n3087, n3092, n3097, n3102, n3107, n3112, n3117, n3122, n3127, n3132, n3137, n3142, n3147, n3152, n3157, n3162, n3167, n3172, n3177, n3181, n3185, n3190, n3194, n3198, n3203, n3208, n3213, n3218, n3223, n3228, n3233, n3238, n3243, n3248, n3253, n3258, n3263, n3268, n3273, n3278, n3283, n3288, n3293, n3298, n3303, n3308, n3313, n3318, n3323, n3328, n3333, n3338, n3343, n3348, n3353, n3358, n3363, n3368, n3373, n3378, n3383, n3388, n3393, n3398, n3403, n3408, n3413, n3418, n3423, n3428, n3433, n3437, n3442, n3446, n3451, n3455, n3460, n3464, n3469, n3473, n3478, n3482, n3487, n3491, n3496, n3500, n3505, n3509, n3514, n3519, n3524, n3529, n3534, n3539, n3544, n3549, n3554, n3559, n3564, n3569, n3574, n3579, n3583, n3588, n3592, n3597, n3601, n3606, n3610, n3615, n3619, n3624, n3628, n3633, n3637, n3642, n3646, n3651, n3655, n3660, n3664, n3669, n3673, n3678, n3682, n3687, n3691, n3695, n3700, n3704, n3708, n3713, n3718, n3723, n3728, n3732, n3736, n3741, n3745, n3750, n3754, n3759, n3763, n3768, n3772, n3777, n3781, n3786, n3790, n3795, n3799, n3803, n3808, n3813, n3818, n3823, n3828, n3833, n3838, n3843, n3848, n3853, n3858, n3863, n3868, n3873, n3878, n3883, n3887, n3891, n3896, n3900, n3905, n3910, n3914, n3919, n3923, n3928, n3933, n3938, n3943, n3948, n3953, n3958, n3963, n3968, n3973, n3978, n3983, n3988, n3993, n3998, n4003, n4008, n4013, n4018, n4023, n4028, n4033, n4038, n4043, n4048, n4053, n4058, n4063, n4068, n4073, n4078, n4083, n4088, n4093, n4098, n4103, n4108, n4113, n4117, n4122, n4127, n4132, n4137, n4142, n4147, n4152, n4157, n4162, n4167, n4172, n4176, n4180, n4185, n4190, n4195, n4200, n4205, n4210, n4215, n4220, n4225, n4230, n4235, n4240, n4245, n4250, n4255, n4260, n4265, n4270, n4275, n4280, n4285, n4290, n4295, n4300, n4305, n4310, n4315, n4320, n4325, n4330, n4335, n4340, n4345, n4350, n4355, n4360, n4365, n4370, n4375, n4380, n4385, n4390, n4395, n4400, n4405, n4410, n4415, n4420, n4425, n4430, n4435, n4440, n4445, n4450, n4455, n4459, n4463, n4468, n4473, n4478, n4483, n4488, n4493, n4498, n4503, n4508, n4513, n4518, n4523, n4528, n4533, n4538, n4543, n4548, n4553, n4558, n4563, n4568, n4573, n4578, n4583, n4588, n4593, n4598, n4603, n4608, n4613, n4618, n4623, n4628, n4633, n4638, n4643, n4648, n4653, n4658, n4663, n4668, n4673, n4678, n4683, n4688, n4693, n4698, n4703, n4708, n4713, n4718, n4723, n4728, n4733, n4738, n4743, n4748, n4753, n4758, n4763, n4768, n4773, n4778, n4783, n4788, n4793, n4798, n4803, n4808, n4813, n4818, n4823, n4828, n4833, n4838, n4843, n4848, n4853, n4858, n4863, n4868, n4873, n4878, n4882, n4886, n4891, n4895, n4899, n4904, n4909, n4914, n4919, n4924, n4929, n4934, n4939, n4944, n4949, n4954, n4959, n4964, n4969, n4974, n4979, n4984, n4989, n4994, n4999, n5004, n5009, n5014, n5019, n5024, n5029, n5034, n5039, n5044, n5049, n5054, n5059, n5064, n5069, n5074, n5079, n5084, n5089, n5094, n5099, n5104, n5109, n5114, n5119, n5124, n5129, n5134, n5138, n5143, n5147, n5152, n5156, n5161, n5165, n5170, n5174, n5179, n5183, n5188, n5192, n5197, n5201, n5206, n5210, n5215, n5220, n5225, n5230, n5235, n5240, n5245, n5250, n5255, n5260, n5265, n5270, n5275, n5280, n5284, n5289, n5293, n5298, n5302, n5307, n5311, n5316, n5320, n5325, n5329, n5334, n5338, n5343, n5347, n5352, n5356, n5361, n5365, n5370, n5374, n5379, n5383, n5388, n5392, n5396, n5401, n5405, n5409, n5414, n5419, n5424, n5429, n5433, n5437, n5442, n5446, n5451, n5455, n5460, n5464, n5469, n5473, n5478, n5482, n5487, n5491, n5496, n5500, n5504, n5509, n5514, n5519, n5524, n5529, n5534, n5539, n5544, n5549, n5554, n5559, n5564, n5569, n5574, n5579, n5584, n5588, n5592, n5597, n5601, n5606, n5611, n5615, n5620, n5624, n5629, n5634, n5639, n5644, n5649, n5654, n5659, n5664, n5669, n5674, n5679, n5684, n5689, n5694, n5699, n5704, n5709, n5714, n5719, n5724, n5729, n5734, n5739, n5744, n5749, n5754, n5759, n5764, n5769, n5774, n5779, n5784, n5789, n5794, n5799, n5804, n5809, n5814, n5818, n5823, n5828, n5833, n5838, n5843, n5848, n5853, n5858, n5863, n5868, n5873, n5877, n5881, n5886, n5891, n5896, n5901, n5906, n5911, n5916, n5921, n5926, n5931, n5936, n5941, n5946, n5951, n5956, n5961, n5966, n5971, n5976, n5981, n5986, n5991, n5996, n6001, n6006, n6011, n6016, n6021, n6026, n6031, n6036, n6041, n6046, n6051, n6056, n6061, n6066, n6071, n6076, n6081, n6086, n6091, n6096, n6101, n6106, n6111, n6116, n6121, n6126, n6131, n6136, n6141, n6146, n6151, n6156, n6160, n6164, n6169, n6174, n6179, n6184, n6189, n6194, n6199, n6204, n6209, n6214, n6219, n6224, n6229, n6234, n6239, n6244, n6249, n6254, n6259, n6264, n6269, n6274, n6279, n6284, n6289, n6294, n6299, n6304, n6309, n6314, n6319, n6324, n6329, n6334, n6339, n6344, n6349, n6354, n6359, n6364, n6369, n6374, n6379, n6384, n6389, n6394, n6399, n6404, n6409, n6414, n6419, n6424, n6429, n6434, n6439, n6444, n6449, n6454, n6459, n6464, n6469, n6474, n6479, n6484, n6489, n6494, n6499, n6504, n6509, n6514, n6519, n6524, n6529, n6534, n6539, n6544, n6549, n6554, n6559, n6564, n6569, n6574, n6579, n6583, n6587, n6592, n6596, n6600, n6605, n6610, n6615, n6620, n6625, n6630, n6635, n6640, n6645, n6650, n6655, n6660, n6665, n6670, n6675, n6680, n6685, n6690, n6695, n6700, n6705, n6710, n6715, n6720, n6725, n6730, n6735, n6740, n6745, n6750, n6755, n6760, n6765, n6770, n6775, n6780, n6785, n6790, n6795, n6800, n6805, n6810, n6815, n6820, n6825, n6830, n6835, n6839, n6844, n6848, n6853, n6857, n6862, n6866, n6871, n6875, n6880, n6884, n6889, n6893, n6898, n6902, n6907, n6911, n6916, n6921, n6926, n6931, n6936, n6941, n6946, n6951, n6956, n6961, n6966, n6971, n6976, n6981, n6985, n6990, n6994, n6999, n7003, n7008, n7012, n7017, n7021, n7026, n7030, n7035, n7039, n7044, n7048, n7053, n7057, n7062, n7066, n7071, n7075, n7080, n7084, n7089, n7093, n7097, n7102, n7106, n7110, n7115, n7120, n7125, n7130, n7134, n7138, n7143, n7147, n7152, n7156, n7161, n7165, n7170, n7174, n7179, n7183, n7188, n7192, n7197, n7201, n7205, n7210, n7215, n7220, n7225, n7230, n7235, n7240, n7245, n7250, n7255, n7260, n7265, n7270, n7275, n7280, n7285, n7289, n7293, n7298, n7302, n7307, n7312, n7316, n7321, n7325, n7330, n7335, n7340, n7345, n7350, n7355, n7360, n7365, n7370, n7375, n7380, n7385, n7390, n7395, n7400, n7405, n7410, n7415, n7420, n7425, n7430, n7435, n7440, n7445, n7450, n7455, n7460, n7465, n7470, n7475, n7480, n7485, n7490, n7495, n7500, n7505, n7510, n7515, n7519, n7524, n7529, n7534, n7539, n7544, n7549, n7554, n7559, n7564, n7569, n7574, n7578, n7582, n7587, n7592, n7597, n7602, n7607, n7612, n7617, n7622, n7627, n7632, n7637, n7642, n7647, n7652, n7657, n7662, n7667, n7672, n7677, n7682, n7687, n7692, n7697, n7702, n7707, n7712, n7717, n7722, n7727, n7732, n7737, n7742, n7747, n7752, n7757, n7762, n7767, n7772, n7777, n7782, n7787, n7792, n7797, n7802, n7807, n7812, n7817, n7822, n7827, n7832, n7837, n7842, n7847, n7852, n7857, n7862, n7867, n7872, n7877, n7882, n7887, n7892, n7897, n7902, n7907, n7912, n7917, n7922, n7927, n7932, n7937, n7942, n7947, n7952, n7957, n7962, n7967, n7972, n7977, n7982, n7987, n7992, n7997, n8002, n8007, n8012, n8017, n8022, n8027, n8032, n8037, n8042, n8047, n8052, n8057, n8062, n8067, n8072, n8077, n8082, n8087, n8092, n8097, n8102, n8107, n8111, n8116, n8121, n8126, n8131, n8136, n8141, n8146, n8151, n8156, n8161, n8166, n8171, n8176, n8181, n8186, n8191, n8196, n8201, n8206, n8211, n8216, n8221, n8226 );
input g290, g288, g286, g284, g282, g26, g1, g23, g20, g17, g11, g14, g5, g2, g8, g48, g45, g42, g39, g27, g30, g33, g36, g291, g289, g287, g285, g283, g281, g294, g295, g296, g297, g308, g298, g309, g56, g79, g321, g323, g322, g314, g313, g312, g317, g316, g315, g320, g319, g318, g219, g216, g150, g147, g149, g148, g51, g563, g1249, g1943, g2637, g3212, g3213, g3214, g3215, g3216, g3217, g3218, g3219, g3220, g3221, g3222, g3223, g3224, g3225, g3226, g3227, g3228, g3229, g3230, g3231, g3232, g3233, g3234, g2814, g2817, g2933, g2950, g2883, g2888, g2896, g2892, g2903, g2900, g2908, g2912, g2917, g2924, g2920, g2984, g2985, g2930, g2929, g2879, g2934, g2935, g2938, g2941, g2944, g2947, g2953, g2956, g2959, g2962, g2963, g2966, g2969, g2972, g2975, g2978, g2981, g2874, g1506, g1501, g1496, g1491, g1486, g1481, g1476, g1471, g2877, g2861, g813, g2864, g809, g2867, g805, g2870, g801, g2818, g797, g2821, g793, g2824, g789, g2827, g785, g2830, g2873, g2833, g125, g2836, g121, g2839, g117, g2842, g113, g2845, g109, g2848, g105, g2851, g101, g2854, g97, g2858, g2857, g2200, g2195, g2190, g2185, g2180, g2175, g2170, g2165, g2878, g3129, g3117, g3109, g3210, g3211, g3084, g3085, g3086, g3087, g3091, g3092, g3093, g3094, g3095, g3096, g3097, g3098, g3099, g3100, g3101, g3102, g3103, g3104, g3105, g3106, g3107, g3108, g3155, g3158, g3161, g3164, g3167, g3170, g3173, g3176, g3179, g3182, g3185, g3088, g3191, g3194, g3197, g3198, g3201, g3204, g3207, g3188, g3133, g3132, g3128, g3127, g3126, g3125, g3124, g3123, g3120, g3114, g3113, g3112, g3110, g3111, g3139, g3136, g3134, g3135, g3151, g3142, g3147, g185, g138, g135, g165, g130, g131, g129, g133, g134, g132, g142, g143, g141, g145, g146, g144, g151, g152, g154, g155, g153, g157, g158, g156, g160, g161, g159, g163, g164, g162, g169, g170, g168, g172, g173, g171, g175, g176, g174, g178, g179, g177, g186, g189, g192, g231, g234, g237, g195, g198, g201, g240, g243, g246, g204, g207, g210, g249, g252, g255, g213, g258, g261, g264, g222, g225, g228, g267, g270, g273, g92, g88, g83, g74, g70, g65, g61, g52, g180, g182, g181, g276, g405, g401, g354, g343, g346, g369, g358, g361, g384, g373, g376, g398, g388, g391, g408, g411, g414, g417, g420, g423, g427, g428, g426, g429, g432, g435, g438, g441, g444, g448, g449, g447, g403, g404, g402, g450, g451, g452, g453, g454, g279, g280, g299, g305, g304, g303, g302, g301, g300, g342, g349, g350, g351, g352, g353, g357, g364, g365, g366, g367, g368, g372, g379, g380, g381, g382, g383, g387, g394, g395, g396, g397, g324, g325, g331, g337, g545, g551, g550, g554, g557, g510, g513, g523, g524, g564, g569, g570, g571, g572, g573, g574, g565, g566, g567, g568, g489, g474, g481, g485, g486, g487, g488, g455, g458, g461, g477, g478, g479, g480, g484, g464, g465, g468, g471, g528, g535, g542, g543, g544, g548, g549, g499, g558, g559, g576, g577, g575, g579, g580, g578, g582, g583, g581, g585, g586, g584, g587, g590, g593, g596, g599, g602, g614, g617, g620, g605, g608, g611, g490, g493, g496, g506, g507, g508, g509, g514, g515, g516, g517, g518, g519, g520, g525, g529, g530, g531, g532, g533, g534, g536, g537, g538, g541, g623, g626, g629, g630, g659, g640, g633, g653, g646, g660, g672, g666, g679, g686, g692, g699, g700, g698, g702, g703, g701, g705, g706, g704, g708, g709, g707, g711, g712, g710, g714, g715, g713, g717, g718, g716, g720, g721, g719, g723, g724, g722, g726, g727, g725, g729, g730, g728, g732, g733, g731, g735, g736, g734, g738, g739, g737, g826, g823, g853, g818, g819, g817, g821, g822, g820, g830, g831, g829, g833, g834, g832, g836, g837, g835, g839, g840, g838, g842, g843, g841, g845, g846, g844, g848, g849, g847, g851, g852, g850, g857, g858, g856, g860, g861, g859, g863, g864, g862, g866, g867, g865, g873, g876, g879, g918, g921, g924, g882, g885, g888, g927, g930, g933, g891, g894, g897, g936, g939, g942, g900, g903, g906, g945, g948, g951, g909, g912, g915, g954, g957, g960, g780, g776, g771, g767, g762, g758, g753, g749, g744, g740, g868, g870, g869, g963, g1092, g1088, g996, g1041, g1030, g1033, g1056, g1045, g1048, g1071, g1060, g1063, g1085, g1075, g1078, g1095, g1098, g1101, g1104, g1107, g1110, g1114, g1115, g1113, g1116, g1119, g1122, g1125, g1128, g1131, g1135, g1136, g1134, g999, g1000, g1001, g1002, g1003, g1004, g1005, g1006, g1007, g1009, g1010, g1008, g1090, g1091, g1089, g1137, g1138, g1139, g1140, g1141, g966, g967, g968, g969, g970, g971, g972, g973, g974, g975, g976, g977, g978, g986, g992, g995, g984, g983, g982, g981, g991, g990, g989, g988, g987, g985, g1029, g1036, g1037, g1038, g1039, g1040, g1044, g1051, g1052, g1053, g1054, g1055, g1059, g1066, g1067, g1068, g1069, g1070, g1074, g1081, g1082, g1083, g1084, g1011, g1012, g1018, g1024, g1231, g1237, g1236, g1240, g1243, g1196, g1199, g1209, g1210, g1250, g1255, g1256, g1257, g1258, g1259, g1260, g1251, g1252, g1253, g1254, g1176, g1161, g1168, g1172, g1173, g1174, g1175, g1142, g1145, g1148, g1164, g1165, g1166, g1167, g1171, g1151, g1152, g1155, g1158, g1214, g1221, g1228, g1229, g1230, g1234, g1235, g1186, g1244, g1245, g1262, g1263, g1261, g1265, g1266, g1264, g1268, g1269, g1267, g1271, g1272, g1270, g1273, g1276, g1279, g1282, g1285, g1288, g1300, g1303, g1306, g1291, g1294, g1297, g1177, g1180, g1183, g1192, g1193, g1194, g1195, g1200, g1201, g1202, g1203, g1204, g1205, g1206, g1211, g1215, g1216, g1217, g1218, g1219, g1220, g1222, g1223, g1224, g1227, g1309, g1312, g1315, g1316, g1345, g1326, g1319, g1339, g1332, g1346, g1358, g1352, g1365, g1372, g1378, g1385, g1386, g1384, g1388, g1389, g1387, g1391, g1392, g1390, g1394, g1395, g1393, g1397, g1398, g1396, g1400, g1401, g1399, g1403, g1404, g1402, g1406, g1407, g1405, g1409, g1410, g1408, g1412, g1413, g1411, g1415, g1416, g1414, g1418, g1419, g1417, g1421, g1422, g1420, g1424, g1425, g1423, g1520, g1517, g1547, g1512, g1513, g1511, g1515, g1516, g1514, g1524, g1525, g1523, g1527, g1528, g1526, g1530, g1531, g1529, g1533, g1534, g1532, g1536, g1537, g1535, g1539, g1540, g1538, g1542, g1543, g1541, g1545, g1546, g1544, g1551, g1552, g1550, g1554, g1555, g1553, g1557, g1558, g1556, g1560, g1561, g1559, g1567, g1570, g1573, g1612, g1615, g1618, g1576, g1579, g1582, g1621, g1624, g1627, g1585, g1588, g1591, g1630, g1633, g1636, g1594, g1597, g1600, g1639, g1642, g1645, g1603, g1606, g1609, g1648, g1651, g1654, g1466, g1462, g1457, g1453, g1448, g1444, g1439, g1435, g1430, g1426, g1562, g1564, g1563, g1657, g1786, g1782, g1690, g1735, g1724, g1727, g1750, g1739, g1742, g1765, g1754, g1757, g1779, g1769, g1772, g1789, g1792, g1795, g1798, g1801, g1804, g1808, g1809, g1807, g1810, g1813, g1816, g1819, g1822, g1825, g1829, g1830, g1828, g1693, g1694, g1695, g1696, g1697, g1698, g1699, g1700, g1701, g1703, g1704, g1702, g1784, g1785, g1783, g1831, g1832, g1833, g1834, g1835, g1660, g1661, g1662, g1663, g1664, g1665, g1666, g1667, g1668, g1669, g1670, g1671, g1672, g1680, g1686, g1689, g1678, g1677, g1676, g1675, g1685, g1684, g1683, g1682, g1681, g1679, g1723, g1730, g1731, g1732, g1733, g1734, g1738, g1745, g1746, g1747, g1748, g1749, g1753, g1760, g1761, g1762, g1763, g1764, g1768, g1775, g1776, g1777, g1778, g1705, g1706, g1712, g1718, g1925, g1931, g1930, g1934, g1937, g1890, g1893, g1903, g1904, g1944, g1949, g1950, g1951, g1952, g1953, g1954, g1945, g1946, g1947, g1948, g1870, g1855, g1862, g1866, g1867, g1868, g1869, g1836, g1839, g1842, g1858, g1859, g1860, g1861, g1865, g1845, g1846, g1849, g1852, g1908, g1915, g1922, g1923, g1924, g1928, g1929, g1880, g1938, g1939, g1956, g1957, g1955, g1959, g1960, g1958, g1962, g1963, g1961, g1965, g1966, g1964, g1967, g1970, g1973, g1976, g1979, g1982, g1994, g1997, g2000, g1985, g1988, g1991, g1871, g1874, g1877, g1886, g1887, g1888, g1889, g1894, g1895, g1896, g1897, g1898, g1899, g1900, g1905, g1909, g1910, g1911, g1912, g1913, g1914, g1916, g1917, g1918, g1921, g2003, g2006, g2009, g2010, g2039, g2020, g2013, g2033, g2026, g2040, g2052, g2046, g2059, g2066, g2072, g2079, g2080, g2078, g2082, g2083, g2081, g2085, g2086, g2084, g2088, g2089, g2087, g2091, g2092, g2090, g2094, g2095, g2093, g2097, g2098, g2096, g2100, g2101, g2099, g2103, g2104, g2102, g2106, g2107, g2105, g2109, g2110, g2108, g2112, g2113, g2111, g2115, g2116, g2114, g2118, g2119, g2117, g2214, g2211, g2241, g2206, g2207, g2205, g2209, g2210, g2208, g2218, g2219, g2217, g2221, g2222, g2220, g2224, g2225, g2223, g2227, g2228, g2226, g2230, g2231, g2229, g2233, g2234, g2232, g2236, g2237, g2235, g2239, g2240, g2238, g2245, g2246, g2244, g2248, g2249, g2247, g2251, g2252, g2250, g2254, g2255, g2253, g2261, g2264, g2267, g2306, g2309, g2312, g2270, g2273, g2276, g2315, g2318, g2321, g2279, g2282, g2285, g2324, g2327, g2330, g2288, g2291, g2294, g2333, g2336, g2339, g2297, g2300, g2303, g2342, g2345, g2348, g2160, g2156, g2151, g2147, g2142, g2138, g2133, g2129, g2124, g2120, g2256, g2258, g2257, g2351, g2480, g2476, g2384, g2429, g2418, g2421, g2444, g2433, g2436, g2459, g2448, g2451, g2473, g2463, g2466, g2483, g2486, g2489, g2492, g2495, g2498, g2502, g2503, g2501, g2504, g2507, g2510, g2513, g2516, g2519, g2523, g2524, g2522, g2387, g2388, g2389, g2390, g2391, g2392, g2393, g2394, g2395, g2397, g2398, g2396, g2478, g2479, g2477, g2525, g2526, g2527, g2528, g2529, g2354, g2355, g2356, g2357, g2358, g2359, g2360, g2361, g2362, g2363, g2364, g2365, g2366, g2374, g2380, g2383, g2372, g2371, g2370, g2369, g2379, g2378, g2377, g2376, g2375, g2373, g2417, g2424, g2425, g2426, g2427, g2428, g2432, g2439, g2440, g2441, g2442, g2443, g2447, g2454, g2455, g2456, g2457, g2458, g2462, g2469, g2470, g2471, g2472, g2399, g2400, g2406, g2412, g2619, g2625, g2624, g2628, g2631, g2584, g2587, g2597, g2598, g2638, g2643, g2644, g2645, g2646, g2647, g2648, g2639, g2640, g2641, g2642, g2564, g2549, g2556, g2560, g2561, g2562, g2563, g2530, g2533, g2536, g2552, g2553, g2554, g2555, g2559, g2539, g2540, g2543, g2546, g2602, g2609, g2616, g2617, g2618, g2622, g2623, g2574, g2632, g2633, g2650, g2651, g2649, g2653, g2654, g2652, g2656, g2657, g2655, g2659, g2660, g2658, g2661, g2664, g2667, g2670, g2673, g2676, g2688, g2691, g2694, g2679, g2682, g2685, g2565, g2568, g2571, g2580, g2581, g2582, g2583, g2588, g2589, g2590, g2591, g2592, g2593, g2594, g2599, g2603, g2604, g2605, g2606, g2607, g2608, g2610, g2611, g2612, g2615, g2697, g2700, g2703, g2704, g2733, g2714, g2707, g2727, g2720, g2734, g2746, g2740, g2753, g2760, g2766, g2773, g2774, g2772, g2776, g2777, g2775, g2779, g2780, g2778, g2782, g2783, g2781, g2785, g2786, g2784, g2788, g2789, g2787, g2791, g2792, g2790, g2794, g2795, g2793, g2797, g2798, g2796, g2800, g2801, g2799, g2803, g2804, g2802, g2806, g2807, g2805, g2809, g2810, g2808, g2812, g2813, g2811, g3054, g3079, g3080, g3043, g3044, g3045, g3046, g3047, g3048, g3049, g3050, g3051, g3052, g3053, g3055, g3056, g3057, g3058, g3059, g3060, g3061, g3062, g3063, g3064, g3065, g3066, g3067, g3068, g3069, g3070, g3071, g3072, g3073, g3074, g3075, g3076, g3077, g3078, g2997, g2993, g2998, g3006, g3002, g3013, g3010, g3024, g3018, g3028, g3036, g3032, g3040, g2986, g2987, g3083, g2992, g2990, g2991;
output g3993, g4088, g4090, g4200, g4321, g4323, g4450, g4590, g5388, g5437, g5472, g5511, g5549, g5555, g5595, g5612, g5629, g5637, g5648, g5657, g5686, g5695, g5738, g5747, g5796, g6225, g6231, g6313, g6368, g6442, g6447, g6485, g6518, g6573, g6642, g6677, g6712, g6750, g6782, g6837, g6895, g6911, g6944, g6979, g7014, g7052, g7084, g7161, g7194, g7229, g7264, g7302, g7334, g7357, g7390, g7425, g7487, g7519, g7909, g7956, g7961, g8007, g8012, g8021, g8023, g8030, g8082, g8087, g8096, g8106, g8167, g8175, g8249, g8251, g8258, g8259, g8260, g8261, g8262, g8263, g8264, g8265, g8266, g8267, g8268, g8269, g8270, g8271, g8272, g8273, g8274, g8275, g16297, g16355, g16399, g16437, g16496, g24734, g25420, g25435, g25442, g25489, g26104, g26135, g26149, g27380, n269, n274, n279, n284, n289, n294, n299, n304, n309, n314, n319, n324, n329, n334, n339, n344, n349, n354, n358, n363, n368, n373, n378, n383, n388, n393, n398, n403, n408, n413, n418, n423, n428, n433, n438, n443, n448, n453, n458, n463, n468, n473, n478, n483, n488, n493, n498, n503, n507, n512, n516, n521, n525, n530, n534, n539, n543, n548, n552, n557, n561, n566, n570, n575, n579, n584, n588, n593, n597, n602, n606, n611, n615, n620, n624, n629, n633, n638, n642, n647, n651, n656, n660, n665, n670, n675, n680, n685, n690, n695, n700, n705, n710, n714, n718, n723, n728, n733, n738, n743, n748, n753, n758, n763, n768, n773, n778, n783, n788, n793, n798, n803, n808, n813, n818, n823, n828, n833, n838, n843, n848, n853, n858, n863, n868, n873, n878, n883, n888, n893, n898, n903, n908, n913, n918, n923, n928, n933, n938, n943, n948, n953, n958, n963, n968, n973, n978, n983, n988, n993, n998, n1003, n1008, n1013, n1018, n1023, n1028, n1033, n1038, n1043, n1048, n1053, n1057, n1061, n1066, n1071, n1076, n1081, n1086, n1091, n1096, n1101, n1106, n1111, n1116, n1121, n1126, n1131, n1136, n1141, n1146, n1151, n1156, n1161, n1166, n1171, n1176, n1181, n1186, n1191, n1196, n1201, n1206, n1211, n1216, n1221, n1226, n1231, n1236, n1241, n1246, n1251, n1256, n1261, n1266, n1271, n1276, n1281, n1286, n1291, n1296, n1301, n1306, n1311, n1316, n1321, n1326, n1331, n1336, n1341, n1346, n1351, n1356, n1361, n1366, n1371, n1376, n1381, n1386, n1391, n1396, n1401, n1406, n1411, n1416, n1421, n1426, n1431, n1436, n1441, n1446, n1451, n1456, n1461, n1466, n1471, n1476, n1480, n1484, n1489, n1493, n1497, n1502, n1507, n1512, n1517, n1522, n1527, n1532, n1537, n1542, n1547, n1552, n1557, n1562, n1567, n1572, n1577, n1582, n1587, n1592, n1597, n1602, n1607, n1612, n1617, n1622, n1627, n1632, n1637, n1642, n1647, n1652, n1657, n1662, n1667, n1672, n1677, n1682, n1687, n1692, n1697, n1702, n1707, n1712, n1717, n1722, n1727, n1732, n1736, n1741, n1745, n1750, n1754, n1759, n1763, n1768, n1772, n1777, n1781, n1786, n1790, n1795, n1799, n1804, n1808, n1813, n1818, n1823, n1828, n1833, n1838, n1843, n1848, n1853, n1858, n1863, n1868, n1873, n1878, n1882, n1887, n1891, n1896, n1900, n1905, n1909, n1914, n1918, n1923, n1927, n1932, n1936, n1941, n1945, n1950, n1954, n1959, n1963, n1968, n1972, n1977, n1981, n1986, n1990, n1994, n1999, n2003, n2007, n2012, n2017, n2022, n2027, n2031, n2035, n2040, n2044, n2049, n2053, n2058, n2062, n2067, n2071, n2076, n2080, n2085, n2089, n2094, n2098, n2102, n2107, n2112, n2117, n2122, n2127, n2132, n2137, n2142, n2147, n2152, n2157, n2162, n2167, n2172, n2177, n2182, n2186, n2190, n2195, n2199, n2204, n2209, n2213, n2218, n2222, n2227, n2232, n2237, n2242, n2247, n2252, n2257, n2262, n2267, n2272, n2277, n2282, n2287, n2292, n2297, n2302, n2307, n2312, n2317, n2322, n2327, n2332, n2337, n2342, n2347, n2352, n2357, n2362, n2367, n2372, n2377, n2382, n2387, n2392, n2397, n2402, n2407, n2412, n2416, n2421, n2426, n2431, n2436, n2441, n2446, n2451, n2456, n2461, n2466, n2471, n2475, n2479, n2484, n2489, n2494, n2499, n2504, n2509, n2514, n2519, n2524, n2529, n2534, n2539, n2544, n2549, n2554, n2559, n2564, n2569, n2574, n2579, n2584, n2589, n2594, n2599, n2604, n2609, n2614, n2619, n2624, n2629, n2634, n2639, n2644, n2649, n2654, n2659, n2664, n2669, n2674, n2679, n2684, n2689, n2694, n2699, n2704, n2709, n2714, n2719, n2724, n2729, n2734, n2739, n2744, n2749, n2754, n2758, n2762, n2767, n2772, n2777, n2782, n2787, n2792, n2797, n2802, n2807, n2812, n2817, n2822, n2827, n2832, n2837, n2842, n2847, n2852, n2857, n2862, n2867, n2872, n2877, n2882, n2887, n2892, n2897, n2902, n2907, n2912, n2917, n2922, n2927, n2932, n2937, n2942, n2947, n2952, n2957, n2962, n2967, n2972, n2977, n2982, n2987, n2992, n2997, n3002, n3007, n3012, n3017, n3022, n3027, n3032, n3037, n3042, n3047, n3052, n3057, n3062, n3067, n3072, n3077, n3082, n3087, n3092, n3097, n3102, n3107, n3112, n3117, n3122, n3127, n3132, n3137, n3142, n3147, n3152, n3157, n3162, n3167, n3172, n3177, n3181, n3185, n3190, n3194, n3198, n3203, n3208, n3213, n3218, n3223, n3228, n3233, n3238, n3243, n3248, n3253, n3258, n3263, n3268, n3273, n3278, n3283, n3288, n3293, n3298, n3303, n3308, n3313, n3318, n3323, n3328, n3333, n3338, n3343, n3348, n3353, n3358, n3363, n3368, n3373, n3378, n3383, n3388, n3393, n3398, n3403, n3408, n3413, n3418, n3423, n3428, n3433, n3437, n3442, n3446, n3451, n3455, n3460, n3464, n3469, n3473, n3478, n3482, n3487, n3491, n3496, n3500, n3505, n3509, n3514, n3519, n3524, n3529, n3534, n3539, n3544, n3549, n3554, n3559, n3564, n3569, n3574, n3579, n3583, n3588, n3592, n3597, n3601, n3606, n3610, n3615, n3619, n3624, n3628, n3633, n3637, n3642, n3646, n3651, n3655, n3660, n3664, n3669, n3673, n3678, n3682, n3687, n3691, n3695, n3700, n3704, n3708, n3713, n3718, n3723, n3728, n3732, n3736, n3741, n3745, n3750, n3754, n3759, n3763, n3768, n3772, n3777, n3781, n3786, n3790, n3795, n3799, n3803, n3808, n3813, n3818, n3823, n3828, n3833, n3838, n3843, n3848, n3853, n3858, n3863, n3868, n3873, n3878, n3883, n3887, n3891, n3896, n3900, n3905, n3910, n3914, n3919, n3923, n3928, n3933, n3938, n3943, n3948, n3953, n3958, n3963, n3968, n3973, n3978, n3983, n3988, n3993, n3998, n4003, n4008, n4013, n4018, n4023, n4028, n4033, n4038, n4043, n4048, n4053, n4058, n4063, n4068, n4073, n4078, n4083, n4088, n4093, n4098, n4103, n4108, n4113, n4117, n4122, n4127, n4132, n4137, n4142, n4147, n4152, n4157, n4162, n4167, n4172, n4176, n4180, n4185, n4190, n4195, n4200, n4205, n4210, n4215, n4220, n4225, n4230, n4235, n4240, n4245, n4250, n4255, n4260, n4265, n4270, n4275, n4280, n4285, n4290, n4295, n4300, n4305, n4310, n4315, n4320, n4325, n4330, n4335, n4340, n4345, n4350, n4355, n4360, n4365, n4370, n4375, n4380, n4385, n4390, n4395, n4400, n4405, n4410, n4415, n4420, n4425, n4430, n4435, n4440, n4445, n4450, n4455, n4459, n4463, n4468, n4473, n4478, n4483, n4488, n4493, n4498, n4503, n4508, n4513, n4518, n4523, n4528, n4533, n4538, n4543, n4548, n4553, n4558, n4563, n4568, n4573, n4578, n4583, n4588, n4593, n4598, n4603, n4608, n4613, n4618, n4623, n4628, n4633, n4638, n4643, n4648, n4653, n4658, n4663, n4668, n4673, n4678, n4683, n4688, n4693, n4698, n4703, n4708, n4713, n4718, n4723, n4728, n4733, n4738, n4743, n4748, n4753, n4758, n4763, n4768, n4773, n4778, n4783, n4788, n4793, n4798, n4803, n4808, n4813, n4818, n4823, n4828, n4833, n4838, n4843, n4848, n4853, n4858, n4863, n4868, n4873, n4878, n4882, n4886, n4891, n4895, n4899, n4904, n4909, n4914, n4919, n4924, n4929, n4934, n4939, n4944, n4949, n4954, n4959, n4964, n4969, n4974, n4979, n4984, n4989, n4994, n4999, n5004, n5009, n5014, n5019, n5024, n5029, n5034, n5039, n5044, n5049, n5054, n5059, n5064, n5069, n5074, n5079, n5084, n5089, n5094, n5099, n5104, n5109, n5114, n5119, n5124, n5129, n5134, n5138, n5143, n5147, n5152, n5156, n5161, n5165, n5170, n5174, n5179, n5183, n5188, n5192, n5197, n5201, n5206, n5210, n5215, n5220, n5225, n5230, n5235, n5240, n5245, n5250, n5255, n5260, n5265, n5270, n5275, n5280, n5284, n5289, n5293, n5298, n5302, n5307, n5311, n5316, n5320, n5325, n5329, n5334, n5338, n5343, n5347, n5352, n5356, n5361, n5365, n5370, n5374, n5379, n5383, n5388, n5392, n5396, n5401, n5405, n5409, n5414, n5419, n5424, n5429, n5433, n5437, n5442, n5446, n5451, n5455, n5460, n5464, n5469, n5473, n5478, n5482, n5487, n5491, n5496, n5500, n5504, n5509, n5514, n5519, n5524, n5529, n5534, n5539, n5544, n5549, n5554, n5559, n5564, n5569, n5574, n5579, n5584, n5588, n5592, n5597, n5601, n5606, n5611, n5615, n5620, n5624, n5629, n5634, n5639, n5644, n5649, n5654, n5659, n5664, n5669, n5674, n5679, n5684, n5689, n5694, n5699, n5704, n5709, n5714, n5719, n5724, n5729, n5734, n5739, n5744, n5749, n5754, n5759, n5764, n5769, n5774, n5779, n5784, n5789, n5794, n5799, n5804, n5809, n5814, n5818, n5823, n5828, n5833, n5838, n5843, n5848, n5853, n5858, n5863, n5868, n5873, n5877, n5881, n5886, n5891, n5896, n5901, n5906, n5911, n5916, n5921, n5926, n5931, n5936, n5941, n5946, n5951, n5956, n5961, n5966, n5971, n5976, n5981, n5986, n5991, n5996, n6001, n6006, n6011, n6016, n6021, n6026, n6031, n6036, n6041, n6046, n6051, n6056, n6061, n6066, n6071, n6076, n6081, n6086, n6091, n6096, n6101, n6106, n6111, n6116, n6121, n6126, n6131, n6136, n6141, n6146, n6151, n6156, n6160, n6164, n6169, n6174, n6179, n6184, n6189, n6194, n6199, n6204, n6209, n6214, n6219, n6224, n6229, n6234, n6239, n6244, n6249, n6254, n6259, n6264, n6269, n6274, n6279, n6284, n6289, n6294, n6299, n6304, n6309, n6314, n6319, n6324, n6329, n6334, n6339, n6344, n6349, n6354, n6359, n6364, n6369, n6374, n6379, n6384, n6389, n6394, n6399, n6404, n6409, n6414, n6419, n6424, n6429, n6434, n6439, n6444, n6449, n6454, n6459, n6464, n6469, n6474, n6479, n6484, n6489, n6494, n6499, n6504, n6509, n6514, n6519, n6524, n6529, n6534, n6539, n6544, n6549, n6554, n6559, n6564, n6569, n6574, n6579, n6583, n6587, n6592, n6596, n6600, n6605, n6610, n6615, n6620, n6625, n6630, n6635, n6640, n6645, n6650, n6655, n6660, n6665, n6670, n6675, n6680, n6685, n6690, n6695, n6700, n6705, n6710, n6715, n6720, n6725, n6730, n6735, n6740, n6745, n6750, n6755, n6760, n6765, n6770, n6775, n6780, n6785, n6790, n6795, n6800, n6805, n6810, n6815, n6820, n6825, n6830, n6835, n6839, n6844, n6848, n6853, n6857, n6862, n6866, n6871, n6875, n6880, n6884, n6889, n6893, n6898, n6902, n6907, n6911, n6916, n6921, n6926, n6931, n6936, n6941, n6946, n6951, n6956, n6961, n6966, n6971, n6976, n6981, n6985, n6990, n6994, n6999, n7003, n7008, n7012, n7017, n7021, n7026, n7030, n7035, n7039, n7044, n7048, n7053, n7057, n7062, n7066, n7071, n7075, n7080, n7084, n7089, n7093, n7097, n7102, n7106, n7110, n7115, n7120, n7125, n7130, n7134, n7138, n7143, n7147, n7152, n7156, n7161, n7165, n7170, n7174, n7179, n7183, n7188, n7192, n7197, n7201, n7205, n7210, n7215, n7220, n7225, n7230, n7235, n7240, n7245, n7250, n7255, n7260, n7265, n7270, n7275, n7280, n7285, n7289, n7293, n7298, n7302, n7307, n7312, n7316, n7321, n7325, n7330, n7335, n7340, n7345, n7350, n7355, n7360, n7365, n7370, n7375, n7380, n7385, n7390, n7395, n7400, n7405, n7410, n7415, n7420, n7425, n7430, n7435, n7440, n7445, n7450, n7455, n7460, n7465, n7470, n7475, n7480, n7485, n7490, n7495, n7500, n7505, n7510, n7515, n7519, n7524, n7529, n7534, n7539, n7544, n7549, n7554, n7559, n7564, n7569, n7574, n7578, n7582, n7587, n7592, n7597, n7602, n7607, n7612, n7617, n7622, n7627, n7632, n7637, n7642, n7647, n7652, n7657, n7662, n7667, n7672, n7677, n7682, n7687, n7692, n7697, n7702, n7707, n7712, n7717, n7722, n7727, n7732, n7737, n7742, n7747, n7752, n7757, n7762, n7767, n7772, n7777, n7782, n7787, n7792, n7797, n7802, n7807, n7812, n7817, n7822, n7827, n7832, n7837, n7842, n7847, n7852, n7857, n7862, n7867, n7872, n7877, n7882, n7887, n7892, n7897, n7902, n7907, n7912, n7917, n7922, n7927, n7932, n7937, n7942, n7947, n7952, n7957, n7962, n7967, n7972, n7977, n7982, n7987, n7992, n7997, n8002, n8007, n8012, n8017, n8022, n8027, n8032, n8037, n8042, n8047, n8052, n8057, n8062, n8067, n8072, n8077, n8082, n8087, n8092, n8097, n8102, n8107, n8111, n8116, n8121, n8126, n8131, n8136, n8141, n8146, n8151, n8156, n8161, n8166, n8171, n8176, n8181, n8186, n8191, n8196, n8201, n8206, n8211, n8216, n8221, n8226;
wire n5042, n5044_1, n5045, n5046, n5047, n5048, n5049_1, n5050, n5051, n5053, n5054_1, n5055, n5056, n5058, n5059_1, n5062, n5064_1, n5065, n5066, n5067, n5068, n5069_1, n5070, n5071, n5072, n5073, n5074_1, n5076, n5077, n5078, n5079_1, n5080, n5081, n5082, n5083, n5084_1, n5085, n5086, n5087, n5088, n5089_1, n5090, n5091, n5092, n5093, n5094_1, n5095, n5096, n5097, n5098, n5099_1, n5100, n5101, n5102, n5103, n5104_1, n5105, n5106, n5107, n5108, n5109_1, n5110, n5111, n5112, n5113, n5114_1, n5115, n5116, n5117, n5118, n5120, n5121, n5122, n5123, n5124_1, n5125, n5126, n5127, n5128, n5129_1, n5130, n5131, n5132, n5133, n5134_1, n5135, n5136, n5137, n5138_1, n5139, n5140, n5141, n5144, n5145, n5146, n5147_1, n5148, n5149, n5150, n5151, n5152_1, n5153, n5154, n5155, n5156_1, n5157, n5158, n5159, n5160, n5161_1, n5162, n5163, n5165_1, n5166, n5167, n5168, n5169, n5170_1, n5171, n5172, n5173, n5174_1, n5177, n5179_1, n5182, n5183_1, n5184, n5185, n5186, n5187, n5188_1, n5190, n5191, n5193, n5194, n5196, n5197_1, n5199, n5200, n5201_1, n5203, n5204, n5206_1, n5207, n5209, n5210_1, n5211, n5212, n5213, n5214, n5216, n5217, n5219, n5220_1, n5222, n5223, n5225_1, n5226, n5227, n5228, n5229, n5230_1, n5231, n5233, n5234, n5235_1, n5236, n5237, n5238, n5239, n5241, n5251, n5252, n5253, n5263, n5264, n5296, n5297, n5298_1, n5303, n5304, n5305, n5306, n5307_1, n5312, n5313, n5314, n5315, n5316_1, n5317, n5318, n5323, n5324, n5325_1, n5326, n5327, n5328, n5329_1, n5348, n5350, n5352_1, n5382, n5383_1, n5384, n5385, n5386, n5387, n5391, n5392_1, n5393, n5397, n5398, n5399, n5400, n5401_1, n5403, n5405_1, n5407, n5415, n5416, n5417, n5418, n5422, n5423, n5424_1, n5425, n5426, n5427, n5428, n5429_1, n5430, n5431, n5432, n5433_1, n5434, n5435, n5436, n5437_1, n5438, n5439, n5440, n5441, n5442_1, n5443, n5444, n5445, n5446_1, n5447, n5448, n5449, n5450, n5451_1, n5452, n5453, n5454, n5455_1, n5456, n5457, n5458, n5459, n5460_1, n5461, n5462, n5463, n5464_1, n5465, n5466, n5467, n5468, n5469_1, n5470, n5471, n5472, n5473_1, n5474, n5475, n5476, n5477, n5478_1, n5479, n5480, n5481, n5482_1, n5483, n5484, n5485, n5486, n5487_1, n5488, n5489, n5490, n5491_1, n5492, n5493, n5494, n5495, n5496_1, n5497, n5498, n5499, n5500_1, n5501, n5502, n5503, n5504_1, n5505, n5506, n5507, n5508, n5509_1, n5510, n5511, n5512, n5513, n5514_1, n5515, n5516, n5517, n5518, n5519_1, n5520, n5521, n5522, n5523, n5524_1, n5525, n5526, n5527, n5528, n5529_1, n5530, n5531, n5532, n5533, n5534_1, n5535, n5536, n5537, n5538, n5539_1, n5540, n5541, n5542, n5543, n5544_1, n5545, n5546, n5547, n5548, n5549_1, n5550, n5551, n5552, n5553, n5554_1, n5555, n5556, n5557, n5558, n5559_1, n5560, n5561, n5562, n5563, n5564_1, n5565, n5566, n5567, n5568, n5569_1, n5570, n5571, n5572, n5573, n5574_1, n5575, n5576, n5577, n5578, n5579_1, n5580, n5581, n5582, n5583, n5584_1, n5585, n5586, n5587, n5588_1, n5589, n5590, n5591, n5592_1, n5593, n5594, n5595, n5596, n5597_1, n5601_1, n5602, n5603, n5604, n5605, n5606_1, n5607, n5611_1, n5612, n5613, n5614, n5615_1, n5619, n5620_1, n5621, n5622, n5623, n5627, n5628, n5629_1, n5630, n5631, n5632, n5636, n5637, n5638, n5639_1, n5640, n5644_1, n5645, n5646, n5647, n5648, n5649_1, n5653, n5654_1, n5655, n5656, n5657, n5661, n5662, n5663, n5664_1, n5665, n5666, n5670, n5671, n5672, n5673, n5674_1, n5678, n5679_1, n5680, n5682, n5683, n5684_1, n5686, n5687, n5688, n5690, n5691, n5693, n5694_1, n5696, n5697, n5698, n5699_1, n5701, n5702, n5703, n5705, n5706, n5707, n5708, n5710, n5711, n5712, n5714_1, n5715, n5716, n5718, n5719_1, n5720, n5721, n5722, n5723, n5724_1, n5725, n5726, n5727, n5728, n5731, n5732, n5733, n5734_1, n5735, n5736, n5737, n5738, n5739_1, n5741, n5743, n5745, n5747, n5748, n5749_1, n5753, n5754_1, n5756, n5757, n5761, n5762, n5763, n5764_1, n5768, n5769_1, n5770, n5771, n5772, n5773, n5774_1, n5775, n5776, n5777, n5778, n5779_1, n5781, n5782, n5783, n5784_1, n5785, n5786, n5787, n5788, n5789_1, n5790, n5794_1, n5795, n5796, n5797, n5798, n5799_1, n5800, n5801, n5805, n5806, n5807, n5808, n5809_1, n5811, n5813, n5815, n5816, n5817, n5818_1, n5819, n5820, n5821, n5822, n5823_1, n5827, n5828_1, n5829, n5830, n5831, n5832, n5833_1, n5834, n5835, n5836, n5837, n5838_1, n5839, n5840, n5844, n5845, n5846, n5847, n5848_1, n5849, n5850, n5852, n5854, n5856, n5857, n5858_1, n5859, n5860, n5864, n5865, n5866, n5867, n5868_1, n5869, n5870, n5871, n5872, n5873_1, n5874, n5875, n5876, n5877_1, n5878, n5879, n5880, n5881_1, n5882, n5883, n5884, n5885, n5886_1, n5887, n5888, n5889, n5890, n5891_1, n5892, n5893, n5894, n5899, n5900, n5901_1, n5902, n5903, n5904, n5905, n5906_1, n5910, n5911_1, n5912, n5913, n5914, n5916_1, n5918, n5920, n5921_1, n5923, n5925, n5927, n5928, n5929, n5930, n5932, n5933, n5934, n5936_1, n5937, n5938, n5940, n5941_1, n5942, n5944, n5945, n5946_1, n5948, n5949, n5950, n5953, n5954, n5955, n5956_1, n5957, n5958, n5959, n5960, n5961_1, n5962, n5963, n5964, n5965, n5966_1, n5967, n5968, n5970, n5971_1, n5972, n5973, n5974, n5975, n5976_1, n5977, n5978, n5979, n5980, n5981_1, n5982, n5984, n5985, n5988, n5989, n6006_1, n6007, n6009, n6010, n6011_1, n6013, n6014, n6016_1, n6017, n6019, n6020, n6021_1, n6022, n6023, n6024, n6025, n6026_1, n6027, n6028, n6031_1, n6032, n6033, n6034, n6035, n6036_1, n6037, n6038, n6039, n6040, n6041_1, n6042, n6043, n6044, n6045, n6046_1, n6047, n6048, n6049, n6050, n6051_1, n6052, n6053, n6055, n6057, n6059, n6061_1, n6062, n6063, n6067, n6068, n6070, n6071_1, n6075, n6076_1, n6077, n6078, n6082, n6083, n6084, n6085, n6086_1, n6087, n6088, n6092, n6093, n6094, n6095, n6096_1, n6097, n6098, n6102, n6103, n6104, n6105, n6106_1, n6107, n6108, n6109, n6110, n6111_1, n6112, n6113, n6115, n6116_1, n6117, n6118, n6119, n6120, n6121_1, n6122, n6123, n6124, n6125, n6126_1, n6127, n6128, n6129, n6130, n6131_1, n6132, n6133, n6134, n6135, n6136_1, n6137, n6138, n6139, n6140, n6141_1, n6142, n6143, n6144, n6145, n6146_1, n6147, n6148, n6149, n6150, n6151_1, n6152, n6153, n6154, n6155, n6156_1, n6157, n6158, n6159, n6160_1, n6161, n6162, n6163, n6164_1, n6165, n6169_1, n6170, n6171, n6172, n6176, n6177, n6181, n6182, n6183, n6184_1, n6186, n6187, n6188, n6190, n6191, n6192, n6194_1, n6195, n6196, n6198, n6199_1, n6213, n6214_1, n6215, n6216, n6217, n6218, n6220, n6221, n6222, n6224_1, n6225, n6226, n6228, n6229_1, n6230, n6232, n6233, n6235, n6236, n6237, n6238, n6240, n6241, n6242, n6244_1, n6245, n6246, n6248, n6249_1, n6250, n6252, n6253, n6255, n6257, n6259_1, n6285, n6289_1, n6292, n6297, n6298, n6299_1, n6300, n6301, n6302, n6303, n6304_1, n6305, n6306, n6307, n6308, n6309_1, n6310, n6311, n6312, n6313, n6314_1, n6315, n6316, n6317, n6318, n6319_1, n6320, n6321, n6322, n6323, n6324_1, n6325, n6326, n6327, n6328, n6329_1, n6330, n6331, n6332, n6333, n6334_1, n6335, n6336, n6337, n6338, n6339_1, n6340, n6341, n6342, n6343, n6344_1, n6345, n6346, n6347, n6348, n6349_1, n6350, n6351, n6352, n6356, n6357, n6358, n6359_1, n6360, n6362, n6364_1, n6367, n6369_1, n6371, n6401, n6402, n6403, n6404_1, n6405, n6406, n6410, n6411, n6412, n6416, n6417, n6419_1, n6421, n6429_1, n6430, n6431, n6432, n6436, n6437, n6438, n6439_1, n6440, n6441, n6442, n6443, n6444_1, n6445, n6446, n6447, n6448, n6449_1, n6450, n6451, n6452, n6453, n6454_1, n6455, n6456, n6457, n6458, n6459_1, n6460, n6461, n6462, n6463, n6464_1, n6465, n6466, n6467, n6468, n6469_1, n6470, n6471, n6472, n6473, n6474_1, n6475, n6476, n6477, n6478, n6479_1, n6480, n6481, n6482, n6483, n6484_1, n6485, n6486, n6487, n6488, n6489_1, n6490, n6491, n6492, n6493, n6494_1, n6495, n6496, n6497, n6498, n6499_1, n6500, n6501, n6502, n6503, n6504_1, n6505, n6506, n6507, n6508, n6509_1, n6510, n6511, n6512, n6513, n6514_1, n6515, n6516, n6517, n6518, n6519_1, n6520, n6521, n6522, n6523, n6524_1, n6525, n6526, n6527, n6528, n6529_1, n6530, n6531, n6532, n6533, n6534_1, n6535, n6536, n6537, n6538, n6539_1, n6540, n6541, n6542, n6543, n6544_1, n6545, n6546, n6547, n6548, n6549_1, n6550, n6551, n6552, n6553, n6554_1, n6555, n6556, n6557, n6558, n6559_1, n6560, n6561, n6562, n6563, n6564_1, n6565, n6566, n6567, n6568, n6569_1, n6570, n6571, n6572, n6573, n6574_1, n6575, n6576, n6577, n6578, n6579_1, n6580, n6581, n6582, n6583_1, n6584, n6585, n6586, n6587_1, n6588, n6589, n6590, n6591, n6592_1, n6593, n6594, n6595, n6596_1, n6597, n6598, n6599, n6600_1, n6601, n6602, n6603, n6604, n6605_1, n6606, n6607, n6608, n6609, n6610_1, n6611, n6615_1, n6616, n6617, n6618, n6619, n6620_1, n6621, n6625_1, n6626, n6627, n6628, n6629, n6633, n6634, n6635_1, n6636, n6637, n6641, n6642, n6643, n6644, n6645_1, n6646, n6650_1, n6651, n6652, n6653, n6654, n6658, n6659, n6660_1, n6661, n6662, n6663, n6667, n6668, n6669, n6670_1, n6671, n6675_1, n6676, n6677, n6678, n6679, n6680_1, n6684, n6685_1, n6686, n6687, n6688, n6692, n6693, n6694, n6696, n6697, n6698, n6700_1, n6701, n6702, n6704, n6705_1, n6707, n6708, n6710_1, n6711, n6712, n6713, n6715_1, n6716, n6717, n6719, n6720_1, n6721, n6722, n6724, n6725_1, n6726, n6728, n6729, n6730_1, n6732, n6733, n6734, n6735_1, n6736, n6737, n6738, n6739, n6740_1, n6741, n6744, n6745_1, n6746, n6747, n6748, n6749, n6750_1, n6751, n6752, n6754, n6756, n6758, n6760_1, n6761, n6762, n6766, n6767, n6769, n6770_1, n6774, n6775_1, n6776, n6777, n6781, n6782, n6783, n6784, n6785_1, n6786, n6787, n6788, n6789, n6790_1, n6791, n6792, n6794, n6795_1, n6796, n6797, n6798, n6799, n6800_1, n6801, n6802, n6803, n6807, n6808, n6809, n6810_1, n6811, n6812, n6813, n6814, n6818, n6819, n6820_1, n6821, n6822, n6824, n6826, n6828, n6829, n6830_1, n6831, n6832, n6833, n6834, n6835_1, n6836, n6840, n6841, n6842, n6843, n6844_1, n6845, n6846, n6847, n6848_1, n6849, n6850, n6851, n6852, n6853_1, n6857_1, n6858, n6859, n6860, n6861, n6862_1, n6863, n6865, n6867, n6869, n6870, n6871_1, n6872, n6873, n6877, n6878, n6879, n6880_1, n6881, n6882, n6883, n6884_1, n6885, n6886, n6887, n6888, n6889_1, n6890, n6891, n6892, n6893_1, n6894, n6895, n6896, n6897, n6898_1, n6899, n6900, n6901, n6902_1, n6903, n6904, n6905, n6906, n6907_1, n6912, n6913, n6914, n6915, n6916_1, n6917, n6918, n6919, n6923, n6924, n6925, n6926_1, n6927, n6929, n6931_1, n6933, n6934, n6936_1, n6938, n6940, n6941_1, n6942, n6944, n6945, n6946_1, n6948, n6949, n6950, n6952, n6953, n6954, n6956_1, n6957, n6958, n6960, n6961_1, n6962, n6965, n6966_1, n6967, n6968, n6969, n6970, n6971_1, n6972, n6973, n6974, n6975, n6976_1, n6977, n6978, n6979, n6980, n6983, n6984, n6987, n6988, n7005, n7006, n7008_1, n7009, n7010, n7011, n7013, n7014, n7016, n7017_1, n7019, n7020, n7021_1, n7022, n7023, n7024, n7025, n7026_1, n7027, n7028, n7031, n7032, n7033, n7034, n7035_1, n7036, n7037, n7038, n7039_1, n7040, n7041, n7042, n7043, n7044_1, n7045, n7046, n7047, n7048_1, n7049, n7050, n7051, n7053_1, n7055, n7057_1, n7059, n7060, n7061, n7065, n7066_1, n7068, n7069, n7073, n7074, n7075_1, n7076, n7080_1, n7081, n7082, n7083, n7084_1, n7085, n7086, n7090, n7091, n7092, n7093_1, n7094, n7095, n7096, n7100, n7101, n7102_1, n7103, n7104, n7105, n7106_1, n7107, n7108, n7109, n7110_1, n7111, n7113, n7114, n7115_1, n7116, n7117, n7118, n7119, n7120_1, n7121, n7122, n7123, n7124, n7125_1, n7126, n7127, n7128, n7129, n7130_1, n7131, n7132, n7133, n7134_1, n7135, n7136, n7137, n7138_1, n7139, n7140, n7141, n7142, n7143_1, n7144, n7145, n7146, n7147_1, n7148, n7149, n7150, n7151, n7152_1, n7153, n7154, n7155, n7156_1, n7157, n7158, n7159, n7160, n7161_1, n7162, n7163, n7167, n7168, n7169, n7170_1, n7174_1, n7175, n7179_1, n7180, n7181, n7182, n7184, n7185, n7186, n7188_1, n7189, n7190, n7192_1, n7193, n7194, n7196, n7197_1, n7198, n7212, n7213, n7214, n7215_1, n7216, n7217, n7219, n7220_1, n7221, n7223, n7224, n7225_1, n7227, n7228, n7229, n7231, n7232, n7234, n7235_1, n7236, n7237, n7239, n7240_1, n7241, n7243, n7244, n7245_1, n7247, n7248, n7249, n7251, n7252, n7254, n7256, n7258, n7284, n7288, n7291, n7296, n7297, n7298_1, n7299, n7300, n7301, n7302_1, n7303, n7304, n7305, n7306, n7307_1, n7308, n7309, n7310, n7311, n7312_1, n7313, n7314, n7315, n7316_1, n7317, n7318, n7319, n7320, n7321_1, n7322, n7323, n7324, n7325_1, n7326, n7327, n7328, n7329, n7330_1, n7331, n7332, n7333, n7334, n7335_1, n7336, n7337, n7338, n7339, n7340_1, n7341, n7342, n7343, n7344, n7345_1, n7346, n7347, n7348, n7349, n7350_1, n7351, n7355_1, n7356, n7357, n7358, n7359, n7361, n7363, n7366, n7368, n7370_1, n7400_1, n7401, n7402, n7403, n7404, n7405_1, n7409, n7410_1, n7411, n7415_1, n7416, n7418, n7420_1, n7428, n7429, n7430_1, n7431, n7435_1, n7436, n7437, n7438, n7439, n7440_1, n7441, n7442, n7443, n7444, n7445_1, n7446, n7447, n7448, n7449, n7450_1, n7451, n7452, n7453, n7454, n7455_1, n7456, n7457, n7458, n7459, n7460_1, n7461, n7462, n7463, n7464, n7465_1, n7466, n7467, n7468, n7469, n7470_1, n7471, n7472, n7473, n7474, n7475_1, n7476, n7477, n7478, n7479, n7480_1, n7481, n7482, n7483, n7484, n7485_1, n7486, n7487, n7488, n7489, n7490_1, n7491, n7492, n7493, n7494, n7495_1, n7496, n7497, n7498, n7499, n7500_1, n7501, n7502, n7503, n7504, n7505_1, n7506, n7507, n7508, n7509, n7510_1, n7511, n7512, n7513, n7514, n7515_1, n7516, n7517, n7518, n7519_1, n7520, n7521, n7522, n7523, n7524_1, n7525, n7526, n7527, n7528, n7529_1, n7530, n7531, n7532, n7533, n7534_1, n7535, n7536, n7537, n7538, n7539_1, n7540, n7541, n7542, n7543, n7544_1, n7545, n7546, n7547, n7548, n7549_1, n7550, n7551, n7552, n7553, n7554_1, n7555, n7556, n7557, n7558, n7559_1, n7560, n7561, n7562, n7563, n7564_1, n7565, n7566, n7567, n7568, n7569_1, n7570, n7571, n7572, n7573, n7574_1, n7575, n7576, n7577, n7578_1, n7579, n7580, n7581, n7582_1, n7583, n7584, n7585, n7586, n7587_1, n7588, n7589, n7590, n7591, n7592_1, n7593, n7594, n7595, n7596, n7597_1, n7598, n7599, n7600, n7601, n7602_1, n7603, n7604, n7605, n7606, n7607_1, n7608, n7609, n7610, n7614, n7615, n7616, n7617_1, n7618, n7619, n7620, n7624, n7625, n7626, n7627_1, n7628, n7632_1, n7633, n7634, n7635, n7636, n7640, n7641, n7642_1, n7643, n7644, n7645, n7649, n7650, n7651, n7652_1, n7653, n7657_1, n7658, n7659, n7660, n7661, n7662_1, n7666, n7667_1, n7668, n7669, n7670, n7674, n7675, n7676, n7677_1, n7678, n7679, n7683, n7684, n7685, n7686, n7687_1, n7691, n7692_1, n7693, n7695, n7696, n7697_1, n7699, n7700, n7701, n7703, n7704, n7706, n7707_1, n7709, n7710, n7711, n7712_1, n7714, n7715, n7716, n7718, n7719, n7720, n7721, n7723, n7724, n7725, n7727_1, n7728, n7729, n7731, n7732_1, n7733, n7734, n7735, n7736, n7737_1, n7738, n7739, n7740, n7743, n7744, n7745, n7746, n7747_1, n7748, n7749, n7750, n7751, n7753, n7755, n7757_1, n7759, n7760, n7761, n7765, n7766, n7768, n7769, n7773, n7774, n7775, n7776, n7780, n7781, n7782_1, n7783, n7784, n7785, n7786, n7787_1, n7788, n7789, n7790, n7791, n7793, n7794, n7795, n7796, n7797_1, n7798, n7799, n7800, n7801, n7802_1, n7806, n7807_1, n7808, n7809, n7810, n7811, n7812_1, n7813, n7817_1, n7818, n7819, n7820, n7821, n7823, n7825, n7827_1, n7828, n7829, n7830, n7831, n7832_1, n7833, n7834, n7835, n7839, n7840, n7841, n7842_1, n7843, n7844, n7845, n7846, n7847_1, n7848, n7849, n7850, n7851, n7852_1, n7856, n7857_1, n7858, n7859, n7860, n7861, n7862_1, n7864, n7866, n7868, n7869, n7870, n7871, n7872_1, n7876, n7877_1, n7878, n7879, n7880, n7881, n7882_1, n7883, n7884, n7885, n7886, n7887_1, n7888, n7889, n7890, n7891, n7892_1, n7893, n7894, n7895, n7896, n7897_1, n7898, n7899, n7900, n7901, n7902_1, n7903, n7904, n7905, n7906, n7911, n7912_1, n7913, n7914, n7915, n7916, n7917_1, n7918, n7922_1, n7923, n7924, n7925, n7926, n7928, n7930, n7932_1, n7933, n7935, n7937_1, n7939, n7940, n7941, n7943, n7944, n7945, n7947_1, n7948, n7949, n7951, n7952_1, n7953, n7955, n7956, n7957_1, n7959, n7960, n7961, n7964, n7965, n7966, n7967_1, n7968, n7969, n7970, n7971, n7972_1, n7973, n7974, n7975, n7976, n7977_1, n7978, n7979, n7982_1, n7983, n7986, n7987_1, n8004, n8005, n8007_1, n8008, n8009, n8011, n8012_1, n8014, n8015, n8017_1, n8018, n8019, n8020, n8021, n8022_1, n8023, n8024, n8025, n8026, n8029, n8030, n8031, n8032_1, n8033, n8034, n8035, n8036, n8037_1, n8038, n8039, n8040, n8041, n8042_1, n8043, n8044, n8045, n8046, n8047_1, n8048, n8049, n8051, n8053, n8055, n8057_1, n8058, n8059, n8063, n8064, n8066, n8067_1, n8071, n8072_1, n8073, n8074, n8078, n8079, n8080, n8081, n8082_1, n8083, n8084, n8088, n8089, n8090, n8091, n8092_1, n8093, n8094, n8098, n8099, n8100, n8101, n8102_1, n8103, n8104, n8105, n8106, n8107_1, n8108, n8109, n8111_1, n8112, n8113, n8114, n8115, n8116_1, n8117, n8118, n8119, n8120, n8121_1, n8122, n8123, n8124, n8125, n8126_1, n8127, n8128, n8129, n8130, n8131_1, n8132, n8133, n8134, n8135, n8136_1, n8137, n8138, n8139, n8140, n8141_1, n8142, n8143, n8144, n8145, n8146_1, n8147, n8148, n8149, n8150, n8151_1, n8152, n8153, n8154, n8155, n8156_1, n8157, n8158, n8159, n8160, n8161_1, n8165, n8166_1, n8167, n8168, n8172, n8173, n8177, n8178, n8179, n8180, n8182, n8183, n8184, n8186_1, n8187, n8188, n8190, n8191_1, n8192, n8194, n8195, n8196_1, n8210, n8211_1, n8212, n8213, n8214, n8215, n8217, n8218, n8219, n8221_1, n8222, n8223, n8225, n8226_1, n8227, n8229, n8230, n8232, n8233, n8234, n8235, n8237, n8238, n8239, n8241, n8242, n8243, n8245, n8246, n8247, n8249, n8250, n8252, n8254, n8256, n8282, n8286, n8289, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8351, n8352, n8353, n8354, n8355, n8357, n8359, n8362, n8364, n8366, n8396, n8397, n8398, n8399, n8400, n8401, n8405, n8406, n8407, n8411, n8412, n8414, n8416, n8424, n8425, n8426, n8427, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8620, n8621, n8622, n8623, n8624, n8628, n8629, n8630, n8631, n8632, n8636, n8637, n8638, n8639, n8640, n8641, n8645, n8646, n8647, n8648, n8649, n8653, n8654, n8655, n8656, n8657, n8658, n8662, n8663, n8664, n8665, n8666, n8670, n8671, n8672, n8673, n8674, n8675, n8679, n8680, n8681, n8682, n8683, n8687, n8688, n8689, n8691, n8692, n8693, n8695, n8696, n8697, n8699, n8700, n8702, n8703, n8705, n8706, n8707, n8708, n8710, n8711, n8712, n8714, n8715, n8716, n8717, n8719, n8720, n8721, n8723, n8724, n8725, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8749, n8751, n8753, n8755, n8756, n8757, n8761, n8762, n8764, n8765, n8769, n8770, n8771, n8772, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8813, n8814, n8815, n8816, n8817, n8819, n8821, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8860, n8862, n8864, n8865, n8866, n8867, n8868, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8918, n8919, n8920, n8921, n8922, n8924, n8926, n8928, n8929, n8931, n8933, n8935, n8936, n8937, n8939, n8940, n8941, n8943, n8944, n8945, n8947, n8948, n8949, n8951, n8952, n8953, n8955, n8956, n8957, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8978, n8979, n8982, n8983, n9000, n9001, n9003, n9004, n9005, n9007, n9008, n9010, n9011, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9047, n9049, n9051, n9053, n9054, n9055, n9059, n9060, n9062, n9063, n9067, n9068, n9069, n9070, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9161, n9162, n9163, n9164, n9168, n9169, n9173, n9174, n9175, n9177, n9178, n9179, n9181, n9182, n9183, n9185, n9186, n9187, n9189, n9190, n9191, n9205, n9206, n9207, n9208, n9209, n9210, n9212, n9213, n9214, n9216, n9217, n9218, n9220, n9221, n9222, n9224, n9225, n9227, n9228, n9229, n9230, n9232, n9233, n9234, n9236, n9237, n9238, n9240, n9241, n9242, n9244, n9245, n9247, n9249, n9251, n9277, n9281, n9284, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9348, n9349, n9350, n9351, n9352, n9354, n9356, n9358, n9360, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9385, n9386, n9387, n9388, n9389, n9390, n9392, n9393, n9395, n9396, n9397, n9398, n9399, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9409, n9410, n9411, n9412, n9413, n9414, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9424, n9425, n9426, n9427, n9428, n9429, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9496, n9497, n9498, n9500, n9501, n9502, n9503, n9505, n9506, n9507, n9508, n9509, n9511, n9512, n9513, n9514, n9515, n9516, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9526, n9527, n9528, n9529, n9530, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9599, n9600, n9601, n9602, n9603, n9604, n9606, n9607, n9608, n9609, n9610, n9612, n9613, n9614, n9615, n9616, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9626, n9627, n9628, n9629, n9630, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9708, n9710, n9711, n9712, n9713, n9714, n9716, n9717, n9718, n9719, n9720, n9721, n9723, n9724, n9725, n9726, n9727, n9728, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9738, n9739, n9740, n9741, n9742, n9743, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9779, n9780, n9781, n9783, n9784, n9786, n9787, n9789, n9790, n9792, n9793, n9795, n9796, n9797, n9799, n9800, n9802, n9803, n9804, n9805, n9807, n9808, n9810, n9811, n9813, n9814, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9844, n9845, n9846, n9847, n9848, n9849, n9850;
INVX1    g0000(.A(g3040), .Y(n5042));
OAI21X1  g0001(.A0(g2986), .A1(n5042), .B0(g2987), .Y(g16496));
INVX1    g0002(.A(g3233), .Y(n5044_1));
NOR2X1   g0003(.A(n5044_1), .B(g3230), .Y(n5045));
INVX1    g0004(.A(g3201), .Y(n5046));
INVX1    g0005(.A(g3207), .Y(n5047));
NOR4X1   g0006(.A(n5047), .B(g3204), .C(n5046), .D(g3188), .Y(n5048));
NOR4X1   g0007(.A(g3197), .B(g3194), .C(g3191), .D(g3198), .Y(n5049_1));
AND2X1   g0008(.A(n5049_1), .B(n5048), .Y(n5050));
INVX1    g0009(.A(n5050), .Y(n5051));
OAI21X1  g0010(.A0(n5051), .A1(g3123), .B0(n5045), .Y(g24734));
INVX1    g0011(.A(g3204), .Y(n5053));
NOR4X1   g0012(.A(g3207), .B(n5053), .C(g3201), .D(g3188), .Y(n5054_1));
AND2X1   g0013(.A(n5054_1), .B(n5049_1), .Y(n5055));
AOI22X1  g0014(.A0(n5050), .A1(g3126), .B0(g3112), .B1(n5055), .Y(n5056));
NAND2X1  g0015(.A(n5056), .B(n5045), .Y(g25420));
INVX1    g0016(.A(g3125), .Y(n5058));
AOI22X1  g0017(.A0(n5050), .A1(n5058), .B0(g3110), .B1(n5055), .Y(n5059_1));
AND2X1   g0018(.A(n5059_1), .B(n5045), .Y(n968));
INVX1    g0019(.A(n968), .Y(g25435));
AOI22X1  g0020(.A0(n5050), .A1(g3124), .B0(g3111), .B1(n5055), .Y(n5062));
NAND2X1  g0021(.A(n5062), .B(n5045), .Y(g25442));
INVX1    g0022(.A(g3151), .Y(n5064_1));
INVX1    g0023(.A(g3142), .Y(n5065));
INVX1    g0024(.A(g3147), .Y(n5066));
NAND3X1  g0025(.A(n5066), .B(n5065), .C(n5064_1), .Y(n5067));
NOR2X1   g0026(.A(g2985), .B(g2984), .Y(n5068));
AOI21X1  g0027(.A0(n5068), .A1(g3151), .B0(g3142), .Y(n5069_1));
NOR2X1   g0028(.A(g2991), .B(g2992), .Y(n5070));
NOR3X1   g0029(.A(n5070), .B(n5065), .C(g3151), .Y(n5071));
NOR3X1   g0030(.A(n5071), .B(n5069_1), .C(g3147), .Y(n5072));
NAND3X1  g0031(.A(g3142), .B(g3151), .C(g3097), .Y(n5073));
AND2X1   g0032(.A(n5073), .B(g3147), .Y(n5074_1));
OAI21X1  g0033(.A0(n5074_1), .A1(n5072), .B0(n5067), .Y(g25489));
INVX1    g0034(.A(n5045), .Y(n5076));
INVX1    g0035(.A(g3092), .Y(n5077));
INVX1    g0036(.A(g3197), .Y(n5078));
NOR4X1   g0037(.A(n5078), .B(g3194), .C(g3191), .D(g3198), .Y(n5079_1));
AND2X1   g0038(.A(g3188), .B(g3207), .Y(n5080));
NAND4X1  g0039(.A(n5079_1), .B(g3204), .C(n5046), .D(n5080), .Y(n5081));
NOR3X1   g0040(.A(g3188), .B(n5047), .C(n5053), .Y(n5082));
NAND3X1  g0041(.A(n5082), .B(n5049_1), .C(g3201), .Y(n5083));
OAI22X1  g0042(.A0(n5081), .A1(n5077), .B0(n5065), .B1(n5083), .Y(n5084_1));
AND2X1   g0043(.A(n5079_1), .B(n5046), .Y(n5085));
INVX1    g0044(.A(n5085), .Y(n5086));
NOR4X1   g0045(.A(g3188), .B(n5047), .C(g3204), .D(n5086), .Y(n5087));
NAND2X1  g0046(.A(n5087), .B(g3084), .Y(n5088));
NOR4X1   g0047(.A(g3207), .B(g3204), .C(g3201), .D(g3188), .Y(n5089_1));
NAND3X1  g0048(.A(n5089_1), .B(n5079_1), .C(g3210), .Y(n5090));
AND2X1   g0049(.A(n5080), .B(n5053), .Y(n5091));
AND2X1   g0050(.A(n5091), .B(n5085), .Y(n5092));
INVX1    g0051(.A(g3188), .Y(n5093));
NOR4X1   g0052(.A(n5093), .B(g3207), .C(g3204), .D(n5086), .Y(n5094_1));
AOI22X1  g0053(.A0(n5092), .A1(g3085), .B0(g3211), .B1(n5094_1), .Y(n5095));
NAND3X1  g0054(.A(n5095), .B(n5090), .C(n5088), .Y(n5096));
NAND4X1  g0055(.A(n5079_1), .B(n5046), .C(g3091), .D(n5082), .Y(n5097));
AND2X1   g0056(.A(n5079_1), .B(n5054_1), .Y(n5098));
INVX1    g0057(.A(n5079_1), .Y(n5099_1));
NAND3X1  g0058(.A(g3188), .B(n5047), .C(g3204), .Y(n5100));
NOR3X1   g0059(.A(n5100), .B(n5099_1), .C(g3201), .Y(n5101));
AOI22X1  g0060(.A0(n5098), .A1(g3086), .B0(g3087), .B1(n5101), .Y(n5102));
NOR4X1   g0061(.A(g3207), .B(g3204), .C(n5046), .D(n5093), .Y(n5103));
NAND3X1  g0062(.A(n5103), .B(n5079_1), .C(g3094), .Y(n5104_1));
NOR4X1   g0063(.A(g3207), .B(n5053), .C(n5046), .D(g3188), .Y(n5105));
NAND3X1  g0064(.A(n5105), .B(n5049_1), .C(g3136), .Y(n5106));
NAND3X1  g0065(.A(n5079_1), .B(n5048), .C(g3095), .Y(n5107));
NAND4X1  g0066(.A(n5079_1), .B(g3201), .C(g3096), .D(n5091), .Y(n5108));
NAND4X1  g0067(.A(n5107), .B(n5106), .C(n5104_1), .D(n5108), .Y(n5109_1));
NAND2X1  g0068(.A(n5089_1), .B(n5049_1), .Y(n5110));
NAND3X1  g0069(.A(n5054_1), .B(n5049_1), .C(g3120), .Y(n5111));
OAI21X1  g0070(.A0(n5110), .A1(n5068), .B0(n5111), .Y(n5112));
NOR4X1   g0071(.A(g3207), .B(g3204), .C(n5046), .D(g3188), .Y(n5113));
NAND3X1  g0072(.A(n5113), .B(n5079_1), .C(g3093), .Y(n5114_1));
NAND3X1  g0073(.A(n5049_1), .B(n5048), .C(g3132), .Y(n5115));
NAND2X1  g0074(.A(n5115), .B(n5114_1), .Y(n5116));
NOR3X1   g0075(.A(n5116), .B(n5112), .C(n5109_1), .Y(n5117));
NAND3X1  g0076(.A(n5117), .B(n5102), .C(n5097), .Y(n5118));
OR4X1    g0077(.A(n5096), .B(n5084_1), .C(n5076), .D(n5118), .Y(g26104));
INVX1    g0078(.A(g3104), .Y(n5120));
OAI22X1  g0079(.A0(n5081), .A1(n5120), .B0(n5066), .B1(n5083), .Y(n5121));
INVX1    g0080(.A(n5121), .Y(n5122));
AND2X1   g0081(.A(n5089_1), .B(n5079_1), .Y(n5123));
AOI22X1  g0082(.A0(n5087), .A1(g3099), .B0(g3097), .B1(n5123), .Y(n5124_1));
AOI22X1  g0083(.A0(n5092), .A1(g3100), .B0(g3098), .B1(n5094_1), .Y(n5125));
NAND3X1  g0084(.A(n5125), .B(n5124_1), .C(n5122), .Y(n5126));
NAND4X1  g0085(.A(n5079_1), .B(n5046), .C(g3103), .D(n5082), .Y(n5127));
AOI22X1  g0086(.A0(n5098), .A1(g3101), .B0(g3102), .B1(n5101), .Y(n5128));
AND2X1   g0087(.A(n5128), .B(n5127), .Y(n5129_1));
INVX1    g0088(.A(n5129_1), .Y(n5130));
NAND3X1  g0089(.A(n5103), .B(n5079_1), .C(g3106), .Y(n5131));
NAND3X1  g0090(.A(n5105), .B(n5049_1), .C(g3134), .Y(n5132));
NAND3X1  g0091(.A(n5079_1), .B(n5048), .C(g3107), .Y(n5133));
NAND4X1  g0092(.A(n5079_1), .B(g3201), .C(g3108), .D(n5091), .Y(n5134_1));
NAND4X1  g0093(.A(n5133), .B(n5132), .C(n5131), .D(n5134_1), .Y(n5135));
NAND3X1  g0094(.A(n5054_1), .B(n5049_1), .C(g3114), .Y(n5136));
OAI21X1  g0095(.A0(n5110), .A1(n5070), .B0(n5136), .Y(n5137));
NAND3X1  g0096(.A(n5113), .B(n5079_1), .C(g3105), .Y(n5138_1));
OAI21X1  g0097(.A0(n5051), .A1(g3128), .B0(n5138_1), .Y(n5139));
NOR3X1   g0098(.A(n5139), .B(n5137), .C(n5135), .Y(n5140));
INVX1    g0099(.A(n5140), .Y(n5141));
NOR4X1   g0100(.A(n5130), .B(n5126), .C(n5076), .D(n5141), .Y(n953));
INVX1    g0101(.A(n953), .Y(g26135));
AOI22X1  g0102(.A0(n5087), .A1(g3161), .B0(g3167), .B1(n5098), .Y(n5144));
NAND3X1  g0103(.A(n5049_1), .B(n5048), .C(g3127), .Y(n5145));
NAND3X1  g0104(.A(n5089_1), .B(n5079_1), .C(g3155), .Y(n5146));
NAND3X1  g0105(.A(n5146), .B(n5145), .C(n5144), .Y(n5147_1));
INVX1    g0106(.A(g3176), .Y(n5148));
NAND3X1  g0107(.A(n5105), .B(n5049_1), .C(g3135), .Y(n5149));
OAI21X1  g0108(.A0(n5081), .A1(n5148), .B0(n5149), .Y(n5150));
AND2X1   g0109(.A(n5092), .B(g3164), .Y(n5151));
AND2X1   g0110(.A(n5094_1), .B(g3158), .Y(n5152_1));
NOR4X1   g0111(.A(n5151), .B(n5150), .C(n5147_1), .D(n5152_1), .Y(n5153));
AND2X1   g0112(.A(n5055), .B(g3113), .Y(n5154));
AND2X1   g0113(.A(n5101), .B(g3170), .Y(n5155));
AND2X1   g0114(.A(n5085), .B(n5082), .Y(n5156_1));
AND2X1   g0115(.A(n5156_1), .B(g3173), .Y(n5157));
NAND3X1  g0116(.A(n5113), .B(n5079_1), .C(g3179), .Y(n5158));
NAND3X1  g0117(.A(n5103), .B(n5079_1), .C(g3182), .Y(n5159));
NAND4X1  g0118(.A(n5079_1), .B(g3201), .C(g3088), .D(n5091), .Y(n5160));
NAND3X1  g0119(.A(n5079_1), .B(n5048), .C(g3185), .Y(n5161_1));
NAND4X1  g0120(.A(n5160), .B(n5159), .C(n5158), .D(n5161_1), .Y(n5162));
NOR4X1   g0121(.A(n5157), .B(n5155), .C(n5154), .D(n5162), .Y(n5163));
NAND3X1  g0122(.A(n5163), .B(n5153), .C(n5045), .Y(g26149));
OAI21X1  g0123(.A0(n5113), .A1(n5089_1), .B0(n5049_1), .Y(n5165_1));
NAND2X1  g0124(.A(n5103), .B(n5049_1), .Y(n5166));
OR4X1    g0125(.A(n5099_1), .B(g185), .C(n5046), .D(n5100), .Y(n5167));
NAND3X1  g0126(.A(n5167), .B(n5166), .C(n5165_1), .Y(n5168));
OAI21X1  g0127(.A0(g2991), .A1(g2992), .B0(g3114), .Y(n5169));
OAI21X1  g0128(.A0(g2985), .A1(g2984), .B0(g3120), .Y(n5170_1));
NAND4X1  g0129(.A(n5169), .B(n5105), .C(n5079_1), .D(n5170_1), .Y(n5171));
NAND3X1  g0130(.A(n5105), .B(n5049_1), .C(g3139), .Y(n5172));
NAND2X1  g0131(.A(n5172), .B(n5171), .Y(n5173));
OAI22X1  g0132(.A0(n5051), .A1(g3133), .B0(n5064_1), .B1(n5083), .Y(n5174_1));
NOR4X1   g0133(.A(n5173), .B(n5168), .C(n5076), .D(n5174_1), .Y(n943));
INVX1    g0134(.A(n943), .Y(g27380));
INVX1    g0135(.A(g2950), .Y(n5177));
NOR2X1   g0136(.A(n5177), .B(g51), .Y(n274));
INVX1    g0137(.A(g2817), .Y(n5179_1));
NOR2X1   g0138(.A(n5179_1), .B(g51), .Y(n279));
OR2X1    g0139(.A(g2933), .B(g51), .Y(n284));
NOR2X1   g0140(.A(g2883), .B(n5177), .Y(n5182));
INVX1    g0141(.A(g2900), .Y(n5183_1));
NAND4X1  g0142(.A(n5183_1), .B(g2892), .C(g2888), .D(g2908), .Y(n5184));
INVX1    g0143(.A(g2903), .Y(n5185));
OR4X1    g0144(.A(g2896), .B(g2883), .C(n5177), .D(n5185), .Y(n5186));
NOR2X1   g0145(.A(n5186), .B(n5184), .Y(n5187));
AND2X1   g0146(.A(g2883), .B(n5177), .Y(n5188_1));
OR4X1    g0147(.A(n5187), .B(n5182), .C(g2814), .D(n5188_1), .Y(n289));
NAND2X1  g0148(.A(g2883), .B(g2950), .Y(n5190));
XOR2X1   g0149(.A(n5190), .B(g2888), .Y(n5191));
NOR3X1   g0150(.A(n5191), .B(n5187), .C(g2814), .Y(n294));
NAND3X1  g0151(.A(g2888), .B(g2883), .C(g2950), .Y(n5193));
XOR2X1   g0152(.A(n5193), .B(g2896), .Y(n5194));
NOR3X1   g0153(.A(n5194), .B(n5187), .C(g2814), .Y(n299));
NAND4X1  g0154(.A(g2888), .B(g2883), .C(g2950), .D(g2896), .Y(n5196));
XOR2X1   g0155(.A(n5196), .B(g2892), .Y(n5197_1));
NOR3X1   g0156(.A(n5197_1), .B(n5187), .C(g2814), .Y(n304));
INVX1    g0157(.A(g2892), .Y(n5199));
NOR2X1   g0158(.A(n5196), .B(n5199), .Y(n5200));
XOR2X1   g0159(.A(n5200), .B(n5185), .Y(n5201_1));
NOR3X1   g0160(.A(n5201_1), .B(n5187), .C(g2814), .Y(n309));
NOR3X1   g0161(.A(n5196), .B(n5185), .C(n5199), .Y(n5203));
XOR2X1   g0162(.A(n5203), .B(n5183_1), .Y(n5204));
NOR3X1   g0163(.A(n5204), .B(n5187), .C(g2814), .Y(n314));
OR4X1    g0164(.A(n5183_1), .B(n5185), .C(n5199), .D(n5196), .Y(n5206_1));
XOR2X1   g0165(.A(n5206_1), .B(g2908), .Y(n5207));
NOR3X1   g0166(.A(n5207), .B(n5187), .C(g2814), .Y(n319));
INVX1    g0167(.A(g2912), .Y(n5209));
NOR4X1   g0168(.A(n5184), .B(g2917), .C(n5209), .D(n5186), .Y(n5210_1));
INVX1    g0169(.A(g2920), .Y(n5211));
NOR2X1   g0170(.A(n5211), .B(g2924), .Y(n5212));
AOI21X1  g0171(.A0(n5212), .A1(n5210_1), .B0(g2814), .Y(n5213));
XOR2X1   g0172(.A(n5187), .B(n5209), .Y(n5214));
NAND2X1  g0173(.A(n5214), .B(n5213), .Y(n324));
NOR3X1   g0174(.A(n5186), .B(n5184), .C(n5209), .Y(n5216));
XOR2X1   g0175(.A(n5216), .B(g2917), .Y(n5217));
AND2X1   g0176(.A(n5217), .B(n5213), .Y(n329));
AND2X1   g0177(.A(n5216), .B(g2917), .Y(n5219));
XOR2X1   g0178(.A(n5219), .B(g2924), .Y(n5220_1));
AND2X1   g0179(.A(n5220_1), .B(n5213), .Y(n334));
NAND3X1  g0180(.A(n5216), .B(g2924), .C(g2917), .Y(n5222));
XOR2X1   g0181(.A(n5222), .B(n5211), .Y(n5223));
AND2X1   g0182(.A(n5223), .B(n5213), .Y(n339));
XOR2X1   g0183(.A(g2938), .B(g2935), .Y(n5225_1));
XOR2X1   g0184(.A(g2944), .B(g2941), .Y(n5226));
XOR2X1   g0185(.A(n5226), .B(n5225_1), .Y(n5227));
XOR2X1   g0186(.A(g2953), .B(g2947), .Y(n5228));
XOR2X1   g0187(.A(g2959), .B(g2956), .Y(n5229));
XOR2X1   g0188(.A(n5229), .B(n5228), .Y(n5230_1));
XOR2X1   g0189(.A(n5230_1), .B(n5227), .Y(n5231));
XOR2X1   g0190(.A(n5231), .B(g2934), .Y(n344));
XOR2X1   g0191(.A(g2966), .B(g2963), .Y(n5233));
XOR2X1   g0192(.A(g2972), .B(g2969), .Y(n5234));
XOR2X1   g0193(.A(n5234), .B(n5233), .Y(n5235_1));
XOR2X1   g0194(.A(g2978), .B(g2975), .Y(n5236));
XOR2X1   g0195(.A(g2874), .B(g2981), .Y(n5237));
XOR2X1   g0196(.A(n5237), .B(n5236), .Y(n5238));
XOR2X1   g0197(.A(n5238), .B(n5235_1), .Y(n5239));
XOR2X1   g0198(.A(n5239), .B(g2962), .Y(n349));
INVX1    g0199(.A(g2930), .Y(n5241));
OAI21X1  g0200(.A0(g2929), .A1(n5241), .B0(g2879), .Y(n363));
MX2X1    g0201(.A(g1506), .B(g2959), .S0(g2879), .Y(n458));
MX2X1    g0202(.A(g1501), .B(g2956), .S0(g2879), .Y(n463));
MX2X1    g0203(.A(g1496), .B(g2953), .S0(g2879), .Y(n468));
MX2X1    g0204(.A(g1491), .B(g2947), .S0(g2879), .Y(n473));
MX2X1    g0205(.A(g1486), .B(g2944), .S0(g2879), .Y(n478));
MX2X1    g0206(.A(g1481), .B(g2941), .S0(g2879), .Y(n483));
MX2X1    g0207(.A(g1476), .B(g2938), .S0(g2879), .Y(n488));
MX2X1    g0208(.A(g1471), .B(g2935), .S0(g2879), .Y(n493));
INVX1    g0209(.A(g3231), .Y(n5251));
NAND2X1  g0210(.A(g3139), .B(n5251), .Y(n5252));
XOR2X1   g0211(.A(n5252), .B(n5231), .Y(n5253));
MX2X1    g0212(.A(g2877), .B(n5253), .S0(g2879), .Y(n498));
MX2X1    g0213(.A(g2874), .B(g2861), .S0(g2879), .Y(n503));
MX2X1    g0214(.A(g2981), .B(g2864), .S0(g2879), .Y(n512));
MX2X1    g0215(.A(g2978), .B(g2867), .S0(g2879), .Y(n521));
MX2X1    g0216(.A(g2975), .B(g2870), .S0(g2879), .Y(n530));
MX2X1    g0217(.A(g2972), .B(g2818), .S0(g2879), .Y(n539));
MX2X1    g0218(.A(g2969), .B(g2821), .S0(g2879), .Y(n548));
MX2X1    g0219(.A(g2966), .B(g2824), .S0(g2879), .Y(n557));
MX2X1    g0220(.A(g2963), .B(g2827), .S0(g2879), .Y(n566));
INVX1    g0221(.A(g2879), .Y(n5263));
XOR2X1   g0222(.A(n5252), .B(n5239), .Y(n5264));
MX2X1    g0223(.A(g2830), .B(n5264), .S0(n5263), .Y(n575));
MX2X1    g0224(.A(g2959), .B(g2833), .S0(g2879), .Y(n584));
MX2X1    g0225(.A(g2956), .B(g2836), .S0(g2879), .Y(n593));
MX2X1    g0226(.A(g2953), .B(g2839), .S0(g2879), .Y(n602));
MX2X1    g0227(.A(g2947), .B(g2842), .S0(g2879), .Y(n611));
MX2X1    g0228(.A(g2944), .B(g2845), .S0(g2879), .Y(n620));
MX2X1    g0229(.A(g2941), .B(g2848), .S0(g2879), .Y(n629));
MX2X1    g0230(.A(g2938), .B(g2851), .S0(g2879), .Y(n638));
MX2X1    g0231(.A(g2935), .B(g2854), .S0(g2879), .Y(n647));
MX2X1    g0232(.A(g2858), .B(n5253), .S0(n5263), .Y(n656));
MX2X1    g0233(.A(g2200), .B(g2874), .S0(g2879), .Y(n665));
MX2X1    g0234(.A(g2195), .B(g2981), .S0(g2879), .Y(n670));
MX2X1    g0235(.A(g2190), .B(g2978), .S0(g2879), .Y(n675));
MX2X1    g0236(.A(g2185), .B(g2975), .S0(g2879), .Y(n680));
MX2X1    g0237(.A(g2180), .B(g2972), .S0(g2879), .Y(n685));
MX2X1    g0238(.A(g2175), .B(g2969), .S0(g2879), .Y(n690));
MX2X1    g0239(.A(g2170), .B(g2966), .S0(g2879), .Y(n695));
MX2X1    g0240(.A(g2165), .B(g2963), .S0(g2879), .Y(n700));
MX2X1    g0241(.A(g2878), .B(n5264), .S0(g2879), .Y(n705));
MX2X1    g0242(.A(g3210), .B(g559), .S0(g3129), .Y(n723));
MX2X1    g0243(.A(g3211), .B(g559), .S0(g3117), .Y(n728));
MX2X1    g0244(.A(g3084), .B(g559), .S0(g3109), .Y(n733));
MX2X1    g0245(.A(g3085), .B(g1245), .S0(g3129), .Y(n738));
MX2X1    g0246(.A(g3086), .B(g1245), .S0(g3117), .Y(n743));
MX2X1    g0247(.A(g3087), .B(g1245), .S0(g3109), .Y(n748));
MX2X1    g0248(.A(g3091), .B(g1939), .S0(g3129), .Y(n753));
MX2X1    g0249(.A(g3092), .B(g1939), .S0(g3117), .Y(n758));
MX2X1    g0250(.A(g3093), .B(g1939), .S0(g3109), .Y(n763));
MX2X1    g0251(.A(g3094), .B(g2633), .S0(g3129), .Y(n768));
MX2X1    g0252(.A(g3095), .B(g2633), .S0(g3117), .Y(n773));
MX2X1    g0253(.A(g3096), .B(g2633), .S0(g3109), .Y(n778));
INVX1    g0254(.A(g499), .Y(n5296));
INVX1    g0255(.A(g545), .Y(n5297));
AND2X1   g0256(.A(g548), .B(n5297), .Y(n5298_1));
MX2X1    g0257(.A(g544), .B(n5298_1), .S0(n5296), .Y(n2204));
MX2X1    g0258(.A(g3097), .B(n2204), .S0(g3129), .Y(n783));
MX2X1    g0259(.A(g3098), .B(n2204), .S0(g3117), .Y(n788));
MX2X1    g0260(.A(g3099), .B(n2204), .S0(g3109), .Y(n793));
INVX1    g0261(.A(g1234), .Y(n5303));
INVX1    g0262(.A(g1186), .Y(n5304));
OAI21X1  g0263(.A0(n5303), .A1(g1231), .B0(n5304), .Y(n5305));
AOI21X1  g0264(.A0(n2204), .A1(g1231), .B0(n5305), .Y(n5306));
NOR2X1   g0265(.A(n5304), .B(g1230), .Y(n5307_1));
NOR2X1   g0266(.A(n5307_1), .B(n5306), .Y(n3905));
MX2X1    g0267(.A(g3100), .B(n3905), .S0(g3129), .Y(n798));
MX2X1    g0268(.A(g3101), .B(n3905), .S0(g3117), .Y(n803));
MX2X1    g0269(.A(g3102), .B(n3905), .S0(g3109), .Y(n808));
INVX1    g0270(.A(g1925), .Y(n5312));
NOR3X1   g0271(.A(n5307_1), .B(n5306), .C(n5312), .Y(n5313));
INVX1    g0272(.A(g1928), .Y(n5314));
INVX1    g0273(.A(g1880), .Y(n5315));
OAI21X1  g0274(.A0(n5314), .A1(g1925), .B0(n5315), .Y(n5316_1));
NOR2X1   g0275(.A(n5316_1), .B(n5313), .Y(n5317));
NOR2X1   g0276(.A(n5315), .B(g1924), .Y(n5318));
NOR2X1   g0277(.A(n5318), .B(n5317), .Y(n5606));
MX2X1    g0278(.A(g3103), .B(n5606), .S0(g3129), .Y(n813));
MX2X1    g0279(.A(g3104), .B(n5606), .S0(g3117), .Y(n818));
MX2X1    g0280(.A(g3105), .B(n5606), .S0(g3109), .Y(n823));
OR2X1    g0281(.A(n5316_1), .B(n5313), .Y(n5323));
INVX1    g0282(.A(n5318), .Y(n5324));
NAND3X1  g0283(.A(n5324), .B(n5323), .C(g2619), .Y(n5325_1));
INVX1    g0284(.A(g2619), .Y(n5326));
AOI21X1  g0285(.A0(g2622), .A1(n5326), .B0(g2574), .Y(n5327));
INVX1    g0286(.A(g2574), .Y(n5328));
NOR2X1   g0287(.A(n5328), .B(g2618), .Y(n5329_1));
AOI21X1  g0288(.A0(n5327), .A1(n5325_1), .B0(n5329_1), .Y(n7307));
MX2X1    g0289(.A(g3106), .B(n7307), .S0(g3129), .Y(n828));
MX2X1    g0290(.A(g3107), .B(n7307), .S0(g3117), .Y(n833));
MX2X1    g0291(.A(g3108), .B(n7307), .S0(g3109), .Y(n838));
MX2X1    g0292(.A(g3155), .B(g499), .S0(g3129), .Y(n843));
MX2X1    g0293(.A(g3158), .B(g499), .S0(g3117), .Y(n848));
MX2X1    g0294(.A(g3161), .B(g499), .S0(g3109), .Y(n853));
MX2X1    g0295(.A(g3164), .B(g1186), .S0(g3129), .Y(n858));
MX2X1    g0296(.A(g3167), .B(g1186), .S0(g3117), .Y(n863));
MX2X1    g0297(.A(g3170), .B(g1186), .S0(g3109), .Y(n868));
MX2X1    g0298(.A(g3173), .B(g1880), .S0(g3129), .Y(n873));
MX2X1    g0299(.A(g3176), .B(g1880), .S0(g3117), .Y(n878));
MX2X1    g0300(.A(g3179), .B(g1880), .S0(g3109), .Y(n883));
MX2X1    g0301(.A(g3182), .B(g2574), .S0(g3129), .Y(n888));
MX2X1    g0302(.A(g3185), .B(g2574), .S0(g3117), .Y(n893));
MX2X1    g0303(.A(g3088), .B(g2574), .S0(g3109), .Y(n898));
INVX1    g0304(.A(g24734), .Y(n978));
INVX1    g0305(.A(g97), .Y(n1795));
NAND2X1  g0306(.A(g181), .B(g138), .Y(n5348));
MX2X1    g0307(.A(n1795), .B(g130), .S0(n5348), .Y(n1066));
NAND2X1  g0308(.A(g181), .B(g135), .Y(n5350));
MX2X1    g0309(.A(n1795), .B(g131), .S0(n5350), .Y(n1071));
AND2X1   g0310(.A(g181), .B(g165), .Y(n5352_1));
MX2X1    g0311(.A(g129), .B(n1795), .S0(n5352_1), .Y(n1076));
INVX1    g0312(.A(g101), .Y(n1786));
MX2X1    g0313(.A(n1786), .B(g133), .S0(n5348), .Y(n1081));
MX2X1    g0314(.A(n1786), .B(g134), .S0(n5350), .Y(n1086));
MX2X1    g0315(.A(g132), .B(n1786), .S0(n5352_1), .Y(n1091));
INVX1    g0316(.A(g105), .Y(n1777));
MX2X1    g0317(.A(n1777), .B(g142), .S0(n5348), .Y(n1096));
MX2X1    g0318(.A(n1777), .B(g143), .S0(n5350), .Y(n1101));
MX2X1    g0319(.A(g141), .B(n1777), .S0(n5352_1), .Y(n1106));
INVX1    g0320(.A(g109), .Y(n1768));
MX2X1    g0321(.A(n1768), .B(g145), .S0(n5348), .Y(n1111));
MX2X1    g0322(.A(n1768), .B(g146), .S0(n5350), .Y(n1116));
MX2X1    g0323(.A(g144), .B(n1768), .S0(n5352_1), .Y(n1121));
INVX1    g0324(.A(g113), .Y(n1759));
MX2X1    g0325(.A(n1759), .B(g148), .S0(n5348), .Y(n1126));
MX2X1    g0326(.A(n1759), .B(g149), .S0(n5350), .Y(n1131));
MX2X1    g0327(.A(g147), .B(n1759), .S0(n5352_1), .Y(n1136));
INVX1    g0328(.A(g117), .Y(n1750));
MX2X1    g0329(.A(n1750), .B(g151), .S0(n5348), .Y(n1141));
MX2X1    g0330(.A(n1750), .B(g152), .S0(n5350), .Y(n1146));
MX2X1    g0331(.A(g150), .B(n1750), .S0(n5352_1), .Y(n1151));
INVX1    g0332(.A(g121), .Y(n1741));
MX2X1    g0333(.A(n1741), .B(g154), .S0(n5348), .Y(n1156));
MX2X1    g0334(.A(n1741), .B(g155), .S0(n5350), .Y(n1161));
MX2X1    g0335(.A(g153), .B(n1741), .S0(n5352_1), .Y(n1166));
INVX1    g0336(.A(g125), .Y(n1732));
MX2X1    g0337(.A(n1732), .B(g157), .S0(n5348), .Y(n1171));
MX2X1    g0338(.A(n1732), .B(g158), .S0(n5350), .Y(n1176));
MX2X1    g0339(.A(g156), .B(n1732), .S0(n5352_1), .Y(n1181));
INVX1    g0340(.A(g138), .Y(n5382));
NOR2X1   g0341(.A(g175), .B(n5382), .Y(n5383_1));
INVX1    g0342(.A(g135), .Y(n5384));
INVX1    g0343(.A(g165), .Y(n5385));
OAI22X1  g0344(.A0(g176), .A1(n5384), .B0(n5385), .B1(g174), .Y(n5386));
NOR2X1   g0345(.A(n5386), .B(n5383_1), .Y(n5387));
MX2X1    g0346(.A(n5387), .B(g160), .S0(n5348), .Y(n1186));
MX2X1    g0347(.A(n5387), .B(g161), .S0(n5350), .Y(n1191));
MX2X1    g0348(.A(g159), .B(n5387), .S0(n5352_1), .Y(n1196));
NOR2X1   g0349(.A(g172), .B(n5382), .Y(n5391));
OAI22X1  g0350(.A0(g173), .A1(n5384), .B0(n5385), .B1(g171), .Y(n5392_1));
NOR2X1   g0351(.A(n5392_1), .B(n5391), .Y(n5393));
MX2X1    g0352(.A(n5393), .B(g163), .S0(n5348), .Y(n1201));
MX2X1    g0353(.A(n5393), .B(g164), .S0(n5350), .Y(n1206));
MX2X1    g0354(.A(g162), .B(n5393), .S0(n5352_1), .Y(n1211));
NOR4X1   g0355(.A(g117), .B(g121), .C(n1732), .D(n1759), .Y(n5397));
OR2X1    g0356(.A(g2900), .B(g2892), .Y(n5398));
NOR4X1   g0357(.A(g2908), .B(g2903), .C(g2896), .D(n5398), .Y(n5399));
NAND4X1  g0358(.A(g2924), .B(n5209), .C(g2883), .D(n5211), .Y(n5400));
NOR3X1   g0359(.A(n5400), .B(g2917), .C(g2888), .Y(n5401_1));
AND2X1   g0360(.A(n5401_1), .B(n5399), .Y(n1476));
AND2X1   g0361(.A(n1476), .B(g138), .Y(n5403));
MX2X1    g0362(.A(g169), .B(n5397), .S0(n5403), .Y(n1216));
AND2X1   g0363(.A(n1476), .B(g135), .Y(n5405_1));
MX2X1    g0364(.A(g170), .B(n5397), .S0(n5405_1), .Y(n1221));
AND2X1   g0365(.A(n1476), .B(g165), .Y(n5407));
MX2X1    g0366(.A(g168), .B(n5397), .S0(n5407), .Y(n1226));
MX2X1    g0367(.A(g172), .B(n1786), .S0(n5403), .Y(n1231));
MX2X1    g0368(.A(g173), .B(n1786), .S0(n5405_1), .Y(n1236));
MX2X1    g0369(.A(g171), .B(n1786), .S0(n5407), .Y(n1241));
MX2X1    g0370(.A(g175), .B(n1795), .S0(n5403), .Y(n1246));
MX2X1    g0371(.A(g176), .B(n1795), .S0(n5405_1), .Y(n1251));
MX2X1    g0372(.A(g174), .B(n1795), .S0(n5407), .Y(n1256));
NAND4X1  g0373(.A(g101), .B(g105), .C(g125), .D(g97), .Y(n5415));
NAND4X1  g0374(.A(g113), .B(g117), .C(g121), .D(g109), .Y(n5416));
NOR2X1   g0375(.A(n5416), .B(n5415), .Y(n5417));
INVX1    g0376(.A(n5417), .Y(n5418));
MX2X1    g0377(.A(g178), .B(n5418), .S0(n5403), .Y(n1261));
MX2X1    g0378(.A(g179), .B(n5418), .S0(n5405_1), .Y(n1266));
MX2X1    g0379(.A(g177), .B(n5418), .S0(n5407), .Y(n1271));
NOR2X1   g0380(.A(g163), .B(n5382), .Y(n5422));
OAI22X1  g0381(.A0(g164), .A1(n5384), .B0(n5385), .B1(g162), .Y(n5423));
OR2X1    g0382(.A(n5423), .B(n5422), .Y(n5424_1));
AND2X1   g0383(.A(n5424_1), .B(n5393), .Y(n5425));
NOR2X1   g0384(.A(g169), .B(n5382), .Y(n5426));
OAI22X1  g0385(.A0(g170), .A1(n5384), .B0(n5385), .B1(g168), .Y(n5427));
OAI21X1  g0386(.A0(n5427), .A1(n5426), .B0(g181), .Y(n5428));
NOR2X1   g0387(.A(g160), .B(n5382), .Y(n5429_1));
OAI22X1  g0388(.A0(g161), .A1(n5384), .B0(n5385), .B1(g159), .Y(n5430));
NOR2X1   g0389(.A(n5430), .B(n5429_1), .Y(n5431));
XOR2X1   g0390(.A(n5431), .B(n5387), .Y(n5432));
NOR2X1   g0391(.A(g154), .B(n5382), .Y(n5433_1));
OAI22X1  g0392(.A0(g155), .A1(n5384), .B0(n5385), .B1(g153), .Y(n5434));
NOR2X1   g0393(.A(n5434), .B(n5433_1), .Y(n5435));
XOR2X1   g0394(.A(n5435), .B(n1741), .Y(n5436));
NOR4X1   g0395(.A(n5432), .B(n5428), .C(n5425), .D(n5436), .Y(n5437_1));
NOR2X1   g0396(.A(g148), .B(n5382), .Y(n5438));
OAI22X1  g0397(.A0(g149), .A1(n5384), .B0(n5385), .B1(g147), .Y(n5439));
NOR2X1   g0398(.A(n5439), .B(n5438), .Y(n5440));
XOR2X1   g0399(.A(n5440), .B(n1759), .Y(n5441));
NOR2X1   g0400(.A(g145), .B(n5382), .Y(n5442_1));
OAI22X1  g0401(.A0(g146), .A1(n5384), .B0(n5385), .B1(g144), .Y(n5443));
NOR2X1   g0402(.A(n5443), .B(n5442_1), .Y(n5444));
XOR2X1   g0403(.A(n5444), .B(n1768), .Y(n5445));
NOR2X1   g0404(.A(g151), .B(n5382), .Y(n5446_1));
OAI22X1  g0405(.A0(g152), .A1(n5384), .B0(n5385), .B1(g150), .Y(n5447));
NOR2X1   g0406(.A(n5447), .B(n5446_1), .Y(n5448));
XOR2X1   g0407(.A(n5448), .B(n1750), .Y(n5449));
NOR2X1   g0408(.A(g157), .B(n5382), .Y(n5450));
OAI22X1  g0409(.A0(g158), .A1(n5384), .B0(n5385), .B1(g156), .Y(n5451_1));
OAI21X1  g0410(.A0(n5451_1), .A1(n5450), .B0(n1732), .Y(n5452));
OAI21X1  g0411(.A0(n5424_1), .A1(n5393), .B0(n5452), .Y(n5453));
NOR4X1   g0412(.A(n5449), .B(n5445), .C(n5441), .D(n5453), .Y(n5454));
NOR3X1   g0413(.A(n5451_1), .B(n5450), .C(n1732), .Y(n5455_1));
NOR2X1   g0414(.A(g142), .B(n5382), .Y(n5456));
OAI22X1  g0415(.A0(g143), .A1(n5384), .B0(n5385), .B1(g141), .Y(n5457));
NOR2X1   g0416(.A(n5457), .B(n5456), .Y(n5458));
XOR2X1   g0417(.A(n5458), .B(n1777), .Y(n5459));
NOR2X1   g0418(.A(g133), .B(n5382), .Y(n5460_1));
OAI22X1  g0419(.A0(g134), .A1(n5384), .B0(n5385), .B1(g132), .Y(n5461));
NOR2X1   g0420(.A(n5461), .B(n5460_1), .Y(n5462));
XOR2X1   g0421(.A(n5462), .B(n1786), .Y(n5463));
NOR2X1   g0422(.A(g130), .B(n5382), .Y(n5464_1));
OAI22X1  g0423(.A0(g131), .A1(n5384), .B0(n5385), .B1(g129), .Y(n5465));
NOR2X1   g0424(.A(n5465), .B(n5464_1), .Y(n5466));
XOR2X1   g0425(.A(n5466), .B(n1795), .Y(n5467));
NOR4X1   g0426(.A(n5463), .B(n5459), .C(n5455_1), .D(n5467), .Y(n5468));
NAND3X1  g0427(.A(n5468), .B(n5454), .C(n5437_1), .Y(n5469_1));
NAND2X1  g0428(.A(g222), .B(g138), .Y(n5470));
AOI22X1  g0429(.A0(g225), .A1(g135), .B0(g165), .B1(g228), .Y(n5471));
AND2X1   g0430(.A(n5471), .B(n5470), .Y(n5472));
NOR3X1   g0431(.A(n5472), .B(n5386), .C(n5383_1), .Y(n5473_1));
OR2X1    g0432(.A(g175), .B(n5382), .Y(n5474));
INVX1    g0433(.A(g176), .Y(n5475));
INVX1    g0434(.A(g174), .Y(n5476));
AOI22X1  g0435(.A0(n5475), .A1(g135), .B0(g165), .B1(n5476), .Y(n5477));
NAND2X1  g0436(.A(n5471), .B(n5470), .Y(n5478_1));
AOI21X1  g0437(.A0(n5477), .A1(n5474), .B0(n5478_1), .Y(n5479));
NAND2X1  g0438(.A(g213), .B(g138), .Y(n5480));
AOI22X1  g0439(.A0(g216), .A1(g135), .B0(g165), .B1(g219), .Y(n5481));
NAND2X1  g0440(.A(n5481), .B(n5480), .Y(n5482_1));
XOR2X1   g0441(.A(n5482_1), .B(g121), .Y(n5483));
NOR3X1   g0442(.A(n5483), .B(n5479), .C(n5473_1), .Y(n5484));
NAND2X1  g0443(.A(g186), .B(g138), .Y(n5485));
AOI22X1  g0444(.A0(g189), .A1(g135), .B0(g165), .B1(g192), .Y(n5486));
NAND2X1  g0445(.A(n5486), .B(n5485), .Y(n5487_1));
XOR2X1   g0446(.A(n5487_1), .B(g97), .Y(n5488));
NAND2X1  g0447(.A(g195), .B(g138), .Y(n5489));
AOI22X1  g0448(.A0(g198), .A1(g135), .B0(g165), .B1(g201), .Y(n5490));
NAND2X1  g0449(.A(n5490), .B(n5489), .Y(n5491_1));
XOR2X1   g0450(.A(n5491_1), .B(g105), .Y(n5492));
NAND2X1  g0451(.A(g204), .B(g138), .Y(n5493));
AOI22X1  g0452(.A0(g207), .A1(g135), .B0(g165), .B1(g210), .Y(n5494));
NAND2X1  g0453(.A(n5494), .B(n5493), .Y(n5495));
XOR2X1   g0454(.A(n5495), .B(g113), .Y(n5496_1));
OAI21X1  g0455(.A0(n5496_1), .A1(n5492), .B0(n5488), .Y(n5497));
NOR2X1   g0456(.A(n5497), .B(n5484), .Y(n5498));
NOR2X1   g0457(.A(n5496_1), .B(n5483), .Y(n5499));
OAI22X1  g0458(.A0(n5488), .A1(n5492), .B0(n5479), .B1(n5473_1), .Y(n5500_1));
NOR2X1   g0459(.A(n5500_1), .B(n5499), .Y(n5501));
XOR2X1   g0460(.A(n5495), .B(n1759), .Y(n5502));
NOR2X1   g0461(.A(n5488), .B(n5483), .Y(n5503));
NOR3X1   g0462(.A(n5492), .B(n5479), .C(n5473_1), .Y(n5504_1));
NOR3X1   g0463(.A(n5504_1), .B(n5503), .C(n5502), .Y(n5505));
NOR3X1   g0464(.A(n5505), .B(n5501), .C(n5498), .Y(n5506));
NAND2X1  g0465(.A(g267), .B(g138), .Y(n5507));
AOI22X1  g0466(.A0(g270), .A1(g135), .B0(g165), .B1(g273), .Y(n5508));
AND2X1   g0467(.A(n5508), .B(n5507), .Y(n5509_1));
NOR3X1   g0468(.A(n5509_1), .B(n5392_1), .C(n5391), .Y(n5510));
OR2X1    g0469(.A(g172), .B(n5382), .Y(n5511));
INVX1    g0470(.A(g173), .Y(n5512));
INVX1    g0471(.A(g171), .Y(n5513));
AOI22X1  g0472(.A0(n5512), .A1(g135), .B0(g165), .B1(n5513), .Y(n5514_1));
NAND2X1  g0473(.A(n5508), .B(n5507), .Y(n5515));
AOI21X1  g0474(.A0(n5514_1), .A1(n5511), .B0(n5515), .Y(n5516));
NAND2X1  g0475(.A(g258), .B(g138), .Y(n5517));
AOI22X1  g0476(.A0(g261), .A1(g135), .B0(g165), .B1(g264), .Y(n5518));
NAND2X1  g0477(.A(n5518), .B(n5517), .Y(n5519_1));
XOR2X1   g0478(.A(n5519_1), .B(g125), .Y(n5520));
NOR3X1   g0479(.A(n5520), .B(n5516), .C(n5510), .Y(n5521));
NAND2X1  g0480(.A(g231), .B(g138), .Y(n5522));
AOI22X1  g0481(.A0(g234), .A1(g135), .B0(g165), .B1(g237), .Y(n5523));
NAND2X1  g0482(.A(n5523), .B(n5522), .Y(n5524_1));
XOR2X1   g0483(.A(n5524_1), .B(g101), .Y(n5525));
NAND2X1  g0484(.A(g240), .B(g138), .Y(n5526));
AOI22X1  g0485(.A0(g243), .A1(g135), .B0(g165), .B1(g246), .Y(n5527));
NAND2X1  g0486(.A(n5527), .B(n5526), .Y(n5528));
XOR2X1   g0487(.A(n5528), .B(g109), .Y(n5529_1));
NAND2X1  g0488(.A(g249), .B(g138), .Y(n5530));
AOI22X1  g0489(.A0(g252), .A1(g135), .B0(g165), .B1(g255), .Y(n5531));
NAND2X1  g0490(.A(n5531), .B(n5530), .Y(n5532));
XOR2X1   g0491(.A(n5532), .B(g117), .Y(n5533));
OAI21X1  g0492(.A0(n5533), .A1(n5529_1), .B0(n5525), .Y(n5534_1));
NOR2X1   g0493(.A(n5534_1), .B(n5521), .Y(n5535));
NOR2X1   g0494(.A(n5533), .B(n5520), .Y(n5536));
OAI22X1  g0495(.A0(n5525), .A1(n5529_1), .B0(n5516), .B1(n5510), .Y(n5537));
NOR2X1   g0496(.A(n5537), .B(n5536), .Y(n5538));
XOR2X1   g0497(.A(n5532), .B(n1750), .Y(n5539_1));
NOR2X1   g0498(.A(n5525), .B(n5520), .Y(n5540));
NOR3X1   g0499(.A(n5529_1), .B(n5516), .C(n5510), .Y(n5541));
NOR3X1   g0500(.A(n5541), .B(n5540), .C(n5539_1), .Y(n5542));
NOR3X1   g0501(.A(n5542), .B(n5538), .C(n5535), .Y(n5543));
AOI21X1  g0502(.A0(n5543), .A1(n5506), .B0(n5428), .Y(n5544_1));
INVX1    g0503(.A(g276), .Y(n5545));
NOR2X1   g0504(.A(g318), .B(n5545), .Y(n5546));
INVX1    g0505(.A(g405), .Y(n5547));
INVX1    g0506(.A(g401), .Y(n5548));
OAI22X1  g0507(.A0(g319), .A1(n5547), .B0(n5548), .B1(g320), .Y(n5549_1));
NOR2X1   g0508(.A(n5549_1), .B(n5546), .Y(n5550));
NOR2X1   g0509(.A(g315), .B(n5545), .Y(n5551));
OAI22X1  g0510(.A0(g316), .A1(n5547), .B0(n5548), .B1(g317), .Y(n5552));
NOR2X1   g0511(.A(n5552), .B(n5551), .Y(n5553));
NOR2X1   g0512(.A(g312), .B(n5545), .Y(n5554_1));
OAI22X1  g0513(.A0(g313), .A1(n5547), .B0(n5548), .B1(g314), .Y(n5555));
NOR2X1   g0514(.A(n5555), .B(n5554_1), .Y(n5556));
INVX1    g0515(.A(n5556), .Y(n5557));
NOR2X1   g0516(.A(g322), .B(n5545), .Y(n5558));
OAI22X1  g0517(.A0(g323), .A1(n5547), .B0(n5548), .B1(g321), .Y(n5559_1));
NOR2X1   g0518(.A(n5559_1), .B(n5558), .Y(n5560));
INVX1    g0519(.A(n5560), .Y(n5561));
NAND4X1  g0520(.A(n5557), .B(n5553), .C(n5550), .D(n5561), .Y(n5562));
NOR3X1   g0521(.A(n5562), .B(n5544_1), .C(n5469_1), .Y(n5563));
NOR4X1   g0522(.A(n5552), .B(n5551), .C(n5550), .D(n5556), .Y(n5564_1));
NAND2X1  g0523(.A(n5564_1), .B(n5561), .Y(n5565));
NOR2X1   g0524(.A(n5565), .B(n5469_1), .Y(n5566));
NOR2X1   g0525(.A(g403), .B(n5545), .Y(n5567));
OAI22X1  g0526(.A0(g404), .A1(n5547), .B0(n5548), .B1(g402), .Y(n5568));
NOR2X1   g0527(.A(n5568), .B(n5567), .Y(n5569_1));
INVX1    g0528(.A(g181), .Y(n5570));
NOR3X1   g0529(.A(n5427), .B(n5426), .C(n5570), .Y(n5571));
INVX1    g0530(.A(n5571), .Y(n5572));
OAI22X1  g0531(.A0(n5569_1), .A1(n5469_1), .B0(n5556), .B1(n5572), .Y(n5573));
OR4X1    g0532(.A(n5551), .B(n5549_1), .C(n5546), .D(n5552), .Y(n5574_1));
NOR3X1   g0533(.A(n5555), .B(n5554_1), .C(n5574_1), .Y(n5575));
INVX1    g0534(.A(n5575), .Y(n5576));
INVX1    g0535(.A(n5553), .Y(n5577));
NAND3X1  g0536(.A(n5556), .B(n5577), .C(n5550), .Y(n5578));
INVX1    g0537(.A(n5550), .Y(n5579_1));
NOR3X1   g0538(.A(n5557), .B(n5553), .C(n5579_1), .Y(n5580));
NAND4X1  g0539(.A(n5493), .B(n5481), .C(n5480), .D(n5494), .Y(n5581));
OR4X1    g0540(.A(n5532), .B(n5519_1), .C(n5487_1), .D(n5581), .Y(n5582));
NAND4X1  g0541(.A(n5489), .B(n5471), .C(n5470), .D(n5490), .Y(n5583));
OR4X1    g0542(.A(n5528), .B(n5524_1), .C(n5515), .D(n5583), .Y(n5584_1));
OR2X1    g0543(.A(n5584_1), .B(n5582), .Y(n5585));
OR2X1    g0544(.A(n5585), .B(n5580), .Y(n5586));
NAND2X1  g0545(.A(n5528), .B(n5515), .Y(n5587));
NAND3X1  g0546(.A(n5524_1), .B(n5491_1), .C(n5478_1), .Y(n5588_1));
OR4X1    g0547(.A(n5587), .B(n5582), .C(n5578), .D(n5588_1), .Y(n5589));
AOI22X1  g0548(.A0(n5586), .A1(n5589), .B0(n5578), .B1(n5576), .Y(n5590));
NOR4X1   g0549(.A(n5573), .B(n5566), .C(n5563), .D(n5590), .Y(n5591));
INVX1    g0550(.A(n5591), .Y(n5592_1));
NAND2X1  g0551(.A(n5578), .B(n5576), .Y(n5593));
XOR2X1   g0552(.A(n5593), .B(n5487_1), .Y(n5594));
NOR3X1   g0553(.A(n5573), .B(n5566), .C(n5563), .Y(n5595));
AOI21X1  g0554(.A0(n5590), .A1(n5595), .B0(n1795), .Y(n5596));
MX2X1    g0555(.A(n5594), .B(n5596), .S0(n5592_1), .Y(n5597_1));
MX2X1    g0556(.A(g186), .B(n5597_1), .S0(g138), .Y(n1276));
MX2X1    g0557(.A(g189), .B(n5597_1), .S0(g135), .Y(n1281));
MX2X1    g0558(.A(g192), .B(n5597_1), .S0(g165), .Y(n1286));
AND2X1   g0559(.A(n5578), .B(n5487_1), .Y(n5601_1));
OAI21X1  g0560(.A0(n5578), .A1(n5487_1), .B0(n5593), .Y(n5602));
OR2X1    g0561(.A(n5602), .B(n5601_1), .Y(n5603));
XOR2X1   g0562(.A(n5603), .B(n5524_1), .Y(n5604));
NAND3X1  g0563(.A(n5590), .B(n5578), .C(n5595), .Y(n5605));
MX2X1    g0564(.A(n1786), .B(n5590), .S0(n5595), .Y(n5606_1));
AOI22X1  g0565(.A0(n5605), .A1(n5606_1), .B0(n5604), .B1(n5591), .Y(n5607));
MX2X1    g0566(.A(g231), .B(n5607), .S0(g138), .Y(n1291));
MX2X1    g0567(.A(g234), .B(n5607), .S0(g135), .Y(n1296));
MX2X1    g0568(.A(g237), .B(n5607), .S0(g165), .Y(n1301));
XOR2X1   g0569(.A(n5580), .B(n5524_1), .Y(n5611_1));
OR2X1    g0570(.A(n5611_1), .B(n5603), .Y(n5612));
XOR2X1   g0571(.A(n5612), .B(n5491_1), .Y(n5613));
MX2X1    g0572(.A(n1777), .B(n5590), .S0(n5595), .Y(n5614));
AOI22X1  g0573(.A0(n5613), .A1(n5591), .B0(n5605), .B1(n5614), .Y(n5615_1));
MX2X1    g0574(.A(g195), .B(n5615_1), .S0(g138), .Y(n1306));
MX2X1    g0575(.A(g198), .B(n5615_1), .S0(g135), .Y(n1311));
MX2X1    g0576(.A(g201), .B(n5615_1), .S0(g165), .Y(n1316));
XOR2X1   g0577(.A(n5580), .B(n5491_1), .Y(n5619));
OR4X1    g0578(.A(n5611_1), .B(n5602), .C(n5601_1), .D(n5619), .Y(n5620_1));
XOR2X1   g0579(.A(n5620_1), .B(n5528), .Y(n5621));
MX2X1    g0580(.A(n1768), .B(n5590), .S0(n5595), .Y(n5622));
AOI22X1  g0581(.A0(n5621), .A1(n5591), .B0(n5605), .B1(n5622), .Y(n5623));
MX2X1    g0582(.A(g240), .B(n5623), .S0(g138), .Y(n1321));
MX2X1    g0583(.A(g243), .B(n5623), .S0(g135), .Y(n1326));
MX2X1    g0584(.A(g246), .B(n5623), .S0(g165), .Y(n1331));
XOR2X1   g0585(.A(n5580), .B(n5528), .Y(n5627));
OR2X1    g0586(.A(n5627), .B(n5619), .Y(n5628));
NOR4X1   g0587(.A(n5611_1), .B(n5602), .C(n5601_1), .D(n5628), .Y(n5629_1));
XOR2X1   g0588(.A(n5629_1), .B(n5495), .Y(n5630));
AOI21X1  g0589(.A0(n5590), .A1(n5595), .B0(n1759), .Y(n5631));
MX2X1    g0590(.A(n5630), .B(n5631), .S0(n5592_1), .Y(n5632));
MX2X1    g0591(.A(g204), .B(n5632), .S0(g138), .Y(n1336));
MX2X1    g0592(.A(g207), .B(n5632), .S0(g135), .Y(n1341));
MX2X1    g0593(.A(g210), .B(n5632), .S0(g165), .Y(n1346));
XOR2X1   g0594(.A(n5578), .B(n5495), .Y(n5636));
AND2X1   g0595(.A(n5636), .B(n5629_1), .Y(n5637));
XOR2X1   g0596(.A(n5637), .B(n5532), .Y(n5638));
AOI21X1  g0597(.A0(n5590), .A1(n5595), .B0(n1750), .Y(n5639_1));
MX2X1    g0598(.A(n5638), .B(n5639_1), .S0(n5592_1), .Y(n5640));
MX2X1    g0599(.A(g249), .B(n5640), .S0(g138), .Y(n1351));
MX2X1    g0600(.A(g252), .B(n5640), .S0(g135), .Y(n1356));
MX2X1    g0601(.A(g255), .B(n5640), .S0(g165), .Y(n1361));
XOR2X1   g0602(.A(n5578), .B(n5532), .Y(n5644_1));
NAND2X1  g0603(.A(n5644_1), .B(n5636), .Y(n5645));
NOR4X1   g0604(.A(n5628), .B(n5611_1), .C(n5603), .D(n5645), .Y(n5646));
XOR2X1   g0605(.A(n5646), .B(n5482_1), .Y(n5647));
AOI21X1  g0606(.A0(n5590), .A1(n5595), .B0(n1741), .Y(n5648));
MX2X1    g0607(.A(n5647), .B(n5648), .S0(n5592_1), .Y(n5649_1));
MX2X1    g0608(.A(g213), .B(n5649_1), .S0(g138), .Y(n1366));
MX2X1    g0609(.A(g216), .B(n5649_1), .S0(g135), .Y(n1371));
MX2X1    g0610(.A(g219), .B(n5649_1), .S0(g165), .Y(n1376));
XOR2X1   g0611(.A(n5578), .B(n5482_1), .Y(n5653));
AND2X1   g0612(.A(n5653), .B(n5646), .Y(n5654_1));
XOR2X1   g0613(.A(n5654_1), .B(n5519_1), .Y(n5655));
AOI21X1  g0614(.A0(n5590), .A1(n5595), .B0(n1732), .Y(n5656));
MX2X1    g0615(.A(n5655), .B(n5656), .S0(n5592_1), .Y(n5657));
MX2X1    g0616(.A(g258), .B(n5657), .S0(g138), .Y(n1381));
MX2X1    g0617(.A(g261), .B(n5657), .S0(g135), .Y(n1386));
MX2X1    g0618(.A(g264), .B(n5657), .S0(g165), .Y(n1391));
XOR2X1   g0619(.A(n5578), .B(n5519_1), .Y(n5661));
NAND4X1  g0620(.A(n5653), .B(n5644_1), .C(n5636), .D(n5661), .Y(n5662));
OR4X1    g0621(.A(n5628), .B(n5611_1), .C(n5603), .D(n5662), .Y(n5663));
XOR2X1   g0622(.A(n5663), .B(n5478_1), .Y(n5664_1));
MX2X1    g0623(.A(n5387), .B(n5590), .S0(n5595), .Y(n5665));
AOI22X1  g0624(.A0(n5664_1), .A1(n5591), .B0(n5605), .B1(n5665), .Y(n5666));
MX2X1    g0625(.A(g222), .B(n5666), .S0(g138), .Y(n1396));
MX2X1    g0626(.A(g225), .B(n5666), .S0(g135), .Y(n1401));
MX2X1    g0627(.A(g228), .B(n5666), .S0(g165), .Y(n1406));
XOR2X1   g0628(.A(n5580), .B(n5478_1), .Y(n5670));
OR2X1    g0629(.A(n5670), .B(n5663), .Y(n5671));
XOR2X1   g0630(.A(n5671), .B(n5515), .Y(n5672));
MX2X1    g0631(.A(n5393), .B(n5590), .S0(n5595), .Y(n5673));
AOI22X1  g0632(.A0(n5672), .A1(n5591), .B0(n5605), .B1(n5673), .Y(n5674_1));
MX2X1    g0633(.A(g267), .B(n5674_1), .S0(g138), .Y(n1411));
MX2X1    g0634(.A(g270), .B(n5674_1), .S0(g135), .Y(n1416));
MX2X1    g0635(.A(g273), .B(n5674_1), .S0(g165), .Y(n1421));
INVX1    g0636(.A(g92), .Y(n5678));
NOR2X1   g0637(.A(n5399), .B(n5385), .Y(n5679_1));
XOR2X1   g0638(.A(n5679_1), .B(n5678), .Y(n5680));
AOI21X1  g0639(.A0(n5399), .A1(n5352_1), .B0(n5680), .Y(n1426));
INVX1    g0640(.A(g88), .Y(n5682));
NOR3X1   g0641(.A(n5399), .B(n5678), .C(n5385), .Y(n5683));
XOR2X1   g0642(.A(n5683), .B(n5682), .Y(n5684_1));
AOI21X1  g0643(.A0(n5399), .A1(n5352_1), .B0(n5684_1), .Y(n1431));
INVX1    g0644(.A(g83), .Y(n5686));
NOR4X1   g0645(.A(n5682), .B(n5678), .C(n5385), .D(n5399), .Y(n5687));
XOR2X1   g0646(.A(n5687), .B(n5686), .Y(n5688));
AOI21X1  g0647(.A0(n5399), .A1(n5352_1), .B0(n5688), .Y(n1436));
NAND2X1  g0648(.A(n5687), .B(g83), .Y(n5690));
XOR2X1   g0649(.A(n5690), .B(g79), .Y(n5691));
AOI21X1  g0650(.A0(n5399), .A1(n5352_1), .B0(n5691), .Y(n1441));
NAND3X1  g0651(.A(n5687), .B(g79), .C(g83), .Y(n5693));
XOR2X1   g0652(.A(n5693), .B(g74), .Y(n5694_1));
AOI21X1  g0653(.A0(n5399), .A1(n5352_1), .B0(n5694_1), .Y(n1446));
INVX1    g0654(.A(g79), .Y(n5696));
INVX1    g0655(.A(g74), .Y(n5697));
OR4X1    g0656(.A(g70), .B(n5697), .C(n5696), .D(n5690), .Y(n5698));
OAI21X1  g0657(.A0(n5693), .A1(n5697), .B0(g70), .Y(n5699_1));
AOI22X1  g0658(.A0(n5698), .A1(n5699_1), .B0(n5399), .B1(n5352_1), .Y(n1451));
INVX1    g0659(.A(g70), .Y(n5701));
OR4X1    g0660(.A(n5701), .B(n5697), .C(n5696), .D(n5690), .Y(n5702));
XOR2X1   g0661(.A(n5702), .B(g65), .Y(n5703));
AOI21X1  g0662(.A0(n5399), .A1(n5352_1), .B0(n5703), .Y(n1456));
INVX1    g0663(.A(g61), .Y(n5705));
INVX1    g0664(.A(g65), .Y(n5706));
NOR4X1   g0665(.A(n5706), .B(n5701), .C(n5697), .D(n5693), .Y(n5707));
XOR2X1   g0666(.A(n5707), .B(n5705), .Y(n5708));
AOI21X1  g0667(.A0(n5399), .A1(n5352_1), .B0(n5708), .Y(n1461));
INVX1    g0668(.A(g56), .Y(n5710));
AND2X1   g0669(.A(n5707), .B(g61), .Y(n5711));
XOR2X1   g0670(.A(n5711), .B(n5710), .Y(n5712));
AOI21X1  g0671(.A0(n5399), .A1(n5352_1), .B0(n5712), .Y(n1466));
INVX1    g0672(.A(g52), .Y(n5714_1));
NOR4X1   g0673(.A(n5710), .B(n5705), .C(n5706), .D(n5702), .Y(n5715));
XOR2X1   g0674(.A(n5715), .B(n5714_1), .Y(n5716));
AOI21X1  g0675(.A0(n5399), .A1(n5352_1), .B0(n5716), .Y(n1471));
INVX1    g0676(.A(g3229), .Y(n5718));
NOR2X1   g0677(.A(g384), .B(n5545), .Y(n5719_1));
OAI22X1  g0678(.A0(g373), .A1(n5547), .B0(n5548), .B1(g376), .Y(n5720));
NOR2X1   g0679(.A(g369), .B(n5545), .Y(n5721));
OAI22X1  g0680(.A0(g358), .A1(n5547), .B0(n5548), .B1(g361), .Y(n5722));
NOR2X1   g0681(.A(n5722), .B(n5721), .Y(n5723));
OR4X1    g0682(.A(n5720), .B(n5719_1), .C(g3229), .D(n5723), .Y(n5724_1));
NOR2X1   g0683(.A(g398), .B(n5545), .Y(n5725));
OAI22X1  g0684(.A0(g388), .A1(n5547), .B0(n5548), .B1(g391), .Y(n5726));
NOR2X1   g0685(.A(n5726), .B(n5725), .Y(n5727));
OAI21X1  g0686(.A0(n5727), .A1(n5718), .B0(n5724_1), .Y(n5728));
INVX1    g0687(.A(n5723), .Y(n1853));
INVX1    g0688(.A(n5727), .Y(n1863));
NOR2X1   g0689(.A(g354), .B(n5545), .Y(n5731));
OAI22X1  g0690(.A0(g343), .A1(n5547), .B0(n5548), .B1(g346), .Y(n5732));
NOR2X1   g0691(.A(n5732), .B(n5731), .Y(n5733));
NOR4X1   g0692(.A(n1863), .B(n1853), .C(n5718), .D(n5733), .Y(n5734_1));
NOR4X1   g0693(.A(n5726), .B(n5725), .C(g3229), .D(n5733), .Y(n5735));
NOR2X1   g0694(.A(n5720), .B(n5719_1), .Y(n5736));
NOR3X1   g0695(.A(n5733), .B(n5736), .C(n5718), .Y(n5737));
NOR4X1   g0696(.A(n5735), .B(n5734_1), .C(n5728), .D(n5737), .Y(n5738));
NOR4X1   g0697(.A(n5554_1), .B(n5553), .C(n5550), .D(n5555), .Y(n5739_1));
AOI21X1  g0698(.A0(n5576), .A1(n5399), .B0(n5739_1), .Y(n1868));
AND2X1   g0699(.A(n1868), .B(g276), .Y(n5741));
MX2X1    g0700(.A(g354), .B(n5738), .S0(n5741), .Y(n1507));
AND2X1   g0701(.A(n1868), .B(g405), .Y(n5743));
MX2X1    g0702(.A(g343), .B(n5738), .S0(n5743), .Y(n1512));
AND2X1   g0703(.A(n1868), .B(g401), .Y(n5745));
MX2X1    g0704(.A(g346), .B(n5738), .S0(n5745), .Y(n1517));
NOR4X1   g0705(.A(n5731), .B(n5736), .C(g3229), .D(n5732), .Y(n5747));
NOR3X1   g0706(.A(n5723), .B(n5720), .C(n5719_1), .Y(n5748));
NOR3X1   g0707(.A(n5748), .B(n5747), .C(n5737), .Y(n5749_1));
MX2X1    g0708(.A(g369), .B(n5749_1), .S0(n5741), .Y(n1522));
MX2X1    g0709(.A(g358), .B(n5749_1), .S0(n5743), .Y(n1527));
MX2X1    g0710(.A(g361), .B(n5749_1), .S0(n5745), .Y(n1532));
NOR4X1   g0711(.A(n5731), .B(n5723), .C(n5718), .D(n5732), .Y(n5753));
NOR3X1   g0712(.A(n5733), .B(n5723), .C(g3229), .Y(n5754_1));
INVX1    g0713(.A(n5733), .Y(n1848));
NOR4X1   g0714(.A(n1863), .B(n1853), .C(g3229), .D(n1848), .Y(n5756));
NOR4X1   g0715(.A(n5754_1), .B(n5753), .C(n5734_1), .D(n5756), .Y(n5757));
MX2X1    g0716(.A(g384), .B(n5757), .S0(n5741), .Y(n1537));
MX2X1    g0717(.A(g373), .B(n5757), .S0(n5743), .Y(n1542));
MX2X1    g0718(.A(g376), .B(n5757), .S0(n5745), .Y(n1547));
NOR2X1   g0719(.A(n5733), .B(g3229), .Y(n5761));
NOR3X1   g0720(.A(n5732), .B(n5731), .C(n5718), .Y(n5762));
NOR4X1   g0721(.A(n5721), .B(n5720), .C(n5719_1), .D(n5722), .Y(n5763));
OAI21X1  g0722(.A0(n5762), .A1(n5761), .B0(n5763), .Y(n5764_1));
MX2X1    g0723(.A(g398), .B(n5764_1), .S0(n5741), .Y(n1552));
MX2X1    g0724(.A(g388), .B(n5764_1), .S0(n5743), .Y(n1557));
MX2X1    g0725(.A(g391), .B(n5764_1), .S0(n5745), .Y(n1562));
NAND2X1  g0726(.A(g408), .B(g276), .Y(n5768));
AOI22X1  g0727(.A0(g411), .A1(g405), .B0(g401), .B1(g414), .Y(n5769_1));
AND2X1   g0728(.A(n5769_1), .B(n5768), .Y(n5770));
INVX1    g0729(.A(n5770), .Y(n5771));
OR4X1    g0730(.A(n5418), .B(n5393), .C(n5387), .D(n5571), .Y(n5772));
NAND2X1  g0731(.A(g417), .B(g276), .Y(n5773));
AOI22X1  g0732(.A0(g420), .A1(g405), .B0(g401), .B1(g423), .Y(n5774_1));
AND2X1   g0733(.A(n5774_1), .B(n5773), .Y(n5775));
AND2X1   g0734(.A(n5775), .B(n5772), .Y(n5776));
NOR3X1   g0735(.A(n5418), .B(n5393), .C(n5387), .Y(n5777));
INVX1    g0736(.A(n5777), .Y(n5778));
OAI21X1  g0737(.A0(n5775), .A1(n5778), .B0(n5770), .Y(n5779_1));
INVX1    g0738(.A(n5775), .Y(n1813));
NOR2X1   g0739(.A(g427), .B(n5545), .Y(n5781));
OAI22X1  g0740(.A0(g428), .A1(n5547), .B0(n5548), .B1(g426), .Y(n5782));
NOR2X1   g0741(.A(n5782), .B(n5781), .Y(n5783));
INVX1    g0742(.A(n5783), .Y(n5784_1));
NOR4X1   g0743(.A(n1813), .B(n5778), .C(n5571), .D(n5784_1), .Y(n5785));
NAND2X1  g0744(.A(n5783), .B(n1813), .Y(n5786));
OAI21X1  g0745(.A0(n5786), .A1(n5777), .B0(n5771), .Y(n5787));
OAI22X1  g0746(.A0(n5785), .A1(n5787), .B0(n5779_1), .B1(n5776), .Y(n5788));
AND2X1   g0747(.A(n5788), .B(g309), .Y(n5789_1));
XOR2X1   g0748(.A(n5789_1), .B(n5771), .Y(n5790));
MX2X1    g0749(.A(g408), .B(n5790), .S0(g276), .Y(n1567));
MX2X1    g0750(.A(g411), .B(n5790), .S0(g405), .Y(n1572));
MX2X1    g0751(.A(g414), .B(n5790), .S0(g401), .Y(n1577));
INVX1    g0752(.A(g309), .Y(n5794_1));
NAND4X1  g0753(.A(n5775), .B(n5777), .C(n5571), .D(n5770), .Y(n5795));
OAI21X1  g0754(.A0(n5784_1), .A1(n5571), .B0(n5777), .Y(n5796));
NAND2X1  g0755(.A(n5796), .B(n5775), .Y(n5797));
OAI21X1  g0756(.A0(n5783), .A1(n5777), .B0(n1813), .Y(n5798));
NAND3X1  g0757(.A(n5798), .B(n5797), .C(n5771), .Y(n5799_1));
AOI21X1  g0758(.A0(n5799_1), .A1(n5795), .B0(n5794_1), .Y(n5800));
XOR2X1   g0759(.A(n5800), .B(n1813), .Y(n5801));
MX2X1    g0760(.A(g417), .B(n5801), .S0(g276), .Y(n1582));
MX2X1    g0761(.A(g420), .B(n5801), .S0(g405), .Y(n1587));
MX2X1    g0762(.A(g423), .B(n5801), .S0(g401), .Y(n1592));
MX2X1    g0763(.A(n5772), .B(n5777), .S0(n1813), .Y(n5805));
OR4X1    g0764(.A(n5784_1), .B(n5770), .C(n5794_1), .D(n5805), .Y(n5806));
NAND3X1  g0765(.A(n5769_1), .B(n5768), .C(g309), .Y(n5807));
OAI21X1  g0766(.A0(n5807), .A1(n5805), .B0(n5806), .Y(n5808));
AND2X1   g0767(.A(n5808), .B(g276), .Y(n5809_1));
MX2X1    g0768(.A(g427), .B(n5806), .S0(n5809_1), .Y(n1597));
AND2X1   g0769(.A(n5808), .B(g405), .Y(n5811));
MX2X1    g0770(.A(g428), .B(n5806), .S0(n5811), .Y(n1602));
AND2X1   g0771(.A(n5808), .B(g401), .Y(n5813));
MX2X1    g0772(.A(g426), .B(n5806), .S0(n5813), .Y(n1607));
NAND2X1  g0773(.A(g429), .B(g276), .Y(n5815));
AOI22X1  g0774(.A0(g432), .A1(g405), .B0(g401), .B1(g435), .Y(n5816));
NAND2X1  g0775(.A(n5816), .B(n5815), .Y(n5817));
OR2X1    g0776(.A(g178), .B(n5382), .Y(n5818_1));
INVX1    g0777(.A(g179), .Y(n5819));
INVX1    g0778(.A(g177), .Y(n5820));
AOI22X1  g0779(.A0(n5819), .A1(g135), .B0(g165), .B1(n5820), .Y(n5821));
AOI21X1  g0780(.A0(n5821), .A1(n5818_1), .B0(n5418), .Y(n5822));
MX2X1    g0781(.A(n5817), .B(n5822), .S0(g309), .Y(n5823_1));
MX2X1    g0782(.A(g429), .B(n5823_1), .S0(g276), .Y(n1612));
MX2X1    g0783(.A(g432), .B(n5823_1), .S0(g405), .Y(n1617));
MX2X1    g0784(.A(g435), .B(n5823_1), .S0(g401), .Y(n1622));
NAND2X1  g0785(.A(g438), .B(g276), .Y(n5827));
AOI22X1  g0786(.A0(g441), .A1(g405), .B0(g401), .B1(g444), .Y(n5828_1));
AND2X1   g0787(.A(n5828_1), .B(n5827), .Y(n5829));
INVX1    g0788(.A(n5829), .Y(n5830));
NOR2X1   g0789(.A(n5829), .B(n5817), .Y(n5831));
INVX1    g0790(.A(n5831), .Y(n5832));
AND2X1   g0791(.A(n5829), .B(n5817), .Y(n5833_1));
INVX1    g0792(.A(n5833_1), .Y(n5834));
MX2X1    g0793(.A(n5832), .B(n5834), .S0(n5822), .Y(n5835));
NOR2X1   g0794(.A(g448), .B(n5545), .Y(n5836));
OAI22X1  g0795(.A0(g449), .A1(n5547), .B0(n5548), .B1(g447), .Y(n5837));
OAI21X1  g0796(.A0(n5837), .A1(n5836), .B0(g309), .Y(n5838_1));
NOR2X1   g0797(.A(n5838_1), .B(n5835), .Y(n5839));
XOR2X1   g0798(.A(n5839), .B(n5830), .Y(n5840));
MX2X1    g0799(.A(g438), .B(n5840), .S0(g276), .Y(n1627));
MX2X1    g0800(.A(g441), .B(n5840), .S0(g405), .Y(n1632));
MX2X1    g0801(.A(g444), .B(n5840), .S0(g401), .Y(n1637));
NOR4X1   g0802(.A(n5836), .B(n5835), .C(n5794_1), .D(n5837), .Y(n5844));
INVX1    g0803(.A(n5844), .Y(n5845));
NOR2X1   g0804(.A(n5830), .B(n5817), .Y(n5846));
AOI22X1  g0805(.A0(n5827), .A1(n5828_1), .B0(n5816), .B1(n5815), .Y(n5847));
MX2X1    g0806(.A(n5847), .B(n5846), .S0(n5822), .Y(n5848_1));
AOI21X1  g0807(.A0(n5848_1), .A1(g309), .B0(n5844), .Y(n5849));
NOR2X1   g0808(.A(n5849), .B(n5545), .Y(n5850));
MX2X1    g0809(.A(g448), .B(n5845), .S0(n5850), .Y(n1642));
NOR2X1   g0810(.A(n5849), .B(n5547), .Y(n5852));
MX2X1    g0811(.A(g449), .B(n5845), .S0(n5852), .Y(n1647));
NOR2X1   g0812(.A(n5849), .B(n5548), .Y(n5854));
MX2X1    g0813(.A(g447), .B(n5845), .S0(n5854), .Y(n1652));
OAI21X1  g0814(.A0(n5577), .A1(n5550), .B0(n5544_1), .Y(n5856));
AOI21X1  g0815(.A0(n5856), .A1(n5557), .B0(n5580), .Y(n5857));
OR2X1    g0816(.A(n5569_1), .B(n5469_1), .Y(n5858_1));
OAI21X1  g0817(.A0(n5857), .A1(n5556), .B0(n5858_1), .Y(n5859));
AOI21X1  g0818(.A0(n5857), .A1(n5556), .B0(n5859), .Y(n5860));
MX2X1    g0819(.A(g312), .B(n5860), .S0(g276), .Y(n1657));
MX2X1    g0820(.A(g313), .B(n5860), .S0(g405), .Y(n1662));
MX2X1    g0821(.A(g314), .B(n5860), .S0(g401), .Y(n1667));
INVX1    g0822(.A(n5428), .Y(n5864));
NAND3X1  g0823(.A(n5539_1), .B(n5502), .C(n5484), .Y(n5865));
NOR2X1   g0824(.A(n5492), .B(n5488), .Y(n5866));
NAND2X1  g0825(.A(n5521), .B(n5866), .Y(n5867));
OR4X1    g0826(.A(n5865), .B(n5529_1), .C(n5525), .D(n5867), .Y(n5868_1));
NAND2X1  g0827(.A(n5868_1), .B(n5864), .Y(n5869));
NOR4X1   g0828(.A(n5560), .B(n5544_1), .C(n5469_1), .D(n5869), .Y(n5870));
NOR2X1   g0829(.A(n5543), .B(n5428), .Y(n5871));
OAI21X1  g0830(.A0(n5868_1), .A1(n5428), .B0(n5572), .Y(n5872));
OR4X1    g0831(.A(n5549_1), .B(n5546), .C(n5871), .D(n5872), .Y(n5873_1));
NAND4X1  g0832(.A(n5468), .B(n5454), .C(n5437_1), .D(n5561), .Y(n5874));
NOR2X1   g0833(.A(n5571), .B(n5550), .Y(n5875));
AOI21X1  g0834(.A0(n5875), .A1(n5874), .B0(n5577), .Y(n5876));
OAI21X1  g0835(.A0(n5873_1), .A1(n5870), .B0(n5876), .Y(n5877_1));
OR2X1    g0836(.A(n5497), .B(n5484), .Y(n5878));
OR2X1    g0837(.A(n5500_1), .B(n5499), .Y(n5879));
OR2X1    g0838(.A(n5488), .B(n5483), .Y(n5880));
NAND3X1  g0839(.A(n5478_1), .B(n5477), .C(n5474), .Y(n5881_1));
OAI21X1  g0840(.A0(n5386), .A1(n5383_1), .B0(n5472), .Y(n5882));
XOR2X1   g0841(.A(n5491_1), .B(n1777), .Y(n5883));
NAND3X1  g0842(.A(n5883), .B(n5882), .C(n5881_1), .Y(n5884));
NAND3X1  g0843(.A(n5884), .B(n5880), .C(n5496_1), .Y(n5885));
NAND3X1  g0844(.A(n5885), .B(n5879), .C(n5878), .Y(n5886_1));
AOI21X1  g0845(.A0(n5886_1), .A1(n5864), .B0(n5579_1), .Y(n5887));
OAI21X1  g0846(.A0(n5869), .A1(n5871), .B0(n5887), .Y(n5888));
AOI21X1  g0847(.A0(n5886_1), .A1(n5864), .B0(n5550), .Y(n5889));
NOR2X1   g0848(.A(n5889), .B(n5553), .Y(n5890));
AOI21X1  g0849(.A0(n5890), .A1(n5888), .B0(n5556), .Y(n5891_1));
AOI22X1  g0850(.A0(n5877_1), .A1(n5891_1), .B0(n5556), .B1(n5574_1), .Y(n5892));
OAI21X1  g0851(.A0(n5892), .A1(n5553), .B0(n5858_1), .Y(n5893));
AOI21X1  g0852(.A0(n5892), .A1(n5553), .B0(n5893), .Y(n5894));
MX2X1    g0853(.A(g315), .B(n5894), .S0(g276), .Y(n1672));
MX2X1    g0854(.A(g316), .B(n5894), .S0(g405), .Y(n1677));
MX2X1    g0855(.A(g317), .B(n5894), .S0(g401), .Y(n1682));
AOI21X1  g0856(.A0(n5872), .A1(n5550), .B0(n5553), .Y(n5899));
OAI21X1  g0857(.A0(n5869), .A1(n5550), .B0(n5899), .Y(n5900));
NOR2X1   g0858(.A(n5506), .B(n5428), .Y(n5901_1));
OR4X1    g0859(.A(n5871), .B(n5901_1), .C(n5794_1), .D(n5579_1), .Y(n5902));
AOI21X1  g0860(.A0(n5902), .A1(n5553), .B0(n5556), .Y(n5903));
AOI22X1  g0861(.A0(n5900), .A1(n5903), .B0(n5556), .B1(n5550), .Y(n5904));
XOR2X1   g0862(.A(n5904), .B(n5579_1), .Y(n5905));
AND2X1   g0863(.A(n5905), .B(n5858_1), .Y(n5906_1));
MX2X1    g0864(.A(g318), .B(n5906_1), .S0(g276), .Y(n1687));
MX2X1    g0865(.A(g319), .B(n5906_1), .S0(g405), .Y(n1692));
MX2X1    g0866(.A(g320), .B(n5906_1), .S0(g401), .Y(n1697));
NOR3X1   g0867(.A(n5579_1), .B(n5544_1), .C(n5469_1), .Y(n5910));
NOR3X1   g0868(.A(n5577), .B(n5550), .C(n5469_1), .Y(n5911_1));
OAI21X1  g0869(.A0(n5911_1), .A1(n5910), .B0(n5557), .Y(n5912));
MX2X1    g0870(.A(n5869), .B(n5794_1), .S0(n5564_1), .Y(n5913));
NOR2X1   g0871(.A(n5913), .B(n5545), .Y(n5914));
MX2X1    g0872(.A(g322), .B(n5912), .S0(n5914), .Y(n1702));
NOR2X1   g0873(.A(n5913), .B(n5547), .Y(n5916_1));
MX2X1    g0874(.A(g323), .B(n5912), .S0(n5916_1), .Y(n1707));
NOR2X1   g0875(.A(n5913), .B(n5548), .Y(n5918));
MX2X1    g0876(.A(g321), .B(n5912), .S0(n5918), .Y(n1712));
NAND4X1  g0877(.A(n5468), .B(n5454), .C(n5437_1), .D(n5569_1), .Y(n5920));
AND2X1   g0878(.A(g309), .B(g276), .Y(n5921_1));
MX2X1    g0879(.A(g403), .B(n5920), .S0(n5921_1), .Y(n1717));
AND2X1   g0880(.A(g309), .B(g405), .Y(n5923));
MX2X1    g0881(.A(g404), .B(n5920), .S0(n5923), .Y(n1722));
AND2X1   g0882(.A(g309), .B(g401), .Y(n5925));
MX2X1    g0883(.A(g402), .B(n5920), .S0(n5925), .Y(n1727));
INVX1    g0884(.A(g305), .Y(n5927));
OAI21X1  g0885(.A0(n5927), .A1(g405), .B0(g299), .Y(n5928));
INVX1    g0886(.A(g298), .Y(n5929));
OR2X1    g0887(.A(n5929), .B(g299), .Y(n5930));
AND2X1   g0888(.A(n5930), .B(n5928), .Y(n1818));
INVX1    g0889(.A(g308), .Y(n5932));
OAI21X1  g0890(.A0(n5932), .A1(g405), .B0(g299), .Y(n5933));
OR2X1    g0891(.A(g300), .B(g299), .Y(n5934));
AND2X1   g0892(.A(n5934), .B(n5933), .Y(n1823));
INVX1    g0893(.A(g297), .Y(n5936_1));
OAI21X1  g0894(.A0(n5936_1), .A1(g405), .B0(g299), .Y(n5937));
OR2X1    g0895(.A(g301), .B(g299), .Y(n5938));
AND2X1   g0896(.A(n5938), .B(n5937), .Y(n1828));
INVX1    g0897(.A(g296), .Y(n5940));
OAI21X1  g0898(.A0(n5940), .A1(g405), .B0(g299), .Y(n5941_1));
OR2X1    g0899(.A(g302), .B(g299), .Y(n5942));
AND2X1   g0900(.A(n5942), .B(n5941_1), .Y(n1833));
INVX1    g0901(.A(g295), .Y(n5944));
OAI21X1  g0902(.A0(n5944), .A1(g405), .B0(g299), .Y(n5945));
OR2X1    g0903(.A(g303), .B(g299), .Y(n5946_1));
AND2X1   g0904(.A(n5946_1), .B(n5945), .Y(n1838));
INVX1    g0905(.A(g294), .Y(n5948));
OAI21X1  g0906(.A0(n5948), .A1(g405), .B0(g299), .Y(n5949));
OR2X1    g0907(.A(g304), .B(g299), .Y(n5950));
AND2X1   g0908(.A(n5950), .B(n5949), .Y(n1843));
INVX1    g0909(.A(n5736), .Y(n1858));
NOR3X1   g0910(.A(n5585), .B(n5557), .C(n5574_1), .Y(n5953));
XOR2X1   g0911(.A(n5495), .B(n5697), .Y(n5954));
XOR2X1   g0912(.A(n5519_1), .B(n5705), .Y(n5955));
XOR2X1   g0913(.A(n5532), .B(n5701), .Y(n5956_1));
NAND3X1  g0914(.A(n5956_1), .B(n5955), .C(n5954), .Y(n5957));
XOR2X1   g0915(.A(n5515), .B(n5714_1), .Y(n5958));
XOR2X1   g0916(.A(n5524_1), .B(n5682), .Y(n5959));
XOR2X1   g0917(.A(n5482_1), .B(n5706), .Y(n5960));
XOR2X1   g0918(.A(n5478_1), .B(n5710), .Y(n5961_1));
NAND4X1  g0919(.A(n5960), .B(n5959), .C(n5958), .D(n5961_1), .Y(n5962));
XOR2X1   g0920(.A(n5528), .B(g79), .Y(n5963));
XOR2X1   g0921(.A(n5491_1), .B(g83), .Y(n5964));
XOR2X1   g0922(.A(n5487_1), .B(g92), .Y(n5965));
OR2X1    g0923(.A(n5965), .B(n5964), .Y(n5966_1));
OR4X1    g0924(.A(n5963), .B(n5739_1), .C(n5399), .D(n5966_1), .Y(n5967));
NOR3X1   g0925(.A(n5967), .B(n5962), .C(n5957), .Y(n5968));
OAI21X1  g0926(.A0(n5968), .A1(n5953), .B0(n1868), .Y(n1873));
INVX1    g0927(.A(g2998), .Y(n5970));
NOR3X1   g0928(.A(g3006), .B(n5970), .C(g2993), .Y(n5971_1));
INVX1    g0929(.A(g3002), .Y(n5972));
INVX1    g0930(.A(g3013), .Y(n5973));
INVX1    g0931(.A(g3024), .Y(n5974));
NOR4X1   g0932(.A(g3010), .B(n5973), .C(n5972), .D(n5974), .Y(n5975));
NAND2X1  g0933(.A(n5975), .B(n5971_1), .Y(n5976_1));
INVX1    g0934(.A(g3018), .Y(n5977));
INVX1    g0935(.A(g3028), .Y(n5978));
NOR4X1   g0936(.A(g3036), .B(n5978), .C(n5977), .D(g3032), .Y(n5979));
INVX1    g0937(.A(n5979), .Y(n5980));
NOR2X1   g0938(.A(n5980), .B(n5976_1), .Y(n5981_1));
INVX1    g0939(.A(n5981_1), .Y(n5982));
MX2X1    g0940(.A(g554), .B(n5982), .S0(g550), .Y(n2012));
INVX1    g0941(.A(g550), .Y(n5984));
INVX1    g0942(.A(g554), .Y(n5985));
MX2X1    g0943(.A(n5985), .B(g557), .S0(n5984), .Y(n2017));
MX2X1    g0944(.A(g510), .B(g557), .S0(g550), .Y(n2022));
NAND2X1  g0945(.A(g569), .B(g545), .Y(n5988));
AOI22X1  g0946(.A0(g571), .A1(g551), .B0(g550), .B1(g573), .Y(n5989));
AND2X1   g0947(.A(n5989), .B(n5988), .Y(n2027));
MX2X1    g0948(.A(g486), .B(n5830), .S0(g474), .Y(n2107));
MX2X1    g0949(.A(g487), .B(n5830), .S0(g481), .Y(n2112));
MX2X1    g0950(.A(g488), .B(n5830), .S0(g485), .Y(n2117));
MX2X1    g0951(.A(g455), .B(n5739_1), .S0(g474), .Y(n2122));
MX2X1    g0952(.A(g458), .B(n5739_1), .S0(g481), .Y(n2127));
MX2X1    g0953(.A(g461), .B(n5739_1), .S0(g485), .Y(n2132));
MX2X1    g0954(.A(g477), .B(n5564_1), .S0(g474), .Y(n2137));
MX2X1    g0955(.A(g478), .B(n5564_1), .S0(g481), .Y(n2142));
MX2X1    g0956(.A(g479), .B(n5564_1), .S0(g485), .Y(n2147));
MX2X1    g0957(.A(g480), .B(n5775), .S0(g474), .Y(n2152));
MX2X1    g0958(.A(g484), .B(n5775), .S0(g481), .Y(n2157));
MX2X1    g0959(.A(g464), .B(n5775), .S0(g485), .Y(n2162));
MX2X1    g0960(.A(g465), .B(n5575), .S0(g474), .Y(n2167));
MX2X1    g0961(.A(g468), .B(n5575), .S0(g481), .Y(n2172));
MX2X1    g0962(.A(g471), .B(n5575), .S0(g485), .Y(n2177));
NAND2X1  g0963(.A(g565), .B(g545), .Y(n6006_1));
AOI22X1  g0964(.A0(g567), .A1(g551), .B0(g550), .B1(g489), .Y(n6007));
AND2X1   g0965(.A(n6007), .B(n6006_1), .Y(n2182));
INVX1    g0966(.A(g551), .Y(n6009));
NOR2X1   g0967(.A(g477), .B(n6009), .Y(n6010));
OAI22X1  g0968(.A0(g478), .A1(n5984), .B0(n5297), .B1(g479), .Y(n6011_1));
NOR2X1   g0969(.A(n6011_1), .B(n6010), .Y(n2195));
NOR2X1   g0970(.A(g480), .B(n6009), .Y(n6013));
OAI22X1  g0971(.A0(g484), .A1(n5984), .B0(n5297), .B1(g464), .Y(n6014));
NOR2X1   g0972(.A(n6014), .B(n6013), .Y(n2209));
NOR2X1   g0973(.A(g486), .B(n6009), .Y(n6016_1));
OAI22X1  g0974(.A0(g487), .A1(n5984), .B0(n5297), .B1(g488), .Y(n6017));
NOR2X1   g0975(.A(n6017), .B(n6016_1), .Y(n2218));
NOR2X1   g0976(.A(g582), .B(n5297), .Y(n6019));
OAI22X1  g0977(.A0(g583), .A1(n6009), .B0(n5984), .B1(g581), .Y(n6020));
NOR2X1   g0978(.A(g579), .B(n5297), .Y(n6021_1));
OAI22X1  g0979(.A0(g580), .A1(n6009), .B0(n5984), .B1(g578), .Y(n6022));
NOR2X1   g0980(.A(n6022), .B(n6021_1), .Y(n6023));
OR4X1    g0981(.A(n6020), .B(n6019), .C(g3229), .D(n6023), .Y(n6024));
NOR2X1   g0982(.A(g585), .B(n5297), .Y(n6025));
OAI22X1  g0983(.A0(g586), .A1(n6009), .B0(n5984), .B1(g584), .Y(n6026_1));
NOR2X1   g0984(.A(n6026_1), .B(n6025), .Y(n6027));
OAI21X1  g0985(.A0(n6027), .A1(n5718), .B0(n6024), .Y(n6028));
INVX1    g0986(.A(n6023), .Y(n2382));
INVX1    g0987(.A(n6027), .Y(n2372));
NOR2X1   g0988(.A(g576), .B(n5297), .Y(n6031_1));
OAI22X1  g0989(.A0(g577), .A1(n6009), .B0(n5984), .B1(g575), .Y(n6032));
NOR2X1   g0990(.A(n6032), .B(n6031_1), .Y(n6033));
NOR4X1   g0991(.A(n2372), .B(n2382), .C(n5718), .D(n6033), .Y(n6034));
NOR4X1   g0992(.A(n6026_1), .B(n6025), .C(g3229), .D(n6033), .Y(n6035));
NOR2X1   g0993(.A(n6020), .B(n6019), .Y(n6036_1));
NOR3X1   g0994(.A(n6033), .B(n6036_1), .C(n5718), .Y(n6037));
NOR4X1   g0995(.A(n6035), .B(n6034), .C(n6028), .D(n6037), .Y(n6038));
NAND2X1  g0996(.A(g490), .B(g545), .Y(n6039));
AOI22X1  g0997(.A0(g493), .A1(g551), .B0(g550), .B1(g496), .Y(n6040));
AND2X1   g0998(.A(n6040), .B(n6039), .Y(n6041_1));
INVX1    g0999(.A(n6041_1), .Y(n6042));
NAND2X1  g1000(.A(g614), .B(g545), .Y(n6043));
AOI22X1  g1001(.A0(g617), .A1(g551), .B0(g550), .B1(g620), .Y(n6044));
AND2X1   g1002(.A(n6044), .B(n6043), .Y(n6045));
INVX1    g1003(.A(n6045), .Y(n6046_1));
NAND3X1  g1004(.A(n6041_1), .B(n6046_1), .C(g510), .Y(n6047));
OR2X1    g1005(.A(g3010), .B(g3002), .Y(n6048));
NOR4X1   g1006(.A(g3024), .B(g3013), .C(g3006), .D(n6048), .Y(n6049));
NAND2X1  g1007(.A(g605), .B(g545), .Y(n6050));
AOI22X1  g1008(.A0(g608), .A1(g551), .B0(g550), .B1(g611), .Y(n6051_1));
AND2X1   g1009(.A(n6051_1), .B(n6050), .Y(n6052));
INVX1    g1010(.A(n6052), .Y(n6053));
AOI22X1  g1011(.A0(n6049), .A1(n6047), .B0(n6042), .B1(n6053), .Y(n2367));
NAND2X1  g1012(.A(n2367), .B(g545), .Y(n6055));
MX2X1    g1013(.A(n6038), .B(g576), .S0(n6055), .Y(n2227));
NAND2X1  g1014(.A(n2367), .B(g551), .Y(n6057));
MX2X1    g1015(.A(n6038), .B(g577), .S0(n6057), .Y(n2232));
NAND2X1  g1016(.A(n2367), .B(g550), .Y(n6059));
MX2X1    g1017(.A(n6038), .B(g575), .S0(n6059), .Y(n2237));
NOR4X1   g1018(.A(n6031_1), .B(n6036_1), .C(g3229), .D(n6032), .Y(n6061_1));
NOR3X1   g1019(.A(n6023), .B(n6020), .C(n6019), .Y(n6062));
NOR3X1   g1020(.A(n6062), .B(n6061_1), .C(n6037), .Y(n6063));
MX2X1    g1021(.A(n6063), .B(g579), .S0(n6055), .Y(n2242));
MX2X1    g1022(.A(n6063), .B(g580), .S0(n6057), .Y(n2247));
MX2X1    g1023(.A(n6063), .B(g578), .S0(n6059), .Y(n2252));
NOR4X1   g1024(.A(n6031_1), .B(n6023), .C(n5718), .D(n6032), .Y(n6067));
NOR3X1   g1025(.A(n6033), .B(n6023), .C(g3229), .Y(n6068));
INVX1    g1026(.A(n6033), .Y(n2387));
NOR4X1   g1027(.A(n2372), .B(n2382), .C(g3229), .D(n2387), .Y(n6070));
NOR4X1   g1028(.A(n6068), .B(n6067), .C(n6034), .D(n6070), .Y(n6071_1));
MX2X1    g1029(.A(n6071_1), .B(g582), .S0(n6055), .Y(n2257));
MX2X1    g1030(.A(n6071_1), .B(g583), .S0(n6057), .Y(n2262));
MX2X1    g1031(.A(n6071_1), .B(g581), .S0(n6059), .Y(n2267));
NOR2X1   g1032(.A(n6033), .B(g3229), .Y(n6075));
NOR3X1   g1033(.A(n6032), .B(n6031_1), .C(n5718), .Y(n6076_1));
NOR4X1   g1034(.A(n6021_1), .B(n6020), .C(n6019), .D(n6022), .Y(n6077));
OAI21X1  g1035(.A0(n6076_1), .A1(n6075), .B0(n6077), .Y(n6078));
MX2X1    g1036(.A(n6078), .B(g585), .S0(n6055), .Y(n2272));
MX2X1    g1037(.A(n6078), .B(g586), .S0(n6057), .Y(n2277));
MX2X1    g1038(.A(n6078), .B(g584), .S0(n6059), .Y(n2282));
INVX1    g1039(.A(n2027), .Y(n6082));
AND2X1   g1040(.A(g524), .B(g185), .Y(n6083));
NAND2X1  g1041(.A(g587), .B(g545), .Y(n6084));
AOI22X1  g1042(.A0(g590), .A1(g551), .B0(g550), .B1(g593), .Y(n6085));
NAND2X1  g1043(.A(n6085), .B(n6084), .Y(n6086_1));
AOI21X1  g1044(.A0(n6083), .A1(n6082), .B0(n6086_1), .Y(n6087));
NOR2X1   g1045(.A(n6087), .B(n5981_1), .Y(n6088));
MX2X1    g1046(.A(g587), .B(n6088), .S0(g545), .Y(n2287));
MX2X1    g1047(.A(g590), .B(n6088), .S0(g551), .Y(n2292));
MX2X1    g1048(.A(g593), .B(n6088), .S0(g550), .Y(n2297));
INVX1    g1049(.A(n2182), .Y(n6092));
AND2X1   g1050(.A(g542), .B(g185), .Y(n6093));
NAND2X1  g1051(.A(g596), .B(g545), .Y(n6094));
AOI22X1  g1052(.A0(g599), .A1(g551), .B0(g550), .B1(g602), .Y(n6095));
NAND2X1  g1053(.A(n6095), .B(n6094), .Y(n6096_1));
AOI21X1  g1054(.A0(n6093), .A1(n6092), .B0(n6096_1), .Y(n6097));
NOR2X1   g1055(.A(n6097), .B(n5981_1), .Y(n6098));
MX2X1    g1056(.A(g596), .B(n6098), .S0(g545), .Y(n2302));
MX2X1    g1057(.A(g599), .B(n6098), .S0(g551), .Y(n2307));
MX2X1    g1058(.A(g602), .B(n6098), .S0(g550), .Y(n2312));
OR4X1    g1059(.A(n6031_1), .B(n6022), .C(n6021_1), .D(n6032), .Y(n6102));
NAND2X1  g1060(.A(g325), .B(g349), .Y(n6103));
AOI22X1  g1061(.A0(g331), .A1(g351), .B0(g353), .B1(g337), .Y(n6104));
AND2X1   g1062(.A(n6104), .B(n6103), .Y(n6105));
INVX1    g1063(.A(n6105), .Y(n6106_1));
NAND2X1  g1064(.A(g325), .B(g364), .Y(n6107));
AOI22X1  g1065(.A0(g331), .A1(g366), .B0(g368), .B1(g337), .Y(n6108));
AND2X1   g1066(.A(n6108), .B(n6107), .Y(n6109));
NAND2X1  g1067(.A(g325), .B(g379), .Y(n6110));
AOI22X1  g1068(.A0(g331), .A1(g381), .B0(g383), .B1(g337), .Y(n6111_1));
AND2X1   g1069(.A(n6111_1), .B(n6110), .Y(n6112));
OR4X1    g1070(.A(n6109), .B(n6106_1), .C(n6102), .D(n6112), .Y(n6113));
INVX1    g1071(.A(n6036_1), .Y(n2377));
INVX1    g1072(.A(n6109), .Y(n6115));
NAND2X1  g1073(.A(g325), .B(g394), .Y(n6116_1));
NAND2X1  g1074(.A(g337), .B(g324), .Y(n6117));
NAND2X1  g1075(.A(g331), .B(g396), .Y(n6118));
NAND3X1  g1076(.A(n6118), .B(n6117), .C(n6116_1), .Y(n6119));
NAND2X1  g1077(.A(n6119), .B(n6115), .Y(n6120));
OR4X1    g1078(.A(n6105), .B(n6023), .C(n2377), .D(n6120), .Y(n6121_1));
AND2X1   g1079(.A(n6112), .B(n6105), .Y(n6122));
NAND3X1  g1080(.A(n6122), .B(n6115), .C(n6077), .Y(n6123));
INVX1    g1081(.A(n6112), .Y(n6124));
NOR4X1   g1082(.A(n6032), .B(n6031_1), .C(n6036_1), .D(n6105), .Y(n6125));
NAND3X1  g1083(.A(n6125), .B(n6124), .C(n6115), .Y(n6126_1));
NAND4X1  g1084(.A(n6123), .B(n6121_1), .C(n6113), .D(n6126_1), .Y(n6127));
OR4X1    g1085(.A(n6105), .B(n2387), .C(n2372), .D(n6119), .Y(n6128));
AND2X1   g1086(.A(n6109), .B(n6105), .Y(n6129));
NAND3X1  g1087(.A(n6129), .B(n2387), .C(n6023), .Y(n6130));
NAND4X1  g1088(.A(n6105), .B(n2387), .C(n2372), .D(n6119), .Y(n6131_1));
OR4X1    g1089(.A(n6115), .B(n6033), .C(n6036_1), .D(n6112), .Y(n6132));
NAND4X1  g1090(.A(n6131_1), .B(n6130), .C(n6128), .D(n6132), .Y(n6133));
OR4X1    g1091(.A(n6105), .B(n6033), .C(n6036_1), .D(n6115), .Y(n6134));
OAI21X1  g1092(.A0(n6026_1), .A1(n6025), .B0(n6122), .Y(n6135));
OR4X1    g1093(.A(n6109), .B(n6105), .C(n6023), .D(n6124), .Y(n6136_1));
OR4X1    g1094(.A(n6032), .B(n6031_1), .C(n6036_1), .D(n6119), .Y(n6137));
NAND4X1  g1095(.A(n6136_1), .B(n6135), .C(n6134), .D(n6137), .Y(n6138));
OR4X1    g1096(.A(n6023), .B(n6020), .C(n6019), .D(n6105), .Y(n6139));
OR2X1    g1097(.A(n6115), .B(n6105), .Y(n6140));
OR4X1    g1098(.A(n6033), .B(n6026_1), .C(n6025), .D(n6112), .Y(n6141_1));
OAI22X1  g1099(.A0(n6140), .A1(n6141_1), .B0(n6139), .B1(n6124), .Y(n6142));
NOR4X1   g1100(.A(n6138), .B(n6133), .C(n6127), .D(n6142), .Y(n6143));
NAND4X1  g1101(.A(n6115), .B(n6105), .C(n6027), .D(n6124), .Y(n6144));
NOR3X1   g1102(.A(n6144), .B(n6033), .C(n2382), .Y(n6145));
NAND4X1  g1103(.A(n6115), .B(n6106_1), .C(n6036_1), .D(n6119), .Y(n6146_1));
NOR2X1   g1104(.A(n6146_1), .B(n6102), .Y(n6147));
NOR4X1   g1105(.A(n6105), .B(n6102), .C(n2372), .D(n6124), .Y(n6148));
NOR4X1   g1106(.A(n6106_1), .B(n6033), .C(n6036_1), .D(n6120), .Y(n6149));
OR4X1    g1107(.A(n6148), .B(n6147), .C(n6145), .D(n6149), .Y(n6150));
NAND4X1  g1108(.A(n6109), .B(n6033), .C(n2382), .D(n6124), .Y(n6151_1));
OR4X1    g1109(.A(n6109), .B(n6105), .C(n6027), .D(n6112), .Y(n6152));
OR4X1    g1110(.A(n6106_1), .B(n6033), .C(n6023), .D(n6124), .Y(n6153));
NAND3X1  g1111(.A(n6153), .B(n6152), .C(n6151_1), .Y(n6154));
NAND2X1  g1112(.A(n6125), .B(n6109), .Y(n6155));
NAND2X1  g1113(.A(n6129), .B(n6062), .Y(n6156_1));
OR4X1    g1114(.A(n6033), .B(n2382), .C(n2377), .D(n6119), .Y(n6157));
NAND3X1  g1115(.A(n6157), .B(n6156_1), .C(n6155), .Y(n6158));
NOR3X1   g1116(.A(n6158), .B(n6154), .C(n6150), .Y(n6159));
NAND2X1  g1117(.A(n6159), .B(n6097), .Y(n6160_1));
OR2X1    g1118(.A(n6160_1), .B(n6143), .Y(n6161));
INVX1    g1119(.A(n6087), .Y(n6162));
NOR2X1   g1120(.A(n6097), .B(n6162), .Y(n6163));
AOI21X1  g1121(.A0(n6163), .A1(n6159), .B0(n5982), .Y(n6164_1));
AOI22X1  g1122(.A0(n6161), .A1(n6164_1), .B0(n6045), .B1(n5982), .Y(n6165));
MX2X1    g1123(.A(g614), .B(n6165), .S0(g545), .Y(n2317));
MX2X1    g1124(.A(g617), .B(n6165), .S0(g551), .Y(n2322));
MX2X1    g1125(.A(g620), .B(n6165), .S0(g550), .Y(n2327));
NAND3X1  g1126(.A(n6143), .B(n6097), .C(n6162), .Y(n6169_1));
NOR2X1   g1127(.A(n6159), .B(n6162), .Y(n6170));
AOI21X1  g1128(.A0(n6170), .A1(n6143), .B0(n5982), .Y(n6171));
AOI22X1  g1129(.A0(n6169_1), .A1(n6171), .B0(n6052), .B1(n5982), .Y(n6172));
MX2X1    g1130(.A(g605), .B(n6172), .S0(g545), .Y(n2332));
MX2X1    g1131(.A(g608), .B(n6172), .S0(g551), .Y(n2337));
MX2X1    g1132(.A(g611), .B(n6172), .S0(g550), .Y(n2342));
INVX1    g1133(.A(g510), .Y(n6176));
NOR3X1   g1134(.A(n6042), .B(n6046_1), .C(n6176), .Y(n6177));
MX2X1    g1135(.A(g490), .B(n6177), .S0(g545), .Y(n2347));
MX2X1    g1136(.A(g493), .B(n6177), .S0(g551), .Y(n2352));
MX2X1    g1137(.A(g496), .B(n6177), .S0(g550), .Y(n2357));
INVX1    g1138(.A(g506), .Y(n6181));
INVX1    g1139(.A(g516), .Y(n6182));
OAI21X1  g1140(.A0(n6182), .A1(g551), .B0(n6181), .Y(n6183));
OR2X1    g1141(.A(g515), .B(n6181), .Y(n6184_1));
AND2X1   g1142(.A(n6184_1), .B(n6183), .Y(n2392));
INVX1    g1143(.A(g517), .Y(n6186));
OAI21X1  g1144(.A0(n6186), .A1(g551), .B0(n6181), .Y(n6187));
OR2X1    g1145(.A(g514), .B(n6181), .Y(n6188));
AND2X1   g1146(.A(n6188), .B(n6187), .Y(n2397));
INVX1    g1147(.A(g518), .Y(n6190));
OAI21X1  g1148(.A0(n6190), .A1(g551), .B0(n6181), .Y(n6191));
OR2X1    g1149(.A(g509), .B(n6181), .Y(n6192));
AND2X1   g1150(.A(n6192), .B(n6191), .Y(n2402));
INVX1    g1151(.A(g519), .Y(n6194_1));
OAI21X1  g1152(.A0(n6194_1), .A1(g551), .B0(n6181), .Y(n6195));
OR2X1    g1153(.A(g508), .B(n6181), .Y(n6196));
AND2X1   g1154(.A(n6196), .B(n6195), .Y(n2407));
INVX1    g1155(.A(g507), .Y(n6198));
NOR3X1   g1156(.A(g520), .B(g506), .C(g551), .Y(n6199_1));
AOI21X1  g1157(.A0(n6198), .A1(g506), .B0(n6199_1), .Y(n2412));
INVX1    g1158(.A(g451), .Y(n2421));
INVX1    g1159(.A(g453), .Y(n2426));
INVX1    g1160(.A(g279), .Y(n2431));
INVX1    g1161(.A(g281), .Y(n2436));
INVX1    g1162(.A(g283), .Y(n2441));
INVX1    g1163(.A(g285), .Y(n2446));
INVX1    g1164(.A(g287), .Y(n2451));
INVX1    g1165(.A(g289), .Y(n2456));
INVX1    g1166(.A(g291), .Y(n2466));
MX2X1    g1167(.A(n2466), .B(g305), .S0(n5718), .Y(n2461));
MX2X1    g1168(.A(g630), .B(g510), .S0(g629), .Y(n2484));
MX2X1    g1169(.A(g659), .B(n6049), .S0(g629), .Y(n2489));
INVX1    g1170(.A(g659), .Y(n6213));
INVX1    g1171(.A(g640), .Y(n6214_1));
NAND3X1  g1172(.A(n6214_1), .B(n6213), .C(g629), .Y(n6215));
INVX1    g1173(.A(g629), .Y(n6216));
OAI21X1  g1174(.A0(g659), .A1(n6216), .B0(g640), .Y(n6217));
AND2X1   g1175(.A(g630), .B(g626), .Y(n6218));
AOI21X1  g1176(.A0(n6217), .A1(n6215), .B0(n6218), .Y(n2494));
INVX1    g1177(.A(g633), .Y(n6220));
NOR3X1   g1178(.A(n6214_1), .B(g659), .C(n6216), .Y(n6221));
XOR2X1   g1179(.A(n6221), .B(n6220), .Y(n6222));
NOR2X1   g1180(.A(n6222), .B(n6218), .Y(n2499));
INVX1    g1181(.A(g653), .Y(n6224_1));
NOR4X1   g1182(.A(n6214_1), .B(g659), .C(n6216), .D(n6220), .Y(n6225));
XOR2X1   g1183(.A(n6225), .B(n6224_1), .Y(n6226));
NOR2X1   g1184(.A(n6226), .B(n6218), .Y(n2504));
INVX1    g1185(.A(g646), .Y(n6228));
AND2X1   g1186(.A(n6225), .B(g653), .Y(n6229_1));
XOR2X1   g1187(.A(n6229_1), .B(n6228), .Y(n6230));
NOR2X1   g1188(.A(n6230), .B(n6218), .Y(n2509));
NAND3X1  g1189(.A(n6225), .B(g646), .C(g653), .Y(n6232));
XOR2X1   g1190(.A(n6232), .B(g660), .Y(n6233));
NOR2X1   g1191(.A(n6233), .B(n6218), .Y(n2514));
INVX1    g1192(.A(g660), .Y(n6235));
OAI21X1  g1193(.A0(n6232), .A1(n6235), .B0(g672), .Y(n6236));
INVX1    g1194(.A(g672), .Y(n6237));
NAND4X1  g1195(.A(n6237), .B(g660), .C(g646), .D(n6229_1), .Y(n6238));
AOI21X1  g1196(.A0(n6238), .A1(n6236), .B0(n6218), .Y(n2519));
INVX1    g1197(.A(g666), .Y(n6240));
NOR3X1   g1198(.A(n6232), .B(n6237), .C(n6235), .Y(n6241));
XOR2X1   g1199(.A(n6241), .B(n6240), .Y(n6242));
NOR2X1   g1200(.A(n6242), .B(n6218), .Y(n2524));
INVX1    g1201(.A(g679), .Y(n6244_1));
NOR4X1   g1202(.A(n6240), .B(n6237), .C(n6235), .D(n6232), .Y(n6245));
XOR2X1   g1203(.A(n6245), .B(n6244_1), .Y(n6246));
NOR2X1   g1204(.A(n6246), .B(n6218), .Y(n2529));
INVX1    g1205(.A(g686), .Y(n6248));
AND2X1   g1206(.A(n6245), .B(g679), .Y(n6249_1));
XOR2X1   g1207(.A(n6249_1), .B(n6248), .Y(n6250));
NOR2X1   g1208(.A(n6250), .B(n6218), .Y(n2534));
NAND3X1  g1209(.A(n6245), .B(g686), .C(g679), .Y(n6252));
XOR2X1   g1210(.A(n6252), .B(g692), .Y(n6253));
NOR2X1   g1211(.A(n6253), .B(n6218), .Y(n2539));
NAND4X1  g1212(.A(g623), .B(g538), .C(g525), .D(n6213), .Y(n6255));
MX2X1    g1213(.A(n6214_1), .B(g699), .S0(n6255), .Y(n2544));
NAND4X1  g1214(.A(g626), .B(g538), .C(g525), .D(n6213), .Y(n6257));
MX2X1    g1215(.A(n6214_1), .B(g700), .S0(n6257), .Y(n2549));
NAND4X1  g1216(.A(g629), .B(g538), .C(g525), .D(n6213), .Y(n6259_1));
MX2X1    g1217(.A(n6214_1), .B(g698), .S0(n6259_1), .Y(n2554));
MX2X1    g1218(.A(n6220), .B(g702), .S0(n6255), .Y(n2559));
MX2X1    g1219(.A(n6220), .B(g703), .S0(n6257), .Y(n2564));
MX2X1    g1220(.A(n6220), .B(g701), .S0(n6259_1), .Y(n2569));
MX2X1    g1221(.A(n6224_1), .B(g705), .S0(n6255), .Y(n2574));
MX2X1    g1222(.A(n6224_1), .B(g706), .S0(n6257), .Y(n2579));
MX2X1    g1223(.A(n6224_1), .B(g704), .S0(n6259_1), .Y(n2584));
MX2X1    g1224(.A(n6228), .B(g708), .S0(n6255), .Y(n2589));
MX2X1    g1225(.A(n6228), .B(g709), .S0(n6257), .Y(n2594));
MX2X1    g1226(.A(n6228), .B(g707), .S0(n6259_1), .Y(n2599));
MX2X1    g1227(.A(n6235), .B(g711), .S0(n6255), .Y(n2604));
MX2X1    g1228(.A(n6235), .B(g712), .S0(n6257), .Y(n2609));
MX2X1    g1229(.A(n6235), .B(g710), .S0(n6259_1), .Y(n2614));
MX2X1    g1230(.A(n6237), .B(g714), .S0(n6255), .Y(n2619));
MX2X1    g1231(.A(n6237), .B(g715), .S0(n6257), .Y(n2624));
MX2X1    g1232(.A(n6237), .B(g713), .S0(n6259_1), .Y(n2629));
MX2X1    g1233(.A(n6240), .B(g717), .S0(n6255), .Y(n2634));
MX2X1    g1234(.A(n6240), .B(g718), .S0(n6257), .Y(n2639));
MX2X1    g1235(.A(n6240), .B(g716), .S0(n6259_1), .Y(n2644));
MX2X1    g1236(.A(n6244_1), .B(g720), .S0(n6255), .Y(n2649));
MX2X1    g1237(.A(n6244_1), .B(g721), .S0(n6257), .Y(n2654));
MX2X1    g1238(.A(n6244_1), .B(g719), .S0(n6259_1), .Y(n2659));
MX2X1    g1239(.A(n6248), .B(g723), .S0(n6255), .Y(n2664));
MX2X1    g1240(.A(n6248), .B(g724), .S0(n6257), .Y(n2669));
MX2X1    g1241(.A(n6248), .B(g722), .S0(n6259_1), .Y(n2674));
INVX1    g1242(.A(g692), .Y(n6285));
MX2X1    g1243(.A(n6285), .B(g726), .S0(n6255), .Y(n2679));
MX2X1    g1244(.A(n6285), .B(g727), .S0(n6257), .Y(n2684));
MX2X1    g1245(.A(n6285), .B(g725), .S0(n6259_1), .Y(n2689));
AND2X1   g1246(.A(g630), .B(g623), .Y(n6289_1));
MX2X1    g1247(.A(g729), .B(n6045), .S0(n6289_1), .Y(n2694));
MX2X1    g1248(.A(g730), .B(n6045), .S0(n6218), .Y(n2699));
AND2X1   g1249(.A(g630), .B(g629), .Y(n6292));
MX2X1    g1250(.A(g728), .B(n6045), .S0(n6292), .Y(n2704));
MX2X1    g1251(.A(g732), .B(n6052), .S0(n6289_1), .Y(n2709));
MX2X1    g1252(.A(g733), .B(n6052), .S0(n6218), .Y(n2714));
MX2X1    g1253(.A(g731), .B(n6052), .S0(n6292), .Y(n2719));
INVX1    g1254(.A(g623), .Y(n6297));
NOR2X1   g1255(.A(g717), .B(n6297), .Y(n6298));
INVX1    g1256(.A(g626), .Y(n6299_1));
OAI22X1  g1257(.A0(g718), .A1(n6299_1), .B0(n6216), .B1(g716), .Y(n6300));
OR2X1    g1258(.A(n6300), .B(n6298), .Y(n6301));
XOR2X1   g1259(.A(n6301), .B(g666), .Y(n6302));
NOR2X1   g1260(.A(g723), .B(n6297), .Y(n6303));
OAI22X1  g1261(.A0(g724), .A1(n6299_1), .B0(n6216), .B1(g722), .Y(n6304_1));
NOR2X1   g1262(.A(n6304_1), .B(n6303), .Y(n6305));
XOR2X1   g1263(.A(n6305), .B(n6248), .Y(n6306));
NOR2X1   g1264(.A(g720), .B(n6297), .Y(n6307));
OAI22X1  g1265(.A0(g721), .A1(n6299_1), .B0(n6216), .B1(g719), .Y(n6308));
NOR2X1   g1266(.A(n6308), .B(n6307), .Y(n6309_1));
XOR2X1   g1267(.A(n6309_1), .B(n6244_1), .Y(n6310));
NOR2X1   g1268(.A(g714), .B(n6297), .Y(n6311));
OAI22X1  g1269(.A0(g715), .A1(n6299_1), .B0(n6216), .B1(g713), .Y(n6312));
NOR2X1   g1270(.A(n6312), .B(n6311), .Y(n6313));
XOR2X1   g1271(.A(n6313), .B(n6237), .Y(n6314_1));
OR4X1    g1272(.A(n6310), .B(n6306), .C(n6302), .D(n6314_1), .Y(n6315));
INVX1    g1273(.A(g709), .Y(n6316));
INVX1    g1274(.A(g707), .Y(n6317));
AOI22X1  g1275(.A0(n6316), .A1(g626), .B0(g629), .B1(n6317), .Y(n6318));
OAI21X1  g1276(.A0(g708), .A1(n6297), .B0(n6318), .Y(n6319_1));
XOR2X1   g1277(.A(n6319_1), .B(n6228), .Y(n6320));
NOR2X1   g1278(.A(g711), .B(n6297), .Y(n6321));
OAI22X1  g1279(.A0(g712), .A1(n6299_1), .B0(n6216), .B1(g710), .Y(n6322));
NOR2X1   g1280(.A(n6322), .B(n6321), .Y(n6323));
XOR2X1   g1281(.A(n6323), .B(g660), .Y(n6324_1));
NAND2X1  g1282(.A(n6324_1), .B(n6320), .Y(n6325));
NOR2X1   g1283(.A(g699), .B(n6297), .Y(n6326));
OAI22X1  g1284(.A0(g700), .A1(n6299_1), .B0(n6216), .B1(g698), .Y(n6327));
NOR2X1   g1285(.A(n6327), .B(n6326), .Y(n6328));
XOR2X1   g1286(.A(n6328), .B(g640), .Y(n6329_1));
INVX1    g1287(.A(g703), .Y(n6330));
INVX1    g1288(.A(g701), .Y(n6331));
AOI22X1  g1289(.A0(n6330), .A1(g626), .B0(g629), .B1(n6331), .Y(n6332));
OAI21X1  g1290(.A0(g702), .A1(n6297), .B0(n6332), .Y(n6333));
XOR2X1   g1291(.A(n6333), .B(n6220), .Y(n6334_1));
NAND2X1  g1292(.A(n6334_1), .B(n6329_1), .Y(n6335));
NOR2X1   g1293(.A(g726), .B(n6297), .Y(n6336));
OAI22X1  g1294(.A0(g727), .A1(n6299_1), .B0(n6216), .B1(g725), .Y(n6337));
NOR2X1   g1295(.A(n6337), .B(n6336), .Y(n6338));
XOR2X1   g1296(.A(n6338), .B(n6285), .Y(n6339_1));
NOR2X1   g1297(.A(g705), .B(n6297), .Y(n6340));
OAI22X1  g1298(.A0(g706), .A1(n6299_1), .B0(n6216), .B1(g704), .Y(n6341));
NOR2X1   g1299(.A(n6341), .B(n6340), .Y(n6342));
XOR2X1   g1300(.A(n6342), .B(n6224_1), .Y(n6343));
OR2X1    g1301(.A(n6343), .B(n6339_1), .Y(n6344_1));
NOR4X1   g1302(.A(n6335), .B(n6325), .C(n6315), .D(n6344_1), .Y(n6345));
INVX1    g1303(.A(g733), .Y(n6346));
INVX1    g1304(.A(g731), .Y(n6347));
AOI22X1  g1305(.A0(n6346), .A1(g626), .B0(g629), .B1(n6347), .Y(n6348));
OAI21X1  g1306(.A0(g732), .A1(n6297), .B0(n6348), .Y(n6349_1));
NOR2X1   g1307(.A(g729), .B(n6297), .Y(n6350));
OAI22X1  g1308(.A0(g730), .A1(n6299_1), .B0(n6216), .B1(g728), .Y(n6351));
NOR4X1   g1309(.A(n6350), .B(n6349_1), .C(n6345), .D(n6351), .Y(n6352));
MX2X1    g1310(.A(n6352), .B(g735), .S0(n6255), .Y(n2724));
MX2X1    g1311(.A(n6352), .B(g736), .S0(n6257), .Y(n2729));
MX2X1    g1312(.A(n6352), .B(g734), .S0(n6259_1), .Y(n2734));
INVX1    g1313(.A(g630), .Y(n6356));
INVX1    g1314(.A(g525), .Y(n6357));
INVX1    g1315(.A(g538), .Y(n6358));
NOR3X1   g1316(.A(g659), .B(n6358), .C(n6357), .Y(n6359_1));
OAI21X1  g1317(.A0(n6359_1), .A1(g630), .B0(g623), .Y(n6360));
MX2X1    g1318(.A(n6356), .B(g738), .S0(n6360), .Y(n2739));
OAI21X1  g1319(.A0(n6359_1), .A1(g630), .B0(g626), .Y(n6362));
MX2X1    g1320(.A(n6356), .B(g739), .S0(n6362), .Y(n2744));
OAI21X1  g1321(.A0(n6359_1), .A1(g630), .B0(g629), .Y(n6364_1));
MX2X1    g1322(.A(n6356), .B(g737), .S0(n6364_1), .Y(n2749));
INVX1    g1323(.A(g785), .Y(n3496));
NAND2X1  g1324(.A(g869), .B(g826), .Y(n6367));
MX2X1    g1325(.A(n3496), .B(g818), .S0(n6367), .Y(n2767));
NAND2X1  g1326(.A(g869), .B(g823), .Y(n6369_1));
MX2X1    g1327(.A(n3496), .B(g819), .S0(n6369_1), .Y(n2772));
AND2X1   g1328(.A(g869), .B(g853), .Y(n6371));
MX2X1    g1329(.A(g817), .B(n3496), .S0(n6371), .Y(n2777));
INVX1    g1330(.A(g789), .Y(n3487));
MX2X1    g1331(.A(n3487), .B(g821), .S0(n6367), .Y(n2782));
MX2X1    g1332(.A(n3487), .B(g822), .S0(n6369_1), .Y(n2787));
MX2X1    g1333(.A(g820), .B(n3487), .S0(n6371), .Y(n2792));
INVX1    g1334(.A(g793), .Y(n3478));
MX2X1    g1335(.A(n3478), .B(g830), .S0(n6367), .Y(n2797));
MX2X1    g1336(.A(n3478), .B(g831), .S0(n6369_1), .Y(n2802));
MX2X1    g1337(.A(g829), .B(n3478), .S0(n6371), .Y(n2807));
INVX1    g1338(.A(g797), .Y(n3469));
MX2X1    g1339(.A(n3469), .B(g833), .S0(n6367), .Y(n2812));
MX2X1    g1340(.A(n3469), .B(g834), .S0(n6369_1), .Y(n2817));
MX2X1    g1341(.A(g832), .B(n3469), .S0(n6371), .Y(n2822));
INVX1    g1342(.A(g801), .Y(n3460));
MX2X1    g1343(.A(n3460), .B(g836), .S0(n6367), .Y(n2827));
MX2X1    g1344(.A(n3460), .B(g837), .S0(n6369_1), .Y(n2832));
MX2X1    g1345(.A(g835), .B(n3460), .S0(n6371), .Y(n2837));
INVX1    g1346(.A(g805), .Y(n3451));
MX2X1    g1347(.A(n3451), .B(g839), .S0(n6367), .Y(n2842));
MX2X1    g1348(.A(n3451), .B(g840), .S0(n6369_1), .Y(n2847));
MX2X1    g1349(.A(g838), .B(n3451), .S0(n6371), .Y(n2852));
INVX1    g1350(.A(g809), .Y(n3442));
MX2X1    g1351(.A(n3442), .B(g842), .S0(n6367), .Y(n2857));
MX2X1    g1352(.A(n3442), .B(g843), .S0(n6369_1), .Y(n2862));
MX2X1    g1353(.A(g841), .B(n3442), .S0(n6371), .Y(n2867));
INVX1    g1354(.A(g813), .Y(n3433));
MX2X1    g1355(.A(n3433), .B(g845), .S0(n6367), .Y(n2872));
MX2X1    g1356(.A(n3433), .B(g846), .S0(n6369_1), .Y(n2877));
MX2X1    g1357(.A(g844), .B(n3433), .S0(n6371), .Y(n2882));
INVX1    g1358(.A(g826), .Y(n6401));
NOR2X1   g1359(.A(g863), .B(n6401), .Y(n6402));
INVX1    g1360(.A(g823), .Y(n6403));
INVX1    g1361(.A(g853), .Y(n6404_1));
OAI22X1  g1362(.A0(g864), .A1(n6403), .B0(n6404_1), .B1(g862), .Y(n6405));
NOR2X1   g1363(.A(n6405), .B(n6402), .Y(n6406));
MX2X1    g1364(.A(n6406), .B(g848), .S0(n6367), .Y(n2887));
MX2X1    g1365(.A(n6406), .B(g849), .S0(n6369_1), .Y(n2892));
MX2X1    g1366(.A(g847), .B(n6406), .S0(n6371), .Y(n2897));
NOR2X1   g1367(.A(g860), .B(n6401), .Y(n6410));
OAI22X1  g1368(.A0(g861), .A1(n6403), .B0(n6404_1), .B1(g859), .Y(n6411));
NOR2X1   g1369(.A(n6411), .B(n6410), .Y(n6412));
MX2X1    g1370(.A(n6412), .B(g851), .S0(n6367), .Y(n2902));
MX2X1    g1371(.A(n6412), .B(g852), .S0(n6369_1), .Y(n2907));
MX2X1    g1372(.A(g850), .B(n6412), .S0(n6371), .Y(n2912));
NOR4X1   g1373(.A(g805), .B(g809), .C(n3433), .D(n3460), .Y(n6416));
AND2X1   g1374(.A(n1476), .B(g826), .Y(n6417));
MX2X1    g1375(.A(g857), .B(n6416), .S0(n6417), .Y(n2917));
AND2X1   g1376(.A(n1476), .B(g823), .Y(n6419_1));
MX2X1    g1377(.A(g858), .B(n6416), .S0(n6419_1), .Y(n2922));
AND2X1   g1378(.A(n1476), .B(g853), .Y(n6421));
MX2X1    g1379(.A(g856), .B(n6416), .S0(n6421), .Y(n2927));
MX2X1    g1380(.A(g860), .B(n3487), .S0(n6417), .Y(n2932));
MX2X1    g1381(.A(g861), .B(n3487), .S0(n6419_1), .Y(n2937));
MX2X1    g1382(.A(g859), .B(n3487), .S0(n6421), .Y(n2942));
MX2X1    g1383(.A(g863), .B(n3496), .S0(n6417), .Y(n2947));
MX2X1    g1384(.A(g864), .B(n3496), .S0(n6419_1), .Y(n2952));
MX2X1    g1385(.A(g862), .B(n3496), .S0(n6421), .Y(n2957));
NAND4X1  g1386(.A(g789), .B(g793), .C(g813), .D(g785), .Y(n6429_1));
NAND4X1  g1387(.A(g801), .B(g805), .C(g809), .D(g797), .Y(n6430));
NOR2X1   g1388(.A(n6430), .B(n6429_1), .Y(n6431));
INVX1    g1389(.A(n6431), .Y(n6432));
MX2X1    g1390(.A(g866), .B(n6432), .S0(n6417), .Y(n2962));
MX2X1    g1391(.A(g867), .B(n6432), .S0(n6419_1), .Y(n2967));
MX2X1    g1392(.A(g865), .B(n6432), .S0(n6421), .Y(n2972));
NOR2X1   g1393(.A(g851), .B(n6401), .Y(n6436));
OAI22X1  g1394(.A0(g852), .A1(n6403), .B0(n6404_1), .B1(g850), .Y(n6437));
OR2X1    g1395(.A(n6437), .B(n6436), .Y(n6438));
AND2X1   g1396(.A(n6438), .B(n6412), .Y(n6439_1));
NOR2X1   g1397(.A(g857), .B(n6401), .Y(n6440));
OAI22X1  g1398(.A0(g858), .A1(n6403), .B0(n6404_1), .B1(g856), .Y(n6441));
OAI21X1  g1399(.A0(n6441), .A1(n6440), .B0(g869), .Y(n6442));
NOR2X1   g1400(.A(g848), .B(n6401), .Y(n6443));
OAI22X1  g1401(.A0(g849), .A1(n6403), .B0(n6404_1), .B1(g847), .Y(n6444_1));
NOR2X1   g1402(.A(n6444_1), .B(n6443), .Y(n6445));
XOR2X1   g1403(.A(n6445), .B(n6406), .Y(n6446));
NOR2X1   g1404(.A(g842), .B(n6401), .Y(n6447));
OAI22X1  g1405(.A0(g843), .A1(n6403), .B0(n6404_1), .B1(g841), .Y(n6448));
NOR2X1   g1406(.A(n6448), .B(n6447), .Y(n6449_1));
XOR2X1   g1407(.A(n6449_1), .B(n3442), .Y(n6450));
NOR4X1   g1408(.A(n6446), .B(n6442), .C(n6439_1), .D(n6450), .Y(n6451));
NOR2X1   g1409(.A(g836), .B(n6401), .Y(n6452));
OAI22X1  g1410(.A0(g837), .A1(n6403), .B0(n6404_1), .B1(g835), .Y(n6453));
NOR2X1   g1411(.A(n6453), .B(n6452), .Y(n6454_1));
XOR2X1   g1412(.A(n6454_1), .B(n3460), .Y(n6455));
NOR2X1   g1413(.A(g833), .B(n6401), .Y(n6456));
OAI22X1  g1414(.A0(g834), .A1(n6403), .B0(n6404_1), .B1(g832), .Y(n6457));
NOR2X1   g1415(.A(n6457), .B(n6456), .Y(n6458));
XOR2X1   g1416(.A(n6458), .B(n3469), .Y(n6459_1));
NOR2X1   g1417(.A(g839), .B(n6401), .Y(n6460));
OAI22X1  g1418(.A0(g840), .A1(n6403), .B0(n6404_1), .B1(g838), .Y(n6461));
NOR2X1   g1419(.A(n6461), .B(n6460), .Y(n6462));
XOR2X1   g1420(.A(n6462), .B(n3451), .Y(n6463));
NOR2X1   g1421(.A(g845), .B(n6401), .Y(n6464_1));
OAI22X1  g1422(.A0(g846), .A1(n6403), .B0(n6404_1), .B1(g844), .Y(n6465));
OAI21X1  g1423(.A0(n6465), .A1(n6464_1), .B0(n3433), .Y(n6466));
OAI21X1  g1424(.A0(n6438), .A1(n6412), .B0(n6466), .Y(n6467));
NOR4X1   g1425(.A(n6463), .B(n6459_1), .C(n6455), .D(n6467), .Y(n6468));
NOR3X1   g1426(.A(n6465), .B(n6464_1), .C(n3433), .Y(n6469_1));
NOR2X1   g1427(.A(g830), .B(n6401), .Y(n6470));
OAI22X1  g1428(.A0(g831), .A1(n6403), .B0(n6404_1), .B1(g829), .Y(n6471));
NOR2X1   g1429(.A(n6471), .B(n6470), .Y(n6472));
XOR2X1   g1430(.A(n6472), .B(n3478), .Y(n6473));
NOR2X1   g1431(.A(g821), .B(n6401), .Y(n6474_1));
OAI22X1  g1432(.A0(g822), .A1(n6403), .B0(n6404_1), .B1(g820), .Y(n6475));
NOR2X1   g1433(.A(n6475), .B(n6474_1), .Y(n6476));
XOR2X1   g1434(.A(n6476), .B(n3487), .Y(n6477));
NOR2X1   g1435(.A(g818), .B(n6401), .Y(n6478));
OAI22X1  g1436(.A0(g819), .A1(n6403), .B0(n6404_1), .B1(g817), .Y(n6479_1));
NOR2X1   g1437(.A(n6479_1), .B(n6478), .Y(n6480));
XOR2X1   g1438(.A(n6480), .B(n3496), .Y(n6481));
NOR4X1   g1439(.A(n6477), .B(n6473), .C(n6469_1), .D(n6481), .Y(n6482));
NAND3X1  g1440(.A(n6482), .B(n6468), .C(n6451), .Y(n6483));
NAND2X1  g1441(.A(g909), .B(g826), .Y(n6484_1));
AOI22X1  g1442(.A0(g912), .A1(g823), .B0(g853), .B1(g915), .Y(n6485));
AND2X1   g1443(.A(n6485), .B(n6484_1), .Y(n6486));
NOR3X1   g1444(.A(n6486), .B(n6405), .C(n6402), .Y(n6487));
OR2X1    g1445(.A(g863), .B(n6401), .Y(n6488));
INVX1    g1446(.A(g864), .Y(n6489_1));
INVX1    g1447(.A(g862), .Y(n6490));
AOI22X1  g1448(.A0(n6489_1), .A1(g823), .B0(g853), .B1(n6490), .Y(n6491));
NAND2X1  g1449(.A(n6485), .B(n6484_1), .Y(n6492));
AOI21X1  g1450(.A0(n6491), .A1(n6488), .B0(n6492), .Y(n6493));
NAND2X1  g1451(.A(g900), .B(g826), .Y(n6494_1));
AOI22X1  g1452(.A0(g903), .A1(g823), .B0(g853), .B1(g906), .Y(n6495));
NAND2X1  g1453(.A(n6495), .B(n6494_1), .Y(n6496));
XOR2X1   g1454(.A(n6496), .B(g809), .Y(n6497));
NOR3X1   g1455(.A(n6497), .B(n6493), .C(n6487), .Y(n6498));
NAND2X1  g1456(.A(g873), .B(g826), .Y(n6499_1));
AOI22X1  g1457(.A0(g876), .A1(g823), .B0(g853), .B1(g879), .Y(n6500));
NAND2X1  g1458(.A(n6500), .B(n6499_1), .Y(n6501));
XOR2X1   g1459(.A(n6501), .B(g785), .Y(n6502));
NAND2X1  g1460(.A(g882), .B(g826), .Y(n6503));
AOI22X1  g1461(.A0(g885), .A1(g823), .B0(g853), .B1(g888), .Y(n6504_1));
NAND2X1  g1462(.A(n6504_1), .B(n6503), .Y(n6505));
XOR2X1   g1463(.A(n6505), .B(g793), .Y(n6506));
NAND2X1  g1464(.A(g891), .B(g826), .Y(n6507));
AOI22X1  g1465(.A0(g894), .A1(g823), .B0(g853), .B1(g897), .Y(n6508));
NAND2X1  g1466(.A(n6508), .B(n6507), .Y(n6509_1));
XOR2X1   g1467(.A(n6509_1), .B(g801), .Y(n6510));
OAI21X1  g1468(.A0(n6510), .A1(n6506), .B0(n6502), .Y(n6511));
NOR2X1   g1469(.A(n6511), .B(n6498), .Y(n6512));
NOR2X1   g1470(.A(n6510), .B(n6497), .Y(n6513));
OAI22X1  g1471(.A0(n6502), .A1(n6506), .B0(n6493), .B1(n6487), .Y(n6514_1));
NOR2X1   g1472(.A(n6514_1), .B(n6513), .Y(n6515));
XOR2X1   g1473(.A(n6509_1), .B(n3460), .Y(n6516));
NOR2X1   g1474(.A(n6502), .B(n6497), .Y(n6517));
NOR3X1   g1475(.A(n6506), .B(n6493), .C(n6487), .Y(n6518));
NOR3X1   g1476(.A(n6518), .B(n6517), .C(n6516), .Y(n6519_1));
NOR3X1   g1477(.A(n6519_1), .B(n6515), .C(n6512), .Y(n6520));
NAND2X1  g1478(.A(g954), .B(g826), .Y(n6521));
AOI22X1  g1479(.A0(g957), .A1(g823), .B0(g853), .B1(g960), .Y(n6522));
AND2X1   g1480(.A(n6522), .B(n6521), .Y(n6523));
NOR3X1   g1481(.A(n6523), .B(n6411), .C(n6410), .Y(n6524_1));
OR2X1    g1482(.A(g860), .B(n6401), .Y(n6525));
INVX1    g1483(.A(g861), .Y(n6526));
INVX1    g1484(.A(g859), .Y(n6527));
AOI22X1  g1485(.A0(n6526), .A1(g823), .B0(g853), .B1(n6527), .Y(n6528));
NAND2X1  g1486(.A(n6522), .B(n6521), .Y(n6529_1));
AOI21X1  g1487(.A0(n6528), .A1(n6525), .B0(n6529_1), .Y(n6530));
NAND2X1  g1488(.A(g945), .B(g826), .Y(n6531));
AOI22X1  g1489(.A0(g948), .A1(g823), .B0(g853), .B1(g951), .Y(n6532));
NAND2X1  g1490(.A(n6532), .B(n6531), .Y(n6533));
XOR2X1   g1491(.A(n6533), .B(g813), .Y(n6534_1));
NOR3X1   g1492(.A(n6534_1), .B(n6530), .C(n6524_1), .Y(n6535));
NAND2X1  g1493(.A(g918), .B(g826), .Y(n6536));
AOI22X1  g1494(.A0(g921), .A1(g823), .B0(g853), .B1(g924), .Y(n6537));
NAND2X1  g1495(.A(n6537), .B(n6536), .Y(n6538));
XOR2X1   g1496(.A(n6538), .B(g789), .Y(n6539_1));
NAND2X1  g1497(.A(g927), .B(g826), .Y(n6540));
AOI22X1  g1498(.A0(g930), .A1(g823), .B0(g853), .B1(g933), .Y(n6541));
NAND2X1  g1499(.A(n6541), .B(n6540), .Y(n6542));
XOR2X1   g1500(.A(n6542), .B(g797), .Y(n6543));
NAND2X1  g1501(.A(g936), .B(g826), .Y(n6544_1));
AOI22X1  g1502(.A0(g939), .A1(g823), .B0(g853), .B1(g942), .Y(n6545));
NAND2X1  g1503(.A(n6545), .B(n6544_1), .Y(n6546));
XOR2X1   g1504(.A(n6546), .B(g805), .Y(n6547));
OAI21X1  g1505(.A0(n6547), .A1(n6543), .B0(n6539_1), .Y(n6548));
NOR2X1   g1506(.A(n6548), .B(n6535), .Y(n6549_1));
NOR2X1   g1507(.A(n6547), .B(n6534_1), .Y(n6550));
OAI22X1  g1508(.A0(n6539_1), .A1(n6543), .B0(n6530), .B1(n6524_1), .Y(n6551));
NOR2X1   g1509(.A(n6551), .B(n6550), .Y(n6552));
XOR2X1   g1510(.A(n6546), .B(n3451), .Y(n6553));
NOR2X1   g1511(.A(n6539_1), .B(n6534_1), .Y(n6554_1));
NOR3X1   g1512(.A(n6543), .B(n6530), .C(n6524_1), .Y(n6555));
NOR3X1   g1513(.A(n6555), .B(n6554_1), .C(n6553), .Y(n6556));
NOR3X1   g1514(.A(n6556), .B(n6552), .C(n6549_1), .Y(n6557));
AOI21X1  g1515(.A0(n6557), .A1(n6520), .B0(n6442), .Y(n6558));
INVX1    g1516(.A(g963), .Y(n6559_1));
NOR2X1   g1517(.A(g1005), .B(n6559_1), .Y(n6560));
INVX1    g1518(.A(g1092), .Y(n6561));
INVX1    g1519(.A(g1088), .Y(n6562));
OAI22X1  g1520(.A0(g1006), .A1(n6561), .B0(n6562), .B1(g1007), .Y(n6563));
NOR2X1   g1521(.A(n6563), .B(n6560), .Y(n6564_1));
NOR2X1   g1522(.A(g1002), .B(n6559_1), .Y(n6565));
OAI22X1  g1523(.A0(g1003), .A1(n6561), .B0(n6562), .B1(g1004), .Y(n6566));
NOR2X1   g1524(.A(n6566), .B(n6565), .Y(n6567));
NOR2X1   g1525(.A(g999), .B(n6559_1), .Y(n6568));
OAI22X1  g1526(.A0(g1000), .A1(n6561), .B0(n6562), .B1(g1001), .Y(n6569_1));
NOR2X1   g1527(.A(n6569_1), .B(n6568), .Y(n6570));
INVX1    g1528(.A(n6570), .Y(n6571));
NOR2X1   g1529(.A(g1009), .B(n6559_1), .Y(n6572));
OAI22X1  g1530(.A0(g1010), .A1(n6561), .B0(n6562), .B1(g1008), .Y(n6573));
NOR2X1   g1531(.A(n6573), .B(n6572), .Y(n6574_1));
INVX1    g1532(.A(n6574_1), .Y(n6575));
NAND4X1  g1533(.A(n6571), .B(n6567), .C(n6564_1), .D(n6575), .Y(n6576));
NOR3X1   g1534(.A(n6576), .B(n6558), .C(n6483), .Y(n6577));
NOR4X1   g1535(.A(n6566), .B(n6565), .C(n6564_1), .D(n6570), .Y(n6578));
NAND2X1  g1536(.A(n6578), .B(n6575), .Y(n6579_1));
NOR2X1   g1537(.A(n6579_1), .B(n6483), .Y(n6580));
NOR2X1   g1538(.A(g1090), .B(n6559_1), .Y(n6581));
OAI22X1  g1539(.A0(g1091), .A1(n6561), .B0(n6562), .B1(g1089), .Y(n6582));
NOR2X1   g1540(.A(n6582), .B(n6581), .Y(n6583_1));
INVX1    g1541(.A(g869), .Y(n6584));
NOR3X1   g1542(.A(n6441), .B(n6440), .C(n6584), .Y(n6585));
INVX1    g1543(.A(n6585), .Y(n6586));
OAI22X1  g1544(.A0(n6583_1), .A1(n6483), .B0(n6570), .B1(n6586), .Y(n6587_1));
OR4X1    g1545(.A(n6565), .B(n6563), .C(n6560), .D(n6566), .Y(n6588));
NOR3X1   g1546(.A(n6569_1), .B(n6568), .C(n6588), .Y(n6589));
INVX1    g1547(.A(n6589), .Y(n6590));
INVX1    g1548(.A(n6567), .Y(n6591));
NAND3X1  g1549(.A(n6570), .B(n6591), .C(n6564_1), .Y(n6592_1));
INVX1    g1550(.A(n6564_1), .Y(n6593));
NOR3X1   g1551(.A(n6571), .B(n6567), .C(n6593), .Y(n6594));
NAND4X1  g1552(.A(n6507), .B(n6495), .C(n6494_1), .D(n6508), .Y(n6595));
OR4X1    g1553(.A(n6546), .B(n6533), .C(n6501), .D(n6595), .Y(n6596_1));
NAND4X1  g1554(.A(n6503), .B(n6485), .C(n6484_1), .D(n6504_1), .Y(n6597));
OR4X1    g1555(.A(n6542), .B(n6538), .C(n6529_1), .D(n6597), .Y(n6598));
OR2X1    g1556(.A(n6598), .B(n6596_1), .Y(n6599));
OR2X1    g1557(.A(n6599), .B(n6594), .Y(n6600_1));
NAND2X1  g1558(.A(n6542), .B(n6529_1), .Y(n6601));
NAND3X1  g1559(.A(n6538), .B(n6505), .C(n6492), .Y(n6602));
OR4X1    g1560(.A(n6601), .B(n6596_1), .C(n6592_1), .D(n6602), .Y(n6603));
AOI22X1  g1561(.A0(n6600_1), .A1(n6603), .B0(n6592_1), .B1(n6590), .Y(n6604));
NOR4X1   g1562(.A(n6587_1), .B(n6580), .C(n6577), .D(n6604), .Y(n6605_1));
INVX1    g1563(.A(n6605_1), .Y(n6606));
NAND2X1  g1564(.A(n6592_1), .B(n6590), .Y(n6607));
XOR2X1   g1565(.A(n6607), .B(n6501), .Y(n6608));
NOR3X1   g1566(.A(n6587_1), .B(n6580), .C(n6577), .Y(n6609));
AOI21X1  g1567(.A0(n6604), .A1(n6609), .B0(n3496), .Y(n6610_1));
MX2X1    g1568(.A(n6608), .B(n6610_1), .S0(n6606), .Y(n6611));
MX2X1    g1569(.A(g873), .B(n6611), .S0(g826), .Y(n2977));
MX2X1    g1570(.A(g876), .B(n6611), .S0(g823), .Y(n2982));
MX2X1    g1571(.A(g879), .B(n6611), .S0(g853), .Y(n2987));
AND2X1   g1572(.A(n6592_1), .B(n6501), .Y(n6615_1));
OAI21X1  g1573(.A0(n6592_1), .A1(n6501), .B0(n6607), .Y(n6616));
OR2X1    g1574(.A(n6616), .B(n6615_1), .Y(n6617));
XOR2X1   g1575(.A(n6617), .B(n6538), .Y(n6618));
NAND3X1  g1576(.A(n6604), .B(n6592_1), .C(n6609), .Y(n6619));
MX2X1    g1577(.A(n3487), .B(n6604), .S0(n6609), .Y(n6620_1));
AOI22X1  g1578(.A0(n6619), .A1(n6620_1), .B0(n6618), .B1(n6605_1), .Y(n6621));
MX2X1    g1579(.A(g918), .B(n6621), .S0(g826), .Y(n2992));
MX2X1    g1580(.A(g921), .B(n6621), .S0(g823), .Y(n2997));
MX2X1    g1581(.A(g924), .B(n6621), .S0(g853), .Y(n3002));
XOR2X1   g1582(.A(n6594), .B(n6538), .Y(n6625_1));
OR2X1    g1583(.A(n6625_1), .B(n6617), .Y(n6626));
XOR2X1   g1584(.A(n6626), .B(n6505), .Y(n6627));
MX2X1    g1585(.A(n3478), .B(n6604), .S0(n6609), .Y(n6628));
AOI22X1  g1586(.A0(n6627), .A1(n6605_1), .B0(n6619), .B1(n6628), .Y(n6629));
MX2X1    g1587(.A(g882), .B(n6629), .S0(g826), .Y(n3007));
MX2X1    g1588(.A(g885), .B(n6629), .S0(g823), .Y(n3012));
MX2X1    g1589(.A(g888), .B(n6629), .S0(g853), .Y(n3017));
XOR2X1   g1590(.A(n6594), .B(n6505), .Y(n6633));
OR4X1    g1591(.A(n6625_1), .B(n6616), .C(n6615_1), .D(n6633), .Y(n6634));
XOR2X1   g1592(.A(n6634), .B(n6542), .Y(n6635_1));
MX2X1    g1593(.A(n3469), .B(n6604), .S0(n6609), .Y(n6636));
AOI22X1  g1594(.A0(n6635_1), .A1(n6605_1), .B0(n6619), .B1(n6636), .Y(n6637));
MX2X1    g1595(.A(g927), .B(n6637), .S0(g826), .Y(n3022));
MX2X1    g1596(.A(g930), .B(n6637), .S0(g823), .Y(n3027));
MX2X1    g1597(.A(g933), .B(n6637), .S0(g853), .Y(n3032));
XOR2X1   g1598(.A(n6594), .B(n6542), .Y(n6641));
OR2X1    g1599(.A(n6641), .B(n6633), .Y(n6642));
NOR4X1   g1600(.A(n6625_1), .B(n6616), .C(n6615_1), .D(n6642), .Y(n6643));
XOR2X1   g1601(.A(n6643), .B(n6509_1), .Y(n6644));
AOI21X1  g1602(.A0(n6604), .A1(n6609), .B0(n3460), .Y(n6645_1));
MX2X1    g1603(.A(n6644), .B(n6645_1), .S0(n6606), .Y(n6646));
MX2X1    g1604(.A(g891), .B(n6646), .S0(g826), .Y(n3037));
MX2X1    g1605(.A(g894), .B(n6646), .S0(g823), .Y(n3042));
MX2X1    g1606(.A(g897), .B(n6646), .S0(g853), .Y(n3047));
XOR2X1   g1607(.A(n6592_1), .B(n6509_1), .Y(n6650_1));
AND2X1   g1608(.A(n6650_1), .B(n6643), .Y(n6651));
XOR2X1   g1609(.A(n6651), .B(n6546), .Y(n6652));
AOI21X1  g1610(.A0(n6604), .A1(n6609), .B0(n3451), .Y(n6653));
MX2X1    g1611(.A(n6652), .B(n6653), .S0(n6606), .Y(n6654));
MX2X1    g1612(.A(g936), .B(n6654), .S0(g826), .Y(n3052));
MX2X1    g1613(.A(g939), .B(n6654), .S0(g823), .Y(n3057));
MX2X1    g1614(.A(g942), .B(n6654), .S0(g853), .Y(n3062));
XOR2X1   g1615(.A(n6592_1), .B(n6546), .Y(n6658));
NAND2X1  g1616(.A(n6658), .B(n6650_1), .Y(n6659));
NOR4X1   g1617(.A(n6642), .B(n6625_1), .C(n6617), .D(n6659), .Y(n6660_1));
XOR2X1   g1618(.A(n6660_1), .B(n6496), .Y(n6661));
AOI21X1  g1619(.A0(n6604), .A1(n6609), .B0(n3442), .Y(n6662));
MX2X1    g1620(.A(n6661), .B(n6662), .S0(n6606), .Y(n6663));
MX2X1    g1621(.A(g900), .B(n6663), .S0(g826), .Y(n3067));
MX2X1    g1622(.A(g903), .B(n6663), .S0(g823), .Y(n3072));
MX2X1    g1623(.A(g906), .B(n6663), .S0(g853), .Y(n3077));
XOR2X1   g1624(.A(n6592_1), .B(n6496), .Y(n6667));
AND2X1   g1625(.A(n6667), .B(n6660_1), .Y(n6668));
XOR2X1   g1626(.A(n6668), .B(n6533), .Y(n6669));
AOI21X1  g1627(.A0(n6604), .A1(n6609), .B0(n3433), .Y(n6670_1));
MX2X1    g1628(.A(n6669), .B(n6670_1), .S0(n6606), .Y(n6671));
MX2X1    g1629(.A(g945), .B(n6671), .S0(g826), .Y(n3082));
MX2X1    g1630(.A(g948), .B(n6671), .S0(g823), .Y(n3087));
MX2X1    g1631(.A(g951), .B(n6671), .S0(g853), .Y(n3092));
XOR2X1   g1632(.A(n6592_1), .B(n6533), .Y(n6675_1));
NAND4X1  g1633(.A(n6667), .B(n6658), .C(n6650_1), .D(n6675_1), .Y(n6676));
OR4X1    g1634(.A(n6642), .B(n6625_1), .C(n6617), .D(n6676), .Y(n6677));
XOR2X1   g1635(.A(n6677), .B(n6492), .Y(n6678));
MX2X1    g1636(.A(n6406), .B(n6604), .S0(n6609), .Y(n6679));
AOI22X1  g1637(.A0(n6678), .A1(n6605_1), .B0(n6619), .B1(n6679), .Y(n6680_1));
MX2X1    g1638(.A(g909), .B(n6680_1), .S0(g826), .Y(n3097));
MX2X1    g1639(.A(g912), .B(n6680_1), .S0(g823), .Y(n3102));
MX2X1    g1640(.A(g915), .B(n6680_1), .S0(g853), .Y(n3107));
XOR2X1   g1641(.A(n6594), .B(n6492), .Y(n6684));
OR2X1    g1642(.A(n6684), .B(n6677), .Y(n6685_1));
XOR2X1   g1643(.A(n6685_1), .B(n6529_1), .Y(n6686));
MX2X1    g1644(.A(n6412), .B(n6604), .S0(n6609), .Y(n6687));
AOI22X1  g1645(.A0(n6686), .A1(n6605_1), .B0(n6619), .B1(n6687), .Y(n6688));
MX2X1    g1646(.A(g954), .B(n6688), .S0(g826), .Y(n3112));
MX2X1    g1647(.A(g957), .B(n6688), .S0(g823), .Y(n3117));
MX2X1    g1648(.A(g960), .B(n6688), .S0(g853), .Y(n3122));
INVX1    g1649(.A(g780), .Y(n6692));
NOR2X1   g1650(.A(n5399), .B(n6404_1), .Y(n6693));
XOR2X1   g1651(.A(n6693), .B(n6692), .Y(n6694));
AOI21X1  g1652(.A0(n6371), .A1(n5399), .B0(n6694), .Y(n3127));
INVX1    g1653(.A(g776), .Y(n6696));
NOR3X1   g1654(.A(n5399), .B(n6692), .C(n6404_1), .Y(n6697));
XOR2X1   g1655(.A(n6697), .B(n6696), .Y(n6698));
AOI21X1  g1656(.A0(n6371), .A1(n5399), .B0(n6698), .Y(n3132));
INVX1    g1657(.A(g771), .Y(n6700_1));
NOR4X1   g1658(.A(n6696), .B(n6692), .C(n6404_1), .D(n5399), .Y(n6701));
XOR2X1   g1659(.A(n6701), .B(n6700_1), .Y(n6702));
AOI21X1  g1660(.A0(n6371), .A1(n5399), .B0(n6702), .Y(n3137));
NAND2X1  g1661(.A(n6701), .B(g771), .Y(n6704));
XOR2X1   g1662(.A(n6704), .B(g767), .Y(n6705_1));
AOI21X1  g1663(.A0(n6371), .A1(n5399), .B0(n6705_1), .Y(n3142));
NAND3X1  g1664(.A(n6701), .B(g767), .C(g771), .Y(n6707));
XOR2X1   g1665(.A(n6707), .B(g762), .Y(n6708));
AOI21X1  g1666(.A0(n6371), .A1(n5399), .B0(n6708), .Y(n3147));
INVX1    g1667(.A(g767), .Y(n6710_1));
INVX1    g1668(.A(g762), .Y(n6711));
OR4X1    g1669(.A(g758), .B(n6711), .C(n6710_1), .D(n6704), .Y(n6712));
OAI21X1  g1670(.A0(n6707), .A1(n6711), .B0(g758), .Y(n6713));
AOI22X1  g1671(.A0(n6712), .A1(n6713), .B0(n6371), .B1(n5399), .Y(n3152));
INVX1    g1672(.A(g758), .Y(n6715_1));
OR4X1    g1673(.A(n6715_1), .B(n6711), .C(n6710_1), .D(n6704), .Y(n6716));
XOR2X1   g1674(.A(n6716), .B(g753), .Y(n6717));
AOI21X1  g1675(.A0(n6371), .A1(n5399), .B0(n6717), .Y(n3157));
INVX1    g1676(.A(g749), .Y(n6719));
INVX1    g1677(.A(g753), .Y(n6720_1));
NOR4X1   g1678(.A(n6720_1), .B(n6715_1), .C(n6711), .D(n6707), .Y(n6721));
XOR2X1   g1679(.A(n6721), .B(n6719), .Y(n6722));
AOI21X1  g1680(.A0(n6371), .A1(n5399), .B0(n6722), .Y(n3162));
INVX1    g1681(.A(g744), .Y(n6724));
AND2X1   g1682(.A(n6721), .B(g749), .Y(n6725_1));
XOR2X1   g1683(.A(n6725_1), .B(n6724), .Y(n6726));
AOI21X1  g1684(.A0(n6371), .A1(n5399), .B0(n6726), .Y(n3167));
INVX1    g1685(.A(g740), .Y(n6728));
NOR4X1   g1686(.A(n6724), .B(n6719), .C(n6720_1), .D(n6716), .Y(n6729));
XOR2X1   g1687(.A(n6729), .B(n6728), .Y(n6730_1));
AOI21X1  g1688(.A0(n6371), .A1(n5399), .B0(n6730_1), .Y(n3172));
NOR2X1   g1689(.A(g1071), .B(n6559_1), .Y(n6732));
OAI22X1  g1690(.A0(g1060), .A1(n6561), .B0(n6562), .B1(g1063), .Y(n6733));
NOR2X1   g1691(.A(g1056), .B(n6559_1), .Y(n6734));
OAI22X1  g1692(.A0(g1045), .A1(n6561), .B0(n6562), .B1(g1048), .Y(n6735_1));
NOR2X1   g1693(.A(n6735_1), .B(n6734), .Y(n6736));
OR4X1    g1694(.A(n6733), .B(n6732), .C(g3229), .D(n6736), .Y(n6737));
NOR2X1   g1695(.A(g1085), .B(n6559_1), .Y(n6738));
OAI22X1  g1696(.A0(g1075), .A1(n6561), .B0(n6562), .B1(g1078), .Y(n6739));
NOR2X1   g1697(.A(n6739), .B(n6738), .Y(n6740_1));
OAI21X1  g1698(.A0(n6740_1), .A1(n5718), .B0(n6737), .Y(n6741));
INVX1    g1699(.A(n6736), .Y(n3554));
INVX1    g1700(.A(n6740_1), .Y(n3564));
NOR2X1   g1701(.A(g1041), .B(n6559_1), .Y(n6744));
OAI22X1  g1702(.A0(g1030), .A1(n6561), .B0(n6562), .B1(g1033), .Y(n6745_1));
NOR2X1   g1703(.A(n6745_1), .B(n6744), .Y(n6746));
NOR4X1   g1704(.A(n3564), .B(n3554), .C(n5718), .D(n6746), .Y(n6747));
NOR4X1   g1705(.A(n6739), .B(n6738), .C(g3229), .D(n6746), .Y(n6748));
NOR2X1   g1706(.A(n6733), .B(n6732), .Y(n6749));
NOR3X1   g1707(.A(n6746), .B(n6749), .C(n5718), .Y(n6750_1));
NOR4X1   g1708(.A(n6748), .B(n6747), .C(n6741), .D(n6750_1), .Y(n6751));
NOR4X1   g1709(.A(n6568), .B(n6567), .C(n6564_1), .D(n6569_1), .Y(n6752));
AOI21X1  g1710(.A0(n6590), .A1(n5399), .B0(n6752), .Y(n3569));
AND2X1   g1711(.A(n3569), .B(g963), .Y(n6754));
MX2X1    g1712(.A(g1041), .B(n6751), .S0(n6754), .Y(n3208));
AND2X1   g1713(.A(n3569), .B(g1092), .Y(n6756));
MX2X1    g1714(.A(g1030), .B(n6751), .S0(n6756), .Y(n3213));
AND2X1   g1715(.A(n3569), .B(g1088), .Y(n6758));
MX2X1    g1716(.A(g1033), .B(n6751), .S0(n6758), .Y(n3218));
NOR4X1   g1717(.A(n6744), .B(n6749), .C(g3229), .D(n6745_1), .Y(n6760_1));
NOR3X1   g1718(.A(n6736), .B(n6733), .C(n6732), .Y(n6761));
NOR3X1   g1719(.A(n6761), .B(n6760_1), .C(n6750_1), .Y(n6762));
MX2X1    g1720(.A(g1056), .B(n6762), .S0(n6754), .Y(n3223));
MX2X1    g1721(.A(g1045), .B(n6762), .S0(n6756), .Y(n3228));
MX2X1    g1722(.A(g1048), .B(n6762), .S0(n6758), .Y(n3233));
NOR4X1   g1723(.A(n6744), .B(n6736), .C(n5718), .D(n6745_1), .Y(n6766));
NOR3X1   g1724(.A(n6746), .B(n6736), .C(g3229), .Y(n6767));
INVX1    g1725(.A(n6746), .Y(n3549));
NOR4X1   g1726(.A(n3564), .B(n3554), .C(g3229), .D(n3549), .Y(n6769));
NOR4X1   g1727(.A(n6767), .B(n6766), .C(n6747), .D(n6769), .Y(n6770_1));
MX2X1    g1728(.A(g1071), .B(n6770_1), .S0(n6754), .Y(n3238));
MX2X1    g1729(.A(g1060), .B(n6770_1), .S0(n6756), .Y(n3243));
MX2X1    g1730(.A(g1063), .B(n6770_1), .S0(n6758), .Y(n3248));
NOR2X1   g1731(.A(n6746), .B(g3229), .Y(n6774));
NOR3X1   g1732(.A(n6745_1), .B(n6744), .C(n5718), .Y(n6775_1));
NOR4X1   g1733(.A(n6734), .B(n6733), .C(n6732), .D(n6735_1), .Y(n6776));
OAI21X1  g1734(.A0(n6775_1), .A1(n6774), .B0(n6776), .Y(n6777));
MX2X1    g1735(.A(g1085), .B(n6777), .S0(n6754), .Y(n3253));
MX2X1    g1736(.A(g1075), .B(n6777), .S0(n6756), .Y(n3258));
MX2X1    g1737(.A(g1078), .B(n6777), .S0(n6758), .Y(n3263));
NAND2X1  g1738(.A(g1095), .B(g963), .Y(n6781));
AOI22X1  g1739(.A0(g1098), .A1(g1092), .B0(g1088), .B1(g1101), .Y(n6782));
AND2X1   g1740(.A(n6782), .B(n6781), .Y(n6783));
INVX1    g1741(.A(n6783), .Y(n6784));
OR4X1    g1742(.A(n6432), .B(n6412), .C(n6406), .D(n6585), .Y(n6785_1));
NAND2X1  g1743(.A(g1104), .B(g963), .Y(n6786));
AOI22X1  g1744(.A0(g1107), .A1(g1092), .B0(g1088), .B1(g1110), .Y(n6787));
AND2X1   g1745(.A(n6787), .B(n6786), .Y(n6788));
AND2X1   g1746(.A(n6788), .B(n6785_1), .Y(n6789));
NOR3X1   g1747(.A(n6432), .B(n6412), .C(n6406), .Y(n6790_1));
INVX1    g1748(.A(n6790_1), .Y(n6791));
OAI21X1  g1749(.A0(n6788), .A1(n6791), .B0(n6783), .Y(n6792));
INVX1    g1750(.A(n6788), .Y(n3514));
NOR2X1   g1751(.A(g1114), .B(n6559_1), .Y(n6794));
OAI22X1  g1752(.A0(g1115), .A1(n6561), .B0(n6562), .B1(g1113), .Y(n6795_1));
NOR2X1   g1753(.A(n6795_1), .B(n6794), .Y(n6796));
INVX1    g1754(.A(n6796), .Y(n6797));
NOR4X1   g1755(.A(n3514), .B(n6791), .C(n6585), .D(n6797), .Y(n6798));
NAND2X1  g1756(.A(n6796), .B(n3514), .Y(n6799));
OAI21X1  g1757(.A0(n6799), .A1(n6790_1), .B0(n6784), .Y(n6800_1));
OAI22X1  g1758(.A0(n6798), .A1(n6800_1), .B0(n6792), .B1(n6789), .Y(n6801));
AND2X1   g1759(.A(n6801), .B(g996), .Y(n6802));
XOR2X1   g1760(.A(n6802), .B(n6784), .Y(n6803));
MX2X1    g1761(.A(g1095), .B(n6803), .S0(g963), .Y(n3268));
MX2X1    g1762(.A(g1098), .B(n6803), .S0(g1092), .Y(n3273));
MX2X1    g1763(.A(g1101), .B(n6803), .S0(g1088), .Y(n3278));
INVX1    g1764(.A(g996), .Y(n6807));
NAND4X1  g1765(.A(n6788), .B(n6790_1), .C(n6585), .D(n6783), .Y(n6808));
OAI21X1  g1766(.A0(n6797), .A1(n6585), .B0(n6790_1), .Y(n6809));
NAND2X1  g1767(.A(n6809), .B(n6788), .Y(n6810_1));
OAI21X1  g1768(.A0(n6796), .A1(n6790_1), .B0(n3514), .Y(n6811));
NAND3X1  g1769(.A(n6811), .B(n6810_1), .C(n6784), .Y(n6812));
AOI21X1  g1770(.A0(n6812), .A1(n6808), .B0(n6807), .Y(n6813));
XOR2X1   g1771(.A(n6813), .B(n3514), .Y(n6814));
MX2X1    g1772(.A(g1104), .B(n6814), .S0(g963), .Y(n3283));
MX2X1    g1773(.A(g1107), .B(n6814), .S0(g1092), .Y(n3288));
MX2X1    g1774(.A(g1110), .B(n6814), .S0(g1088), .Y(n3293));
MX2X1    g1775(.A(n6785_1), .B(n6790_1), .S0(n3514), .Y(n6818));
OR4X1    g1776(.A(n6797), .B(n6783), .C(n6807), .D(n6818), .Y(n6819));
NAND3X1  g1777(.A(n6782), .B(n6781), .C(g996), .Y(n6820_1));
OAI21X1  g1778(.A0(n6820_1), .A1(n6818), .B0(n6819), .Y(n6821));
AND2X1   g1779(.A(n6821), .B(g963), .Y(n6822));
MX2X1    g1780(.A(g1114), .B(n6819), .S0(n6822), .Y(n3298));
AND2X1   g1781(.A(n6821), .B(g1092), .Y(n6824));
MX2X1    g1782(.A(g1115), .B(n6819), .S0(n6824), .Y(n3303));
AND2X1   g1783(.A(n6821), .B(g1088), .Y(n6826));
MX2X1    g1784(.A(g1113), .B(n6819), .S0(n6826), .Y(n3308));
NAND2X1  g1785(.A(g1116), .B(g963), .Y(n6828));
AOI22X1  g1786(.A0(g1119), .A1(g1092), .B0(g1088), .B1(g1122), .Y(n6829));
NAND2X1  g1787(.A(n6829), .B(n6828), .Y(n6830_1));
OR2X1    g1788(.A(g866), .B(n6401), .Y(n6831));
INVX1    g1789(.A(g867), .Y(n6832));
INVX1    g1790(.A(g865), .Y(n6833));
AOI22X1  g1791(.A0(n6832), .A1(g823), .B0(g853), .B1(n6833), .Y(n6834));
AOI21X1  g1792(.A0(n6834), .A1(n6831), .B0(n6432), .Y(n6835_1));
MX2X1    g1793(.A(n6830_1), .B(n6835_1), .S0(g996), .Y(n6836));
MX2X1    g1794(.A(g1116), .B(n6836), .S0(g963), .Y(n3313));
MX2X1    g1795(.A(g1119), .B(n6836), .S0(g1092), .Y(n3318));
MX2X1    g1796(.A(g1122), .B(n6836), .S0(g1088), .Y(n3323));
NAND2X1  g1797(.A(g1125), .B(g963), .Y(n6840));
AOI22X1  g1798(.A0(g1128), .A1(g1092), .B0(g1088), .B1(g1131), .Y(n6841));
AND2X1   g1799(.A(n6841), .B(n6840), .Y(n6842));
INVX1    g1800(.A(n6842), .Y(n6843));
NOR2X1   g1801(.A(n6842), .B(n6830_1), .Y(n6844_1));
INVX1    g1802(.A(n6844_1), .Y(n6845));
AND2X1   g1803(.A(n6842), .B(n6830_1), .Y(n6846));
INVX1    g1804(.A(n6846), .Y(n6847));
MX2X1    g1805(.A(n6845), .B(n6847), .S0(n6835_1), .Y(n6848_1));
NOR2X1   g1806(.A(g1135), .B(n6559_1), .Y(n6849));
OAI22X1  g1807(.A0(g1136), .A1(n6561), .B0(n6562), .B1(g1134), .Y(n6850));
OAI21X1  g1808(.A0(n6850), .A1(n6849), .B0(g996), .Y(n6851));
NOR2X1   g1809(.A(n6851), .B(n6848_1), .Y(n6852));
XOR2X1   g1810(.A(n6852), .B(n6843), .Y(n6853_1));
MX2X1    g1811(.A(g1125), .B(n6853_1), .S0(g963), .Y(n3328));
MX2X1    g1812(.A(g1128), .B(n6853_1), .S0(g1092), .Y(n3333));
MX2X1    g1813(.A(g1131), .B(n6853_1), .S0(g1088), .Y(n3338));
NOR4X1   g1814(.A(n6849), .B(n6848_1), .C(n6807), .D(n6850), .Y(n6857_1));
INVX1    g1815(.A(n6857_1), .Y(n6858));
NOR2X1   g1816(.A(n6843), .B(n6830_1), .Y(n6859));
AOI22X1  g1817(.A0(n6840), .A1(n6841), .B0(n6829), .B1(n6828), .Y(n6860));
MX2X1    g1818(.A(n6860), .B(n6859), .S0(n6835_1), .Y(n6861));
AOI21X1  g1819(.A0(n6861), .A1(g996), .B0(n6857_1), .Y(n6862_1));
NOR2X1   g1820(.A(n6862_1), .B(n6559_1), .Y(n6863));
MX2X1    g1821(.A(g1135), .B(n6858), .S0(n6863), .Y(n3343));
NOR2X1   g1822(.A(n6862_1), .B(n6561), .Y(n6865));
MX2X1    g1823(.A(g1136), .B(n6858), .S0(n6865), .Y(n3348));
NOR2X1   g1824(.A(n6862_1), .B(n6562), .Y(n6867));
MX2X1    g1825(.A(g1134), .B(n6858), .S0(n6867), .Y(n3353));
OAI21X1  g1826(.A0(n6591), .A1(n6564_1), .B0(n6558), .Y(n6869));
AOI21X1  g1827(.A0(n6869), .A1(n6571), .B0(n6594), .Y(n6870));
OR2X1    g1828(.A(n6583_1), .B(n6483), .Y(n6871_1));
OAI21X1  g1829(.A0(n6870), .A1(n6570), .B0(n6871_1), .Y(n6872));
AOI21X1  g1830(.A0(n6870), .A1(n6570), .B0(n6872), .Y(n6873));
MX2X1    g1831(.A(g999), .B(n6873), .S0(g963), .Y(n3358));
MX2X1    g1832(.A(g1000), .B(n6873), .S0(g1092), .Y(n3363));
MX2X1    g1833(.A(g1001), .B(n6873), .S0(g1088), .Y(n3368));
INVX1    g1834(.A(n6442), .Y(n6877));
NAND3X1  g1835(.A(n6553), .B(n6516), .C(n6498), .Y(n6878));
NOR2X1   g1836(.A(n6506), .B(n6502), .Y(n6879));
NAND2X1  g1837(.A(n6535), .B(n6879), .Y(n6880_1));
OR4X1    g1838(.A(n6878), .B(n6543), .C(n6539_1), .D(n6880_1), .Y(n6881));
NAND2X1  g1839(.A(n6881), .B(n6877), .Y(n6882));
NOR4X1   g1840(.A(n6574_1), .B(n6558), .C(n6483), .D(n6882), .Y(n6883));
NOR2X1   g1841(.A(n6557), .B(n6442), .Y(n6884_1));
OAI21X1  g1842(.A0(n6881), .A1(n6442), .B0(n6586), .Y(n6885));
OR4X1    g1843(.A(n6563), .B(n6560), .C(n6884_1), .D(n6885), .Y(n6886));
NAND4X1  g1844(.A(n6482), .B(n6468), .C(n6451), .D(n6575), .Y(n6887));
NOR2X1   g1845(.A(n6585), .B(n6564_1), .Y(n6888));
AOI21X1  g1846(.A0(n6888), .A1(n6887), .B0(n6591), .Y(n6889_1));
OAI21X1  g1847(.A0(n6886), .A1(n6883), .B0(n6889_1), .Y(n6890));
OR2X1    g1848(.A(n6511), .B(n6498), .Y(n6891));
OR2X1    g1849(.A(n6514_1), .B(n6513), .Y(n6892));
OR2X1    g1850(.A(n6502), .B(n6497), .Y(n6893_1));
NAND3X1  g1851(.A(n6492), .B(n6491), .C(n6488), .Y(n6894));
OAI21X1  g1852(.A0(n6405), .A1(n6402), .B0(n6486), .Y(n6895));
XOR2X1   g1853(.A(n6505), .B(n3478), .Y(n6896));
NAND3X1  g1854(.A(n6896), .B(n6895), .C(n6894), .Y(n6897));
NAND3X1  g1855(.A(n6897), .B(n6893_1), .C(n6510), .Y(n6898_1));
NAND3X1  g1856(.A(n6898_1), .B(n6892), .C(n6891), .Y(n6899));
AOI21X1  g1857(.A0(n6899), .A1(n6877), .B0(n6593), .Y(n6900));
OAI21X1  g1858(.A0(n6882), .A1(n6884_1), .B0(n6900), .Y(n6901));
AOI21X1  g1859(.A0(n6899), .A1(n6877), .B0(n6564_1), .Y(n6902_1));
NOR2X1   g1860(.A(n6902_1), .B(n6567), .Y(n6903));
AOI21X1  g1861(.A0(n6903), .A1(n6901), .B0(n6570), .Y(n6904));
AOI22X1  g1862(.A0(n6890), .A1(n6904), .B0(n6570), .B1(n6588), .Y(n6905));
OAI21X1  g1863(.A0(n6905), .A1(n6567), .B0(n6871_1), .Y(n6906));
AOI21X1  g1864(.A0(n6905), .A1(n6567), .B0(n6906), .Y(n6907_1));
MX2X1    g1865(.A(g1002), .B(n6907_1), .S0(g963), .Y(n3373));
MX2X1    g1866(.A(g1003), .B(n6907_1), .S0(g1092), .Y(n3378));
MX2X1    g1867(.A(g1004), .B(n6907_1), .S0(g1088), .Y(n3383));
AOI21X1  g1868(.A0(n6885), .A1(n6564_1), .B0(n6567), .Y(n6912));
OAI21X1  g1869(.A0(n6882), .A1(n6564_1), .B0(n6912), .Y(n6913));
NOR2X1   g1870(.A(n6520), .B(n6442), .Y(n6914));
OR4X1    g1871(.A(n6884_1), .B(n6914), .C(n6807), .D(n6593), .Y(n6915));
AOI21X1  g1872(.A0(n6915), .A1(n6567), .B0(n6570), .Y(n6916_1));
AOI22X1  g1873(.A0(n6913), .A1(n6916_1), .B0(n6570), .B1(n6564_1), .Y(n6917));
XOR2X1   g1874(.A(n6917), .B(n6593), .Y(n6918));
AND2X1   g1875(.A(n6918), .B(n6871_1), .Y(n6919));
MX2X1    g1876(.A(g1005), .B(n6919), .S0(g963), .Y(n3388));
MX2X1    g1877(.A(g1006), .B(n6919), .S0(g1092), .Y(n3393));
MX2X1    g1878(.A(g1007), .B(n6919), .S0(g1088), .Y(n3398));
NOR3X1   g1879(.A(n6593), .B(n6558), .C(n6483), .Y(n6923));
NOR3X1   g1880(.A(n6591), .B(n6564_1), .C(n6483), .Y(n6924));
OAI21X1  g1881(.A0(n6924), .A1(n6923), .B0(n6571), .Y(n6925));
MX2X1    g1882(.A(n6882), .B(n6807), .S0(n6578), .Y(n6926_1));
NOR2X1   g1883(.A(n6926_1), .B(n6559_1), .Y(n6927));
MX2X1    g1884(.A(g1009), .B(n6925), .S0(n6927), .Y(n3403));
NOR2X1   g1885(.A(n6926_1), .B(n6561), .Y(n6929));
MX2X1    g1886(.A(g1010), .B(n6925), .S0(n6929), .Y(n3408));
NOR2X1   g1887(.A(n6926_1), .B(n6562), .Y(n6931_1));
MX2X1    g1888(.A(g1008), .B(n6925), .S0(n6931_1), .Y(n3413));
NAND4X1  g1889(.A(n6482), .B(n6468), .C(n6451), .D(n6583_1), .Y(n6933));
AND2X1   g1890(.A(g996), .B(g963), .Y(n6934));
MX2X1    g1891(.A(g1090), .B(n6933), .S0(n6934), .Y(n3418));
AND2X1   g1892(.A(g996), .B(g1092), .Y(n6936_1));
MX2X1    g1893(.A(g1091), .B(n6933), .S0(n6936_1), .Y(n3423));
AND2X1   g1894(.A(g996), .B(g1088), .Y(n6938));
MX2X1    g1895(.A(g1089), .B(n6933), .S0(n6938), .Y(n3428));
INVX1    g1896(.A(g986), .Y(n6940));
NAND3X1  g1897(.A(n5930), .B(n5928), .C(g1092), .Y(n6941_1));
AOI21X1  g1898(.A0(g992), .A1(n6561), .B0(n6940), .Y(n6942));
AOI22X1  g1899(.A0(n6941_1), .A1(n6942), .B0(g985), .B1(n6940), .Y(n3519));
NAND3X1  g1900(.A(n5934), .B(n5933), .C(g1092), .Y(n6944));
AOI21X1  g1901(.A0(g995), .A1(n6561), .B0(n6940), .Y(n6945));
NOR2X1   g1902(.A(g987), .B(g986), .Y(n6946_1));
AOI21X1  g1903(.A0(n6945), .A1(n6944), .B0(n6946_1), .Y(n3524));
NAND3X1  g1904(.A(n5938), .B(n5937), .C(g1092), .Y(n6948));
AOI21X1  g1905(.A0(g984), .A1(n6561), .B0(n6940), .Y(n6949));
NOR2X1   g1906(.A(g988), .B(g986), .Y(n6950));
AOI21X1  g1907(.A0(n6949), .A1(n6948), .B0(n6950), .Y(n3529));
NAND3X1  g1908(.A(n5942), .B(n5941_1), .C(g1092), .Y(n6952));
AOI21X1  g1909(.A0(g983), .A1(n6561), .B0(n6940), .Y(n6953));
NOR2X1   g1910(.A(g989), .B(g986), .Y(n6954));
AOI21X1  g1911(.A0(n6953), .A1(n6952), .B0(n6954), .Y(n3534));
NAND3X1  g1912(.A(n5946_1), .B(n5945), .C(g1092), .Y(n6956_1));
AOI21X1  g1913(.A0(g982), .A1(n6561), .B0(n6940), .Y(n6957));
NOR2X1   g1914(.A(g990), .B(g986), .Y(n6958));
AOI21X1  g1915(.A0(n6957), .A1(n6956_1), .B0(n6958), .Y(n3539));
NAND3X1  g1916(.A(n5950), .B(n5949), .C(g1092), .Y(n6960));
AOI21X1  g1917(.A0(g981), .A1(n6561), .B0(n6940), .Y(n6961_1));
NOR2X1   g1918(.A(g991), .B(g986), .Y(n6962));
AOI21X1  g1919(.A0(n6961_1), .A1(n6960), .B0(n6962), .Y(n3544));
INVX1    g1920(.A(n6749), .Y(n3559));
NOR3X1   g1921(.A(n6599), .B(n6571), .C(n6588), .Y(n6965));
XOR2X1   g1922(.A(n6509_1), .B(n6711), .Y(n6966_1));
XOR2X1   g1923(.A(n6533), .B(n6719), .Y(n6967));
XOR2X1   g1924(.A(n6546), .B(n6715_1), .Y(n6968));
NAND3X1  g1925(.A(n6968), .B(n6967), .C(n6966_1), .Y(n6969));
XOR2X1   g1926(.A(n6529_1), .B(n6728), .Y(n6970));
XOR2X1   g1927(.A(n6538), .B(n6696), .Y(n6971_1));
XOR2X1   g1928(.A(n6496), .B(n6720_1), .Y(n6972));
XOR2X1   g1929(.A(n6492), .B(n6724), .Y(n6973));
NAND4X1  g1930(.A(n6972), .B(n6971_1), .C(n6970), .D(n6973), .Y(n6974));
XOR2X1   g1931(.A(n6542), .B(g767), .Y(n6975));
XOR2X1   g1932(.A(n6505), .B(g771), .Y(n6976_1));
XOR2X1   g1933(.A(n6501), .B(g780), .Y(n6977));
OR2X1    g1934(.A(n6977), .B(n6976_1), .Y(n6978));
OR4X1    g1935(.A(n6975), .B(n6752), .C(n5399), .D(n6978), .Y(n6979));
NOR3X1   g1936(.A(n6979), .B(n6974), .C(n6969), .Y(n6980));
OAI21X1  g1937(.A0(n6980), .A1(n6965), .B0(n3569), .Y(n3574));
MX2X1    g1938(.A(g1240), .B(n5982), .S0(g1236), .Y(n3713));
INVX1    g1939(.A(g1236), .Y(n6983));
INVX1    g1940(.A(g1240), .Y(n6984));
MX2X1    g1941(.A(n6984), .B(g1243), .S0(n6983), .Y(n3718));
MX2X1    g1942(.A(g1196), .B(g1243), .S0(g1236), .Y(n3723));
NAND2X1  g1943(.A(g1255), .B(g1231), .Y(n6987));
AOI22X1  g1944(.A0(g1257), .A1(g1237), .B0(g1236), .B1(g1259), .Y(n6988));
AND2X1   g1945(.A(n6988), .B(n6987), .Y(n3728));
MX2X1    g1946(.A(g1173), .B(n6843), .S0(g1161), .Y(n3808));
MX2X1    g1947(.A(g1174), .B(n6843), .S0(g1168), .Y(n3813));
MX2X1    g1948(.A(g1175), .B(n6843), .S0(g1172), .Y(n3818));
MX2X1    g1949(.A(g1142), .B(n6752), .S0(g1161), .Y(n3823));
MX2X1    g1950(.A(g1145), .B(n6752), .S0(g1168), .Y(n3828));
MX2X1    g1951(.A(g1148), .B(n6752), .S0(g1172), .Y(n3833));
MX2X1    g1952(.A(g1164), .B(n6578), .S0(g1161), .Y(n3838));
MX2X1    g1953(.A(g1165), .B(n6578), .S0(g1168), .Y(n3843));
MX2X1    g1954(.A(g1166), .B(n6578), .S0(g1172), .Y(n3848));
MX2X1    g1955(.A(g1167), .B(n6788), .S0(g1161), .Y(n3853));
MX2X1    g1956(.A(g1171), .B(n6788), .S0(g1168), .Y(n3858));
MX2X1    g1957(.A(g1151), .B(n6788), .S0(g1172), .Y(n3863));
MX2X1    g1958(.A(g1152), .B(n6589), .S0(g1161), .Y(n3868));
MX2X1    g1959(.A(g1155), .B(n6589), .S0(g1168), .Y(n3873));
MX2X1    g1960(.A(g1158), .B(n6589), .S0(g1172), .Y(n3878));
NAND2X1  g1961(.A(g1251), .B(g1231), .Y(n7005));
AOI22X1  g1962(.A0(g1253), .A1(g1237), .B0(g1236), .B1(g1176), .Y(n7006));
AND2X1   g1963(.A(n7006), .B(n7005), .Y(n3883));
INVX1    g1964(.A(g1237), .Y(n7008_1));
NOR2X1   g1965(.A(g1164), .B(n7008_1), .Y(n7009));
INVX1    g1966(.A(g1231), .Y(n7010));
OAI22X1  g1967(.A0(g1165), .A1(n6983), .B0(n7010), .B1(g1166), .Y(n7011));
NOR2X1   g1968(.A(n7011), .B(n7009), .Y(n3896));
NOR2X1   g1969(.A(g1167), .B(n7008_1), .Y(n7013));
OAI22X1  g1970(.A0(g1171), .A1(n6983), .B0(n7010), .B1(g1151), .Y(n7014));
NOR2X1   g1971(.A(n7014), .B(n7013), .Y(n3910));
NOR2X1   g1972(.A(g1173), .B(n7008_1), .Y(n7016));
OAI22X1  g1973(.A0(g1174), .A1(n6983), .B0(n7010), .B1(g1175), .Y(n7017_1));
NOR2X1   g1974(.A(n7017_1), .B(n7016), .Y(n3919));
NOR2X1   g1975(.A(g1268), .B(n7010), .Y(n7019));
OAI22X1  g1976(.A0(g1269), .A1(n7008_1), .B0(n6983), .B1(g1267), .Y(n7020));
NOR2X1   g1977(.A(g1265), .B(n7010), .Y(n7021_1));
OAI22X1  g1978(.A0(g1266), .A1(n7008_1), .B0(n6983), .B1(g1264), .Y(n7022));
NOR2X1   g1979(.A(n7022), .B(n7021_1), .Y(n7023));
OR4X1    g1980(.A(n7020), .B(n7019), .C(g3229), .D(n7023), .Y(n7024));
NOR2X1   g1981(.A(g1271), .B(n7010), .Y(n7025));
OAI22X1  g1982(.A0(g1272), .A1(n7008_1), .B0(n6983), .B1(g1270), .Y(n7026_1));
NOR2X1   g1983(.A(n7026_1), .B(n7025), .Y(n7027));
OAI21X1  g1984(.A0(n7027), .A1(n5718), .B0(n7024), .Y(n7028));
INVX1    g1985(.A(n7023), .Y(n4083));
INVX1    g1986(.A(n7027), .Y(n4073));
NOR2X1   g1987(.A(g1262), .B(n7010), .Y(n7031));
OAI22X1  g1988(.A0(g1263), .A1(n7008_1), .B0(n6983), .B1(g1261), .Y(n7032));
NOR2X1   g1989(.A(n7032), .B(n7031), .Y(n7033));
NOR4X1   g1990(.A(n4073), .B(n4083), .C(n5718), .D(n7033), .Y(n7034));
NOR4X1   g1991(.A(n7026_1), .B(n7025), .C(g3229), .D(n7033), .Y(n7035_1));
NOR2X1   g1992(.A(n7020), .B(n7019), .Y(n7036));
NOR3X1   g1993(.A(n7033), .B(n7036), .C(n5718), .Y(n7037));
NOR4X1   g1994(.A(n7035_1), .B(n7034), .C(n7028), .D(n7037), .Y(n7038));
NAND2X1  g1995(.A(g1177), .B(g1231), .Y(n7039_1));
AOI22X1  g1996(.A0(g1180), .A1(g1237), .B0(g1236), .B1(g1183), .Y(n7040));
AND2X1   g1997(.A(n7040), .B(n7039_1), .Y(n7041));
INVX1    g1998(.A(n7041), .Y(n7042));
NAND2X1  g1999(.A(g1300), .B(g1231), .Y(n7043));
AOI22X1  g2000(.A0(g1303), .A1(g1237), .B0(g1236), .B1(g1306), .Y(n7044_1));
AND2X1   g2001(.A(n7044_1), .B(n7043), .Y(n7045));
INVX1    g2002(.A(n7045), .Y(n7046));
NAND3X1  g2003(.A(n7041), .B(n7046), .C(g1196), .Y(n7047));
NAND2X1  g2004(.A(g1291), .B(g1231), .Y(n7048_1));
AOI22X1  g2005(.A0(g1294), .A1(g1237), .B0(g1236), .B1(g1297), .Y(n7049));
AND2X1   g2006(.A(n7049), .B(n7048_1), .Y(n7050));
INVX1    g2007(.A(n7050), .Y(n7051));
AOI22X1  g2008(.A0(n7047), .A1(n6049), .B0(n7042), .B1(n7051), .Y(n4068));
NAND2X1  g2009(.A(n4068), .B(g1231), .Y(n7053_1));
MX2X1    g2010(.A(n7038), .B(g1262), .S0(n7053_1), .Y(n3928));
NAND2X1  g2011(.A(n4068), .B(g1237), .Y(n7055));
MX2X1    g2012(.A(n7038), .B(g1263), .S0(n7055), .Y(n3933));
NAND2X1  g2013(.A(n4068), .B(g1236), .Y(n7057_1));
MX2X1    g2014(.A(n7038), .B(g1261), .S0(n7057_1), .Y(n3938));
NOR4X1   g2015(.A(n7031), .B(n7036), .C(g3229), .D(n7032), .Y(n7059));
NOR3X1   g2016(.A(n7023), .B(n7020), .C(n7019), .Y(n7060));
NOR3X1   g2017(.A(n7060), .B(n7059), .C(n7037), .Y(n7061));
MX2X1    g2018(.A(n7061), .B(g1265), .S0(n7053_1), .Y(n3943));
MX2X1    g2019(.A(n7061), .B(g1266), .S0(n7055), .Y(n3948));
MX2X1    g2020(.A(n7061), .B(g1264), .S0(n7057_1), .Y(n3953));
NOR4X1   g2021(.A(n7031), .B(n7023), .C(n5718), .D(n7032), .Y(n7065));
NOR3X1   g2022(.A(n7033), .B(n7023), .C(g3229), .Y(n7066_1));
INVX1    g2023(.A(n7033), .Y(n4088));
NOR4X1   g2024(.A(n4073), .B(n4083), .C(g3229), .D(n4088), .Y(n7068));
NOR4X1   g2025(.A(n7066_1), .B(n7065), .C(n7034), .D(n7068), .Y(n7069));
MX2X1    g2026(.A(n7069), .B(g1268), .S0(n7053_1), .Y(n3958));
MX2X1    g2027(.A(n7069), .B(g1269), .S0(n7055), .Y(n3963));
MX2X1    g2028(.A(n7069), .B(g1267), .S0(n7057_1), .Y(n3968));
NOR2X1   g2029(.A(n7033), .B(g3229), .Y(n7073));
NOR3X1   g2030(.A(n7032), .B(n7031), .C(n5718), .Y(n7074));
NOR4X1   g2031(.A(n7021_1), .B(n7020), .C(n7019), .D(n7022), .Y(n7075_1));
OAI21X1  g2032(.A0(n7074), .A1(n7073), .B0(n7075_1), .Y(n7076));
MX2X1    g2033(.A(n7076), .B(g1271), .S0(n7053_1), .Y(n3973));
MX2X1    g2034(.A(n7076), .B(g1272), .S0(n7055), .Y(n3978));
MX2X1    g2035(.A(n7076), .B(g1270), .S0(n7057_1), .Y(n3983));
INVX1    g2036(.A(n3728), .Y(n7080_1));
AND2X1   g2037(.A(g1210), .B(g185), .Y(n7081));
NAND2X1  g2038(.A(g1273), .B(g1231), .Y(n7082));
AOI22X1  g2039(.A0(g1276), .A1(g1237), .B0(g1236), .B1(g1279), .Y(n7083));
NAND2X1  g2040(.A(n7083), .B(n7082), .Y(n7084_1));
AOI21X1  g2041(.A0(n7081), .A1(n7080_1), .B0(n7084_1), .Y(n7085));
NOR2X1   g2042(.A(n7085), .B(n5981_1), .Y(n7086));
MX2X1    g2043(.A(g1273), .B(n7086), .S0(g1231), .Y(n3988));
MX2X1    g2044(.A(g1276), .B(n7086), .S0(g1237), .Y(n3993));
MX2X1    g2045(.A(g1279), .B(n7086), .S0(g1236), .Y(n3998));
INVX1    g2046(.A(n3883), .Y(n7090));
AND2X1   g2047(.A(g1228), .B(g185), .Y(n7091));
NAND2X1  g2048(.A(g1282), .B(g1231), .Y(n7092));
AOI22X1  g2049(.A0(g1285), .A1(g1237), .B0(g1236), .B1(g1288), .Y(n7093_1));
NAND2X1  g2050(.A(n7093_1), .B(n7092), .Y(n7094));
AOI21X1  g2051(.A0(n7091), .A1(n7090), .B0(n7094), .Y(n7095));
NOR2X1   g2052(.A(n7095), .B(n5981_1), .Y(n7096));
MX2X1    g2053(.A(g1282), .B(n7096), .S0(g1231), .Y(n4003));
MX2X1    g2054(.A(g1285), .B(n7096), .S0(g1237), .Y(n4008));
MX2X1    g2055(.A(g1288), .B(n7096), .S0(g1236), .Y(n4013));
OR4X1    g2056(.A(n7031), .B(n7022), .C(n7021_1), .D(n7032), .Y(n7100));
NAND2X1  g2057(.A(g1012), .B(g1036), .Y(n7101));
AOI22X1  g2058(.A0(g1018), .A1(g1038), .B0(g1040), .B1(g1024), .Y(n7102_1));
AND2X1   g2059(.A(n7102_1), .B(n7101), .Y(n7103));
INVX1    g2060(.A(n7103), .Y(n7104));
NAND2X1  g2061(.A(g1012), .B(g1051), .Y(n7105));
AOI22X1  g2062(.A0(g1018), .A1(g1053), .B0(g1055), .B1(g1024), .Y(n7106_1));
AND2X1   g2063(.A(n7106_1), .B(n7105), .Y(n7107));
NAND2X1  g2064(.A(g1012), .B(g1066), .Y(n7108));
AOI22X1  g2065(.A0(g1018), .A1(g1068), .B0(g1070), .B1(g1024), .Y(n7109));
AND2X1   g2066(.A(n7109), .B(n7108), .Y(n7110_1));
OR4X1    g2067(.A(n7107), .B(n7104), .C(n7100), .D(n7110_1), .Y(n7111));
INVX1    g2068(.A(n7036), .Y(n4078));
INVX1    g2069(.A(n7107), .Y(n7113));
NAND2X1  g2070(.A(g1012), .B(g1081), .Y(n7114));
NAND2X1  g2071(.A(g1024), .B(g1011), .Y(n7115_1));
NAND2X1  g2072(.A(g1018), .B(g1083), .Y(n7116));
NAND3X1  g2073(.A(n7116), .B(n7115_1), .C(n7114), .Y(n7117));
NAND2X1  g2074(.A(n7117), .B(n7113), .Y(n7118));
OR4X1    g2075(.A(n7103), .B(n7023), .C(n4078), .D(n7118), .Y(n7119));
AND2X1   g2076(.A(n7110_1), .B(n7103), .Y(n7120_1));
NAND3X1  g2077(.A(n7120_1), .B(n7113), .C(n7075_1), .Y(n7121));
INVX1    g2078(.A(n7110_1), .Y(n7122));
NOR4X1   g2079(.A(n7032), .B(n7031), .C(n7036), .D(n7103), .Y(n7123));
NAND3X1  g2080(.A(n7123), .B(n7122), .C(n7113), .Y(n7124));
NAND4X1  g2081(.A(n7121), .B(n7119), .C(n7111), .D(n7124), .Y(n7125_1));
OR4X1    g2082(.A(n7103), .B(n4088), .C(n4073), .D(n7117), .Y(n7126));
AND2X1   g2083(.A(n7107), .B(n7103), .Y(n7127));
NAND3X1  g2084(.A(n7127), .B(n4088), .C(n7023), .Y(n7128));
NAND4X1  g2085(.A(n7103), .B(n4088), .C(n4073), .D(n7117), .Y(n7129));
OR4X1    g2086(.A(n7113), .B(n7033), .C(n7036), .D(n7110_1), .Y(n7130_1));
NAND4X1  g2087(.A(n7129), .B(n7128), .C(n7126), .D(n7130_1), .Y(n7131));
OR4X1    g2088(.A(n7103), .B(n7033), .C(n7036), .D(n7113), .Y(n7132));
OAI21X1  g2089(.A0(n7026_1), .A1(n7025), .B0(n7120_1), .Y(n7133));
OR4X1    g2090(.A(n7107), .B(n7103), .C(n7023), .D(n7122), .Y(n7134_1));
OR4X1    g2091(.A(n7032), .B(n7031), .C(n7036), .D(n7117), .Y(n7135));
NAND4X1  g2092(.A(n7134_1), .B(n7133), .C(n7132), .D(n7135), .Y(n7136));
OR4X1    g2093(.A(n7023), .B(n7020), .C(n7019), .D(n7103), .Y(n7137));
OR2X1    g2094(.A(n7113), .B(n7103), .Y(n7138_1));
OR4X1    g2095(.A(n7033), .B(n7026_1), .C(n7025), .D(n7110_1), .Y(n7139));
OAI22X1  g2096(.A0(n7138_1), .A1(n7139), .B0(n7137), .B1(n7122), .Y(n7140));
NOR4X1   g2097(.A(n7136), .B(n7131), .C(n7125_1), .D(n7140), .Y(n7141));
NAND4X1  g2098(.A(n7113), .B(n7103), .C(n7027), .D(n7122), .Y(n7142));
NOR3X1   g2099(.A(n7142), .B(n7033), .C(n4083), .Y(n7143_1));
NAND4X1  g2100(.A(n7113), .B(n7104), .C(n7036), .D(n7117), .Y(n7144));
NOR2X1   g2101(.A(n7144), .B(n7100), .Y(n7145));
NOR4X1   g2102(.A(n7103), .B(n7100), .C(n4073), .D(n7122), .Y(n7146));
NOR4X1   g2103(.A(n7104), .B(n7033), .C(n7036), .D(n7118), .Y(n7147_1));
OR4X1    g2104(.A(n7146), .B(n7145), .C(n7143_1), .D(n7147_1), .Y(n7148));
NAND4X1  g2105(.A(n7107), .B(n7033), .C(n4083), .D(n7122), .Y(n7149));
OR4X1    g2106(.A(n7107), .B(n7103), .C(n7027), .D(n7110_1), .Y(n7150));
OR4X1    g2107(.A(n7104), .B(n7033), .C(n7023), .D(n7122), .Y(n7151));
NAND3X1  g2108(.A(n7151), .B(n7150), .C(n7149), .Y(n7152_1));
NAND2X1  g2109(.A(n7123), .B(n7107), .Y(n7153));
NAND2X1  g2110(.A(n7127), .B(n7060), .Y(n7154));
OR4X1    g2111(.A(n7033), .B(n4083), .C(n4078), .D(n7117), .Y(n7155));
NAND3X1  g2112(.A(n7155), .B(n7154), .C(n7153), .Y(n7156_1));
NOR3X1   g2113(.A(n7156_1), .B(n7152_1), .C(n7148), .Y(n7157));
NAND2X1  g2114(.A(n7157), .B(n7095), .Y(n7158));
OR2X1    g2115(.A(n7158), .B(n7141), .Y(n7159));
INVX1    g2116(.A(n7085), .Y(n7160));
NOR2X1   g2117(.A(n7095), .B(n7160), .Y(n7161_1));
AOI21X1  g2118(.A0(n7161_1), .A1(n7157), .B0(n5982), .Y(n7162));
AOI22X1  g2119(.A0(n7159), .A1(n7162), .B0(n7045), .B1(n5982), .Y(n7163));
MX2X1    g2120(.A(g1300), .B(n7163), .S0(g1231), .Y(n4018));
MX2X1    g2121(.A(g1303), .B(n7163), .S0(g1237), .Y(n4023));
MX2X1    g2122(.A(g1306), .B(n7163), .S0(g1236), .Y(n4028));
NAND3X1  g2123(.A(n7141), .B(n7095), .C(n7160), .Y(n7167));
NOR2X1   g2124(.A(n7157), .B(n7160), .Y(n7168));
AOI21X1  g2125(.A0(n7168), .A1(n7141), .B0(n5982), .Y(n7169));
AOI22X1  g2126(.A0(n7167), .A1(n7169), .B0(n7050), .B1(n5982), .Y(n7170_1));
MX2X1    g2127(.A(g1291), .B(n7170_1), .S0(g1231), .Y(n4033));
MX2X1    g2128(.A(g1294), .B(n7170_1), .S0(g1237), .Y(n4038));
MX2X1    g2129(.A(g1297), .B(n7170_1), .S0(g1236), .Y(n4043));
INVX1    g2130(.A(g1196), .Y(n7174_1));
NOR3X1   g2131(.A(n7042), .B(n7046), .C(n7174_1), .Y(n7175));
MX2X1    g2132(.A(g1177), .B(n7175), .S0(g1231), .Y(n4048));
MX2X1    g2133(.A(g1180), .B(n7175), .S0(g1237), .Y(n4053));
MX2X1    g2134(.A(g1183), .B(n7175), .S0(g1236), .Y(n4058));
NAND3X1  g2135(.A(n6184_1), .B(n6183), .C(g1237), .Y(n7179_1));
AOI21X1  g2136(.A0(g1202), .A1(n7008_1), .B0(g1192), .Y(n7180));
INVX1    g2137(.A(g1192), .Y(n7181));
NOR2X1   g2138(.A(g1201), .B(n7181), .Y(n7182));
AOI21X1  g2139(.A0(n7180), .A1(n7179_1), .B0(n7182), .Y(n4093));
NAND3X1  g2140(.A(n6188), .B(n6187), .C(g1237), .Y(n7184));
AOI21X1  g2141(.A0(g1203), .A1(n7008_1), .B0(g1192), .Y(n7185));
NOR2X1   g2142(.A(g1200), .B(n7181), .Y(n7186));
AOI21X1  g2143(.A0(n7185), .A1(n7184), .B0(n7186), .Y(n4098));
NAND3X1  g2144(.A(n6192), .B(n6191), .C(g1237), .Y(n7188_1));
AOI21X1  g2145(.A0(g1204), .A1(n7008_1), .B0(g1192), .Y(n7189));
NOR2X1   g2146(.A(g1195), .B(n7181), .Y(n7190));
AOI21X1  g2147(.A0(n7189), .A1(n7188_1), .B0(n7190), .Y(n4103));
NAND3X1  g2148(.A(n6196), .B(n6195), .C(g1237), .Y(n7192_1));
AOI21X1  g2149(.A0(g1205), .A1(n7008_1), .B0(g1192), .Y(n7193));
NOR2X1   g2150(.A(g1194), .B(n7181), .Y(n7194));
AOI21X1  g2151(.A0(n7193), .A1(n7192_1), .B0(n7194), .Y(n4108));
NAND2X1  g2152(.A(n2412), .B(g1237), .Y(n7196));
AOI21X1  g2153(.A0(g1206), .A1(n7008_1), .B0(g1192), .Y(n7197_1));
NOR2X1   g2154(.A(g1193), .B(n7181), .Y(n7198));
AOI21X1  g2155(.A0(n7197_1), .A1(n7196), .B0(n7198), .Y(n4113));
INVX1    g2156(.A(g1138), .Y(n4122));
INVX1    g2157(.A(g1140), .Y(n4127));
INVX1    g2158(.A(g966), .Y(n4132));
INVX1    g2159(.A(g968), .Y(n4137));
INVX1    g2160(.A(g970), .Y(n4142));
INVX1    g2161(.A(g972), .Y(n4147));
INVX1    g2162(.A(g974), .Y(n4152));
INVX1    g2163(.A(g976), .Y(n4157));
INVX1    g2164(.A(g978), .Y(n4167));
MX2X1    g2165(.A(n4167), .B(g992), .S0(n5718), .Y(n4162));
MX2X1    g2166(.A(g1316), .B(g1196), .S0(g1315), .Y(n4185));
MX2X1    g2167(.A(g1345), .B(n6049), .S0(g1315), .Y(n4190));
INVX1    g2168(.A(g1345), .Y(n7212));
INVX1    g2169(.A(g1326), .Y(n7213));
NAND3X1  g2170(.A(n7213), .B(n7212), .C(g1315), .Y(n7214));
INVX1    g2171(.A(g1315), .Y(n7215_1));
OAI21X1  g2172(.A0(g1345), .A1(n7215_1), .B0(g1326), .Y(n7216));
AND2X1   g2173(.A(g1316), .B(g1312), .Y(n7217));
AOI21X1  g2174(.A0(n7216), .A1(n7214), .B0(n7217), .Y(n4195));
INVX1    g2175(.A(g1319), .Y(n7219));
NOR3X1   g2176(.A(n7213), .B(g1345), .C(n7215_1), .Y(n7220_1));
XOR2X1   g2177(.A(n7220_1), .B(n7219), .Y(n7221));
NOR2X1   g2178(.A(n7221), .B(n7217), .Y(n4200));
INVX1    g2179(.A(g1339), .Y(n7223));
NOR4X1   g2180(.A(n7213), .B(g1345), .C(n7215_1), .D(n7219), .Y(n7224));
XOR2X1   g2181(.A(n7224), .B(n7223), .Y(n7225_1));
NOR2X1   g2182(.A(n7225_1), .B(n7217), .Y(n4205));
INVX1    g2183(.A(g1332), .Y(n7227));
AND2X1   g2184(.A(n7224), .B(g1339), .Y(n7228));
XOR2X1   g2185(.A(n7228), .B(n7227), .Y(n7229));
NOR2X1   g2186(.A(n7229), .B(n7217), .Y(n4210));
NAND3X1  g2187(.A(n7224), .B(g1332), .C(g1339), .Y(n7231));
XOR2X1   g2188(.A(n7231), .B(g1346), .Y(n7232));
NOR2X1   g2189(.A(n7232), .B(n7217), .Y(n4215));
INVX1    g2190(.A(g1346), .Y(n7234));
OAI21X1  g2191(.A0(n7231), .A1(n7234), .B0(g1358), .Y(n7235_1));
INVX1    g2192(.A(g1358), .Y(n7236));
NAND4X1  g2193(.A(n7236), .B(g1346), .C(g1332), .D(n7228), .Y(n7237));
AOI21X1  g2194(.A0(n7237), .A1(n7235_1), .B0(n7217), .Y(n4220));
INVX1    g2195(.A(g1352), .Y(n7239));
NOR3X1   g2196(.A(n7231), .B(n7236), .C(n7234), .Y(n7240_1));
XOR2X1   g2197(.A(n7240_1), .B(n7239), .Y(n7241));
NOR2X1   g2198(.A(n7241), .B(n7217), .Y(n4225));
INVX1    g2199(.A(g1365), .Y(n7243));
NOR4X1   g2200(.A(n7239), .B(n7236), .C(n7234), .D(n7231), .Y(n7244));
XOR2X1   g2201(.A(n7244), .B(n7243), .Y(n7245_1));
NOR2X1   g2202(.A(n7245_1), .B(n7217), .Y(n4230));
INVX1    g2203(.A(g1372), .Y(n7247));
AND2X1   g2204(.A(n7244), .B(g1365), .Y(n7248));
XOR2X1   g2205(.A(n7248), .B(n7247), .Y(n7249));
NOR2X1   g2206(.A(n7249), .B(n7217), .Y(n4235));
NAND3X1  g2207(.A(n7244), .B(g1372), .C(g1365), .Y(n7251));
XOR2X1   g2208(.A(n7251), .B(g1378), .Y(n7252));
NOR2X1   g2209(.A(n7252), .B(n7217), .Y(n4240));
NAND4X1  g2210(.A(g1309), .B(g1224), .C(g1211), .D(n7212), .Y(n7254));
MX2X1    g2211(.A(n7213), .B(g1385), .S0(n7254), .Y(n4245));
NAND4X1  g2212(.A(g1312), .B(g1224), .C(g1211), .D(n7212), .Y(n7256));
MX2X1    g2213(.A(n7213), .B(g1386), .S0(n7256), .Y(n4250));
NAND4X1  g2214(.A(g1315), .B(g1224), .C(g1211), .D(n7212), .Y(n7258));
MX2X1    g2215(.A(n7213), .B(g1384), .S0(n7258), .Y(n4255));
MX2X1    g2216(.A(n7219), .B(g1388), .S0(n7254), .Y(n4260));
MX2X1    g2217(.A(n7219), .B(g1389), .S0(n7256), .Y(n4265));
MX2X1    g2218(.A(n7219), .B(g1387), .S0(n7258), .Y(n4270));
MX2X1    g2219(.A(n7223), .B(g1391), .S0(n7254), .Y(n4275));
MX2X1    g2220(.A(n7223), .B(g1392), .S0(n7256), .Y(n4280));
MX2X1    g2221(.A(n7223), .B(g1390), .S0(n7258), .Y(n4285));
MX2X1    g2222(.A(n7227), .B(g1394), .S0(n7254), .Y(n4290));
MX2X1    g2223(.A(n7227), .B(g1395), .S0(n7256), .Y(n4295));
MX2X1    g2224(.A(n7227), .B(g1393), .S0(n7258), .Y(n4300));
MX2X1    g2225(.A(n7234), .B(g1397), .S0(n7254), .Y(n4305));
MX2X1    g2226(.A(n7234), .B(g1398), .S0(n7256), .Y(n4310));
MX2X1    g2227(.A(n7234), .B(g1396), .S0(n7258), .Y(n4315));
MX2X1    g2228(.A(n7236), .B(g1400), .S0(n7254), .Y(n4320));
MX2X1    g2229(.A(n7236), .B(g1401), .S0(n7256), .Y(n4325));
MX2X1    g2230(.A(n7236), .B(g1399), .S0(n7258), .Y(n4330));
MX2X1    g2231(.A(n7239), .B(g1403), .S0(n7254), .Y(n4335));
MX2X1    g2232(.A(n7239), .B(g1404), .S0(n7256), .Y(n4340));
MX2X1    g2233(.A(n7239), .B(g1402), .S0(n7258), .Y(n4345));
MX2X1    g2234(.A(n7243), .B(g1406), .S0(n7254), .Y(n4350));
MX2X1    g2235(.A(n7243), .B(g1407), .S0(n7256), .Y(n4355));
MX2X1    g2236(.A(n7243), .B(g1405), .S0(n7258), .Y(n4360));
MX2X1    g2237(.A(n7247), .B(g1409), .S0(n7254), .Y(n4365));
MX2X1    g2238(.A(n7247), .B(g1410), .S0(n7256), .Y(n4370));
MX2X1    g2239(.A(n7247), .B(g1408), .S0(n7258), .Y(n4375));
INVX1    g2240(.A(g1378), .Y(n7284));
MX2X1    g2241(.A(n7284), .B(g1412), .S0(n7254), .Y(n4380));
MX2X1    g2242(.A(n7284), .B(g1413), .S0(n7256), .Y(n4385));
MX2X1    g2243(.A(n7284), .B(g1411), .S0(n7258), .Y(n4390));
AND2X1   g2244(.A(g1316), .B(g1309), .Y(n7288));
MX2X1    g2245(.A(g1415), .B(n7045), .S0(n7288), .Y(n4395));
MX2X1    g2246(.A(g1416), .B(n7045), .S0(n7217), .Y(n4400));
AND2X1   g2247(.A(g1316), .B(g1315), .Y(n7291));
MX2X1    g2248(.A(g1414), .B(n7045), .S0(n7291), .Y(n4405));
MX2X1    g2249(.A(g1418), .B(n7050), .S0(n7288), .Y(n4410));
MX2X1    g2250(.A(g1419), .B(n7050), .S0(n7217), .Y(n4415));
MX2X1    g2251(.A(g1417), .B(n7050), .S0(n7291), .Y(n4420));
INVX1    g2252(.A(g1309), .Y(n7296));
NOR2X1   g2253(.A(g1403), .B(n7296), .Y(n7297));
INVX1    g2254(.A(g1312), .Y(n7298_1));
OAI22X1  g2255(.A0(g1404), .A1(n7298_1), .B0(n7215_1), .B1(g1402), .Y(n7299));
OR2X1    g2256(.A(n7299), .B(n7297), .Y(n7300));
XOR2X1   g2257(.A(n7300), .B(g1352), .Y(n7301));
NOR2X1   g2258(.A(g1409), .B(n7296), .Y(n7302_1));
OAI22X1  g2259(.A0(g1410), .A1(n7298_1), .B0(n7215_1), .B1(g1408), .Y(n7303));
NOR2X1   g2260(.A(n7303), .B(n7302_1), .Y(n7304));
XOR2X1   g2261(.A(n7304), .B(n7247), .Y(n7305));
NOR2X1   g2262(.A(g1406), .B(n7296), .Y(n7306));
OAI22X1  g2263(.A0(g1407), .A1(n7298_1), .B0(n7215_1), .B1(g1405), .Y(n7307_1));
NOR2X1   g2264(.A(n7307_1), .B(n7306), .Y(n7308));
XOR2X1   g2265(.A(n7308), .B(n7243), .Y(n7309));
NOR2X1   g2266(.A(g1400), .B(n7296), .Y(n7310));
OAI22X1  g2267(.A0(g1401), .A1(n7298_1), .B0(n7215_1), .B1(g1399), .Y(n7311));
NOR2X1   g2268(.A(n7311), .B(n7310), .Y(n7312_1));
XOR2X1   g2269(.A(n7312_1), .B(n7236), .Y(n7313));
OR4X1    g2270(.A(n7309), .B(n7305), .C(n7301), .D(n7313), .Y(n7314));
INVX1    g2271(.A(g1395), .Y(n7315));
INVX1    g2272(.A(g1393), .Y(n7316_1));
AOI22X1  g2273(.A0(n7315), .A1(g1312), .B0(g1315), .B1(n7316_1), .Y(n7317));
OAI21X1  g2274(.A0(g1394), .A1(n7296), .B0(n7317), .Y(n7318));
XOR2X1   g2275(.A(n7318), .B(n7227), .Y(n7319));
NOR2X1   g2276(.A(g1397), .B(n7296), .Y(n7320));
OAI22X1  g2277(.A0(g1398), .A1(n7298_1), .B0(n7215_1), .B1(g1396), .Y(n7321_1));
NOR2X1   g2278(.A(n7321_1), .B(n7320), .Y(n7322));
XOR2X1   g2279(.A(n7322), .B(g1346), .Y(n7323));
NAND2X1  g2280(.A(n7323), .B(n7319), .Y(n7324));
NOR2X1   g2281(.A(g1385), .B(n7296), .Y(n7325_1));
OAI22X1  g2282(.A0(g1386), .A1(n7298_1), .B0(n7215_1), .B1(g1384), .Y(n7326));
NOR2X1   g2283(.A(n7326), .B(n7325_1), .Y(n7327));
XOR2X1   g2284(.A(n7327), .B(g1326), .Y(n7328));
INVX1    g2285(.A(g1389), .Y(n7329));
INVX1    g2286(.A(g1387), .Y(n7330_1));
AOI22X1  g2287(.A0(n7329), .A1(g1312), .B0(g1315), .B1(n7330_1), .Y(n7331));
OAI21X1  g2288(.A0(g1388), .A1(n7296), .B0(n7331), .Y(n7332));
XOR2X1   g2289(.A(n7332), .B(n7219), .Y(n7333));
NAND2X1  g2290(.A(n7333), .B(n7328), .Y(n7334));
NOR2X1   g2291(.A(g1412), .B(n7296), .Y(n7335_1));
OAI22X1  g2292(.A0(g1413), .A1(n7298_1), .B0(n7215_1), .B1(g1411), .Y(n7336));
NOR2X1   g2293(.A(n7336), .B(n7335_1), .Y(n7337));
XOR2X1   g2294(.A(n7337), .B(n7284), .Y(n7338));
NOR2X1   g2295(.A(g1391), .B(n7296), .Y(n7339));
OAI22X1  g2296(.A0(g1392), .A1(n7298_1), .B0(n7215_1), .B1(g1390), .Y(n7340_1));
NOR2X1   g2297(.A(n7340_1), .B(n7339), .Y(n7341));
XOR2X1   g2298(.A(n7341), .B(n7223), .Y(n7342));
OR2X1    g2299(.A(n7342), .B(n7338), .Y(n7343));
NOR4X1   g2300(.A(n7334), .B(n7324), .C(n7314), .D(n7343), .Y(n7344));
INVX1    g2301(.A(g1419), .Y(n7345_1));
INVX1    g2302(.A(g1417), .Y(n7346));
AOI22X1  g2303(.A0(n7345_1), .A1(g1312), .B0(g1315), .B1(n7346), .Y(n7347));
OAI21X1  g2304(.A0(g1418), .A1(n7296), .B0(n7347), .Y(n7348));
NOR2X1   g2305(.A(g1415), .B(n7296), .Y(n7349));
OAI22X1  g2306(.A0(g1416), .A1(n7298_1), .B0(n7215_1), .B1(g1414), .Y(n7350_1));
NOR4X1   g2307(.A(n7349), .B(n7348), .C(n7344), .D(n7350_1), .Y(n7351));
MX2X1    g2308(.A(n7351), .B(g1421), .S0(n7254), .Y(n4425));
MX2X1    g2309(.A(n7351), .B(g1422), .S0(n7256), .Y(n4430));
MX2X1    g2310(.A(n7351), .B(g1420), .S0(n7258), .Y(n4435));
INVX1    g2311(.A(g1316), .Y(n7355_1));
INVX1    g2312(.A(g1211), .Y(n7356));
INVX1    g2313(.A(g1224), .Y(n7357));
NOR3X1   g2314(.A(g1345), .B(n7357), .C(n7356), .Y(n7358));
OAI21X1  g2315(.A0(n7358), .A1(g1316), .B0(g1309), .Y(n7359));
MX2X1    g2316(.A(n7355_1), .B(g1424), .S0(n7359), .Y(n4440));
OAI21X1  g2317(.A0(n7358), .A1(g1316), .B0(g1312), .Y(n7361));
MX2X1    g2318(.A(n7355_1), .B(g1425), .S0(n7361), .Y(n4445));
OAI21X1  g2319(.A0(n7358), .A1(g1316), .B0(g1315), .Y(n7363));
MX2X1    g2320(.A(n7355_1), .B(g1423), .S0(n7363), .Y(n4450));
INVX1    g2321(.A(g1471), .Y(n5197));
NAND2X1  g2322(.A(g1563), .B(g1520), .Y(n7366));
MX2X1    g2323(.A(n5197), .B(g1512), .S0(n7366), .Y(n4468));
NAND2X1  g2324(.A(g1563), .B(g1517), .Y(n7368));
MX2X1    g2325(.A(n5197), .B(g1513), .S0(n7368), .Y(n4473));
AND2X1   g2326(.A(g1563), .B(g1547), .Y(n7370_1));
MX2X1    g2327(.A(g1511), .B(n5197), .S0(n7370_1), .Y(n4478));
INVX1    g2328(.A(g1476), .Y(n5188));
MX2X1    g2329(.A(n5188), .B(g1515), .S0(n7366), .Y(n4483));
MX2X1    g2330(.A(n5188), .B(g1516), .S0(n7368), .Y(n4488));
MX2X1    g2331(.A(g1514), .B(n5188), .S0(n7370_1), .Y(n4493));
INVX1    g2332(.A(g1481), .Y(n5179));
MX2X1    g2333(.A(n5179), .B(g1524), .S0(n7366), .Y(n4498));
MX2X1    g2334(.A(n5179), .B(g1525), .S0(n7368), .Y(n4503));
MX2X1    g2335(.A(g1523), .B(n5179), .S0(n7370_1), .Y(n4508));
INVX1    g2336(.A(g1486), .Y(n5170));
MX2X1    g2337(.A(n5170), .B(g1527), .S0(n7366), .Y(n4513));
MX2X1    g2338(.A(n5170), .B(g1528), .S0(n7368), .Y(n4518));
MX2X1    g2339(.A(g1526), .B(n5170), .S0(n7370_1), .Y(n4523));
INVX1    g2340(.A(g1491), .Y(n5161));
MX2X1    g2341(.A(n5161), .B(g1530), .S0(n7366), .Y(n4528));
MX2X1    g2342(.A(n5161), .B(g1531), .S0(n7368), .Y(n4533));
MX2X1    g2343(.A(g1529), .B(n5161), .S0(n7370_1), .Y(n4538));
INVX1    g2344(.A(g1496), .Y(n5152));
MX2X1    g2345(.A(n5152), .B(g1533), .S0(n7366), .Y(n4543));
MX2X1    g2346(.A(n5152), .B(g1534), .S0(n7368), .Y(n4548));
MX2X1    g2347(.A(g1532), .B(n5152), .S0(n7370_1), .Y(n4553));
INVX1    g2348(.A(g1501), .Y(n5143));
MX2X1    g2349(.A(n5143), .B(g1536), .S0(n7366), .Y(n4558));
MX2X1    g2350(.A(n5143), .B(g1537), .S0(n7368), .Y(n4563));
MX2X1    g2351(.A(g1535), .B(n5143), .S0(n7370_1), .Y(n4568));
INVX1    g2352(.A(g1506), .Y(n5134));
MX2X1    g2353(.A(n5134), .B(g1539), .S0(n7366), .Y(n4573));
MX2X1    g2354(.A(n5134), .B(g1540), .S0(n7368), .Y(n4578));
MX2X1    g2355(.A(g1538), .B(n5134), .S0(n7370_1), .Y(n4583));
INVX1    g2356(.A(g1520), .Y(n7400_1));
NOR2X1   g2357(.A(g1557), .B(n7400_1), .Y(n7401));
INVX1    g2358(.A(g1517), .Y(n7402));
INVX1    g2359(.A(g1547), .Y(n7403));
OAI22X1  g2360(.A0(g1558), .A1(n7402), .B0(n7403), .B1(g1556), .Y(n7404));
NOR2X1   g2361(.A(n7404), .B(n7401), .Y(n7405_1));
MX2X1    g2362(.A(n7405_1), .B(g1542), .S0(n7366), .Y(n4588));
MX2X1    g2363(.A(n7405_1), .B(g1543), .S0(n7368), .Y(n4593));
MX2X1    g2364(.A(g1541), .B(n7405_1), .S0(n7370_1), .Y(n4598));
NOR2X1   g2365(.A(g1554), .B(n7400_1), .Y(n7409));
OAI22X1  g2366(.A0(g1555), .A1(n7402), .B0(n7403), .B1(g1553), .Y(n7410_1));
NOR2X1   g2367(.A(n7410_1), .B(n7409), .Y(n7411));
MX2X1    g2368(.A(n7411), .B(g1545), .S0(n7366), .Y(n4603));
MX2X1    g2369(.A(n7411), .B(g1546), .S0(n7368), .Y(n4608));
MX2X1    g2370(.A(g1544), .B(n7411), .S0(n7370_1), .Y(n4613));
NOR4X1   g2371(.A(g1496), .B(g1501), .C(n5134), .D(n5161), .Y(n7415_1));
AND2X1   g2372(.A(n1476), .B(g1520), .Y(n7416));
MX2X1    g2373(.A(g1551), .B(n7415_1), .S0(n7416), .Y(n4618));
AND2X1   g2374(.A(n1476), .B(g1517), .Y(n7418));
MX2X1    g2375(.A(g1552), .B(n7415_1), .S0(n7418), .Y(n4623));
AND2X1   g2376(.A(n1476), .B(g1547), .Y(n7420_1));
MX2X1    g2377(.A(g1550), .B(n7415_1), .S0(n7420_1), .Y(n4628));
MX2X1    g2378(.A(g1554), .B(n5188), .S0(n7416), .Y(n4633));
MX2X1    g2379(.A(g1555), .B(n5188), .S0(n7418), .Y(n4638));
MX2X1    g2380(.A(g1553), .B(n5188), .S0(n7420_1), .Y(n4643));
MX2X1    g2381(.A(g1557), .B(n5197), .S0(n7416), .Y(n4648));
MX2X1    g2382(.A(g1558), .B(n5197), .S0(n7418), .Y(n4653));
MX2X1    g2383(.A(g1556), .B(n5197), .S0(n7420_1), .Y(n4658));
NAND4X1  g2384(.A(g1476), .B(g1481), .C(g1506), .D(g1471), .Y(n7428));
NAND4X1  g2385(.A(g1491), .B(g1496), .C(g1501), .D(g1486), .Y(n7429));
NOR2X1   g2386(.A(n7429), .B(n7428), .Y(n7430_1));
INVX1    g2387(.A(n7430_1), .Y(n7431));
MX2X1    g2388(.A(g1560), .B(n7431), .S0(n7416), .Y(n4663));
MX2X1    g2389(.A(g1561), .B(n7431), .S0(n7418), .Y(n4668));
MX2X1    g2390(.A(g1559), .B(n7431), .S0(n7420_1), .Y(n4673));
NOR2X1   g2391(.A(g1545), .B(n7400_1), .Y(n7435_1));
OAI22X1  g2392(.A0(g1546), .A1(n7402), .B0(n7403), .B1(g1544), .Y(n7436));
OR2X1    g2393(.A(n7436), .B(n7435_1), .Y(n7437));
AND2X1   g2394(.A(n7437), .B(n7411), .Y(n7438));
NOR2X1   g2395(.A(g1551), .B(n7400_1), .Y(n7439));
OAI22X1  g2396(.A0(g1552), .A1(n7402), .B0(n7403), .B1(g1550), .Y(n7440_1));
OAI21X1  g2397(.A0(n7440_1), .A1(n7439), .B0(g1563), .Y(n7441));
NOR2X1   g2398(.A(g1542), .B(n7400_1), .Y(n7442));
OAI22X1  g2399(.A0(g1543), .A1(n7402), .B0(n7403), .B1(g1541), .Y(n7443));
NOR2X1   g2400(.A(n7443), .B(n7442), .Y(n7444));
XOR2X1   g2401(.A(n7444), .B(n7405_1), .Y(n7445_1));
NOR2X1   g2402(.A(g1536), .B(n7400_1), .Y(n7446));
OAI22X1  g2403(.A0(g1537), .A1(n7402), .B0(n7403), .B1(g1535), .Y(n7447));
NOR2X1   g2404(.A(n7447), .B(n7446), .Y(n7448));
XOR2X1   g2405(.A(n7448), .B(n5143), .Y(n7449));
NOR4X1   g2406(.A(n7445_1), .B(n7441), .C(n7438), .D(n7449), .Y(n7450_1));
NOR2X1   g2407(.A(g1530), .B(n7400_1), .Y(n7451));
OAI22X1  g2408(.A0(g1531), .A1(n7402), .B0(n7403), .B1(g1529), .Y(n7452));
NOR2X1   g2409(.A(n7452), .B(n7451), .Y(n7453));
XOR2X1   g2410(.A(n7453), .B(n5161), .Y(n7454));
NOR2X1   g2411(.A(g1527), .B(n7400_1), .Y(n7455_1));
OAI22X1  g2412(.A0(g1528), .A1(n7402), .B0(n7403), .B1(g1526), .Y(n7456));
NOR2X1   g2413(.A(n7456), .B(n7455_1), .Y(n7457));
XOR2X1   g2414(.A(n7457), .B(n5170), .Y(n7458));
NOR2X1   g2415(.A(g1533), .B(n7400_1), .Y(n7459));
OAI22X1  g2416(.A0(g1534), .A1(n7402), .B0(n7403), .B1(g1532), .Y(n7460_1));
NOR2X1   g2417(.A(n7460_1), .B(n7459), .Y(n7461));
XOR2X1   g2418(.A(n7461), .B(n5152), .Y(n7462));
NOR2X1   g2419(.A(g1539), .B(n7400_1), .Y(n7463));
OAI22X1  g2420(.A0(g1540), .A1(n7402), .B0(n7403), .B1(g1538), .Y(n7464));
OAI21X1  g2421(.A0(n7464), .A1(n7463), .B0(n5134), .Y(n7465_1));
OAI21X1  g2422(.A0(n7437), .A1(n7411), .B0(n7465_1), .Y(n7466));
NOR4X1   g2423(.A(n7462), .B(n7458), .C(n7454), .D(n7466), .Y(n7467));
NOR3X1   g2424(.A(n7464), .B(n7463), .C(n5134), .Y(n7468));
NOR2X1   g2425(.A(g1524), .B(n7400_1), .Y(n7469));
OAI22X1  g2426(.A0(g1525), .A1(n7402), .B0(n7403), .B1(g1523), .Y(n7470_1));
NOR2X1   g2427(.A(n7470_1), .B(n7469), .Y(n7471));
XOR2X1   g2428(.A(n7471), .B(n5179), .Y(n7472));
NOR2X1   g2429(.A(g1515), .B(n7400_1), .Y(n7473));
OAI22X1  g2430(.A0(g1516), .A1(n7402), .B0(n7403), .B1(g1514), .Y(n7474));
NOR2X1   g2431(.A(n7474), .B(n7473), .Y(n7475_1));
XOR2X1   g2432(.A(n7475_1), .B(n5188), .Y(n7476));
NOR2X1   g2433(.A(g1512), .B(n7400_1), .Y(n7477));
OAI22X1  g2434(.A0(g1513), .A1(n7402), .B0(n7403), .B1(g1511), .Y(n7478));
NOR2X1   g2435(.A(n7478), .B(n7477), .Y(n7479));
XOR2X1   g2436(.A(n7479), .B(n5197), .Y(n7480_1));
NOR4X1   g2437(.A(n7476), .B(n7472), .C(n7468), .D(n7480_1), .Y(n7481));
NAND3X1  g2438(.A(n7481), .B(n7467), .C(n7450_1), .Y(n7482));
NAND2X1  g2439(.A(g1603), .B(g1520), .Y(n7483));
AOI22X1  g2440(.A0(g1606), .A1(g1517), .B0(g1547), .B1(g1609), .Y(n7484));
AND2X1   g2441(.A(n7484), .B(n7483), .Y(n7485_1));
NOR3X1   g2442(.A(n7485_1), .B(n7404), .C(n7401), .Y(n7486));
OR2X1    g2443(.A(g1557), .B(n7400_1), .Y(n7487));
INVX1    g2444(.A(g1558), .Y(n7488));
INVX1    g2445(.A(g1556), .Y(n7489));
AOI22X1  g2446(.A0(n7488), .A1(g1517), .B0(g1547), .B1(n7489), .Y(n7490_1));
NAND2X1  g2447(.A(n7484), .B(n7483), .Y(n7491));
AOI21X1  g2448(.A0(n7490_1), .A1(n7487), .B0(n7491), .Y(n7492));
NAND2X1  g2449(.A(g1594), .B(g1520), .Y(n7493));
AOI22X1  g2450(.A0(g1597), .A1(g1517), .B0(g1547), .B1(g1600), .Y(n7494));
NAND2X1  g2451(.A(n7494), .B(n7493), .Y(n7495_1));
XOR2X1   g2452(.A(n7495_1), .B(g1501), .Y(n7496));
NOR3X1   g2453(.A(n7496), .B(n7492), .C(n7486), .Y(n7497));
NAND2X1  g2454(.A(g1567), .B(g1520), .Y(n7498));
AOI22X1  g2455(.A0(g1570), .A1(g1517), .B0(g1547), .B1(g1573), .Y(n7499));
NAND2X1  g2456(.A(n7499), .B(n7498), .Y(n7500_1));
XOR2X1   g2457(.A(n7500_1), .B(g1471), .Y(n7501));
NAND2X1  g2458(.A(g1576), .B(g1520), .Y(n7502));
AOI22X1  g2459(.A0(g1579), .A1(g1517), .B0(g1547), .B1(g1582), .Y(n7503));
NAND2X1  g2460(.A(n7503), .B(n7502), .Y(n7504));
XOR2X1   g2461(.A(n7504), .B(g1481), .Y(n7505_1));
NAND2X1  g2462(.A(g1585), .B(g1520), .Y(n7506));
AOI22X1  g2463(.A0(g1588), .A1(g1517), .B0(g1547), .B1(g1591), .Y(n7507));
NAND2X1  g2464(.A(n7507), .B(n7506), .Y(n7508));
XOR2X1   g2465(.A(n7508), .B(g1491), .Y(n7509));
OAI21X1  g2466(.A0(n7509), .A1(n7505_1), .B0(n7501), .Y(n7510_1));
NOR2X1   g2467(.A(n7510_1), .B(n7497), .Y(n7511));
NOR2X1   g2468(.A(n7509), .B(n7496), .Y(n7512));
OAI22X1  g2469(.A0(n7501), .A1(n7505_1), .B0(n7492), .B1(n7486), .Y(n7513));
NOR2X1   g2470(.A(n7513), .B(n7512), .Y(n7514));
XOR2X1   g2471(.A(n7508), .B(n5161), .Y(n7515_1));
NOR2X1   g2472(.A(n7501), .B(n7496), .Y(n7516));
NOR3X1   g2473(.A(n7505_1), .B(n7492), .C(n7486), .Y(n7517));
NOR3X1   g2474(.A(n7517), .B(n7516), .C(n7515_1), .Y(n7518));
NOR3X1   g2475(.A(n7518), .B(n7514), .C(n7511), .Y(n7519_1));
NAND2X1  g2476(.A(g1648), .B(g1520), .Y(n7520));
AOI22X1  g2477(.A0(g1651), .A1(g1517), .B0(g1547), .B1(g1654), .Y(n7521));
AND2X1   g2478(.A(n7521), .B(n7520), .Y(n7522));
NOR3X1   g2479(.A(n7522), .B(n7410_1), .C(n7409), .Y(n7523));
OR2X1    g2480(.A(g1554), .B(n7400_1), .Y(n7524_1));
INVX1    g2481(.A(g1555), .Y(n7525));
INVX1    g2482(.A(g1553), .Y(n7526));
AOI22X1  g2483(.A0(n7525), .A1(g1517), .B0(g1547), .B1(n7526), .Y(n7527));
NAND2X1  g2484(.A(n7521), .B(n7520), .Y(n7528));
AOI21X1  g2485(.A0(n7527), .A1(n7524_1), .B0(n7528), .Y(n7529_1));
NAND2X1  g2486(.A(g1639), .B(g1520), .Y(n7530));
AOI22X1  g2487(.A0(g1642), .A1(g1517), .B0(g1547), .B1(g1645), .Y(n7531));
NAND2X1  g2488(.A(n7531), .B(n7530), .Y(n7532));
XOR2X1   g2489(.A(n7532), .B(g1506), .Y(n7533));
NOR3X1   g2490(.A(n7533), .B(n7529_1), .C(n7523), .Y(n7534_1));
NAND2X1  g2491(.A(g1612), .B(g1520), .Y(n7535));
AOI22X1  g2492(.A0(g1615), .A1(g1517), .B0(g1547), .B1(g1618), .Y(n7536));
NAND2X1  g2493(.A(n7536), .B(n7535), .Y(n7537));
XOR2X1   g2494(.A(n7537), .B(g1476), .Y(n7538));
NAND2X1  g2495(.A(g1621), .B(g1520), .Y(n7539_1));
AOI22X1  g2496(.A0(g1624), .A1(g1517), .B0(g1547), .B1(g1627), .Y(n7540));
NAND2X1  g2497(.A(n7540), .B(n7539_1), .Y(n7541));
XOR2X1   g2498(.A(n7541), .B(g1486), .Y(n7542));
NAND2X1  g2499(.A(g1630), .B(g1520), .Y(n7543));
AOI22X1  g2500(.A0(g1633), .A1(g1517), .B0(g1547), .B1(g1636), .Y(n7544_1));
NAND2X1  g2501(.A(n7544_1), .B(n7543), .Y(n7545));
XOR2X1   g2502(.A(n7545), .B(g1496), .Y(n7546));
OAI21X1  g2503(.A0(n7546), .A1(n7542), .B0(n7538), .Y(n7547));
NOR2X1   g2504(.A(n7547), .B(n7534_1), .Y(n7548));
NOR2X1   g2505(.A(n7546), .B(n7533), .Y(n7549_1));
OAI22X1  g2506(.A0(n7538), .A1(n7542), .B0(n7529_1), .B1(n7523), .Y(n7550));
NOR2X1   g2507(.A(n7550), .B(n7549_1), .Y(n7551));
XOR2X1   g2508(.A(n7545), .B(n5152), .Y(n7552));
NOR2X1   g2509(.A(n7538), .B(n7533), .Y(n7553));
NOR3X1   g2510(.A(n7542), .B(n7529_1), .C(n7523), .Y(n7554_1));
NOR3X1   g2511(.A(n7554_1), .B(n7553), .C(n7552), .Y(n7555));
NOR3X1   g2512(.A(n7555), .B(n7551), .C(n7548), .Y(n7556));
AOI21X1  g2513(.A0(n7556), .A1(n7519_1), .B0(n7441), .Y(n7557));
INVX1    g2514(.A(g1657), .Y(n7558));
NOR2X1   g2515(.A(g1699), .B(n7558), .Y(n7559_1));
INVX1    g2516(.A(g1786), .Y(n7560));
INVX1    g2517(.A(g1782), .Y(n7561));
OAI22X1  g2518(.A0(g1700), .A1(n7560), .B0(n7561), .B1(g1701), .Y(n7562));
NOR2X1   g2519(.A(n7562), .B(n7559_1), .Y(n7563));
NOR2X1   g2520(.A(g1696), .B(n7558), .Y(n7564_1));
OAI22X1  g2521(.A0(g1697), .A1(n7560), .B0(n7561), .B1(g1698), .Y(n7565));
NOR2X1   g2522(.A(n7565), .B(n7564_1), .Y(n7566));
NOR2X1   g2523(.A(g1693), .B(n7558), .Y(n7567));
OAI22X1  g2524(.A0(g1694), .A1(n7560), .B0(n7561), .B1(g1695), .Y(n7568));
NOR2X1   g2525(.A(n7568), .B(n7567), .Y(n7569_1));
INVX1    g2526(.A(n7569_1), .Y(n7570));
NOR2X1   g2527(.A(g1703), .B(n7558), .Y(n7571));
OAI22X1  g2528(.A0(g1704), .A1(n7560), .B0(n7561), .B1(g1702), .Y(n7572));
NOR2X1   g2529(.A(n7572), .B(n7571), .Y(n7573));
INVX1    g2530(.A(n7573), .Y(n7574_1));
NAND4X1  g2531(.A(n7570), .B(n7566), .C(n7563), .D(n7574_1), .Y(n7575));
NOR3X1   g2532(.A(n7575), .B(n7557), .C(n7482), .Y(n7576));
NOR4X1   g2533(.A(n7565), .B(n7564_1), .C(n7563), .D(n7569_1), .Y(n7577));
NAND2X1  g2534(.A(n7577), .B(n7574_1), .Y(n7578_1));
NOR2X1   g2535(.A(n7578_1), .B(n7482), .Y(n7579));
NOR2X1   g2536(.A(g1784), .B(n7558), .Y(n7580));
OAI22X1  g2537(.A0(g1785), .A1(n7560), .B0(n7561), .B1(g1783), .Y(n7581));
NOR2X1   g2538(.A(n7581), .B(n7580), .Y(n7582_1));
INVX1    g2539(.A(g1563), .Y(n7583));
NOR3X1   g2540(.A(n7440_1), .B(n7439), .C(n7583), .Y(n7584));
INVX1    g2541(.A(n7584), .Y(n7585));
OAI22X1  g2542(.A0(n7582_1), .A1(n7482), .B0(n7569_1), .B1(n7585), .Y(n7586));
OR4X1    g2543(.A(n7564_1), .B(n7562), .C(n7559_1), .D(n7565), .Y(n7587_1));
NOR3X1   g2544(.A(n7568), .B(n7567), .C(n7587_1), .Y(n7588));
INVX1    g2545(.A(n7588), .Y(n7589));
INVX1    g2546(.A(n7566), .Y(n7590));
NAND3X1  g2547(.A(n7569_1), .B(n7590), .C(n7563), .Y(n7591));
INVX1    g2548(.A(n7563), .Y(n7592_1));
NOR3X1   g2549(.A(n7570), .B(n7566), .C(n7592_1), .Y(n7593));
NAND4X1  g2550(.A(n7506), .B(n7494), .C(n7493), .D(n7507), .Y(n7594));
OR4X1    g2551(.A(n7545), .B(n7532), .C(n7500_1), .D(n7594), .Y(n7595));
NAND4X1  g2552(.A(n7502), .B(n7484), .C(n7483), .D(n7503), .Y(n7596));
OR4X1    g2553(.A(n7541), .B(n7537), .C(n7528), .D(n7596), .Y(n7597_1));
OR2X1    g2554(.A(n7597_1), .B(n7595), .Y(n7598));
OR2X1    g2555(.A(n7598), .B(n7593), .Y(n7599));
NAND2X1  g2556(.A(n7541), .B(n7528), .Y(n7600));
NAND3X1  g2557(.A(n7537), .B(n7504), .C(n7491), .Y(n7601));
OR4X1    g2558(.A(n7600), .B(n7595), .C(n7591), .D(n7601), .Y(n7602_1));
AOI22X1  g2559(.A0(n7599), .A1(n7602_1), .B0(n7591), .B1(n7589), .Y(n7603));
NOR4X1   g2560(.A(n7586), .B(n7579), .C(n7576), .D(n7603), .Y(n7604));
INVX1    g2561(.A(n7604), .Y(n7605));
NAND2X1  g2562(.A(n7591), .B(n7589), .Y(n7606));
XOR2X1   g2563(.A(n7606), .B(n7500_1), .Y(n7607_1));
NOR3X1   g2564(.A(n7586), .B(n7579), .C(n7576), .Y(n7608));
AOI21X1  g2565(.A0(n7603), .A1(n7608), .B0(n5197), .Y(n7609));
MX2X1    g2566(.A(n7607_1), .B(n7609), .S0(n7605), .Y(n7610));
MX2X1    g2567(.A(g1567), .B(n7610), .S0(g1520), .Y(n4678));
MX2X1    g2568(.A(g1570), .B(n7610), .S0(g1517), .Y(n4683));
MX2X1    g2569(.A(g1573), .B(n7610), .S0(g1547), .Y(n4688));
AND2X1   g2570(.A(n7591), .B(n7500_1), .Y(n7614));
OAI21X1  g2571(.A0(n7591), .A1(n7500_1), .B0(n7606), .Y(n7615));
OR2X1    g2572(.A(n7615), .B(n7614), .Y(n7616));
XOR2X1   g2573(.A(n7616), .B(n7537), .Y(n7617_1));
NAND3X1  g2574(.A(n7603), .B(n7591), .C(n7608), .Y(n7618));
MX2X1    g2575(.A(n5188), .B(n7603), .S0(n7608), .Y(n7619));
AOI22X1  g2576(.A0(n7618), .A1(n7619), .B0(n7617_1), .B1(n7604), .Y(n7620));
MX2X1    g2577(.A(g1612), .B(n7620), .S0(g1520), .Y(n4693));
MX2X1    g2578(.A(g1615), .B(n7620), .S0(g1517), .Y(n4698));
MX2X1    g2579(.A(g1618), .B(n7620), .S0(g1547), .Y(n4703));
XOR2X1   g2580(.A(n7593), .B(n7537), .Y(n7624));
OR2X1    g2581(.A(n7624), .B(n7616), .Y(n7625));
XOR2X1   g2582(.A(n7625), .B(n7504), .Y(n7626));
MX2X1    g2583(.A(n5179), .B(n7603), .S0(n7608), .Y(n7627_1));
AOI22X1  g2584(.A0(n7626), .A1(n7604), .B0(n7618), .B1(n7627_1), .Y(n7628));
MX2X1    g2585(.A(g1576), .B(n7628), .S0(g1520), .Y(n4708));
MX2X1    g2586(.A(g1579), .B(n7628), .S0(g1517), .Y(n4713));
MX2X1    g2587(.A(g1582), .B(n7628), .S0(g1547), .Y(n4718));
XOR2X1   g2588(.A(n7593), .B(n7504), .Y(n7632_1));
OR4X1    g2589(.A(n7624), .B(n7615), .C(n7614), .D(n7632_1), .Y(n7633));
XOR2X1   g2590(.A(n7633), .B(n7541), .Y(n7634));
MX2X1    g2591(.A(n5170), .B(n7603), .S0(n7608), .Y(n7635));
AOI22X1  g2592(.A0(n7634), .A1(n7604), .B0(n7618), .B1(n7635), .Y(n7636));
MX2X1    g2593(.A(g1621), .B(n7636), .S0(g1520), .Y(n4723));
MX2X1    g2594(.A(g1624), .B(n7636), .S0(g1517), .Y(n4728));
MX2X1    g2595(.A(g1627), .B(n7636), .S0(g1547), .Y(n4733));
XOR2X1   g2596(.A(n7593), .B(n7541), .Y(n7640));
OR2X1    g2597(.A(n7640), .B(n7632_1), .Y(n7641));
NOR4X1   g2598(.A(n7624), .B(n7615), .C(n7614), .D(n7641), .Y(n7642_1));
XOR2X1   g2599(.A(n7642_1), .B(n7508), .Y(n7643));
AOI21X1  g2600(.A0(n7603), .A1(n7608), .B0(n5161), .Y(n7644));
MX2X1    g2601(.A(n7643), .B(n7644), .S0(n7605), .Y(n7645));
MX2X1    g2602(.A(g1585), .B(n7645), .S0(g1520), .Y(n4738));
MX2X1    g2603(.A(g1588), .B(n7645), .S0(g1517), .Y(n4743));
MX2X1    g2604(.A(g1591), .B(n7645), .S0(g1547), .Y(n4748));
XOR2X1   g2605(.A(n7591), .B(n7508), .Y(n7649));
AND2X1   g2606(.A(n7649), .B(n7642_1), .Y(n7650));
XOR2X1   g2607(.A(n7650), .B(n7545), .Y(n7651));
AOI21X1  g2608(.A0(n7603), .A1(n7608), .B0(n5152), .Y(n7652_1));
MX2X1    g2609(.A(n7651), .B(n7652_1), .S0(n7605), .Y(n7653));
MX2X1    g2610(.A(g1630), .B(n7653), .S0(g1520), .Y(n4753));
MX2X1    g2611(.A(g1633), .B(n7653), .S0(g1517), .Y(n4758));
MX2X1    g2612(.A(g1636), .B(n7653), .S0(g1547), .Y(n4763));
XOR2X1   g2613(.A(n7591), .B(n7545), .Y(n7657_1));
NAND2X1  g2614(.A(n7657_1), .B(n7649), .Y(n7658));
NOR4X1   g2615(.A(n7641), .B(n7624), .C(n7616), .D(n7658), .Y(n7659));
XOR2X1   g2616(.A(n7659), .B(n7495_1), .Y(n7660));
AOI21X1  g2617(.A0(n7603), .A1(n7608), .B0(n5143), .Y(n7661));
MX2X1    g2618(.A(n7660), .B(n7661), .S0(n7605), .Y(n7662_1));
MX2X1    g2619(.A(g1594), .B(n7662_1), .S0(g1520), .Y(n4768));
MX2X1    g2620(.A(g1597), .B(n7662_1), .S0(g1517), .Y(n4773));
MX2X1    g2621(.A(g1600), .B(n7662_1), .S0(g1547), .Y(n4778));
XOR2X1   g2622(.A(n7591), .B(n7495_1), .Y(n7666));
AND2X1   g2623(.A(n7666), .B(n7659), .Y(n7667_1));
XOR2X1   g2624(.A(n7667_1), .B(n7532), .Y(n7668));
AOI21X1  g2625(.A0(n7603), .A1(n7608), .B0(n5134), .Y(n7669));
MX2X1    g2626(.A(n7668), .B(n7669), .S0(n7605), .Y(n7670));
MX2X1    g2627(.A(g1639), .B(n7670), .S0(g1520), .Y(n4783));
MX2X1    g2628(.A(g1642), .B(n7670), .S0(g1517), .Y(n4788));
MX2X1    g2629(.A(g1645), .B(n7670), .S0(g1547), .Y(n4793));
XOR2X1   g2630(.A(n7591), .B(n7532), .Y(n7674));
NAND4X1  g2631(.A(n7666), .B(n7657_1), .C(n7649), .D(n7674), .Y(n7675));
OR4X1    g2632(.A(n7641), .B(n7624), .C(n7616), .D(n7675), .Y(n7676));
XOR2X1   g2633(.A(n7676), .B(n7491), .Y(n7677_1));
MX2X1    g2634(.A(n7405_1), .B(n7603), .S0(n7608), .Y(n7678));
AOI22X1  g2635(.A0(n7677_1), .A1(n7604), .B0(n7618), .B1(n7678), .Y(n7679));
MX2X1    g2636(.A(g1603), .B(n7679), .S0(g1520), .Y(n4798));
MX2X1    g2637(.A(g1606), .B(n7679), .S0(g1517), .Y(n4803));
MX2X1    g2638(.A(g1609), .B(n7679), .S0(g1547), .Y(n4808));
XOR2X1   g2639(.A(n7593), .B(n7491), .Y(n7683));
OR2X1    g2640(.A(n7683), .B(n7676), .Y(n7684));
XOR2X1   g2641(.A(n7684), .B(n7528), .Y(n7685));
MX2X1    g2642(.A(n7411), .B(n7603), .S0(n7608), .Y(n7686));
AOI22X1  g2643(.A0(n7685), .A1(n7604), .B0(n7618), .B1(n7686), .Y(n7687_1));
MX2X1    g2644(.A(g1648), .B(n7687_1), .S0(g1520), .Y(n4813));
MX2X1    g2645(.A(g1651), .B(n7687_1), .S0(g1517), .Y(n4818));
MX2X1    g2646(.A(g1654), .B(n7687_1), .S0(g1547), .Y(n4823));
INVX1    g2647(.A(g1466), .Y(n7691));
NOR2X1   g2648(.A(n5399), .B(n7403), .Y(n7692_1));
XOR2X1   g2649(.A(n7692_1), .B(n7691), .Y(n7693));
AOI21X1  g2650(.A0(n7370_1), .A1(n5399), .B0(n7693), .Y(n4828));
INVX1    g2651(.A(g1462), .Y(n7695));
NOR3X1   g2652(.A(n5399), .B(n7691), .C(n7403), .Y(n7696));
XOR2X1   g2653(.A(n7696), .B(n7695), .Y(n7697_1));
AOI21X1  g2654(.A0(n7370_1), .A1(n5399), .B0(n7697_1), .Y(n4833));
INVX1    g2655(.A(g1457), .Y(n7699));
NOR4X1   g2656(.A(n7695), .B(n7691), .C(n7403), .D(n5399), .Y(n7700));
XOR2X1   g2657(.A(n7700), .B(n7699), .Y(n7701));
AOI21X1  g2658(.A0(n7370_1), .A1(n5399), .B0(n7701), .Y(n4838));
NAND2X1  g2659(.A(n7700), .B(g1457), .Y(n7703));
XOR2X1   g2660(.A(n7703), .B(g1453), .Y(n7704));
AOI21X1  g2661(.A0(n7370_1), .A1(n5399), .B0(n7704), .Y(n4843));
NAND3X1  g2662(.A(n7700), .B(g1453), .C(g1457), .Y(n7706));
XOR2X1   g2663(.A(n7706), .B(g1448), .Y(n7707_1));
AOI21X1  g2664(.A0(n7370_1), .A1(n5399), .B0(n7707_1), .Y(n4848));
INVX1    g2665(.A(g1453), .Y(n7709));
INVX1    g2666(.A(g1448), .Y(n7710));
OR4X1    g2667(.A(g1444), .B(n7710), .C(n7709), .D(n7703), .Y(n7711));
OAI21X1  g2668(.A0(n7706), .A1(n7710), .B0(g1444), .Y(n7712_1));
AOI22X1  g2669(.A0(n7711), .A1(n7712_1), .B0(n7370_1), .B1(n5399), .Y(n4853));
INVX1    g2670(.A(g1444), .Y(n7714));
OR4X1    g2671(.A(n7714), .B(n7710), .C(n7709), .D(n7703), .Y(n7715));
XOR2X1   g2672(.A(n7715), .B(g1439), .Y(n7716));
AOI21X1  g2673(.A0(n7370_1), .A1(n5399), .B0(n7716), .Y(n4858));
INVX1    g2674(.A(g1435), .Y(n7718));
INVX1    g2675(.A(g1439), .Y(n7719));
NOR4X1   g2676(.A(n7719), .B(n7714), .C(n7710), .D(n7706), .Y(n7720));
XOR2X1   g2677(.A(n7720), .B(n7718), .Y(n7721));
AOI21X1  g2678(.A0(n7370_1), .A1(n5399), .B0(n7721), .Y(n4863));
INVX1    g2679(.A(g1430), .Y(n7723));
AND2X1   g2680(.A(n7720), .B(g1435), .Y(n7724));
XOR2X1   g2681(.A(n7724), .B(n7723), .Y(n7725));
AOI21X1  g2682(.A0(n7370_1), .A1(n5399), .B0(n7725), .Y(n4868));
INVX1    g2683(.A(g1426), .Y(n7727_1));
NOR4X1   g2684(.A(n7723), .B(n7718), .C(n7719), .D(n7715), .Y(n7728));
XOR2X1   g2685(.A(n7728), .B(n7727_1), .Y(n7729));
AOI21X1  g2686(.A0(n7370_1), .A1(n5399), .B0(n7729), .Y(n4873));
NOR2X1   g2687(.A(g1765), .B(n7558), .Y(n7731));
OAI22X1  g2688(.A0(g1754), .A1(n7560), .B0(n7561), .B1(g1757), .Y(n7732_1));
NOR2X1   g2689(.A(g1750), .B(n7558), .Y(n7733));
OAI22X1  g2690(.A0(g1739), .A1(n7560), .B0(n7561), .B1(g1742), .Y(n7734));
NOR2X1   g2691(.A(n7734), .B(n7733), .Y(n7735));
OR4X1    g2692(.A(n7732_1), .B(n7731), .C(g3229), .D(n7735), .Y(n7736));
NOR2X1   g2693(.A(g1779), .B(n7558), .Y(n7737_1));
OAI22X1  g2694(.A0(g1769), .A1(n7560), .B0(n7561), .B1(g1772), .Y(n7738));
NOR2X1   g2695(.A(n7738), .B(n7737_1), .Y(n7739));
OAI21X1  g2696(.A0(n7739), .A1(n5718), .B0(n7736), .Y(n7740));
INVX1    g2697(.A(n7735), .Y(n5255));
INVX1    g2698(.A(n7739), .Y(n5265));
NOR2X1   g2699(.A(g1735), .B(n7558), .Y(n7743));
OAI22X1  g2700(.A0(g1724), .A1(n7560), .B0(n7561), .B1(g1727), .Y(n7744));
NOR2X1   g2701(.A(n7744), .B(n7743), .Y(n7745));
NOR4X1   g2702(.A(n5265), .B(n5255), .C(n5718), .D(n7745), .Y(n7746));
NOR4X1   g2703(.A(n7738), .B(n7737_1), .C(g3229), .D(n7745), .Y(n7747_1));
NOR2X1   g2704(.A(n7732_1), .B(n7731), .Y(n7748));
NOR3X1   g2705(.A(n7745), .B(n7748), .C(n5718), .Y(n7749));
NOR4X1   g2706(.A(n7747_1), .B(n7746), .C(n7740), .D(n7749), .Y(n7750));
NOR4X1   g2707(.A(n7567), .B(n7566), .C(n7563), .D(n7568), .Y(n7751));
AOI21X1  g2708(.A0(n7589), .A1(n5399), .B0(n7751), .Y(n5270));
AND2X1   g2709(.A(n5270), .B(g1657), .Y(n7753));
MX2X1    g2710(.A(g1735), .B(n7750), .S0(n7753), .Y(n4909));
AND2X1   g2711(.A(n5270), .B(g1786), .Y(n7755));
MX2X1    g2712(.A(g1724), .B(n7750), .S0(n7755), .Y(n4914));
AND2X1   g2713(.A(n5270), .B(g1782), .Y(n7757_1));
MX2X1    g2714(.A(g1727), .B(n7750), .S0(n7757_1), .Y(n4919));
NOR4X1   g2715(.A(n7743), .B(n7748), .C(g3229), .D(n7744), .Y(n7759));
NOR3X1   g2716(.A(n7735), .B(n7732_1), .C(n7731), .Y(n7760));
NOR3X1   g2717(.A(n7760), .B(n7759), .C(n7749), .Y(n7761));
MX2X1    g2718(.A(g1750), .B(n7761), .S0(n7753), .Y(n4924));
MX2X1    g2719(.A(g1739), .B(n7761), .S0(n7755), .Y(n4929));
MX2X1    g2720(.A(g1742), .B(n7761), .S0(n7757_1), .Y(n4934));
NOR4X1   g2721(.A(n7743), .B(n7735), .C(n5718), .D(n7744), .Y(n7765));
NOR3X1   g2722(.A(n7745), .B(n7735), .C(g3229), .Y(n7766));
INVX1    g2723(.A(n7745), .Y(n5250));
NOR4X1   g2724(.A(n5265), .B(n5255), .C(g3229), .D(n5250), .Y(n7768));
NOR4X1   g2725(.A(n7766), .B(n7765), .C(n7746), .D(n7768), .Y(n7769));
MX2X1    g2726(.A(g1765), .B(n7769), .S0(n7753), .Y(n4939));
MX2X1    g2727(.A(g1754), .B(n7769), .S0(n7755), .Y(n4944));
MX2X1    g2728(.A(g1757), .B(n7769), .S0(n7757_1), .Y(n4949));
NOR2X1   g2729(.A(n7745), .B(g3229), .Y(n7773));
NOR3X1   g2730(.A(n7744), .B(n7743), .C(n5718), .Y(n7774));
NOR4X1   g2731(.A(n7733), .B(n7732_1), .C(n7731), .D(n7734), .Y(n7775));
OAI21X1  g2732(.A0(n7774), .A1(n7773), .B0(n7775), .Y(n7776));
MX2X1    g2733(.A(g1779), .B(n7776), .S0(n7753), .Y(n4954));
MX2X1    g2734(.A(g1769), .B(n7776), .S0(n7755), .Y(n4959));
MX2X1    g2735(.A(g1772), .B(n7776), .S0(n7757_1), .Y(n4964));
NAND2X1  g2736(.A(g1789), .B(g1657), .Y(n7780));
AOI22X1  g2737(.A0(g1792), .A1(g1786), .B0(g1782), .B1(g1795), .Y(n7781));
AND2X1   g2738(.A(n7781), .B(n7780), .Y(n7782_1));
INVX1    g2739(.A(n7782_1), .Y(n7783));
OR4X1    g2740(.A(n7431), .B(n7411), .C(n7405_1), .D(n7584), .Y(n7784));
NAND2X1  g2741(.A(g1798), .B(g1657), .Y(n7785));
AOI22X1  g2742(.A0(g1801), .A1(g1786), .B0(g1782), .B1(g1804), .Y(n7786));
AND2X1   g2743(.A(n7786), .B(n7785), .Y(n7787_1));
AND2X1   g2744(.A(n7787_1), .B(n7784), .Y(n7788));
NOR3X1   g2745(.A(n7431), .B(n7411), .C(n7405_1), .Y(n7789));
INVX1    g2746(.A(n7789), .Y(n7790));
OAI21X1  g2747(.A0(n7787_1), .A1(n7790), .B0(n7782_1), .Y(n7791));
INVX1    g2748(.A(n7787_1), .Y(n5215));
NOR2X1   g2749(.A(g1808), .B(n7558), .Y(n7793));
OAI22X1  g2750(.A0(g1809), .A1(n7560), .B0(n7561), .B1(g1807), .Y(n7794));
NOR2X1   g2751(.A(n7794), .B(n7793), .Y(n7795));
INVX1    g2752(.A(n7795), .Y(n7796));
NOR4X1   g2753(.A(n5215), .B(n7790), .C(n7584), .D(n7796), .Y(n7797_1));
NAND2X1  g2754(.A(n7795), .B(n5215), .Y(n7798));
OAI21X1  g2755(.A0(n7798), .A1(n7789), .B0(n7783), .Y(n7799));
OAI22X1  g2756(.A0(n7797_1), .A1(n7799), .B0(n7791), .B1(n7788), .Y(n7800));
AND2X1   g2757(.A(n7800), .B(g1690), .Y(n7801));
XOR2X1   g2758(.A(n7801), .B(n7783), .Y(n7802_1));
MX2X1    g2759(.A(g1789), .B(n7802_1), .S0(g1657), .Y(n4969));
MX2X1    g2760(.A(g1792), .B(n7802_1), .S0(g1786), .Y(n4974));
MX2X1    g2761(.A(g1795), .B(n7802_1), .S0(g1782), .Y(n4979));
INVX1    g2762(.A(g1690), .Y(n7806));
NAND4X1  g2763(.A(n7787_1), .B(n7789), .C(n7584), .D(n7782_1), .Y(n7807_1));
OAI21X1  g2764(.A0(n7796), .A1(n7584), .B0(n7789), .Y(n7808));
NAND2X1  g2765(.A(n7808), .B(n7787_1), .Y(n7809));
OAI21X1  g2766(.A0(n7795), .A1(n7789), .B0(n5215), .Y(n7810));
NAND3X1  g2767(.A(n7810), .B(n7809), .C(n7783), .Y(n7811));
AOI21X1  g2768(.A0(n7811), .A1(n7807_1), .B0(n7806), .Y(n7812_1));
XOR2X1   g2769(.A(n7812_1), .B(n5215), .Y(n7813));
MX2X1    g2770(.A(g1798), .B(n7813), .S0(g1657), .Y(n4984));
MX2X1    g2771(.A(g1801), .B(n7813), .S0(g1786), .Y(n4989));
MX2X1    g2772(.A(g1804), .B(n7813), .S0(g1782), .Y(n4994));
MX2X1    g2773(.A(n7784), .B(n7789), .S0(n5215), .Y(n7817_1));
OR4X1    g2774(.A(n7796), .B(n7782_1), .C(n7806), .D(n7817_1), .Y(n7818));
NAND3X1  g2775(.A(n7781), .B(n7780), .C(g1690), .Y(n7819));
OAI21X1  g2776(.A0(n7819), .A1(n7817_1), .B0(n7818), .Y(n7820));
AND2X1   g2777(.A(n7820), .B(g1657), .Y(n7821));
MX2X1    g2778(.A(g1808), .B(n7818), .S0(n7821), .Y(n4999));
AND2X1   g2779(.A(n7820), .B(g1786), .Y(n7823));
MX2X1    g2780(.A(g1809), .B(n7818), .S0(n7823), .Y(n5004));
AND2X1   g2781(.A(n7820), .B(g1782), .Y(n7825));
MX2X1    g2782(.A(g1807), .B(n7818), .S0(n7825), .Y(n5009));
NAND2X1  g2783(.A(g1810), .B(g1657), .Y(n7827_1));
AOI22X1  g2784(.A0(g1813), .A1(g1786), .B0(g1782), .B1(g1816), .Y(n7828));
NAND2X1  g2785(.A(n7828), .B(n7827_1), .Y(n7829));
OR2X1    g2786(.A(g1560), .B(n7400_1), .Y(n7830));
INVX1    g2787(.A(g1561), .Y(n7831));
INVX1    g2788(.A(g1559), .Y(n7832_1));
AOI22X1  g2789(.A0(n7831), .A1(g1517), .B0(g1547), .B1(n7832_1), .Y(n7833));
AOI21X1  g2790(.A0(n7833), .A1(n7830), .B0(n7431), .Y(n7834));
MX2X1    g2791(.A(n7829), .B(n7834), .S0(g1690), .Y(n7835));
MX2X1    g2792(.A(g1810), .B(n7835), .S0(g1657), .Y(n5014));
MX2X1    g2793(.A(g1813), .B(n7835), .S0(g1786), .Y(n5019));
MX2X1    g2794(.A(g1816), .B(n7835), .S0(g1782), .Y(n5024));
NAND2X1  g2795(.A(g1819), .B(g1657), .Y(n7839));
AOI22X1  g2796(.A0(g1822), .A1(g1786), .B0(g1782), .B1(g1825), .Y(n7840));
AND2X1   g2797(.A(n7840), .B(n7839), .Y(n7841));
INVX1    g2798(.A(n7841), .Y(n7842_1));
NOR2X1   g2799(.A(n7841), .B(n7829), .Y(n7843));
INVX1    g2800(.A(n7843), .Y(n7844));
AND2X1   g2801(.A(n7841), .B(n7829), .Y(n7845));
INVX1    g2802(.A(n7845), .Y(n7846));
MX2X1    g2803(.A(n7844), .B(n7846), .S0(n7834), .Y(n7847_1));
NOR2X1   g2804(.A(g1829), .B(n7558), .Y(n7848));
OAI22X1  g2805(.A0(g1830), .A1(n7560), .B0(n7561), .B1(g1828), .Y(n7849));
OAI21X1  g2806(.A0(n7849), .A1(n7848), .B0(g1690), .Y(n7850));
NOR2X1   g2807(.A(n7850), .B(n7847_1), .Y(n7851));
XOR2X1   g2808(.A(n7851), .B(n7842_1), .Y(n7852_1));
MX2X1    g2809(.A(g1819), .B(n7852_1), .S0(g1657), .Y(n5029));
MX2X1    g2810(.A(g1822), .B(n7852_1), .S0(g1786), .Y(n5034));
MX2X1    g2811(.A(g1825), .B(n7852_1), .S0(g1782), .Y(n5039));
NOR4X1   g2812(.A(n7848), .B(n7847_1), .C(n7806), .D(n7849), .Y(n7856));
INVX1    g2813(.A(n7856), .Y(n7857_1));
NOR2X1   g2814(.A(n7842_1), .B(n7829), .Y(n7858));
AOI22X1  g2815(.A0(n7839), .A1(n7840), .B0(n7828), .B1(n7827_1), .Y(n7859));
MX2X1    g2816(.A(n7859), .B(n7858), .S0(n7834), .Y(n7860));
AOI21X1  g2817(.A0(n7860), .A1(g1690), .B0(n7856), .Y(n7861));
NOR2X1   g2818(.A(n7861), .B(n7558), .Y(n7862_1));
MX2X1    g2819(.A(g1829), .B(n7857_1), .S0(n7862_1), .Y(n5044));
NOR2X1   g2820(.A(n7861), .B(n7560), .Y(n7864));
MX2X1    g2821(.A(g1830), .B(n7857_1), .S0(n7864), .Y(n5049));
NOR2X1   g2822(.A(n7861), .B(n7561), .Y(n7866));
MX2X1    g2823(.A(g1828), .B(n7857_1), .S0(n7866), .Y(n5054));
OAI21X1  g2824(.A0(n7590), .A1(n7563), .B0(n7557), .Y(n7868));
AOI21X1  g2825(.A0(n7868), .A1(n7570), .B0(n7593), .Y(n7869));
OR2X1    g2826(.A(n7582_1), .B(n7482), .Y(n7870));
OAI21X1  g2827(.A0(n7869), .A1(n7569_1), .B0(n7870), .Y(n7871));
AOI21X1  g2828(.A0(n7869), .A1(n7569_1), .B0(n7871), .Y(n7872_1));
MX2X1    g2829(.A(g1693), .B(n7872_1), .S0(g1657), .Y(n5059));
MX2X1    g2830(.A(g1694), .B(n7872_1), .S0(g1786), .Y(n5064));
MX2X1    g2831(.A(g1695), .B(n7872_1), .S0(g1782), .Y(n5069));
INVX1    g2832(.A(n7441), .Y(n7876));
NAND3X1  g2833(.A(n7552), .B(n7515_1), .C(n7497), .Y(n7877_1));
NOR2X1   g2834(.A(n7505_1), .B(n7501), .Y(n7878));
NAND2X1  g2835(.A(n7534_1), .B(n7878), .Y(n7879));
OR4X1    g2836(.A(n7877_1), .B(n7542), .C(n7538), .D(n7879), .Y(n7880));
NAND2X1  g2837(.A(n7880), .B(n7876), .Y(n7881));
NOR4X1   g2838(.A(n7573), .B(n7557), .C(n7482), .D(n7881), .Y(n7882_1));
NOR2X1   g2839(.A(n7556), .B(n7441), .Y(n7883));
OAI21X1  g2840(.A0(n7880), .A1(n7441), .B0(n7585), .Y(n7884));
OR4X1    g2841(.A(n7562), .B(n7559_1), .C(n7883), .D(n7884), .Y(n7885));
NAND4X1  g2842(.A(n7481), .B(n7467), .C(n7450_1), .D(n7574_1), .Y(n7886));
NOR2X1   g2843(.A(n7584), .B(n7563), .Y(n7887_1));
AOI21X1  g2844(.A0(n7887_1), .A1(n7886), .B0(n7590), .Y(n7888));
OAI21X1  g2845(.A0(n7885), .A1(n7882_1), .B0(n7888), .Y(n7889));
OR2X1    g2846(.A(n7510_1), .B(n7497), .Y(n7890));
OR2X1    g2847(.A(n7513), .B(n7512), .Y(n7891));
OR2X1    g2848(.A(n7501), .B(n7496), .Y(n7892_1));
NAND3X1  g2849(.A(n7491), .B(n7490_1), .C(n7487), .Y(n7893));
OAI21X1  g2850(.A0(n7404), .A1(n7401), .B0(n7485_1), .Y(n7894));
XOR2X1   g2851(.A(n7504), .B(n5179), .Y(n7895));
NAND3X1  g2852(.A(n7895), .B(n7894), .C(n7893), .Y(n7896));
NAND3X1  g2853(.A(n7896), .B(n7892_1), .C(n7509), .Y(n7897_1));
NAND3X1  g2854(.A(n7897_1), .B(n7891), .C(n7890), .Y(n7898));
AOI21X1  g2855(.A0(n7898), .A1(n7876), .B0(n7592_1), .Y(n7899));
OAI21X1  g2856(.A0(n7881), .A1(n7883), .B0(n7899), .Y(n7900));
AOI21X1  g2857(.A0(n7898), .A1(n7876), .B0(n7563), .Y(n7901));
NOR2X1   g2858(.A(n7901), .B(n7566), .Y(n7902_1));
AOI21X1  g2859(.A0(n7902_1), .A1(n7900), .B0(n7569_1), .Y(n7903));
AOI22X1  g2860(.A0(n7889), .A1(n7903), .B0(n7569_1), .B1(n7587_1), .Y(n7904));
OAI21X1  g2861(.A0(n7904), .A1(n7566), .B0(n7870), .Y(n7905));
AOI21X1  g2862(.A0(n7904), .A1(n7566), .B0(n7905), .Y(n7906));
MX2X1    g2863(.A(g1696), .B(n7906), .S0(g1657), .Y(n5074));
MX2X1    g2864(.A(g1697), .B(n7906), .S0(g1786), .Y(n5079));
MX2X1    g2865(.A(g1698), .B(n7906), .S0(g1782), .Y(n5084));
AOI21X1  g2866(.A0(n7884), .A1(n7563), .B0(n7566), .Y(n7911));
OAI21X1  g2867(.A0(n7881), .A1(n7563), .B0(n7911), .Y(n7912_1));
NOR2X1   g2868(.A(n7519_1), .B(n7441), .Y(n7913));
OR4X1    g2869(.A(n7883), .B(n7913), .C(n7806), .D(n7592_1), .Y(n7914));
AOI21X1  g2870(.A0(n7914), .A1(n7566), .B0(n7569_1), .Y(n7915));
AOI22X1  g2871(.A0(n7912_1), .A1(n7915), .B0(n7569_1), .B1(n7563), .Y(n7916));
XOR2X1   g2872(.A(n7916), .B(n7592_1), .Y(n7917_1));
AND2X1   g2873(.A(n7917_1), .B(n7870), .Y(n7918));
MX2X1    g2874(.A(g1699), .B(n7918), .S0(g1657), .Y(n5089));
MX2X1    g2875(.A(g1700), .B(n7918), .S0(g1786), .Y(n5094));
MX2X1    g2876(.A(g1701), .B(n7918), .S0(g1782), .Y(n5099));
NOR3X1   g2877(.A(n7592_1), .B(n7557), .C(n7482), .Y(n7922_1));
NOR3X1   g2878(.A(n7590), .B(n7563), .C(n7482), .Y(n7923));
OAI21X1  g2879(.A0(n7923), .A1(n7922_1), .B0(n7570), .Y(n7924));
MX2X1    g2880(.A(n7881), .B(n7806), .S0(n7577), .Y(n7925));
NOR2X1   g2881(.A(n7925), .B(n7558), .Y(n7926));
MX2X1    g2882(.A(g1703), .B(n7924), .S0(n7926), .Y(n5104));
NOR2X1   g2883(.A(n7925), .B(n7560), .Y(n7928));
MX2X1    g2884(.A(g1704), .B(n7924), .S0(n7928), .Y(n5109));
NOR2X1   g2885(.A(n7925), .B(n7561), .Y(n7930));
MX2X1    g2886(.A(g1702), .B(n7924), .S0(n7930), .Y(n5114));
NAND4X1  g2887(.A(n7481), .B(n7467), .C(n7450_1), .D(n7582_1), .Y(n7932_1));
AND2X1   g2888(.A(g1690), .B(g1657), .Y(n7933));
MX2X1    g2889(.A(g1784), .B(n7932_1), .S0(n7933), .Y(n5119));
AND2X1   g2890(.A(g1690), .B(g1786), .Y(n7935));
MX2X1    g2891(.A(g1785), .B(n7932_1), .S0(n7935), .Y(n5124));
AND2X1   g2892(.A(g1690), .B(g1782), .Y(n7937_1));
MX2X1    g2893(.A(g1783), .B(n7932_1), .S0(n7937_1), .Y(n5129));
INVX1    g2894(.A(g1680), .Y(n7939));
NAND2X1  g2895(.A(n3519), .B(g1786), .Y(n7940));
AOI21X1  g2896(.A0(g1686), .A1(n7560), .B0(n7939), .Y(n7941));
AOI22X1  g2897(.A0(n7940), .A1(n7941), .B0(g1679), .B1(n7939), .Y(n5220));
NAND2X1  g2898(.A(n3524), .B(g1786), .Y(n7943));
AOI21X1  g2899(.A0(g1689), .A1(n7560), .B0(n7939), .Y(n7944));
NOR2X1   g2900(.A(g1681), .B(g1680), .Y(n7945));
AOI21X1  g2901(.A0(n7944), .A1(n7943), .B0(n7945), .Y(n5225));
NAND2X1  g2902(.A(n3529), .B(g1786), .Y(n7947_1));
AOI21X1  g2903(.A0(g1678), .A1(n7560), .B0(n7939), .Y(n7948));
NOR2X1   g2904(.A(g1682), .B(g1680), .Y(n7949));
AOI21X1  g2905(.A0(n7948), .A1(n7947_1), .B0(n7949), .Y(n5230));
NAND2X1  g2906(.A(n3534), .B(g1786), .Y(n7951));
AOI21X1  g2907(.A0(g1677), .A1(n7560), .B0(n7939), .Y(n7952_1));
NOR2X1   g2908(.A(g1683), .B(g1680), .Y(n7953));
AOI21X1  g2909(.A0(n7952_1), .A1(n7951), .B0(n7953), .Y(n5235));
NAND2X1  g2910(.A(n3539), .B(g1786), .Y(n7955));
AOI21X1  g2911(.A0(g1676), .A1(n7560), .B0(n7939), .Y(n7956));
NOR2X1   g2912(.A(g1684), .B(g1680), .Y(n7957_1));
AOI21X1  g2913(.A0(n7956), .A1(n7955), .B0(n7957_1), .Y(n5240));
NAND2X1  g2914(.A(n3544), .B(g1786), .Y(n7959));
AOI21X1  g2915(.A0(g1675), .A1(n7560), .B0(n7939), .Y(n7960));
NOR2X1   g2916(.A(g1685), .B(g1680), .Y(n7961));
AOI21X1  g2917(.A0(n7960), .A1(n7959), .B0(n7961), .Y(n5245));
INVX1    g2918(.A(n7748), .Y(n5260));
NOR3X1   g2919(.A(n7598), .B(n7570), .C(n7587_1), .Y(n7964));
XOR2X1   g2920(.A(n7508), .B(n7710), .Y(n7965));
XOR2X1   g2921(.A(n7532), .B(n7718), .Y(n7966));
XOR2X1   g2922(.A(n7545), .B(n7714), .Y(n7967_1));
NAND3X1  g2923(.A(n7967_1), .B(n7966), .C(n7965), .Y(n7968));
XOR2X1   g2924(.A(n7528), .B(n7727_1), .Y(n7969));
XOR2X1   g2925(.A(n7537), .B(n7695), .Y(n7970));
XOR2X1   g2926(.A(n7495_1), .B(n7719), .Y(n7971));
XOR2X1   g2927(.A(n7491), .B(n7723), .Y(n7972_1));
NAND4X1  g2928(.A(n7971), .B(n7970), .C(n7969), .D(n7972_1), .Y(n7973));
XOR2X1   g2929(.A(n7541), .B(g1453), .Y(n7974));
XOR2X1   g2930(.A(n7504), .B(g1457), .Y(n7975));
XOR2X1   g2931(.A(n7500_1), .B(g1466), .Y(n7976));
OR2X1    g2932(.A(n7976), .B(n7975), .Y(n7977_1));
OR4X1    g2933(.A(n7974), .B(n7751), .C(n5399), .D(n7977_1), .Y(n7978));
NOR3X1   g2934(.A(n7978), .B(n7973), .C(n7968), .Y(n7979));
OAI21X1  g2935(.A0(n7979), .A1(n7964), .B0(n5270), .Y(n5275));
MX2X1    g2936(.A(g1934), .B(n5982), .S0(g1930), .Y(n5414));
INVX1    g2937(.A(g1930), .Y(n7982_1));
INVX1    g2938(.A(g1934), .Y(n7983));
MX2X1    g2939(.A(n7983), .B(g1937), .S0(n7982_1), .Y(n5419));
MX2X1    g2940(.A(g1890), .B(g1937), .S0(g1930), .Y(n5424));
NAND2X1  g2941(.A(g1949), .B(g1925), .Y(n7986));
AOI22X1  g2942(.A0(g1951), .A1(g1931), .B0(g1930), .B1(g1953), .Y(n7987_1));
AND2X1   g2943(.A(n7987_1), .B(n7986), .Y(n5429));
MX2X1    g2944(.A(g1867), .B(n7842_1), .S0(g1855), .Y(n5509));
MX2X1    g2945(.A(g1868), .B(n7842_1), .S0(g1862), .Y(n5514));
MX2X1    g2946(.A(g1869), .B(n7842_1), .S0(g1866), .Y(n5519));
MX2X1    g2947(.A(g1836), .B(n7751), .S0(g1855), .Y(n5524));
MX2X1    g2948(.A(g1839), .B(n7751), .S0(g1862), .Y(n5529));
MX2X1    g2949(.A(g1842), .B(n7751), .S0(g1866), .Y(n5534));
MX2X1    g2950(.A(g1858), .B(n7577), .S0(g1855), .Y(n5539));
MX2X1    g2951(.A(g1859), .B(n7577), .S0(g1862), .Y(n5544));
MX2X1    g2952(.A(g1860), .B(n7577), .S0(g1866), .Y(n5549));
MX2X1    g2953(.A(g1861), .B(n7787_1), .S0(g1855), .Y(n5554));
MX2X1    g2954(.A(g1865), .B(n7787_1), .S0(g1862), .Y(n5559));
MX2X1    g2955(.A(g1845), .B(n7787_1), .S0(g1866), .Y(n5564));
MX2X1    g2956(.A(g1846), .B(n7588), .S0(g1855), .Y(n5569));
MX2X1    g2957(.A(g1849), .B(n7588), .S0(g1862), .Y(n5574));
MX2X1    g2958(.A(g1852), .B(n7588), .S0(g1866), .Y(n5579));
NAND2X1  g2959(.A(g1945), .B(g1925), .Y(n8004));
AOI22X1  g2960(.A0(g1947), .A1(g1931), .B0(g1930), .B1(g1870), .Y(n8005));
AND2X1   g2961(.A(n8005), .B(n8004), .Y(n5584));
INVX1    g2962(.A(g1931), .Y(n8007_1));
NOR2X1   g2963(.A(g1858), .B(n8007_1), .Y(n8008));
OAI22X1  g2964(.A0(g1859), .A1(n7982_1), .B0(n5312), .B1(g1860), .Y(n8009));
NOR2X1   g2965(.A(n8009), .B(n8008), .Y(n5597));
NOR2X1   g2966(.A(g1861), .B(n8007_1), .Y(n8011));
OAI22X1  g2967(.A0(g1865), .A1(n7982_1), .B0(n5312), .B1(g1845), .Y(n8012_1));
NOR2X1   g2968(.A(n8012_1), .B(n8011), .Y(n5611));
NOR2X1   g2969(.A(g1867), .B(n8007_1), .Y(n8014));
OAI22X1  g2970(.A0(g1868), .A1(n7982_1), .B0(n5312), .B1(g1869), .Y(n8015));
NOR2X1   g2971(.A(n8015), .B(n8014), .Y(n5620));
NOR2X1   g2972(.A(g1962), .B(n5312), .Y(n8017_1));
OAI22X1  g2973(.A0(g1963), .A1(n8007_1), .B0(n7982_1), .B1(g1961), .Y(n8018));
NOR2X1   g2974(.A(g1959), .B(n5312), .Y(n8019));
OAI22X1  g2975(.A0(g1960), .A1(n8007_1), .B0(n7982_1), .B1(g1958), .Y(n8020));
NOR2X1   g2976(.A(n8020), .B(n8019), .Y(n8021));
OR4X1    g2977(.A(n8018), .B(n8017_1), .C(g3229), .D(n8021), .Y(n8022_1));
NOR2X1   g2978(.A(g1965), .B(n5312), .Y(n8023));
OAI22X1  g2979(.A0(g1966), .A1(n8007_1), .B0(n7982_1), .B1(g1964), .Y(n8024));
NOR2X1   g2980(.A(n8024), .B(n8023), .Y(n8025));
OAI21X1  g2981(.A0(n8025), .A1(n5718), .B0(n8022_1), .Y(n8026));
INVX1    g2982(.A(n8021), .Y(n5784));
INVX1    g2983(.A(n8025), .Y(n5774));
NOR2X1   g2984(.A(g1956), .B(n5312), .Y(n8029));
OAI22X1  g2985(.A0(g1957), .A1(n8007_1), .B0(n7982_1), .B1(g1955), .Y(n8030));
NOR2X1   g2986(.A(n8030), .B(n8029), .Y(n8031));
NOR4X1   g2987(.A(n5774), .B(n5784), .C(n5718), .D(n8031), .Y(n8032_1));
NOR4X1   g2988(.A(n8024), .B(n8023), .C(g3229), .D(n8031), .Y(n8033));
NOR2X1   g2989(.A(n8018), .B(n8017_1), .Y(n8034));
NOR3X1   g2990(.A(n8031), .B(n8034), .C(n5718), .Y(n8035));
NOR4X1   g2991(.A(n8033), .B(n8032_1), .C(n8026), .D(n8035), .Y(n8036));
NAND2X1  g2992(.A(g1871), .B(g1925), .Y(n8037_1));
AOI22X1  g2993(.A0(g1874), .A1(g1931), .B0(g1930), .B1(g1877), .Y(n8038));
AND2X1   g2994(.A(n8038), .B(n8037_1), .Y(n8039));
INVX1    g2995(.A(n8039), .Y(n8040));
NAND2X1  g2996(.A(g1994), .B(g1925), .Y(n8041));
AOI22X1  g2997(.A0(g1997), .A1(g1931), .B0(g1930), .B1(g2000), .Y(n8042_1));
AND2X1   g2998(.A(n8042_1), .B(n8041), .Y(n8043));
INVX1    g2999(.A(n8043), .Y(n8044));
NAND3X1  g3000(.A(n8039), .B(n8044), .C(g1890), .Y(n8045));
NAND2X1  g3001(.A(g1985), .B(g1925), .Y(n8046));
AOI22X1  g3002(.A0(g1988), .A1(g1931), .B0(g1930), .B1(g1991), .Y(n8047_1));
AND2X1   g3003(.A(n8047_1), .B(n8046), .Y(n8048));
INVX1    g3004(.A(n8048), .Y(n8049));
AOI22X1  g3005(.A0(n8045), .A1(n6049), .B0(n8040), .B1(n8049), .Y(n5769));
NAND2X1  g3006(.A(n5769), .B(g1925), .Y(n8051));
MX2X1    g3007(.A(n8036), .B(g1956), .S0(n8051), .Y(n5629));
NAND2X1  g3008(.A(n5769), .B(g1931), .Y(n8053));
MX2X1    g3009(.A(n8036), .B(g1957), .S0(n8053), .Y(n5634));
NAND2X1  g3010(.A(n5769), .B(g1930), .Y(n8055));
MX2X1    g3011(.A(n8036), .B(g1955), .S0(n8055), .Y(n5639));
NOR4X1   g3012(.A(n8029), .B(n8034), .C(g3229), .D(n8030), .Y(n8057_1));
NOR3X1   g3013(.A(n8021), .B(n8018), .C(n8017_1), .Y(n8058));
NOR3X1   g3014(.A(n8058), .B(n8057_1), .C(n8035), .Y(n8059));
MX2X1    g3015(.A(n8059), .B(g1959), .S0(n8051), .Y(n5644));
MX2X1    g3016(.A(n8059), .B(g1960), .S0(n8053), .Y(n5649));
MX2X1    g3017(.A(n8059), .B(g1958), .S0(n8055), .Y(n5654));
NOR4X1   g3018(.A(n8029), .B(n8021), .C(n5718), .D(n8030), .Y(n8063));
NOR3X1   g3019(.A(n8031), .B(n8021), .C(g3229), .Y(n8064));
INVX1    g3020(.A(n8031), .Y(n5789));
NOR4X1   g3021(.A(n5774), .B(n5784), .C(g3229), .D(n5789), .Y(n8066));
NOR4X1   g3022(.A(n8064), .B(n8063), .C(n8032_1), .D(n8066), .Y(n8067_1));
MX2X1    g3023(.A(n8067_1), .B(g1962), .S0(n8051), .Y(n5659));
MX2X1    g3024(.A(n8067_1), .B(g1963), .S0(n8053), .Y(n5664));
MX2X1    g3025(.A(n8067_1), .B(g1961), .S0(n8055), .Y(n5669));
NOR2X1   g3026(.A(n8031), .B(g3229), .Y(n8071));
NOR3X1   g3027(.A(n8030), .B(n8029), .C(n5718), .Y(n8072_1));
NOR4X1   g3028(.A(n8019), .B(n8018), .C(n8017_1), .D(n8020), .Y(n8073));
OAI21X1  g3029(.A0(n8072_1), .A1(n8071), .B0(n8073), .Y(n8074));
MX2X1    g3030(.A(n8074), .B(g1965), .S0(n8051), .Y(n5674));
MX2X1    g3031(.A(n8074), .B(g1966), .S0(n8053), .Y(n5679));
MX2X1    g3032(.A(n8074), .B(g1964), .S0(n8055), .Y(n5684));
INVX1    g3033(.A(n5429), .Y(n8078));
AND2X1   g3034(.A(g1904), .B(g185), .Y(n8079));
NAND2X1  g3035(.A(g1967), .B(g1925), .Y(n8080));
AOI22X1  g3036(.A0(g1970), .A1(g1931), .B0(g1930), .B1(g1973), .Y(n8081));
NAND2X1  g3037(.A(n8081), .B(n8080), .Y(n8082_1));
AOI21X1  g3038(.A0(n8079), .A1(n8078), .B0(n8082_1), .Y(n8083));
NOR2X1   g3039(.A(n8083), .B(n5981_1), .Y(n8084));
MX2X1    g3040(.A(g1967), .B(n8084), .S0(g1925), .Y(n5689));
MX2X1    g3041(.A(g1970), .B(n8084), .S0(g1931), .Y(n5694));
MX2X1    g3042(.A(g1973), .B(n8084), .S0(g1930), .Y(n5699));
INVX1    g3043(.A(n5584), .Y(n8088));
AND2X1   g3044(.A(g1922), .B(g185), .Y(n8089));
NAND2X1  g3045(.A(g1976), .B(g1925), .Y(n8090));
AOI22X1  g3046(.A0(g1979), .A1(g1931), .B0(g1930), .B1(g1982), .Y(n8091));
NAND2X1  g3047(.A(n8091), .B(n8090), .Y(n8092_1));
AOI21X1  g3048(.A0(n8089), .A1(n8088), .B0(n8092_1), .Y(n8093));
NOR2X1   g3049(.A(n8093), .B(n5981_1), .Y(n8094));
MX2X1    g3050(.A(g1976), .B(n8094), .S0(g1925), .Y(n5704));
MX2X1    g3051(.A(g1979), .B(n8094), .S0(g1931), .Y(n5709));
MX2X1    g3052(.A(g1982), .B(n8094), .S0(g1930), .Y(n5714));
OR4X1    g3053(.A(n8029), .B(n8020), .C(n8019), .D(n8030), .Y(n8098));
NAND2X1  g3054(.A(g1706), .B(g1730), .Y(n8099));
AOI22X1  g3055(.A0(g1712), .A1(g1732), .B0(g1734), .B1(g1718), .Y(n8100));
AND2X1   g3056(.A(n8100), .B(n8099), .Y(n8101));
INVX1    g3057(.A(n8101), .Y(n8102_1));
NAND2X1  g3058(.A(g1706), .B(g1745), .Y(n8103));
AOI22X1  g3059(.A0(g1712), .A1(g1747), .B0(g1749), .B1(g1718), .Y(n8104));
AND2X1   g3060(.A(n8104), .B(n8103), .Y(n8105));
NAND2X1  g3061(.A(g1706), .B(g1760), .Y(n8106));
AOI22X1  g3062(.A0(g1712), .A1(g1762), .B0(g1764), .B1(g1718), .Y(n8107_1));
AND2X1   g3063(.A(n8107_1), .B(n8106), .Y(n8108));
OR4X1    g3064(.A(n8105), .B(n8102_1), .C(n8098), .D(n8108), .Y(n8109));
INVX1    g3065(.A(n8034), .Y(n5779));
INVX1    g3066(.A(n8105), .Y(n8111_1));
NAND2X1  g3067(.A(g1706), .B(g1775), .Y(n8112));
NAND2X1  g3068(.A(g1718), .B(g1705), .Y(n8113));
NAND2X1  g3069(.A(g1712), .B(g1777), .Y(n8114));
NAND3X1  g3070(.A(n8114), .B(n8113), .C(n8112), .Y(n8115));
NAND2X1  g3071(.A(n8115), .B(n8111_1), .Y(n8116_1));
OR4X1    g3072(.A(n8101), .B(n8021), .C(n5779), .D(n8116_1), .Y(n8117));
AND2X1   g3073(.A(n8108), .B(n8101), .Y(n8118));
NAND3X1  g3074(.A(n8118), .B(n8111_1), .C(n8073), .Y(n8119));
INVX1    g3075(.A(n8108), .Y(n8120));
NOR4X1   g3076(.A(n8030), .B(n8029), .C(n8034), .D(n8101), .Y(n8121_1));
NAND3X1  g3077(.A(n8121_1), .B(n8120), .C(n8111_1), .Y(n8122));
NAND4X1  g3078(.A(n8119), .B(n8117), .C(n8109), .D(n8122), .Y(n8123));
OR4X1    g3079(.A(n8101), .B(n5789), .C(n5774), .D(n8115), .Y(n8124));
AND2X1   g3080(.A(n8105), .B(n8101), .Y(n8125));
NAND3X1  g3081(.A(n8125), .B(n5789), .C(n8021), .Y(n8126_1));
NAND4X1  g3082(.A(n8101), .B(n5789), .C(n5774), .D(n8115), .Y(n8127));
OR4X1    g3083(.A(n8111_1), .B(n8031), .C(n8034), .D(n8108), .Y(n8128));
NAND4X1  g3084(.A(n8127), .B(n8126_1), .C(n8124), .D(n8128), .Y(n8129));
OR4X1    g3085(.A(n8101), .B(n8031), .C(n8034), .D(n8111_1), .Y(n8130));
OAI21X1  g3086(.A0(n8024), .A1(n8023), .B0(n8118), .Y(n8131_1));
OR4X1    g3087(.A(n8105), .B(n8101), .C(n8021), .D(n8120), .Y(n8132));
OR4X1    g3088(.A(n8030), .B(n8029), .C(n8034), .D(n8115), .Y(n8133));
NAND4X1  g3089(.A(n8132), .B(n8131_1), .C(n8130), .D(n8133), .Y(n8134));
OR4X1    g3090(.A(n8021), .B(n8018), .C(n8017_1), .D(n8101), .Y(n8135));
OR2X1    g3091(.A(n8111_1), .B(n8101), .Y(n8136_1));
OR4X1    g3092(.A(n8031), .B(n8024), .C(n8023), .D(n8108), .Y(n8137));
OAI22X1  g3093(.A0(n8136_1), .A1(n8137), .B0(n8135), .B1(n8120), .Y(n8138));
NOR4X1   g3094(.A(n8134), .B(n8129), .C(n8123), .D(n8138), .Y(n8139));
NAND4X1  g3095(.A(n8111_1), .B(n8101), .C(n8025), .D(n8120), .Y(n8140));
NOR3X1   g3096(.A(n8140), .B(n8031), .C(n5784), .Y(n8141_1));
NAND4X1  g3097(.A(n8111_1), .B(n8102_1), .C(n8034), .D(n8115), .Y(n8142));
NOR2X1   g3098(.A(n8142), .B(n8098), .Y(n8143));
NOR4X1   g3099(.A(n8101), .B(n8098), .C(n5774), .D(n8120), .Y(n8144));
NOR4X1   g3100(.A(n8102_1), .B(n8031), .C(n8034), .D(n8116_1), .Y(n8145));
OR4X1    g3101(.A(n8144), .B(n8143), .C(n8141_1), .D(n8145), .Y(n8146_1));
NAND4X1  g3102(.A(n8105), .B(n8031), .C(n5784), .D(n8120), .Y(n8147));
OR4X1    g3103(.A(n8105), .B(n8101), .C(n8025), .D(n8108), .Y(n8148));
OR4X1    g3104(.A(n8102_1), .B(n8031), .C(n8021), .D(n8120), .Y(n8149));
NAND3X1  g3105(.A(n8149), .B(n8148), .C(n8147), .Y(n8150));
NAND2X1  g3106(.A(n8121_1), .B(n8105), .Y(n8151_1));
NAND2X1  g3107(.A(n8125), .B(n8058), .Y(n8152));
OR4X1    g3108(.A(n8031), .B(n5784), .C(n5779), .D(n8115), .Y(n8153));
NAND3X1  g3109(.A(n8153), .B(n8152), .C(n8151_1), .Y(n8154));
NOR3X1   g3110(.A(n8154), .B(n8150), .C(n8146_1), .Y(n8155));
NAND2X1  g3111(.A(n8155), .B(n8093), .Y(n8156_1));
OR2X1    g3112(.A(n8156_1), .B(n8139), .Y(n8157));
INVX1    g3113(.A(n8083), .Y(n8158));
NOR2X1   g3114(.A(n8093), .B(n8158), .Y(n8159));
AOI21X1  g3115(.A0(n8159), .A1(n8155), .B0(n5982), .Y(n8160));
AOI22X1  g3116(.A0(n8157), .A1(n8160), .B0(n8043), .B1(n5982), .Y(n8161_1));
MX2X1    g3117(.A(g1994), .B(n8161_1), .S0(g1925), .Y(n5719));
MX2X1    g3118(.A(g1997), .B(n8161_1), .S0(g1931), .Y(n5724));
MX2X1    g3119(.A(g2000), .B(n8161_1), .S0(g1930), .Y(n5729));
NAND3X1  g3120(.A(n8139), .B(n8093), .C(n8158), .Y(n8165));
NOR2X1   g3121(.A(n8155), .B(n8158), .Y(n8166_1));
AOI21X1  g3122(.A0(n8166_1), .A1(n8139), .B0(n5982), .Y(n8167));
AOI22X1  g3123(.A0(n8165), .A1(n8167), .B0(n8048), .B1(n5982), .Y(n8168));
MX2X1    g3124(.A(g1985), .B(n8168), .S0(g1925), .Y(n5734));
MX2X1    g3125(.A(g1988), .B(n8168), .S0(g1931), .Y(n5739));
MX2X1    g3126(.A(g1991), .B(n8168), .S0(g1930), .Y(n5744));
INVX1    g3127(.A(g1890), .Y(n8172));
NOR3X1   g3128(.A(n8040), .B(n8044), .C(n8172), .Y(n8173));
MX2X1    g3129(.A(g1871), .B(n8173), .S0(g1925), .Y(n5749));
MX2X1    g3130(.A(g1874), .B(n8173), .S0(g1931), .Y(n5754));
MX2X1    g3131(.A(g1877), .B(n8173), .S0(g1930), .Y(n5759));
NAND2X1  g3132(.A(n4093), .B(g1931), .Y(n8177));
AOI21X1  g3133(.A0(g1896), .A1(n8007_1), .B0(g1886), .Y(n8178));
INVX1    g3134(.A(g1886), .Y(n8179));
NOR2X1   g3135(.A(g1895), .B(n8179), .Y(n8180));
AOI21X1  g3136(.A0(n8178), .A1(n8177), .B0(n8180), .Y(n5794));
NAND2X1  g3137(.A(n4098), .B(g1931), .Y(n8182));
AOI21X1  g3138(.A0(g1897), .A1(n8007_1), .B0(g1886), .Y(n8183));
NOR2X1   g3139(.A(g1894), .B(n8179), .Y(n8184));
AOI21X1  g3140(.A0(n8183), .A1(n8182), .B0(n8184), .Y(n5799));
NAND2X1  g3141(.A(n4103), .B(g1931), .Y(n8186_1));
AOI21X1  g3142(.A0(g1898), .A1(n8007_1), .B0(g1886), .Y(n8187));
NOR2X1   g3143(.A(g1889), .B(n8179), .Y(n8188));
AOI21X1  g3144(.A0(n8187), .A1(n8186_1), .B0(n8188), .Y(n5804));
NAND2X1  g3145(.A(n4108), .B(g1931), .Y(n8190));
AOI21X1  g3146(.A0(g1899), .A1(n8007_1), .B0(g1886), .Y(n8191_1));
NOR2X1   g3147(.A(g1888), .B(n8179), .Y(n8192));
AOI21X1  g3148(.A0(n8191_1), .A1(n8190), .B0(n8192), .Y(n5809));
NAND2X1  g3149(.A(n4113), .B(g1931), .Y(n8194));
AOI21X1  g3150(.A0(g1900), .A1(n8007_1), .B0(g1886), .Y(n8195));
NOR2X1   g3151(.A(g1887), .B(n8179), .Y(n8196_1));
AOI21X1  g3152(.A0(n8195), .A1(n8194), .B0(n8196_1), .Y(n5814));
INVX1    g3153(.A(g1832), .Y(n5823));
INVX1    g3154(.A(g1834), .Y(n5828));
INVX1    g3155(.A(g1660), .Y(n5833));
INVX1    g3156(.A(g1662), .Y(n5838));
INVX1    g3157(.A(g1664), .Y(n5843));
INVX1    g3158(.A(g1666), .Y(n5848));
INVX1    g3159(.A(g1668), .Y(n5853));
INVX1    g3160(.A(g1670), .Y(n5858));
INVX1    g3161(.A(g1672), .Y(n5868));
MX2X1    g3162(.A(n5868), .B(g1686), .S0(n5718), .Y(n5863));
MX2X1    g3163(.A(g2010), .B(g1890), .S0(g2009), .Y(n5886));
MX2X1    g3164(.A(g2039), .B(n6049), .S0(g2009), .Y(n5891));
INVX1    g3165(.A(g2039), .Y(n8210));
INVX1    g3166(.A(g2020), .Y(n8211_1));
NAND3X1  g3167(.A(n8211_1), .B(n8210), .C(g2009), .Y(n8212));
INVX1    g3168(.A(g2009), .Y(n8213));
OAI21X1  g3169(.A0(g2039), .A1(n8213), .B0(g2020), .Y(n8214));
AND2X1   g3170(.A(g2010), .B(g2006), .Y(n8215));
AOI21X1  g3171(.A0(n8214), .A1(n8212), .B0(n8215), .Y(n5896));
INVX1    g3172(.A(g2013), .Y(n8217));
NOR3X1   g3173(.A(n8211_1), .B(g2039), .C(n8213), .Y(n8218));
XOR2X1   g3174(.A(n8218), .B(n8217), .Y(n8219));
NOR2X1   g3175(.A(n8219), .B(n8215), .Y(n5901));
INVX1    g3176(.A(g2033), .Y(n8221_1));
NOR4X1   g3177(.A(n8211_1), .B(g2039), .C(n8213), .D(n8217), .Y(n8222));
XOR2X1   g3178(.A(n8222), .B(n8221_1), .Y(n8223));
NOR2X1   g3179(.A(n8223), .B(n8215), .Y(n5906));
INVX1    g3180(.A(g2026), .Y(n8225));
AND2X1   g3181(.A(n8222), .B(g2033), .Y(n8226_1));
XOR2X1   g3182(.A(n8226_1), .B(n8225), .Y(n8227));
NOR2X1   g3183(.A(n8227), .B(n8215), .Y(n5911));
NAND3X1  g3184(.A(n8222), .B(g2026), .C(g2033), .Y(n8229));
XOR2X1   g3185(.A(n8229), .B(g2040), .Y(n8230));
NOR2X1   g3186(.A(n8230), .B(n8215), .Y(n5916));
INVX1    g3187(.A(g2040), .Y(n8232));
OAI21X1  g3188(.A0(n8229), .A1(n8232), .B0(g2052), .Y(n8233));
INVX1    g3189(.A(g2052), .Y(n8234));
NAND4X1  g3190(.A(n8234), .B(g2040), .C(g2026), .D(n8226_1), .Y(n8235));
AOI21X1  g3191(.A0(n8235), .A1(n8233), .B0(n8215), .Y(n5921));
INVX1    g3192(.A(g2046), .Y(n8237));
NOR3X1   g3193(.A(n8229), .B(n8234), .C(n8232), .Y(n8238));
XOR2X1   g3194(.A(n8238), .B(n8237), .Y(n8239));
NOR2X1   g3195(.A(n8239), .B(n8215), .Y(n5926));
INVX1    g3196(.A(g2059), .Y(n8241));
NOR4X1   g3197(.A(n8237), .B(n8234), .C(n8232), .D(n8229), .Y(n8242));
XOR2X1   g3198(.A(n8242), .B(n8241), .Y(n8243));
NOR2X1   g3199(.A(n8243), .B(n8215), .Y(n5931));
INVX1    g3200(.A(g2066), .Y(n8245));
AND2X1   g3201(.A(n8242), .B(g2059), .Y(n8246));
XOR2X1   g3202(.A(n8246), .B(n8245), .Y(n8247));
NOR2X1   g3203(.A(n8247), .B(n8215), .Y(n5936));
NAND3X1  g3204(.A(n8242), .B(g2066), .C(g2059), .Y(n8249));
XOR2X1   g3205(.A(n8249), .B(g2072), .Y(n8250));
NOR2X1   g3206(.A(n8250), .B(n8215), .Y(n5941));
NAND4X1  g3207(.A(g2003), .B(g1918), .C(g1905), .D(n8210), .Y(n8252));
MX2X1    g3208(.A(n8211_1), .B(g2079), .S0(n8252), .Y(n5946));
NAND4X1  g3209(.A(g2006), .B(g1918), .C(g1905), .D(n8210), .Y(n8254));
MX2X1    g3210(.A(n8211_1), .B(g2080), .S0(n8254), .Y(n5951));
NAND4X1  g3211(.A(g2009), .B(g1918), .C(g1905), .D(n8210), .Y(n8256));
MX2X1    g3212(.A(n8211_1), .B(g2078), .S0(n8256), .Y(n5956));
MX2X1    g3213(.A(n8217), .B(g2082), .S0(n8252), .Y(n5961));
MX2X1    g3214(.A(n8217), .B(g2083), .S0(n8254), .Y(n5966));
MX2X1    g3215(.A(n8217), .B(g2081), .S0(n8256), .Y(n5971));
MX2X1    g3216(.A(n8221_1), .B(g2085), .S0(n8252), .Y(n5976));
MX2X1    g3217(.A(n8221_1), .B(g2086), .S0(n8254), .Y(n5981));
MX2X1    g3218(.A(n8221_1), .B(g2084), .S0(n8256), .Y(n5986));
MX2X1    g3219(.A(n8225), .B(g2088), .S0(n8252), .Y(n5991));
MX2X1    g3220(.A(n8225), .B(g2089), .S0(n8254), .Y(n5996));
MX2X1    g3221(.A(n8225), .B(g2087), .S0(n8256), .Y(n6001));
MX2X1    g3222(.A(n8232), .B(g2091), .S0(n8252), .Y(n6006));
MX2X1    g3223(.A(n8232), .B(g2092), .S0(n8254), .Y(n6011));
MX2X1    g3224(.A(n8232), .B(g2090), .S0(n8256), .Y(n6016));
MX2X1    g3225(.A(n8234), .B(g2094), .S0(n8252), .Y(n6021));
MX2X1    g3226(.A(n8234), .B(g2095), .S0(n8254), .Y(n6026));
MX2X1    g3227(.A(n8234), .B(g2093), .S0(n8256), .Y(n6031));
MX2X1    g3228(.A(n8237), .B(g2097), .S0(n8252), .Y(n6036));
MX2X1    g3229(.A(n8237), .B(g2098), .S0(n8254), .Y(n6041));
MX2X1    g3230(.A(n8237), .B(g2096), .S0(n8256), .Y(n6046));
MX2X1    g3231(.A(n8241), .B(g2100), .S0(n8252), .Y(n6051));
MX2X1    g3232(.A(n8241), .B(g2101), .S0(n8254), .Y(n6056));
MX2X1    g3233(.A(n8241), .B(g2099), .S0(n8256), .Y(n6061));
MX2X1    g3234(.A(n8245), .B(g2103), .S0(n8252), .Y(n6066));
MX2X1    g3235(.A(n8245), .B(g2104), .S0(n8254), .Y(n6071));
MX2X1    g3236(.A(n8245), .B(g2102), .S0(n8256), .Y(n6076));
INVX1    g3237(.A(g2072), .Y(n8282));
MX2X1    g3238(.A(n8282), .B(g2106), .S0(n8252), .Y(n6081));
MX2X1    g3239(.A(n8282), .B(g2107), .S0(n8254), .Y(n6086));
MX2X1    g3240(.A(n8282), .B(g2105), .S0(n8256), .Y(n6091));
AND2X1   g3241(.A(g2010), .B(g2003), .Y(n8286));
MX2X1    g3242(.A(g2109), .B(n8043), .S0(n8286), .Y(n6096));
MX2X1    g3243(.A(g2110), .B(n8043), .S0(n8215), .Y(n6101));
AND2X1   g3244(.A(g2010), .B(g2009), .Y(n8289));
MX2X1    g3245(.A(g2108), .B(n8043), .S0(n8289), .Y(n6106));
MX2X1    g3246(.A(g2112), .B(n8048), .S0(n8286), .Y(n6111));
MX2X1    g3247(.A(g2113), .B(n8048), .S0(n8215), .Y(n6116));
MX2X1    g3248(.A(g2111), .B(n8048), .S0(n8289), .Y(n6121));
INVX1    g3249(.A(g2003), .Y(n8294));
NOR2X1   g3250(.A(g2097), .B(n8294), .Y(n8295));
INVX1    g3251(.A(g2006), .Y(n8296));
OAI22X1  g3252(.A0(g2098), .A1(n8296), .B0(n8213), .B1(g2096), .Y(n8297));
NOR2X1   g3253(.A(n8297), .B(n8295), .Y(n8298));
XOR2X1   g3254(.A(n8298), .B(n8237), .Y(n8299));
NOR2X1   g3255(.A(g2103), .B(n8294), .Y(n8300));
OAI22X1  g3256(.A0(g2104), .A1(n8296), .B0(n8213), .B1(g2102), .Y(n8301));
NOR2X1   g3257(.A(n8301), .B(n8300), .Y(n8302));
XOR2X1   g3258(.A(n8302), .B(n8245), .Y(n8303));
NOR2X1   g3259(.A(g2100), .B(n8294), .Y(n8304));
OAI22X1  g3260(.A0(g2101), .A1(n8296), .B0(n8213), .B1(g2099), .Y(n8305));
NOR2X1   g3261(.A(n8305), .B(n8304), .Y(n8306));
XOR2X1   g3262(.A(n8306), .B(n8241), .Y(n8307));
NOR2X1   g3263(.A(g2094), .B(n8294), .Y(n8308));
OAI22X1  g3264(.A0(g2095), .A1(n8296), .B0(n8213), .B1(g2093), .Y(n8309));
NOR2X1   g3265(.A(n8309), .B(n8308), .Y(n8310));
XOR2X1   g3266(.A(n8310), .B(n8234), .Y(n8311));
OR4X1    g3267(.A(n8307), .B(n8303), .C(n8299), .D(n8311), .Y(n8312));
NOR2X1   g3268(.A(g2088), .B(n8294), .Y(n8313));
OAI22X1  g3269(.A0(g2089), .A1(n8296), .B0(n8213), .B1(g2087), .Y(n8314));
OR2X1    g3270(.A(n8314), .B(n8313), .Y(n8315));
XOR2X1   g3271(.A(n8315), .B(n8225), .Y(n8316));
NOR2X1   g3272(.A(g2091), .B(n8294), .Y(n8317));
OAI22X1  g3273(.A0(g2092), .A1(n8296), .B0(n8213), .B1(g2090), .Y(n8318));
NOR2X1   g3274(.A(n8318), .B(n8317), .Y(n8319));
XOR2X1   g3275(.A(n8319), .B(g2040), .Y(n8320));
NAND2X1  g3276(.A(n8320), .B(n8316), .Y(n8321));
NOR2X1   g3277(.A(g2079), .B(n8294), .Y(n8322));
OAI22X1  g3278(.A0(g2080), .A1(n8296), .B0(n8213), .B1(g2078), .Y(n8323));
NOR2X1   g3279(.A(n8323), .B(n8322), .Y(n8324));
XOR2X1   g3280(.A(n8324), .B(g2020), .Y(n8325));
NOR2X1   g3281(.A(g2082), .B(n8294), .Y(n8326));
OAI22X1  g3282(.A0(g2083), .A1(n8296), .B0(n8213), .B1(g2081), .Y(n8327));
NOR2X1   g3283(.A(n8327), .B(n8326), .Y(n8328));
XOR2X1   g3284(.A(n8328), .B(g2013), .Y(n8329));
NAND2X1  g3285(.A(n8329), .B(n8325), .Y(n8330));
NOR2X1   g3286(.A(g2106), .B(n8294), .Y(n8331));
OAI22X1  g3287(.A0(g2107), .A1(n8296), .B0(n8213), .B1(g2105), .Y(n8332));
NOR2X1   g3288(.A(n8332), .B(n8331), .Y(n8333));
XOR2X1   g3289(.A(n8333), .B(n8282), .Y(n8334));
NOR2X1   g3290(.A(g2085), .B(n8294), .Y(n8335));
OAI22X1  g3291(.A0(g2086), .A1(n8296), .B0(n8213), .B1(g2084), .Y(n8336));
NOR2X1   g3292(.A(n8336), .B(n8335), .Y(n8337));
XOR2X1   g3293(.A(n8337), .B(n8221_1), .Y(n8338));
OR2X1    g3294(.A(n8338), .B(n8334), .Y(n8339));
NOR4X1   g3295(.A(n8330), .B(n8321), .C(n8312), .D(n8339), .Y(n8340));
INVX1    g3296(.A(g2113), .Y(n8341));
INVX1    g3297(.A(g2111), .Y(n8342));
AOI22X1  g3298(.A0(n8341), .A1(g2006), .B0(g2009), .B1(n8342), .Y(n8343));
OAI21X1  g3299(.A0(g2112), .A1(n8294), .B0(n8343), .Y(n8344));
NOR2X1   g3300(.A(g2109), .B(n8294), .Y(n8345));
OAI22X1  g3301(.A0(g2110), .A1(n8296), .B0(n8213), .B1(g2108), .Y(n8346));
NOR4X1   g3302(.A(n8345), .B(n8344), .C(n8340), .D(n8346), .Y(n8347));
MX2X1    g3303(.A(n8347), .B(g2115), .S0(n8252), .Y(n6126));
MX2X1    g3304(.A(n8347), .B(g2116), .S0(n8254), .Y(n6131));
MX2X1    g3305(.A(n8347), .B(g2114), .S0(n8256), .Y(n6136));
INVX1    g3306(.A(g2010), .Y(n8351));
INVX1    g3307(.A(g1905), .Y(n8352));
INVX1    g3308(.A(g1918), .Y(n8353));
NOR3X1   g3309(.A(g2039), .B(n8353), .C(n8352), .Y(n8354));
OAI21X1  g3310(.A0(n8354), .A1(g2010), .B0(g2003), .Y(n8355));
MX2X1    g3311(.A(n8351), .B(g2118), .S0(n8355), .Y(n6141));
OAI21X1  g3312(.A0(n8354), .A1(g2010), .B0(g2006), .Y(n8357));
MX2X1    g3313(.A(n8351), .B(g2119), .S0(n8357), .Y(n6146));
OAI21X1  g3314(.A0(n8354), .A1(g2010), .B0(g2009), .Y(n8359));
MX2X1    g3315(.A(n8351), .B(g2117), .S0(n8359), .Y(n6151));
INVX1    g3316(.A(g2165), .Y(n6898));
NAND2X1  g3317(.A(g2257), .B(g2214), .Y(n8362));
MX2X1    g3318(.A(n6898), .B(g2206), .S0(n8362), .Y(n6169));
NAND2X1  g3319(.A(g2257), .B(g2211), .Y(n8364));
MX2X1    g3320(.A(n6898), .B(g2207), .S0(n8364), .Y(n6174));
AND2X1   g3321(.A(g2257), .B(g2241), .Y(n8366));
MX2X1    g3322(.A(g2205), .B(n6898), .S0(n8366), .Y(n6179));
INVX1    g3323(.A(g2170), .Y(n6889));
MX2X1    g3324(.A(n6889), .B(g2209), .S0(n8362), .Y(n6184));
MX2X1    g3325(.A(n6889), .B(g2210), .S0(n8364), .Y(n6189));
MX2X1    g3326(.A(g2208), .B(n6889), .S0(n8366), .Y(n6194));
INVX1    g3327(.A(g2175), .Y(n6880));
MX2X1    g3328(.A(n6880), .B(g2218), .S0(n8362), .Y(n6199));
MX2X1    g3329(.A(n6880), .B(g2219), .S0(n8364), .Y(n6204));
MX2X1    g3330(.A(g2217), .B(n6880), .S0(n8366), .Y(n6209));
INVX1    g3331(.A(g2180), .Y(n6871));
MX2X1    g3332(.A(n6871), .B(g2221), .S0(n8362), .Y(n6214));
MX2X1    g3333(.A(n6871), .B(g2222), .S0(n8364), .Y(n6219));
MX2X1    g3334(.A(g2220), .B(n6871), .S0(n8366), .Y(n6224));
INVX1    g3335(.A(g2185), .Y(n6862));
MX2X1    g3336(.A(n6862), .B(g2224), .S0(n8362), .Y(n6229));
MX2X1    g3337(.A(n6862), .B(g2225), .S0(n8364), .Y(n6234));
MX2X1    g3338(.A(g2223), .B(n6862), .S0(n8366), .Y(n6239));
INVX1    g3339(.A(g2190), .Y(n6853));
MX2X1    g3340(.A(n6853), .B(g2227), .S0(n8362), .Y(n6244));
MX2X1    g3341(.A(n6853), .B(g2228), .S0(n8364), .Y(n6249));
MX2X1    g3342(.A(g2226), .B(n6853), .S0(n8366), .Y(n6254));
INVX1    g3343(.A(g2195), .Y(n6844));
MX2X1    g3344(.A(n6844), .B(g2230), .S0(n8362), .Y(n6259));
MX2X1    g3345(.A(n6844), .B(g2231), .S0(n8364), .Y(n6264));
MX2X1    g3346(.A(g2229), .B(n6844), .S0(n8366), .Y(n6269));
INVX1    g3347(.A(g2200), .Y(n6835));
MX2X1    g3348(.A(n6835), .B(g2233), .S0(n8362), .Y(n6274));
MX2X1    g3349(.A(n6835), .B(g2234), .S0(n8364), .Y(n6279));
MX2X1    g3350(.A(g2232), .B(n6835), .S0(n8366), .Y(n6284));
INVX1    g3351(.A(g2214), .Y(n8396));
NOR2X1   g3352(.A(g2251), .B(n8396), .Y(n8397));
INVX1    g3353(.A(g2211), .Y(n8398));
INVX1    g3354(.A(g2241), .Y(n8399));
OAI22X1  g3355(.A0(g2252), .A1(n8398), .B0(n8399), .B1(g2250), .Y(n8400));
NOR2X1   g3356(.A(n8400), .B(n8397), .Y(n8401));
MX2X1    g3357(.A(n8401), .B(g2236), .S0(n8362), .Y(n6289));
MX2X1    g3358(.A(n8401), .B(g2237), .S0(n8364), .Y(n6294));
MX2X1    g3359(.A(g2235), .B(n8401), .S0(n8366), .Y(n6299));
NOR2X1   g3360(.A(g2248), .B(n8396), .Y(n8405));
OAI22X1  g3361(.A0(g2249), .A1(n8398), .B0(n8399), .B1(g2247), .Y(n8406));
NOR2X1   g3362(.A(n8406), .B(n8405), .Y(n8407));
MX2X1    g3363(.A(n8407), .B(g2239), .S0(n8362), .Y(n6304));
MX2X1    g3364(.A(n8407), .B(g2240), .S0(n8364), .Y(n6309));
MX2X1    g3365(.A(g2238), .B(n8407), .S0(n8366), .Y(n6314));
NOR4X1   g3366(.A(g2190), .B(g2195), .C(n6835), .D(n6862), .Y(n8411));
AND2X1   g3367(.A(n1476), .B(g2214), .Y(n8412));
MX2X1    g3368(.A(g2245), .B(n8411), .S0(n8412), .Y(n6319));
AND2X1   g3369(.A(n1476), .B(g2211), .Y(n8414));
MX2X1    g3370(.A(g2246), .B(n8411), .S0(n8414), .Y(n6324));
AND2X1   g3371(.A(n1476), .B(g2241), .Y(n8416));
MX2X1    g3372(.A(g2244), .B(n8411), .S0(n8416), .Y(n6329));
MX2X1    g3373(.A(g2248), .B(n6889), .S0(n8412), .Y(n6334));
MX2X1    g3374(.A(g2249), .B(n6889), .S0(n8414), .Y(n6339));
MX2X1    g3375(.A(g2247), .B(n6889), .S0(n8416), .Y(n6344));
MX2X1    g3376(.A(g2251), .B(n6898), .S0(n8412), .Y(n6349));
MX2X1    g3377(.A(g2252), .B(n6898), .S0(n8414), .Y(n6354));
MX2X1    g3378(.A(g2250), .B(n6898), .S0(n8416), .Y(n6359));
NAND4X1  g3379(.A(g2170), .B(g2175), .C(g2200), .D(g2165), .Y(n8424));
NAND4X1  g3380(.A(g2185), .B(g2190), .C(g2195), .D(g2180), .Y(n8425));
NOR2X1   g3381(.A(n8425), .B(n8424), .Y(n8426));
INVX1    g3382(.A(n8426), .Y(n8427));
MX2X1    g3383(.A(g2254), .B(n8427), .S0(n8412), .Y(n6364));
MX2X1    g3384(.A(g2255), .B(n8427), .S0(n8414), .Y(n6369));
MX2X1    g3385(.A(g2253), .B(n8427), .S0(n8416), .Y(n6374));
NOR2X1   g3386(.A(g2239), .B(n8396), .Y(n8431));
OAI22X1  g3387(.A0(g2240), .A1(n8398), .B0(n8399), .B1(g2238), .Y(n8432));
OR2X1    g3388(.A(n8432), .B(n8431), .Y(n8433));
AND2X1   g3389(.A(n8433), .B(n8407), .Y(n8434));
NOR2X1   g3390(.A(g2245), .B(n8396), .Y(n8435));
OAI22X1  g3391(.A0(g2246), .A1(n8398), .B0(n8399), .B1(g2244), .Y(n8436));
OAI21X1  g3392(.A0(n8436), .A1(n8435), .B0(g2257), .Y(n8437));
NOR2X1   g3393(.A(g2236), .B(n8396), .Y(n8438));
OAI22X1  g3394(.A0(g2237), .A1(n8398), .B0(n8399), .B1(g2235), .Y(n8439));
NOR2X1   g3395(.A(n8439), .B(n8438), .Y(n8440));
XOR2X1   g3396(.A(n8440), .B(n8401), .Y(n8441));
NOR2X1   g3397(.A(g2230), .B(n8396), .Y(n8442));
OAI22X1  g3398(.A0(g2231), .A1(n8398), .B0(n8399), .B1(g2229), .Y(n8443));
NOR2X1   g3399(.A(n8443), .B(n8442), .Y(n8444));
XOR2X1   g3400(.A(n8444), .B(n6844), .Y(n8445));
NOR4X1   g3401(.A(n8441), .B(n8437), .C(n8434), .D(n8445), .Y(n8446));
NOR2X1   g3402(.A(g2224), .B(n8396), .Y(n8447));
OAI22X1  g3403(.A0(g2225), .A1(n8398), .B0(n8399), .B1(g2223), .Y(n8448));
NOR2X1   g3404(.A(n8448), .B(n8447), .Y(n8449));
XOR2X1   g3405(.A(n8449), .B(n6862), .Y(n8450));
NOR2X1   g3406(.A(g2221), .B(n8396), .Y(n8451));
OAI22X1  g3407(.A0(g2222), .A1(n8398), .B0(n8399), .B1(g2220), .Y(n8452));
NOR2X1   g3408(.A(n8452), .B(n8451), .Y(n8453));
XOR2X1   g3409(.A(n8453), .B(n6871), .Y(n8454));
NOR2X1   g3410(.A(g2227), .B(n8396), .Y(n8455));
OAI22X1  g3411(.A0(g2228), .A1(n8398), .B0(n8399), .B1(g2226), .Y(n8456));
NOR2X1   g3412(.A(n8456), .B(n8455), .Y(n8457));
XOR2X1   g3413(.A(n8457), .B(n6853), .Y(n8458));
NOR2X1   g3414(.A(g2233), .B(n8396), .Y(n8459));
OAI22X1  g3415(.A0(g2234), .A1(n8398), .B0(n8399), .B1(g2232), .Y(n8460));
OAI21X1  g3416(.A0(n8460), .A1(n8459), .B0(n6835), .Y(n8461));
OAI21X1  g3417(.A0(n8433), .A1(n8407), .B0(n8461), .Y(n8462));
NOR4X1   g3418(.A(n8458), .B(n8454), .C(n8450), .D(n8462), .Y(n8463));
NOR3X1   g3419(.A(n8460), .B(n8459), .C(n6835), .Y(n8464));
NOR2X1   g3420(.A(g2218), .B(n8396), .Y(n8465));
OAI22X1  g3421(.A0(g2219), .A1(n8398), .B0(n8399), .B1(g2217), .Y(n8466));
NOR2X1   g3422(.A(n8466), .B(n8465), .Y(n8467));
XOR2X1   g3423(.A(n8467), .B(n6880), .Y(n8468));
NOR2X1   g3424(.A(g2209), .B(n8396), .Y(n8469));
OAI22X1  g3425(.A0(g2210), .A1(n8398), .B0(n8399), .B1(g2208), .Y(n8470));
NOR2X1   g3426(.A(n8470), .B(n8469), .Y(n8471));
XOR2X1   g3427(.A(n8471), .B(n6889), .Y(n8472));
NOR2X1   g3428(.A(g2206), .B(n8396), .Y(n8473));
OAI22X1  g3429(.A0(g2207), .A1(n8398), .B0(n8399), .B1(g2205), .Y(n8474));
NOR2X1   g3430(.A(n8474), .B(n8473), .Y(n8475));
XOR2X1   g3431(.A(n8475), .B(n6898), .Y(n8476));
NOR4X1   g3432(.A(n8472), .B(n8468), .C(n8464), .D(n8476), .Y(n8477));
NAND3X1  g3433(.A(n8477), .B(n8463), .C(n8446), .Y(n8478));
NAND2X1  g3434(.A(g2297), .B(g2214), .Y(n8479));
AOI22X1  g3435(.A0(g2300), .A1(g2211), .B0(g2241), .B1(g2303), .Y(n8480));
AND2X1   g3436(.A(n8480), .B(n8479), .Y(n8481));
NOR3X1   g3437(.A(n8481), .B(n8400), .C(n8397), .Y(n8482));
OR2X1    g3438(.A(g2251), .B(n8396), .Y(n8483));
INVX1    g3439(.A(g2252), .Y(n8484));
INVX1    g3440(.A(g2250), .Y(n8485));
AOI22X1  g3441(.A0(n8484), .A1(g2211), .B0(g2241), .B1(n8485), .Y(n8486));
NAND2X1  g3442(.A(n8480), .B(n8479), .Y(n8487));
AOI21X1  g3443(.A0(n8486), .A1(n8483), .B0(n8487), .Y(n8488));
NAND2X1  g3444(.A(g2288), .B(g2214), .Y(n8489));
AOI22X1  g3445(.A0(g2291), .A1(g2211), .B0(g2241), .B1(g2294), .Y(n8490));
NAND2X1  g3446(.A(n8490), .B(n8489), .Y(n8491));
XOR2X1   g3447(.A(n8491), .B(g2195), .Y(n8492));
NOR3X1   g3448(.A(n8492), .B(n8488), .C(n8482), .Y(n8493));
NAND2X1  g3449(.A(g2261), .B(g2214), .Y(n8494));
AOI22X1  g3450(.A0(g2264), .A1(g2211), .B0(g2241), .B1(g2267), .Y(n8495));
NAND2X1  g3451(.A(n8495), .B(n8494), .Y(n8496));
XOR2X1   g3452(.A(n8496), .B(g2165), .Y(n8497));
NAND2X1  g3453(.A(g2270), .B(g2214), .Y(n8498));
AOI22X1  g3454(.A0(g2273), .A1(g2211), .B0(g2241), .B1(g2276), .Y(n8499));
NAND2X1  g3455(.A(n8499), .B(n8498), .Y(n8500));
XOR2X1   g3456(.A(n8500), .B(g2175), .Y(n8501));
NAND2X1  g3457(.A(g2279), .B(g2214), .Y(n8502));
AOI22X1  g3458(.A0(g2282), .A1(g2211), .B0(g2241), .B1(g2285), .Y(n8503));
NAND2X1  g3459(.A(n8503), .B(n8502), .Y(n8504));
XOR2X1   g3460(.A(n8504), .B(g2185), .Y(n8505));
OAI21X1  g3461(.A0(n8505), .A1(n8501), .B0(n8497), .Y(n8506));
NOR2X1   g3462(.A(n8506), .B(n8493), .Y(n8507));
NOR2X1   g3463(.A(n8505), .B(n8492), .Y(n8508));
OAI22X1  g3464(.A0(n8497), .A1(n8501), .B0(n8488), .B1(n8482), .Y(n8509));
NOR2X1   g3465(.A(n8509), .B(n8508), .Y(n8510));
XOR2X1   g3466(.A(n8504), .B(n6862), .Y(n8511));
NOR2X1   g3467(.A(n8497), .B(n8492), .Y(n8512));
NOR3X1   g3468(.A(n8501), .B(n8488), .C(n8482), .Y(n8513));
NOR3X1   g3469(.A(n8513), .B(n8512), .C(n8511), .Y(n8514));
NOR3X1   g3470(.A(n8514), .B(n8510), .C(n8507), .Y(n8515));
NAND2X1  g3471(.A(g2342), .B(g2214), .Y(n8516));
AOI22X1  g3472(.A0(g2345), .A1(g2211), .B0(g2241), .B1(g2348), .Y(n8517));
AND2X1   g3473(.A(n8517), .B(n8516), .Y(n8518));
NOR3X1   g3474(.A(n8518), .B(n8406), .C(n8405), .Y(n8519));
OR2X1    g3475(.A(g2248), .B(n8396), .Y(n8520));
INVX1    g3476(.A(g2249), .Y(n8521));
INVX1    g3477(.A(g2247), .Y(n8522));
AOI22X1  g3478(.A0(n8521), .A1(g2211), .B0(g2241), .B1(n8522), .Y(n8523));
NAND2X1  g3479(.A(n8517), .B(n8516), .Y(n8524));
AOI21X1  g3480(.A0(n8523), .A1(n8520), .B0(n8524), .Y(n8525));
NAND2X1  g3481(.A(g2333), .B(g2214), .Y(n8526));
AOI22X1  g3482(.A0(g2336), .A1(g2211), .B0(g2241), .B1(g2339), .Y(n8527));
NAND2X1  g3483(.A(n8527), .B(n8526), .Y(n8528));
XOR2X1   g3484(.A(n8528), .B(g2200), .Y(n8529));
NOR3X1   g3485(.A(n8529), .B(n8525), .C(n8519), .Y(n8530));
NAND2X1  g3486(.A(g2306), .B(g2214), .Y(n8531));
AOI22X1  g3487(.A0(g2309), .A1(g2211), .B0(g2241), .B1(g2312), .Y(n8532));
NAND2X1  g3488(.A(n8532), .B(n8531), .Y(n8533));
XOR2X1   g3489(.A(n8533), .B(g2170), .Y(n8534));
NAND2X1  g3490(.A(g2315), .B(g2214), .Y(n8535));
AOI22X1  g3491(.A0(g2318), .A1(g2211), .B0(g2241), .B1(g2321), .Y(n8536));
NAND2X1  g3492(.A(n8536), .B(n8535), .Y(n8537));
XOR2X1   g3493(.A(n8537), .B(g2180), .Y(n8538));
NAND2X1  g3494(.A(g2324), .B(g2214), .Y(n8539));
AOI22X1  g3495(.A0(g2327), .A1(g2211), .B0(g2241), .B1(g2330), .Y(n8540));
NAND2X1  g3496(.A(n8540), .B(n8539), .Y(n8541));
XOR2X1   g3497(.A(n8541), .B(g2190), .Y(n8542));
OAI21X1  g3498(.A0(n8542), .A1(n8538), .B0(n8534), .Y(n8543));
NOR2X1   g3499(.A(n8543), .B(n8530), .Y(n8544));
NOR2X1   g3500(.A(n8542), .B(n8529), .Y(n8545));
OAI22X1  g3501(.A0(n8534), .A1(n8538), .B0(n8525), .B1(n8519), .Y(n8546));
NOR2X1   g3502(.A(n8546), .B(n8545), .Y(n8547));
XOR2X1   g3503(.A(n8541), .B(n6853), .Y(n8548));
NOR2X1   g3504(.A(n8534), .B(n8529), .Y(n8549));
NOR3X1   g3505(.A(n8538), .B(n8525), .C(n8519), .Y(n8550));
NOR3X1   g3506(.A(n8550), .B(n8549), .C(n8548), .Y(n8551));
NOR3X1   g3507(.A(n8551), .B(n8547), .C(n8544), .Y(n8552));
AOI21X1  g3508(.A0(n8552), .A1(n8515), .B0(n8437), .Y(n8553));
INVX1    g3509(.A(g2351), .Y(n8554));
NOR2X1   g3510(.A(g2393), .B(n8554), .Y(n8555));
INVX1    g3511(.A(g2480), .Y(n8556));
INVX1    g3512(.A(g2476), .Y(n8557));
OAI22X1  g3513(.A0(g2394), .A1(n8556), .B0(n8557), .B1(g2395), .Y(n8558));
NOR2X1   g3514(.A(n8558), .B(n8555), .Y(n8559));
NOR2X1   g3515(.A(g2390), .B(n8554), .Y(n8560));
OAI22X1  g3516(.A0(g2391), .A1(n8556), .B0(n8557), .B1(g2392), .Y(n8561));
NOR2X1   g3517(.A(n8561), .B(n8560), .Y(n8562));
NOR2X1   g3518(.A(g2387), .B(n8554), .Y(n8563));
OAI22X1  g3519(.A0(g2388), .A1(n8556), .B0(n8557), .B1(g2389), .Y(n8564));
NOR2X1   g3520(.A(n8564), .B(n8563), .Y(n8565));
INVX1    g3521(.A(n8565), .Y(n8566));
NOR2X1   g3522(.A(g2397), .B(n8554), .Y(n8567));
OAI22X1  g3523(.A0(g2398), .A1(n8556), .B0(n8557), .B1(g2396), .Y(n8568));
NOR2X1   g3524(.A(n8568), .B(n8567), .Y(n8569));
INVX1    g3525(.A(n8569), .Y(n8570));
NAND4X1  g3526(.A(n8566), .B(n8562), .C(n8559), .D(n8570), .Y(n8571));
NOR3X1   g3527(.A(n8571), .B(n8553), .C(n8478), .Y(n8572));
NOR4X1   g3528(.A(n8561), .B(n8560), .C(n8559), .D(n8565), .Y(n8573));
NAND2X1  g3529(.A(n8573), .B(n8570), .Y(n8574));
NOR2X1   g3530(.A(n8574), .B(n8478), .Y(n8575));
NOR2X1   g3531(.A(g2478), .B(n8554), .Y(n8576));
OAI22X1  g3532(.A0(g2479), .A1(n8556), .B0(n8557), .B1(g2477), .Y(n8577));
NOR2X1   g3533(.A(n8577), .B(n8576), .Y(n8578));
INVX1    g3534(.A(g2257), .Y(n8579));
NOR3X1   g3535(.A(n8436), .B(n8435), .C(n8579), .Y(n8580));
INVX1    g3536(.A(n8580), .Y(n8581));
OAI22X1  g3537(.A0(n8578), .A1(n8478), .B0(n8565), .B1(n8581), .Y(n8582));
OR4X1    g3538(.A(n8560), .B(n8558), .C(n8555), .D(n8561), .Y(n8583));
NOR3X1   g3539(.A(n8564), .B(n8563), .C(n8583), .Y(n8584));
INVX1    g3540(.A(n8584), .Y(n8585));
INVX1    g3541(.A(n8562), .Y(n8586));
NAND3X1  g3542(.A(n8565), .B(n8586), .C(n8559), .Y(n8587));
INVX1    g3543(.A(n8559), .Y(n8588));
NOR3X1   g3544(.A(n8566), .B(n8562), .C(n8588), .Y(n8589));
NAND4X1  g3545(.A(n8502), .B(n8490), .C(n8489), .D(n8503), .Y(n8590));
OR4X1    g3546(.A(n8541), .B(n8528), .C(n8496), .D(n8590), .Y(n8591));
NAND4X1  g3547(.A(n8498), .B(n8480), .C(n8479), .D(n8499), .Y(n8592));
OR4X1    g3548(.A(n8537), .B(n8533), .C(n8524), .D(n8592), .Y(n8593));
OR2X1    g3549(.A(n8593), .B(n8591), .Y(n8594));
OR2X1    g3550(.A(n8594), .B(n8589), .Y(n8595));
NAND2X1  g3551(.A(n8537), .B(n8524), .Y(n8596));
NAND3X1  g3552(.A(n8533), .B(n8500), .C(n8487), .Y(n8597));
OR4X1    g3553(.A(n8596), .B(n8591), .C(n8587), .D(n8597), .Y(n8598));
AOI22X1  g3554(.A0(n8595), .A1(n8598), .B0(n8587), .B1(n8585), .Y(n8599));
NOR4X1   g3555(.A(n8582), .B(n8575), .C(n8572), .D(n8599), .Y(n8600));
INVX1    g3556(.A(n8600), .Y(n8601));
NAND2X1  g3557(.A(n8587), .B(n8585), .Y(n8602));
XOR2X1   g3558(.A(n8602), .B(n8496), .Y(n8603));
NOR3X1   g3559(.A(n8582), .B(n8575), .C(n8572), .Y(n8604));
AOI21X1  g3560(.A0(n8599), .A1(n8604), .B0(n6898), .Y(n8605));
MX2X1    g3561(.A(n8603), .B(n8605), .S0(n8601), .Y(n8606));
MX2X1    g3562(.A(g2261), .B(n8606), .S0(g2214), .Y(n6379));
MX2X1    g3563(.A(g2264), .B(n8606), .S0(g2211), .Y(n6384));
MX2X1    g3564(.A(g2267), .B(n8606), .S0(g2241), .Y(n6389));
AND2X1   g3565(.A(n8587), .B(n8496), .Y(n8610));
OAI21X1  g3566(.A0(n8587), .A1(n8496), .B0(n8602), .Y(n8611));
OR2X1    g3567(.A(n8611), .B(n8610), .Y(n8612));
XOR2X1   g3568(.A(n8612), .B(n8533), .Y(n8613));
NAND3X1  g3569(.A(n8599), .B(n8587), .C(n8604), .Y(n8614));
MX2X1    g3570(.A(n6889), .B(n8599), .S0(n8604), .Y(n8615));
AOI22X1  g3571(.A0(n8614), .A1(n8615), .B0(n8613), .B1(n8600), .Y(n8616));
MX2X1    g3572(.A(g2306), .B(n8616), .S0(g2214), .Y(n6394));
MX2X1    g3573(.A(g2309), .B(n8616), .S0(g2211), .Y(n6399));
MX2X1    g3574(.A(g2312), .B(n8616), .S0(g2241), .Y(n6404));
XOR2X1   g3575(.A(n8589), .B(n8533), .Y(n8620));
OR2X1    g3576(.A(n8620), .B(n8612), .Y(n8621));
XOR2X1   g3577(.A(n8621), .B(n8500), .Y(n8622));
MX2X1    g3578(.A(n6880), .B(n8599), .S0(n8604), .Y(n8623));
AOI22X1  g3579(.A0(n8622), .A1(n8600), .B0(n8614), .B1(n8623), .Y(n8624));
MX2X1    g3580(.A(g2270), .B(n8624), .S0(g2214), .Y(n6409));
MX2X1    g3581(.A(g2273), .B(n8624), .S0(g2211), .Y(n6414));
MX2X1    g3582(.A(g2276), .B(n8624), .S0(g2241), .Y(n6419));
XOR2X1   g3583(.A(n8589), .B(n8500), .Y(n8628));
OR4X1    g3584(.A(n8620), .B(n8611), .C(n8610), .D(n8628), .Y(n8629));
XOR2X1   g3585(.A(n8629), .B(n8537), .Y(n8630));
MX2X1    g3586(.A(n6871), .B(n8599), .S0(n8604), .Y(n8631));
AOI22X1  g3587(.A0(n8630), .A1(n8600), .B0(n8614), .B1(n8631), .Y(n8632));
MX2X1    g3588(.A(g2315), .B(n8632), .S0(g2214), .Y(n6424));
MX2X1    g3589(.A(g2318), .B(n8632), .S0(g2211), .Y(n6429));
MX2X1    g3590(.A(g2321), .B(n8632), .S0(g2241), .Y(n6434));
XOR2X1   g3591(.A(n8589), .B(n8537), .Y(n8636));
OR2X1    g3592(.A(n8636), .B(n8628), .Y(n8637));
NOR4X1   g3593(.A(n8620), .B(n8611), .C(n8610), .D(n8637), .Y(n8638));
XOR2X1   g3594(.A(n8638), .B(n8504), .Y(n8639));
AOI21X1  g3595(.A0(n8599), .A1(n8604), .B0(n6862), .Y(n8640));
MX2X1    g3596(.A(n8639), .B(n8640), .S0(n8601), .Y(n8641));
MX2X1    g3597(.A(g2279), .B(n8641), .S0(g2214), .Y(n6439));
MX2X1    g3598(.A(g2282), .B(n8641), .S0(g2211), .Y(n6444));
MX2X1    g3599(.A(g2285), .B(n8641), .S0(g2241), .Y(n6449));
XOR2X1   g3600(.A(n8587), .B(n8504), .Y(n8645));
AND2X1   g3601(.A(n8645), .B(n8638), .Y(n8646));
XOR2X1   g3602(.A(n8646), .B(n8541), .Y(n8647));
AOI21X1  g3603(.A0(n8599), .A1(n8604), .B0(n6853), .Y(n8648));
MX2X1    g3604(.A(n8647), .B(n8648), .S0(n8601), .Y(n8649));
MX2X1    g3605(.A(g2324), .B(n8649), .S0(g2214), .Y(n6454));
MX2X1    g3606(.A(g2327), .B(n8649), .S0(g2211), .Y(n6459));
MX2X1    g3607(.A(g2330), .B(n8649), .S0(g2241), .Y(n6464));
XOR2X1   g3608(.A(n8587), .B(n8541), .Y(n8653));
NAND2X1  g3609(.A(n8653), .B(n8645), .Y(n8654));
NOR4X1   g3610(.A(n8637), .B(n8620), .C(n8612), .D(n8654), .Y(n8655));
XOR2X1   g3611(.A(n8655), .B(n8491), .Y(n8656));
AOI21X1  g3612(.A0(n8599), .A1(n8604), .B0(n6844), .Y(n8657));
MX2X1    g3613(.A(n8656), .B(n8657), .S0(n8601), .Y(n8658));
MX2X1    g3614(.A(g2288), .B(n8658), .S0(g2214), .Y(n6469));
MX2X1    g3615(.A(g2291), .B(n8658), .S0(g2211), .Y(n6474));
MX2X1    g3616(.A(g2294), .B(n8658), .S0(g2241), .Y(n6479));
XOR2X1   g3617(.A(n8587), .B(n8491), .Y(n8662));
AND2X1   g3618(.A(n8662), .B(n8655), .Y(n8663));
XOR2X1   g3619(.A(n8663), .B(n8528), .Y(n8664));
AOI21X1  g3620(.A0(n8599), .A1(n8604), .B0(n6835), .Y(n8665));
MX2X1    g3621(.A(n8664), .B(n8665), .S0(n8601), .Y(n8666));
MX2X1    g3622(.A(g2333), .B(n8666), .S0(g2214), .Y(n6484));
MX2X1    g3623(.A(g2336), .B(n8666), .S0(g2211), .Y(n6489));
MX2X1    g3624(.A(g2339), .B(n8666), .S0(g2241), .Y(n6494));
XOR2X1   g3625(.A(n8587), .B(n8528), .Y(n8670));
NAND4X1  g3626(.A(n8662), .B(n8653), .C(n8645), .D(n8670), .Y(n8671));
OR4X1    g3627(.A(n8637), .B(n8620), .C(n8612), .D(n8671), .Y(n8672));
XOR2X1   g3628(.A(n8672), .B(n8487), .Y(n8673));
MX2X1    g3629(.A(n8401), .B(n8599), .S0(n8604), .Y(n8674));
AOI22X1  g3630(.A0(n8673), .A1(n8600), .B0(n8614), .B1(n8674), .Y(n8675));
MX2X1    g3631(.A(g2297), .B(n8675), .S0(g2214), .Y(n6499));
MX2X1    g3632(.A(g2300), .B(n8675), .S0(g2211), .Y(n6504));
MX2X1    g3633(.A(g2303), .B(n8675), .S0(g2241), .Y(n6509));
XOR2X1   g3634(.A(n8589), .B(n8487), .Y(n8679));
OR2X1    g3635(.A(n8679), .B(n8672), .Y(n8680));
XOR2X1   g3636(.A(n8680), .B(n8524), .Y(n8681));
MX2X1    g3637(.A(n8407), .B(n8599), .S0(n8604), .Y(n8682));
AOI22X1  g3638(.A0(n8681), .A1(n8600), .B0(n8614), .B1(n8682), .Y(n8683));
MX2X1    g3639(.A(g2342), .B(n8683), .S0(g2214), .Y(n6514));
MX2X1    g3640(.A(g2345), .B(n8683), .S0(g2211), .Y(n6519));
MX2X1    g3641(.A(g2348), .B(n8683), .S0(g2241), .Y(n6524));
INVX1    g3642(.A(g2160), .Y(n8687));
NOR2X1   g3643(.A(n5399), .B(n8399), .Y(n8688));
XOR2X1   g3644(.A(n8688), .B(n8687), .Y(n8689));
AOI21X1  g3645(.A0(n8366), .A1(n5399), .B0(n8689), .Y(n6529));
INVX1    g3646(.A(g2156), .Y(n8691));
NOR3X1   g3647(.A(n5399), .B(n8687), .C(n8399), .Y(n8692));
XOR2X1   g3648(.A(n8692), .B(n8691), .Y(n8693));
AOI21X1  g3649(.A0(n8366), .A1(n5399), .B0(n8693), .Y(n6534));
INVX1    g3650(.A(g2151), .Y(n8695));
NOR4X1   g3651(.A(n8691), .B(n8687), .C(n8399), .D(n5399), .Y(n8696));
XOR2X1   g3652(.A(n8696), .B(n8695), .Y(n8697));
AOI21X1  g3653(.A0(n8366), .A1(n5399), .B0(n8697), .Y(n6539));
NAND2X1  g3654(.A(n8696), .B(g2151), .Y(n8699));
XOR2X1   g3655(.A(n8699), .B(g2147), .Y(n8700));
AOI21X1  g3656(.A0(n8366), .A1(n5399), .B0(n8700), .Y(n6544));
NAND3X1  g3657(.A(n8696), .B(g2147), .C(g2151), .Y(n8702));
XOR2X1   g3658(.A(n8702), .B(g2142), .Y(n8703));
AOI21X1  g3659(.A0(n8366), .A1(n5399), .B0(n8703), .Y(n6549));
INVX1    g3660(.A(g2147), .Y(n8705));
INVX1    g3661(.A(g2142), .Y(n8706));
OR4X1    g3662(.A(g2138), .B(n8706), .C(n8705), .D(n8699), .Y(n8707));
OAI21X1  g3663(.A0(n8702), .A1(n8706), .B0(g2138), .Y(n8708));
AOI22X1  g3664(.A0(n8707), .A1(n8708), .B0(n8366), .B1(n5399), .Y(n6554));
INVX1    g3665(.A(g2138), .Y(n8710));
OR4X1    g3666(.A(n8710), .B(n8706), .C(n8705), .D(n8699), .Y(n8711));
XOR2X1   g3667(.A(n8711), .B(g2133), .Y(n8712));
AOI21X1  g3668(.A0(n8366), .A1(n5399), .B0(n8712), .Y(n6559));
INVX1    g3669(.A(g2129), .Y(n8714));
INVX1    g3670(.A(g2133), .Y(n8715));
NOR4X1   g3671(.A(n8715), .B(n8710), .C(n8706), .D(n8702), .Y(n8716));
XOR2X1   g3672(.A(n8716), .B(n8714), .Y(n8717));
AOI21X1  g3673(.A0(n8366), .A1(n5399), .B0(n8717), .Y(n6564));
INVX1    g3674(.A(g2124), .Y(n8719));
AND2X1   g3675(.A(n8716), .B(g2129), .Y(n8720));
XOR2X1   g3676(.A(n8720), .B(n8719), .Y(n8721));
AOI21X1  g3677(.A0(n8366), .A1(n5399), .B0(n8721), .Y(n6569));
INVX1    g3678(.A(g2120), .Y(n8723));
NOR4X1   g3679(.A(n8719), .B(n8714), .C(n8715), .D(n8711), .Y(n8724));
XOR2X1   g3680(.A(n8724), .B(n8723), .Y(n8725));
AOI21X1  g3681(.A0(n8366), .A1(n5399), .B0(n8725), .Y(n6574));
NOR2X1   g3682(.A(g2459), .B(n8554), .Y(n8727));
OAI22X1  g3683(.A0(g2448), .A1(n8556), .B0(n8557), .B1(g2451), .Y(n8728));
NOR2X1   g3684(.A(g2444), .B(n8554), .Y(n8729));
OAI22X1  g3685(.A0(g2433), .A1(n8556), .B0(n8557), .B1(g2436), .Y(n8730));
NOR2X1   g3686(.A(n8730), .B(n8729), .Y(n8731));
OR4X1    g3687(.A(n8728), .B(n8727), .C(g3229), .D(n8731), .Y(n8732));
NOR2X1   g3688(.A(g2473), .B(n8554), .Y(n8733));
OAI22X1  g3689(.A0(g2463), .A1(n8556), .B0(n8557), .B1(g2466), .Y(n8734));
NOR2X1   g3690(.A(n8734), .B(n8733), .Y(n8735));
OAI21X1  g3691(.A0(n8735), .A1(n5718), .B0(n8732), .Y(n8736));
INVX1    g3692(.A(n8731), .Y(n6956));
INVX1    g3693(.A(n8735), .Y(n6966));
NOR2X1   g3694(.A(g2429), .B(n8554), .Y(n8739));
OAI22X1  g3695(.A0(g2418), .A1(n8556), .B0(n8557), .B1(g2421), .Y(n8740));
NOR2X1   g3696(.A(n8740), .B(n8739), .Y(n8741));
NOR4X1   g3697(.A(n6966), .B(n6956), .C(n5718), .D(n8741), .Y(n8742));
NOR4X1   g3698(.A(n8734), .B(n8733), .C(g3229), .D(n8741), .Y(n8743));
NOR2X1   g3699(.A(n8728), .B(n8727), .Y(n8744));
NOR3X1   g3700(.A(n8741), .B(n8744), .C(n5718), .Y(n8745));
NOR4X1   g3701(.A(n8743), .B(n8742), .C(n8736), .D(n8745), .Y(n8746));
NOR4X1   g3702(.A(n8563), .B(n8562), .C(n8559), .D(n8564), .Y(n8747));
AOI21X1  g3703(.A0(n8585), .A1(n5399), .B0(n8747), .Y(n6971));
AND2X1   g3704(.A(n6971), .B(g2351), .Y(n8749));
MX2X1    g3705(.A(g2429), .B(n8746), .S0(n8749), .Y(n6610));
AND2X1   g3706(.A(n6971), .B(g2480), .Y(n8751));
MX2X1    g3707(.A(g2418), .B(n8746), .S0(n8751), .Y(n6615));
AND2X1   g3708(.A(n6971), .B(g2476), .Y(n8753));
MX2X1    g3709(.A(g2421), .B(n8746), .S0(n8753), .Y(n6620));
NOR4X1   g3710(.A(n8739), .B(n8744), .C(g3229), .D(n8740), .Y(n8755));
NOR3X1   g3711(.A(n8731), .B(n8728), .C(n8727), .Y(n8756));
NOR3X1   g3712(.A(n8756), .B(n8755), .C(n8745), .Y(n8757));
MX2X1    g3713(.A(g2444), .B(n8757), .S0(n8749), .Y(n6625));
MX2X1    g3714(.A(g2433), .B(n8757), .S0(n8751), .Y(n6630));
MX2X1    g3715(.A(g2436), .B(n8757), .S0(n8753), .Y(n6635));
NOR4X1   g3716(.A(n8739), .B(n8731), .C(n5718), .D(n8740), .Y(n8761));
NOR3X1   g3717(.A(n8741), .B(n8731), .C(g3229), .Y(n8762));
INVX1    g3718(.A(n8741), .Y(n6951));
NOR4X1   g3719(.A(n6966), .B(n6956), .C(g3229), .D(n6951), .Y(n8764));
NOR4X1   g3720(.A(n8762), .B(n8761), .C(n8742), .D(n8764), .Y(n8765));
MX2X1    g3721(.A(g2459), .B(n8765), .S0(n8749), .Y(n6640));
MX2X1    g3722(.A(g2448), .B(n8765), .S0(n8751), .Y(n6645));
MX2X1    g3723(.A(g2451), .B(n8765), .S0(n8753), .Y(n6650));
NOR2X1   g3724(.A(n8741), .B(g3229), .Y(n8769));
NOR3X1   g3725(.A(n8740), .B(n8739), .C(n5718), .Y(n8770));
NOR4X1   g3726(.A(n8729), .B(n8728), .C(n8727), .D(n8730), .Y(n8771));
OAI21X1  g3727(.A0(n8770), .A1(n8769), .B0(n8771), .Y(n8772));
MX2X1    g3728(.A(g2473), .B(n8772), .S0(n8749), .Y(n6655));
MX2X1    g3729(.A(g2463), .B(n8772), .S0(n8751), .Y(n6660));
MX2X1    g3730(.A(g2466), .B(n8772), .S0(n8753), .Y(n6665));
NAND2X1  g3731(.A(g2483), .B(g2351), .Y(n8776));
AOI22X1  g3732(.A0(g2486), .A1(g2480), .B0(g2476), .B1(g2489), .Y(n8777));
AND2X1   g3733(.A(n8777), .B(n8776), .Y(n8778));
INVX1    g3734(.A(n8778), .Y(n8779));
OR4X1    g3735(.A(n8427), .B(n8407), .C(n8401), .D(n8580), .Y(n8780));
NAND2X1  g3736(.A(g2492), .B(g2351), .Y(n8781));
AOI22X1  g3737(.A0(g2495), .A1(g2480), .B0(g2476), .B1(g2498), .Y(n8782));
AND2X1   g3738(.A(n8782), .B(n8781), .Y(n8783));
AND2X1   g3739(.A(n8783), .B(n8780), .Y(n8784));
NOR3X1   g3740(.A(n8427), .B(n8407), .C(n8401), .Y(n8785));
INVX1    g3741(.A(n8785), .Y(n8786));
OAI21X1  g3742(.A0(n8783), .A1(n8786), .B0(n8778), .Y(n8787));
INVX1    g3743(.A(n8783), .Y(n6916));
NOR2X1   g3744(.A(g2502), .B(n8554), .Y(n8789));
OAI22X1  g3745(.A0(g2503), .A1(n8556), .B0(n8557), .B1(g2501), .Y(n8790));
NOR2X1   g3746(.A(n8790), .B(n8789), .Y(n8791));
INVX1    g3747(.A(n8791), .Y(n8792));
NOR4X1   g3748(.A(n6916), .B(n8786), .C(n8580), .D(n8792), .Y(n8793));
NAND2X1  g3749(.A(n8791), .B(n6916), .Y(n8794));
OAI21X1  g3750(.A0(n8794), .A1(n8785), .B0(n8779), .Y(n8795));
OAI22X1  g3751(.A0(n8793), .A1(n8795), .B0(n8787), .B1(n8784), .Y(n8796));
AND2X1   g3752(.A(n8796), .B(g2384), .Y(n8797));
XOR2X1   g3753(.A(n8797), .B(n8779), .Y(n8798));
MX2X1    g3754(.A(g2483), .B(n8798), .S0(g2351), .Y(n6670));
MX2X1    g3755(.A(g2486), .B(n8798), .S0(g2480), .Y(n6675));
MX2X1    g3756(.A(g2489), .B(n8798), .S0(g2476), .Y(n6680));
INVX1    g3757(.A(g2384), .Y(n8802));
NAND4X1  g3758(.A(n8783), .B(n8785), .C(n8580), .D(n8778), .Y(n8803));
OAI21X1  g3759(.A0(n8792), .A1(n8580), .B0(n8785), .Y(n8804));
NAND2X1  g3760(.A(n8804), .B(n8783), .Y(n8805));
OAI21X1  g3761(.A0(n8791), .A1(n8785), .B0(n6916), .Y(n8806));
NAND3X1  g3762(.A(n8806), .B(n8805), .C(n8779), .Y(n8807));
AOI21X1  g3763(.A0(n8807), .A1(n8803), .B0(n8802), .Y(n8808));
XOR2X1   g3764(.A(n8808), .B(n6916), .Y(n8809));
MX2X1    g3765(.A(g2492), .B(n8809), .S0(g2351), .Y(n6685));
MX2X1    g3766(.A(g2495), .B(n8809), .S0(g2480), .Y(n6690));
MX2X1    g3767(.A(g2498), .B(n8809), .S0(g2476), .Y(n6695));
MX2X1    g3768(.A(n8780), .B(n8785), .S0(n6916), .Y(n8813));
OR4X1    g3769(.A(n8792), .B(n8778), .C(n8802), .D(n8813), .Y(n8814));
NAND3X1  g3770(.A(n8777), .B(n8776), .C(g2384), .Y(n8815));
OAI21X1  g3771(.A0(n8815), .A1(n8813), .B0(n8814), .Y(n8816));
AND2X1   g3772(.A(n8816), .B(g2351), .Y(n8817));
MX2X1    g3773(.A(g2502), .B(n8814), .S0(n8817), .Y(n6700));
AND2X1   g3774(.A(n8816), .B(g2480), .Y(n8819));
MX2X1    g3775(.A(g2503), .B(n8814), .S0(n8819), .Y(n6705));
AND2X1   g3776(.A(n8816), .B(g2476), .Y(n8821));
MX2X1    g3777(.A(g2501), .B(n8814), .S0(n8821), .Y(n6710));
NAND2X1  g3778(.A(g2504), .B(g2351), .Y(n8823));
AOI22X1  g3779(.A0(g2507), .A1(g2480), .B0(g2476), .B1(g2510), .Y(n8824));
NAND2X1  g3780(.A(n8824), .B(n8823), .Y(n8825));
OR2X1    g3781(.A(g2254), .B(n8396), .Y(n8826));
INVX1    g3782(.A(g2255), .Y(n8827));
INVX1    g3783(.A(g2253), .Y(n8828));
AOI22X1  g3784(.A0(n8827), .A1(g2211), .B0(g2241), .B1(n8828), .Y(n8829));
AOI21X1  g3785(.A0(n8829), .A1(n8826), .B0(n8427), .Y(n8830));
MX2X1    g3786(.A(n8825), .B(n8830), .S0(g2384), .Y(n8831));
MX2X1    g3787(.A(g2504), .B(n8831), .S0(g2351), .Y(n6715));
MX2X1    g3788(.A(g2507), .B(n8831), .S0(g2480), .Y(n6720));
MX2X1    g3789(.A(g2510), .B(n8831), .S0(g2476), .Y(n6725));
NAND2X1  g3790(.A(g2513), .B(g2351), .Y(n8835));
AOI22X1  g3791(.A0(g2516), .A1(g2480), .B0(g2476), .B1(g2519), .Y(n8836));
AND2X1   g3792(.A(n8836), .B(n8835), .Y(n8837));
INVX1    g3793(.A(n8837), .Y(n8838));
NOR2X1   g3794(.A(n8837), .B(n8825), .Y(n8839));
INVX1    g3795(.A(n8839), .Y(n8840));
AND2X1   g3796(.A(n8837), .B(n8825), .Y(n8841));
INVX1    g3797(.A(n8841), .Y(n8842));
MX2X1    g3798(.A(n8840), .B(n8842), .S0(n8830), .Y(n8843));
NOR2X1   g3799(.A(g2523), .B(n8554), .Y(n8844));
OAI22X1  g3800(.A0(g2524), .A1(n8556), .B0(n8557), .B1(g2522), .Y(n8845));
OAI21X1  g3801(.A0(n8845), .A1(n8844), .B0(g2384), .Y(n8846));
NOR2X1   g3802(.A(n8846), .B(n8843), .Y(n8847));
XOR2X1   g3803(.A(n8847), .B(n8838), .Y(n8848));
MX2X1    g3804(.A(g2513), .B(n8848), .S0(g2351), .Y(n6730));
MX2X1    g3805(.A(g2516), .B(n8848), .S0(g2480), .Y(n6735));
MX2X1    g3806(.A(g2519), .B(n8848), .S0(g2476), .Y(n6740));
NOR4X1   g3807(.A(n8844), .B(n8843), .C(n8802), .D(n8845), .Y(n8852));
INVX1    g3808(.A(n8852), .Y(n8853));
NOR2X1   g3809(.A(n8838), .B(n8825), .Y(n8854));
AOI22X1  g3810(.A0(n8835), .A1(n8836), .B0(n8824), .B1(n8823), .Y(n8855));
MX2X1    g3811(.A(n8855), .B(n8854), .S0(n8830), .Y(n8856));
AOI21X1  g3812(.A0(n8856), .A1(g2384), .B0(n8852), .Y(n8857));
NOR2X1   g3813(.A(n8857), .B(n8554), .Y(n8858));
MX2X1    g3814(.A(g2523), .B(n8853), .S0(n8858), .Y(n6745));
NOR2X1   g3815(.A(n8857), .B(n8556), .Y(n8860));
MX2X1    g3816(.A(g2524), .B(n8853), .S0(n8860), .Y(n6750));
NOR2X1   g3817(.A(n8857), .B(n8557), .Y(n8862));
MX2X1    g3818(.A(g2522), .B(n8853), .S0(n8862), .Y(n6755));
OAI21X1  g3819(.A0(n8586), .A1(n8559), .B0(n8553), .Y(n8864));
AOI21X1  g3820(.A0(n8864), .A1(n8566), .B0(n8589), .Y(n8865));
OR2X1    g3821(.A(n8578), .B(n8478), .Y(n8866));
OAI21X1  g3822(.A0(n8865), .A1(n8565), .B0(n8866), .Y(n8867));
AOI21X1  g3823(.A0(n8865), .A1(n8565), .B0(n8867), .Y(n8868));
MX2X1    g3824(.A(g2387), .B(n8868), .S0(g2351), .Y(n6760));
MX2X1    g3825(.A(g2388), .B(n8868), .S0(g2480), .Y(n6765));
MX2X1    g3826(.A(g2389), .B(n8868), .S0(g2476), .Y(n6770));
INVX1    g3827(.A(n8437), .Y(n8872));
NAND3X1  g3828(.A(n8548), .B(n8511), .C(n8493), .Y(n8873));
NOR2X1   g3829(.A(n8501), .B(n8497), .Y(n8874));
NAND2X1  g3830(.A(n8530), .B(n8874), .Y(n8875));
OR4X1    g3831(.A(n8873), .B(n8538), .C(n8534), .D(n8875), .Y(n8876));
NAND2X1  g3832(.A(n8876), .B(n8872), .Y(n8877));
NOR4X1   g3833(.A(n8569), .B(n8553), .C(n8478), .D(n8877), .Y(n8878));
NOR2X1   g3834(.A(n8552), .B(n8437), .Y(n8879));
OAI21X1  g3835(.A0(n8876), .A1(n8437), .B0(n8581), .Y(n8880));
OR4X1    g3836(.A(n8558), .B(n8555), .C(n8879), .D(n8880), .Y(n8881));
NAND4X1  g3837(.A(n8477), .B(n8463), .C(n8446), .D(n8570), .Y(n8882));
NOR2X1   g3838(.A(n8580), .B(n8559), .Y(n8883));
AOI21X1  g3839(.A0(n8883), .A1(n8882), .B0(n8586), .Y(n8884));
OAI21X1  g3840(.A0(n8881), .A1(n8878), .B0(n8884), .Y(n8885));
OR2X1    g3841(.A(n8506), .B(n8493), .Y(n8886));
OR2X1    g3842(.A(n8509), .B(n8508), .Y(n8887));
OR2X1    g3843(.A(n8497), .B(n8492), .Y(n8888));
NAND3X1  g3844(.A(n8487), .B(n8486), .C(n8483), .Y(n8889));
OAI21X1  g3845(.A0(n8400), .A1(n8397), .B0(n8481), .Y(n8890));
XOR2X1   g3846(.A(n8500), .B(n6880), .Y(n8891));
NAND3X1  g3847(.A(n8891), .B(n8890), .C(n8889), .Y(n8892));
NAND3X1  g3848(.A(n8892), .B(n8888), .C(n8505), .Y(n8893));
NAND3X1  g3849(.A(n8893), .B(n8887), .C(n8886), .Y(n8894));
AOI21X1  g3850(.A0(n8894), .A1(n8872), .B0(n8588), .Y(n8895));
OAI21X1  g3851(.A0(n8877), .A1(n8879), .B0(n8895), .Y(n8896));
AOI21X1  g3852(.A0(n8894), .A1(n8872), .B0(n8559), .Y(n8897));
NOR2X1   g3853(.A(n8897), .B(n8562), .Y(n8898));
AOI21X1  g3854(.A0(n8898), .A1(n8896), .B0(n8565), .Y(n8899));
AOI22X1  g3855(.A0(n8885), .A1(n8899), .B0(n8565), .B1(n8583), .Y(n8900));
OAI21X1  g3856(.A0(n8900), .A1(n8562), .B0(n8866), .Y(n8901));
AOI21X1  g3857(.A0(n8900), .A1(n8562), .B0(n8901), .Y(n8902));
MX2X1    g3858(.A(g2390), .B(n8902), .S0(g2351), .Y(n6775));
MX2X1    g3859(.A(g2391), .B(n8902), .S0(g2480), .Y(n6780));
MX2X1    g3860(.A(g2392), .B(n8902), .S0(g2476), .Y(n6785));
AOI21X1  g3861(.A0(n8880), .A1(n8559), .B0(n8562), .Y(n8907));
OAI21X1  g3862(.A0(n8877), .A1(n8559), .B0(n8907), .Y(n8908));
NOR2X1   g3863(.A(n8515), .B(n8437), .Y(n8909));
OR4X1    g3864(.A(n8879), .B(n8909), .C(n8802), .D(n8588), .Y(n8910));
AOI21X1  g3865(.A0(n8910), .A1(n8562), .B0(n8565), .Y(n8911));
AOI22X1  g3866(.A0(n8908), .A1(n8911), .B0(n8565), .B1(n8559), .Y(n8912));
XOR2X1   g3867(.A(n8912), .B(n8588), .Y(n8913));
AND2X1   g3868(.A(n8913), .B(n8866), .Y(n8914));
MX2X1    g3869(.A(g2393), .B(n8914), .S0(g2351), .Y(n6790));
MX2X1    g3870(.A(g2394), .B(n8914), .S0(g2480), .Y(n6795));
MX2X1    g3871(.A(g2395), .B(n8914), .S0(g2476), .Y(n6800));
NOR3X1   g3872(.A(n8588), .B(n8553), .C(n8478), .Y(n8918));
NOR3X1   g3873(.A(n8586), .B(n8559), .C(n8478), .Y(n8919));
OAI21X1  g3874(.A0(n8919), .A1(n8918), .B0(n8566), .Y(n8920));
MX2X1    g3875(.A(n8877), .B(n8802), .S0(n8573), .Y(n8921));
NOR2X1   g3876(.A(n8921), .B(n8554), .Y(n8922));
MX2X1    g3877(.A(g2397), .B(n8920), .S0(n8922), .Y(n6805));
NOR2X1   g3878(.A(n8921), .B(n8556), .Y(n8924));
MX2X1    g3879(.A(g2398), .B(n8920), .S0(n8924), .Y(n6810));
NOR2X1   g3880(.A(n8921), .B(n8557), .Y(n8926));
MX2X1    g3881(.A(g2396), .B(n8920), .S0(n8926), .Y(n6815));
NAND4X1  g3882(.A(n8477), .B(n8463), .C(n8446), .D(n8578), .Y(n8928));
AND2X1   g3883(.A(g2384), .B(g2351), .Y(n8929));
MX2X1    g3884(.A(g2478), .B(n8928), .S0(n8929), .Y(n6820));
AND2X1   g3885(.A(g2384), .B(g2480), .Y(n8931));
MX2X1    g3886(.A(g2479), .B(n8928), .S0(n8931), .Y(n6825));
AND2X1   g3887(.A(g2384), .B(g2476), .Y(n8933));
MX2X1    g3888(.A(g2477), .B(n8928), .S0(n8933), .Y(n6830));
INVX1    g3889(.A(g2374), .Y(n8935));
NAND2X1  g3890(.A(n5220), .B(g2480), .Y(n8936));
AOI21X1  g3891(.A0(g2380), .A1(n8556), .B0(n8935), .Y(n8937));
AOI22X1  g3892(.A0(n8936), .A1(n8937), .B0(g2373), .B1(n8935), .Y(n6921));
NAND2X1  g3893(.A(n5225), .B(g2480), .Y(n8939));
AOI21X1  g3894(.A0(g2383), .A1(n8556), .B0(n8935), .Y(n8940));
NOR2X1   g3895(.A(g2375), .B(g2374), .Y(n8941));
AOI21X1  g3896(.A0(n8940), .A1(n8939), .B0(n8941), .Y(n6926));
NAND2X1  g3897(.A(n5230), .B(g2480), .Y(n8943));
AOI21X1  g3898(.A0(g2372), .A1(n8556), .B0(n8935), .Y(n8944));
NOR2X1   g3899(.A(g2376), .B(g2374), .Y(n8945));
AOI21X1  g3900(.A0(n8944), .A1(n8943), .B0(n8945), .Y(n6931));
NAND2X1  g3901(.A(n5235), .B(g2480), .Y(n8947));
AOI21X1  g3902(.A0(g2371), .A1(n8556), .B0(n8935), .Y(n8948));
NOR2X1   g3903(.A(g2377), .B(g2374), .Y(n8949));
AOI21X1  g3904(.A0(n8948), .A1(n8947), .B0(n8949), .Y(n6936));
NAND2X1  g3905(.A(n5240), .B(g2480), .Y(n8951));
AOI21X1  g3906(.A0(g2370), .A1(n8556), .B0(n8935), .Y(n8952));
NOR2X1   g3907(.A(g2378), .B(g2374), .Y(n8953));
AOI21X1  g3908(.A0(n8952), .A1(n8951), .B0(n8953), .Y(n6941));
NAND2X1  g3909(.A(n5245), .B(g2480), .Y(n8955));
AOI21X1  g3910(.A0(g2369), .A1(n8556), .B0(n8935), .Y(n8956));
NOR2X1   g3911(.A(g2379), .B(g2374), .Y(n8957));
AOI21X1  g3912(.A0(n8956), .A1(n8955), .B0(n8957), .Y(n6946));
INVX1    g3913(.A(n8744), .Y(n6961));
NOR3X1   g3914(.A(n8594), .B(n8566), .C(n8583), .Y(n8960));
XOR2X1   g3915(.A(n8504), .B(n8706), .Y(n8961));
XOR2X1   g3916(.A(n8528), .B(n8714), .Y(n8962));
XOR2X1   g3917(.A(n8541), .B(n8710), .Y(n8963));
NAND3X1  g3918(.A(n8963), .B(n8962), .C(n8961), .Y(n8964));
XOR2X1   g3919(.A(n8524), .B(n8723), .Y(n8965));
XOR2X1   g3920(.A(n8533), .B(n8691), .Y(n8966));
XOR2X1   g3921(.A(n8491), .B(n8715), .Y(n8967));
XOR2X1   g3922(.A(n8487), .B(n8719), .Y(n8968));
NAND4X1  g3923(.A(n8967), .B(n8966), .C(n8965), .D(n8968), .Y(n8969));
XOR2X1   g3924(.A(n8537), .B(g2147), .Y(n8970));
XOR2X1   g3925(.A(n8500), .B(g2151), .Y(n8971));
XOR2X1   g3926(.A(n8496), .B(g2160), .Y(n8972));
OR2X1    g3927(.A(n8972), .B(n8971), .Y(n8973));
OR4X1    g3928(.A(n8970), .B(n8747), .C(n5399), .D(n8973), .Y(n8974));
NOR3X1   g3929(.A(n8974), .B(n8969), .C(n8964), .Y(n8975));
OAI21X1  g3930(.A0(n8975), .A1(n8960), .B0(n6971), .Y(n6976));
MX2X1    g3931(.A(g2628), .B(n5982), .S0(g2624), .Y(n7115));
INVX1    g3932(.A(g2624), .Y(n8978));
INVX1    g3933(.A(g2628), .Y(n8979));
MX2X1    g3934(.A(n8979), .B(g2631), .S0(n8978), .Y(n7120));
MX2X1    g3935(.A(g2584), .B(g2631), .S0(g2624), .Y(n7125));
NAND2X1  g3936(.A(g2643), .B(g2619), .Y(n8982));
AOI22X1  g3937(.A0(g2645), .A1(g2625), .B0(g2624), .B1(g2647), .Y(n8983));
AND2X1   g3938(.A(n8983), .B(n8982), .Y(n7130));
MX2X1    g3939(.A(g2561), .B(n8838), .S0(g2549), .Y(n7210));
MX2X1    g3940(.A(g2562), .B(n8838), .S0(g2556), .Y(n7215));
MX2X1    g3941(.A(g2563), .B(n8838), .S0(g2560), .Y(n7220));
MX2X1    g3942(.A(g2530), .B(n8747), .S0(g2549), .Y(n7225));
MX2X1    g3943(.A(g2533), .B(n8747), .S0(g2556), .Y(n7230));
MX2X1    g3944(.A(g2536), .B(n8747), .S0(g2560), .Y(n7235));
MX2X1    g3945(.A(g2552), .B(n8573), .S0(g2549), .Y(n7240));
MX2X1    g3946(.A(g2553), .B(n8573), .S0(g2556), .Y(n7245));
MX2X1    g3947(.A(g2554), .B(n8573), .S0(g2560), .Y(n7250));
MX2X1    g3948(.A(g2555), .B(n8783), .S0(g2549), .Y(n7255));
MX2X1    g3949(.A(g2559), .B(n8783), .S0(g2556), .Y(n7260));
MX2X1    g3950(.A(g2539), .B(n8783), .S0(g2560), .Y(n7265));
MX2X1    g3951(.A(g2540), .B(n8584), .S0(g2549), .Y(n7270));
MX2X1    g3952(.A(g2543), .B(n8584), .S0(g2556), .Y(n7275));
MX2X1    g3953(.A(g2546), .B(n8584), .S0(g2560), .Y(n7280));
NAND2X1  g3954(.A(g2639), .B(g2619), .Y(n9000));
AOI22X1  g3955(.A0(g2641), .A1(g2625), .B0(g2624), .B1(g2564), .Y(n9001));
AND2X1   g3956(.A(n9001), .B(n9000), .Y(n7285));
INVX1    g3957(.A(g2625), .Y(n9003));
NOR2X1   g3958(.A(g2552), .B(n9003), .Y(n9004));
OAI22X1  g3959(.A0(g2553), .A1(n8978), .B0(n5326), .B1(g2554), .Y(n9005));
NOR2X1   g3960(.A(n9005), .B(n9004), .Y(n7298));
NOR2X1   g3961(.A(g2555), .B(n9003), .Y(n9007));
OAI22X1  g3962(.A0(g2559), .A1(n8978), .B0(n5326), .B1(g2539), .Y(n9008));
NOR2X1   g3963(.A(n9008), .B(n9007), .Y(n7312));
NOR2X1   g3964(.A(g2561), .B(n9003), .Y(n9010));
OAI22X1  g3965(.A0(g2562), .A1(n8978), .B0(n5326), .B1(g2563), .Y(n9011));
NOR2X1   g3966(.A(n9011), .B(n9010), .Y(n7321));
NOR2X1   g3967(.A(g2656), .B(n5326), .Y(n9013));
OAI22X1  g3968(.A0(g2657), .A1(n9003), .B0(n8978), .B1(g2655), .Y(n9014));
NOR2X1   g3969(.A(g2653), .B(n5326), .Y(n9015));
OAI22X1  g3970(.A0(g2654), .A1(n9003), .B0(n8978), .B1(g2652), .Y(n9016));
NOR2X1   g3971(.A(n9016), .B(n9015), .Y(n9017));
OR4X1    g3972(.A(n9014), .B(n9013), .C(g3229), .D(n9017), .Y(n9018));
NOR2X1   g3973(.A(g2659), .B(n5326), .Y(n9019));
OAI22X1  g3974(.A0(g2660), .A1(n9003), .B0(n8978), .B1(g2658), .Y(n9020));
NOR2X1   g3975(.A(n9020), .B(n9019), .Y(n9021));
OAI21X1  g3976(.A0(n9021), .A1(n5718), .B0(n9018), .Y(n9022));
INVX1    g3977(.A(n9017), .Y(n7485));
INVX1    g3978(.A(n9021), .Y(n7475));
NOR2X1   g3979(.A(g2650), .B(n5326), .Y(n9025));
OAI22X1  g3980(.A0(g2651), .A1(n9003), .B0(n8978), .B1(g2649), .Y(n9026));
NOR2X1   g3981(.A(n9026), .B(n9025), .Y(n9027));
NOR4X1   g3982(.A(n7475), .B(n7485), .C(n5718), .D(n9027), .Y(n9028));
NOR4X1   g3983(.A(n9020), .B(n9019), .C(g3229), .D(n9027), .Y(n9029));
NOR2X1   g3984(.A(n9014), .B(n9013), .Y(n9030));
NOR3X1   g3985(.A(n9027), .B(n9030), .C(n5718), .Y(n9031));
NOR4X1   g3986(.A(n9029), .B(n9028), .C(n9022), .D(n9031), .Y(n9032));
NAND2X1  g3987(.A(g2565), .B(g2619), .Y(n9033));
AOI22X1  g3988(.A0(g2568), .A1(g2625), .B0(g2624), .B1(g2571), .Y(n9034));
AND2X1   g3989(.A(n9034), .B(n9033), .Y(n9035));
INVX1    g3990(.A(n9035), .Y(n9036));
NAND2X1  g3991(.A(g2688), .B(g2619), .Y(n9037));
AOI22X1  g3992(.A0(g2691), .A1(g2625), .B0(g2624), .B1(g2694), .Y(n9038));
AND2X1   g3993(.A(n9038), .B(n9037), .Y(n9039));
INVX1    g3994(.A(n9039), .Y(n9040));
NAND3X1  g3995(.A(n9035), .B(n9040), .C(g2584), .Y(n9041));
NAND2X1  g3996(.A(g2679), .B(g2619), .Y(n9042));
AOI22X1  g3997(.A0(g2682), .A1(g2625), .B0(g2624), .B1(g2685), .Y(n9043));
AND2X1   g3998(.A(n9043), .B(n9042), .Y(n9044));
INVX1    g3999(.A(n9044), .Y(n9045));
AOI22X1  g4000(.A0(n9041), .A1(n6049), .B0(n9036), .B1(n9045), .Y(n7470));
NAND2X1  g4001(.A(n7470), .B(g2619), .Y(n9047));
MX2X1    g4002(.A(n9032), .B(g2650), .S0(n9047), .Y(n7330));
NAND2X1  g4003(.A(n7470), .B(g2625), .Y(n9049));
MX2X1    g4004(.A(n9032), .B(g2651), .S0(n9049), .Y(n7335));
NAND2X1  g4005(.A(n7470), .B(g2624), .Y(n9051));
MX2X1    g4006(.A(n9032), .B(g2649), .S0(n9051), .Y(n7340));
NOR4X1   g4007(.A(n9025), .B(n9030), .C(g3229), .D(n9026), .Y(n9053));
NOR3X1   g4008(.A(n9017), .B(n9014), .C(n9013), .Y(n9054));
NOR3X1   g4009(.A(n9054), .B(n9053), .C(n9031), .Y(n9055));
MX2X1    g4010(.A(n9055), .B(g2653), .S0(n9047), .Y(n7345));
MX2X1    g4011(.A(n9055), .B(g2654), .S0(n9049), .Y(n7350));
MX2X1    g4012(.A(n9055), .B(g2652), .S0(n9051), .Y(n7355));
NOR4X1   g4013(.A(n9025), .B(n9017), .C(n5718), .D(n9026), .Y(n9059));
NOR3X1   g4014(.A(n9027), .B(n9017), .C(g3229), .Y(n9060));
INVX1    g4015(.A(n9027), .Y(n7490));
NOR4X1   g4016(.A(n7475), .B(n7485), .C(g3229), .D(n7490), .Y(n9062));
NOR4X1   g4017(.A(n9060), .B(n9059), .C(n9028), .D(n9062), .Y(n9063));
MX2X1    g4018(.A(n9063), .B(g2656), .S0(n9047), .Y(n7360));
MX2X1    g4019(.A(n9063), .B(g2657), .S0(n9049), .Y(n7365));
MX2X1    g4020(.A(n9063), .B(g2655), .S0(n9051), .Y(n7370));
NOR2X1   g4021(.A(n9027), .B(g3229), .Y(n9067));
NOR3X1   g4022(.A(n9026), .B(n9025), .C(n5718), .Y(n9068));
NOR4X1   g4023(.A(n9015), .B(n9014), .C(n9013), .D(n9016), .Y(n9069));
OAI21X1  g4024(.A0(n9068), .A1(n9067), .B0(n9069), .Y(n9070));
MX2X1    g4025(.A(n9070), .B(g2659), .S0(n9047), .Y(n7375));
MX2X1    g4026(.A(n9070), .B(g2660), .S0(n9049), .Y(n7380));
MX2X1    g4027(.A(n9070), .B(g2658), .S0(n9051), .Y(n7385));
INVX1    g4028(.A(n7130), .Y(n9074));
AND2X1   g4029(.A(g2598), .B(g185), .Y(n9075));
NAND2X1  g4030(.A(g2661), .B(g2619), .Y(n9076));
AOI22X1  g4031(.A0(g2664), .A1(g2625), .B0(g2624), .B1(g2667), .Y(n9077));
NAND2X1  g4032(.A(n9077), .B(n9076), .Y(n9078));
AOI21X1  g4033(.A0(n9075), .A1(n9074), .B0(n9078), .Y(n9079));
NOR2X1   g4034(.A(n9079), .B(n5981_1), .Y(n9080));
MX2X1    g4035(.A(g2661), .B(n9080), .S0(g2619), .Y(n7390));
MX2X1    g4036(.A(g2664), .B(n9080), .S0(g2625), .Y(n7395));
MX2X1    g4037(.A(g2667), .B(n9080), .S0(g2624), .Y(n7400));
INVX1    g4038(.A(n7285), .Y(n9084));
AND2X1   g4039(.A(g2616), .B(g185), .Y(n9085));
NAND2X1  g4040(.A(g2670), .B(g2619), .Y(n9086));
AOI22X1  g4041(.A0(g2673), .A1(g2625), .B0(g2624), .B1(g2676), .Y(n9087));
NAND2X1  g4042(.A(n9087), .B(n9086), .Y(n9088));
AOI21X1  g4043(.A0(n9085), .A1(n9084), .B0(n9088), .Y(n9089));
NOR2X1   g4044(.A(n9089), .B(n5981_1), .Y(n9090));
MX2X1    g4045(.A(g2670), .B(n9090), .S0(g2619), .Y(n7405));
MX2X1    g4046(.A(g2673), .B(n9090), .S0(g2625), .Y(n7410));
MX2X1    g4047(.A(g2676), .B(n9090), .S0(g2624), .Y(n7415));
OR4X1    g4048(.A(n9025), .B(n9016), .C(n9015), .D(n9026), .Y(n9094));
NAND2X1  g4049(.A(g2400), .B(g2424), .Y(n9095));
AOI22X1  g4050(.A0(g2406), .A1(g2426), .B0(g2428), .B1(g2412), .Y(n9096));
AND2X1   g4051(.A(n9096), .B(n9095), .Y(n9097));
INVX1    g4052(.A(n9097), .Y(n9098));
NAND2X1  g4053(.A(g2400), .B(g2439), .Y(n9099));
AOI22X1  g4054(.A0(g2406), .A1(g2441), .B0(g2443), .B1(g2412), .Y(n9100));
AND2X1   g4055(.A(n9100), .B(n9099), .Y(n9101));
NAND2X1  g4056(.A(g2400), .B(g2454), .Y(n9102));
AOI22X1  g4057(.A0(g2406), .A1(g2456), .B0(g2458), .B1(g2412), .Y(n9103));
AND2X1   g4058(.A(n9103), .B(n9102), .Y(n9104));
OR4X1    g4059(.A(n9101), .B(n9098), .C(n9094), .D(n9104), .Y(n9105));
INVX1    g4060(.A(n9030), .Y(n7480));
INVX1    g4061(.A(n9101), .Y(n9107));
NAND2X1  g4062(.A(g2400), .B(g2469), .Y(n9108));
NAND2X1  g4063(.A(g2412), .B(g2399), .Y(n9109));
NAND2X1  g4064(.A(g2406), .B(g2471), .Y(n9110));
NAND3X1  g4065(.A(n9110), .B(n9109), .C(n9108), .Y(n9111));
NAND2X1  g4066(.A(n9111), .B(n9107), .Y(n9112));
OR4X1    g4067(.A(n9097), .B(n9017), .C(n7480), .D(n9112), .Y(n9113));
AND2X1   g4068(.A(n9104), .B(n9097), .Y(n9114));
NAND3X1  g4069(.A(n9114), .B(n9107), .C(n9069), .Y(n9115));
INVX1    g4070(.A(n9104), .Y(n9116));
NOR4X1   g4071(.A(n9026), .B(n9025), .C(n9030), .D(n9097), .Y(n9117));
NAND3X1  g4072(.A(n9117), .B(n9116), .C(n9107), .Y(n9118));
NAND4X1  g4073(.A(n9115), .B(n9113), .C(n9105), .D(n9118), .Y(n9119));
OR4X1    g4074(.A(n9097), .B(n7490), .C(n7475), .D(n9111), .Y(n9120));
AND2X1   g4075(.A(n9101), .B(n9097), .Y(n9121));
NAND3X1  g4076(.A(n9121), .B(n7490), .C(n9017), .Y(n9122));
NAND4X1  g4077(.A(n9097), .B(n7490), .C(n7475), .D(n9111), .Y(n9123));
OR4X1    g4078(.A(n9107), .B(n9027), .C(n9030), .D(n9104), .Y(n9124));
NAND4X1  g4079(.A(n9123), .B(n9122), .C(n9120), .D(n9124), .Y(n9125));
OR4X1    g4080(.A(n9097), .B(n9027), .C(n9030), .D(n9107), .Y(n9126));
OAI21X1  g4081(.A0(n9020), .A1(n9019), .B0(n9114), .Y(n9127));
OR4X1    g4082(.A(n9101), .B(n9097), .C(n9017), .D(n9116), .Y(n9128));
OR4X1    g4083(.A(n9026), .B(n9025), .C(n9030), .D(n9111), .Y(n9129));
NAND4X1  g4084(.A(n9128), .B(n9127), .C(n9126), .D(n9129), .Y(n9130));
OR4X1    g4085(.A(n9017), .B(n9014), .C(n9013), .D(n9097), .Y(n9131));
OR2X1    g4086(.A(n9107), .B(n9097), .Y(n9132));
OR4X1    g4087(.A(n9027), .B(n9020), .C(n9019), .D(n9104), .Y(n9133));
OAI22X1  g4088(.A0(n9132), .A1(n9133), .B0(n9131), .B1(n9116), .Y(n9134));
NOR4X1   g4089(.A(n9130), .B(n9125), .C(n9119), .D(n9134), .Y(n9135));
NAND4X1  g4090(.A(n9107), .B(n9097), .C(n9021), .D(n9116), .Y(n9136));
NOR3X1   g4091(.A(n9136), .B(n9027), .C(n7485), .Y(n9137));
NAND4X1  g4092(.A(n9107), .B(n9098), .C(n9030), .D(n9111), .Y(n9138));
NOR2X1   g4093(.A(n9138), .B(n9094), .Y(n9139));
NOR4X1   g4094(.A(n9097), .B(n9094), .C(n7475), .D(n9116), .Y(n9140));
NOR4X1   g4095(.A(n9098), .B(n9027), .C(n9030), .D(n9112), .Y(n9141));
OR4X1    g4096(.A(n9140), .B(n9139), .C(n9137), .D(n9141), .Y(n9142));
NAND4X1  g4097(.A(n9101), .B(n9027), .C(n7485), .D(n9116), .Y(n9143));
OR4X1    g4098(.A(n9101), .B(n9097), .C(n9021), .D(n9104), .Y(n9144));
OR4X1    g4099(.A(n9098), .B(n9027), .C(n9017), .D(n9116), .Y(n9145));
NAND3X1  g4100(.A(n9145), .B(n9144), .C(n9143), .Y(n9146));
NAND2X1  g4101(.A(n9117), .B(n9101), .Y(n9147));
NAND2X1  g4102(.A(n9121), .B(n9054), .Y(n9148));
OR4X1    g4103(.A(n9027), .B(n7485), .C(n7480), .D(n9111), .Y(n9149));
NAND3X1  g4104(.A(n9149), .B(n9148), .C(n9147), .Y(n9150));
NOR3X1   g4105(.A(n9150), .B(n9146), .C(n9142), .Y(n9151));
NAND2X1  g4106(.A(n9151), .B(n9089), .Y(n9152));
OR2X1    g4107(.A(n9152), .B(n9135), .Y(n9153));
INVX1    g4108(.A(n9079), .Y(n9154));
NOR2X1   g4109(.A(n9089), .B(n9154), .Y(n9155));
AOI21X1  g4110(.A0(n9155), .A1(n9151), .B0(n5982), .Y(n9156));
AOI22X1  g4111(.A0(n9153), .A1(n9156), .B0(n9039), .B1(n5982), .Y(n9157));
MX2X1    g4112(.A(g2688), .B(n9157), .S0(g2619), .Y(n7420));
MX2X1    g4113(.A(g2691), .B(n9157), .S0(g2625), .Y(n7425));
MX2X1    g4114(.A(g2694), .B(n9157), .S0(g2624), .Y(n7430));
NAND3X1  g4115(.A(n9135), .B(n9089), .C(n9154), .Y(n9161));
NOR2X1   g4116(.A(n9151), .B(n9154), .Y(n9162));
AOI21X1  g4117(.A0(n9162), .A1(n9135), .B0(n5982), .Y(n9163));
AOI22X1  g4118(.A0(n9161), .A1(n9163), .B0(n9044), .B1(n5982), .Y(n9164));
MX2X1    g4119(.A(g2679), .B(n9164), .S0(g2619), .Y(n7435));
MX2X1    g4120(.A(g2682), .B(n9164), .S0(g2625), .Y(n7440));
MX2X1    g4121(.A(g2685), .B(n9164), .S0(g2624), .Y(n7445));
INVX1    g4122(.A(g2584), .Y(n9168));
NOR3X1   g4123(.A(n9036), .B(n9040), .C(n9168), .Y(n9169));
MX2X1    g4124(.A(g2565), .B(n9169), .S0(g2619), .Y(n7450));
MX2X1    g4125(.A(g2568), .B(n9169), .S0(g2625), .Y(n7455));
MX2X1    g4126(.A(g2571), .B(n9169), .S0(g2624), .Y(n7460));
INVX1    g4127(.A(g2589), .Y(n9173));
NAND2X1  g4128(.A(n5794), .B(g2625), .Y(n9174));
AOI21X1  g4129(.A0(g2590), .A1(n9003), .B0(g2580), .Y(n9175));
AOI22X1  g4130(.A0(n9174), .A1(n9175), .B0(n9173), .B1(g2580), .Y(n7495));
INVX1    g4131(.A(g2588), .Y(n9177));
NAND2X1  g4132(.A(n5799), .B(g2625), .Y(n9178));
AOI21X1  g4133(.A0(g2591), .A1(n9003), .B0(g2580), .Y(n9179));
AOI22X1  g4134(.A0(n9178), .A1(n9179), .B0(n9177), .B1(g2580), .Y(n7500));
INVX1    g4135(.A(g2583), .Y(n9181));
NAND2X1  g4136(.A(n5804), .B(g2625), .Y(n9182));
AOI21X1  g4137(.A0(g2592), .A1(n9003), .B0(g2580), .Y(n9183));
AOI22X1  g4138(.A0(n9182), .A1(n9183), .B0(n9181), .B1(g2580), .Y(n7505));
INVX1    g4139(.A(g2582), .Y(n9185));
NAND2X1  g4140(.A(n5809), .B(g2625), .Y(n9186));
AOI21X1  g4141(.A0(g2593), .A1(n9003), .B0(g2580), .Y(n9187));
AOI22X1  g4142(.A0(n9186), .A1(n9187), .B0(n9185), .B1(g2580), .Y(n7510));
INVX1    g4143(.A(g2581), .Y(n9189));
NAND2X1  g4144(.A(n5814), .B(g2625), .Y(n9190));
AOI21X1  g4145(.A0(g2594), .A1(n9003), .B0(g2580), .Y(n9191));
AOI22X1  g4146(.A0(n9190), .A1(n9191), .B0(n9189), .B1(g2580), .Y(n7515));
INVX1    g4147(.A(g2526), .Y(n7524));
INVX1    g4148(.A(g2528), .Y(n7529));
INVX1    g4149(.A(g2354), .Y(n7534));
INVX1    g4150(.A(g2356), .Y(n7539));
INVX1    g4151(.A(g2358), .Y(n7544));
INVX1    g4152(.A(g2360), .Y(n7549));
INVX1    g4153(.A(g2362), .Y(n7554));
INVX1    g4154(.A(g2364), .Y(n7559));
INVX1    g4155(.A(g2366), .Y(n7569));
MX2X1    g4156(.A(n7569), .B(g2380), .S0(n5718), .Y(n7564));
MX2X1    g4157(.A(g2704), .B(g2584), .S0(g2703), .Y(n7587));
MX2X1    g4158(.A(g2733), .B(n6049), .S0(g2703), .Y(n7592));
INVX1    g4159(.A(g2733), .Y(n9205));
INVX1    g4160(.A(g2714), .Y(n9206));
NAND3X1  g4161(.A(n9206), .B(n9205), .C(g2703), .Y(n9207));
INVX1    g4162(.A(g2703), .Y(n9208));
OAI21X1  g4163(.A0(g2733), .A1(n9208), .B0(g2714), .Y(n9209));
AND2X1   g4164(.A(g2704), .B(g2700), .Y(n9210));
AOI21X1  g4165(.A0(n9209), .A1(n9207), .B0(n9210), .Y(n7597));
INVX1    g4166(.A(g2707), .Y(n9212));
NOR3X1   g4167(.A(n9206), .B(g2733), .C(n9208), .Y(n9213));
XOR2X1   g4168(.A(n9213), .B(n9212), .Y(n9214));
NOR2X1   g4169(.A(n9214), .B(n9210), .Y(n7602));
INVX1    g4170(.A(g2727), .Y(n9216));
NOR4X1   g4171(.A(n9206), .B(g2733), .C(n9208), .D(n9212), .Y(n9217));
XOR2X1   g4172(.A(n9217), .B(n9216), .Y(n9218));
NOR2X1   g4173(.A(n9218), .B(n9210), .Y(n7607));
INVX1    g4174(.A(g2720), .Y(n9220));
AND2X1   g4175(.A(n9217), .B(g2727), .Y(n9221));
XOR2X1   g4176(.A(n9221), .B(n9220), .Y(n9222));
NOR2X1   g4177(.A(n9222), .B(n9210), .Y(n7612));
NAND3X1  g4178(.A(n9217), .B(g2720), .C(g2727), .Y(n9224));
XOR2X1   g4179(.A(n9224), .B(g2734), .Y(n9225));
NOR2X1   g4180(.A(n9225), .B(n9210), .Y(n7617));
INVX1    g4181(.A(g2734), .Y(n9227));
OAI21X1  g4182(.A0(n9224), .A1(n9227), .B0(g2746), .Y(n9228));
INVX1    g4183(.A(g2746), .Y(n9229));
NAND4X1  g4184(.A(n9229), .B(g2734), .C(g2720), .D(n9221), .Y(n9230));
AOI21X1  g4185(.A0(n9230), .A1(n9228), .B0(n9210), .Y(n7622));
INVX1    g4186(.A(g2740), .Y(n9232));
NOR3X1   g4187(.A(n9224), .B(n9229), .C(n9227), .Y(n9233));
XOR2X1   g4188(.A(n9233), .B(n9232), .Y(n9234));
NOR2X1   g4189(.A(n9234), .B(n9210), .Y(n7627));
INVX1    g4190(.A(g2753), .Y(n9236));
NOR4X1   g4191(.A(n9232), .B(n9229), .C(n9227), .D(n9224), .Y(n9237));
XOR2X1   g4192(.A(n9237), .B(n9236), .Y(n9238));
NOR2X1   g4193(.A(n9238), .B(n9210), .Y(n7632));
INVX1    g4194(.A(g2760), .Y(n9240));
AND2X1   g4195(.A(n9237), .B(g2753), .Y(n9241));
XOR2X1   g4196(.A(n9241), .B(n9240), .Y(n9242));
NOR2X1   g4197(.A(n9242), .B(n9210), .Y(n7637));
NAND3X1  g4198(.A(n9237), .B(g2760), .C(g2753), .Y(n9244));
XOR2X1   g4199(.A(n9244), .B(g2766), .Y(n9245));
NOR2X1   g4200(.A(n9245), .B(n9210), .Y(n7642));
NAND4X1  g4201(.A(g2697), .B(g2612), .C(g2599), .D(n9205), .Y(n9247));
MX2X1    g4202(.A(n9206), .B(g2773), .S0(n9247), .Y(n7647));
NAND4X1  g4203(.A(g2700), .B(g2612), .C(g2599), .D(n9205), .Y(n9249));
MX2X1    g4204(.A(n9206), .B(g2774), .S0(n9249), .Y(n7652));
NAND4X1  g4205(.A(g2703), .B(g2612), .C(g2599), .D(n9205), .Y(n9251));
MX2X1    g4206(.A(n9206), .B(g2772), .S0(n9251), .Y(n7657));
MX2X1    g4207(.A(n9212), .B(g2776), .S0(n9247), .Y(n7662));
MX2X1    g4208(.A(n9212), .B(g2777), .S0(n9249), .Y(n7667));
MX2X1    g4209(.A(n9212), .B(g2775), .S0(n9251), .Y(n7672));
MX2X1    g4210(.A(n9216), .B(g2779), .S0(n9247), .Y(n7677));
MX2X1    g4211(.A(n9216), .B(g2780), .S0(n9249), .Y(n7682));
MX2X1    g4212(.A(n9216), .B(g2778), .S0(n9251), .Y(n7687));
MX2X1    g4213(.A(n9220), .B(g2782), .S0(n9247), .Y(n7692));
MX2X1    g4214(.A(n9220), .B(g2783), .S0(n9249), .Y(n7697));
MX2X1    g4215(.A(n9220), .B(g2781), .S0(n9251), .Y(n7702));
MX2X1    g4216(.A(n9227), .B(g2785), .S0(n9247), .Y(n7707));
MX2X1    g4217(.A(n9227), .B(g2786), .S0(n9249), .Y(n7712));
MX2X1    g4218(.A(n9227), .B(g2784), .S0(n9251), .Y(n7717));
MX2X1    g4219(.A(n9229), .B(g2788), .S0(n9247), .Y(n7722));
MX2X1    g4220(.A(n9229), .B(g2789), .S0(n9249), .Y(n7727));
MX2X1    g4221(.A(n9229), .B(g2787), .S0(n9251), .Y(n7732));
MX2X1    g4222(.A(n9232), .B(g2791), .S0(n9247), .Y(n7737));
MX2X1    g4223(.A(n9232), .B(g2792), .S0(n9249), .Y(n7742));
MX2X1    g4224(.A(n9232), .B(g2790), .S0(n9251), .Y(n7747));
MX2X1    g4225(.A(n9236), .B(g2794), .S0(n9247), .Y(n7752));
MX2X1    g4226(.A(n9236), .B(g2795), .S0(n9249), .Y(n7757));
MX2X1    g4227(.A(n9236), .B(g2793), .S0(n9251), .Y(n7762));
MX2X1    g4228(.A(n9240), .B(g2797), .S0(n9247), .Y(n7767));
MX2X1    g4229(.A(n9240), .B(g2798), .S0(n9249), .Y(n7772));
MX2X1    g4230(.A(n9240), .B(g2796), .S0(n9251), .Y(n7777));
INVX1    g4231(.A(g2766), .Y(n9277));
MX2X1    g4232(.A(n9277), .B(g2800), .S0(n9247), .Y(n7782));
MX2X1    g4233(.A(n9277), .B(g2801), .S0(n9249), .Y(n7787));
MX2X1    g4234(.A(n9277), .B(g2799), .S0(n9251), .Y(n7792));
AND2X1   g4235(.A(g2704), .B(g2697), .Y(n9281));
MX2X1    g4236(.A(g2803), .B(n9039), .S0(n9281), .Y(n7797));
MX2X1    g4237(.A(g2804), .B(n9039), .S0(n9210), .Y(n7802));
AND2X1   g4238(.A(g2704), .B(g2703), .Y(n9284));
MX2X1    g4239(.A(g2802), .B(n9039), .S0(n9284), .Y(n7807));
MX2X1    g4240(.A(g2806), .B(n9044), .S0(n9281), .Y(n7812));
MX2X1    g4241(.A(g2807), .B(n9044), .S0(n9210), .Y(n7817));
MX2X1    g4242(.A(g2805), .B(n9044), .S0(n9284), .Y(n7822));
INVX1    g4243(.A(g2697), .Y(n9289));
NOR2X1   g4244(.A(g2791), .B(n9289), .Y(n9290));
INVX1    g4245(.A(g2700), .Y(n9291));
OAI22X1  g4246(.A0(g2792), .A1(n9291), .B0(n9208), .B1(g2790), .Y(n9292));
OR2X1    g4247(.A(n9292), .B(n9290), .Y(n9293));
XOR2X1   g4248(.A(n9293), .B(g2740), .Y(n9294));
NOR2X1   g4249(.A(g2797), .B(n9289), .Y(n9295));
OAI22X1  g4250(.A0(g2798), .A1(n9291), .B0(n9208), .B1(g2796), .Y(n9296));
NOR2X1   g4251(.A(n9296), .B(n9295), .Y(n9297));
XOR2X1   g4252(.A(n9297), .B(n9240), .Y(n9298));
NOR2X1   g4253(.A(g2794), .B(n9289), .Y(n9299));
OAI22X1  g4254(.A0(g2795), .A1(n9291), .B0(n9208), .B1(g2793), .Y(n9300));
NOR2X1   g4255(.A(n9300), .B(n9299), .Y(n9301));
XOR2X1   g4256(.A(n9301), .B(n9236), .Y(n9302));
NOR2X1   g4257(.A(g2788), .B(n9289), .Y(n9303));
OAI22X1  g4258(.A0(g2789), .A1(n9291), .B0(n9208), .B1(g2787), .Y(n9304));
NOR2X1   g4259(.A(n9304), .B(n9303), .Y(n9305));
XOR2X1   g4260(.A(n9305), .B(n9229), .Y(n9306));
OR4X1    g4261(.A(n9302), .B(n9298), .C(n9294), .D(n9306), .Y(n9307));
INVX1    g4262(.A(g2783), .Y(n9308));
INVX1    g4263(.A(g2781), .Y(n9309));
AOI22X1  g4264(.A0(n9308), .A1(g2700), .B0(g2703), .B1(n9309), .Y(n9310));
OAI21X1  g4265(.A0(g2782), .A1(n9289), .B0(n9310), .Y(n9311));
XOR2X1   g4266(.A(n9311), .B(n9220), .Y(n9312));
NOR2X1   g4267(.A(g2785), .B(n9289), .Y(n9313));
OAI22X1  g4268(.A0(g2786), .A1(n9291), .B0(n9208), .B1(g2784), .Y(n9314));
NOR2X1   g4269(.A(n9314), .B(n9313), .Y(n9315));
XOR2X1   g4270(.A(n9315), .B(g2734), .Y(n9316));
NAND2X1  g4271(.A(n9316), .B(n9312), .Y(n9317));
NOR2X1   g4272(.A(g2773), .B(n9289), .Y(n9318));
OAI22X1  g4273(.A0(g2774), .A1(n9291), .B0(n9208), .B1(g2772), .Y(n9319));
NOR2X1   g4274(.A(n9319), .B(n9318), .Y(n9320));
XOR2X1   g4275(.A(n9320), .B(g2714), .Y(n9321));
INVX1    g4276(.A(g2777), .Y(n9322));
INVX1    g4277(.A(g2775), .Y(n9323));
AOI22X1  g4278(.A0(n9322), .A1(g2700), .B0(g2703), .B1(n9323), .Y(n9324));
OAI21X1  g4279(.A0(g2776), .A1(n9289), .B0(n9324), .Y(n9325));
XOR2X1   g4280(.A(n9325), .B(n9212), .Y(n9326));
NAND2X1  g4281(.A(n9326), .B(n9321), .Y(n9327));
NOR2X1   g4282(.A(g2800), .B(n9289), .Y(n9328));
OAI22X1  g4283(.A0(g2801), .A1(n9291), .B0(n9208), .B1(g2799), .Y(n9329));
NOR2X1   g4284(.A(n9329), .B(n9328), .Y(n9330));
XOR2X1   g4285(.A(n9330), .B(n9277), .Y(n9331));
NOR2X1   g4286(.A(g2779), .B(n9289), .Y(n9332));
OAI22X1  g4287(.A0(g2780), .A1(n9291), .B0(n9208), .B1(g2778), .Y(n9333));
NOR2X1   g4288(.A(n9333), .B(n9332), .Y(n9334));
XOR2X1   g4289(.A(n9334), .B(n9216), .Y(n9335));
OR2X1    g4290(.A(n9335), .B(n9331), .Y(n9336));
NOR4X1   g4291(.A(n9327), .B(n9317), .C(n9307), .D(n9336), .Y(n9337));
INVX1    g4292(.A(g2807), .Y(n9338));
INVX1    g4293(.A(g2805), .Y(n9339));
AOI22X1  g4294(.A0(n9338), .A1(g2700), .B0(g2703), .B1(n9339), .Y(n9340));
OAI21X1  g4295(.A0(g2806), .A1(n9289), .B0(n9340), .Y(n9341));
NOR2X1   g4296(.A(g2803), .B(n9289), .Y(n9342));
OAI22X1  g4297(.A0(g2804), .A1(n9291), .B0(n9208), .B1(g2802), .Y(n9343));
NOR4X1   g4298(.A(n9342), .B(n9341), .C(n9337), .D(n9343), .Y(n9344));
MX2X1    g4299(.A(n9344), .B(g2809), .S0(n9247), .Y(n7827));
MX2X1    g4300(.A(n9344), .B(g2810), .S0(n9249), .Y(n7832));
MX2X1    g4301(.A(n9344), .B(g2808), .S0(n9251), .Y(n7837));
INVX1    g4302(.A(g2704), .Y(n9348));
INVX1    g4303(.A(g2599), .Y(n9349));
INVX1    g4304(.A(g2612), .Y(n9350));
NOR3X1   g4305(.A(g2733), .B(n9350), .C(n9349), .Y(n9351));
OAI21X1  g4306(.A0(n9351), .A1(g2704), .B0(g2697), .Y(n9352));
MX2X1    g4307(.A(n9348), .B(g2812), .S0(n9352), .Y(n7842));
OAI21X1  g4308(.A0(n9351), .A1(g2704), .B0(g2700), .Y(n9354));
MX2X1    g4309(.A(n9348), .B(g2813), .S0(n9354), .Y(n7847));
OAI21X1  g4310(.A0(n9351), .A1(g2704), .B0(g2703), .Y(n9356));
MX2X1    g4311(.A(n9348), .B(g2811), .S0(n9356), .Y(n7852));
INVX1    g4312(.A(g3080), .Y(n9358));
NOR2X1   g4313(.A(n9358), .B(g3234), .Y(n7857));
INVX1    g4314(.A(g3234), .Y(n9360));
AND2X1   g4315(.A(g3054), .B(n9360), .Y(n7862));
OR2X1    g4316(.A(g3079), .B(g3234), .Y(n7867));
NOR2X1   g4317(.A(g499), .B(n5297), .Y(n9363));
NOR4X1   g4318(.A(n2204), .B(g559), .C(g563), .D(n9363), .Y(n9364));
OR4X1    g4319(.A(n6311), .B(n6308), .C(n6307), .D(n6312), .Y(n9365));
NOR3X1   g4320(.A(n9365), .B(n6305), .C(n6301), .Y(n9366));
NAND2X1  g4321(.A(n6333), .B(n6328), .Y(n9367));
NOR2X1   g4322(.A(g738), .B(n6297), .Y(n9368));
OAI22X1  g4323(.A0(g739), .A1(n6299_1), .B0(n6216), .B1(g737), .Y(n9369));
OR2X1    g4324(.A(n9369), .B(n9368), .Y(n9370));
NAND4X1  g4325(.A(n6349_1), .B(n6323), .C(n6319_1), .D(n9370), .Y(n9371));
NOR4X1   g4326(.A(n9367), .B(n6342), .C(n6338), .D(n9371), .Y(n9372));
NAND2X1  g4327(.A(n9372), .B(n9366), .Y(n9373));
NOR2X1   g4328(.A(g736), .B(n6299_1), .Y(n9374));
OAI22X1  g4329(.A0(g735), .A1(n6297), .B0(n6216), .B1(g734), .Y(n9375));
NOR2X1   g4330(.A(n9375), .B(n9374), .Y(n9376));
AOI21X1  g4331(.A0(n9376), .A1(n9373), .B0(n5296), .Y(n9377));
NAND2X1  g4332(.A(n9377), .B(n9364), .Y(n9378));
INVX1    g4333(.A(g557), .Y(n9379));
NOR2X1   g4334(.A(g510), .B(n9379), .Y(n9380));
NAND2X1  g4335(.A(n9380), .B(n9378), .Y(n9381));
OAI21X1  g4336(.A0(g525), .A1(g557), .B0(n6176), .Y(n9382));
INVX1    g4337(.A(n9382), .Y(n9383));
XOR2X1   g4338(.A(n6309_1), .B(n6053), .Y(n9385));
NAND3X1  g4339(.A(n9385), .B(n9364), .C(g499), .Y(n9386));
OAI21X1  g4340(.A0(g525), .A1(g510), .B0(n9379), .Y(n9387));
NOR2X1   g4341(.A(n9382), .B(g529), .Y(n9388));
AOI21X1  g4342(.A0(n9388), .A1(n9364), .B0(n9387), .Y(n9389));
OAI21X1  g4343(.A0(n9386), .A1(n9383), .B0(n9389), .Y(n9390));
NAND2X1  g4344(.A(n9390), .B(n9381), .Y(n7872));
INVX1    g4345(.A(n9364), .Y(n9392));
OAI21X1  g4346(.A0(n9377), .A1(n9392), .B0(n9380), .Y(n9393));
XOR2X1   g4347(.A(n6301), .B(n6045), .Y(n9395));
NAND4X1  g4348(.A(n9382), .B(n9364), .C(g499), .D(n9395), .Y(n9396));
NOR2X1   g4349(.A(n9382), .B(g530), .Y(n9397));
AOI21X1  g4350(.A0(n9397), .A1(n9364), .B0(n9387), .Y(n9398));
NAND2X1  g4351(.A(n9398), .B(n9396), .Y(n9399));
NAND2X1  g4352(.A(n9399), .B(n9393), .Y(n7877));
AND2X1   g4353(.A(n9364), .B(g499), .Y(n9401));
AOI21X1  g4354(.A0(n9372), .A1(n9366), .B0(n6313), .Y(n9402));
XOR2X1   g4355(.A(n9402), .B(n6052), .Y(n9403));
NAND2X1  g4356(.A(n9403), .B(n9401), .Y(n9404));
NOR2X1   g4357(.A(n9382), .B(g531), .Y(n9405));
AOI21X1  g4358(.A0(n9405), .A1(n9364), .B0(n9387), .Y(n9406));
OAI21X1  g4359(.A0(n9404), .A1(n9383), .B0(n9406), .Y(n9407));
NAND2X1  g4360(.A(n9407), .B(n9393), .Y(n7882));
AOI21X1  g4361(.A0(n9372), .A1(n9366), .B0(n6323), .Y(n9409));
XOR2X1   g4362(.A(n9409), .B(n6045), .Y(n9410));
NAND2X1  g4363(.A(n9410), .B(n9401), .Y(n9411));
NOR2X1   g4364(.A(n9382), .B(g532), .Y(n9412));
AOI21X1  g4365(.A0(n9412), .A1(n9364), .B0(n9387), .Y(n9413));
OAI21X1  g4366(.A0(n9411), .A1(n9383), .B0(n9413), .Y(n9414));
NAND2X1  g4367(.A(n9414), .B(n9381), .Y(n7887));
INVX1    g4368(.A(n9380), .Y(n9416));
NAND2X1  g4369(.A(n9373), .B(n6319_1), .Y(n9417));
XOR2X1   g4370(.A(n9417), .B(n6053), .Y(n9418));
NAND2X1  g4371(.A(n9418), .B(n9401), .Y(n9419));
NOR2X1   g4372(.A(n9382), .B(g533), .Y(n9420));
AOI21X1  g4373(.A0(n9420), .A1(n9364), .B0(n9387), .Y(n9421));
OAI21X1  g4374(.A0(n9419), .A1(n9383), .B0(n9421), .Y(n9422));
OAI21X1  g4375(.A0(n9416), .A1(n9364), .B0(n9422), .Y(n7892));
INVX1    g4376(.A(n9401), .Y(n9424));
AOI21X1  g4377(.A0(n9372), .A1(n9366), .B0(n6342), .Y(n9425));
XOR2X1   g4378(.A(n9425), .B(n6046_1), .Y(n9426));
NOR3X1   g4379(.A(n9426), .B(n9424), .C(n9383), .Y(n9427));
NOR3X1   g4380(.A(n9382), .B(n9392), .C(g534), .Y(n9428));
OR2X1    g4381(.A(n9428), .B(n9387), .Y(n9429));
OAI22X1  g4382(.A0(n9427), .A1(n9429), .B0(n9416), .B1(n9364), .Y(n7897));
AOI21X1  g4383(.A0(n9372), .A1(n9366), .B0(n6338), .Y(n9431));
XOR2X1   g4384(.A(n9431), .B(n6053), .Y(n9432));
NOR2X1   g4385(.A(n9432), .B(n9424), .Y(n9433));
NAND2X1  g4386(.A(n9373), .B(n6333), .Y(n9434));
XOR2X1   g4387(.A(n9434), .B(n6053), .Y(n9435));
NAND2X1  g4388(.A(n9435), .B(n9401), .Y(n9436));
NOR2X1   g4389(.A(n9382), .B(g536), .Y(n9437));
AOI21X1  g4390(.A0(n9437), .A1(n9364), .B0(n9387), .Y(n9438));
OAI21X1  g4391(.A0(n9436), .A1(n9383), .B0(n9438), .Y(n9439));
OAI21X1  g4392(.A0(n9433), .A1(n9416), .B0(n9439), .Y(n7902));
AOI21X1  g4393(.A0(n9372), .A1(n9366), .B0(n6305), .Y(n9441));
XOR2X1   g4394(.A(n9441), .B(n6046_1), .Y(n9442));
NOR2X1   g4395(.A(n9442), .B(n9424), .Y(n9443));
AOI21X1  g4396(.A0(n9372), .A1(n9366), .B0(n6328), .Y(n9444));
XOR2X1   g4397(.A(n9444), .B(n6046_1), .Y(n9445));
NOR3X1   g4398(.A(n9445), .B(n9424), .C(n9383), .Y(n9446));
NOR3X1   g4399(.A(n9382), .B(n9392), .C(g537), .Y(n9447));
OR2X1    g4400(.A(n9447), .B(n9387), .Y(n9448));
OAI22X1  g4401(.A0(n9446), .A1(n9448), .B0(n9443), .B1(n9416), .Y(n7907));
NOR2X1   g4402(.A(n9445), .B(n9424), .Y(n9450));
XOR2X1   g4403(.A(n9450), .B(n9436), .Y(n9451));
NOR2X1   g4404(.A(n9426), .B(n9424), .Y(n9452));
XOR2X1   g4405(.A(n9452), .B(n9419), .Y(n9453));
XOR2X1   g4406(.A(n9453), .B(n9451), .Y(n9454));
XOR2X1   g4407(.A(n9411), .B(n9404), .Y(n9455));
AND2X1   g4408(.A(n9395), .B(n9401), .Y(n9456));
XOR2X1   g4409(.A(n9456), .B(n9386), .Y(n9457));
XOR2X1   g4410(.A(n9457), .B(n9455), .Y(n9458));
XOR2X1   g4411(.A(n9458), .B(n9454), .Y(n9459));
NOR2X1   g4412(.A(g541), .B(g3229), .Y(n9460));
NOR3X1   g4413(.A(n9460), .B(g510), .C(g557), .Y(n9461));
OAI21X1  g4414(.A0(g538), .A1(n5718), .B0(n9461), .Y(n9462));
NOR4X1   g4415(.A(n9382), .B(n9387), .C(n9392), .D(n9462), .Y(n9463));
XOR2X1   g4416(.A(n9443), .B(n9433), .Y(n9464));
AOI21X1  g4417(.A0(n9464), .A1(g557), .B0(n9463), .Y(n9465));
OAI21X1  g4418(.A0(n9459), .A1(n6176), .B0(n9465), .Y(n7912));
NOR3X1   g4419(.A(n3905), .B(g1245), .C(g1249), .Y(n9467));
OR4X1    g4420(.A(n7310), .B(n7307_1), .C(n7306), .D(n7311), .Y(n9468));
NOR3X1   g4421(.A(n9468), .B(n7304), .C(n7300), .Y(n9469));
NAND2X1  g4422(.A(n7332), .B(n7327), .Y(n9470));
NOR2X1   g4423(.A(g1424), .B(n7296), .Y(n9471));
OAI22X1  g4424(.A0(g1425), .A1(n7298_1), .B0(n7215_1), .B1(g1423), .Y(n9472));
OR2X1    g4425(.A(n9472), .B(n9471), .Y(n9473));
NAND4X1  g4426(.A(n7348), .B(n7322), .C(n7318), .D(n9473), .Y(n9474));
NOR4X1   g4427(.A(n9470), .B(n7341), .C(n7337), .D(n9474), .Y(n9475));
NAND2X1  g4428(.A(n9475), .B(n9469), .Y(n9476));
NOR2X1   g4429(.A(g1422), .B(n7298_1), .Y(n9477));
OAI22X1  g4430(.A0(g1421), .A1(n7296), .B0(n7215_1), .B1(g1420), .Y(n9478));
NOR2X1   g4431(.A(n9478), .B(n9477), .Y(n9479));
AOI21X1  g4432(.A0(n9479), .A1(n9476), .B0(n5304), .Y(n9480));
NAND2X1  g4433(.A(n9480), .B(n9467), .Y(n9481));
INVX1    g4434(.A(g1243), .Y(n9482));
NOR2X1   g4435(.A(g1196), .B(n9482), .Y(n9483));
NAND2X1  g4436(.A(n9483), .B(n9481), .Y(n9484));
OAI21X1  g4437(.A0(g1211), .A1(g1243), .B0(n7174_1), .Y(n9485));
INVX1    g4438(.A(n9485), .Y(n9486));
XOR2X1   g4439(.A(n7308), .B(n7051), .Y(n9488));
NOR4X1   g4440(.A(g1245), .B(n5304), .C(g1249), .D(n3905), .Y(n9489));
NAND2X1  g4441(.A(n9489), .B(n9488), .Y(n9490));
OAI21X1  g4442(.A0(g1211), .A1(g1196), .B0(n9482), .Y(n9491));
NOR2X1   g4443(.A(n9485), .B(g1215), .Y(n9492));
AOI21X1  g4444(.A0(n9492), .A1(n9467), .B0(n9491), .Y(n9493));
OAI21X1  g4445(.A0(n9490), .A1(n9486), .B0(n9493), .Y(n9494));
NAND2X1  g4446(.A(n9494), .B(n9484), .Y(n7917));
INVX1    g4447(.A(n9467), .Y(n9496));
OAI21X1  g4448(.A0(n9480), .A1(n9496), .B0(n9483), .Y(n9497));
INVX1    g4449(.A(n9489), .Y(n9498));
XOR2X1   g4450(.A(n7300), .B(n7046), .Y(n9500));
NOR3X1   g4451(.A(n9500), .B(n9498), .C(n9486), .Y(n9501));
NOR3X1   g4452(.A(n9485), .B(n9496), .C(g1216), .Y(n9502));
OR2X1    g4453(.A(n9502), .B(n9491), .Y(n9503));
OAI21X1  g4454(.A0(n9503), .A1(n9501), .B0(n9497), .Y(n7922));
AOI21X1  g4455(.A0(n9475), .A1(n9469), .B0(n7312_1), .Y(n9505));
XOR2X1   g4456(.A(n9505), .B(n7051), .Y(n9506));
NOR3X1   g4457(.A(n9506), .B(n9498), .C(n9486), .Y(n9507));
NOR3X1   g4458(.A(n9485), .B(n9496), .C(g1217), .Y(n9508));
OR2X1    g4459(.A(n9508), .B(n9491), .Y(n9509));
OAI21X1  g4460(.A0(n9509), .A1(n9507), .B0(n9497), .Y(n7927));
AOI21X1  g4461(.A0(n9475), .A1(n9469), .B0(n7322), .Y(n9511));
XOR2X1   g4462(.A(n9511), .B(n7046), .Y(n9512));
OR4X1    g4463(.A(n9486), .B(n9496), .C(n5304), .D(n9512), .Y(n9513));
NOR2X1   g4464(.A(n9485), .B(g1218), .Y(n9514));
AOI21X1  g4465(.A0(n9514), .A1(n9467), .B0(n9491), .Y(n9515));
NAND2X1  g4466(.A(n9515), .B(n9513), .Y(n9516));
NAND2X1  g4467(.A(n9516), .B(n9484), .Y(n7932));
INVX1    g4468(.A(n9483), .Y(n9518));
NAND2X1  g4469(.A(n9476), .B(n7318), .Y(n9519));
XOR2X1   g4470(.A(n9519), .B(n7051), .Y(n9520));
NAND2X1  g4471(.A(n9520), .B(n9489), .Y(n9521));
NOR2X1   g4472(.A(n9485), .B(g1219), .Y(n9522));
AOI21X1  g4473(.A0(n9522), .A1(n9467), .B0(n9491), .Y(n9523));
OAI21X1  g4474(.A0(n9521), .A1(n9486), .B0(n9523), .Y(n9524));
OAI21X1  g4475(.A0(n9518), .A1(n9467), .B0(n9524), .Y(n7937));
AOI21X1  g4476(.A0(n9475), .A1(n9469), .B0(n7341), .Y(n9526));
XOR2X1   g4477(.A(n9526), .B(n7046), .Y(n9527));
NOR3X1   g4478(.A(n9527), .B(n9498), .C(n9486), .Y(n9528));
NOR3X1   g4479(.A(n9485), .B(n9496), .C(g1220), .Y(n9529));
OR2X1    g4480(.A(n9529), .B(n9491), .Y(n9530));
OAI22X1  g4481(.A0(n9528), .A1(n9530), .B0(n9518), .B1(n9467), .Y(n7942));
AOI21X1  g4482(.A0(n9475), .A1(n9469), .B0(n7337), .Y(n9532));
XOR2X1   g4483(.A(n9532), .B(n7051), .Y(n9533));
NOR2X1   g4484(.A(n9533), .B(n9498), .Y(n9534));
NAND2X1  g4485(.A(n9476), .B(n7332), .Y(n9535));
XOR2X1   g4486(.A(n9535), .B(n7051), .Y(n9536));
NAND2X1  g4487(.A(n9536), .B(n9489), .Y(n9537));
NOR2X1   g4488(.A(n9485), .B(g1222), .Y(n9538));
AOI21X1  g4489(.A0(n9538), .A1(n9467), .B0(n9491), .Y(n9539));
OAI21X1  g4490(.A0(n9537), .A1(n9486), .B0(n9539), .Y(n9540));
OAI21X1  g4491(.A0(n9534), .A1(n9518), .B0(n9540), .Y(n7947));
AOI21X1  g4492(.A0(n9475), .A1(n9469), .B0(n7304), .Y(n9542));
XOR2X1   g4493(.A(n9542), .B(n7046), .Y(n9543));
NOR2X1   g4494(.A(n9543), .B(n9498), .Y(n9544));
AOI21X1  g4495(.A0(n9475), .A1(n9469), .B0(n7327), .Y(n9545));
XOR2X1   g4496(.A(n9545), .B(n7046), .Y(n9546));
NOR3X1   g4497(.A(n9546), .B(n9498), .C(n9486), .Y(n9547));
NOR3X1   g4498(.A(n9485), .B(n9496), .C(g1223), .Y(n9548));
OR2X1    g4499(.A(n9548), .B(n9491), .Y(n9549));
OAI22X1  g4500(.A0(n9547), .A1(n9549), .B0(n9544), .B1(n9518), .Y(n7952));
NOR2X1   g4501(.A(n9546), .B(n9498), .Y(n9551));
XOR2X1   g4502(.A(n9551), .B(n9537), .Y(n9552));
NOR2X1   g4503(.A(n9527), .B(n9498), .Y(n9553));
XOR2X1   g4504(.A(n9553), .B(n9521), .Y(n9554));
XOR2X1   g4505(.A(n9554), .B(n9552), .Y(n9555));
NOR2X1   g4506(.A(n9506), .B(n9498), .Y(n9556));
NOR2X1   g4507(.A(n9512), .B(n9498), .Y(n9557));
XOR2X1   g4508(.A(n9557), .B(n9556), .Y(n9558));
NOR2X1   g4509(.A(n9500), .B(n9498), .Y(n9559));
XOR2X1   g4510(.A(n9559), .B(n9490), .Y(n9560));
XOR2X1   g4511(.A(n9560), .B(n9558), .Y(n9561));
XOR2X1   g4512(.A(n9561), .B(n9555), .Y(n9562));
NOR2X1   g4513(.A(g1224), .B(n5718), .Y(n9563));
NOR2X1   g4514(.A(g1196), .B(g1243), .Y(n9564));
OAI21X1  g4515(.A0(g1227), .A1(g3229), .B0(n9564), .Y(n9565));
NOR4X1   g4516(.A(n9563), .B(n9485), .C(n9491), .D(n9565), .Y(n9566));
XOR2X1   g4517(.A(n9544), .B(n9534), .Y(n9567));
AOI22X1  g4518(.A0(n9566), .A1(n9467), .B0(g1243), .B1(n9567), .Y(n9568));
OAI21X1  g4519(.A0(n9562), .A1(n7174_1), .B0(n9568), .Y(n7957));
NOR2X1   g4520(.A(g1939), .B(g1943), .Y(n9570));
OAI21X1  g4521(.A0(n5318), .A1(n5317), .B0(n9570), .Y(n9571));
NOR3X1   g4522(.A(n8302), .B(n8297), .C(n8295), .Y(n9572));
NOR4X1   g4523(.A(n8308), .B(n8305), .C(n8304), .D(n8309), .Y(n9573));
AND2X1   g4524(.A(n9573), .B(n9572), .Y(n9574));
OAI21X1  g4525(.A0(n8327), .A1(n8326), .B0(n8324), .Y(n9575));
NOR2X1   g4526(.A(g2118), .B(n8294), .Y(n9576));
OAI22X1  g4527(.A0(g2119), .A1(n8296), .B0(n8213), .B1(g2117), .Y(n9577));
OR2X1    g4528(.A(n9577), .B(n9576), .Y(n9578));
NAND4X1  g4529(.A(n8344), .B(n8319), .C(n8315), .D(n9578), .Y(n9579));
NOR4X1   g4530(.A(n9575), .B(n8337), .C(n8333), .D(n9579), .Y(n9580));
NOR2X1   g4531(.A(g2116), .B(n8296), .Y(n9581));
OAI22X1  g4532(.A0(g2115), .A1(n8294), .B0(n8213), .B1(g2114), .Y(n9582));
NOR2X1   g4533(.A(n9582), .B(n9581), .Y(n9583));
INVX1    g4534(.A(n9583), .Y(n9584));
AOI21X1  g4535(.A0(n9580), .A1(n9574), .B0(n9584), .Y(n9585));
NOR3X1   g4536(.A(n9585), .B(n9571), .C(n5315), .Y(n9586));
INVX1    g4537(.A(g1937), .Y(n9587));
NOR2X1   g4538(.A(g1890), .B(n9587), .Y(n9588));
INVX1    g4539(.A(n9588), .Y(n9589));
OAI21X1  g4540(.A0(g1905), .A1(g1937), .B0(n8172), .Y(n9590));
INVX1    g4541(.A(n9590), .Y(n9591));
XOR2X1   g4542(.A(n8306), .B(n8048), .Y(n9592));
NOR4X1   g4543(.A(n9591), .B(n9571), .C(n5315), .D(n9592), .Y(n9593));
OAI21X1  g4544(.A0(g1905), .A1(g1890), .B0(n9587), .Y(n9594));
INVX1    g4545(.A(n9594), .Y(n9595));
OR2X1    g4546(.A(n9590), .B(g1909), .Y(n9596));
OAI21X1  g4547(.A0(n9596), .A1(n9571), .B0(n9595), .Y(n9597));
OAI22X1  g4548(.A0(n9593), .A1(n9597), .B0(n9589), .B1(n9586), .Y(n7962));
NOR2X1   g4549(.A(n9585), .B(n5315), .Y(n9599));
OAI21X1  g4550(.A0(n9599), .A1(n9571), .B0(n9588), .Y(n9600));
XOR2X1   g4551(.A(n8298), .B(n8043), .Y(n9601));
NOR4X1   g4552(.A(n9591), .B(n9571), .C(n5315), .D(n9601), .Y(n9602));
OR2X1    g4553(.A(n9590), .B(g1910), .Y(n9603));
OAI21X1  g4554(.A0(n9603), .A1(n9571), .B0(n9595), .Y(n9604));
OAI21X1  g4555(.A0(n9604), .A1(n9602), .B0(n9600), .Y(n7967));
AOI21X1  g4556(.A0(n9580), .A1(n9574), .B0(n8310), .Y(n9606));
XOR2X1   g4557(.A(n9606), .B(n8049), .Y(n9607));
NOR4X1   g4558(.A(n9591), .B(n9571), .C(n5315), .D(n9607), .Y(n9608));
OR2X1    g4559(.A(n9590), .B(g1911), .Y(n9609));
OAI21X1  g4560(.A0(n9609), .A1(n9571), .B0(n9595), .Y(n9610));
OAI21X1  g4561(.A0(n9610), .A1(n9608), .B0(n9600), .Y(n7972));
AOI21X1  g4562(.A0(n9580), .A1(n9574), .B0(n8319), .Y(n9612));
XOR2X1   g4563(.A(n9612), .B(n8044), .Y(n9613));
NOR4X1   g4564(.A(n9591), .B(n9571), .C(n5315), .D(n9613), .Y(n9614));
OR2X1    g4565(.A(n9590), .B(g1912), .Y(n9615));
OAI21X1  g4566(.A0(n9615), .A1(n9571), .B0(n9595), .Y(n9616));
OAI22X1  g4567(.A0(n9614), .A1(n9616), .B0(n9589), .B1(n9586), .Y(n7977));
INVX1    g4568(.A(n9571), .Y(n9618));
INVX1    g4569(.A(n8315), .Y(n9619));
AOI21X1  g4570(.A0(n9580), .A1(n9574), .B0(n9619), .Y(n9620));
XOR2X1   g4571(.A(n9620), .B(n8049), .Y(n9621));
NOR4X1   g4572(.A(n9591), .B(n9571), .C(n5315), .D(n9621), .Y(n9622));
OR2X1    g4573(.A(n9590), .B(g1913), .Y(n9623));
OAI21X1  g4574(.A0(n9623), .A1(n9571), .B0(n9595), .Y(n9624));
OAI22X1  g4575(.A0(n9622), .A1(n9624), .B0(n9589), .B1(n9618), .Y(n7982));
AOI21X1  g4576(.A0(n9580), .A1(n9574), .B0(n8337), .Y(n9626));
XOR2X1   g4577(.A(n9626), .B(n8044), .Y(n9627));
NOR4X1   g4578(.A(n9591), .B(n9571), .C(n5315), .D(n9627), .Y(n9628));
OR2X1    g4579(.A(n9590), .B(g1914), .Y(n9629));
OAI21X1  g4580(.A0(n9629), .A1(n9571), .B0(n9595), .Y(n9630));
OAI22X1  g4581(.A0(n9628), .A1(n9630), .B0(n9589), .B1(n9618), .Y(n7987));
AOI21X1  g4582(.A0(n9580), .A1(n9574), .B0(n8333), .Y(n9632));
XOR2X1   g4583(.A(n9632), .B(n8049), .Y(n9633));
NOR3X1   g4584(.A(n9633), .B(n9571), .C(n5315), .Y(n9634));
AOI21X1  g4585(.A0(n9580), .A1(n9574), .B0(n8328), .Y(n9635));
XOR2X1   g4586(.A(n9635), .B(n8049), .Y(n9636));
NOR4X1   g4587(.A(n9591), .B(n9571), .C(n5315), .D(n9636), .Y(n9637));
OR2X1    g4588(.A(n9590), .B(g1916), .Y(n9638));
OAI21X1  g4589(.A0(n9638), .A1(n9571), .B0(n9595), .Y(n9639));
OAI22X1  g4590(.A0(n9637), .A1(n9639), .B0(n9634), .B1(n9589), .Y(n7992));
AOI21X1  g4591(.A0(n9580), .A1(n9574), .B0(n8302), .Y(n9641));
XOR2X1   g4592(.A(n9641), .B(n8044), .Y(n9642));
NOR3X1   g4593(.A(n9642), .B(n9571), .C(n5315), .Y(n9643));
AOI21X1  g4594(.A0(n9580), .A1(n9574), .B0(n8324), .Y(n9644));
XOR2X1   g4595(.A(n9644), .B(n8044), .Y(n9645));
NOR4X1   g4596(.A(n9591), .B(n9571), .C(n5315), .D(n9645), .Y(n9646));
OR2X1    g4597(.A(n9590), .B(g1917), .Y(n9647));
OAI21X1  g4598(.A0(n9647), .A1(n9571), .B0(n9595), .Y(n9648));
OAI22X1  g4599(.A0(n9646), .A1(n9648), .B0(n9643), .B1(n9589), .Y(n7997));
NOR3X1   g4600(.A(n9636), .B(n9571), .C(n5315), .Y(n9650));
NOR3X1   g4601(.A(n9645), .B(n9571), .C(n5315), .Y(n9651));
XOR2X1   g4602(.A(n9651), .B(n9650), .Y(n9652));
NOR3X1   g4603(.A(n9621), .B(n9571), .C(n5315), .Y(n9653));
NOR3X1   g4604(.A(n9627), .B(n9571), .C(n5315), .Y(n9654));
XOR2X1   g4605(.A(n9654), .B(n9653), .Y(n9655));
XOR2X1   g4606(.A(n9655), .B(n9652), .Y(n9656));
NOR3X1   g4607(.A(n9607), .B(n9571), .C(n5315), .Y(n9657));
NOR3X1   g4608(.A(n9613), .B(n9571), .C(n5315), .Y(n9658));
XOR2X1   g4609(.A(n9658), .B(n9657), .Y(n9659));
INVX1    g4610(.A(n9570), .Y(n9660));
OR4X1    g4611(.A(n9660), .B(n5606), .C(n5315), .D(n9592), .Y(n9661));
NOR3X1   g4612(.A(n9601), .B(n9571), .C(n5315), .Y(n9662));
XOR2X1   g4613(.A(n9662), .B(n9661), .Y(n9663));
XOR2X1   g4614(.A(n9663), .B(n9659), .Y(n9664));
XOR2X1   g4615(.A(n9664), .B(n9656), .Y(n9665));
NOR2X1   g4616(.A(g1921), .B(g3229), .Y(n9666));
NOR3X1   g4617(.A(n9666), .B(g1890), .C(g1937), .Y(n9667));
OAI21X1  g4618(.A0(g1918), .A1(n5718), .B0(n9667), .Y(n9668));
NOR4X1   g4619(.A(n9590), .B(n9594), .C(n9571), .D(n9668), .Y(n9669));
XOR2X1   g4620(.A(n9643), .B(n9634), .Y(n9670));
AOI21X1  g4621(.A0(n9670), .A1(g1937), .B0(n9669), .Y(n9671));
OAI21X1  g4622(.A0(n9665), .A1(n8172), .B0(n9671), .Y(n8002));
NOR3X1   g4623(.A(n5318), .B(n5317), .C(n5326), .Y(n9673));
INVX1    g4624(.A(n5327), .Y(n9674));
OAI22X1  g4625(.A0(n9673), .A1(n9674), .B0(n5328), .B1(g2618), .Y(n9675));
NOR2X1   g4626(.A(g2633), .B(g2637), .Y(n9676));
OR4X1    g4627(.A(n9303), .B(n9300), .C(n9299), .D(n9304), .Y(n9677));
NOR3X1   g4628(.A(n9677), .B(n9297), .C(n9293), .Y(n9678));
NAND2X1  g4629(.A(n9325), .B(n9320), .Y(n9679));
NOR2X1   g4630(.A(g2812), .B(n9289), .Y(n9680));
OAI22X1  g4631(.A0(g2813), .A1(n9291), .B0(n9208), .B1(g2811), .Y(n9681));
OR2X1    g4632(.A(n9681), .B(n9680), .Y(n9682));
NAND4X1  g4633(.A(n9341), .B(n9315), .C(n9311), .D(n9682), .Y(n9683));
NOR4X1   g4634(.A(n9679), .B(n9334), .C(n9330), .D(n9683), .Y(n9684));
NAND2X1  g4635(.A(n9684), .B(n9678), .Y(n9685));
NOR2X1   g4636(.A(g2810), .B(n9291), .Y(n9686));
OAI22X1  g4637(.A0(g2809), .A1(n9289), .B0(n9208), .B1(g2808), .Y(n9687));
NOR2X1   g4638(.A(n9687), .B(n9686), .Y(n9688));
AOI21X1  g4639(.A0(n9688), .A1(n9685), .B0(n5328), .Y(n9689));
NAND3X1  g4640(.A(n9689), .B(n9676), .C(n9675), .Y(n9690));
INVX1    g4641(.A(g2631), .Y(n9691));
NOR2X1   g4642(.A(g2584), .B(n9691), .Y(n9692));
NAND2X1  g4643(.A(n9692), .B(n9690), .Y(n9693));
OAI21X1  g4644(.A0(g2599), .A1(g2631), .B0(n9168), .Y(n9694));
INVX1    g4645(.A(n9694), .Y(n9695));
XOR2X1   g4646(.A(n9301), .B(n9045), .Y(n9697));
NAND4X1  g4647(.A(n9676), .B(n9675), .C(g2574), .D(n9697), .Y(n9698));
NOR2X1   g4648(.A(n9698), .B(n9695), .Y(n9699));
INVX1    g4649(.A(n9676), .Y(n9700));
NOR2X1   g4650(.A(n9700), .B(n7307), .Y(n9701));
INVX1    g4651(.A(n9701), .Y(n9702));
OAI21X1  g4652(.A0(g2599), .A1(g2584), .B0(n9691), .Y(n9703));
INVX1    g4653(.A(n9703), .Y(n9704));
OR2X1    g4654(.A(n9694), .B(g2603), .Y(n9705));
OAI21X1  g4655(.A0(n9705), .A1(n9702), .B0(n9704), .Y(n9706));
OAI21X1  g4656(.A0(n9706), .A1(n9699), .B0(n9693), .Y(n8007));
OAI21X1  g4657(.A0(n9689), .A1(n9702), .B0(n9692), .Y(n9708));
XOR2X1   g4658(.A(n9293), .B(n9040), .Y(n9710));
NOR4X1   g4659(.A(n9700), .B(n7307), .C(n5328), .D(n9710), .Y(n9711));
AND2X1   g4660(.A(n9711), .B(n9694), .Y(n9712));
OR2X1    g4661(.A(n9694), .B(g2604), .Y(n9713));
OAI21X1  g4662(.A0(n9713), .A1(n9702), .B0(n9704), .Y(n9714));
OAI21X1  g4663(.A0(n9714), .A1(n9712), .B0(n9708), .Y(n8012));
AOI21X1  g4664(.A0(n9684), .A1(n9678), .B0(n9305), .Y(n9716));
XOR2X1   g4665(.A(n9716), .B(n9045), .Y(n9717));
NOR4X1   g4666(.A(n9700), .B(n7307), .C(n5328), .D(n9717), .Y(n9718));
AND2X1   g4667(.A(n9718), .B(n9694), .Y(n9719));
OR2X1    g4668(.A(n9694), .B(g2605), .Y(n9720));
OAI21X1  g4669(.A0(n9720), .A1(n9702), .B0(n9704), .Y(n9721));
OAI21X1  g4670(.A0(n9721), .A1(n9719), .B0(n9708), .Y(n8017));
AOI21X1  g4671(.A0(n9684), .A1(n9678), .B0(n9315), .Y(n9723));
XOR2X1   g4672(.A(n9723), .B(n9040), .Y(n9724));
NOR4X1   g4673(.A(n9700), .B(n7307), .C(n5328), .D(n9724), .Y(n9725));
AND2X1   g4674(.A(n9725), .B(n9694), .Y(n9726));
OR2X1    g4675(.A(n9694), .B(g2606), .Y(n9727));
OAI21X1  g4676(.A0(n9727), .A1(n9702), .B0(n9704), .Y(n9728));
OAI21X1  g4677(.A0(n9728), .A1(n9726), .B0(n9693), .Y(n8022));
INVX1    g4678(.A(n9692), .Y(n9730));
NAND2X1  g4679(.A(n9685), .B(n9311), .Y(n9731));
XOR2X1   g4680(.A(n9731), .B(n9045), .Y(n9732));
NAND4X1  g4681(.A(n9676), .B(n9675), .C(g2574), .D(n9732), .Y(n9733));
NOR2X1   g4682(.A(n9733), .B(n9695), .Y(n9734));
OR2X1    g4683(.A(n9694), .B(g2607), .Y(n9735));
OAI21X1  g4684(.A0(n9735), .A1(n9702), .B0(n9704), .Y(n9736));
OAI22X1  g4685(.A0(n9734), .A1(n9736), .B0(n9730), .B1(n9701), .Y(n8027));
AOI21X1  g4686(.A0(n9684), .A1(n9678), .B0(n9334), .Y(n9738));
XOR2X1   g4687(.A(n9738), .B(n9040), .Y(n9739));
NOR4X1   g4688(.A(n9700), .B(n7307), .C(n5328), .D(n9739), .Y(n9740));
AND2X1   g4689(.A(n9740), .B(n9694), .Y(n9741));
OR2X1    g4690(.A(n9694), .B(g2608), .Y(n9742));
OAI21X1  g4691(.A0(n9742), .A1(n9702), .B0(n9704), .Y(n9743));
OAI22X1  g4692(.A0(n9741), .A1(n9743), .B0(n9730), .B1(n9701), .Y(n8032));
AOI21X1  g4693(.A0(n9684), .A1(n9678), .B0(n9330), .Y(n9745));
XOR2X1   g4694(.A(n9745), .B(n9045), .Y(n9746));
NOR4X1   g4695(.A(n9700), .B(n7307), .C(n5328), .D(n9746), .Y(n9747));
NAND2X1  g4696(.A(n9685), .B(n9325), .Y(n9748));
XOR2X1   g4697(.A(n9748), .B(n9045), .Y(n9749));
NAND4X1  g4698(.A(n9676), .B(n9675), .C(g2574), .D(n9749), .Y(n9750));
NOR2X1   g4699(.A(n9750), .B(n9695), .Y(n9751));
OR2X1    g4700(.A(n9694), .B(g2610), .Y(n9752));
OAI21X1  g4701(.A0(n9752), .A1(n9702), .B0(n9704), .Y(n9753));
OAI22X1  g4702(.A0(n9751), .A1(n9753), .B0(n9747), .B1(n9730), .Y(n8037));
AOI21X1  g4703(.A0(n9684), .A1(n9678), .B0(n9297), .Y(n9755));
XOR2X1   g4704(.A(n9755), .B(n9040), .Y(n9756));
NOR4X1   g4705(.A(n9700), .B(n7307), .C(n5328), .D(n9756), .Y(n9757));
AOI21X1  g4706(.A0(n9684), .A1(n9678), .B0(n9320), .Y(n9758));
XOR2X1   g4707(.A(n9758), .B(n9040), .Y(n9759));
NOR4X1   g4708(.A(n9700), .B(n7307), .C(n5328), .D(n9759), .Y(n9760));
AND2X1   g4709(.A(n9760), .B(n9694), .Y(n9761));
OR2X1    g4710(.A(n9694), .B(g2611), .Y(n9762));
OAI21X1  g4711(.A0(n9762), .A1(n9702), .B0(n9704), .Y(n9763));
OAI22X1  g4712(.A0(n9761), .A1(n9763), .B0(n9757), .B1(n9730), .Y(n8042));
XOR2X1   g4713(.A(n9760), .B(n9750), .Y(n9765));
XOR2X1   g4714(.A(n9740), .B(n9733), .Y(n9766));
XOR2X1   g4715(.A(n9766), .B(n9765), .Y(n9767));
XOR2X1   g4716(.A(n9725), .B(n9718), .Y(n9768));
XOR2X1   g4717(.A(n9711), .B(n9698), .Y(n9769));
XOR2X1   g4718(.A(n9769), .B(n9768), .Y(n9770));
XOR2X1   g4719(.A(n9770), .B(n9767), .Y(n9771));
NOR2X1   g4720(.A(g2612), .B(n5718), .Y(n9772));
NOR2X1   g4721(.A(g2584), .B(g2631), .Y(n9773));
OAI21X1  g4722(.A0(g2615), .A1(g3229), .B0(n9773), .Y(n9774));
NOR4X1   g4723(.A(n9772), .B(n9694), .C(n9703), .D(n9774), .Y(n9775));
XOR2X1   g4724(.A(n9757), .B(n9747), .Y(n9776));
AOI22X1  g4725(.A0(n9775), .A1(n9701), .B0(g2631), .B1(n9776), .Y(n9777));
OAI21X1  g4726(.A0(n9771), .A1(n9168), .B0(n9777), .Y(n8047));
NOR2X1   g4727(.A(n5976_1), .B(n9358), .Y(n9779));
NOR2X1   g4728(.A(n9779), .B(g3234), .Y(n9780));
XOR2X1   g4729(.A(g2993), .B(g3080), .Y(n9781));
MX2X1    g4730(.A(n9360), .B(n9781), .S0(n9780), .Y(n8052));
AND2X1   g4731(.A(g2993), .B(g3080), .Y(n9783));
XOR2X1   g4732(.A(n9783), .B(n5970), .Y(n9784));
OAI21X1  g4733(.A0(n9784), .A1(n9779), .B0(n9360), .Y(n8057));
NAND3X1  g4734(.A(g2998), .B(g2993), .C(g3080), .Y(n9786));
XOR2X1   g4735(.A(n9786), .B(g3006), .Y(n9787));
NOR3X1   g4736(.A(n9787), .B(n9779), .C(g3234), .Y(n8062));
NAND4X1  g4737(.A(g2998), .B(g2993), .C(g3080), .D(g3006), .Y(n9789));
XOR2X1   g4738(.A(n9789), .B(g3002), .Y(n9790));
NOR3X1   g4739(.A(n9790), .B(n9779), .C(g3234), .Y(n8067));
NOR2X1   g4740(.A(n9789), .B(n5972), .Y(n9792));
XOR2X1   g4741(.A(n9792), .B(n5973), .Y(n9793));
NOR3X1   g4742(.A(n9793), .B(n9779), .C(g3234), .Y(n8072));
INVX1    g4743(.A(g3010), .Y(n9795));
NOR3X1   g4744(.A(n9789), .B(n5973), .C(n5972), .Y(n9796));
XOR2X1   g4745(.A(n9796), .B(n9795), .Y(n9797));
NOR3X1   g4746(.A(n9797), .B(n9779), .C(g3234), .Y(n8077));
NOR4X1   g4747(.A(n9795), .B(n5973), .C(n5972), .D(n9789), .Y(n9799));
XOR2X1   g4748(.A(n9799), .B(n5974), .Y(n9800));
NOR3X1   g4749(.A(n9800), .B(n9779), .C(g3234), .Y(n8082));
INVX1    g4750(.A(g3036), .Y(n9802));
NOR3X1   g4751(.A(n5976_1), .B(n5977), .C(n9358), .Y(n9803));
NAND4X1  g4752(.A(g3032), .B(n9802), .C(n5978), .D(n9803), .Y(n9804));
XOR2X1   g4753(.A(n9779), .B(n5977), .Y(n9805));
NAND3X1  g4754(.A(n9805), .B(n9804), .C(n9360), .Y(n8087));
AND2X1   g4755(.A(n9804), .B(n9360), .Y(n9807));
XOR2X1   g4756(.A(n9803), .B(g3028), .Y(n9808));
AND2X1   g4757(.A(n9808), .B(n9807), .Y(n8092));
NOR4X1   g4758(.A(n5978), .B(n5977), .C(n9358), .D(n5976_1), .Y(n9810));
XOR2X1   g4759(.A(n9810), .B(g3036), .Y(n9811));
AND2X1   g4760(.A(n9811), .B(n9807), .Y(n8097));
AND2X1   g4761(.A(n9810), .B(g3036), .Y(n9813));
XOR2X1   g4762(.A(n9813), .B(g3032), .Y(n9814));
AND2X1   g4763(.A(n9814), .B(n9807), .Y(n8102));
MX2X1    g4764(.A(g3043), .B(g3062), .S0(g2987), .Y(n8121));
MX2X1    g4765(.A(g3044), .B(g3063), .S0(g2987), .Y(n8126));
MX2X1    g4766(.A(g3045), .B(g3064), .S0(g2987), .Y(n8131));
MX2X1    g4767(.A(g3046), .B(g3065), .S0(g2987), .Y(n8136));
MX2X1    g4768(.A(g3047), .B(g3066), .S0(g2987), .Y(n8141));
MX2X1    g4769(.A(g3048), .B(g3067), .S0(g2987), .Y(n8146));
MX2X1    g4770(.A(g3049), .B(g3068), .S0(g2987), .Y(n8151));
MX2X1    g4771(.A(g3050), .B(g3069), .S0(g2987), .Y(n8156));
MX2X1    g4772(.A(g3051), .B(g3070), .S0(g2987), .Y(n8161));
XOR2X1   g4773(.A(g36), .B(g33), .Y(n9825));
XOR2X1   g4774(.A(g30), .B(g27), .Y(n9826));
XOR2X1   g4775(.A(n9826), .B(n9825), .Y(n9827));
XOR2X1   g4776(.A(g39), .B(g42), .Y(n9828));
XOR2X1   g4777(.A(g45), .B(g48), .Y(n9829));
XOR2X1   g4778(.A(n9829), .B(n9828), .Y(n9830));
XOR2X1   g4779(.A(n9830), .B(n9827), .Y(n9831));
AND2X1   g4780(.A(g3136), .B(n5251), .Y(n9832));
XOR2X1   g4781(.A(n9832), .B(n9831), .Y(n8166));
XOR2X1   g4782(.A(n9831), .B(g3083), .Y(n8171));
MX2X1    g4783(.A(g3052), .B(g3071), .S0(g2987), .Y(n8176));
MX2X1    g4784(.A(g3053), .B(g3072), .S0(g2987), .Y(n8181));
MX2X1    g4785(.A(g3055), .B(g3073), .S0(g2987), .Y(n8186));
MX2X1    g4786(.A(g3056), .B(g3074), .S0(g2987), .Y(n8191));
MX2X1    g4787(.A(g3057), .B(g3075), .S0(g2987), .Y(n8196));
MX2X1    g4788(.A(g3058), .B(g3076), .S0(g2987), .Y(n8201));
MX2X1    g4789(.A(g3059), .B(g3077), .S0(g2987), .Y(n8206));
MX2X1    g4790(.A(g3060), .B(g3078), .S0(g2987), .Y(n8211));
MX2X1    g4791(.A(g3061), .B(g2997), .S0(g2987), .Y(n8216));
XOR2X1   g4792(.A(g2), .B(g8), .Y(n9844));
XOR2X1   g4793(.A(g5), .B(g14), .Y(n9845));
XOR2X1   g4794(.A(n9845), .B(n9844), .Y(n9846));
XOR2X1   g4795(.A(g11), .B(g17), .Y(n9847));
XOR2X1   g4796(.A(g20), .B(g23), .Y(n9848));
XOR2X1   g4797(.A(n9848), .B(n9847), .Y(n9849));
XOR2X1   g4798(.A(n9849), .B(n9846), .Y(n9850));
XOR2X1   g4799(.A(n9850), .B(g2990), .Y(n8221));
XOR2X1   g4800(.A(n9850), .B(n9832), .Y(n8226));
BUFX1    g4801(.A(g2848), .Y(g3993));
BUFX1    g4802(.A(g2836), .Y(g4088));
BUFX1    g4803(.A(g2864), .Y(g4090));
BUFX1    g4804(.A(g2851), .Y(g4200));
BUFX1    g4805(.A(g2839), .Y(g4321));
BUFX1    g4806(.A(g2867), .Y(g4323));
BUFX1    g4807(.A(g2854), .Y(g4450));
BUFX1    g4808(.A(g2870), .Y(g4590));
BUFX1    g4809(.A(g3040), .Y(g5388));
BUFX1    g4810(.A(g276), .Y(g5437));
BUFX1    g4811(.A(g963), .Y(g5472));
BUFX1    g4812(.A(g1657), .Y(g5511));
BUFX1    g4813(.A(g182), .Y(g5549));
BUFX1    g4814(.A(g2351), .Y(g5555));
BUFX1    g4815(.A(g870), .Y(g5595));
BUFX1    g4816(.A(g1564), .Y(g5612));
BUFX1    g4817(.A(g325), .Y(g5629));
BUFX1    g4818(.A(g2258), .Y(g5637));
BUFX1    g4819(.A(g331), .Y(g5648));
BUFX1    g4820(.A(g1012), .Y(g5657));
BUFX1    g4821(.A(g1018), .Y(g5686));
BUFX1    g4822(.A(g1706), .Y(g5695));
BUFX1    g4823(.A(g1712), .Y(g5738));
BUFX1    g4824(.A(g2400), .Y(g5747));
BUFX1    g4825(.A(g2406), .Y(g5796));
BUFX1    g4826(.A(g2818), .Y(g6225));
BUFX1    g4827(.A(g138), .Y(g6231));
BUFX1    g4828(.A(g135), .Y(g6313));
BUFX1    g4829(.A(g826), .Y(g6368));
BUFX1    g4830(.A(g2821), .Y(g6442));
BUFX1    g4831(.A(g405), .Y(g6447));
BUFX1    g4832(.A(g545), .Y(g6485));
BUFX1    g4833(.A(g823), .Y(g6518));
BUFX1    g4834(.A(g1520), .Y(g6573));
BUFX1    g4835(.A(g551), .Y(g6642));
BUFX1    g4836(.A(g623), .Y(g6677));
BUFX1    g4837(.A(g1092), .Y(g6712));
BUFX1    g4838(.A(g1231), .Y(g6750));
BUFX1    g4839(.A(g1517), .Y(g6782));
BUFX1    g4840(.A(g2214), .Y(g6837));
BUFX1    g4841(.A(g2824), .Y(g6895));
BUFX1    g4842(.A(g626), .Y(g6911));
BUFX1    g4843(.A(g1237), .Y(g6944));
BUFX1    g4844(.A(g1309), .Y(g6979));
BUFX1    g4845(.A(g1786), .Y(g7014));
BUFX1    g4846(.A(g1925), .Y(g7052));
BUFX1    g4847(.A(g2211), .Y(g7084));
BUFX1    g4848(.A(g1312), .Y(g7161));
BUFX1    g4849(.A(g1931), .Y(g7194));
BUFX1    g4850(.A(g2003), .Y(g7229));
BUFX1    g4851(.A(g2480), .Y(g7264));
BUFX1    g4852(.A(g2619), .Y(g7302));
BUFX1    g4853(.A(g2827), .Y(g7334));
BUFX1    g4854(.A(g2006), .Y(g7357));
BUFX1    g4855(.A(g2625), .Y(g7390));
BUFX1    g4856(.A(g2697), .Y(g7425));
BUFX1    g4857(.A(g2700), .Y(g7487));
BUFX1    g4858(.A(g2830), .Y(g7519));
BUFX1    g4859(.A(g474), .Y(g7909));
BUFX1    g4860(.A(g481), .Y(g7956));
BUFX1    g4861(.A(g1161), .Y(g7961));
BUFX1    g4862(.A(g1168), .Y(g8007));
BUFX1    g4863(.A(g1855), .Y(g8012));
BUFX1    g4864(.A(g2930), .Y(g8021));
BUFX1    g4865(.A(g2842), .Y(g8023));
BUFX1    g4866(.A(g3117), .Y(g8030));
BUFX1    g4867(.A(g1862), .Y(g8082));
BUFX1    g4868(.A(g2549), .Y(g8087));
BUFX1    g4869(.A(g2858), .Y(g8096));
BUFX1    g4870(.A(g3129), .Y(g8106));
BUFX1    g4871(.A(g2556), .Y(g8167));
BUFX1    g4872(.A(g2845), .Y(g8175));
BUFX1    g4873(.A(g2833), .Y(g8249));
BUFX1    g4874(.A(g2861), .Y(g8251));
BUFX1    g4875(.A(g1), .Y(g8258));
BUFX1    g4876(.A(g2), .Y(g8259));
BUFX1    g4877(.A(g5), .Y(g8260));
BUFX1    g4878(.A(g8), .Y(g8261));
BUFX1    g4879(.A(g11), .Y(g8262));
BUFX1    g4880(.A(g14), .Y(g8263));
BUFX1    g4881(.A(g17), .Y(g8264));
BUFX1    g4882(.A(g20), .Y(g8265));
BUFX1    g4883(.A(g23), .Y(g8266));
BUFX1    g4884(.A(g26), .Y(g8267));
BUFX1    g4885(.A(g27), .Y(g8268));
BUFX1    g4886(.A(g30), .Y(g8269));
BUFX1    g4887(.A(g33), .Y(g8270));
BUFX1    g4888(.A(g36), .Y(g8271));
BUFX1    g4889(.A(g39), .Y(g8272));
BUFX1    g4890(.A(g42), .Y(g8273));
BUFX1    g4891(.A(g45), .Y(g8274));
BUFX1    g4892(.A(g48), .Y(g8275));
BUFX1    g4893(.A(g520), .Y(g16297));
BUFX1    g4894(.A(g1206), .Y(g16355));
BUFX1    g4895(.A(g1900), .Y(g16399));
BUFX1    g4896(.A(g2594), .Y(g16437));
BUFX1    g4897(.A(g51), .Y(n269));
BUFX1    g4898(.A(g51), .Y(n354));
BUFX1    g4899(.A(g2930), .Y(n358));
BUFX1    g4900(.A(g3212), .Y(n368));
BUFX1    g4901(.A(g3228), .Y(n373));
BUFX1    g4902(.A(g3227), .Y(n378));
BUFX1    g4903(.A(g3226), .Y(n383));
BUFX1    g4904(.A(g3225), .Y(n388));
BUFX1    g4905(.A(g3224), .Y(n393));
BUFX1    g4906(.A(g3223), .Y(n398));
BUFX1    g4907(.A(g3222), .Y(n403));
BUFX1    g4908(.A(g3221), .Y(n408));
BUFX1    g4909(.A(g3232), .Y(n413));
BUFX1    g4910(.A(g3220), .Y(n418));
BUFX1    g4911(.A(g3219), .Y(n423));
BUFX1    g4912(.A(g3218), .Y(n428));
BUFX1    g4913(.A(g3217), .Y(n433));
BUFX1    g4914(.A(g3216), .Y(n438));
BUFX1    g4915(.A(g3215), .Y(n443));
BUFX1    g4916(.A(g3214), .Y(n448));
BUFX1    g4917(.A(g3213), .Y(n453));
BUFX1    g4918(.A(g2861), .Y(n507));
BUFX1    g4919(.A(g2864), .Y(n516));
BUFX1    g4920(.A(g2867), .Y(n525));
BUFX1    g4921(.A(g2870), .Y(n534));
BUFX1    g4922(.A(g2818), .Y(n543));
BUFX1    g4923(.A(g2821), .Y(n552));
BUFX1    g4924(.A(g2824), .Y(n561));
BUFX1    g4925(.A(g2827), .Y(n570));
BUFX1    g4926(.A(g2830), .Y(n579));
BUFX1    g4927(.A(g2833), .Y(n588));
BUFX1    g4928(.A(g2836), .Y(n597));
BUFX1    g4929(.A(g2839), .Y(n606));
BUFX1    g4930(.A(g2842), .Y(n615));
BUFX1    g4931(.A(g2845), .Y(n624));
BUFX1    g4932(.A(g2848), .Y(n633));
BUFX1    g4933(.A(g2851), .Y(n642));
BUFX1    g4934(.A(g2854), .Y(n651));
BUFX1    g4935(.A(g2858), .Y(n660));
BUFX1    g4936(.A(g3080), .Y(n710));
BUFX1    g4937(.A(g3129), .Y(n714));
BUFX1    g4938(.A(g3117), .Y(n718));
OAI21X1  g4939(.A0(n5051), .A1(g3123), .B0(n5045), .Y(n903));
NAND2X1  g4940(.A(n5062), .B(n5045), .Y(n908));
INVX1    g4941(.A(n968), .Y(n913));
NAND2X1  g4942(.A(n5056), .B(n5045), .Y(n918));
NAND3X1  g4943(.A(n5163), .B(n5153), .C(n5045), .Y(n923));
INVX1    g4944(.A(n953), .Y(n928));
OR4X1    g4945(.A(n5096), .B(n5084_1), .C(n5076), .D(n5118), .Y(n933));
INVX1    g4946(.A(n943), .Y(n938));
OR4X1    g4947(.A(n5096), .B(n5084_1), .C(n5076), .D(n5118), .Y(n948));
NAND3X1  g4948(.A(n5163), .B(n5153), .C(n5045), .Y(n958));
NAND2X1  g4949(.A(n5056), .B(n5045), .Y(n963));
NAND2X1  g4950(.A(n5062), .B(n5045), .Y(n973));
OR4X1    g4951(.A(n5096), .B(n5084_1), .C(n5076), .D(n5118), .Y(n983));
INVX1    g4952(.A(n953), .Y(n988));
NAND3X1  g4953(.A(n5163), .B(n5153), .C(n5045), .Y(n993));
NAND2X1  g4954(.A(n5056), .B(n5045), .Y(n998));
INVX1    g4955(.A(n968), .Y(n1003));
NAND2X1  g4956(.A(n5062), .B(n5045), .Y(n1008));
INVX1    g4957(.A(n943), .Y(n1013));
OR4X1    g4958(.A(n5096), .B(n5084_1), .C(n5076), .D(n5118), .Y(n1018));
INVX1    g4959(.A(n953), .Y(n1023));
NAND3X1  g4960(.A(n5163), .B(n5153), .C(n5045), .Y(n1028));
INVX1    g4961(.A(n943), .Y(n1033));
OR4X1    g4962(.A(n5096), .B(n5084_1), .C(n5076), .D(n5118), .Y(n1038));
INVX1    g4963(.A(n953), .Y(n1043));
NOR4X1   g4964(.A(n5173), .B(n5168), .C(n5076), .D(n5174_1), .Y(n1048));
BUFX1    g4965(.A(g2950), .Y(n1053));
BUFX1    g4966(.A(g138), .Y(n1057));
BUFX1    g4967(.A(g135), .Y(n1061));
BUFX1    g4968(.A(g180), .Y(n1480));
BUFX1    g4969(.A(g182), .Y(n1484));
BUFX1    g4970(.A(g2950), .Y(n1489));
BUFX1    g4971(.A(g276), .Y(n1493));
BUFX1    g4972(.A(g405), .Y(n1497));
BUFX1    g4973(.A(g182), .Y(n1502));
BUFX1    g4974(.A(g450), .Y(n1736));
BUFX1    g4975(.A(g452), .Y(n1745));
BUFX1    g4976(.A(g454), .Y(n1754));
BUFX1    g4977(.A(g280), .Y(n1763));
BUFX1    g4978(.A(g282), .Y(n1772));
BUFX1    g4979(.A(g284), .Y(n1781));
BUFX1    g4980(.A(g286), .Y(n1790));
BUFX1    g4981(.A(g288), .Y(n1799));
BUFX1    g4982(.A(g2857), .Y(n1804));
BUFX1    g4983(.A(g290), .Y(n1808));
BUFX1    g4984(.A(g354), .Y(n1878));
BUFX1    g4985(.A(g342), .Y(n1882));
BUFX1    g4986(.A(g343), .Y(n1887));
BUFX1    g4987(.A(g350), .Y(n1891));
BUFX1    g4988(.A(g346), .Y(n1896));
BUFX1    g4989(.A(g352), .Y(n1900));
BUFX1    g4990(.A(g369), .Y(n1905));
BUFX1    g4991(.A(g357), .Y(n1909));
BUFX1    g4992(.A(g358), .Y(n1914));
BUFX1    g4993(.A(g365), .Y(n1918));
BUFX1    g4994(.A(g361), .Y(n1923));
BUFX1    g4995(.A(g367), .Y(n1927));
BUFX1    g4996(.A(g384), .Y(n1932));
BUFX1    g4997(.A(g372), .Y(n1936));
BUFX1    g4998(.A(g373), .Y(n1941));
BUFX1    g4999(.A(g380), .Y(n1945));
BUFX1    g5000(.A(g376), .Y(n1950));
BUFX1    g5001(.A(g382), .Y(n1954));
BUFX1    g5002(.A(g398), .Y(n1959));
BUFX1    g5003(.A(g387), .Y(n1963));
BUFX1    g5004(.A(g388), .Y(n1968));
BUFX1    g5005(.A(g395), .Y(n1972));
BUFX1    g5006(.A(g391), .Y(n1977));
BUFX1    g5007(.A(g397), .Y(n1981));
BUFX1    g5008(.A(g3080), .Y(n1986));
BUFX1    g5009(.A(g325), .Y(n1990));
BUFX1    g5010(.A(g331), .Y(n1994));
BUFX1    g5011(.A(g3080), .Y(n1999));
BUFX1    g5012(.A(g545), .Y(n2003));
BUFX1    g5013(.A(g551), .Y(n2007));
BUFX1    g5014(.A(g513), .Y(n2031));
BUFX1    g5015(.A(g523), .Y(n2035));
BUFX1    g5016(.A(g455), .Y(n2040));
BUFX1    g5017(.A(g564), .Y(n2044));
BUFX1    g5018(.A(g458), .Y(n2049));
BUFX1    g5019(.A(g570), .Y(n2053));
BUFX1    g5020(.A(g461), .Y(n2058));
BUFX1    g5021(.A(g572), .Y(n2062));
BUFX1    g5022(.A(g465), .Y(n2067));
BUFX1    g5023(.A(g574), .Y(n2071));
BUFX1    g5024(.A(g468), .Y(n2076));
BUFX1    g5025(.A(g566), .Y(n2080));
BUFX1    g5026(.A(g471), .Y(n2085));
BUFX1    g5027(.A(g568), .Y(n2089));
BUFX1    g5028(.A(g2950), .Y(n2094));
BUFX1    g5029(.A(g474), .Y(n2098));
BUFX1    g5030(.A(g481), .Y(n2102));
BUFX1    g5031(.A(g528), .Y(n2186));
BUFX1    g5032(.A(g535), .Y(n2190));
BUFX1    g5033(.A(g543), .Y(n2199));
BUFX1    g5034(.A(g549), .Y(n2213));
BUFX1    g5035(.A(g558), .Y(n2222));
BUFX1    g5036(.A(g499), .Y(n2362));
BUFX1    g5037(.A(g520), .Y(n2416));
BUFX1    g5038(.A(g3080), .Y(n2471));
BUFX1    g5039(.A(g623), .Y(n2475));
BUFX1    g5040(.A(g626), .Y(n2479));
BUFX1    g5041(.A(g2950), .Y(n2754));
BUFX1    g5042(.A(g826), .Y(n2758));
BUFX1    g5043(.A(g823), .Y(n2762));
AND2X1   g5044(.A(n5401_1), .B(n5399), .Y(n3177));
BUFX1    g5045(.A(g868), .Y(n3181));
BUFX1    g5046(.A(g870), .Y(n3185));
BUFX1    g5047(.A(g2950), .Y(n3190));
BUFX1    g5048(.A(g963), .Y(n3194));
BUFX1    g5049(.A(g1092), .Y(n3198));
BUFX1    g5050(.A(g870), .Y(n3203));
BUFX1    g5051(.A(g1137), .Y(n3437));
BUFX1    g5052(.A(g1139), .Y(n3446));
BUFX1    g5053(.A(g1141), .Y(n3455));
BUFX1    g5054(.A(g967), .Y(n3464));
BUFX1    g5055(.A(g969), .Y(n3473));
BUFX1    g5056(.A(g971), .Y(n3482));
BUFX1    g5057(.A(g973), .Y(n3491));
BUFX1    g5058(.A(g975), .Y(n3500));
BUFX1    g5059(.A(g2873), .Y(n3505));
BUFX1    g5060(.A(g977), .Y(n3509));
BUFX1    g5061(.A(g1041), .Y(n3579));
BUFX1    g5062(.A(g1029), .Y(n3583));
BUFX1    g5063(.A(g1030), .Y(n3588));
BUFX1    g5064(.A(g1037), .Y(n3592));
BUFX1    g5065(.A(g1033), .Y(n3597));
BUFX1    g5066(.A(g1039), .Y(n3601));
BUFX1    g5067(.A(g1056), .Y(n3606));
BUFX1    g5068(.A(g1044), .Y(n3610));
BUFX1    g5069(.A(g1045), .Y(n3615));
BUFX1    g5070(.A(g1052), .Y(n3619));
BUFX1    g5071(.A(g1048), .Y(n3624));
BUFX1    g5072(.A(g1054), .Y(n3628));
BUFX1    g5073(.A(g1071), .Y(n3633));
BUFX1    g5074(.A(g1059), .Y(n3637));
BUFX1    g5075(.A(g1060), .Y(n3642));
BUFX1    g5076(.A(g1067), .Y(n3646));
BUFX1    g5077(.A(g1063), .Y(n3651));
BUFX1    g5078(.A(g1069), .Y(n3655));
BUFX1    g5079(.A(g1085), .Y(n3660));
BUFX1    g5080(.A(g1074), .Y(n3664));
BUFX1    g5081(.A(g1075), .Y(n3669));
BUFX1    g5082(.A(g1082), .Y(n3673));
BUFX1    g5083(.A(g1078), .Y(n3678));
BUFX1    g5084(.A(g1084), .Y(n3682));
BUFX1    g5085(.A(g3080), .Y(n3687));
BUFX1    g5086(.A(g1012), .Y(n3691));
BUFX1    g5087(.A(g1018), .Y(n3695));
BUFX1    g5088(.A(g3080), .Y(n3700));
BUFX1    g5089(.A(g1231), .Y(n3704));
BUFX1    g5090(.A(g1237), .Y(n3708));
BUFX1    g5091(.A(g1199), .Y(n3732));
BUFX1    g5092(.A(g1209), .Y(n3736));
BUFX1    g5093(.A(g1142), .Y(n3741));
BUFX1    g5094(.A(g1250), .Y(n3745));
BUFX1    g5095(.A(g1145), .Y(n3750));
BUFX1    g5096(.A(g1256), .Y(n3754));
BUFX1    g5097(.A(g1148), .Y(n3759));
BUFX1    g5098(.A(g1258), .Y(n3763));
BUFX1    g5099(.A(g1152), .Y(n3768));
BUFX1    g5100(.A(g1260), .Y(n3772));
BUFX1    g5101(.A(g1155), .Y(n3777));
BUFX1    g5102(.A(g1252), .Y(n3781));
BUFX1    g5103(.A(g1158), .Y(n3786));
BUFX1    g5104(.A(g1254), .Y(n3790));
BUFX1    g5105(.A(g2950), .Y(n3795));
BUFX1    g5106(.A(g1161), .Y(n3799));
BUFX1    g5107(.A(g1168), .Y(n3803));
BUFX1    g5108(.A(g1214), .Y(n3887));
BUFX1    g5109(.A(g1221), .Y(n3891));
BUFX1    g5110(.A(g1229), .Y(n3900));
BUFX1    g5111(.A(g1235), .Y(n3914));
BUFX1    g5112(.A(g1244), .Y(n3923));
BUFX1    g5113(.A(g1186), .Y(n4063));
BUFX1    g5114(.A(g1206), .Y(n4117));
BUFX1    g5115(.A(g3080), .Y(n4172));
BUFX1    g5116(.A(g1309), .Y(n4176));
BUFX1    g5117(.A(g1312), .Y(n4180));
BUFX1    g5118(.A(g2950), .Y(n4455));
BUFX1    g5119(.A(g1520), .Y(n4459));
BUFX1    g5120(.A(g1517), .Y(n4463));
AND2X1   g5121(.A(n5401_1), .B(n5399), .Y(n4878));
BUFX1    g5122(.A(g1562), .Y(n4882));
BUFX1    g5123(.A(g1564), .Y(n4886));
BUFX1    g5124(.A(g2950), .Y(n4891));
BUFX1    g5125(.A(g1657), .Y(n4895));
BUFX1    g5126(.A(g1786), .Y(n4899));
BUFX1    g5127(.A(g1564), .Y(n4904));
BUFX1    g5128(.A(g1831), .Y(n5138));
BUFX1    g5129(.A(g1833), .Y(n5147));
BUFX1    g5130(.A(g1835), .Y(n5156));
BUFX1    g5131(.A(g1661), .Y(n5165));
BUFX1    g5132(.A(g1663), .Y(n5174));
BUFX1    g5133(.A(g1665), .Y(n5183));
BUFX1    g5134(.A(g1667), .Y(n5192));
BUFX1    g5135(.A(g1669), .Y(n5201));
BUFX1    g5136(.A(g2877), .Y(n5206));
BUFX1    g5137(.A(g1671), .Y(n5210));
BUFX1    g5138(.A(g1735), .Y(n5280));
BUFX1    g5139(.A(g1723), .Y(n5284));
BUFX1    g5140(.A(g1724), .Y(n5289));
BUFX1    g5141(.A(g1731), .Y(n5293));
BUFX1    g5142(.A(g1727), .Y(n5298));
BUFX1    g5143(.A(g1733), .Y(n5302));
BUFX1    g5144(.A(g1750), .Y(n5307));
BUFX1    g5145(.A(g1738), .Y(n5311));
BUFX1    g5146(.A(g1739), .Y(n5316));
BUFX1    g5147(.A(g1746), .Y(n5320));
BUFX1    g5148(.A(g1742), .Y(n5325));
BUFX1    g5149(.A(g1748), .Y(n5329));
BUFX1    g5150(.A(g1765), .Y(n5334));
BUFX1    g5151(.A(g1753), .Y(n5338));
BUFX1    g5152(.A(g1754), .Y(n5343));
BUFX1    g5153(.A(g1761), .Y(n5347));
BUFX1    g5154(.A(g1757), .Y(n5352));
BUFX1    g5155(.A(g1763), .Y(n5356));
BUFX1    g5156(.A(g1779), .Y(n5361));
BUFX1    g5157(.A(g1768), .Y(n5365));
BUFX1    g5158(.A(g1769), .Y(n5370));
BUFX1    g5159(.A(g1776), .Y(n5374));
BUFX1    g5160(.A(g1772), .Y(n5379));
BUFX1    g5161(.A(g1778), .Y(n5383));
BUFX1    g5162(.A(g3080), .Y(n5388));
BUFX1    g5163(.A(g1706), .Y(n5392));
BUFX1    g5164(.A(g1712), .Y(n5396));
BUFX1    g5165(.A(g3080), .Y(n5401));
BUFX1    g5166(.A(g1925), .Y(n5405));
BUFX1    g5167(.A(g1931), .Y(n5409));
BUFX1    g5168(.A(g1893), .Y(n5433));
BUFX1    g5169(.A(g1903), .Y(n5437));
BUFX1    g5170(.A(g1836), .Y(n5442));
BUFX1    g5171(.A(g1944), .Y(n5446));
BUFX1    g5172(.A(g1839), .Y(n5451));
BUFX1    g5173(.A(g1950), .Y(n5455));
BUFX1    g5174(.A(g1842), .Y(n5460));
BUFX1    g5175(.A(g1952), .Y(n5464));
BUFX1    g5176(.A(g1846), .Y(n5469));
BUFX1    g5177(.A(g1954), .Y(n5473));
BUFX1    g5178(.A(g1849), .Y(n5478));
BUFX1    g5179(.A(g1946), .Y(n5482));
BUFX1    g5180(.A(g1852), .Y(n5487));
BUFX1    g5181(.A(g1948), .Y(n5491));
BUFX1    g5182(.A(g2950), .Y(n5496));
BUFX1    g5183(.A(g1855), .Y(n5500));
BUFX1    g5184(.A(g1862), .Y(n5504));
BUFX1    g5185(.A(g1908), .Y(n5588));
BUFX1    g5186(.A(g1915), .Y(n5592));
BUFX1    g5187(.A(g1923), .Y(n5601));
BUFX1    g5188(.A(g1929), .Y(n5615));
BUFX1    g5189(.A(g1938), .Y(n5624));
BUFX1    g5190(.A(g1880), .Y(n5764));
BUFX1    g5191(.A(g1900), .Y(n5818));
BUFX1    g5192(.A(g3080), .Y(n5873));
BUFX1    g5193(.A(g2003), .Y(n5877));
BUFX1    g5194(.A(g2006), .Y(n5881));
BUFX1    g5195(.A(g2950), .Y(n6156));
BUFX1    g5196(.A(g2214), .Y(n6160));
BUFX1    g5197(.A(g2211), .Y(n6164));
AND2X1   g5198(.A(n5401_1), .B(n5399), .Y(n6579));
BUFX1    g5199(.A(g2256), .Y(n6583));
BUFX1    g5200(.A(g2258), .Y(n6587));
BUFX1    g5201(.A(g2950), .Y(n6592));
BUFX1    g5202(.A(g2351), .Y(n6596));
BUFX1    g5203(.A(g2480), .Y(n6600));
BUFX1    g5204(.A(g2258), .Y(n6605));
BUFX1    g5205(.A(g2525), .Y(n6839));
BUFX1    g5206(.A(g2527), .Y(n6848));
BUFX1    g5207(.A(g2529), .Y(n6857));
BUFX1    g5208(.A(g2355), .Y(n6866));
BUFX1    g5209(.A(g2357), .Y(n6875));
BUFX1    g5210(.A(g2359), .Y(n6884));
BUFX1    g5211(.A(g2361), .Y(n6893));
BUFX1    g5212(.A(g2363), .Y(n6902));
BUFX1    g5213(.A(g2878), .Y(n6907));
BUFX1    g5214(.A(g2365), .Y(n6911));
BUFX1    g5215(.A(g2429), .Y(n6981));
BUFX1    g5216(.A(g2417), .Y(n6985));
BUFX1    g5217(.A(g2418), .Y(n6990));
BUFX1    g5218(.A(g2425), .Y(n6994));
BUFX1    g5219(.A(g2421), .Y(n6999));
BUFX1    g5220(.A(g2427), .Y(n7003));
BUFX1    g5221(.A(g2444), .Y(n7008));
BUFX1    g5222(.A(g2432), .Y(n7012));
BUFX1    g5223(.A(g2433), .Y(n7017));
BUFX1    g5224(.A(g2440), .Y(n7021));
BUFX1    g5225(.A(g2436), .Y(n7026));
BUFX1    g5226(.A(g2442), .Y(n7030));
BUFX1    g5227(.A(g2459), .Y(n7035));
BUFX1    g5228(.A(g2447), .Y(n7039));
BUFX1    g5229(.A(g2448), .Y(n7044));
BUFX1    g5230(.A(g2455), .Y(n7048));
BUFX1    g5231(.A(g2451), .Y(n7053));
BUFX1    g5232(.A(g2457), .Y(n7057));
BUFX1    g5233(.A(g2473), .Y(n7062));
BUFX1    g5234(.A(g2462), .Y(n7066));
BUFX1    g5235(.A(g2463), .Y(n7071));
BUFX1    g5236(.A(g2470), .Y(n7075));
BUFX1    g5237(.A(g2466), .Y(n7080));
BUFX1    g5238(.A(g2472), .Y(n7084));
BUFX1    g5239(.A(g3080), .Y(n7089));
BUFX1    g5240(.A(g2400), .Y(n7093));
BUFX1    g5241(.A(g2406), .Y(n7097));
BUFX1    g5242(.A(g3080), .Y(n7102));
BUFX1    g5243(.A(g2619), .Y(n7106));
BUFX1    g5244(.A(g2625), .Y(n7110));
BUFX1    g5245(.A(g2587), .Y(n7134));
BUFX1    g5246(.A(g2597), .Y(n7138));
BUFX1    g5247(.A(g2530), .Y(n7143));
BUFX1    g5248(.A(g2638), .Y(n7147));
BUFX1    g5249(.A(g2533), .Y(n7152));
BUFX1    g5250(.A(g2644), .Y(n7156));
BUFX1    g5251(.A(g2536), .Y(n7161));
BUFX1    g5252(.A(g2646), .Y(n7165));
BUFX1    g5253(.A(g2540), .Y(n7170));
BUFX1    g5254(.A(g2648), .Y(n7174));
BUFX1    g5255(.A(g2543), .Y(n7179));
BUFX1    g5256(.A(g2640), .Y(n7183));
BUFX1    g5257(.A(g2546), .Y(n7188));
BUFX1    g5258(.A(g2642), .Y(n7192));
BUFX1    g5259(.A(g2950), .Y(n7197));
BUFX1    g5260(.A(g2549), .Y(n7201));
BUFX1    g5261(.A(g2556), .Y(n7205));
BUFX1    g5262(.A(g2602), .Y(n7289));
BUFX1    g5263(.A(g2609), .Y(n7293));
BUFX1    g5264(.A(g2617), .Y(n7302));
BUFX1    g5265(.A(g2623), .Y(n7316));
BUFX1    g5266(.A(g2632), .Y(n7325));
BUFX1    g5267(.A(g2574), .Y(n7465));
BUFX1    g5268(.A(g2594), .Y(n7519));
BUFX1    g5269(.A(g3080), .Y(n7574));
BUFX1    g5270(.A(g2697), .Y(n7578));
BUFX1    g5271(.A(g2700), .Y(n7582));
BUFX1    g5272(.A(g3234), .Y(n8107));
BUFX1    g5273(.A(g3040), .Y(n8111));
OAI21X1  g5274(.A0(g2986), .A1(n5042), .B0(g2987), .Y(n8116));
endmodule
