//Converted to Combinational , Module name: s953 , Timestamp: 2018-12-03T15:51:02.154841 
module s953 ( Rdy1RtHS1, Rdy2RtHS1, Rdy1BmHS1, Rdy2BmHS1, InDoneHS1, RtTSHS1, TpArrayHS1, OutputHS1, WantBmHS1, WantRtHS1, OutAvHS1, FullOHS1, FullIHS1, Prog_2, Prog_1, Prog_0, State_5, State_4, State_3, State_2, State_1, State_0, ReWhBufHS1, TgWhBufHS1, SeOutAvHS1, LdProgHS1, Mode2HS1, ReRtTSHS1, ShftIRHS1, NewTrHS1, Mode1HS1, ShftORHS1, ActRtHS1, Mode0HS1, TxHInHS1, LxHInHS1, NewLineHS1, ActBmHS1, GoBmHS1, LoadOHHS1, DumpIHS1, SeFullOHS1, GoRtHS1, LoadIHHS1, SeFullIHS1, n79, n84, n89, n94, n99, n104 );
input Rdy1RtHS1, Rdy2RtHS1, Rdy1BmHS1, Rdy2BmHS1, InDoneHS1, RtTSHS1, TpArrayHS1, OutputHS1, WantBmHS1, WantRtHS1, OutAvHS1, FullOHS1, FullIHS1, Prog_2, Prog_1, Prog_0, State_5, State_4, State_3, State_2, State_1, State_0;
output ReWhBufHS1, TgWhBufHS1, SeOutAvHS1, LdProgHS1, Mode2HS1, ReRtTSHS1, ShftIRHS1, NewTrHS1, Mode1HS1, ShftORHS1, ActRtHS1, Mode0HS1, TxHInHS1, LxHInHS1, NewLineHS1, ActBmHS1, GoBmHS1, LoadOHHS1, DumpIHS1, SeFullOHS1, GoRtHS1, LoadIHHS1, SeFullIHS1, n79, n84, n89, n94, n99, n104;
wire n126, n127, n128, n129_1, n130, n131, n132, n133_1, n134, n135, n136, n137_1, n138, n139, n140, n141_1, n142, n143, n144, n145_1, n146, n147, n148, n149_1, n150, n151, n152, n153_1, n154, n155, n156, n157_1, n158, n159, n160, n161_1, n162, n164, n165_1, n167, n168, n169_1, n170, n171, n172, n173_1, n174, n175, n176, n177_1, n178, n179, n180, n181_1, n182, n183, n185_1, n186, n187, n188, n189_1, n190, n191, n192, n193_1, n194, n195, n196, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n253, n254, n255, n256, n257, n258, n259, n261, n262, n263, n264, n265, n267, n268, n269, n270, n271, n272, n273, n274, n275, n277, n278, n279, n280, n281, n282, n283, n284, n286, n289, n290, n291, n293, n295, n296, n297, n298, n299, n300, n301, n303, n304, n305, n306, n307, n310, n311, n312, n313, n314, n315, n316, n317, n318, n320, n321, n322, n323, n324, n325, n326, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n343, n344, n345, n346, n347, n348, n349, n350, n353, n354, n355, n356, n358, n359, n363, n365;
INVX1    g000(.A(Rdy1RtHS1), .Y(n126));
INVX1    g001(.A(State_3), .Y(n127));
INVX1    g002(.A(State_2), .Y(n128));
NAND3X1  g003(.A(n128), .B(n127), .C(State_5), .Y(n129_1));
NOR3X1   g004(.A(n129_1), .B(State_4), .C(Rdy1BmHS1), .Y(n130));
INVX1    g005(.A(Prog_2), .Y(n131));
INVX1    g006(.A(State_1), .Y(n132));
NAND4X1  g007(.A(n128), .B(n127), .C(State_5), .D(n132), .Y(n133_1));
NOR3X1   g008(.A(n133_1), .B(State_0), .C(n131), .Y(n134));
INVX1    g009(.A(State_0), .Y(n135));
NOR2X1   g010(.A(FullIHS1), .B(FullOHS1), .Y(n136));
NOR4X1   g011(.A(n129_1), .B(n135), .C(State_4), .D(n136), .Y(n137_1));
XOR2X1   g012(.A(State_0), .B(State_1), .Y(n138));
INVX1    g013(.A(State_5), .Y(n139));
NOR3X1   g014(.A(n128), .B(State_3), .C(n139), .Y(n140));
AND2X1   g015(.A(n140), .B(n138), .Y(n141_1));
NAND2X1  g016(.A(n127), .B(State_5), .Y(n142));
XOR2X1   g017(.A(State_0), .B(n132), .Y(n143));
NOR4X1   g018(.A(n142), .B(State_4), .C(Prog_2), .D(n143), .Y(n144));
OR4X1    g019(.A(n141_1), .B(n137_1), .C(n134), .D(n144), .Y(n145_1));
AOI21X1  g020(.A0(n130), .A1(n126), .B0(n145_1), .Y(n146));
INVX1    g021(.A(Rdy1BmHS1), .Y(n147));
INVX1    g022(.A(Rdy2BmHS1), .Y(n148));
NAND2X1  g023(.A(State_0), .B(n132), .Y(n149_1));
OAI22X1  g024(.A0(n133_1), .A1(Prog_0), .B0(n142), .B1(n149_1), .Y(n150));
OAI21X1  g025(.A0(n148), .A1(n147), .B0(n150), .Y(n151));
AND2X1   g026(.A(Rdy2RtHS1), .B(Rdy1RtHS1), .Y(n152));
NOR4X1   g027(.A(State_2), .B(State_3), .C(n139), .D(State_0), .Y(n153_1));
NOR4X1   g028(.A(n132), .B(State_3), .C(n139), .D(State_0), .Y(n154));
AOI21X1  g029(.A0(n153_1), .A1(Prog_0), .B0(n154), .Y(n155));
OR2X1    g030(.A(n155), .B(n152), .Y(n156));
NOR2X1   g031(.A(Prog_1), .B(Prog_2), .Y(n157_1));
NOR2X1   g032(.A(State_4), .B(State_5), .Y(n158));
NAND3X1  g033(.A(n158), .B(n135), .C(State_2), .Y(n159));
NAND3X1  g034(.A(n132), .B(n127), .C(RtTSHS1), .Y(n160));
NOR3X1   g035(.A(n160), .B(n159), .C(n157_1), .Y(n161_1));
INVX1    g036(.A(State_4), .Y(n162));
NOR3X1   g037(.A(n133_1), .B(State_0), .C(n162), .Y(Mode2HS1));
NOR4X1   g038(.A(n129_1), .B(State_4), .C(n131), .D(n136), .Y(n164));
NOR3X1   g039(.A(n164), .B(Mode2HS1), .C(n161_1), .Y(n165_1));
NAND4X1  g040(.A(n156), .B(n151), .C(n146), .D(n165_1), .Y(n79));
NAND2X1  g041(.A(n136), .B(n162), .Y(n167));
NOR4X1   g042(.A(n133_1), .B(State_0), .C(n131), .D(n167), .Y(n168));
INVX1    g043(.A(WantBmHS1), .Y(n169_1));
AOI21X1  g044(.A0(n148), .A1(Rdy1BmHS1), .B0(n169_1), .Y(n170));
INVX1    g045(.A(n170), .Y(n171));
NAND4X1  g046(.A(n168), .B(Prog_0), .C(Rdy2RtHS1), .D(n171), .Y(n172));
OAI21X1  g047(.A0(Rdy2RtHS1), .A1(n126), .B0(WantRtHS1), .Y(n173_1));
INVX1    g048(.A(Prog_1), .Y(n174));
XOR2X1   g049(.A(Prog_0), .B(n174), .Y(n175));
OAI21X1  g050(.A0(n175), .A1(n148), .B0(n170), .Y(n176));
NAND3X1  g051(.A(n176), .B(n173_1), .C(n168), .Y(n177_1));
INVX1    g052(.A(Rdy2RtHS1), .Y(n178));
NAND3X1  g053(.A(n135), .B(State_1), .C(n178), .Y(n179));
NAND3X1  g054(.A(State_0), .B(n132), .C(n148), .Y(n180));
AOI21X1  g055(.A0(n180), .A1(n179), .B0(n142), .Y(n181_1));
OAI21X1  g056(.A0(n181_1), .A1(n141_1), .B0(State_4), .Y(n182));
OR4X1    g057(.A(State_0), .B(n162), .C(InDoneHS1), .D(n133_1), .Y(n183));
NAND4X1  g058(.A(n182), .B(n177_1), .C(n172), .D(n183), .Y(n84));
NAND4X1  g059(.A(State_0), .B(n128), .C(State_3), .D(n158), .Y(n185_1));
OR2X1    g060(.A(n185_1), .B(TpArrayHS1), .Y(n186));
OR2X1    g061(.A(FullIHS1), .B(FullOHS1), .Y(n187));
NOR4X1   g062(.A(State_0), .B(n148), .C(n147), .D(n187), .Y(n188));
NOR4X1   g063(.A(State_2), .B(State_4), .C(State_5), .D(State_1), .Y(n189_1));
OAI21X1  g064(.A0(n188), .A1(State_3), .B0(n189_1), .Y(n190));
NOR2X1   g065(.A(n135), .B(State_1), .Y(n191));
NAND2X1  g066(.A(n158), .B(State_3), .Y(n192));
INVX1    g067(.A(n192), .Y(n193_1));
NAND4X1  g068(.A(n135), .B(State_1), .C(State_2), .D(n158), .Y(n194));
INVX1    g069(.A(n194), .Y(n195));
AOI22X1  g070(.A0(n193_1), .A1(n191), .B0(State_3), .B1(n195), .Y(n196));
NAND3X1  g071(.A(n196), .B(n190), .C(n186), .Y(n89));
OR2X1    g072(.A(n185_1), .B(n132), .Y(n198));
OR4X1    g073(.A(State_2), .B(State_3), .C(State_4), .D(State_1), .Y(n199));
NOR2X1   g074(.A(n199), .B(State_5), .Y(n200));
AND2X1   g075(.A(n200), .B(n188), .Y(n201));
NOR4X1   g076(.A(n142), .B(n128), .C(InDoneHS1), .D(n143), .Y(n202));
AOI21X1  g077(.A0(n127), .A1(RtTSHS1), .B0(n159), .Y(n203));
NOR4X1   g078(.A(n202), .B(n201), .C(n195), .D(n203), .Y(n204));
NOR2X1   g079(.A(Rdy2RtHS1), .B(n126), .Y(n205));
NAND4X1  g080(.A(n128), .B(n127), .C(State_5), .D(n135), .Y(n206));
NOR3X1   g081(.A(n131), .B(FullIHS1), .C(FullOHS1), .Y(n207));
NOR2X1   g082(.A(n207), .B(State_4), .Y(n208));
NOR3X1   g083(.A(n208), .B(n206), .C(n132), .Y(n209));
NAND2X1  g084(.A(n209), .B(n205), .Y(n210));
NAND2X1  g085(.A(n148), .B(Rdy1BmHS1), .Y(n211));
OR4X1    g086(.A(n211), .B(n133_1), .C(n135), .D(n208), .Y(n212));
NAND4X1  g087(.A(n210), .B(n204), .C(n198), .D(n212), .Y(n94));
AND2X1   g088(.A(WantBmHS1), .B(Rdy2BmHS1), .Y(n214));
INVX1    g089(.A(n214), .Y(n215));
NOR4X1   g090(.A(n206), .B(n131), .C(n126), .D(n167), .Y(n216));
AOI22X1  g091(.A0(n168), .A1(Rdy2RtHS1), .B0(n132), .B1(n216), .Y(n217));
OR2X1    g092(.A(n217), .B(n215), .Y(n218));
INVX1    g093(.A(WantRtHS1), .Y(n219));
NAND3X1  g094(.A(n214), .B(n168), .C(n219), .Y(n220));
NAND2X1  g095(.A(Rdy2BmHS1), .B(n147), .Y(n221));
NOR4X1   g096(.A(n208), .B(n133_1), .C(n135), .D(n221), .Y(n222));
OR4X1    g097(.A(n129_1), .B(n135), .C(State_4), .D(n136), .Y(n223));
OAI21X1  g098(.A0(n223), .A1(n132), .B0(n185_1), .Y(n224));
NOR3X1   g099(.A(n194), .B(n127), .C(InDoneHS1), .Y(n225));
NAND4X1  g100(.A(State_1), .B(n127), .C(n162), .D(n135), .Y(n226));
NOR3X1   g101(.A(n226), .B(n152), .C(n128), .Y(n227));
NOR4X1   g102(.A(n225), .B(n224), .C(n222), .D(n227), .Y(n228));
MX2X1    g103(.A(InDoneHS1), .B(n136), .S0(Prog_2), .Y(n229));
OAI21X1  g104(.A0(n229), .A1(State_4), .B0(n128), .Y(n230));
NOR2X1   g105(.A(State_4), .B(Prog_2), .Y(n231));
NOR2X1   g106(.A(n152), .B(n231), .Y(n232));
OR2X1    g107(.A(n232), .B(n230), .Y(n233));
NOR2X1   g108(.A(Rdy2BmHS1), .B(n147), .Y(n234));
MX2X1    g109(.A(n234), .B(n205), .S0(Prog_0), .Y(n235));
NOR2X1   g110(.A(State_1), .B(State_4), .Y(n236));
NAND2X1  g111(.A(n236), .B(FullOHS1), .Y(n237));
NOR4X1   g112(.A(n206), .B(Prog_2), .C(FullIHS1), .D(n237), .Y(n238));
AOI22X1  g113(.A0(n235), .A1(n238), .B0(n233), .B1(n154), .Y(n239));
NAND4X1  g114(.A(n228), .B(n220), .C(n218), .D(n239), .Y(n99));
NAND3X1  g115(.A(WantBmHS1), .B(n148), .C(n147), .Y(n241));
NAND4X1  g116(.A(n168), .B(WantRtHS1), .C(Rdy2RtHS1), .D(n241), .Y(n242));
NAND3X1  g117(.A(n236), .B(n153_1), .C(n131), .Y(n243));
NOR2X1   g118(.A(n243), .B(FullOHS1), .Y(n244));
NAND2X1  g119(.A(n244), .B(n235), .Y(n245));
NOR4X1   g120(.A(State_1), .B(State_3), .C(n139), .D(n135), .Y(n246));
AOI21X1  g121(.A0(Rdy2BmHS1), .A1(Rdy1BmHS1), .B0(n231), .Y(n247));
OAI21X1  g122(.A0(n247), .A1(n230), .B0(n246), .Y(n248));
NOR2X1   g123(.A(n178), .B(Rdy1RtHS1), .Y(n249));
OAI21X1  g124(.A0(n223), .A1(n132), .B0(n190), .Y(n250));
AOI21X1  g125(.A0(n249), .A1(n209), .B0(n250), .Y(n251));
NAND4X1  g126(.A(n248), .B(n245), .C(n242), .D(n251), .Y(n104));
NOR4X1   g127(.A(State_2), .B(State_3), .C(n139), .D(State_1), .Y(n253));
NAND3X1  g128(.A(n253), .B(n135), .C(State_4), .Y(n254));
NOR4X1   g129(.A(n132), .B(State_3), .C(State_4), .D(State_0), .Y(n255));
NAND4X1  g130(.A(State_5), .B(Prog_0), .C(n131), .D(n255), .Y(n256));
NOR4X1   g131(.A(n142), .B(State_4), .C(Prog_2), .D(n149_1), .Y(n257));
NAND3X1  g132(.A(n257), .B(n128), .C(Prog_0), .Y(n258));
NAND3X1  g133(.A(n140), .B(n135), .C(State_1), .Y(n259));
NAND4X1  g134(.A(n258), .B(n256), .C(n254), .D(n259), .Y(ActRtHS1));
INVX1    g135(.A(Prog_0), .Y(n261));
NOR4X1   g136(.A(State_2), .B(n139), .C(Prog_2), .D(n226), .Y(n262));
OAI21X1  g137(.A0(n262), .A1(n257), .B0(n261), .Y(n263));
AOI21X1  g138(.A0(State_1), .A1(n128), .B0(State_0), .Y(n264));
AOI22X1  g139(.A0(n193_1), .A1(n264), .B0(n191), .B1(n140), .Y(n265));
NAND4X1  g140(.A(n263), .B(n185_1), .C(n254), .D(n265), .Y(ActBmHS1));
NAND4X1  g141(.A(n171), .B(WantRtHS1), .C(n178), .D(n216), .Y(n267));
XOR2X1   g142(.A(Rdy2RtHS1), .B(n126), .Y(n268));
AND2X1   g143(.A(FullIHS1), .B(FullOHS1), .Y(n269));
OR4X1    g144(.A(n268), .B(n243), .C(n261), .D(n269), .Y(n270));
OR2X1    g145(.A(FullOHS1), .B(Rdy1RtHS1), .Y(n271));
OR4X1    g146(.A(n135), .B(n132), .C(Rdy1BmHS1), .D(n271), .Y(n272));
NOR4X1   g147(.A(n129_1), .B(State_4), .C(FullIHS1), .D(n272), .Y(n273));
NOR4X1   g148(.A(State_3), .B(n178), .C(n126), .D(n194), .Y(n274));
NOR2X1   g149(.A(n274), .B(n273), .Y(n275));
NAND4X1  g150(.A(n270), .B(n267), .C(n210), .D(n275), .Y(GoRtHS1));
INVX1    g151(.A(FullOHS1), .Y(n277));
INVX1    g152(.A(FullIHS1), .Y(n278));
NAND4X1  g153(.A(n253), .B(n135), .C(n261), .D(n231), .Y(n279));
AOI21X1  g154(.A0(n221), .A1(n211), .B0(n279), .Y(n280));
OAI21X1  g155(.A0(n278), .A1(n277), .B0(n280), .Y(n281));
NOR3X1   g156(.A(n167), .B(n133_1), .C(n131), .Y(n282));
NAND4X1  g157(.A(n234), .B(n282), .C(WantBmHS1), .D(n173_1), .Y(n283));
NOR2X1   g158(.A(n273), .B(n201), .Y(n284));
NAND4X1  g159(.A(n283), .B(n281), .C(n212), .D(n284), .Y(GoBmHS1));
NAND3X1  g160(.A(n264), .B(n158), .C(State_3), .Y(n286));
NAND2X1  g161(.A(n286), .B(n185_1), .Y(NewTrHS1));
NOR2X1   g162(.A(n160), .B(n159), .Y(ReRtTSHS1));
NAND3X1  g163(.A(n255), .B(State_2), .C(State_5), .Y(n289));
NAND3X1  g164(.A(n255), .B(State_5), .C(n131), .Y(n290));
MX2X1    g165(.A(n254), .B(n290), .S0(n261), .Y(n291));
NAND3X1  g166(.A(n291), .B(n289), .C(n258), .Y(Mode0HS1));
AOI21X1  g167(.A0(n141_1), .A1(n162), .B0(n144), .Y(n293));
OAI21X1  g168(.A0(n254), .A1(n174), .B0(n293), .Y(Mode1HS1));
INVX1    g169(.A(n273), .Y(n295));
NOR3X1   g170(.A(n129_1), .B(State_4), .C(FullIHS1), .Y(n296));
NOR4X1   g171(.A(n132), .B(Rdy2RtHS1), .C(n126), .D(State_0), .Y(n297));
NOR4X1   g172(.A(State_1), .B(Rdy2BmHS1), .C(n147), .D(n135), .Y(n298));
OR2X1    g173(.A(n298), .B(n297), .Y(n299));
NAND4X1  g174(.A(n296), .B(Prog_2), .C(n277), .D(n299), .Y(n300));
AOI21X1  g175(.A0(ReRtTSHS1), .A1(Prog_2), .B0(n201), .Y(n301));
NAND4X1  g176(.A(n300), .B(n295), .C(n243), .D(n301), .Y(NewLineHS1));
INVX1    g177(.A(n185_1), .Y(n303));
AOI22X1  g178(.A0(n138), .A1(State_2), .B0(n131), .B1(n191), .Y(n304));
NOR3X1   g179(.A(n304), .B(n142), .C(State_4), .Y(n305));
NAND4X1  g180(.A(n132), .B(n128), .C(State_3), .D(n158), .Y(n306));
OAI21X1  g181(.A0(n194), .A1(n127), .B0(n306), .Y(n307));
OR4X1    g182(.A(n305), .B(n303), .C(Mode2HS1), .D(n307), .Y(ShftORHS1));
OR2X1    g183(.A(n262), .B(Mode2HS1), .Y(ShftIRHS1));
NOR2X1   g184(.A(n133_1), .B(n131), .Y(n310));
NOR3X1   g185(.A(n269), .B(n133_1), .C(Prog_0), .Y(n311));
OAI21X1  g186(.A0(n311), .A1(n310), .B0(n148), .Y(n312));
NOR2X1   g187(.A(n206), .B(n131), .Y(n313));
NOR3X1   g188(.A(n269), .B(n206), .C(n261), .Y(n314));
OAI21X1  g189(.A0(n314), .A1(n313), .B0(n178), .Y(n315));
NOR3X1   g190(.A(n199), .B(State_0), .C(n131), .Y(n316));
NOR4X1   g191(.A(State_1), .B(State_4), .C(State_5), .D(State_0), .Y(n317));
NOR3X1   g192(.A(n317), .B(n316), .C(n303), .Y(n318));
NAND3X1  g193(.A(n318), .B(n315), .C(n312), .Y(LxHInHS1));
MX2X1    g194(.A(Rdy2RtHS1), .B(n147), .S0(n261), .Y(n320));
NAND4X1  g195(.A(n153_1), .B(n131), .C(n278), .D(n320), .Y(n321));
NAND3X1  g196(.A(n261), .B(n277), .C(Rdy2BmHS1), .Y(n322));
NOR3X1   g197(.A(n322), .B(n206), .C(Prog_2), .Y(n323));
NOR3X1   g198(.A(n323), .B(n317), .C(n303), .Y(n324));
NOR4X1   g199(.A(n206), .B(n261), .C(Prog_2), .D(n271), .Y(n325));
AOI21X1  g200(.A0(n130), .A1(State_0), .B0(n325), .Y(n326));
NAND3X1  g201(.A(n326), .B(n324), .C(n321), .Y(TxHInHS1));
AOI22X1  g202(.A0(n168), .A1(n219), .B0(n178), .B1(n216), .Y(n328));
NOR2X1   g203(.A(n328), .B(WantBmHS1), .Y(n329));
NOR4X1   g204(.A(n243), .B(n261), .C(FullOHS1), .D(n268), .Y(n330));
NOR2X1   g205(.A(State_0), .B(State_1), .Y(n331));
NAND2X1  g206(.A(n331), .B(State_2), .Y(n332));
NAND4X1  g207(.A(State_1), .B(n128), .C(TpArrayHS1), .D(State_0), .Y(n333));
AOI21X1  g208(.A0(n333), .A1(n332), .B0(n192), .Y(n334));
NOR2X1   g209(.A(n334), .B(n273), .Y(n335));
NAND2X1  g210(.A(n335), .B(n300), .Y(n336));
OR4X1    g211(.A(n133_1), .B(State_4), .C(n131), .D(n187), .Y(n337));
NAND2X1  g212(.A(n173_1), .B(n234), .Y(n338));
XOR2X1   g213(.A(Rdy2BmHS1), .B(Rdy1BmHS1), .Y(n339));
NAND2X1  g214(.A(n339), .B(n277), .Y(n340));
OAI22X1  g215(.A0(n338), .A1(n337), .B0(n279), .B1(n340), .Y(n341));
OR4X1    g216(.A(n336), .B(n330), .C(n329), .D(n341), .Y(LoadOHHS1));
NAND4X1  g217(.A(n175), .B(n168), .C(n219), .D(n214), .Y(n343));
NAND4X1  g218(.A(n131), .B(FullOHS1), .C(n126), .D(Prog_0), .Y(n344));
OR2X1    g219(.A(Prog_0), .B(WantBmHS1), .Y(n345));
OR4X1    g220(.A(n131), .B(FullOHS1), .C(n219), .D(n345), .Y(n346));
NAND2X1  g221(.A(n346), .B(n344), .Y(n347));
NAND4X1  g222(.A(n296), .B(n331), .C(Rdy2RtHS1), .D(n347), .Y(n348));
MX2X1    g223(.A(n205), .B(n339), .S0(n261), .Y(n349));
NAND2X1  g224(.A(n349), .B(n238), .Y(n350));
NAND3X1  g225(.A(n350), .B(n348), .C(n343), .Y(LoadIHHS1));
NOR2X1   g226(.A(n136), .B(OutAvHS1), .Y(SeOutAvHS1));
NAND3X1  g227(.A(n249), .B(n244), .C(Prog_0), .Y(n353));
AND2X1   g228(.A(Mode2HS1), .B(OutputHS1), .Y(n354));
OAI21X1  g229(.A0(n354), .A1(n305), .B0(InDoneHS1), .Y(n355));
OR4X1    g230(.A(FullOHS1), .B(n148), .C(Rdy1BmHS1), .D(n279), .Y(n356));
NAND4X1  g231(.A(n355), .B(n353), .C(n335), .D(n356), .Y(SeFullOHS1));
OR4X1    g232(.A(n221), .B(FullIHS1), .C(n277), .D(n279), .Y(n358));
NAND2X1  g233(.A(n262), .B(InDoneHS1), .Y(n359));
NAND4X1  g234(.A(n358), .B(n348), .C(n343), .D(n359), .Y(SeFullIHS1));
NOR2X1   g235(.A(n278), .B(OutAvHS1), .Y(TgWhBufHS1));
NOR2X1   g236(.A(FullIHS1), .B(OutAvHS1), .Y(ReWhBufHS1));
NOR2X1   g237(.A(State_2), .B(n127), .Y(n363));
AND2X1   g238(.A(n363), .B(n317), .Y(LdProgHS1));
NAND3X1  g239(.A(n168), .B(WantRtHS1), .C(Rdy2RtHS1), .Y(n365));
OAI21X1  g240(.A0(n345), .A1(n365), .B0(n343), .Y(DumpIHS1));
endmodule
