// Benchmark "b20_C" written by ABC on Wed Aug 05 14:44:27 2020

module b20_C ( 
    P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
    SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_, SI_17_,
    SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_, SI_8_,
    SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
    P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
    P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
    P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
    P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
    P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
    P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
    P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
    P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
    P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
    P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN,
    P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN,
    P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN,
    P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN,
    P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN,
    P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
    P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
    P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
    P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
    P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
    P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
    P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
    P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
    P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
    P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
    P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
    P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
    P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN,
    P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
    P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
    P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
    P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
    P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
    P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
    P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
    P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
    P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
    P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
    P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
    P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
    P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
    P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
    P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
    P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
    P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
    P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
    P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
    P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
    P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
    P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
    P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
    P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
    P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
    P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
    P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
    P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
    P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
    P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
    P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
    P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
    P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
    P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
    P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
    P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
    P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
    P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
    P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
    P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
    P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
    P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
    P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
    P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
    P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
    P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
    P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
    P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
    P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
    P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
    P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
    P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
    P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
    P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
    P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
    P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
    P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
    P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
    P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
    P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
    P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
    P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
    P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
    P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
    P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
    P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
    P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
    P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
    P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
    P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
    P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
    P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
    P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
    P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
    P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
    P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
    P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
    P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
    P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
    P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
    P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
    P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
    P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
    P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
    P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
    P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
    P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
    P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
    P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
    P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
    P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
    P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
    P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
    P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
    P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
    P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
    P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
    P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
    P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
    P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
    P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
    P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
    P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
    P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
    P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
    P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
    P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
    P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
    P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
    P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
    P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
    P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
    P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
    P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
    P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
    P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
    P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
    P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
    P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
    P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
    P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
    P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
    P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
    P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
    P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
    P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
    P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
    P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
    P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
    P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
    P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
    P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
    P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
    P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
    P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
    P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
    P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
    P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
    P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
    P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
    P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
    P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
    P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
    P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
    P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
    P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
    P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
    P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
    P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
    P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
    P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
    P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
    P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
    P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
    P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
    P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
    P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
    P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
    P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
    P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
    P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
    P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
    P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
    P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
    P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
    P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
    P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
    P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
    P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
    P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
    P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
    P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
    P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
    P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
    P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
    P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
    P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
    P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
    P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
    P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
    P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
    ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
    ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
    ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
    ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
    U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
    P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
    P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
    P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
    P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440,
    P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
    P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
    P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
    P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
    P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465,
    P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486,
    P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507,
    P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
    P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
    P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
    P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
    P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
    P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
    P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
    P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
    P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
    P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
    P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
    P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
    P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
    P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554,
    P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
    P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
    P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
    P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
    P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
    P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
    P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
    P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
    P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
    P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290,
    P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283,
    P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276,
    P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269,
    P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377,
    P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257,
    P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250,
    P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243,
    P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236,
    P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402,
    P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423,
    P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444,
    P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452,
    P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459,
    P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466,
    P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473,
    P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480,
    P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487,
    P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230,
    P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223,
    P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216,
    P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209,
    P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202,
    P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195,
    P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188,
    P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491,
    P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498,
    P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505,
    P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
    P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
    P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179,
    P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
    P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
    P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
    P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150,
    P2_U3893  );
  input  P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_,
    SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
    SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
    SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
    P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, P2_REG3_REG_7__SCAN_IN,
    P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
    P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
    P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
    P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
    P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
    P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
    P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
    P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
    P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN,
    P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN,
    P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN,
    P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN,
    P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN,
    P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
    P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
    P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
    P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
    P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
    P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
    P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
    P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
    P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
    P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
    P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
    P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
    P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, P1_IR_REG_0__SCAN_IN,
    P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
    P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
    P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
    P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
    P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
    P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
    P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
    P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
    P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
    P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
    P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
    P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
    P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
    P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
    P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
    P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
    P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
    P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
    P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
    P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
    P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
    P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
    P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
    P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
    P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
    P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
    P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
    P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
    P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
    P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
    P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
    P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
    P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
    P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
    P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
    P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
    P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
    P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
    P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
    P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
    P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
    P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
    P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
    P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
    P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
    P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
    P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
    P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
    P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
    P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
    P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
    P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
    P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
    P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
    P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
    P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
    P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
    P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
    P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
    P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
    P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
    P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
    P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
    P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
    P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
    P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
    P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
    P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
    P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
    P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
    P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
    P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
    P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
    P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
    P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
    P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
    P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
    P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
    P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
    P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
    P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
    P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
    P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
    P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
    P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
    P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
    P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
    P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
    P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
    P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
    P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
    P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
    P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
    P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
    P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
    P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
    P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
    P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
    P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
    P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
    P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
    P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
    P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
    P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
    P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
    P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
    P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
    P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
    P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
    P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
    P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
    P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
    P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
    P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
    P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
    P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
    P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
    P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
    P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
    P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
    P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
    P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
    P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
    P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
    P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
    P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
    P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
    P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
    P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
    P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
    P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
    P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
    P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
    P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
    P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
    P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
    P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
    P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
    P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
    P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
    P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
    P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
    P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
    P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
    P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
    P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
    P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
    P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
    P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
    P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
    P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
    P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
    P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
    P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
    P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
    P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
    P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
    P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
    P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
    P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
    P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
    P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
    P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
    P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
    P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
    P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
    P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
    P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
    P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
    P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
    P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
    P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
    P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
    P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
    P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
    P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
    P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
    P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
    P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
    P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
    P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN;
  output ADD_1068_U4, ADD_1068_U55, ADD_1068_U56, ADD_1068_U57, ADD_1068_U58,
    ADD_1068_U59, ADD_1068_U60, ADD_1068_U61, ADD_1068_U62, ADD_1068_U63,
    ADD_1068_U47, ADD_1068_U48, ADD_1068_U49, ADD_1068_U50, ADD_1068_U51,
    ADD_1068_U52, ADD_1068_U53, ADD_1068_U54, ADD_1068_U5, ADD_1068_U46,
    U126, U123, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
    P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
    P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
    P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
    P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3439, P1_U3440,
    P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
    P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
    P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
    P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
    P1_U3295, P1_U3294, P1_U3453, P1_U3456, P1_U3459, P1_U3462, P1_U3465,
    P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486,
    P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507,
    P1_U3509, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
    P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
    P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
    P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
    P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
    P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
    P1_U3551, P1_U3552, P1_U3553, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
    P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
    P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
    P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
    P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
    P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
    P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
    P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3554,
    P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
    P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
    P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
    P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
    P1_U3583, P1_U3584, P1_U3585, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
    P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
    P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
    P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
    P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
    P1_U3973, P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290,
    P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283,
    P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276,
    P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269,
    P2_U3268, P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3376, P2_U3377,
    P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257,
    P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250,
    P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243,
    P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236,
    P2_U3235, P2_U3234, P2_U3390, P2_U3393, P2_U3396, P2_U3399, P2_U3402,
    P2_U3405, P2_U3408, P2_U3411, P2_U3414, P2_U3417, P2_U3420, P2_U3423,
    P2_U3426, P2_U3429, P2_U3432, P2_U3435, P2_U3438, P2_U3441, P2_U3444,
    P2_U3446, P2_U3447, P2_U3448, P2_U3449, P2_U3450, P2_U3451, P2_U3452,
    P2_U3453, P2_U3454, P2_U3455, P2_U3456, P2_U3457, P2_U3458, P2_U3459,
    P2_U3460, P2_U3461, P2_U3462, P2_U3463, P2_U3464, P2_U3465, P2_U3466,
    P2_U3467, P2_U3468, P2_U3469, P2_U3470, P2_U3471, P2_U3472, P2_U3473,
    P2_U3474, P2_U3475, P2_U3476, P2_U3477, P2_U3478, P2_U3479, P2_U3480,
    P2_U3481, P2_U3482, P2_U3483, P2_U3484, P2_U3485, P2_U3486, P2_U3487,
    P2_U3488, P2_U3489, P2_U3490, P2_U3233, P2_U3232, P2_U3231, P2_U3230,
    P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223,
    P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216,
    P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209,
    P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202,
    P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195,
    P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188,
    P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3491,
    P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498,
    P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505,
    P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
    P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
    P2_U3520, P2_U3521, P2_U3522, P2_U3296, P2_U3181, P2_U3180, P2_U3179,
    P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
    P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
    P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
    P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3151, P2_U3150,
    P2_U3893;
  wire n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
    n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
    n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
    n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
    n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
    n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1094,
    n1096, n1097, n1099, n1100, n1102, n1104, n1106, n1108, n1110, n1112,
    n1114, n1116, n1118, n1120, n1122, n1124, n1126, n1128, n1130, n1131,
    n1132, n1133, n1134, n1135, n1138, n1140, n1142, n1143, n1144, n1145,
    n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
    n1156, n1158, n1159, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
    n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
    n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1186, n1187, n1188,
    n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
    n1199, n1200, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
    n1210, n1211, n1212, n1213, n1214, n1215, n1217, n1218, n1219, n1220,
    n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
    n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
    n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
    n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1261, n1262,
    n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
    n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
    n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
    n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
    n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
    n1314, n1315, n1316, n1317, n1318, n1320, n1321, n1322, n1323, n1324,
    n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
    n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1345,
    n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
    n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1365, n1366,
    n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
    n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1387,
    n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
    n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
    n1408, n1409, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
    n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
    n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
    n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1448, n1449, n1450,
    n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
    n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1469, n1470, n1471,
    n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
    n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
    n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
    n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
    n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
    n1523, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
    n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1543, n1544,
    n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
    n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
    n1565, n1566, n1567, n1568, n1569, n1571, n1572, n1573, n1574, n1575,
    n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
    n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1594, n1595, n1596,
    n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
    n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
    n1617, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
    n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1637, n1638,
    n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
    n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
    n1659, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
    n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
    n1680, n1681, n1682, n1683, n1684, n1685, n1687, n1688, n1689, n1690,
    n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
    n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1709, n1710, n1711,
    n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
    n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1731, n1732,
    n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
    n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
    n1753, n1754, n1755, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
    n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
    n1774, n1775, n1776, n1777, n1778, n1780, n1781, n1782, n1783, n1784,
    n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
    n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
    n1805, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
    n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
    n1826, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
    n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
    n1847, n1848, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
    n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
    n1868, n1869, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
    n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
    n1889, n1890, n1891, n1892, n1893, n1895, n1896, n1898, n1900, n1902,
    n1904, n1906, n1908, n1910, n1912, n1914, n1916, n1918, n1920, n1922,
    n1924, n1926, n1928, n1930, n1932, n1934, n1936, n1938, n1940, n1942,
    n1944, n1946, n1948, n1950, n1952, n1954, n1956, n1958, n1959, n1960,
    n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
    n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
    n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
    n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
    n2001, n2002, n2003, n2004, n2005, n2006, n2008, n2009, n2010, n2011,
    n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
    n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
    n2032, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
    n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
    n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
    n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2071, n2072, n2073,
    n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
    n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
    n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
    n2104, n2105, n2106, n2107, n2108, n2110, n2111, n2112, n2113, n2114,
    n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2123, n2124, n2125,
    n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
    n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
    n2146, n2147, n2148, n2149, n2150, n2151, n2153, n2154, n2155, n2156,
    n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
    n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
    n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
    n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
    n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
    n2208, n2209, n2211, n2212, n2213, n2215, n2218, n2219, n2220, n2221,
    n2222, n2223, n2224, n2225, n2226, n2227, n2229, n2230, n2231, n2232,
    n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
    n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
    n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
    n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
    n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2283, n2284,
    n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
    n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
    n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
    n2315, n2316, n2317, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
    n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
    n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2345, n2346,
    n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
    n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
    n2367, n2368, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
    n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
    n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
    n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
    n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2416, n2417, n2418,
    n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2427, n2428, n2429,
    n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
    n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
    n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
    n2460, n2461, n2462, n2463, n2465, n2466, n2467, n2468, n2469, n2470,
    n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
    n2481, n2482, n2483, n2484, n2485, n2486, n2488, n2489, n2490, n2491,
    n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
    n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2511, n2512,
    n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
    n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
    n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
    n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
    n2554, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
    n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
    n2575, n2576, n2577, n2578, n2579, n2580, n2582, n2583, n2584, n2585,
    n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
    n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
    n2606, n2607, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
    n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
    n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2637,
    n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
    n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2657, n2658,
    n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
    n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
    n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
    n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
    n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2709,
    n2710, n2711, n2712, n2713, n2714, n2715, n2717, n2718, n2719, n2720,
    n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
    n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
    n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
    n2751, n2752, n2753, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
    n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
    n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
    n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
    n2792, n2793, n2794, n2795, n2796, n2798, n2799, n2801, n2802, n2803,
    n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
    n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2823, n2824, n2825,
    n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
    n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
    n2846, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
    n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
    n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
    n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
    n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
    n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
    n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
    n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
    n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2940,
    n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
    n2951, n2952, n2953, n2954, n2956, n2957, n2958, n2959, n2960, n2961,
    n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
    n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
    n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
    n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
    n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
    n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
    n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
    n3033, n3034, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
    n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
    n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
    n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
    n3074, n3075, n3076, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
    n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
    n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
    n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
    n3115, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
    n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
    n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
    n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
    n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
    n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
    n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
    n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
    n3197, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
    n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3218,
    n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
    n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
    n3239, n3240, n3241, n3243, n3244, n3245, n3246, n3247, n3249, n3250,
    n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
    n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
    n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
    n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3289, n3290, n3291,
    n3292, n3293, n3294, n3295, n3297, n3298, n3299, n3300, n3301, n3302,
    n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
    n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
    n3323, n3324, n3325, n3326, n3327, n3329, n3330, n3331, n3332, n3333,
    n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
    n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
    n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
    n3364, n3365, n3366, n3367, n3368, n3369, n3371, n3372, n3373, n3374,
    n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
    n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
    n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
    n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
    n3415, n3416, n3417, n3418, n3420, n3421, n3422, n3423, n3424, n3425,
    n3426, n3427, n3428, n3429, n3430, n3432, n3433, n3434, n3435, n3436,
    n3437, n3439, n3440, n3441, n3443, n3445, n3447, n3449, n3451, n3453,
    n3455, n3457, n3459, n3461, n3463, n3465, n3467, n3469, n3471, n3473,
    n3475, n3477, n3479, n3481, n3483, n3485, n3487, n3489, n3491, n3493,
    n3495, n3497, n3499, n3501, n3503, n3505, n3506, n3507, n3508, n3509,
    n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
    n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3528, n3529, n3530,
    n3531, n3532, n3534, n3535, n3536, n3537, n3538, n3539, n3541, n3542,
    n3543, n3544, n3545, n3546, n3547, n3549, n3550, n3551, n3552, n3553,
    n3554, n3555, n3556, n3557, n3558, n3560, n3561, n3562, n3563, n3564,
    n3565, n3567, n3568, n3569, n3570, n3572, n3573, n3574, n3575, n3576,
    n3577, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3587, n3588,
    n3589, n3590, n3591, n3592, n3593, n3595, n3596, n3597, n3598, n3599,
    n3600, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3610, n3611,
    n3612, n3613, n3614, n3615, n3616, n3617, n3619, n3620, n3621, n3622,
    n3623, n3624, n3626, n3627, n3628, n3629, n3630, n3631, n3633, n3634,
    n3635, n3636, n3637, n3638, n3640, n3641, n3642, n3643, n3644, n3646,
    n3647, n3648, n3649, n3650, n3651, n3653, n3654, n3655, n3656, n3657,
    n3658, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3668, n3669,
    n3670, n3671, n3672, n3673, n3675, n3676, n3677, n3678, n3679, n3680,
    n3681, n3682, n3683, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
    n3692, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3702, n3703,
    n3704, n3705, n3706, n3707, n3708, n3709, n3711, n3712, n3713, n3714,
    n3715, n3716, n3717, n3718, n3720, n3721, n3722, n3723, n3724, n3725,
    n3726, n3727, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
    n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3746, n3747, n3748,
    n3749, n3750, n3751, n3752, n3753, n3755, n3756, n3757, n3758, n3759,
    n3760, n3761, n3762, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
    n3771, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
    n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
    n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
    n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
    n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
    n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
    n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
    n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
    n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3862, n3863,
    n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
    n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
    n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
    n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
    n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
    n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
    n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
    n3934, n3935, n3936, n3937, n3938, n3939, n3941, n3943, n3944, n3945,
    n3946, n3947, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
    n3957, n3958, n3960, n3961, n3962, n3963, n3966, n3967, n3968, n3969,
    n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3978, n3979, n3980,
    n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
    n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4001,
    n4002, n4003, n4004, n4005, n4007, n4008, n4009, n4010, n4011, n4012,
    n4013, n4014, n4015, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
    n4024, n4025, n4026, n4027, n4028, n4030, n4031, n4032, n4033, n4034,
    n4035, n4036, n4037, n4038, n4039, n4040, n4042, n4043, n4044, n4045,
    n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
    n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
    n4066, n4067, n4068, n4069, n4073, n4074, n4075, n4076, n4077, n4079,
    n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4088, n4089, n4090,
    n4091, n4092, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
    n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
    n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
    n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4132, n4134,
    n4135, n4136, n4137, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
    n4146, n4148, n4149, n4150, n4152, n4153, n4154, n4156, n4157, n4158,
    n4159, n4160, n4161, n4162, n4164, n4165, n4166, n4167, n4168, n4169,
    n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
    n4180, n4181, n4182, n4183, n4184, n4186, n4187, n4189, n4190, n4191,
    n4192, n4193, n4195, n4196, n4197, n4198, n4199, n4201, n4202, n4203,
    n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
    n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
    n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
    n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
    n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
    n4256, n4257, n4258, n4260, n4261, n4262, n4263, n4264, n4265, n4267,
    n4268, n4269, n4270, n4271, n4272, n4274, n4275, n4276, n4277, n4278,
    n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4289,
    n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
    n4300, n4301, n4302, n4303, n4304, n4305, n4307, n4308, n4309, n4310,
    n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4319, n4320, n4321,
    n4322, n4323, n4324, n4325, n4326, n4328, n4330, n4332, n4334, n4336,
    n4338, n4340, n4342, n4344, n4346, n4348, n4350, n4352, n4354, n4356,
    n4358, n4360, n4362, n4364, n4366, n4368, n4370, n4372, n4374, n4376,
    n4378, n4380, n4382, n4384, n4386, n4388, n4390, n4391, n4392, n4394,
    n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
    n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
    n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
    n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
    n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
    n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
    n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
    n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
    n4475, n4476, n4477, n4478, n4482, n4483, n4484, n4485, n4486, n4487,
    n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
    n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
    n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
    n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
    n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
    n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
    n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
    n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
    n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
    n4578, n4580, n4581, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
    n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
    n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
    n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
    n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
    n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
    n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
    n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
    n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
    n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
    n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
    n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
    n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
    n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
    n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
    n4730, n4731, n4732, n4733, n4735, n4736, n4740, n4742, n4744, n4748,
    n4749, n4750, n4752, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
    n4763, n4766, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4776,
    n4778, n4779, n4780, n4781, n4782, n4784, n4785, n4786, n4787, n4788,
    n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
    n4800, n4803, n4804, n4805, n4806, n4808, n4809, n4810, n4811, n4812,
    n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4824,
    n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4834, n4835, n4839,
    n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
    n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
    n4860, n4861, n4862, n4863, n4864, n4865, n4867, n4868, n4869, n4870,
    n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
    n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
    n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
    n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
    n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
    n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
    n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
    n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
    n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
    n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
    n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
    n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
    n4991, n4992, n4993, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
    n5002, n5004, n5005, n5006, n5008, n5009, n5010, n5011, n5012, n5013,
    n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
    n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
    n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
    n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
    n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
    n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
    n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
    n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
    n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
    n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
    n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
    n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
    n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
    n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
    n5154, n5155, n5156, n5157, n5158, n5160, n5161, n5162, n5163, n5164,
    n5165, n5166, n5167, n5168, n5169, n5170, n5172, n5173, n5174, n5175,
    n5176, n5177, n5178, n5180, n5181, n5182, n5183, n5184, n5185, n5186,
    n5187, n5188, n5189, n5190, n5191, n5193, n5194, n5195, n5196, n5197,
    n5198, n5199, n5200, n5201, n5202, n5204, n5205, n5207, n5208, n5209,
    n5210, n5211, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
    n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5229, n5230, n5231,
    n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5241, n5242, n5243,
    n5244, n5245, n5246, n5247, n5249, n5250, n5251, n5252, n5253, n5254,
    n5255, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5266,
    n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5276, n5277,
    n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
    n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5297, n5298, n5299,
    n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5309, n5310,
    n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5321,
    n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
    n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
    n5343, n5344, n5345, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
    n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5363, n5364, n5365,
    n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
    n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
    n5386, n5387, n5388, n5390, n5391, n5392, n5393, n5394, n5395, n5396,
    n5397, n5398, n5399, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
    n5408, n5409, n5410, n5411, n5413, n5414, n5415, n5416, n5417, n5418,
    n5419, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
    n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5439, n5440, n5441,
    n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
    n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
    n5463, n5465, n5466, n5467, n5469, n5470, n5472, n5473, n5474, n5475,
    n5476, n5478, n5479, n5480, n5481, n5482, n5483, n5485, n5486, n5487,
    n5488, n5489, n5490, n5492, n5493, n5494, n5495, n5496, n5497, n5499,
    n5500, n5501, n5502, n5503, n5505, n5506, n5507, n5508, n5509, n5510,
    n5511, n5512, n5513, n5515, n5516, n5517, n5518, n5519, n5521, n5522,
    n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5532, n5533,
    n5534, n5535, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5545,
    n5546, n5547, n5548, n5549, n5551, n5552, n5553, n5554, n5555, n5556,
    n5557, n5558, n5559, n5560, n5562, n5563, n5564, n5565, n5567, n5568,
    n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5577, n5578, n5579,
    n5580, n5581, n5582, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
    n5591, n5592, n5593, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
    n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
    n5614, n5615, n5616, n5617, n5618, n5619, n5621, n5622, n5623, n5624,
    n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5633, n5634, n5635,
    n5636, n5637, n5638, n5640, n5641, n5642, n5643, n5644, n5645, n5646,
    n5647, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5657, n5658,
    n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5667, n5668, n5669,
    n5670, n5671, n5672, n5673, n5675, n5676, n5677, n5678, n5679, n5680,
    n5681, n5682, n5683, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
    n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
    n5704, n5705, n5706, n5707, n5708, n5709, n5711, n5712, n5713, n5714,
    n5715, n5716, n5717, n5719, n5720, n5721, n5722, n5723, n5724, n5726,
    n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736,
    n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746,
    n5747, n5748, n5750, n5751, n5752, n5754, n5756, n5758, n5760, n5762,
    n5764, n5766, n5768, n5770, n5772, n5774, n5776, n5778, n5780, n5782,
    n5784, n5786, n5788, n5790, n5792, n5794, n5796, n5798, n5800, n5802,
    n5804, n5806, n5808, n5810, n5812, n5814, n5815, n5816, n5817, n5818,
    n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
    n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
    n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
    n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
    n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
    n5869, n5870, n5871, n5872, n5873, n5874, n5876, n5877, n5878, n5879,
    n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
    n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
    n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
    n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
    n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
    n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
    n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
    n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
    n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
    n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
    n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
    n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
    n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
    n6013, n6014, n6015, n6016, n6018, n6019, n6020, n6021, n6022, n6023,
    n6024, n6025, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
    n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
    n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
    n6055, n6056, n6057, n6058, n6059, n6060, n6062, n6063, n6064, n6065,
    n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
    n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
    n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
    n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6104, n6105, n6106,
    n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116,
    n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126,
    n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136,
    n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146,
    n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6156, n6157,
    n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167,
    n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177,
    n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187,
    n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197,
    n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6206, n6207, n6208,
    n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
    n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
    n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
    n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6248, n6249,
    n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6259, n6260,
    n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
    n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
    n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6290, n6291,
    n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
    n6302, n6303, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
    n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
    n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
    n6333, n6334, n6335, n6336, n6337, n6338, n6340, n6341, n6342, n6343,
    n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
    n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
    n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
    n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
    n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
    n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
    n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
    n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
    n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6435, n6436,
    n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446,
    n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456,
    n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466,
    n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6476, n6477,
    n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487,
    n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497,
    n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
    n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
    n6518, n6519, n6520, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
    n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
    n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
    n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
    n6559, n6560, n6561, n6562, n6563, n6565, n6566, n6567, n6568, n6569,
    n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
    n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
    n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6599, n6600,
    n6601, n6602, n6603, n6604, n6605, n6607, n6608, n6609, n6610, n6611,
    n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
    n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
    n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
    n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6651, n6652,
    n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
    n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
    n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
    n6683, n6684, n6685, n6686, n6687, n6688, n6690, n6691, n6692, n6693,
    n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
    n6705, n6706, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
    n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
    n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6735, n6736,
    n6737, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
    n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
    n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
    n6769, n6770, n6771, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
    n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
    n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
    n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
    n6810, n6812, n6813, n6814, n6815, n6816, n6818, n6819, n6820, n6821,
    n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
    n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
    n6842, n6843, n6844, n6845, n6846, n6848, n6849, n6850, n6851, n6852,
    n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
    n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
    n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
    n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
    n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
    n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
    n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6922, n6923, n6924,
    n6925, n6926, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
    n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
    n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
    n6956, n6957, n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966,
    n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976,
    n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986,
    n6987, n6988, n6989, n6990, n6991, n6993, n6994, n6995, n6996, n6997,
    n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007,
    n7008, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
    n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7029, n7030,
    n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7039, n7040, n7041,
    n7042, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
    n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
    n7063, n7064, n7065, n7066, n7067, n7068, n7070, n7071, n7072, n7073,
    n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
    n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
    n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
    n7104, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
    n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
    n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
    n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7144, n7145,
    n7146, n7147, n7148, n7149, n7150, n7151, n7153, n7154, n7155, n7157,
    n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
    n7169, n7170, n7172, n7173, n7175, n7177, n7179, n7181, n7183, n7185,
    n7187, n7189, n7191, n7193, n7195, n7197, n7199, n7201, n7203, n7205,
    n7207, n7209, n7211, n7213, n7215, n7217, n7219, n7221, n7223, n7225,
    n7227, n7229, n7231, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
    n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
    n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7258, n7259, n7260,
    n7261, n7262, n7263, n7264, n7266, n7267, n7268, n7269, n7270, n7271,
    n7272, n7273, n7275, n7276, n7277, n7278, n7279, n7280, n7282, n7283,
    n7284, n7285, n7286, n7287, n7289, n7290, n7291, n7292, n7293, n7295,
    n7296, n7297, n7298, n7299, n7300, n7301, n7303, n7304, n7305, n7306,
    n7308, n7309, n7310, n7311, n7312, n7313, n7315, n7316, n7317, n7318,
    n7319, n7321, n7322, n7323, n7324, n7325, n7326, n7328, n7329, n7330,
    n7331, n7333, n7334, n7335, n7336, n7337, n7339, n7340, n7341, n7342,
    n7343, n7344, n7346, n7347, n7348, n7349, n7351, n7352, n7353, n7354,
    n7355, n7357, n7358, n7359, n7360, n7361, n7363, n7364, n7365, n7366,
    n7367, n7368, n7369, n7371, n7372, n7373, n7374, n7376, n7377, n7378,
    n7379, n7380, n7382, n7383, n7384, n7385, n7386, n7388, n7389, n7390,
    n7391, n7392, n7394, n7395, n7396, n7397, n7398, n7400, n7401, n7402,
    n7403, n7404, n7405, n7406, n7408, n7409, n7410, n7411, n7412, n7413,
    n7415, n7416, n7417, n7418, n7419, n7420, n7422, n7423, n7424, n7425,
    n7426, n7427, n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7437,
    n7438, n7439, n7440, n7441, n7443, n7444, n7445, n7446, n7448, n7449,
    n7450, n7451, n7453, n7454, n7456, n7457, n7458, n7459, n7460, n7461,
    n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471,
    n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481,
    n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491,
    n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501,
    n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511,
    n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521,
    n7524, n7525, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
    n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
    n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
    n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
    n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
    n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
    n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7596, n7599,
    n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
    n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
    n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
    n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
    n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
    n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
    n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
    n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
    n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
    n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
    n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
    n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
    n7720, n7721, n7722, n7723, n7724, n7725, n7727, n7728, n7729, n7730,
    n7731, n7732, n7733, n7734, n7736, n7737, n7738, n7739, n7740, n7741,
    n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751,
    n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
    n7763, n7764, n7765, n7766, n7767, n7768, n7770, n7771, n7772, n7773,
    n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
    n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
    n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
    n7805, n7806, n7807, n7808, n7810, n7811, n7812, n7813, n7814, n7815,
    n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7825, n7826,
    n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836,
    n7837, n7838, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847,
    n7848, n7849, n7850, n7851, n7852, n7853, n7855, n7856, n7857, n7858,
    n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
    n7869, n7870, n7871, n7872, n7873, n7874, n7876, n7877, n7878, n7879,
    n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
    n7890, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
    n7901, n7902, n7903, n7904, n7905, n7906, n7908, n7909, n7910, n7911,
    n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921,
    n7922, n7923, n7924, n7925, n7926, n7928, n7929, n7930, n7931, n7932,
    n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
    n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
    n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
    n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
    n7975, n7976, n7977, n7978, n7979, n7981, n7982, n7983, n7984, n7985,
    n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
    n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
    n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016,
    n8017, n8018, n8019, n8020, n8022, n8023, n8024, n8025, n8026, n8027,
    n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8037, n8038,
    n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
    n8049, n8050, n8051, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
    n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8068, n8070, n8072,
    n8074, n8076, n8078, n8080, n8082, n8084, n8086, n8088, n8090, n8092,
    n8094, n8096, n8098, n8100, n8102, n8104, n8106, n8108, n8110, n8112,
    n8114, n8116, n8118, n8120, n8122, n8124, n8126, n8128, n8129, n8131,
    n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
    n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
    n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
    n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
    n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
    n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
    n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
    n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
    n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
    n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
    n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
    n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
    n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
    n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
    n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
    n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
    n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303,
    n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
    n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323,
    n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333,
    n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343,
    n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353,
    n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363,
    n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373,
    n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383,
    n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393,
    n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
    n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
    n8414, n8415, n8416, n8417, n8421, n8422, n8423, n8424, n8425, n8426,
    n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436,
    n8439, n8441, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451,
    n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8462,
    n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
    n8474, n8475, n8476, n8477, n8478, n8480, n8481, n8482, n8483, n8487,
    n8488, n8489, n8490, n8492, n8494, n8495, n8496, n8497, n8498, n8499,
    n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511,
    n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8524,
    n8528, n8529, n8530, n8531, n8532, n8533, n8536, n8537, n8538, n8540,
    n8541, n8542, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
    n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8562, n8563,
    n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
    n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583,
    n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
    n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603,
    n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
    n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
    n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
    n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
    n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
    n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
    n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8674,
    n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
    n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
    n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
    n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
    n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
    n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
    n8735, n8736, n8737, n8738, n8739, n8740, n8745, n8746, n8747, n8748,
    n8749, n8751, n8752, n8753, n8755, n8756, n8757, n8758, n8759, n8760,
    n8761, n8762, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771,
    n8772, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
    n8783, n8784, n8785, n8787, n8788, n8789, n8790, n8792, n8793, n8794,
    n8795, n8796, n8797, n8798, n8800, n8801, n8802, n8803, n8804, n8805,
    n8806, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816,
    n8817, n8818, n8819, n8820, n8821, n8822, n8824, n8825, n8827, n8828,
    n8829, n8830, n8831, n8832, n8833, n8835, n8837, n8838, n8839, n8840,
    n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8851, n8852,
    n8853, n8854, n8855, n8856, n8857, n8859, n8860, n8861, n8862, n8863,
    n8864, n8865, n8866, n8867, n8869, n8870, n8871, n8872, n8873, n8874,
    n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8883, n8884, n8885,
    n8886, n8887, n8888, n8889, n8890, n8892, n8894, n8895, n8896, n8897,
    n8898, n8899, n8900, n8902, n8903, n8904, n8906, n8907, n8908, n8909,
    n8910, n8911, n8912, n8914, n8916, n8917, n8918, n8919, n8920, n8921,
    n8922, n8923, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
    n8933, n8934, n8935, n8936, n8938, n8939, n8940, n8941, n8942, n8943,
    n8944, n8945, n8946, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
    n8955, n8956, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
    n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
    n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8986,
    n8987, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8997, n8998,
    n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
    n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9019, n9020,
    n9021, n9022, n9023, n9024, n9025, n9027, n9028, n9029, n9030, n9031,
    n9032, n9033, n9034, n9035, n9036, n9038, n9039, n9040, n9041, n9042,
    n9043, n9044, n9045, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
    n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9062, n9063;
  NAND2X1 g0000(.A(P2_ADDR_REG_17__SCAN_IN), .B(P1_ADDR_REG_17__SCAN_IN), .Y(n1034));
  NOR2X1  g0001(.A(P2_ADDR_REG_17__SCAN_IN), .B(P1_ADDR_REG_17__SCAN_IN), .Y(n1035));
  NOR2X1  g0002(.A(P2_ADDR_REG_16__SCAN_IN), .B(P1_ADDR_REG_16__SCAN_IN), .Y(n1036));
  NAND2X1 g0003(.A(P2_ADDR_REG_15__SCAN_IN), .B(P1_ADDR_REG_15__SCAN_IN), .Y(n1037));
  NAND2X1 g0004(.A(P2_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), .Y(n1038));
  NAND2X1 g0005(.A(P2_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), .Y(n1039));
  NAND2X1 g0006(.A(P2_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), .Y(n1040));
  NAND2X1 g0007(.A(P2_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), .Y(n1041));
  NAND2X1 g0008(.A(P2_ADDR_REG_10__SCAN_IN), .B(P1_ADDR_REG_10__SCAN_IN), .Y(n1042));
  NAND2X1 g0009(.A(P2_ADDR_REG_9__SCAN_IN), .B(P1_ADDR_REG_9__SCAN_IN), .Y(n1043));
  NAND2X1 g0010(.A(P2_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), .Y(n1044));
  NAND2X1 g0011(.A(P2_ADDR_REG_7__SCAN_IN), .B(P1_ADDR_REG_7__SCAN_IN), .Y(n1045));
  NAND2X1 g0012(.A(P2_ADDR_REG_6__SCAN_IN), .B(P1_ADDR_REG_6__SCAN_IN), .Y(n1046));
  NAND2X1 g0013(.A(P2_ADDR_REG_5__SCAN_IN), .B(P1_ADDR_REG_5__SCAN_IN), .Y(n1047));
  NAND2X1 g0014(.A(P2_ADDR_REG_4__SCAN_IN), .B(P1_ADDR_REG_4__SCAN_IN), .Y(n1048));
  NAND2X1 g0015(.A(P2_ADDR_REG_3__SCAN_IN), .B(P1_ADDR_REG_3__SCAN_IN), .Y(n1049));
  NAND2X1 g0016(.A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Y(n1050));
  INVX1   g0017(.A(P2_ADDR_REG_1__SCAN_IN), .Y(n1051));
  NAND3X1 g0018(.A(P2_ADDR_REG_0__SCAN_IN), .B(P1_ADDR_REG_0__SCAN_IN), .C(P1_ADDR_REG_1__SCAN_IN), .Y(n1052));
  AOI21X1 g0019(.A0(P2_ADDR_REG_0__SCAN_IN), .A1(P1_ADDR_REG_0__SCAN_IN), .B0(P1_ADDR_REG_1__SCAN_IN), .Y(n1053));
  OAI21X1 g0020(.A0(n1053), .A1(n1051), .B0(n1052), .Y(n1054));
  OAI21X1 g0021(.A0(P2_ADDR_REG_2__SCAN_IN), .A1(P1_ADDR_REG_2__SCAN_IN), .B0(n1054), .Y(n1055));
  NAND2X1 g0022(.A(n1055), .B(n1050), .Y(n1056));
  OAI21X1 g0023(.A0(P2_ADDR_REG_3__SCAN_IN), .A1(P1_ADDR_REG_3__SCAN_IN), .B0(n1056), .Y(n1057));
  NAND2X1 g0024(.A(n1057), .B(n1049), .Y(n1058));
  OAI21X1 g0025(.A0(P2_ADDR_REG_4__SCAN_IN), .A1(P1_ADDR_REG_4__SCAN_IN), .B0(n1058), .Y(n1059));
  NAND2X1 g0026(.A(n1059), .B(n1048), .Y(n1060));
  OAI21X1 g0027(.A0(P2_ADDR_REG_5__SCAN_IN), .A1(P1_ADDR_REG_5__SCAN_IN), .B0(n1060), .Y(n1061));
  NAND2X1 g0028(.A(n1061), .B(n1047), .Y(n1062));
  OAI21X1 g0029(.A0(P2_ADDR_REG_6__SCAN_IN), .A1(P1_ADDR_REG_6__SCAN_IN), .B0(n1062), .Y(n1063));
  NAND2X1 g0030(.A(n1063), .B(n1046), .Y(n1064));
  OAI21X1 g0031(.A0(P2_ADDR_REG_7__SCAN_IN), .A1(P1_ADDR_REG_7__SCAN_IN), .B0(n1064), .Y(n1065));
  NAND2X1 g0032(.A(n1065), .B(n1045), .Y(n1066));
  OAI21X1 g0033(.A0(P2_ADDR_REG_8__SCAN_IN), .A1(P1_ADDR_REG_8__SCAN_IN), .B0(n1066), .Y(n1067));
  NAND2X1 g0034(.A(n1067), .B(n1044), .Y(n1068));
  OAI21X1 g0035(.A0(P2_ADDR_REG_9__SCAN_IN), .A1(P1_ADDR_REG_9__SCAN_IN), .B0(n1068), .Y(n1069));
  NAND2X1 g0036(.A(n1069), .B(n1043), .Y(n1070));
  OAI21X1 g0037(.A0(P2_ADDR_REG_10__SCAN_IN), .A1(P1_ADDR_REG_10__SCAN_IN), .B0(n1070), .Y(n1071));
  NAND2X1 g0038(.A(n1071), .B(n1042), .Y(n1072));
  OAI21X1 g0039(.A0(P2_ADDR_REG_11__SCAN_IN), .A1(P1_ADDR_REG_11__SCAN_IN), .B0(n1072), .Y(n1073));
  NAND2X1 g0040(.A(n1073), .B(n1041), .Y(n1074));
  OAI21X1 g0041(.A0(P2_ADDR_REG_12__SCAN_IN), .A1(P1_ADDR_REG_12__SCAN_IN), .B0(n1074), .Y(n1075));
  NAND2X1 g0042(.A(n1075), .B(n1040), .Y(n1076));
  OAI21X1 g0043(.A0(P2_ADDR_REG_13__SCAN_IN), .A1(P1_ADDR_REG_13__SCAN_IN), .B0(n1076), .Y(n1077));
  NAND2X1 g0044(.A(n1077), .B(n1039), .Y(n1078));
  OAI21X1 g0045(.A0(P2_ADDR_REG_14__SCAN_IN), .A1(P1_ADDR_REG_14__SCAN_IN), .B0(n1078), .Y(n1079));
  NAND2X1 g0046(.A(n1079), .B(n1038), .Y(n1080));
  OAI21X1 g0047(.A0(P2_ADDR_REG_15__SCAN_IN), .A1(P1_ADDR_REG_15__SCAN_IN), .B0(n1080), .Y(n1081));
  AOI21X1 g0048(.A0(n1081), .A1(n1037), .B0(n1036), .Y(n1082));
  AOI21X1 g0049(.A0(P2_ADDR_REG_16__SCAN_IN), .A1(P1_ADDR_REG_16__SCAN_IN), .B0(n1082), .Y(n1083));
  OAI21X1 g0050(.A0(n1083), .A1(n1035), .B0(n1034), .Y(n1084));
  AOI21X1 g0051(.A0(P2_ADDR_REG_18__SCAN_IN), .A1(P1_ADDR_REG_18__SCAN_IN), .B0(n1084), .Y(n1085));
  INVX1   g0052(.A(P1_ADDR_REG_19__SCAN_IN), .Y(n1086));
  XOR2X1  g0053(.A(P2_ADDR_REG_19__SCAN_IN), .B(n1086), .Y(n1087));
  INVX1   g0054(.A(n1087), .Y(n1088));
  OAI21X1 g0055(.A0(P2_ADDR_REG_18__SCAN_IN), .A1(P1_ADDR_REG_18__SCAN_IN), .B0(n1088), .Y(n1089));
  NOR2X1  g0056(.A(n1089), .B(n1085), .Y(n1090));
  OAI21X1 g0057(.A0(P2_ADDR_REG_18__SCAN_IN), .A1(P1_ADDR_REG_18__SCAN_IN), .B0(n1084), .Y(n1091));
  AOI21X1 g0058(.A0(P2_ADDR_REG_18__SCAN_IN), .A1(P1_ADDR_REG_18__SCAN_IN), .B0(n1088), .Y(n1092));
  AOI21X1 g0059(.A0(n1092), .A1(n1091), .B0(n1090), .Y(ADD_1068_U4));
  XOR2X1  g0060(.A(P2_ADDR_REG_18__SCAN_IN), .B(P1_ADDR_REG_18__SCAN_IN), .Y(n1094));
  XOR2X1  g0061(.A(n1094), .B(n1084), .Y(ADD_1068_U55));
  INVX1   g0062(.A(P1_ADDR_REG_17__SCAN_IN), .Y(n1096));
  XOR2X1  g0063(.A(P2_ADDR_REG_17__SCAN_IN), .B(n1096), .Y(n1097));
  XOR2X1  g0064(.A(n1097), .B(n1083), .Y(ADD_1068_U56));
  NAND2X1 g0065(.A(n1081), .B(n1037), .Y(n1099));
  XOR2X1  g0066(.A(P2_ADDR_REG_16__SCAN_IN), .B(P1_ADDR_REG_16__SCAN_IN), .Y(n1100));
  XOR2X1  g0067(.A(n1100), .B(n1099), .Y(ADD_1068_U57));
  XOR2X1  g0068(.A(P2_ADDR_REG_15__SCAN_IN), .B(P1_ADDR_REG_15__SCAN_IN), .Y(n1102));
  XOR2X1  g0069(.A(n1102), .B(n1080), .Y(ADD_1068_U58));
  XOR2X1  g0070(.A(P2_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), .Y(n1104));
  XOR2X1  g0071(.A(n1104), .B(n1078), .Y(ADD_1068_U59));
  XOR2X1  g0072(.A(P2_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), .Y(n1106));
  XOR2X1  g0073(.A(n1106), .B(n1076), .Y(ADD_1068_U60));
  XOR2X1  g0074(.A(P2_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), .Y(n1108));
  XOR2X1  g0075(.A(n1108), .B(n1074), .Y(ADD_1068_U61));
  XOR2X1  g0076(.A(P2_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), .Y(n1110));
  XOR2X1  g0077(.A(n1110), .B(n1072), .Y(ADD_1068_U62));
  XOR2X1  g0078(.A(P2_ADDR_REG_10__SCAN_IN), .B(P1_ADDR_REG_10__SCAN_IN), .Y(n1112));
  XOR2X1  g0079(.A(n1112), .B(n1070), .Y(ADD_1068_U63));
  XOR2X1  g0080(.A(P2_ADDR_REG_9__SCAN_IN), .B(P1_ADDR_REG_9__SCAN_IN), .Y(n1114));
  XOR2X1  g0081(.A(n1114), .B(n1068), .Y(ADD_1068_U47));
  XOR2X1  g0082(.A(P2_ADDR_REG_8__SCAN_IN), .B(P1_ADDR_REG_8__SCAN_IN), .Y(n1116));
  XOR2X1  g0083(.A(n1116), .B(n1066), .Y(ADD_1068_U48));
  XOR2X1  g0084(.A(P2_ADDR_REG_7__SCAN_IN), .B(P1_ADDR_REG_7__SCAN_IN), .Y(n1118));
  XOR2X1  g0085(.A(n1118), .B(n1064), .Y(ADD_1068_U49));
  XOR2X1  g0086(.A(P2_ADDR_REG_6__SCAN_IN), .B(P1_ADDR_REG_6__SCAN_IN), .Y(n1120));
  XOR2X1  g0087(.A(n1120), .B(n1062), .Y(ADD_1068_U50));
  XOR2X1  g0088(.A(P2_ADDR_REG_5__SCAN_IN), .B(P1_ADDR_REG_5__SCAN_IN), .Y(n1122));
  XOR2X1  g0089(.A(n1122), .B(n1060), .Y(ADD_1068_U51));
  XOR2X1  g0090(.A(P2_ADDR_REG_4__SCAN_IN), .B(P1_ADDR_REG_4__SCAN_IN), .Y(n1124));
  XOR2X1  g0091(.A(n1124), .B(n1058), .Y(ADD_1068_U52));
  XOR2X1  g0092(.A(P2_ADDR_REG_3__SCAN_IN), .B(P1_ADDR_REG_3__SCAN_IN), .Y(n1126));
  XOR2X1  g0093(.A(n1126), .B(n1056), .Y(ADD_1068_U53));
  XOR2X1  g0094(.A(P2_ADDR_REG_2__SCAN_IN), .B(P1_ADDR_REG_2__SCAN_IN), .Y(n1128));
  XOR2X1  g0095(.A(n1128), .B(n1054), .Y(ADD_1068_U54));
  NAND2X1 g0096(.A(P2_ADDR_REG_0__SCAN_IN), .B(P1_ADDR_REG_0__SCAN_IN), .Y(n1130));
  XOR2X1  g0097(.A(n1130), .B(P2_ADDR_REG_1__SCAN_IN), .Y(n1131));
  NOR2X1  g0098(.A(n1052), .B(n1051), .Y(n1132));
  INVX1   g0099(.A(P1_ADDR_REG_1__SCAN_IN), .Y(n1133));
  NOR2X1  g0100(.A(P2_ADDR_REG_1__SCAN_IN), .B(n1133), .Y(n1134));
  AOI21X1 g0101(.A0(n1134), .A1(n1130), .B0(n1132), .Y(n1135));
  OAI21X1 g0102(.A0(n1131), .A1(P1_ADDR_REG_1__SCAN_IN), .B0(n1135), .Y(ADD_1068_U5));
  XOR2X1  g0103(.A(P2_ADDR_REG_0__SCAN_IN), .B(P1_ADDR_REG_0__SCAN_IN), .Y(ADD_1068_U46));
  INVX1   g0104(.A(P2_RD_REG_SCAN_IN), .Y(n1138));
  XOR2X1  g0105(.A(P1_RD_REG_SCAN_IN), .B(n1138), .Y(U126));
  INVX1   g0106(.A(P2_WR_REG_SCAN_IN), .Y(n1140));
  XOR2X1  g0107(.A(P1_WR_REG_SCAN_IN), .B(n1140), .Y(U123));
  NAND3X1 g0108(.A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), .C(n1138), .Y(n1142));
  NOR2X1  g0109(.A(P2_ADDR_REG_19__SCAN_IN), .B(P1_RD_REG_SCAN_IN), .Y(n1143));
  NAND2X1 g0110(.A(n1143), .B(n1086), .Y(n1144));
  NAND2X1 g0111(.A(n1144), .B(n1142), .Y(n1145));
  INVX1   g0112(.A(P2_DATAO_REG_0__SCAN_IN), .Y(n1146));
  INVX1   g0113(.A(P2_ADDR_REG_19__SCAN_IN), .Y(n1147));
  NOR3X1  g0114(.A(n1147), .B(n1086), .C(P2_RD_REG_SCAN_IN), .Y(n1148));
  NOR3X1  g0115(.A(P2_ADDR_REG_19__SCAN_IN), .B(P1_RD_REG_SCAN_IN), .C(P1_ADDR_REG_19__SCAN_IN), .Y(n1149));
  NOR3X1  g0116(.A(n1149), .B(n1148), .C(n1146), .Y(n1150));
  INVX1   g0117(.A(SI_0_), .Y(n1151));
  NOR2X1  g0118(.A(n1149), .B(n1148), .Y(n1152));
  AOI21X1 g0119(.A0(n1144), .A1(n1142), .B0(n1146), .Y(n1153));
  AOI21X1 g0120(.A0(n1152), .A1(P1_DATAO_REG_0__SCAN_IN), .B0(n1153), .Y(n1154));
  XOR2X1  g0121(.A(n1154), .B(n1151), .Y(n1155));
  AOI21X1 g0122(.A0(n1155), .A1(n1145), .B0(n1150), .Y(n1156));
  INVX1   g0123(.A(P1_STATE_REG_SCAN_IN), .Y(P1_U3086));
  NOR2X1  g0124(.A(P1_U3086), .B(P1_IR_REG_31__SCAN_IN), .Y(n1158));
  OAI21X1 g0125(.A0(n1158), .A1(P1_STATE_REG_SCAN_IN), .B0(P1_IR_REG_0__SCAN_IN), .Y(n1159));
  OAI21X1 g0126(.A0(n1156), .A1(P1_STATE_REG_SCAN_IN), .B0(n1159), .Y(P1_U3355));
  INVX1   g0127(.A(P2_DATAO_REG_1__SCAN_IN), .Y(n1161));
  NOR3X1  g0128(.A(n1149), .B(n1148), .C(n1161), .Y(n1162));
  INVX1   g0129(.A(P1_DATAO_REG_1__SCAN_IN), .Y(n1163));
  OAI21X1 g0130(.A0(n1149), .A1(n1148), .B0(P2_DATAO_REG_1__SCAN_IN), .Y(n1164));
  OAI21X1 g0131(.A0(n1145), .A1(n1163), .B0(n1164), .Y(n1165));
  INVX1   g0132(.A(P1_DATAO_REG_0__SCAN_IN), .Y(n1166));
  OAI21X1 g0133(.A0(n1149), .A1(n1148), .B0(P2_DATAO_REG_0__SCAN_IN), .Y(n1167));
  OAI21X1 g0134(.A0(n1145), .A1(n1166), .B0(n1167), .Y(n1168));
  NAND2X1 g0135(.A(n1168), .B(SI_0_), .Y(n1169));
  XOR2X1  g0136(.A(n1169), .B(n1165), .Y(n1170));
  AOI21X1 g0137(.A0(n1144), .A1(n1142), .B0(n1161), .Y(n1171));
  AOI21X1 g0138(.A0(n1152), .A1(P1_DATAO_REG_1__SCAN_IN), .B0(n1171), .Y(n1172));
  INVX1   g0139(.A(SI_1_), .Y(n1173));
  NOR2X1  g0140(.A(n1151), .B(n1173), .Y(n1174));
  INVX1   g0141(.A(n1174), .Y(n1175));
  NOR3X1  g0142(.A(n1175), .B(n1172), .C(n1154), .Y(n1176));
  NOR2X1  g0143(.A(n1165), .B(n1173), .Y(n1177));
  AOI21X1 g0144(.A0(n1177), .A1(n1169), .B0(n1176), .Y(n1178));
  OAI21X1 g0145(.A0(n1170), .A1(SI_1_), .B0(n1178), .Y(n1179));
  AOI21X1 g0146(.A0(n1179), .A1(n1145), .B0(n1162), .Y(n1180));
  INVX1   g0147(.A(P1_IR_REG_31__SCAN_IN), .Y(n1181));
  NOR2X1  g0148(.A(P1_U3086), .B(n1181), .Y(n1182));
  XOR2X1  g0149(.A(P1_IR_REG_1__SCAN_IN), .B(P1_IR_REG_0__SCAN_IN), .Y(n1183));
  AOI22X1 g0150(.A0(n1182), .A1(n1183), .B0(n1158), .B1(P1_IR_REG_1__SCAN_IN), .Y(n1184));
  OAI21X1 g0151(.A0(n1180), .A1(P1_STATE_REG_SCAN_IN), .B0(n1184), .Y(P1_U3354));
  INVX1   g0152(.A(P2_DATAO_REG_2__SCAN_IN), .Y(n1186));
  NOR3X1  g0153(.A(n1149), .B(n1148), .C(n1186), .Y(n1187));
  NAND3X1 g0154(.A(n1165), .B(n1168), .C(SI_0_), .Y(n1188));
  AOI22X1 g0155(.A0(n1165), .A1(SI_1_), .B0(n1168), .B1(n1174), .Y(n1189));
  NAND2X1 g0156(.A(n1189), .B(n1188), .Y(n1190));
  INVX1   g0157(.A(SI_2_), .Y(n1191));
  AOI21X1 g0158(.A0(n1144), .A1(n1142), .B0(n1186), .Y(n1192));
  AOI21X1 g0159(.A0(n1152), .A1(P1_DATAO_REG_2__SCAN_IN), .B0(n1192), .Y(n1193));
  XOR2X1  g0160(.A(n1193), .B(n1191), .Y(n1194));
  XOR2X1  g0161(.A(n1194), .B(n1190), .Y(n1195));
  AOI21X1 g0162(.A0(n1195), .A1(n1145), .B0(n1187), .Y(n1196));
  INVX1   g0163(.A(P1_IR_REG_2__SCAN_IN), .Y(n1197));
  NOR2X1  g0164(.A(P1_IR_REG_1__SCAN_IN), .B(P1_IR_REG_0__SCAN_IN), .Y(n1198));
  XOR2X1  g0165(.A(n1198), .B(n1197), .Y(n1199));
  AOI22X1 g0166(.A0(n1182), .A1(n1199), .B0(n1158), .B1(P1_IR_REG_2__SCAN_IN), .Y(n1200));
  OAI21X1 g0167(.A0(n1196), .A1(P1_STATE_REG_SCAN_IN), .B0(n1200), .Y(P1_U3353));
  INVX1   g0168(.A(P2_DATAO_REG_3__SCAN_IN), .Y(n1202));
  NOR3X1  g0169(.A(n1149), .B(n1148), .C(n1202), .Y(n1203));
  NOR2X1  g0170(.A(n1193), .B(n1191), .Y(n1204));
  AOI22X1 g0171(.A0(n1189), .A1(n1188), .B0(n1191), .B1(n1193), .Y(n1205));
  NOR2X1  g0172(.A(n1205), .B(n1204), .Y(n1206));
  AOI21X1 g0173(.A0(n1144), .A1(n1142), .B0(n1202), .Y(n1207));
  AOI21X1 g0174(.A0(n1152), .A1(P1_DATAO_REG_3__SCAN_IN), .B0(n1207), .Y(n1208));
  XOR2X1  g0175(.A(n1208), .B(SI_3_), .Y(n1209));
  XOR2X1  g0176(.A(n1209), .B(n1206), .Y(n1210));
  AOI21X1 g0177(.A0(n1210), .A1(n1145), .B0(n1203), .Y(n1211));
  INVX1   g0178(.A(P1_IR_REG_3__SCAN_IN), .Y(n1212));
  NOR3X1  g0179(.A(P1_IR_REG_2__SCAN_IN), .B(P1_IR_REG_1__SCAN_IN), .C(P1_IR_REG_0__SCAN_IN), .Y(n1213));
  XOR2X1  g0180(.A(n1213), .B(n1212), .Y(n1214));
  AOI22X1 g0181(.A0(n1182), .A1(n1214), .B0(n1158), .B1(P1_IR_REG_3__SCAN_IN), .Y(n1215));
  OAI21X1 g0182(.A0(n1211), .A1(P1_STATE_REG_SCAN_IN), .B0(n1215), .Y(P1_U3352));
  INVX1   g0183(.A(P2_DATAO_REG_4__SCAN_IN), .Y(n1217));
  NOR3X1  g0184(.A(n1149), .B(n1148), .C(n1217), .Y(n1218));
  NOR3X1  g0185(.A(n1172), .B(n1154), .C(n1151), .Y(n1219));
  OAI22X1 g0186(.A0(n1172), .A1(n1173), .B0(n1154), .B1(n1175), .Y(n1220));
  INVX1   g0187(.A(SI_3_), .Y(n1221));
  AOI22X1 g0188(.A0(n1193), .A1(n1191), .B0(n1221), .B1(n1208), .Y(n1222));
  OAI21X1 g0189(.A0(n1220), .A1(n1219), .B0(n1222), .Y(n1223));
  NAND2X1 g0190(.A(n1208), .B(n1221), .Y(n1224));
  NOR2X1  g0191(.A(n1208), .B(n1221), .Y(n1225));
  AOI21X1 g0192(.A0(n1224), .A1(n1204), .B0(n1225), .Y(n1226));
  NAND2X1 g0193(.A(n1226), .B(n1223), .Y(n1227));
  INVX1   g0194(.A(SI_4_), .Y(n1228));
  INVX1   g0195(.A(P1_DATAO_REG_4__SCAN_IN), .Y(n1229));
  NOR3X1  g0196(.A(n1149), .B(n1148), .C(n1229), .Y(n1230));
  AOI21X1 g0197(.A0(n1144), .A1(n1142), .B0(n1217), .Y(n1231));
  NOR2X1  g0198(.A(n1231), .B(n1230), .Y(n1232));
  XOR2X1  g0199(.A(n1232), .B(n1228), .Y(n1233));
  XOR2X1  g0200(.A(n1233), .B(n1227), .Y(n1234));
  AOI21X1 g0201(.A0(n1234), .A1(n1145), .B0(n1218), .Y(n1235));
  NAND2X1 g0202(.A(n1213), .B(n1212), .Y(n1236));
  INVX1   g0203(.A(n1213), .Y(n1237));
  NOR3X1  g0204(.A(n1237), .B(P1_IR_REG_4__SCAN_IN), .C(P1_IR_REG_3__SCAN_IN), .Y(n1238));
  AOI21X1 g0205(.A0(n1236), .A1(P1_IR_REG_4__SCAN_IN), .B0(n1238), .Y(n1239));
  AOI22X1 g0206(.A0(n1182), .A1(n1239), .B0(n1158), .B1(P1_IR_REG_4__SCAN_IN), .Y(n1240));
  OAI21X1 g0207(.A0(n1235), .A1(P1_STATE_REG_SCAN_IN), .B0(n1240), .Y(P1_U3351));
  INVX1   g0208(.A(P2_DATAO_REG_5__SCAN_IN), .Y(n1242));
  NOR3X1  g0209(.A(n1149), .B(n1148), .C(n1242), .Y(n1243));
  NAND3X1 g0210(.A(n1144), .B(n1142), .C(P1_DATAO_REG_4__SCAN_IN), .Y(n1244));
  OAI21X1 g0211(.A0(n1149), .A1(n1148), .B0(P2_DATAO_REG_4__SCAN_IN), .Y(n1245));
  NAND3X1 g0212(.A(n1245), .B(n1244), .C(n1228), .Y(n1246));
  OAI21X1 g0213(.A0(n1231), .A1(n1230), .B0(SI_4_), .Y(n1247));
  INVX1   g0214(.A(n1247), .Y(n1248));
  AOI21X1 g0215(.A0(n1246), .A1(n1227), .B0(n1248), .Y(n1249));
  INVX1   g0216(.A(P1_DATAO_REG_5__SCAN_IN), .Y(n1250));
  NOR3X1  g0217(.A(n1149), .B(n1148), .C(n1250), .Y(n1251));
  AOI21X1 g0218(.A0(n1144), .A1(n1142), .B0(n1242), .Y(n1252));
  NOR2X1  g0219(.A(n1252), .B(n1251), .Y(n1253));
  XOR2X1  g0220(.A(n1253), .B(SI_5_), .Y(n1254));
  XOR2X1  g0221(.A(n1254), .B(n1249), .Y(n1255));
  AOI21X1 g0222(.A0(n1255), .A1(n1145), .B0(n1243), .Y(n1256));
  INVX1   g0223(.A(P1_IR_REG_5__SCAN_IN), .Y(n1257));
  XOR2X1  g0224(.A(n1238), .B(n1257), .Y(n1258));
  AOI22X1 g0225(.A0(n1182), .A1(n1258), .B0(n1158), .B1(P1_IR_REG_5__SCAN_IN), .Y(n1259));
  OAI21X1 g0226(.A0(n1256), .A1(P1_STATE_REG_SCAN_IN), .B0(n1259), .Y(P1_U3350));
  INVX1   g0227(.A(P2_DATAO_REG_6__SCAN_IN), .Y(n1261));
  NOR3X1  g0228(.A(n1149), .B(n1148), .C(n1261), .Y(n1262));
  NOR3X1  g0229(.A(n1252), .B(n1251), .C(SI_5_), .Y(n1263));
  OAI21X1 g0230(.A0(n1252), .A1(n1251), .B0(SI_5_), .Y(n1264));
  OAI21X1 g0231(.A0(n1263), .A1(n1247), .B0(n1264), .Y(n1265));
  NOR3X1  g0232(.A(n1231), .B(n1230), .C(SI_4_), .Y(n1266));
  NOR2X1  g0233(.A(n1263), .B(n1266), .Y(n1267));
  AOI21X1 g0234(.A0(n1267), .A1(n1227), .B0(n1265), .Y(n1268));
  INVX1   g0235(.A(P1_DATAO_REG_6__SCAN_IN), .Y(n1269));
  NOR3X1  g0236(.A(n1149), .B(n1148), .C(n1269), .Y(n1270));
  AOI21X1 g0237(.A0(n1144), .A1(n1142), .B0(n1261), .Y(n1271));
  NOR2X1  g0238(.A(n1271), .B(n1270), .Y(n1272));
  XOR2X1  g0239(.A(n1272), .B(SI_6_), .Y(n1273));
  XOR2X1  g0240(.A(n1273), .B(n1268), .Y(n1274));
  AOI21X1 g0241(.A0(n1274), .A1(n1145), .B0(n1262), .Y(n1275));
  INVX1   g0242(.A(P1_IR_REG_4__SCAN_IN), .Y(n1276));
  NAND4X1 g0243(.A(n1257), .B(n1276), .C(n1212), .D(n1213), .Y(n1277));
  INVX1   g0244(.A(P1_IR_REG_6__SCAN_IN), .Y(n1278));
  NAND2X1 g0245(.A(n1278), .B(n1257), .Y(n1279));
  NOR4X1  g0246(.A(n1237), .B(P1_IR_REG_4__SCAN_IN), .C(P1_IR_REG_3__SCAN_IN), .D(n1279), .Y(n1280));
  AOI21X1 g0247(.A0(n1277), .A1(P1_IR_REG_6__SCAN_IN), .B0(n1280), .Y(n1281));
  AOI22X1 g0248(.A0(n1182), .A1(n1281), .B0(n1158), .B1(P1_IR_REG_6__SCAN_IN), .Y(n1282));
  OAI21X1 g0249(.A0(n1275), .A1(P1_STATE_REG_SCAN_IN), .B0(n1282), .Y(P1_U3349));
  INVX1   g0250(.A(P2_DATAO_REG_7__SCAN_IN), .Y(n1284));
  NOR3X1  g0251(.A(n1149), .B(n1148), .C(n1284), .Y(n1285));
  INVX1   g0252(.A(P1_DATAO_REG_2__SCAN_IN), .Y(n1286));
  OAI21X1 g0253(.A0(n1149), .A1(n1148), .B0(P2_DATAO_REG_2__SCAN_IN), .Y(n1287));
  OAI21X1 g0254(.A0(n1145), .A1(n1286), .B0(n1287), .Y(n1288));
  INVX1   g0255(.A(P1_DATAO_REG_3__SCAN_IN), .Y(n1289));
  OAI21X1 g0256(.A0(n1149), .A1(n1148), .B0(P2_DATAO_REG_3__SCAN_IN), .Y(n1290));
  OAI21X1 g0257(.A0(n1145), .A1(n1289), .B0(n1290), .Y(n1291));
  OAI22X1 g0258(.A0(n1288), .A1(SI_2_), .B0(SI_3_), .B1(n1291), .Y(n1292));
  AOI21X1 g0259(.A0(n1189), .A1(n1188), .B0(n1292), .Y(n1293));
  NAND2X1 g0260(.A(n1288), .B(SI_2_), .Y(n1294));
  NOR2X1  g0261(.A(n1291), .B(SI_3_), .Y(n1295));
  NAND2X1 g0262(.A(n1291), .B(SI_3_), .Y(n1296));
  OAI21X1 g0263(.A0(n1295), .A1(n1294), .B0(n1296), .Y(n1297));
  NOR3X1  g0264(.A(n1271), .B(n1270), .C(SI_6_), .Y(n1298));
  NOR3X1  g0265(.A(n1298), .B(n1263), .C(n1266), .Y(n1299));
  OAI21X1 g0266(.A0(n1297), .A1(n1293), .B0(n1299), .Y(n1300));
  INVX1   g0267(.A(SI_6_), .Y(n1301));
  NAND3X1 g0268(.A(n1144), .B(n1142), .C(P1_DATAO_REG_6__SCAN_IN), .Y(n1302));
  OAI21X1 g0269(.A0(n1149), .A1(n1148), .B0(P2_DATAO_REG_6__SCAN_IN), .Y(n1303));
  NAND3X1 g0270(.A(n1303), .B(n1302), .C(n1301), .Y(n1304));
  AOI21X1 g0271(.A0(n1303), .A1(n1302), .B0(n1301), .Y(n1305));
  AOI21X1 g0272(.A0(n1304), .A1(n1265), .B0(n1305), .Y(n1306));
  NAND2X1 g0273(.A(n1306), .B(n1300), .Y(n1307));
  INVX1   g0274(.A(SI_7_), .Y(n1308));
  INVX1   g0275(.A(P1_DATAO_REG_7__SCAN_IN), .Y(n1309));
  NOR3X1  g0276(.A(n1149), .B(n1148), .C(n1309), .Y(n1310));
  AOI21X1 g0277(.A0(n1144), .A1(n1142), .B0(n1284), .Y(n1311));
  NOR2X1  g0278(.A(n1311), .B(n1310), .Y(n1312));
  XOR2X1  g0279(.A(n1312), .B(n1308), .Y(n1313));
  XOR2X1  g0280(.A(n1313), .B(n1307), .Y(n1314));
  AOI21X1 g0281(.A0(n1314), .A1(n1145), .B0(n1285), .Y(n1315));
  INVX1   g0282(.A(P1_IR_REG_7__SCAN_IN), .Y(n1316));
  XOR2X1  g0283(.A(n1280), .B(n1316), .Y(n1317));
  AOI22X1 g0284(.A0(n1182), .A1(n1317), .B0(n1158), .B1(P1_IR_REG_7__SCAN_IN), .Y(n1318));
  OAI21X1 g0285(.A0(n1315), .A1(P1_STATE_REG_SCAN_IN), .B0(n1318), .Y(P1_U3348));
  INVX1   g0286(.A(P2_DATAO_REG_8__SCAN_IN), .Y(n1320));
  NOR3X1  g0287(.A(n1149), .B(n1148), .C(n1320), .Y(n1321));
  NAND2X1 g0288(.A(n1304), .B(n1267), .Y(n1322));
  AOI21X1 g0289(.A0(n1226), .A1(n1223), .B0(n1322), .Y(n1323));
  NAND2X1 g0290(.A(n1304), .B(n1265), .Y(n1324));
  OAI21X1 g0291(.A0(n1272), .A1(n1301), .B0(n1324), .Y(n1325));
  NAND3X1 g0292(.A(n1144), .B(n1142), .C(P1_DATAO_REG_7__SCAN_IN), .Y(n1326));
  OAI21X1 g0293(.A0(n1149), .A1(n1148), .B0(P2_DATAO_REG_7__SCAN_IN), .Y(n1327));
  NAND2X1 g0294(.A(n1327), .B(n1326), .Y(n1328));
  OAI22X1 g0295(.A0(n1325), .A1(n1323), .B0(SI_7_), .B1(n1328), .Y(n1329));
  OAI21X1 g0296(.A0(n1312), .A1(n1308), .B0(n1329), .Y(n1330));
  INVX1   g0297(.A(SI_8_), .Y(n1331));
  AOI21X1 g0298(.A0(n1144), .A1(n1142), .B0(n1320), .Y(n1332));
  AOI21X1 g0299(.A0(n1152), .A1(P1_DATAO_REG_8__SCAN_IN), .B0(n1332), .Y(n1333));
  XOR2X1  g0300(.A(n1333), .B(n1331), .Y(n1334));
  XOR2X1  g0301(.A(n1334), .B(n1330), .Y(n1335));
  AOI21X1 g0302(.A0(n1335), .A1(n1145), .B0(n1321), .Y(n1336));
  INVX1   g0303(.A(P1_IR_REG_8__SCAN_IN), .Y(n1337));
  AOI21X1 g0304(.A0(n1280), .A1(n1316), .B0(n1337), .Y(n1338));
  NOR2X1  g0305(.A(P1_IR_REG_6__SCAN_IN), .B(P1_IR_REG_5__SCAN_IN), .Y(n1339));
  NAND3X1 g0306(.A(n1339), .B(n1276), .C(n1212), .Y(n1340));
  NOR4X1  g0307(.A(n1237), .B(P1_IR_REG_8__SCAN_IN), .C(P1_IR_REG_7__SCAN_IN), .D(n1340), .Y(n1341));
  NOR2X1  g0308(.A(n1341), .B(n1338), .Y(n1342));
  AOI22X1 g0309(.A0(n1182), .A1(n1342), .B0(n1158), .B1(P1_IR_REG_8__SCAN_IN), .Y(n1343));
  OAI21X1 g0310(.A0(n1336), .A1(P1_STATE_REG_SCAN_IN), .B0(n1343), .Y(P1_U3347));
  INVX1   g0311(.A(P2_DATAO_REG_9__SCAN_IN), .Y(n1345));
  NOR3X1  g0312(.A(n1149), .B(n1148), .C(n1345), .Y(n1346));
  AOI21X1 g0313(.A0(n1327), .A1(n1326), .B0(n1308), .Y(n1347));
  NAND3X1 g0314(.A(n1144), .B(n1142), .C(P1_DATAO_REG_8__SCAN_IN), .Y(n1348));
  OAI21X1 g0315(.A0(n1149), .A1(n1148), .B0(P2_DATAO_REG_8__SCAN_IN), .Y(n1349));
  NAND3X1 g0316(.A(n1349), .B(n1348), .C(n1331), .Y(n1350));
  AOI21X1 g0317(.A0(n1349), .A1(n1348), .B0(n1331), .Y(n1351));
  AOI21X1 g0318(.A0(n1350), .A1(n1347), .B0(n1351), .Y(n1352));
  INVX1   g0319(.A(n1352), .Y(n1353));
  AOI22X1 g0320(.A0(n1312), .A1(n1308), .B0(n1331), .B1(n1333), .Y(n1354));
  AOI21X1 g0321(.A0(n1354), .A1(n1307), .B0(n1353), .Y(n1355));
  AOI21X1 g0322(.A0(n1144), .A1(n1142), .B0(n1345), .Y(n1356));
  AOI21X1 g0323(.A0(n1152), .A1(P1_DATAO_REG_9__SCAN_IN), .B0(n1356), .Y(n1357));
  XOR2X1  g0324(.A(n1357), .B(SI_9_), .Y(n1358));
  XOR2X1  g0325(.A(n1358), .B(n1355), .Y(n1359));
  AOI21X1 g0326(.A0(n1359), .A1(n1145), .B0(n1346), .Y(n1360));
  INVX1   g0327(.A(P1_IR_REG_9__SCAN_IN), .Y(n1361));
  XOR2X1  g0328(.A(n1341), .B(n1361), .Y(n1362));
  AOI22X1 g0329(.A0(n1182), .A1(n1362), .B0(n1158), .B1(P1_IR_REG_9__SCAN_IN), .Y(n1363));
  OAI21X1 g0330(.A0(n1360), .A1(P1_STATE_REG_SCAN_IN), .B0(n1363), .Y(P1_U3346));
  INVX1   g0331(.A(P2_DATAO_REG_10__SCAN_IN), .Y(n1365));
  NOR3X1  g0332(.A(n1149), .B(n1148), .C(n1365), .Y(n1366));
  INVX1   g0333(.A(P1_DATAO_REG_9__SCAN_IN), .Y(n1367));
  OAI21X1 g0334(.A0(n1149), .A1(n1148), .B0(P2_DATAO_REG_9__SCAN_IN), .Y(n1368));
  OAI21X1 g0335(.A0(n1145), .A1(n1367), .B0(n1368), .Y(n1369));
  NOR2X1  g0336(.A(n1369), .B(SI_9_), .Y(n1370));
  NAND2X1 g0337(.A(n1369), .B(SI_9_), .Y(n1371));
  OAI21X1 g0338(.A0(n1370), .A1(n1352), .B0(n1371), .Y(n1372));
  OAI21X1 g0339(.A0(n1328), .A1(SI_7_), .B0(n1350), .Y(n1373));
  NOR2X1  g0340(.A(n1370), .B(n1373), .Y(n1374));
  AOI21X1 g0341(.A0(n1374), .A1(n1307), .B0(n1372), .Y(n1375));
  AOI21X1 g0342(.A0(n1144), .A1(n1142), .B0(n1365), .Y(n1376));
  AOI21X1 g0343(.A0(n1152), .A1(P1_DATAO_REG_10__SCAN_IN), .B0(n1376), .Y(n1377));
  XOR2X1  g0344(.A(n1377), .B(SI_10_), .Y(n1378));
  XOR2X1  g0345(.A(n1378), .B(n1375), .Y(n1379));
  AOI21X1 g0346(.A0(n1379), .A1(n1145), .B0(n1366), .Y(n1380));
  INVX1   g0347(.A(P1_IR_REG_10__SCAN_IN), .Y(n1381));
  AOI21X1 g0348(.A0(n1341), .A1(n1361), .B0(n1381), .Y(n1382));
  NOR2X1  g0349(.A(P1_IR_REG_10__SCAN_IN), .B(P1_IR_REG_9__SCAN_IN), .Y(n1383));
  AOI21X1 g0350(.A0(n1383), .A1(n1341), .B0(n1382), .Y(n1384));
  AOI22X1 g0351(.A0(n1182), .A1(n1384), .B0(n1158), .B1(P1_IR_REG_10__SCAN_IN), .Y(n1385));
  OAI21X1 g0352(.A0(n1380), .A1(P1_STATE_REG_SCAN_IN), .B0(n1385), .Y(P1_U3345));
  INVX1   g0353(.A(P2_DATAO_REG_11__SCAN_IN), .Y(n1387));
  NOR3X1  g0354(.A(n1149), .B(n1148), .C(n1387), .Y(n1388));
  INVX1   g0355(.A(P1_DATAO_REG_10__SCAN_IN), .Y(n1389));
  NOR3X1  g0356(.A(n1149), .B(n1148), .C(n1389), .Y(n1390));
  NOR3X1  g0357(.A(n1376), .B(n1390), .C(SI_10_), .Y(n1391));
  INVX1   g0358(.A(n1391), .Y(n1392));
  NAND2X1 g0359(.A(n1392), .B(n1374), .Y(n1393));
  AOI21X1 g0360(.A0(n1306), .A1(n1300), .B0(n1393), .Y(n1394));
  INVX1   g0361(.A(SI_10_), .Y(n1395));
  NAND2X1 g0362(.A(n1392), .B(n1372), .Y(n1396));
  OAI21X1 g0363(.A0(n1377), .A1(n1395), .B0(n1396), .Y(n1397));
  NOR2X1  g0364(.A(n1397), .B(n1394), .Y(n1398));
  AOI21X1 g0365(.A0(n1144), .A1(n1142), .B0(n1387), .Y(n1399));
  AOI21X1 g0366(.A0(n1152), .A1(P1_DATAO_REG_11__SCAN_IN), .B0(n1399), .Y(n1400));
  XOR2X1  g0367(.A(n1400), .B(SI_11_), .Y(n1401));
  XOR2X1  g0368(.A(n1401), .B(n1398), .Y(n1402));
  AOI21X1 g0369(.A0(n1402), .A1(n1145), .B0(n1388), .Y(n1403));
  INVX1   g0370(.A(P1_IR_REG_11__SCAN_IN), .Y(n1404));
  INVX1   g0371(.A(n1341), .Y(n1405));
  INVX1   g0372(.A(n1383), .Y(n1406));
  NOR2X1  g0373(.A(n1406), .B(n1405), .Y(n1407));
  XOR2X1  g0374(.A(n1407), .B(n1404), .Y(n1408));
  AOI22X1 g0375(.A0(n1182), .A1(n1408), .B0(n1158), .B1(P1_IR_REG_11__SCAN_IN), .Y(n1409));
  OAI21X1 g0376(.A0(n1403), .A1(P1_STATE_REG_SCAN_IN), .B0(n1409), .Y(P1_U3344));
  INVX1   g0377(.A(P2_DATAO_REG_12__SCAN_IN), .Y(n1411));
  NOR3X1  g0378(.A(n1149), .B(n1148), .C(n1411), .Y(n1412));
  INVX1   g0379(.A(SI_11_), .Y(n1413));
  INVX1   g0380(.A(P1_DATAO_REG_11__SCAN_IN), .Y(n1414));
  OAI21X1 g0381(.A0(n1149), .A1(n1148), .B0(P2_DATAO_REG_11__SCAN_IN), .Y(n1415));
  OAI21X1 g0382(.A0(n1145), .A1(n1414), .B0(n1415), .Y(n1416));
  OAI22X1 g0383(.A0(n1397), .A1(n1394), .B0(SI_11_), .B1(n1416), .Y(n1417));
  OAI21X1 g0384(.A0(n1400), .A1(n1413), .B0(n1417), .Y(n1418));
  INVX1   g0385(.A(SI_12_), .Y(n1419));
  AOI21X1 g0386(.A0(n1144), .A1(n1142), .B0(n1411), .Y(n1420));
  AOI21X1 g0387(.A0(n1152), .A1(P1_DATAO_REG_12__SCAN_IN), .B0(n1420), .Y(n1421));
  XOR2X1  g0388(.A(n1421), .B(n1419), .Y(n1422));
  XOR2X1  g0389(.A(n1422), .B(n1418), .Y(n1423));
  AOI21X1 g0390(.A0(n1423), .A1(n1145), .B0(n1412), .Y(n1424));
  NAND3X1 g0391(.A(n1383), .B(n1341), .C(n1404), .Y(n1425));
  NOR4X1  g0392(.A(n1405), .B(P1_IR_REG_12__SCAN_IN), .C(P1_IR_REG_11__SCAN_IN), .D(n1406), .Y(n1426));
  AOI21X1 g0393(.A0(n1425), .A1(P1_IR_REG_12__SCAN_IN), .B0(n1426), .Y(n1427));
  AOI22X1 g0394(.A0(n1182), .A1(n1427), .B0(n1158), .B1(P1_IR_REG_12__SCAN_IN), .Y(n1428));
  OAI21X1 g0395(.A0(n1424), .A1(P1_STATE_REG_SCAN_IN), .B0(n1428), .Y(P1_U3343));
  INVX1   g0396(.A(P2_DATAO_REG_13__SCAN_IN), .Y(n1430));
  NOR3X1  g0397(.A(n1149), .B(n1148), .C(n1430), .Y(n1431));
  NOR2X1  g0398(.A(n1400), .B(n1413), .Y(n1432));
  NAND2X1 g0399(.A(n1421), .B(n1419), .Y(n1433));
  NOR2X1  g0400(.A(n1421), .B(n1419), .Y(n1434));
  AOI21X1 g0401(.A0(n1433), .A1(n1432), .B0(n1434), .Y(n1435));
  OAI21X1 g0402(.A0(n1416), .A1(SI_11_), .B0(n1433), .Y(n1436));
  OAI21X1 g0403(.A0(n1436), .A1(n1398), .B0(n1435), .Y(n1437));
  INVX1   g0404(.A(P1_DATAO_REG_13__SCAN_IN), .Y(n1438));
  OAI21X1 g0405(.A0(n1149), .A1(n1148), .B0(P2_DATAO_REG_13__SCAN_IN), .Y(n1439));
  OAI21X1 g0406(.A0(n1145), .A1(n1438), .B0(n1439), .Y(n1440));
  XOR2X1  g0407(.A(n1440), .B(SI_13_), .Y(n1441));
  XOR2X1  g0408(.A(n1441), .B(n1437), .Y(n1442));
  AOI21X1 g0409(.A0(n1442), .A1(n1145), .B0(n1431), .Y(n1443));
  INVX1   g0410(.A(P1_IR_REG_13__SCAN_IN), .Y(n1444));
  XOR2X1  g0411(.A(n1426), .B(n1444), .Y(n1445));
  AOI22X1 g0412(.A0(n1182), .A1(n1445), .B0(n1158), .B1(P1_IR_REG_13__SCAN_IN), .Y(n1446));
  OAI21X1 g0413(.A0(n1443), .A1(P1_STATE_REG_SCAN_IN), .B0(n1446), .Y(P1_U3342));
  INVX1   g0414(.A(P2_DATAO_REG_14__SCAN_IN), .Y(n1448));
  NOR3X1  g0415(.A(n1149), .B(n1148), .C(n1448), .Y(n1449));
  NOR2X1  g0416(.A(n1440), .B(SI_13_), .Y(n1450));
  NOR2X1  g0417(.A(n1450), .B(n1435), .Y(n1451));
  AOI21X1 g0418(.A0(n1440), .A1(SI_13_), .B0(n1451), .Y(n1452));
  AOI22X1 g0419(.A0(n1400), .A1(n1413), .B0(n1419), .B1(n1421), .Y(n1453));
  OAI21X1 g0420(.A0(n1440), .A1(SI_13_), .B0(n1453), .Y(n1454));
  OAI21X1 g0421(.A0(n1454), .A1(n1398), .B0(n1452), .Y(n1455));
  INVX1   g0422(.A(SI_14_), .Y(n1456));
  AOI21X1 g0423(.A0(n1144), .A1(n1142), .B0(n1448), .Y(n1457));
  AOI21X1 g0424(.A0(n1152), .A1(P1_DATAO_REG_14__SCAN_IN), .B0(n1457), .Y(n1458));
  XOR2X1  g0425(.A(n1458), .B(n1456), .Y(n1459));
  XOR2X1  g0426(.A(n1459), .B(n1455), .Y(n1460));
  AOI21X1 g0427(.A0(n1460), .A1(n1145), .B0(n1449), .Y(n1461));
  INVX1   g0428(.A(P1_IR_REG_14__SCAN_IN), .Y(n1462));
  AOI21X1 g0429(.A0(n1426), .A1(n1444), .B0(n1462), .Y(n1463));
  INVX1   g0430(.A(n1426), .Y(n1464));
  NOR3X1  g0431(.A(n1464), .B(P1_IR_REG_14__SCAN_IN), .C(P1_IR_REG_13__SCAN_IN), .Y(n1465));
  NOR2X1  g0432(.A(n1465), .B(n1463), .Y(n1466));
  AOI22X1 g0433(.A0(n1182), .A1(n1466), .B0(n1158), .B1(P1_IR_REG_14__SCAN_IN), .Y(n1467));
  OAI21X1 g0434(.A0(n1461), .A1(P1_STATE_REG_SCAN_IN), .B0(n1467), .Y(P1_U3341));
  INVX1   g0435(.A(P2_DATAO_REG_15__SCAN_IN), .Y(n1469));
  NOR3X1  g0436(.A(n1149), .B(n1148), .C(n1469), .Y(n1470));
  NOR3X1  g0437(.A(n1391), .B(n1370), .C(n1373), .Y(n1471));
  OAI21X1 g0438(.A0(n1325), .A1(n1323), .B0(n1471), .Y(n1472));
  NOR2X1  g0439(.A(n1377), .B(n1395), .Y(n1473));
  AOI21X1 g0440(.A0(n1392), .A1(n1372), .B0(n1473), .Y(n1474));
  NOR2X1  g0441(.A(n1450), .B(n1436), .Y(n1475));
  NAND2X1 g0442(.A(n1458), .B(n1456), .Y(n1476));
  NAND2X1 g0443(.A(n1476), .B(n1475), .Y(n1477));
  AOI21X1 g0444(.A0(n1474), .A1(n1472), .B0(n1477), .Y(n1478));
  INVX1   g0445(.A(n1476), .Y(n1479));
  NOR2X1  g0446(.A(n1458), .B(n1456), .Y(n1480));
  INVX1   g0447(.A(n1480), .Y(n1481));
  OAI21X1 g0448(.A0(n1479), .A1(n1452), .B0(n1481), .Y(n1482));
  NOR2X1  g0449(.A(n1482), .B(n1478), .Y(n1483));
  AOI21X1 g0450(.A0(n1144), .A1(n1142), .B0(n1469), .Y(n1484));
  AOI21X1 g0451(.A0(n1152), .A1(P1_DATAO_REG_15__SCAN_IN), .B0(n1484), .Y(n1485));
  XOR2X1  g0452(.A(n1485), .B(SI_15_), .Y(n1486));
  XOR2X1  g0453(.A(n1486), .B(n1483), .Y(n1487));
  AOI21X1 g0454(.A0(n1487), .A1(n1145), .B0(n1470), .Y(n1488));
  INVX1   g0455(.A(P1_IR_REG_15__SCAN_IN), .Y(n1489));
  XOR2X1  g0456(.A(n1465), .B(n1489), .Y(n1490));
  AOI22X1 g0457(.A0(n1182), .A1(n1490), .B0(n1158), .B1(P1_IR_REG_15__SCAN_IN), .Y(n1491));
  OAI21X1 g0458(.A0(n1488), .A1(P1_STATE_REG_SCAN_IN), .B0(n1491), .Y(P1_U3340));
  INVX1   g0459(.A(P2_DATAO_REG_16__SCAN_IN), .Y(n1493));
  NOR3X1  g0460(.A(n1149), .B(n1148), .C(n1493), .Y(n1494));
  INVX1   g0461(.A(SI_15_), .Y(n1495));
  NOR2X1  g0462(.A(n1485), .B(n1495), .Y(n1496));
  NOR2X1  g0463(.A(n1479), .B(n1454), .Y(n1497));
  OAI21X1 g0464(.A0(n1397), .A1(n1394), .B0(n1497), .Y(n1498));
  NAND2X1 g0465(.A(n1440), .B(SI_13_), .Y(n1499));
  OAI21X1 g0466(.A0(n1450), .A1(n1435), .B0(n1499), .Y(n1500));
  AOI21X1 g0467(.A0(n1476), .A1(n1500), .B0(n1480), .Y(n1501));
  AOI22X1 g0468(.A0(n1501), .A1(n1498), .B0(n1495), .B1(n1485), .Y(n1502));
  NOR2X1  g0469(.A(n1502), .B(n1496), .Y(n1503));
  AOI21X1 g0470(.A0(n1144), .A1(n1142), .B0(n1493), .Y(n1504));
  AOI21X1 g0471(.A0(n1152), .A1(P1_DATAO_REG_16__SCAN_IN), .B0(n1504), .Y(n1505));
  XOR2X1  g0472(.A(n1505), .B(SI_16_), .Y(n1506));
  XOR2X1  g0473(.A(n1506), .B(n1503), .Y(n1507));
  AOI21X1 g0474(.A0(n1507), .A1(n1145), .B0(n1494), .Y(n1508));
  INVX1   g0475(.A(P1_IR_REG_16__SCAN_IN), .Y(n1509));
  NOR4X1  g0476(.A(P1_IR_REG_15__SCAN_IN), .B(P1_IR_REG_14__SCAN_IN), .C(P1_IR_REG_13__SCAN_IN), .D(n1464), .Y(n1510));
  NOR4X1  g0477(.A(P1_IR_REG_12__SCAN_IN), .B(P1_IR_REG_11__SCAN_IN), .C(P1_IR_REG_10__SCAN_IN), .D(P1_IR_REG_13__SCAN_IN), .Y(n1511));
  NAND2X1 g0478(.A(n1511), .B(n1462), .Y(n1512));
  NOR2X1  g0479(.A(P1_IR_REG_16__SCAN_IN), .B(P1_IR_REG_15__SCAN_IN), .Y(n1513));
  NAND3X1 g0480(.A(n1513), .B(n1198), .C(n1257), .Y(n1514));
  NOR4X1  g0481(.A(P1_IR_REG_8__SCAN_IN), .B(P1_IR_REG_7__SCAN_IN), .C(P1_IR_REG_6__SCAN_IN), .D(P1_IR_REG_9__SCAN_IN), .Y(n1515));
  INVX1   g0482(.A(n1515), .Y(n1516));
  NOR2X1  g0483(.A(P1_IR_REG_3__SCAN_IN), .B(P1_IR_REG_2__SCAN_IN), .Y(n1517));
  NAND2X1 g0484(.A(n1517), .B(n1276), .Y(n1518));
  NOR4X1  g0485(.A(n1516), .B(n1514), .C(n1512), .D(n1518), .Y(n1519));
  INVX1   g0486(.A(n1519), .Y(n1520));
  OAI21X1 g0487(.A0(n1510), .A1(n1509), .B0(n1520), .Y(n1521));
  INVX1   g0488(.A(n1521), .Y(n1522));
  AOI22X1 g0489(.A0(n1182), .A1(n1522), .B0(n1158), .B1(P1_IR_REG_16__SCAN_IN), .Y(n1523));
  OAI21X1 g0490(.A0(n1508), .A1(P1_STATE_REG_SCAN_IN), .B0(n1523), .Y(P1_U3339));
  INVX1   g0491(.A(P2_DATAO_REG_17__SCAN_IN), .Y(n1525));
  NOR3X1  g0492(.A(n1149), .B(n1148), .C(n1525), .Y(n1526));
  INVX1   g0493(.A(SI_16_), .Y(n1527));
  NOR2X1  g0494(.A(n1505), .B(n1527), .Y(n1528));
  INVX1   g0495(.A(n1496), .Y(n1529));
  NAND2X1 g0496(.A(n1485), .B(n1495), .Y(n1530));
  OAI21X1 g0497(.A0(n1482), .A1(n1478), .B0(n1530), .Y(n1531));
  AOI22X1 g0498(.A0(n1531), .A1(n1529), .B0(n1527), .B1(n1505), .Y(n1532));
  NOR2X1  g0499(.A(n1532), .B(n1528), .Y(n1533));
  AOI21X1 g0500(.A0(n1144), .A1(n1142), .B0(n1525), .Y(n1534));
  AOI21X1 g0501(.A0(n1152), .A1(P1_DATAO_REG_17__SCAN_IN), .B0(n1534), .Y(n1535));
  XOR2X1  g0502(.A(n1535), .B(SI_17_), .Y(n1536));
  XOR2X1  g0503(.A(n1536), .B(n1533), .Y(n1537));
  AOI21X1 g0504(.A0(n1537), .A1(n1145), .B0(n1526), .Y(n1538));
  INVX1   g0505(.A(P1_IR_REG_17__SCAN_IN), .Y(n1539));
  XOR2X1  g0506(.A(n1519), .B(n1539), .Y(n1540));
  AOI22X1 g0507(.A0(n1182), .A1(n1540), .B0(n1158), .B1(P1_IR_REG_17__SCAN_IN), .Y(n1541));
  OAI21X1 g0508(.A0(n1538), .A1(P1_STATE_REG_SCAN_IN), .B0(n1541), .Y(P1_U3338));
  INVX1   g0509(.A(P2_DATAO_REG_18__SCAN_IN), .Y(n1543));
  NOR3X1  g0510(.A(n1149), .B(n1148), .C(n1543), .Y(n1544));
  INVX1   g0511(.A(SI_17_), .Y(n1545));
  NOR2X1  g0512(.A(n1535), .B(n1545), .Y(n1546));
  INVX1   g0513(.A(n1528), .Y(n1547));
  INVX1   g0514(.A(n1505), .Y(n1548));
  OAI22X1 g0515(.A0(n1502), .A1(n1496), .B0(SI_16_), .B1(n1548), .Y(n1549));
  AOI22X1 g0516(.A0(n1549), .A1(n1547), .B0(n1545), .B1(n1535), .Y(n1550));
  NOR2X1  g0517(.A(n1550), .B(n1546), .Y(n1551));
  AOI21X1 g0518(.A0(n1144), .A1(n1142), .B0(n1543), .Y(n1552));
  AOI21X1 g0519(.A0(n1152), .A1(P1_DATAO_REG_18__SCAN_IN), .B0(n1552), .Y(n1553));
  XOR2X1  g0520(.A(n1553), .B(SI_18_), .Y(n1554));
  XOR2X1  g0521(.A(n1554), .B(n1551), .Y(n1555));
  AOI21X1 g0522(.A0(n1555), .A1(n1145), .B0(n1544), .Y(n1556));
  OAI21X1 g0523(.A0(n1520), .A1(P1_IR_REG_17__SCAN_IN), .B0(P1_IR_REG_18__SCAN_IN), .Y(n1557));
  NOR3X1  g0524(.A(P1_IR_REG_12__SCAN_IN), .B(P1_IR_REG_11__SCAN_IN), .C(P1_IR_REG_10__SCAN_IN), .Y(n1558));
  NAND2X1 g0525(.A(n1558), .B(n1444), .Y(n1559));
  NOR2X1  g0526(.A(n1559), .B(P1_IR_REG_14__SCAN_IN), .Y(n1560));
  INVX1   g0527(.A(P1_IR_REG_1__SCAN_IN), .Y(n1561));
  INVX1   g0528(.A(P1_IR_REG_18__SCAN_IN), .Y(n1562));
  NAND4X1 g0529(.A(n1539), .B(n1257), .C(n1561), .D(n1562), .Y(n1563));
  NOR3X1  g0530(.A(n1563), .B(P1_IR_REG_16__SCAN_IN), .C(P1_IR_REG_15__SCAN_IN), .Y(n1564));
  NOR4X1  g0531(.A(P1_IR_REG_3__SCAN_IN), .B(P1_IR_REG_2__SCAN_IN), .C(P1_IR_REG_0__SCAN_IN), .D(P1_IR_REG_4__SCAN_IN), .Y(n1565));
  NAND4X1 g0532(.A(n1564), .B(n1515), .C(n1560), .D(n1565), .Y(n1566));
  NAND2X1 g0533(.A(n1566), .B(n1557), .Y(n1567));
  INVX1   g0534(.A(n1567), .Y(n1568));
  AOI22X1 g0535(.A0(n1182), .A1(n1568), .B0(n1158), .B1(P1_IR_REG_18__SCAN_IN), .Y(n1569));
  OAI21X1 g0536(.A0(n1556), .A1(P1_STATE_REG_SCAN_IN), .B0(n1569), .Y(P1_U3337));
  INVX1   g0537(.A(P2_DATAO_REG_19__SCAN_IN), .Y(n1571));
  NOR3X1  g0538(.A(n1149), .B(n1148), .C(n1571), .Y(n1572));
  INVX1   g0539(.A(SI_18_), .Y(n1573));
  NOR2X1  g0540(.A(n1553), .B(n1573), .Y(n1574));
  INVX1   g0541(.A(n1546), .Y(n1575));
  INVX1   g0542(.A(n1535), .Y(n1576));
  OAI22X1 g0543(.A0(n1532), .A1(n1528), .B0(SI_17_), .B1(n1576), .Y(n1577));
  AOI22X1 g0544(.A0(n1577), .A1(n1575), .B0(n1573), .B1(n1553), .Y(n1578));
  NOR2X1  g0545(.A(n1578), .B(n1574), .Y(n1579));
  AOI21X1 g0546(.A0(n1144), .A1(n1142), .B0(n1571), .Y(n1580));
  AOI21X1 g0547(.A0(n1152), .A1(P1_DATAO_REG_19__SCAN_IN), .B0(n1580), .Y(n1581));
  XOR2X1  g0548(.A(n1581), .B(SI_19_), .Y(n1582));
  XOR2X1  g0549(.A(n1582), .B(n1579), .Y(n1583));
  AOI21X1 g0550(.A0(n1583), .A1(n1145), .B0(n1572), .Y(n1584));
  NOR4X1  g0551(.A(P1_IR_REG_9__SCAN_IN), .B(P1_IR_REG_8__SCAN_IN), .C(P1_IR_REG_7__SCAN_IN), .D(n1279), .Y(n1585));
  INVX1   g0552(.A(P1_IR_REG_19__SCAN_IN), .Y(n1586));
  NAND4X1 g0553(.A(n1562), .B(n1509), .C(n1276), .D(n1586), .Y(n1587));
  NOR4X1  g0554(.A(n1236), .B(P1_IR_REG_17__SCAN_IN), .C(P1_IR_REG_15__SCAN_IN), .D(n1587), .Y(n1588));
  NAND2X1 g0555(.A(n1588), .B(n1585), .Y(n1589));
  NOR2X1  g0556(.A(n1589), .B(n1512), .Y(n1590));
  AOI21X1 g0557(.A0(n1566), .A1(P1_IR_REG_19__SCAN_IN), .B0(n1590), .Y(n1591));
  AOI22X1 g0558(.A0(n1182), .A1(n1591), .B0(n1158), .B1(P1_IR_REG_19__SCAN_IN), .Y(n1592));
  OAI21X1 g0559(.A0(n1584), .A1(P1_STATE_REG_SCAN_IN), .B0(n1592), .Y(P1_U3336));
  INVX1   g0560(.A(P2_DATAO_REG_20__SCAN_IN), .Y(n1594));
  NOR3X1  g0561(.A(n1149), .B(n1148), .C(n1594), .Y(n1595));
  INVX1   g0562(.A(SI_19_), .Y(n1596));
  NOR2X1  g0563(.A(n1581), .B(n1596), .Y(n1597));
  INVX1   g0564(.A(n1574), .Y(n1598));
  INVX1   g0565(.A(n1553), .Y(n1599));
  OAI22X1 g0566(.A0(n1550), .A1(n1546), .B0(SI_18_), .B1(n1599), .Y(n1600));
  AOI22X1 g0567(.A0(n1600), .A1(n1598), .B0(n1596), .B1(n1581), .Y(n1601));
  NOR2X1  g0568(.A(n1601), .B(n1597), .Y(n1602));
  AOI21X1 g0569(.A0(n1144), .A1(n1142), .B0(n1594), .Y(n1603));
  AOI21X1 g0570(.A0(n1152), .A1(P1_DATAO_REG_20__SCAN_IN), .B0(n1603), .Y(n1604));
  XOR2X1  g0571(.A(n1604), .B(SI_20_), .Y(n1605));
  XOR2X1  g0572(.A(n1605), .B(n1602), .Y(n1606));
  AOI21X1 g0573(.A0(n1606), .A1(n1145), .B0(n1595), .Y(n1607));
  NAND3X1 g0574(.A(n1588), .B(n1585), .C(n1560), .Y(n1608));
  NAND4X1 g0575(.A(n1489), .B(n1462), .C(n1444), .D(n1558), .Y(n1609));
  INVX1   g0576(.A(P1_IR_REG_20__SCAN_IN), .Y(n1610));
  NAND2X1 g0577(.A(n1565), .B(n1610), .Y(n1611));
  NAND3X1 g0578(.A(n1562), .B(n1539), .C(n1561), .Y(n1612));
  NOR3X1  g0579(.A(n1612), .B(P1_IR_REG_19__SCAN_IN), .C(P1_IR_REG_16__SCAN_IN), .Y(n1613));
  NAND2X1 g0580(.A(n1613), .B(n1585), .Y(n1614));
  NOR3X1  g0581(.A(n1614), .B(n1611), .C(n1609), .Y(n1615));
  AOI21X1 g0582(.A0(n1608), .A1(P1_IR_REG_20__SCAN_IN), .B0(n1615), .Y(n1616));
  AOI22X1 g0583(.A0(n1182), .A1(n1616), .B0(n1158), .B1(P1_IR_REG_20__SCAN_IN), .Y(n1617));
  OAI21X1 g0584(.A0(n1607), .A1(P1_STATE_REG_SCAN_IN), .B0(n1617), .Y(P1_U3335));
  INVX1   g0585(.A(P2_DATAO_REG_21__SCAN_IN), .Y(n1619));
  NOR3X1  g0586(.A(n1149), .B(n1148), .C(n1619), .Y(n1620));
  INVX1   g0587(.A(SI_20_), .Y(n1621));
  NOR2X1  g0588(.A(n1604), .B(n1621), .Y(n1622));
  INVX1   g0589(.A(n1597), .Y(n1623));
  INVX1   g0590(.A(n1581), .Y(n1624));
  OAI22X1 g0591(.A0(n1578), .A1(n1574), .B0(SI_19_), .B1(n1624), .Y(n1625));
  AOI22X1 g0592(.A0(n1625), .A1(n1623), .B0(n1621), .B1(n1604), .Y(n1626));
  NOR2X1  g0593(.A(n1626), .B(n1622), .Y(n1627));
  AOI21X1 g0594(.A0(n1144), .A1(n1142), .B0(n1619), .Y(n1628));
  AOI21X1 g0595(.A0(n1152), .A1(P1_DATAO_REG_21__SCAN_IN), .B0(n1628), .Y(n1629));
  XOR2X1  g0596(.A(n1629), .B(SI_21_), .Y(n1630));
  XOR2X1  g0597(.A(n1630), .B(n1627), .Y(n1631));
  AOI21X1 g0598(.A0(n1631), .A1(n1145), .B0(n1620), .Y(n1632));
  INVX1   g0599(.A(P1_IR_REG_21__SCAN_IN), .Y(n1633));
  XOR2X1  g0600(.A(n1615), .B(n1633), .Y(n1634));
  AOI22X1 g0601(.A0(n1182), .A1(n1634), .B0(n1158), .B1(P1_IR_REG_21__SCAN_IN), .Y(n1635));
  OAI21X1 g0602(.A0(n1632), .A1(P1_STATE_REG_SCAN_IN), .B0(n1635), .Y(P1_U3334));
  INVX1   g0603(.A(P2_DATAO_REG_22__SCAN_IN), .Y(n1637));
  NOR3X1  g0604(.A(n1149), .B(n1148), .C(n1637), .Y(n1638));
  INVX1   g0605(.A(SI_21_), .Y(n1639));
  NOR2X1  g0606(.A(n1629), .B(n1639), .Y(n1640));
  INVX1   g0607(.A(n1622), .Y(n1641));
  INVX1   g0608(.A(n1604), .Y(n1642));
  OAI22X1 g0609(.A0(n1601), .A1(n1597), .B0(SI_20_), .B1(n1642), .Y(n1643));
  AOI22X1 g0610(.A0(n1643), .A1(n1641), .B0(n1639), .B1(n1629), .Y(n1644));
  NOR2X1  g0611(.A(n1644), .B(n1640), .Y(n1645));
  AOI21X1 g0612(.A0(n1144), .A1(n1142), .B0(n1637), .Y(n1646));
  AOI21X1 g0613(.A0(n1152), .A1(P1_DATAO_REG_22__SCAN_IN), .B0(n1646), .Y(n1647));
  XOR2X1  g0614(.A(n1647), .B(SI_22_), .Y(n1648));
  XOR2X1  g0615(.A(n1648), .B(n1645), .Y(n1649));
  AOI21X1 g0616(.A0(n1649), .A1(n1145), .B0(n1638), .Y(n1650));
  NOR3X1  g0617(.A(P1_IR_REG_21__SCAN_IN), .B(P1_IR_REG_20__SCAN_IN), .C(P1_IR_REG_0__SCAN_IN), .Y(n1651));
  NAND3X1 g0618(.A(n1651), .B(n1517), .C(n1276), .Y(n1652));
  NOR2X1  g0619(.A(n1652), .B(n1609), .Y(n1653));
  NAND3X1 g0620(.A(n1653), .B(n1613), .C(n1585), .Y(n1654));
  INVX1   g0621(.A(P1_IR_REG_22__SCAN_IN), .Y(n1655));
  NAND4X1 g0622(.A(n1633), .B(n1610), .C(n1586), .D(n1655), .Y(n1656));
  NOR3X1  g0623(.A(n1656), .B(P1_IR_REG_18__SCAN_IN), .C(P1_IR_REG_17__SCAN_IN), .Y(n1657));
  AOI22X1 g0624(.A0(n1654), .A1(P1_IR_REG_22__SCAN_IN), .B0(n1519), .B1(n1657), .Y(n1658));
  AOI22X1 g0625(.A0(n1182), .A1(n1658), .B0(n1158), .B1(P1_IR_REG_22__SCAN_IN), .Y(n1659));
  OAI21X1 g0626(.A0(n1650), .A1(P1_STATE_REG_SCAN_IN), .B0(n1659), .Y(P1_U3333));
  INVX1   g0627(.A(P2_DATAO_REG_23__SCAN_IN), .Y(n1661));
  NOR3X1  g0628(.A(n1149), .B(n1148), .C(n1661), .Y(n1662));
  INVX1   g0629(.A(SI_22_), .Y(n1663));
  NOR2X1  g0630(.A(n1647), .B(n1663), .Y(n1664));
  INVX1   g0631(.A(n1664), .Y(n1665));
  INVX1   g0632(.A(n1647), .Y(n1666));
  OAI22X1 g0633(.A0(n1644), .A1(n1640), .B0(SI_22_), .B1(n1666), .Y(n1667));
  NAND2X1 g0634(.A(n1667), .B(n1665), .Y(n1668));
  AOI21X1 g0635(.A0(n1144), .A1(n1142), .B0(n1661), .Y(n1669));
  AOI21X1 g0636(.A0(n1152), .A1(P1_DATAO_REG_23__SCAN_IN), .B0(n1669), .Y(n1670));
  XOR2X1  g0637(.A(n1670), .B(SI_23_), .Y(n1671));
  XOR2X1  g0638(.A(n1671), .B(n1668), .Y(n1672));
  NOR2X1  g0639(.A(n1672), .B(n1152), .Y(n1673));
  NOR2X1  g0640(.A(n1673), .B(n1662), .Y(n1674));
  INVX1   g0641(.A(P1_IR_REG_23__SCAN_IN), .Y(n1675));
  AOI21X1 g0642(.A0(n1657), .A1(n1519), .B0(n1675), .Y(n1676));
  NAND3X1 g0643(.A(n1655), .B(n1633), .C(n1610), .Y(n1677));
  NAND3X1 g0644(.A(n1586), .B(n1562), .C(n1509), .Y(n1678));
  NOR3X1  g0645(.A(n1678), .B(n1677), .C(n1609), .Y(n1679));
  NOR3X1  g0646(.A(P1_IR_REG_9__SCAN_IN), .B(P1_IR_REG_8__SCAN_IN), .C(P1_IR_REG_7__SCAN_IN), .Y(n1680));
  NAND3X1 g0647(.A(n1680), .B(n1339), .C(n1276), .Y(n1681));
  NAND4X1 g0648(.A(n1198), .B(n1675), .C(n1539), .D(n1517), .Y(n1682));
  NOR2X1  g0649(.A(n1682), .B(n1681), .Y(n1683));
  AOI21X1 g0650(.A0(n1683), .A1(n1679), .B0(n1676), .Y(n1684));
  AOI22X1 g0651(.A0(n1182), .A1(n1684), .B0(n1158), .B1(P1_IR_REG_23__SCAN_IN), .Y(n1685));
  OAI21X1 g0652(.A0(n1674), .A1(P1_STATE_REG_SCAN_IN), .B0(n1685), .Y(P1_U3332));
  INVX1   g0653(.A(P2_DATAO_REG_24__SCAN_IN), .Y(n1687));
  NOR3X1  g0654(.A(n1149), .B(n1148), .C(n1687), .Y(n1688));
  INVX1   g0655(.A(SI_23_), .Y(n1689));
  NOR2X1  g0656(.A(n1670), .B(n1689), .Y(n1690));
  AOI22X1 g0657(.A0(n1667), .A1(n1665), .B0(n1689), .B1(n1670), .Y(n1691));
  NOR2X1  g0658(.A(n1691), .B(n1690), .Y(n1692));
  AOI21X1 g0659(.A0(n1144), .A1(n1142), .B0(n1687), .Y(n1693));
  AOI21X1 g0660(.A0(n1152), .A1(P1_DATAO_REG_24__SCAN_IN), .B0(n1693), .Y(n1694));
  XOR2X1  g0661(.A(n1694), .B(SI_24_), .Y(n1695));
  XOR2X1  g0662(.A(n1695), .B(n1692), .Y(n1696));
  AOI21X1 g0663(.A0(n1696), .A1(n1145), .B0(n1688), .Y(n1697));
  INVX1   g0664(.A(P1_IR_REG_24__SCAN_IN), .Y(n1698));
  AOI21X1 g0665(.A0(n1683), .A1(n1679), .B0(n1698), .Y(n1699));
  NOR3X1  g0666(.A(P1_IR_REG_16__SCAN_IN), .B(P1_IR_REG_15__SCAN_IN), .C(P1_IR_REG_14__SCAN_IN), .Y(n1700));
  NOR4X1  g0667(.A(P1_IR_REG_19__SCAN_IN), .B(P1_IR_REG_18__SCAN_IN), .C(P1_IR_REG_17__SCAN_IN), .D(P1_IR_REG_20__SCAN_IN), .Y(n1701));
  NAND3X1 g0668(.A(n1701), .B(n1700), .C(n1198), .Y(n1702));
  NOR3X1  g0669(.A(P1_IR_REG_23__SCAN_IN), .B(P1_IR_REG_22__SCAN_IN), .C(P1_IR_REG_21__SCAN_IN), .Y(n1703));
  NAND3X1 g0670(.A(n1703), .B(n1517), .C(n1698), .Y(n1704));
  NOR4X1  g0671(.A(n1702), .B(n1681), .C(n1559), .D(n1704), .Y(n1705));
  NOR2X1  g0672(.A(n1705), .B(n1699), .Y(n1706));
  AOI22X1 g0673(.A0(n1182), .A1(n1706), .B0(n1158), .B1(P1_IR_REG_24__SCAN_IN), .Y(n1707));
  OAI21X1 g0674(.A0(n1697), .A1(P1_STATE_REG_SCAN_IN), .B0(n1707), .Y(P1_U3331));
  INVX1   g0675(.A(P2_DATAO_REG_25__SCAN_IN), .Y(n1709));
  NOR3X1  g0676(.A(n1149), .B(n1148), .C(n1709), .Y(n1710));
  INVX1   g0677(.A(SI_24_), .Y(n1711));
  NOR2X1  g0678(.A(n1694), .B(n1711), .Y(n1712));
  INVX1   g0679(.A(n1690), .Y(n1713));
  INVX1   g0680(.A(n1640), .Y(n1714));
  INVX1   g0681(.A(n1629), .Y(n1715));
  OAI22X1 g0682(.A0(n1626), .A1(n1622), .B0(SI_21_), .B1(n1715), .Y(n1716));
  AOI22X1 g0683(.A0(n1716), .A1(n1714), .B0(n1663), .B1(n1647), .Y(n1717));
  INVX1   g0684(.A(n1670), .Y(n1718));
  OAI22X1 g0685(.A0(n1717), .A1(n1664), .B0(SI_23_), .B1(n1718), .Y(n1719));
  AOI22X1 g0686(.A0(n1719), .A1(n1713), .B0(n1711), .B1(n1694), .Y(n1720));
  NOR2X1  g0687(.A(n1720), .B(n1712), .Y(n1721));
  AOI21X1 g0688(.A0(n1144), .A1(n1142), .B0(n1709), .Y(n1722));
  AOI21X1 g0689(.A0(n1152), .A1(P1_DATAO_REG_25__SCAN_IN), .B0(n1722), .Y(n1723));
  XOR2X1  g0690(.A(n1723), .B(SI_25_), .Y(n1724));
  XOR2X1  g0691(.A(n1724), .B(n1721), .Y(n1725));
  AOI21X1 g0692(.A0(n1725), .A1(n1145), .B0(n1710), .Y(n1726));
  INVX1   g0693(.A(P1_IR_REG_25__SCAN_IN), .Y(n1727));
  XOR2X1  g0694(.A(n1705), .B(n1727), .Y(n1728));
  AOI22X1 g0695(.A0(n1182), .A1(n1728), .B0(n1158), .B1(P1_IR_REG_25__SCAN_IN), .Y(n1729));
  OAI21X1 g0696(.A0(n1726), .A1(P1_STATE_REG_SCAN_IN), .B0(n1729), .Y(P1_U3330));
  INVX1   g0697(.A(P2_DATAO_REG_26__SCAN_IN), .Y(n1731));
  NOR3X1  g0698(.A(n1149), .B(n1148), .C(n1731), .Y(n1732));
  INVX1   g0699(.A(SI_25_), .Y(n1733));
  NOR2X1  g0700(.A(n1723), .B(n1733), .Y(n1734));
  INVX1   g0701(.A(n1712), .Y(n1735));
  INVX1   g0702(.A(n1694), .Y(n1736));
  OAI22X1 g0703(.A0(n1691), .A1(n1690), .B0(SI_24_), .B1(n1736), .Y(n1737));
  AOI22X1 g0704(.A0(n1737), .A1(n1735), .B0(n1733), .B1(n1723), .Y(n1738));
  NOR2X1  g0705(.A(n1738), .B(n1734), .Y(n1739));
  AOI21X1 g0706(.A0(n1144), .A1(n1142), .B0(n1731), .Y(n1740));
  AOI21X1 g0707(.A0(n1152), .A1(P1_DATAO_REG_26__SCAN_IN), .B0(n1740), .Y(n1741));
  XOR2X1  g0708(.A(n1741), .B(SI_26_), .Y(n1742));
  XOR2X1  g0709(.A(n1742), .B(n1739), .Y(n1743));
  AOI21X1 g0710(.A0(n1743), .A1(n1145), .B0(n1732), .Y(n1744));
  INVX1   g0711(.A(P1_IR_REG_26__SCAN_IN), .Y(n1745));
  NAND4X1 g0712(.A(n1517), .B(n1727), .C(n1698), .D(n1703), .Y(n1746));
  NOR4X1  g0713(.A(n1702), .B(n1681), .C(n1559), .D(n1746), .Y(n1747));
  NOR2X1  g0714(.A(n1747), .B(n1745), .Y(n1748));
  NOR4X1  g0715(.A(P1_IR_REG_18__SCAN_IN), .B(P1_IR_REG_17__SCAN_IN), .C(P1_IR_REG_1__SCAN_IN), .D(P1_IR_REG_19__SCAN_IN), .Y(n1749));
  NAND4X1 g0716(.A(n1700), .B(n1651), .C(n1511), .D(n1749), .Y(n1750));
  NOR4X1  g0717(.A(P1_IR_REG_24__SCAN_IN), .B(P1_IR_REG_23__SCAN_IN), .C(P1_IR_REG_22__SCAN_IN), .D(P1_IR_REG_25__SCAN_IN), .Y(n1751));
  NAND3X1 g0718(.A(n1751), .B(n1517), .C(n1745), .Y(n1752));
  NOR3X1  g0719(.A(n1752), .B(n1750), .C(n1681), .Y(n1753));
  NOR2X1  g0720(.A(n1753), .B(n1748), .Y(n1754));
  AOI22X1 g0721(.A0(n1182), .A1(n1754), .B0(n1158), .B1(P1_IR_REG_26__SCAN_IN), .Y(n1755));
  OAI21X1 g0722(.A0(n1744), .A1(P1_STATE_REG_SCAN_IN), .B0(n1755), .Y(P1_U3329));
  INVX1   g0723(.A(P2_DATAO_REG_27__SCAN_IN), .Y(n1757));
  NOR3X1  g0724(.A(n1149), .B(n1148), .C(n1757), .Y(n1758));
  INVX1   g0725(.A(SI_26_), .Y(n1759));
  NOR2X1  g0726(.A(n1741), .B(n1759), .Y(n1760));
  INVX1   g0727(.A(n1760), .Y(n1761));
  INVX1   g0728(.A(n1741), .Y(n1762));
  OAI22X1 g0729(.A0(n1738), .A1(n1734), .B0(SI_26_), .B1(n1762), .Y(n1763));
  AOI21X1 g0730(.A0(n1144), .A1(n1142), .B0(n1757), .Y(n1764));
  AOI21X1 g0731(.A0(n1152), .A1(P1_DATAO_REG_27__SCAN_IN), .B0(n1764), .Y(n1765));
  XOR2X1  g0732(.A(n1765), .B(SI_27_), .Y(n1766));
  INVX1   g0733(.A(n1766), .Y(n1767));
  NAND3X1 g0734(.A(n1767), .B(n1763), .C(n1761), .Y(n1768));
  INVX1   g0735(.A(n1734), .Y(n1769));
  INVX1   g0736(.A(n1723), .Y(n1770));
  OAI22X1 g0737(.A0(n1720), .A1(n1712), .B0(SI_25_), .B1(n1770), .Y(n1771));
  AOI22X1 g0738(.A0(n1771), .A1(n1769), .B0(n1759), .B1(n1741), .Y(n1772));
  OAI21X1 g0739(.A0(n1772), .A1(n1760), .B0(n1766), .Y(n1773));
  AOI21X1 g0740(.A0(n1773), .A1(n1768), .B0(n1152), .Y(n1774));
  NOR2X1  g0741(.A(n1774), .B(n1758), .Y(n1775));
  XOR2X1  g0742(.A(n1753), .B(P1_IR_REG_27__SCAN_IN), .Y(n1776));
  INVX1   g0743(.A(n1776), .Y(n1777));
  AOI22X1 g0744(.A0(n1182), .A1(n1777), .B0(n1158), .B1(P1_IR_REG_27__SCAN_IN), .Y(n1778));
  OAI21X1 g0745(.A0(n1775), .A1(P1_STATE_REG_SCAN_IN), .B0(n1778), .Y(P1_U3328));
  INVX1   g0746(.A(P2_DATAO_REG_28__SCAN_IN), .Y(n1780));
  NOR3X1  g0747(.A(n1149), .B(n1148), .C(n1780), .Y(n1781));
  INVX1   g0748(.A(SI_27_), .Y(n1782));
  NOR2X1  g0749(.A(n1765), .B(n1782), .Y(n1783));
  AOI22X1 g0750(.A0(n1763), .A1(n1761), .B0(n1782), .B1(n1765), .Y(n1784));
  NOR2X1  g0751(.A(n1784), .B(n1783), .Y(n1785));
  AOI21X1 g0752(.A0(n1144), .A1(n1142), .B0(n1780), .Y(n1786));
  AOI21X1 g0753(.A0(n1152), .A1(P1_DATAO_REG_28__SCAN_IN), .B0(n1786), .Y(n1787));
  XOR2X1  g0754(.A(n1787), .B(SI_28_), .Y(n1788));
  XOR2X1  g0755(.A(n1788), .B(n1785), .Y(n1789));
  AOI21X1 g0756(.A0(n1789), .A1(n1145), .B0(n1781), .Y(n1790));
  INVX1   g0757(.A(P1_IR_REG_28__SCAN_IN), .Y(n1791));
  NAND4X1 g0758(.A(n1339), .B(n1276), .C(n1212), .D(n1680), .Y(n1792));
  INVX1   g0759(.A(P1_IR_REG_27__SCAN_IN), .Y(n1793));
  NAND4X1 g0760(.A(n1793), .B(n1745), .C(n1197), .D(n1751), .Y(n1794));
  NOR3X1  g0761(.A(n1794), .B(n1792), .C(n1750), .Y(n1795));
  NAND4X1 g0762(.A(n1586), .B(n1562), .C(n1539), .D(n1198), .Y(n1796));
  NAND4X1 g0763(.A(n1655), .B(n1633), .C(n1610), .D(n1700), .Y(n1797));
  NOR3X1  g0764(.A(n1797), .B(n1796), .C(n1559), .Y(n1798));
  NAND4X1 g0765(.A(n1727), .B(n1698), .C(n1675), .D(n1745), .Y(n1799));
  NAND3X1 g0766(.A(n1791), .B(n1793), .C(n1197), .Y(n1800));
  NOR3X1  g0767(.A(n1800), .B(n1799), .C(n1792), .Y(n1801));
  NAND2X1 g0768(.A(n1801), .B(n1798), .Y(n1802));
  OAI21X1 g0769(.A0(n1795), .A1(n1791), .B0(n1802), .Y(n1803));
  NOR3X1  g0770(.A(n1803), .B(P1_U3086), .C(n1181), .Y(n1804));
  AOI21X1 g0771(.A0(n1158), .A1(P1_IR_REG_28__SCAN_IN), .B0(n1804), .Y(n1805));
  OAI21X1 g0772(.A0(n1790), .A1(P1_STATE_REG_SCAN_IN), .B0(n1805), .Y(P1_U3327));
  INVX1   g0773(.A(P2_DATAO_REG_29__SCAN_IN), .Y(n1807));
  NOR3X1  g0774(.A(n1149), .B(n1148), .C(n1807), .Y(n1808));
  INVX1   g0775(.A(SI_28_), .Y(n1809));
  NOR2X1  g0776(.A(n1787), .B(n1809), .Y(n1810));
  INVX1   g0777(.A(n1783), .Y(n1811));
  INVX1   g0778(.A(n1765), .Y(n1812));
  OAI22X1 g0779(.A0(n1772), .A1(n1760), .B0(SI_27_), .B1(n1812), .Y(n1813));
  AOI22X1 g0780(.A0(n1813), .A1(n1811), .B0(n1809), .B1(n1787), .Y(n1814));
  NOR2X1  g0781(.A(n1814), .B(n1810), .Y(n1815));
  AOI21X1 g0782(.A0(n1144), .A1(n1142), .B0(n1807), .Y(n1816));
  AOI21X1 g0783(.A0(n1152), .A1(P1_DATAO_REG_29__SCAN_IN), .B0(n1816), .Y(n1817));
  XOR2X1  g0784(.A(n1817), .B(SI_29_), .Y(n1818));
  XOR2X1  g0785(.A(n1818), .B(n1815), .Y(n1819));
  AOI21X1 g0786(.A0(n1819), .A1(n1145), .B0(n1808), .Y(n1820));
  NAND2X1 g0787(.A(n1802), .B(P1_IR_REG_29__SCAN_IN), .Y(n1821));
  NOR4X1  g0788(.A(n1799), .B(n1792), .C(P1_IR_REG_29__SCAN_IN), .D(n1800), .Y(n1822));
  NAND2X1 g0789(.A(n1822), .B(n1798), .Y(n1823));
  NAND2X1 g0790(.A(n1823), .B(n1821), .Y(n1824));
  NOR3X1  g0791(.A(n1824), .B(P1_U3086), .C(n1181), .Y(n1825));
  AOI21X1 g0792(.A0(n1158), .A1(P1_IR_REG_29__SCAN_IN), .B0(n1825), .Y(n1826));
  OAI21X1 g0793(.A0(n1820), .A1(P1_STATE_REG_SCAN_IN), .B0(n1826), .Y(P1_U3326));
  INVX1   g0794(.A(P2_DATAO_REG_30__SCAN_IN), .Y(n1828));
  NOR3X1  g0795(.A(n1149), .B(n1148), .C(n1828), .Y(n1829));
  INVX1   g0796(.A(SI_29_), .Y(n1830));
  NOR2X1  g0797(.A(n1817), .B(n1830), .Y(n1831));
  INVX1   g0798(.A(n1831), .Y(n1832));
  INVX1   g0799(.A(n1817), .Y(n1833));
  OAI22X1 g0800(.A0(n1814), .A1(n1810), .B0(SI_29_), .B1(n1833), .Y(n1834));
  AOI21X1 g0801(.A0(n1144), .A1(n1142), .B0(n1828), .Y(n1835));
  AOI21X1 g0802(.A0(n1152), .A1(P1_DATAO_REG_30__SCAN_IN), .B0(n1835), .Y(n1836));
  XOR2X1  g0803(.A(n1836), .B(SI_30_), .Y(n1837));
  INVX1   g0804(.A(n1837), .Y(n1838));
  NAND3X1 g0805(.A(n1838), .B(n1834), .C(n1832), .Y(n1839));
  INVX1   g0806(.A(n1810), .Y(n1840));
  INVX1   g0807(.A(n1787), .Y(n1841));
  OAI22X1 g0808(.A0(n1784), .A1(n1783), .B0(SI_28_), .B1(n1841), .Y(n1842));
  AOI22X1 g0809(.A0(n1842), .A1(n1840), .B0(n1830), .B1(n1817), .Y(n1843));
  OAI21X1 g0810(.A0(n1843), .A1(n1831), .B0(n1837), .Y(n1844));
  AOI21X1 g0811(.A0(n1844), .A1(n1839), .B0(n1152), .Y(n1845));
  NOR2X1  g0812(.A(n1845), .B(n1829), .Y(n1846));
  XOR2X1  g0813(.A(n1823), .B(P1_IR_REG_30__SCAN_IN), .Y(n1847));
  AOI22X1 g0814(.A0(n1182), .A1(n1847), .B0(n1158), .B1(P1_IR_REG_30__SCAN_IN), .Y(n1848));
  OAI21X1 g0815(.A0(n1846), .A1(P1_STATE_REG_SCAN_IN), .B0(n1848), .Y(P1_U3325));
  INVX1   g0816(.A(P2_DATAO_REG_31__SCAN_IN), .Y(n1850));
  NOR3X1  g0817(.A(n1149), .B(n1148), .C(n1850), .Y(n1851));
  INVX1   g0818(.A(SI_30_), .Y(n1852));
  AOI21X1 g0819(.A0(n1144), .A1(n1142), .B0(n1850), .Y(n1853));
  AOI21X1 g0820(.A0(n1152), .A1(P1_DATAO_REG_31__SCAN_IN), .B0(n1853), .Y(n1854));
  XOR2X1  g0821(.A(n1854), .B(SI_31_), .Y(n1855));
  AOI21X1 g0822(.A0(n1836), .A1(n1852), .B0(n1855), .Y(n1856));
  INVX1   g0823(.A(n1856), .Y(n1857));
  AOI21X1 g0824(.A0(n1834), .A1(n1832), .B0(n1857), .Y(n1858));
  NOR2X1  g0825(.A(n1836), .B(n1852), .Y(n1859));
  INVX1   g0826(.A(n1859), .Y(n1860));
  NAND3X1 g0827(.A(n1860), .B(n1855), .C(n1832), .Y(n1861));
  NAND3X1 g0828(.A(n1855), .B(n1836), .C(n1852), .Y(n1862));
  OAI21X1 g0829(.A0(n1860), .A1(n1855), .B0(n1862), .Y(n1863));
  INVX1   g0830(.A(n1863), .Y(n1864));
  OAI21X1 g0831(.A0(n1861), .A1(n1843), .B0(n1864), .Y(n1865));
  NOR3X1  g0832(.A(n1865), .B(n1858), .C(n1152), .Y(n1866));
  OAI21X1 g0833(.A0(n1866), .A1(n1851), .B0(P1_U3086), .Y(n1867));
  NOR2X1  g0834(.A(n1823), .B(P1_IR_REG_30__SCAN_IN), .Y(n1868));
  NAND3X1 g0835(.A(n1868), .B(P1_STATE_REG_SCAN_IN), .C(P1_IR_REG_31__SCAN_IN), .Y(n1869));
  NAND2X1 g0836(.A(n1869), .B(n1867), .Y(P1_U3324));
  NOR2X1  g0837(.A(P1_IR_REG_31__SCAN_IN), .B(n1675), .Y(n1871));
  AOI21X1 g0838(.A0(n1684), .A1(P1_IR_REG_31__SCAN_IN), .B0(n1871), .Y(n1872));
  INVX1   g0839(.A(n1872), .Y(n1873));
  NAND2X1 g0840(.A(n1706), .B(P1_IR_REG_31__SCAN_IN), .Y(n1874));
  OAI21X1 g0841(.A0(P1_IR_REG_31__SCAN_IN), .A1(n1698), .B0(n1874), .Y(n1875));
  INVX1   g0842(.A(n1875), .Y(n1876));
  NAND2X1 g0843(.A(n1754), .B(P1_IR_REG_31__SCAN_IN), .Y(n1877));
  OAI21X1 g0844(.A0(P1_IR_REG_31__SCAN_IN), .A1(n1745), .B0(n1877), .Y(n1878));
  INVX1   g0845(.A(n1878), .Y(n1879));
  NOR2X1  g0846(.A(P1_IR_REG_31__SCAN_IN), .B(n1727), .Y(n1880));
  AOI21X1 g0847(.A0(n1728), .A1(P1_IR_REG_31__SCAN_IN), .B0(n1880), .Y(n1881));
  NOR3X1  g0848(.A(n1881), .B(n1879), .C(n1876), .Y(n1882));
  INVX1   g0849(.A(P1_B_REG_SCAN_IN), .Y(n1883));
  INVX1   g0850(.A(n1881), .Y(n1884));
  NOR4X1  g0851(.A(n1879), .B(n1875), .C(n1883), .D(n1884), .Y(n1885));
  OAI21X1 g0852(.A0(n1876), .A1(P1_B_REG_SCAN_IN), .B0(n1878), .Y(n1886));
  NOR2X1  g0853(.A(n1886), .B(n1885), .Y(n1887));
  NOR4X1  g0854(.A(n1882), .B(n1873), .C(P1_U3086), .D(n1887), .Y(n1888));
  OAI21X1 g0855(.A0(n1884), .A1(n1879), .B0(n1876), .Y(n1889));
  NAND2X1 g0856(.A(n1889), .B(n1888), .Y(n1890));
  NOR3X1  g0857(.A(n1882), .B(n1873), .C(P1_U3086), .Y(n1891));
  INVX1   g0858(.A(n1891), .Y(n1892));
  OAI21X1 g0859(.A0(n1887), .A1(n1892), .B0(P1_D_REG_0__SCAN_IN), .Y(n1893));
  NAND2X1 g0860(.A(n1893), .B(n1890), .Y(P1_U3439));
  OAI21X1 g0861(.A0(n1884), .A1(n1878), .B0(n1888), .Y(n1895));
  OAI21X1 g0862(.A0(n1887), .A1(n1892), .B0(P1_D_REG_1__SCAN_IN), .Y(n1896));
  NAND2X1 g0863(.A(n1896), .B(n1895), .Y(P1_U3440));
  INVX1   g0864(.A(P1_D_REG_2__SCAN_IN), .Y(n1898));
  NOR2X1  g0865(.A(n1888), .B(n1898), .Y(P1_U3323));
  INVX1   g0866(.A(P1_D_REG_3__SCAN_IN), .Y(n1900));
  NOR2X1  g0867(.A(n1888), .B(n1900), .Y(P1_U3322));
  INVX1   g0868(.A(P1_D_REG_4__SCAN_IN), .Y(n1902));
  NOR2X1  g0869(.A(n1888), .B(n1902), .Y(P1_U3321));
  INVX1   g0870(.A(P1_D_REG_5__SCAN_IN), .Y(n1904));
  NOR2X1  g0871(.A(n1888), .B(n1904), .Y(P1_U3320));
  INVX1   g0872(.A(P1_D_REG_6__SCAN_IN), .Y(n1906));
  NOR2X1  g0873(.A(n1888), .B(n1906), .Y(P1_U3319));
  INVX1   g0874(.A(P1_D_REG_7__SCAN_IN), .Y(n1908));
  NOR2X1  g0875(.A(n1888), .B(n1908), .Y(P1_U3318));
  INVX1   g0876(.A(P1_D_REG_8__SCAN_IN), .Y(n1910));
  NOR2X1  g0877(.A(n1888), .B(n1910), .Y(P1_U3317));
  INVX1   g0878(.A(P1_D_REG_9__SCAN_IN), .Y(n1912));
  NOR2X1  g0879(.A(n1888), .B(n1912), .Y(P1_U3316));
  INVX1   g0880(.A(P1_D_REG_10__SCAN_IN), .Y(n1914));
  NOR2X1  g0881(.A(n1888), .B(n1914), .Y(P1_U3315));
  INVX1   g0882(.A(P1_D_REG_11__SCAN_IN), .Y(n1916));
  NOR2X1  g0883(.A(n1888), .B(n1916), .Y(P1_U3314));
  INVX1   g0884(.A(P1_D_REG_12__SCAN_IN), .Y(n1918));
  NOR2X1  g0885(.A(n1888), .B(n1918), .Y(P1_U3313));
  INVX1   g0886(.A(P1_D_REG_13__SCAN_IN), .Y(n1920));
  NOR2X1  g0887(.A(n1888), .B(n1920), .Y(P1_U3312));
  INVX1   g0888(.A(P1_D_REG_14__SCAN_IN), .Y(n1922));
  NOR2X1  g0889(.A(n1888), .B(n1922), .Y(P1_U3311));
  INVX1   g0890(.A(P1_D_REG_15__SCAN_IN), .Y(n1924));
  NOR2X1  g0891(.A(n1888), .B(n1924), .Y(P1_U3310));
  INVX1   g0892(.A(P1_D_REG_16__SCAN_IN), .Y(n1926));
  NOR2X1  g0893(.A(n1888), .B(n1926), .Y(P1_U3309));
  INVX1   g0894(.A(P1_D_REG_17__SCAN_IN), .Y(n1928));
  NOR2X1  g0895(.A(n1888), .B(n1928), .Y(P1_U3308));
  INVX1   g0896(.A(P1_D_REG_18__SCAN_IN), .Y(n1930));
  NOR2X1  g0897(.A(n1888), .B(n1930), .Y(P1_U3307));
  INVX1   g0898(.A(P1_D_REG_19__SCAN_IN), .Y(n1932));
  NOR2X1  g0899(.A(n1888), .B(n1932), .Y(P1_U3306));
  INVX1   g0900(.A(P1_D_REG_20__SCAN_IN), .Y(n1934));
  NOR2X1  g0901(.A(n1888), .B(n1934), .Y(P1_U3305));
  INVX1   g0902(.A(P1_D_REG_21__SCAN_IN), .Y(n1936));
  NOR2X1  g0903(.A(n1888), .B(n1936), .Y(P1_U3304));
  INVX1   g0904(.A(P1_D_REG_22__SCAN_IN), .Y(n1938));
  NOR2X1  g0905(.A(n1888), .B(n1938), .Y(P1_U3303));
  INVX1   g0906(.A(P1_D_REG_23__SCAN_IN), .Y(n1940));
  NOR2X1  g0907(.A(n1888), .B(n1940), .Y(P1_U3302));
  INVX1   g0908(.A(P1_D_REG_24__SCAN_IN), .Y(n1942));
  NOR2X1  g0909(.A(n1888), .B(n1942), .Y(P1_U3301));
  INVX1   g0910(.A(P1_D_REG_25__SCAN_IN), .Y(n1944));
  NOR2X1  g0911(.A(n1888), .B(n1944), .Y(P1_U3300));
  INVX1   g0912(.A(P1_D_REG_26__SCAN_IN), .Y(n1946));
  NOR2X1  g0913(.A(n1888), .B(n1946), .Y(P1_U3299));
  INVX1   g0914(.A(P1_D_REG_27__SCAN_IN), .Y(n1948));
  NOR2X1  g0915(.A(n1888), .B(n1948), .Y(P1_U3298));
  INVX1   g0916(.A(P1_D_REG_28__SCAN_IN), .Y(n1950));
  NOR2X1  g0917(.A(n1888), .B(n1950), .Y(P1_U3297));
  INVX1   g0918(.A(P1_D_REG_29__SCAN_IN), .Y(n1952));
  NOR2X1  g0919(.A(n1888), .B(n1952), .Y(P1_U3296));
  INVX1   g0920(.A(P1_D_REG_30__SCAN_IN), .Y(n1954));
  NOR2X1  g0921(.A(n1888), .B(n1954), .Y(P1_U3295));
  INVX1   g0922(.A(P1_D_REG_31__SCAN_IN), .Y(n1956));
  NOR2X1  g0923(.A(n1888), .B(n1956), .Y(P1_U3294));
  OAI21X1 g0924(.A0(P1_D_REG_7__SCAN_IN), .A1(P1_D_REG_3__SCAN_IN), .B0(n1887), .Y(n1958));
  OAI21X1 g0925(.A0(P1_D_REG_9__SCAN_IN), .A1(P1_D_REG_8__SCAN_IN), .B0(n1887), .Y(n1959));
  OAI21X1 g0926(.A0(P1_D_REG_10__SCAN_IN), .A1(P1_D_REG_5__SCAN_IN), .B0(n1887), .Y(n1960));
  OAI21X1 g0927(.A0(P1_D_REG_6__SCAN_IN), .A1(P1_D_REG_4__SCAN_IN), .B0(n1887), .Y(n1961));
  NAND4X1 g0928(.A(n1960), .B(n1959), .C(n1958), .D(n1961), .Y(n1962));
  OAI21X1 g0929(.A0(P1_D_REG_28__SCAN_IN), .A1(P1_D_REG_27__SCAN_IN), .B0(n1887), .Y(n1963));
  OAI21X1 g0930(.A0(P1_D_REG_26__SCAN_IN), .A1(P1_D_REG_25__SCAN_IN), .B0(n1887), .Y(n1964));
  OAI21X1 g0931(.A0(P1_D_REG_31__SCAN_IN), .A1(P1_D_REG_30__SCAN_IN), .B0(n1887), .Y(n1965));
  OAI21X1 g0932(.A0(P1_D_REG_29__SCAN_IN), .A1(P1_D_REG_2__SCAN_IN), .B0(n1887), .Y(n1966));
  NAND4X1 g0933(.A(n1965), .B(n1964), .C(n1963), .D(n1966), .Y(n1967));
  OAI21X1 g0934(.A0(P1_D_REG_21__SCAN_IN), .A1(P1_D_REG_20__SCAN_IN), .B0(n1887), .Y(n1968));
  OAI21X1 g0935(.A0(P1_D_REG_19__SCAN_IN), .A1(P1_D_REG_18__SCAN_IN), .B0(n1887), .Y(n1969));
  OAI21X1 g0936(.A0(P1_D_REG_23__SCAN_IN), .A1(P1_D_REG_22__SCAN_IN), .B0(n1887), .Y(n1970));
  NAND3X1 g0937(.A(n1970), .B(n1969), .C(n1968), .Y(n1971));
  OAI21X1 g0938(.A0(P1_D_REG_14__SCAN_IN), .A1(P1_D_REG_12__SCAN_IN), .B0(n1887), .Y(n1972));
  OAI21X1 g0939(.A0(P1_D_REG_13__SCAN_IN), .A1(P1_D_REG_11__SCAN_IN), .B0(n1887), .Y(n1973));
  OAI21X1 g0940(.A0(P1_D_REG_24__SCAN_IN), .A1(P1_D_REG_16__SCAN_IN), .B0(n1887), .Y(n1974));
  OAI21X1 g0941(.A0(P1_D_REG_17__SCAN_IN), .A1(P1_D_REG_15__SCAN_IN), .B0(n1887), .Y(n1975));
  NAND4X1 g0942(.A(n1974), .B(n1973), .C(n1972), .D(n1975), .Y(n1976));
  NOR4X1  g0943(.A(n1971), .B(n1967), .C(n1962), .D(n1976), .Y(n1977));
  INVX1   g0944(.A(n1977), .Y(n1978));
  AOI21X1 g0945(.A0(n1881), .A1(n1879), .B0(n1887), .Y(n1979));
  AOI21X1 g0946(.A0(n1887), .A1(P1_D_REG_1__SCAN_IN), .B0(n1979), .Y(n1980));
  NOR2X1  g0947(.A(P1_IR_REG_31__SCAN_IN), .B(n1655), .Y(n1981));
  AOI21X1 g0948(.A0(n1658), .A1(P1_IR_REG_31__SCAN_IN), .B0(n1981), .Y(n1982));
  INVX1   g0949(.A(n1982), .Y(n1983));
  NOR2X1  g0950(.A(P1_IR_REG_31__SCAN_IN), .B(n1610), .Y(n1984));
  AOI21X1 g0951(.A0(n1616), .A1(P1_IR_REG_31__SCAN_IN), .B0(n1984), .Y(n1985));
  NOR2X1  g0952(.A(P1_IR_REG_31__SCAN_IN), .B(n1633), .Y(n1986));
  AOI21X1 g0953(.A0(n1634), .A1(P1_IR_REG_31__SCAN_IN), .B0(n1986), .Y(n1987));
  AOI21X1 g0954(.A0(n1987), .A1(n1985), .B0(n1983), .Y(n1988));
  INVX1   g0955(.A(n1987), .Y(n1989));
  NOR2X1  g0956(.A(P1_IR_REG_31__SCAN_IN), .B(n1586), .Y(n1990));
  AOI21X1 g0957(.A0(n1591), .A1(P1_IR_REG_31__SCAN_IN), .B0(n1990), .Y(n1991));
  NAND2X1 g0958(.A(n1991), .B(n1985), .Y(n1992));
  OAI21X1 g0959(.A0(n1989), .A1(n1982), .B0(n1992), .Y(n1993));
  OAI21X1 g0960(.A0(n1993), .A1(n1988), .B0(n1980), .Y(n1994));
  NOR2X1  g0961(.A(n1994), .B(n1978), .Y(n1995));
  AOI21X1 g0962(.A0(n1879), .A1(n1876), .B0(n1887), .Y(n1996));
  AOI21X1 g0963(.A0(n1887), .A1(P1_D_REG_0__SCAN_IN), .B0(n1996), .Y(n1997));
  NAND3X1 g0964(.A(n1997), .B(n1995), .C(n1891), .Y(n1998));
  NOR2X1  g0965(.A(n1803), .B(n1181), .Y(n1999));
  NOR2X1  g0966(.A(P1_IR_REG_31__SCAN_IN), .B(n1791), .Y(n2000));
  NAND2X1 g0967(.A(n1181), .B(P1_IR_REG_27__SCAN_IN), .Y(n2001));
  OAI21X1 g0968(.A0(n1776), .A1(n1181), .B0(n2001), .Y(n2002));
  NOR3X1  g0969(.A(n2002), .B(n2000), .C(n1999), .Y(n2003));
  INVX1   g0970(.A(P1_IR_REG_0__SCAN_IN), .Y(n2004));
  NOR2X1  g0971(.A(n1181), .B(n2004), .Y(n2005));
  NOR2X1  g0972(.A(P1_IR_REG_31__SCAN_IN), .B(n2004), .Y(n2006));
  INVX1   g0973(.A(n2004), .Y(n2008));
  NAND2X1 g0974(.A(n2008), .B(n2003), .Y(n2009));
  OAI21X1 g0975(.A0(n2003), .A1(n1156), .B0(n2009), .Y(n2010));
  INVX1   g0976(.A(n2010), .Y(n2011));
  INVX1   g0977(.A(P1_REG0_REG_0__SCAN_IN), .Y(n2012));
  INVX1   g0978(.A(P1_IR_REG_30__SCAN_IN), .Y(n2013));
  NAND2X1 g0979(.A(n1847), .B(P1_IR_REG_31__SCAN_IN), .Y(n2014));
  OAI21X1 g0980(.A0(P1_IR_REG_31__SCAN_IN), .A1(n2013), .B0(n2014), .Y(n2015));
  NAND2X1 g0981(.A(n1181), .B(P1_IR_REG_29__SCAN_IN), .Y(n2016));
  OAI21X1 g0982(.A0(n1824), .A1(n1181), .B0(n2016), .Y(n2017));
  NOR3X1  g0983(.A(n2017), .B(n2015), .C(n2012), .Y(n2018));
  INVX1   g0984(.A(P1_REG2_REG_0__SCAN_IN), .Y(n2019));
  NOR2X1  g0985(.A(P1_IR_REG_31__SCAN_IN), .B(n2013), .Y(n2020));
  AOI21X1 g0986(.A0(n1847), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2020), .Y(n2021));
  NOR3X1  g0987(.A(n2017), .B(n2021), .C(n2019), .Y(n2022));
  NOR2X1  g0988(.A(n2022), .B(n2018), .Y(n2023));
  NAND3X1 g0989(.A(n2017), .B(n2021), .C(P1_REG1_REG_0__SCAN_IN), .Y(n2024));
  NAND3X1 g0990(.A(n2017), .B(n2015), .C(P1_REG3_REG_0__SCAN_IN), .Y(n2025));
  NAND3X1 g0991(.A(n2025), .B(n2024), .C(n2023), .Y(n2026));
  XOR2X1  g0992(.A(n2026), .B(n2011), .Y(n2027));
  INVX1   g0993(.A(n1985), .Y(n2028));
  NOR3X1  g0994(.A(n1991), .B(n2028), .C(n1982), .Y(n2029));
  INVX1   g0995(.A(n2029), .Y(n2030));
  NOR2X1  g0996(.A(n2030), .B(n2027), .Y(n2031));
  INVX1   g0997(.A(n2031), .Y(n2032));
  NOR3X1  g0998(.A(n1991), .B(n1987), .C(n1985), .Y(n2034));
  NAND2X1 g0999(.A(n1566), .B(P1_IR_REG_19__SCAN_IN), .Y(n2035));
  NAND3X1 g1000(.A(n1608), .B(n2035), .C(P1_IR_REG_31__SCAN_IN), .Y(n2036));
  OAI21X1 g1001(.A0(P1_IR_REG_31__SCAN_IN), .A1(n1586), .B0(n2036), .Y(n2037));
  NOR3X1  g1002(.A(n2037), .B(n1985), .C(n1982), .Y(n2038));
  OAI21X1 g1003(.A0(n2038), .A1(n2034), .B0(n4841), .Y(n2039));
  NOR3X1  g1004(.A(n1991), .B(n1985), .C(n1982), .Y(n2040));
  NOR3X1  g1005(.A(n2037), .B(n1987), .C(n1985), .Y(n2041));
  OAI21X1 g1006(.A0(n2041), .A1(n2040), .B0(n4841), .Y(n2042));
  NOR3X1  g1007(.A(n1992), .B(n1987), .C(n1983), .Y(n2043));
  NAND3X1 g1008(.A(n1991), .B(n1985), .C(n1983), .Y(n2044));
  NOR2X1  g1009(.A(n2044), .B(n1989), .Y(n2045));
  OAI21X1 g1010(.A0(n2045), .A1(n2043), .B0(n4841), .Y(n2046));
  NAND4X1 g1011(.A(n2042), .B(n2039), .C(n2032), .D(n2046), .Y(n2047));
  NOR3X1  g1012(.A(n1991), .B(n2028), .C(n1983), .Y(n2048));
  INVX1   g1013(.A(n2048), .Y(n2049));
  NOR4X1  g1014(.A(n1999), .B(n1987), .C(n1982), .D(n2000), .Y(n2050));
  INVX1   g1015(.A(P1_REG2_REG_1__SCAN_IN), .Y(n2051));
  NOR3X1  g1016(.A(n2017), .B(n2021), .C(n2051), .Y(n2052));
  INVX1   g1017(.A(P1_REG0_REG_1__SCAN_IN), .Y(n2053));
  NOR3X1  g1018(.A(n2017), .B(n2015), .C(n2053), .Y(n2054));
  NOR2X1  g1019(.A(n2054), .B(n2052), .Y(n2055));
  NAND3X1 g1020(.A(n2017), .B(n2021), .C(P1_REG1_REG_1__SCAN_IN), .Y(n2056));
  NAND3X1 g1021(.A(n2017), .B(n2015), .C(P1_REG3_REG_1__SCAN_IN), .Y(n2057));
  NAND3X1 g1022(.A(n2057), .B(n2056), .C(n2055), .Y(n2058));
  NOR2X1  g1023(.A(n2037), .B(n1985), .Y(n2059));
  NOR2X1  g1024(.A(n1991), .B(n1983), .Y(n2060));
  NOR2X1  g1025(.A(n1989), .B(n1983), .Y(n2061));
  AOI22X1 g1026(.A0(n2060), .A1(n1987), .B0(n2059), .B1(n2061), .Y(n2062));
  NOR3X1  g1027(.A(n1989), .B(n2028), .C(n1983), .Y(n2063));
  INVX1   g1028(.A(n2063), .Y(n2064));
  AOI21X1 g1029(.A0(n2064), .A1(n2062), .B0(n2011), .Y(n2065));
  AOI21X1 g1030(.A0(n2058), .A1(n2050), .B0(n2065), .Y(n2066));
  OAI21X1 g1031(.A0(n2049), .A1(n2027), .B0(n2066), .Y(n2067));
  NOR2X1  g1032(.A(n2067), .B(n2047), .Y(n2068));
  NAND2X1 g1033(.A(n1998), .B(P1_REG0_REG_0__SCAN_IN), .Y(n2069));
  OAI21X1 g1034(.A0(n2068), .A1(n1998), .B0(n2069), .Y(P1_U3453));
  NOR2X1  g1035(.A(P1_IR_REG_31__SCAN_IN), .B(n1561), .Y(n2071));
  AOI21X1 g1036(.A0(n1183), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2071), .Y(n2072));
  INVX1   g1037(.A(n2072), .Y(n2073));
  NAND2X1 g1038(.A(n2073), .B(n2003), .Y(n2074));
  OAI21X1 g1039(.A0(n2003), .A1(n1180), .B0(n2074), .Y(n2075));
  XOR2X1  g1040(.A(n2075), .B(n2058), .Y(n2076));
  NAND2X1 g1041(.A(n2026), .B(n2010), .Y(n2077));
  XOR2X1  g1042(.A(n2077), .B(n2076), .Y(n2078));
  INVX1   g1043(.A(n2078), .Y(n2079));
  NOR2X1  g1044(.A(n2000), .B(n1999), .Y(n2080));
  NOR3X1  g1045(.A(n2080), .B(n1987), .C(n1982), .Y(n2081));
  AOI22X1 g1046(.A0(n2079), .A1(n2043), .B0(n2026), .B1(n2081), .Y(n2082));
  OAI21X1 g1047(.A0(n2045), .A1(n2038), .B0(n2079), .Y(n2083));
  NAND4X1 g1048(.A(n2024), .B(n2023), .C(n2010), .D(n2025), .Y(n2084));
  XOR2X1  g1049(.A(n2058), .B(n2084), .Y(n2085));
  XOR2X1  g1050(.A(n2085), .B(n2075), .Y(n2086));
  INVX1   g1051(.A(n2086), .Y(n2087));
  OAI21X1 g1052(.A0(n2041), .A1(n2040), .B0(n2087), .Y(n2088));
  OAI21X1 g1053(.A0(n2034), .A1(n2029), .B0(n2087), .Y(n2089));
  NAND4X1 g1054(.A(n2088), .B(n2083), .C(n2082), .D(n2089), .Y(n2090));
  XOR2X1  g1055(.A(n2075), .B(n2010), .Y(n2091));
  INVX1   g1056(.A(n2050), .Y(n2092));
  INVX1   g1057(.A(n2075), .Y(n2093));
  NOR2X1  g1058(.A(n2017), .B(n2015), .Y(n2094));
  NOR2X1  g1059(.A(n2017), .B(n2021), .Y(n2095));
  AOI22X1 g1060(.A0(n2094), .A1(P1_REG0_REG_2__SCAN_IN), .B0(P1_REG2_REG_2__SCAN_IN), .B1(n2095), .Y(n2096));
  NOR2X1  g1061(.A(n1824), .B(n1181), .Y(n2097));
  AOI21X1 g1062(.A0(n1181), .A1(P1_IR_REG_29__SCAN_IN), .B0(n2097), .Y(n2098));
  NOR2X1  g1063(.A(n2098), .B(n2015), .Y(n2099));
  NOR2X1  g1064(.A(n2098), .B(n2021), .Y(n2100));
  AOI22X1 g1065(.A0(n2099), .A1(P1_REG1_REG_2__SCAN_IN), .B0(P1_REG3_REG_2__SCAN_IN), .B1(n2100), .Y(n2101));
  NAND2X1 g1066(.A(n2101), .B(n2096), .Y(n2102));
  INVX1   g1067(.A(n2102), .Y(n2103));
  OAI22X1 g1068(.A0(n2093), .A1(n2062), .B0(n2092), .B1(n2103), .Y(n2104));
  AOI21X1 g1069(.A0(n2091), .A1(n2063), .B0(n2104), .Y(n2105));
  OAI21X1 g1070(.A0(n2078), .A1(n2049), .B0(n2105), .Y(n2106));
  NOR2X1  g1071(.A(n2106), .B(n2090), .Y(n2107));
  NAND2X1 g1072(.A(n1998), .B(P1_REG0_REG_1__SCAN_IN), .Y(n2108));
  OAI21X1 g1073(.A0(n2107), .A1(n1998), .B0(n2108), .Y(P1_U3456));
  NOR2X1  g1074(.A(P1_IR_REG_31__SCAN_IN), .B(n1197), .Y(n2110));
  AOI21X1 g1075(.A0(n1199), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2110), .Y(n2111));
  INVX1   g1076(.A(n2111), .Y(n2112));
  NAND2X1 g1077(.A(n2112), .B(n2003), .Y(n2113));
  OAI21X1 g1078(.A0(n2003), .A1(n1196), .B0(n2113), .Y(n2114));
  XOR2X1  g1079(.A(n2114), .B(n2102), .Y(n2115));
  NAND2X1 g1080(.A(n2057), .B(n2056), .Y(n2116));
  NOR3X1  g1081(.A(n2116), .B(n2054), .C(n2052), .Y(n2117));
  NOR2X1  g1082(.A(n2093), .B(n2117), .Y(n2118));
  AOI21X1 g1083(.A0(n2093), .A1(n2117), .B0(n2077), .Y(n2119));
  NOR2X1  g1084(.A(n2119), .B(n2118), .Y(n2120));
  INVX1   g1085(.A(n2120), .Y(n2121));
  NOR3X1  g1086(.A(n2115), .B(n2119), .C(n2118), .Y(n2123));
  AOI21X1 g1087(.A0(n2121), .A1(n2115), .B0(n2123), .Y(n2124));
  AOI22X1 g1088(.A0(n2081), .A1(n2058), .B0(n2043), .B1(n2124), .Y(n2125));
  OAI21X1 g1089(.A0(n2045), .A1(n2038), .B0(n2124), .Y(n2126));
  NAND2X1 g1090(.A(n2025), .B(n2024), .Y(n2127));
  NOR3X1  g1091(.A(n2127), .B(n2022), .C(n2018), .Y(n2128));
  AOI21X1 g1092(.A0(n2128), .A1(n2010), .B0(n2117), .Y(n2129));
  NAND3X1 g1093(.A(n2117), .B(n2128), .C(n2010), .Y(n2130));
  AOI21X1 g1094(.A0(n2130), .A1(n2093), .B0(n2129), .Y(n2131));
  XOR2X1  g1095(.A(n2131), .B(n2115), .Y(n2132));
  OAI21X1 g1096(.A0(n2041), .A1(n2040), .B0(n2132), .Y(n2133));
  OAI21X1 g1097(.A0(n2034), .A1(n2029), .B0(n2132), .Y(n2134));
  NAND4X1 g1098(.A(n2133), .B(n2126), .C(n2125), .D(n2134), .Y(n2135));
  NAND2X1 g1099(.A(n2124), .B(n2048), .Y(n2136));
  INVX1   g1100(.A(n2114), .Y(n2137));
  NOR2X1  g1101(.A(n2075), .B(n2010), .Y(n2138));
  XOR2X1  g1102(.A(n2138), .B(n2137), .Y(n2139));
  AOI22X1 g1103(.A0(n2094), .A1(P1_REG0_REG_3__SCAN_IN), .B0(P1_REG2_REG_3__SCAN_IN), .B1(n2095), .Y(n2140));
  INVX1   g1104(.A(n2140), .Y(n2141));
  INVX1   g1105(.A(P1_REG1_REG_3__SCAN_IN), .Y(n2142));
  NAND2X1 g1106(.A(n2017), .B(n2021), .Y(n2143));
  NAND2X1 g1107(.A(n2017), .B(n2015), .Y(n2144));
  OAI22X1 g1108(.A0(n2143), .A1(n2142), .B0(P1_REG3_REG_3__SCAN_IN), .B1(n2144), .Y(n2145));
  NOR2X1  g1109(.A(n2145), .B(n2141), .Y(n2146));
  OAI22X1 g1110(.A0(n2137), .A1(n2062), .B0(n2092), .B1(n2146), .Y(n2147));
  AOI21X1 g1111(.A0(n2139), .A1(n2063), .B0(n2147), .Y(n2148));
  NAND2X1 g1112(.A(n2148), .B(n2136), .Y(n2149));
  NOR2X1  g1113(.A(n2149), .B(n2135), .Y(n2150));
  NAND2X1 g1114(.A(n1998), .B(P1_REG0_REG_2__SCAN_IN), .Y(n2151));
  OAI21X1 g1115(.A0(n2150), .A1(n1998), .B0(n2151), .Y(P1_U3459));
  NAND3X1 g1116(.A(n2137), .B(n2101), .C(n2096), .Y(n2153));
  AOI21X1 g1117(.A0(n2101), .A1(n2096), .B0(n2137), .Y(n2154));
  AOI21X1 g1118(.A0(n2153), .A1(n2118), .B0(n2154), .Y(n2155));
  INVX1   g1119(.A(n2155), .Y(n2156));
  AOI21X1 g1120(.A0(n2119), .A1(n2153), .B0(n2156), .Y(n2157));
  INVX1   g1121(.A(P1_REG3_REG_3__SCAN_IN), .Y(n2158));
  AOI22X1 g1122(.A0(n2099), .A1(P1_REG1_REG_3__SCAN_IN), .B0(n2158), .B1(n2100), .Y(n2159));
  NAND2X1 g1123(.A(n2159), .B(n2140), .Y(n2160));
  NOR2X1  g1124(.A(P1_IR_REG_31__SCAN_IN), .B(n1212), .Y(n2161));
  AOI21X1 g1125(.A0(n1214), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2161), .Y(n2162));
  INVX1   g1126(.A(n2162), .Y(n2163));
  NOR2X1  g1127(.A(n2003), .B(n1211), .Y(n2164));
  AOI21X1 g1128(.A0(n2163), .A1(n2003), .B0(n2164), .Y(n2165));
  XOR2X1  g1129(.A(n2165), .B(n2160), .Y(n2166));
  NAND2X1 g1130(.A(n2163), .B(n2003), .Y(n2168));
  OAI21X1 g1131(.A0(n2003), .A1(n1211), .B0(n2168), .Y(n2169));
  XOR2X1  g1132(.A(n2169), .B(n2160), .Y(n2170));
  NOR2X1  g1133(.A(n2170), .B(n2157), .Y(n2171));
  AOI21X1 g1134(.A0(n2170), .A1(n2157), .B0(n2171), .Y(n2172));
  INVX1   g1135(.A(n2172), .Y(n2173));
  AOI22X1 g1136(.A0(n2102), .A1(n2081), .B0(n2043), .B1(n2173), .Y(n2174));
  OAI21X1 g1137(.A0(n2045), .A1(n2038), .B0(n2173), .Y(n2175));
  INVX1   g1138(.A(n2040), .Y(n2176));
  INVX1   g1139(.A(n2041), .Y(n2177));
  AOI21X1 g1140(.A0(n2101), .A1(n2096), .B0(n2114), .Y(n2178));
  NAND2X1 g1141(.A(n2058), .B(n2084), .Y(n2179));
  OAI21X1 g1142(.A0(n2058), .A1(n2084), .B0(n2093), .Y(n2180));
  NAND2X1 g1143(.A(n2180), .B(n2179), .Y(n2181));
  INVX1   g1144(.A(n2096), .Y(n2182));
  INVX1   g1145(.A(P1_REG1_REG_2__SCAN_IN), .Y(n2183));
  INVX1   g1146(.A(P1_REG3_REG_2__SCAN_IN), .Y(n2184));
  OAI22X1 g1147(.A0(n2143), .A1(n2183), .B0(n2184), .B1(n2144), .Y(n2185));
  NOR3X1  g1148(.A(n2137), .B(n2185), .C(n2182), .Y(n2186));
  NOR2X1  g1149(.A(n2166), .B(n2186), .Y(n2187));
  OAI21X1 g1150(.A0(n2181), .A1(n2178), .B0(n2187), .Y(n2188));
  NOR2X1  g1151(.A(n2170), .B(n2178), .Y(n2189));
  OAI21X1 g1152(.A0(n2131), .A1(n2186), .B0(n2189), .Y(n2190));
  AOI22X1 g1153(.A0(n2188), .A1(n2190), .B0(n2177), .B1(n2176), .Y(n2191));
  INVX1   g1154(.A(n2034), .Y(n2192));
  AOI22X1 g1155(.A0(n2188), .A1(n2190), .B0(n2192), .B1(n2030), .Y(n2193));
  NOR2X1  g1156(.A(n2193), .B(n2191), .Y(n2194));
  NAND3X1 g1157(.A(n2194), .B(n2175), .C(n2174), .Y(n2195));
  NAND2X1 g1158(.A(n2138), .B(n2137), .Y(n2196));
  XOR2X1  g1159(.A(n2169), .B(n2196), .Y(n2197));
  AOI22X1 g1160(.A0(n2094), .A1(P1_REG0_REG_4__SCAN_IN), .B0(P1_REG2_REG_4__SCAN_IN), .B1(n2095), .Y(n2198));
  INVX1   g1161(.A(n2198), .Y(n2199));
  INVX1   g1162(.A(P1_REG1_REG_4__SCAN_IN), .Y(n2200));
  INVX1   g1163(.A(P1_REG3_REG_4__SCAN_IN), .Y(n2201));
  XOR2X1  g1164(.A(P1_REG3_REG_3__SCAN_IN), .B(n2201), .Y(n2202));
  OAI22X1 g1165(.A0(n2144), .A1(n2202), .B0(n2143), .B1(n2200), .Y(n2203));
  NOR2X1  g1166(.A(n2203), .B(n2199), .Y(n2204));
  OAI22X1 g1167(.A0(n2165), .A1(n2062), .B0(n2092), .B1(n2204), .Y(n2205));
  AOI21X1 g1168(.A0(n2197), .A1(n2063), .B0(n2205), .Y(n2206));
  OAI21X1 g1169(.A0(n2172), .A1(n2049), .B0(n2206), .Y(n2207));
  NOR2X1  g1170(.A(n2207), .B(n2195), .Y(n2208));
  NAND2X1 g1171(.A(n1998), .B(P1_REG0_REG_3__SCAN_IN), .Y(n2209));
  OAI21X1 g1172(.A0(n2208), .A1(n1998), .B0(n2209), .Y(P1_U3462));
  INVX1   g1173(.A(n2043), .Y(n2211));
  INVX1   g1174(.A(n2081), .Y(n2212));
  NAND2X1 g1175(.A(n2165), .B(n2146), .Y(n2213));
  NOR2X1  g1176(.A(n2165), .B(n2146), .Y(n2215));
  INVX1   g1177(.A(n2203), .Y(n2218));
  NAND2X1 g1178(.A(n2218), .B(n2198), .Y(n2219));
  NOR2X1  g1179(.A(P1_IR_REG_31__SCAN_IN), .B(n1276), .Y(n2220));
  AOI21X1 g1180(.A0(n1239), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2220), .Y(n2221));
  INVX1   g1181(.A(n2221), .Y(n2222));
  NAND2X1 g1182(.A(n2222), .B(n2003), .Y(n2223));
  OAI21X1 g1183(.A0(n2003), .A1(n1235), .B0(n2223), .Y(n2224));
  INVX1   g1184(.A(n2224), .Y(n2225));
  XOR2X1  g1185(.A(n2225), .B(n2219), .Y(n2226));
  NOR2X1  g1186(.A(n2337), .B(n2226), .Y(n2227));
  AOI21X1 g1187(.A0(n2226), .A1(n2337), .B0(n2227), .Y(n2229));
  OAI22X1 g1188(.A0(n2146), .A1(n2212), .B0(n2211), .B1(n2229), .Y(n2230));
  INVX1   g1189(.A(n2038), .Y(n2231));
  INVX1   g1190(.A(n2045), .Y(n2232));
  AOI21X1 g1191(.A0(n2232), .A1(n2231), .B0(n2229), .Y(n2233));
  NAND3X1 g1192(.A(n2169), .B(n2159), .C(n2140), .Y(n2234));
  AOI21X1 g1193(.A0(n2180), .A1(n2179), .B0(n2186), .Y(n2235));
  OAI21X1 g1194(.A0(n2160), .A1(n2178), .B0(n2165), .Y(n2236));
  NAND2X1 g1195(.A(n2160), .B(n2178), .Y(n2237));
  NAND2X1 g1196(.A(n2237), .B(n2236), .Y(n2238));
  AOI21X1 g1197(.A0(n2235), .A1(n2234), .B0(n2238), .Y(n2239));
  XOR2X1  g1198(.A(n2239), .B(n2226), .Y(n2240));
  INVX1   g1199(.A(n2240), .Y(n2241));
  OAI21X1 g1200(.A0(n2041), .A1(n2040), .B0(n2241), .Y(n2242));
  OAI21X1 g1201(.A0(n2034), .A1(n2029), .B0(n2241), .Y(n2243));
  NAND2X1 g1202(.A(n2243), .B(n2242), .Y(n2244));
  NOR4X1  g1203(.A(n2114), .B(n2075), .C(n2010), .D(n2169), .Y(n2245));
  XOR2X1  g1204(.A(n2225), .B(n2245), .Y(n2246));
  INVX1   g1205(.A(P1_REG2_REG_5__SCAN_IN), .Y(n2247));
  NAND2X1 g1206(.A(n2098), .B(n2015), .Y(n2248));
  NAND2X1 g1207(.A(n2094), .B(P1_REG0_REG_5__SCAN_IN), .Y(n2249));
  OAI21X1 g1208(.A0(n2248), .A1(n2247), .B0(n2249), .Y(n2250));
  NAND3X1 g1209(.A(n2017), .B(n2021), .C(P1_REG1_REG_5__SCAN_IN), .Y(n2251));
  NAND2X1 g1210(.A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), .Y(n2252));
  XOR2X1  g1211(.A(n2252), .B(P1_REG3_REG_5__SCAN_IN), .Y(n2253));
  INVX1   g1212(.A(n2253), .Y(n2254));
  NAND3X1 g1213(.A(n2254), .B(n2017), .C(n2015), .Y(n2255));
  NAND2X1 g1214(.A(n2255), .B(n2251), .Y(n2256));
  NOR2X1  g1215(.A(n2256), .B(n2250), .Y(n2257));
  OAI22X1 g1216(.A0(n2225), .A1(n2062), .B0(n2092), .B1(n2257), .Y(n2258));
  AOI21X1 g1217(.A0(n2246), .A1(n2063), .B0(n2258), .Y(n2259));
  OAI21X1 g1218(.A0(n2229), .A1(n2049), .B0(n2259), .Y(n2260));
  NOR4X1  g1219(.A(n2244), .B(n2233), .C(n2230), .D(n2260), .Y(n2261));
  NAND2X1 g1220(.A(n1998), .B(P1_REG0_REG_4__SCAN_IN), .Y(n2262));
  OAI21X1 g1221(.A0(n2261), .A1(n1998), .B0(n2262), .Y(P1_U3465));
  NOR2X1  g1222(.A(P1_IR_REG_31__SCAN_IN), .B(n1257), .Y(n2264));
  AOI21X1 g1223(.A0(n1258), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2264), .Y(n2265));
  INVX1   g1224(.A(n2265), .Y(n2266));
  NAND2X1 g1225(.A(n2266), .B(n2003), .Y(n2267));
  OAI21X1 g1226(.A0(n2003), .A1(n1256), .B0(n2267), .Y(n2268));
  XOR2X1  g1227(.A(n2268), .B(n2257), .Y(n2269));
  NOR2X1  g1228(.A(n2225), .B(n2219), .Y(n2270));
  INVX1   g1229(.A(n2270), .Y(n2271));
  AOI21X1 g1230(.A0(n2218), .A1(n2198), .B0(n2224), .Y(n2272));
  NAND2X1 g1231(.A(n2235), .B(n2234), .Y(n2273));
  NAND3X1 g1232(.A(n2237), .B(n2236), .C(n2273), .Y(n2274));
  AOI21X1 g1233(.A0(n2274), .A1(n2271), .B0(n2272), .Y(n2275));
  XOR2X1  g1234(.A(n2275), .B(n2269), .Y(n2276));
  INVX1   g1235(.A(n2276), .Y(n2277));
  NAND2X1 g1236(.A(n2277), .B(n2041), .Y(n2278));
  NOR2X1  g1237(.A(n2225), .B(n2204), .Y(n2279));
  NOR2X1  g1238(.A(n2279), .B(n2337), .Y(n2280));
  INVX1   g1239(.A(n2280), .Y(n2281));
  INVX1   g1240(.A(n2268), .Y(n2283));
  AOI22X1 g1241(.A0(n2257), .A1(n2283), .B0(n2225), .B1(n2204), .Y(n2284));
  INVX1   g1242(.A(n2284), .Y(n2285));
  AOI21X1 g1243(.A0(n2268), .A1(n4594), .B0(n2285), .Y(n2286));
  OAI21X1 g1244(.A0(n2224), .A1(n2219), .B0(n2337), .Y(n2287));
  NAND2X1 g1245(.A(n2268), .B(n2257), .Y(n2288));
  INVX1   g1246(.A(n2288), .Y(n2289));
  NOR2X1  g1247(.A(n2268), .B(n2257), .Y(n2290));
  NOR3X1  g1248(.A(n2290), .B(n2289), .C(n2279), .Y(n2291));
  AOI22X1 g1249(.A0(n2287), .A1(n2291), .B0(n2286), .B1(n2281), .Y(n2292));
  AOI22X1 g1250(.A0(n2219), .A1(n2081), .B0(n2043), .B1(n2292), .Y(n2293));
  OAI21X1 g1251(.A0(n2045), .A1(n2038), .B0(n2292), .Y(n2294));
  NAND3X1 g1252(.A(n2294), .B(n2293), .C(n2278), .Y(n2295));
  OAI21X1 g1253(.A0(n2040), .A1(n2029), .B0(n2277), .Y(n2296));
  OAI21X1 g1254(.A0(n2276), .A1(n2192), .B0(n2296), .Y(n2297));
  INVX1   g1255(.A(n2292), .Y(n2298));
  NOR2X1  g1256(.A(n2298), .B(n2049), .Y(n2299));
  NOR3X1  g1257(.A(n2224), .B(n2169), .C(n2196), .Y(n2300));
  XOR2X1  g1258(.A(n2268), .B(n2300), .Y(n2301));
  INVX1   g1259(.A(n2062), .Y(n2302));
  INVX1   g1260(.A(P1_REG2_REG_6__SCAN_IN), .Y(n2303));
  NAND2X1 g1261(.A(n2094), .B(P1_REG0_REG_6__SCAN_IN), .Y(n2304));
  OAI21X1 g1262(.A0(n2248), .A1(n2303), .B0(n2304), .Y(n2305));
  NAND3X1 g1263(.A(n2017), .B(n2021), .C(P1_REG1_REG_6__SCAN_IN), .Y(n2306));
  NAND3X1 g1264(.A(P1_REG3_REG_3__SCAN_IN), .B(P1_REG3_REG_5__SCAN_IN), .C(P1_REG3_REG_4__SCAN_IN), .Y(n2307));
  XOR2X1  g1265(.A(n2307), .B(P1_REG3_REG_6__SCAN_IN), .Y(n2308));
  INVX1   g1266(.A(n2308), .Y(n2309));
  NAND3X1 g1267(.A(n2309), .B(n2017), .C(n2015), .Y(n2310));
  NAND2X1 g1268(.A(n2310), .B(n2306), .Y(n2311));
  NOR2X1  g1269(.A(n2311), .B(n2305), .Y(n2312));
  INVX1   g1270(.A(n2312), .Y(n2313));
  AOI22X1 g1271(.A0(n2268), .A1(n2302), .B0(n2050), .B1(n2313), .Y(n2314));
  OAI21X1 g1272(.A0(n2301), .A1(n2064), .B0(n2314), .Y(n2315));
  NOR4X1  g1273(.A(n2299), .B(n2297), .C(n2295), .D(n2315), .Y(n2316));
  NAND2X1 g1274(.A(n1998), .B(P1_REG0_REG_5__SCAN_IN), .Y(n2317));
  OAI21X1 g1275(.A0(n2316), .A1(n1998), .B0(n2317), .Y(P1_U3468));
  INVX1   g1276(.A(n2275), .Y(n2319));
  NOR2X1  g1277(.A(P1_IR_REG_31__SCAN_IN), .B(n1278), .Y(n2320));
  AOI21X1 g1278(.A0(n1281), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2320), .Y(n2321));
  INVX1   g1279(.A(n2321), .Y(n2322));
  NAND2X1 g1280(.A(n2322), .B(n2003), .Y(n2323));
  OAI21X1 g1281(.A0(n2003), .A1(n1275), .B0(n2323), .Y(n2324));
  XOR2X1  g1282(.A(n2324), .B(n2312), .Y(n2325));
  AOI21X1 g1283(.A0(n2268), .A1(n2257), .B0(n2325), .Y(n2326));
  OAI21X1 g1284(.A0(n2319), .A1(n2290), .B0(n2326), .Y(n2327));
  NAND2X1 g1285(.A(n2324), .B(n2312), .Y(n2328));
  INVX1   g1286(.A(n2328), .Y(n2329));
  NOR2X1  g1287(.A(n2324), .B(n2312), .Y(n2330));
  NOR3X1  g1288(.A(n2330), .B(n2329), .C(n2290), .Y(n2331));
  OAI21X1 g1289(.A0(n2275), .A1(n2289), .B0(n2331), .Y(n2332));
  AOI21X1 g1290(.A0(n2332), .A1(n2327), .B0(n2177), .Y(n2333));
  INVX1   g1291(.A(n2333), .Y(n2334));
  OAI21X1 g1292(.A0(n2169), .A1(n2160), .B0(n2153), .Y(n2335));
  AOI21X1 g1293(.A0(n2213), .A1(n2154), .B0(n2215), .Y(n2336));
  OAI21X1 g1294(.A0(n2335), .A1(n2120), .B0(n2336), .Y(n2337));
  NAND3X1 g1295(.A(n2268), .B(n2224), .C(n2219), .Y(n2338));
  AOI21X1 g1296(.A0(n2224), .A1(n2219), .B0(n2268), .Y(n2339));
  OAI21X1 g1297(.A0(n2339), .A1(n2257), .B0(n2338), .Y(n2340));
  AOI21X1 g1298(.A0(n2337), .A1(n2284), .B0(n2340), .Y(n2341));
  INVX1   g1299(.A(n2341), .Y(n2342));
  NOR2X1  g1300(.A(n2342), .B(n2325), .Y(n2343));
  AOI21X1 g1301(.A0(n2325), .A1(n2342), .B0(n2343), .Y(n2345));
  INVX1   g1302(.A(n2345), .Y(n2346));
  AOI22X1 g1303(.A0(n4594), .A1(n2081), .B0(n2043), .B1(n2346), .Y(n2347));
  OAI21X1 g1304(.A0(n2045), .A1(n2038), .B0(n2346), .Y(n2348));
  AOI21X1 g1305(.A0(n2332), .A1(n2327), .B0(n2192), .Y(n2349));
  AOI21X1 g1306(.A0(n2332), .A1(n2327), .B0(n2176), .Y(n2350));
  AOI21X1 g1307(.A0(n2332), .A1(n2327), .B0(n2030), .Y(n2351));
  NOR3X1  g1308(.A(n2351), .B(n2350), .C(n2349), .Y(n2352));
  NAND4X1 g1309(.A(n2348), .B(n2347), .C(n2334), .D(n2352), .Y(n2353));
  NOR4X1  g1310(.A(n2224), .B(n2169), .C(n2196), .D(n2268), .Y(n2354));
  INVX1   g1311(.A(n2324), .Y(n2355));
  XOR2X1  g1312(.A(n2355), .B(n2354), .Y(n2356));
  AOI22X1 g1313(.A0(n2094), .A1(P1_REG0_REG_7__SCAN_IN), .B0(P1_REG2_REG_7__SCAN_IN), .B1(n2095), .Y(n2357));
  NAND4X1 g1314(.A(P1_REG3_REG_5__SCAN_IN), .B(P1_REG3_REG_4__SCAN_IN), .C(P1_REG3_REG_6__SCAN_IN), .D(P1_REG3_REG_3__SCAN_IN), .Y(n2358));
  XOR2X1  g1315(.A(n2358), .B(P1_REG3_REG_7__SCAN_IN), .Y(n2359));
  INVX1   g1316(.A(n2359), .Y(n2360));
  AOI22X1 g1317(.A0(n2100), .A1(n2360), .B0(n2099), .B1(P1_REG1_REG_7__SCAN_IN), .Y(n2361));
  NAND2X1 g1318(.A(n2361), .B(n2357), .Y(n2362));
  INVX1   g1319(.A(n2362), .Y(n2363));
  OAI22X1 g1320(.A0(n2355), .A1(n2062), .B0(n2092), .B1(n2363), .Y(n2364));
  AOI21X1 g1321(.A0(n2356), .A1(n2063), .B0(n2364), .Y(n2365));
  OAI21X1 g1322(.A0(n2345), .A1(n2049), .B0(n2365), .Y(n2366));
  NOR2X1  g1323(.A(n2366), .B(n2353), .Y(n2367));
  NAND2X1 g1324(.A(n1998), .B(P1_REG0_REG_6__SCAN_IN), .Y(n2368));
  OAI21X1 g1325(.A0(n2367), .A1(n1998), .B0(n2368), .Y(P1_U3471));
  OAI21X1 g1326(.A0(n2311), .A1(n2305), .B0(n2324), .Y(n2370));
  INVX1   g1327(.A(n2370), .Y(n2371));
  NOR2X1  g1328(.A(P1_IR_REG_31__SCAN_IN), .B(n1316), .Y(n2372));
  AOI21X1 g1329(.A0(n1317), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2372), .Y(n2373));
  INVX1   g1330(.A(n2373), .Y(n2374));
  NAND2X1 g1331(.A(n2374), .B(n2003), .Y(n2375));
  OAI21X1 g1332(.A0(n2003), .A1(n1315), .B0(n2375), .Y(n2376));
  OAI22X1 g1333(.A0(n2362), .A1(n2376), .B0(n2324), .B1(n2313), .Y(n2377));
  AOI21X1 g1334(.A0(n2376), .A1(n2362), .B0(n2377), .Y(n2378));
  OAI21X1 g1335(.A0(n2371), .A1(n2342), .B0(n2378), .Y(n2379));
  AOI21X1 g1336(.A0(n2355), .A1(n2312), .B0(n2341), .Y(n2380));
  XOR2X1  g1337(.A(n2376), .B(n2363), .Y(n2381));
  NAND2X1 g1338(.A(n2381), .B(n2370), .Y(n2382));
  OAI21X1 g1339(.A0(n2382), .A1(n2380), .B0(n2379), .Y(n2383));
  AOI21X1 g1340(.A0(n2232), .A1(n2231), .B0(n2383), .Y(n2384));
  NOR2X1  g1341(.A(n2330), .B(n2290), .Y(n2385));
  NAND2X1 g1342(.A(n2288), .B(n2272), .Y(n2386));
  AOI21X1 g1343(.A0(n2386), .A1(n2385), .B0(n2329), .Y(n2387));
  NAND3X1 g1344(.A(n2328), .B(n2288), .C(n2271), .Y(n2388));
  NOR2X1  g1345(.A(n2388), .B(n2239), .Y(n2389));
  NOR2X1  g1346(.A(n2389), .B(n2387), .Y(n2390));
  XOR2X1  g1347(.A(n2390), .B(n2381), .Y(n2391));
  OAI22X1 g1348(.A0(n2383), .A1(n2211), .B0(n2192), .B1(n2391), .Y(n2392));
  INVX1   g1349(.A(n2391), .Y(n2393));
  AOI22X1 g1350(.A0(n2313), .A1(n2081), .B0(n2041), .B1(n2393), .Y(n2394));
  OAI21X1 g1351(.A0(n2040), .A1(n2029), .B0(n2393), .Y(n2395));
  NAND2X1 g1352(.A(n2395), .B(n2394), .Y(n2396));
  NAND3X1 g1353(.A(n2355), .B(n2283), .C(n2300), .Y(n2397));
  XOR2X1  g1354(.A(n2376), .B(n2397), .Y(n2398));
  INVX1   g1355(.A(n2376), .Y(n2399));
  AOI22X1 g1356(.A0(n2094), .A1(P1_REG0_REG_8__SCAN_IN), .B0(P1_REG2_REG_8__SCAN_IN), .B1(n2095), .Y(n2400));
  NAND3X1 g1357(.A(n2017), .B(n2021), .C(P1_REG1_REG_8__SCAN_IN), .Y(n2401));
  INVX1   g1358(.A(P1_REG3_REG_8__SCAN_IN), .Y(n2402));
  INVX1   g1359(.A(P1_REG3_REG_7__SCAN_IN), .Y(n2403));
  NOR2X1  g1360(.A(n2358), .B(n2403), .Y(n2404));
  XOR2X1  g1361(.A(n2404), .B(n2402), .Y(n2405));
  INVX1   g1362(.A(n2405), .Y(n2406));
  NAND3X1 g1363(.A(n2406), .B(n2017), .C(n2015), .Y(n2407));
  NAND3X1 g1364(.A(n2407), .B(n2401), .C(n2400), .Y(n2408));
  INVX1   g1365(.A(n2408), .Y(n2409));
  OAI22X1 g1366(.A0(n2399), .A1(n2062), .B0(n2092), .B1(n2409), .Y(n2410));
  AOI21X1 g1367(.A0(n2398), .A1(n2063), .B0(n2410), .Y(n2411));
  OAI21X1 g1368(.A0(n2383), .A1(n2049), .B0(n2411), .Y(n2412));
  NOR4X1  g1369(.A(n2396), .B(n2392), .C(n2384), .D(n2412), .Y(n2413));
  NAND2X1 g1370(.A(n1998), .B(P1_REG0_REG_7__SCAN_IN), .Y(n2414));
  OAI21X1 g1371(.A0(n2413), .A1(n1998), .B0(n2414), .Y(P1_U3474));
  AOI21X1 g1372(.A0(n2399), .A1(n2370), .B0(n2363), .Y(n2416));
  AOI21X1 g1373(.A0(n2376), .A1(n2371), .B0(n2416), .Y(n2417));
  OAI21X1 g1374(.A0(n2377), .A1(n2341), .B0(n2417), .Y(n2418));
  INVX1   g1375(.A(n2418), .Y(n2419));
  NOR2X1  g1376(.A(P1_IR_REG_31__SCAN_IN), .B(n1337), .Y(n2420));
  AOI21X1 g1377(.A0(n1342), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2420), .Y(n2421));
  INVX1   g1378(.A(n2421), .Y(n2422));
  NAND2X1 g1379(.A(n2422), .B(n2003), .Y(n2423));
  OAI21X1 g1380(.A0(n2003), .A1(n1336), .B0(n2423), .Y(n2424));
  XOR2X1  g1381(.A(n2424), .B(n2409), .Y(n2425));
  XOR2X1  g1382(.A(n2424), .B(n2408), .Y(n2427));
  NOR2X1  g1383(.A(n2427), .B(n2419), .Y(n2428));
  AOI21X1 g1384(.A0(n2427), .A1(n2419), .B0(n2428), .Y(n2429));
  AOI21X1 g1385(.A0(n2232), .A1(n2231), .B0(n2429), .Y(n2430));
  NOR2X1  g1386(.A(n2399), .B(n2362), .Y(n2431));
  AOI21X1 g1387(.A0(n2361), .A1(n2357), .B0(n2376), .Y(n2432));
  NOR3X1  g1388(.A(n2389), .B(n2387), .C(n2432), .Y(n2433));
  NOR3X1  g1389(.A(n2433), .B(n2425), .C(n2431), .Y(n2434));
  NAND2X1 g1390(.A(n2386), .B(n2385), .Y(n2435));
  NAND2X1 g1391(.A(n2435), .B(n2328), .Y(n2436));
  NAND4X1 g1392(.A(n2288), .B(n2274), .C(n2271), .D(n2328), .Y(n2437));
  AOI21X1 g1393(.A0(n2437), .A1(n2436), .B0(n2431), .Y(n2438));
  NOR3X1  g1394(.A(n2438), .B(n2427), .C(n2432), .Y(n2439));
  NOR2X1  g1395(.A(n2439), .B(n2434), .Y(n2440));
  OAI22X1 g1396(.A0(n2429), .A1(n2211), .B0(n2192), .B1(n2440), .Y(n2441));
  OAI21X1 g1397(.A0(n2439), .A1(n2434), .B0(n2041), .Y(n2442));
  NAND2X1 g1398(.A(n2362), .B(n2081), .Y(n2443));
  OAI22X1 g1399(.A0(n2434), .A1(n2439), .B0(n2040), .B1(n2029), .Y(n2444));
  NAND3X1 g1400(.A(n2444), .B(n2443), .C(n2442), .Y(n2445));
  NOR2X1  g1401(.A(n2376), .B(n2397), .Y(n2446));
  INVX1   g1402(.A(n2424), .Y(n2447));
  XOR2X1  g1403(.A(n2447), .B(n2446), .Y(n2448));
  INVX1   g1404(.A(P1_REG3_REG_9__SCAN_IN), .Y(n2449));
  NOR3X1  g1405(.A(n2358), .B(n2403), .C(n2402), .Y(n2450));
  XOR2X1  g1406(.A(n2450), .B(n2449), .Y(n2451));
  NOR2X1  g1407(.A(n2451), .B(n2144), .Y(n2452));
  INVX1   g1408(.A(P1_REG0_REG_9__SCAN_IN), .Y(n2453));
  NOR3X1  g1409(.A(n2017), .B(n2015), .C(n2453), .Y(n2454));
  NOR2X1  g1410(.A(n2454), .B(n2452), .Y(n2455));
  AOI22X1 g1411(.A0(n2095), .A1(P1_REG2_REG_9__SCAN_IN), .B0(P1_REG1_REG_9__SCAN_IN), .B1(n2099), .Y(n2456));
  NAND2X1 g1412(.A(n2456), .B(n2455), .Y(n2457));
  INVX1   g1413(.A(n2457), .Y(n2458));
  OAI22X1 g1414(.A0(n2447), .A1(n2062), .B0(n2092), .B1(n2458), .Y(n2459));
  AOI21X1 g1415(.A0(n2448), .A1(n2063), .B0(n2459), .Y(n2460));
  OAI21X1 g1416(.A0(n2429), .A1(n2049), .B0(n2460), .Y(n2461));
  NOR4X1  g1417(.A(n2445), .B(n2441), .C(n2430), .D(n2461), .Y(n2462));
  NAND2X1 g1418(.A(n1998), .B(P1_REG0_REG_8__SCAN_IN), .Y(n2463));
  OAI21X1 g1419(.A0(n2462), .A1(n1998), .B0(n2463), .Y(P1_U3477));
  NOR2X1  g1420(.A(P1_IR_REG_31__SCAN_IN), .B(n1361), .Y(n2465));
  AOI21X1 g1421(.A0(n1362), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2465), .Y(n2466));
  INVX1   g1422(.A(n2466), .Y(n2467));
  NAND2X1 g1423(.A(n2467), .B(n2003), .Y(n2468));
  OAI21X1 g1424(.A0(n2003), .A1(n1360), .B0(n2468), .Y(n2469));
  XOR2X1  g1425(.A(n2469), .B(n2458), .Y(n2470));
  AOI22X1 g1426(.A0(n2409), .A1(n2424), .B0(n2376), .B1(n2363), .Y(n2471));
  INVX1   g1427(.A(n2471), .Y(n2472));
  AOI21X1 g1428(.A0(n2437), .A1(n2436), .B0(n2472), .Y(n2473));
  INVX1   g1429(.A(n2432), .Y(n2474));
  OAI21X1 g1430(.A0(n2408), .A1(n2432), .B0(n2447), .Y(n2475));
  OAI21X1 g1431(.A0(n2409), .A1(n2474), .B0(n2475), .Y(n2476));
  NOR2X1  g1432(.A(n2476), .B(n2473), .Y(n2477));
  XOR2X1  g1433(.A(n2477), .B(n2470), .Y(n2478));
  INVX1   g1434(.A(n2478), .Y(n2479));
  OAI21X1 g1435(.A0(n2040), .A1(n2029), .B0(n2479), .Y(n2480));
  OAI21X1 g1436(.A0(n2478), .A1(n2192), .B0(n2480), .Y(n2481));
  NOR2X1  g1437(.A(n2424), .B(n2408), .Y(n2482));
  NAND2X1 g1438(.A(n2424), .B(n2408), .Y(n2483));
  OAI21X1 g1439(.A0(n2482), .A1(n2419), .B0(n2483), .Y(n2484));
  NOR2X1  g1440(.A(n2484), .B(n2470), .Y(n2485));
  XOR2X1  g1441(.A(n2469), .B(n2457), .Y(n2486));
  AOI21X1 g1442(.A0(n2470), .A1(n2484), .B0(n2485), .Y(n2488));
  AOI22X1 g1443(.A0(n2408), .A1(n2081), .B0(n2041), .B1(n2479), .Y(n2489));
  OAI21X1 g1444(.A0(n2488), .A1(n2231), .B0(n2489), .Y(n2490));
  INVX1   g1445(.A(n2488), .Y(n2491));
  OAI21X1 g1446(.A0(n2045), .A1(n2043), .B0(n2491), .Y(n2492));
  INVX1   g1447(.A(n2492), .Y(n2493));
  NAND4X1 g1448(.A(n2399), .B(n2355), .C(n2354), .D(n2447), .Y(n2494));
  XOR2X1  g1449(.A(n2469), .B(n2494), .Y(n2495));
  INVX1   g1450(.A(n2469), .Y(n2496));
  INVX1   g1451(.A(P1_REG3_REG_10__SCAN_IN), .Y(n2497));
  NOR4X1  g1452(.A(n2403), .B(n2402), .C(n2449), .D(n2358), .Y(n2498));
  XOR2X1  g1453(.A(n2498), .B(n2497), .Y(n2499));
  INVX1   g1454(.A(n2499), .Y(n2500));
  AOI22X1 g1455(.A0(n2100), .A1(n2500), .B0(n2094), .B1(P1_REG0_REG_10__SCAN_IN), .Y(n2501));
  AOI22X1 g1456(.A0(n2095), .A1(P1_REG2_REG_10__SCAN_IN), .B0(P1_REG1_REG_10__SCAN_IN), .B1(n2099), .Y(n2502));
  NAND2X1 g1457(.A(n2502), .B(n2501), .Y(n2503));
  INVX1   g1458(.A(n2503), .Y(n2504));
  OAI22X1 g1459(.A0(n2496), .A1(n2062), .B0(n2092), .B1(n2504), .Y(n2505));
  AOI21X1 g1460(.A0(n2495), .A1(n2063), .B0(n2505), .Y(n2506));
  OAI21X1 g1461(.A0(n2488), .A1(n2049), .B0(n2506), .Y(n2507));
  NOR4X1  g1462(.A(n2493), .B(n2490), .C(n2481), .D(n2507), .Y(n2508));
  NAND2X1 g1463(.A(n1998), .B(P1_REG0_REG_9__SCAN_IN), .Y(n2509));
  OAI21X1 g1464(.A0(n2508), .A1(n1998), .B0(n2509), .Y(P1_U3480));
  AOI21X1 g1465(.A0(n2469), .A1(n2457), .B0(n2484), .Y(n2511));
  NOR2X1  g1466(.A(P1_IR_REG_31__SCAN_IN), .B(n1381), .Y(n2512));
  AOI21X1 g1467(.A0(n1384), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2512), .Y(n2513));
  INVX1   g1468(.A(n2513), .Y(n2514));
  NAND2X1 g1469(.A(n2514), .B(n2003), .Y(n2515));
  OAI21X1 g1470(.A0(n2003), .A1(n1380), .B0(n2515), .Y(n2516));
  INVX1   g1471(.A(n2516), .Y(n2517));
  NOR2X1  g1472(.A(n2517), .B(n2504), .Y(n2518));
  OAI22X1 g1473(.A0(n2503), .A1(n2516), .B0(n2469), .B1(n2457), .Y(n2519));
  NOR3X1  g1474(.A(n2519), .B(n2518), .C(n2511), .Y(n2520));
  OAI21X1 g1475(.A0(n2469), .A1(n2457), .B0(n2484), .Y(n2521));
  XOR2X1  g1476(.A(n2516), .B(n2504), .Y(n2522));
  AOI21X1 g1477(.A0(n2469), .A1(n2457), .B0(n4840), .Y(n2524));
  AOI21X1 g1478(.A0(n2524), .A1(n2521), .B0(n2520), .Y(n2525));
  INVX1   g1479(.A(n2525), .Y(n2526));
  AOI21X1 g1480(.A0(n2232), .A1(n2231), .B0(n2526), .Y(n2527));
  NAND2X1 g1481(.A(n2469), .B(n2458), .Y(n2528));
  NOR2X1  g1482(.A(n2469), .B(n2458), .Y(n2529));
  INVX1   g1483(.A(n2477), .Y(n2530));
  AOI21X1 g1484(.A0(n2530), .A1(n2528), .B0(n2529), .Y(n2531));
  XOR2X1  g1485(.A(n2531), .B(n2522), .Y(n2532));
  OAI22X1 g1486(.A0(n2526), .A1(n2211), .B0(n2192), .B1(n2532), .Y(n2533));
  INVX1   g1487(.A(n2532), .Y(n2534));
  AOI22X1 g1488(.A0(n2457), .A1(n2081), .B0(n2041), .B1(n2534), .Y(n2535));
  OAI21X1 g1489(.A0(n2040), .A1(n2029), .B0(n2534), .Y(n2536));
  NAND2X1 g1490(.A(n2536), .B(n2535), .Y(n2537));
  NOR4X1  g1491(.A(n2424), .B(n2376), .C(n2397), .D(n2469), .Y(n2538));
  NOR2X1  g1492(.A(n2517), .B(n2538), .Y(n2539));
  NOR3X1  g1493(.A(n2516), .B(n2469), .C(n2494), .Y(n2540));
  NOR2X1  g1494(.A(n2540), .B(n2539), .Y(n2541));
  NAND2X1 g1495(.A(n2498), .B(P1_REG3_REG_10__SCAN_IN), .Y(n2542));
  XOR2X1  g1496(.A(n2542), .B(P1_REG3_REG_11__SCAN_IN), .Y(n2543));
  NOR2X1  g1497(.A(n2543), .B(n2144), .Y(n2544));
  INVX1   g1498(.A(P1_REG0_REG_11__SCAN_IN), .Y(n2545));
  NOR3X1  g1499(.A(n2017), .B(n2015), .C(n2545), .Y(n2546));
  AOI22X1 g1500(.A0(n2095), .A1(P1_REG2_REG_11__SCAN_IN), .B0(P1_REG1_REG_11__SCAN_IN), .B1(n2099), .Y(n2547));
  INVX1   g1501(.A(n2547), .Y(n2548));
  NOR3X1  g1502(.A(n2548), .B(n2546), .C(n2544), .Y(n2549));
  OAI22X1 g1503(.A0(n2517), .A1(n2062), .B0(n2092), .B1(n2549), .Y(n2550));
  AOI21X1 g1504(.A0(n2541), .A1(n2063), .B0(n2550), .Y(n2551));
  OAI21X1 g1505(.A0(n2526), .A1(n2049), .B0(n2551), .Y(n2552));
  NOR4X1  g1506(.A(n2537), .B(n2533), .C(n2527), .D(n2552), .Y(n2553));
  NAND2X1 g1507(.A(n1998), .B(P1_REG0_REG_10__SCAN_IN), .Y(n2554));
  OAI21X1 g1508(.A0(n2553), .A1(n1998), .B0(n2554), .Y(P1_U3483));
  NOR2X1  g1509(.A(n2516), .B(n2504), .Y(n2556));
  INVX1   g1510(.A(n2531), .Y(n2557));
  NOR2X1  g1511(.A(P1_IR_REG_31__SCAN_IN), .B(n1404), .Y(n2558));
  AOI21X1 g1512(.A0(n1408), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2558), .Y(n2559));
  INVX1   g1513(.A(n2559), .Y(n2560));
  NAND2X1 g1514(.A(n2560), .B(n2003), .Y(n2561));
  OAI21X1 g1515(.A0(n2003), .A1(n1403), .B0(n2561), .Y(n2562));
  XOR2X1  g1516(.A(n2562), .B(n2549), .Y(n2563));
  AOI21X1 g1517(.A0(n2516), .A1(n2504), .B0(n2563), .Y(n2564));
  OAI21X1 g1518(.A0(n2557), .A1(n2556), .B0(n2564), .Y(n2565));
  NAND2X1 g1519(.A(n2516), .B(n2504), .Y(n2566));
  INVX1   g1520(.A(n2566), .Y(n2567));
  NAND2X1 g1521(.A(n2562), .B(n2549), .Y(n2568));
  INVX1   g1522(.A(n2568), .Y(n2569));
  NOR2X1  g1523(.A(n2562), .B(n2549), .Y(n2570));
  NOR3X1  g1524(.A(n2570), .B(n2569), .C(n2556), .Y(n2571));
  OAI21X1 g1525(.A0(n2531), .A1(n2567), .B0(n2571), .Y(n2572));
  AOI21X1 g1526(.A0(n2572), .A1(n2565), .B0(n2177), .Y(n2573));
  INVX1   g1527(.A(n2563), .Y(n2574));
  NAND2X1 g1528(.A(n2517), .B(n2504), .Y(n2575));
  AOI22X1 g1529(.A0(n2503), .A1(n2516), .B0(n2469), .B1(n2457), .Y(n2576));
  OAI21X1 g1530(.A0(n2519), .A1(n2483), .B0(n2576), .Y(n2577));
  NOR2X1  g1531(.A(n2519), .B(n2482), .Y(n2578));
  AOI22X1 g1532(.A0(n2577), .A1(n2575), .B0(n2418), .B1(n2578), .Y(n2579));
  INVX1   g1533(.A(n2549), .Y(n2580));
  NOR2X1  g1534(.A(n2574), .B(n2579), .Y(n2582));
  AOI21X1 g1535(.A0(n2579), .A1(n2574), .B0(n2582), .Y(n2583));
  OAI22X1 g1536(.A0(n2504), .A1(n2212), .B0(n2211), .B1(n2583), .Y(n2584));
  NOR2X1  g1537(.A(n2583), .B(n2232), .Y(n2585));
  NOR2X1  g1538(.A(n2583), .B(n2231), .Y(n2586));
  NOR3X1  g1539(.A(n2586), .B(n2585), .C(n2584), .Y(n2587));
  INVX1   g1540(.A(n2587), .Y(n2588));
  AOI21X1 g1541(.A0(n2572), .A1(n2565), .B0(n2192), .Y(n2589));
  AOI22X1 g1542(.A0(n2565), .A1(n2572), .B0(n2176), .B1(n2030), .Y(n2590));
  NOR4X1  g1543(.A(n2589), .B(n2588), .C(n2573), .D(n2590), .Y(n2591));
  INVX1   g1544(.A(n2591), .Y(n2592));
  INVX1   g1545(.A(n2562), .Y(n2593));
  XOR2X1  g1546(.A(n2593), .B(n2540), .Y(n2594));
  NAND3X1 g1547(.A(n2498), .B(P1_REG3_REG_10__SCAN_IN), .C(P1_REG3_REG_11__SCAN_IN), .Y(n2595));
  XOR2X1  g1548(.A(n2595), .B(P1_REG3_REG_12__SCAN_IN), .Y(n2596));
  NOR2X1  g1549(.A(n2596), .B(n2144), .Y(n2597));
  INVX1   g1550(.A(P1_REG0_REG_12__SCAN_IN), .Y(n2598));
  NOR3X1  g1551(.A(n2017), .B(n2015), .C(n2598), .Y(n2599));
  AOI22X1 g1552(.A0(n2095), .A1(P1_REG2_REG_12__SCAN_IN), .B0(P1_REG1_REG_12__SCAN_IN), .B1(n2099), .Y(n2600));
  INVX1   g1553(.A(n2600), .Y(n2601));
  NOR3X1  g1554(.A(n2601), .B(n2599), .C(n2597), .Y(n2602));
  OAI22X1 g1555(.A0(n2593), .A1(n2062), .B0(n2092), .B1(n2602), .Y(n2603));
  AOI21X1 g1556(.A0(n2594), .A1(n2063), .B0(n2603), .Y(n2604));
  OAI21X1 g1557(.A0(n2583), .A1(n2049), .B0(n2604), .Y(n2605));
  NOR2X1  g1558(.A(n2605), .B(n2592), .Y(n2606));
  NAND2X1 g1559(.A(n1998), .B(P1_REG0_REG_11__SCAN_IN), .Y(n2607));
  OAI21X1 g1560(.A0(n2606), .A1(n1998), .B0(n2607), .Y(P1_U3486));
  INVX1   g1561(.A(P1_IR_REG_12__SCAN_IN), .Y(n2609));
  NOR2X1  g1562(.A(P1_IR_REG_31__SCAN_IN), .B(n2609), .Y(n2610));
  AOI21X1 g1563(.A0(n1427), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2610), .Y(n2611));
  INVX1   g1564(.A(n2611), .Y(n2612));
  NAND2X1 g1565(.A(n2612), .B(n2003), .Y(n2613));
  OAI21X1 g1566(.A0(n2003), .A1(n1424), .B0(n2613), .Y(n2614));
  XOR2X1  g1567(.A(n2614), .B(n2602), .Y(n2615));
  NOR2X1  g1568(.A(n2570), .B(n2556), .Y(n2616));
  NAND2X1 g1569(.A(n2566), .B(n2529), .Y(n2617));
  AOI21X1 g1570(.A0(n2617), .A1(n2616), .B0(n2569), .Y(n2618));
  OAI21X1 g1571(.A0(n2389), .A1(n2387), .B0(n2471), .Y(n2619));
  AOI21X1 g1572(.A0(n2409), .A1(n2474), .B0(n2424), .Y(n2620));
  AOI21X1 g1573(.A0(n2408), .A1(n2432), .B0(n2620), .Y(n2621));
  NAND3X1 g1574(.A(n2568), .B(n2566), .C(n2528), .Y(n2622));
  AOI21X1 g1575(.A0(n2621), .A1(n2619), .B0(n2622), .Y(n2623));
  NOR2X1  g1576(.A(n2623), .B(n2618), .Y(n2624));
  XOR2X1  g1577(.A(n2624), .B(n2615), .Y(n2625));
  INVX1   g1578(.A(n2625), .Y(n2626));
  OAI21X1 g1579(.A0(n2040), .A1(n2029), .B0(n2626), .Y(n2627));
  OAI21X1 g1580(.A0(n2625), .A1(n2192), .B0(n2627), .Y(n2628));
  NOR4X1  g1581(.A(n2548), .B(n2546), .C(n2544), .D(n2562), .Y(n2629));
  NOR2X1  g1582(.A(n2593), .B(n2549), .Y(n2630));
  INVX1   g1583(.A(n2630), .Y(n2631));
  OAI21X1 g1584(.A0(n2629), .A1(n2579), .B0(n2631), .Y(n2632));
  NOR2X1  g1585(.A(n2632), .B(n2615), .Y(n2633));
  INVX1   g1586(.A(n2602), .Y(n2634));
  XOR2X1  g1587(.A(n2614), .B(n2634), .Y(n2635));
  AOI21X1 g1588(.A0(n2615), .A1(n2632), .B0(n2633), .Y(n2637));
  AOI22X1 g1589(.A0(n2580), .A1(n2081), .B0(n2041), .B1(n2626), .Y(n2638));
  OAI21X1 g1590(.A0(n2637), .A1(n2231), .B0(n2638), .Y(n2639));
  AOI21X1 g1591(.A0(n2232), .A1(n2211), .B0(n2637), .Y(n2640));
  NOR4X1  g1592(.A(n2516), .B(n2469), .C(n2494), .D(n2562), .Y(n2641));
  INVX1   g1593(.A(n2614), .Y(n2642));
  XOR2X1  g1594(.A(n2642), .B(n2641), .Y(n2643));
  NAND4X1 g1595(.A(P1_REG3_REG_10__SCAN_IN), .B(P1_REG3_REG_12__SCAN_IN), .C(P1_REG3_REG_11__SCAN_IN), .D(n2498), .Y(n2644));
  XOR2X1  g1596(.A(n2644), .B(P1_REG3_REG_13__SCAN_IN), .Y(n2645));
  INVX1   g1597(.A(n2645), .Y(n2646));
  AOI22X1 g1598(.A0(n2100), .A1(n2646), .B0(n2094), .B1(P1_REG0_REG_13__SCAN_IN), .Y(n2647));
  AOI22X1 g1599(.A0(n2095), .A1(P1_REG2_REG_13__SCAN_IN), .B0(P1_REG1_REG_13__SCAN_IN), .B1(n2099), .Y(n2648));
  NAND2X1 g1600(.A(n2648), .B(n2647), .Y(n2649));
  INVX1   g1601(.A(n2649), .Y(n2650));
  OAI22X1 g1602(.A0(n2642), .A1(n2062), .B0(n2092), .B1(n2650), .Y(n2651));
  AOI21X1 g1603(.A0(n2643), .A1(n2063), .B0(n2651), .Y(n2652));
  OAI21X1 g1604(.A0(n2637), .A1(n2049), .B0(n2652), .Y(n2653));
  NOR4X1  g1605(.A(n2640), .B(n2639), .C(n2628), .D(n2653), .Y(n2654));
  NAND2X1 g1606(.A(n1998), .B(P1_REG0_REG_12__SCAN_IN), .Y(n2655));
  OAI21X1 g1607(.A0(n2654), .A1(n1998), .B0(n2655), .Y(P1_U3489));
  NAND2X1 g1608(.A(n2614), .B(n2634), .Y(n2657));
  INVX1   g1609(.A(n2657), .Y(n2658));
  NOR2X1  g1610(.A(n2658), .B(n2632), .Y(n2659));
  INVX1   g1611(.A(n2659), .Y(n2660));
  NOR2X1  g1612(.A(P1_IR_REG_31__SCAN_IN), .B(n1444), .Y(n2661));
  AOI21X1 g1613(.A0(n1445), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2661), .Y(n2662));
  INVX1   g1614(.A(n2662), .Y(n2663));
  NAND2X1 g1615(.A(n2663), .B(n2003), .Y(n2664));
  OAI21X1 g1616(.A0(n2003), .A1(n1443), .B0(n2664), .Y(n2665));
  NOR2X1  g1617(.A(n2665), .B(n2649), .Y(n2666));
  AOI21X1 g1618(.A0(n2642), .A1(n2602), .B0(n2666), .Y(n2667));
  INVX1   g1619(.A(n2667), .Y(n2668));
  AOI21X1 g1620(.A0(n2665), .A1(n2649), .B0(n2668), .Y(n2669));
  OAI21X1 g1621(.A0(n2614), .A1(n2634), .B0(n2632), .Y(n2670));
  INVX1   g1622(.A(n2665), .Y(n2671));
  NOR2X1  g1623(.A(n2671), .B(n2649), .Y(n2672));
  NOR2X1  g1624(.A(n2665), .B(n2650), .Y(n2673));
  NOR3X1  g1625(.A(n2673), .B(n2672), .C(n2658), .Y(n2674));
  AOI22X1 g1626(.A0(n2670), .A1(n2674), .B0(n2669), .B1(n2660), .Y(n2675));
  INVX1   g1627(.A(n2675), .Y(n2676));
  AOI21X1 g1628(.A0(n2232), .A1(n2231), .B0(n2676), .Y(n2677));
  XOR2X1  g1629(.A(n2665), .B(n2650), .Y(n2678));
  NOR2X1  g1630(.A(n2614), .B(n2602), .Y(n2679));
  INVX1   g1631(.A(n2618), .Y(n2680));
  INVX1   g1632(.A(n2622), .Y(n2681));
  OAI21X1 g1633(.A0(n2476), .A1(n2473), .B0(n2681), .Y(n2682));
  AOI22X1 g1634(.A0(n2680), .A1(n2682), .B0(n2614), .B1(n2602), .Y(n2683));
  NOR2X1  g1635(.A(n2683), .B(n2679), .Y(n2684));
  XOR2X1  g1636(.A(n2684), .B(n2678), .Y(n2685));
  OAI22X1 g1637(.A0(n2676), .A1(n2211), .B0(n2192), .B1(n2685), .Y(n2686));
  INVX1   g1638(.A(n2685), .Y(n2687));
  AOI22X1 g1639(.A0(n2634), .A1(n2081), .B0(n2041), .B1(n2687), .Y(n2688));
  OAI21X1 g1640(.A0(n2040), .A1(n2029), .B0(n2687), .Y(n2689));
  NAND2X1 g1641(.A(n2689), .B(n2688), .Y(n2690));
  INVX1   g1642(.A(n2641), .Y(n2691));
  NOR2X1  g1643(.A(n2614), .B(n2691), .Y(n2692));
  XOR2X1  g1644(.A(n2671), .B(n2692), .Y(n2693));
  INVX1   g1645(.A(P1_REG3_REG_14__SCAN_IN), .Y(n2694));
  INVX1   g1646(.A(P1_REG3_REG_13__SCAN_IN), .Y(n2695));
  NOR2X1  g1647(.A(n2644), .B(n2695), .Y(n2696));
  XOR2X1  g1648(.A(n2696), .B(n2694), .Y(n2697));
  INVX1   g1649(.A(n2697), .Y(n2698));
  INVX1   g1650(.A(P1_REG1_REG_14__SCAN_IN), .Y(n2699));
  AOI22X1 g1651(.A0(n2094), .A1(P1_REG0_REG_14__SCAN_IN), .B0(P1_REG2_REG_14__SCAN_IN), .B1(n2095), .Y(n2700));
  OAI21X1 g1652(.A0(n2143), .A1(n2699), .B0(n2700), .Y(n2701));
  AOI21X1 g1653(.A0(n2698), .A1(n2100), .B0(n2701), .Y(n2702));
  OAI22X1 g1654(.A0(n2671), .A1(n2062), .B0(n2092), .B1(n2702), .Y(n2703));
  AOI21X1 g1655(.A0(n2693), .A1(n2063), .B0(n2703), .Y(n2704));
  OAI21X1 g1656(.A0(n2676), .A1(n2049), .B0(n2704), .Y(n2705));
  NOR4X1  g1657(.A(n2690), .B(n2686), .C(n2677), .D(n2705), .Y(n2706));
  NAND2X1 g1658(.A(n1998), .B(P1_REG0_REG_13__SCAN_IN), .Y(n2707));
  OAI21X1 g1659(.A0(n2706), .A1(n1998), .B0(n2707), .Y(P1_U3492));
  INVX1   g1660(.A(n2702), .Y(n2709));
  NOR2X1  g1661(.A(P1_IR_REG_31__SCAN_IN), .B(n1462), .Y(n2710));
  AOI21X1 g1662(.A0(n1466), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2710), .Y(n2711));
  INVX1   g1663(.A(n2711), .Y(n2712));
  NOR2X1  g1664(.A(n2003), .B(n1461), .Y(n2713));
  AOI21X1 g1665(.A0(n2712), .A1(n2003), .B0(n2713), .Y(n2714));
  XOR2X1  g1666(.A(n2714), .B(n2709), .Y(n2715));
  INVX1   g1667(.A(n2673), .Y(n2717));
  OAI22X1 g1668(.A0(n2671), .A1(n2649), .B0(n2679), .B1(n2683), .Y(n2718));
  NAND2X1 g1669(.A(n2718), .B(n2717), .Y(n2719));
  XOR2X1  g1670(.A(n2719), .B(n4850), .Y(n2720));
  NOR2X1  g1671(.A(n2720), .B(n2177), .Y(n2721));
  OAI21X1 g1672(.A0(n2671), .A1(n2650), .B0(n2657), .Y(n2722));
  AOI21X1 g1673(.A0(n2667), .A1(n2630), .B0(n2722), .Y(n2723));
  OAI21X1 g1674(.A0(n2562), .A1(n2580), .B0(n2667), .Y(n2724));
  OAI22X1 g1675(.A0(n2723), .A1(n2666), .B0(n2579), .B1(n2724), .Y(n2725));
  XOR2X1  g1676(.A(n2725), .B(n2715), .Y(n2726));
  INVX1   g1677(.A(n2726), .Y(n2727));
  AOI22X1 g1678(.A0(n2649), .A1(n2081), .B0(n2043), .B1(n2727), .Y(n2728));
  INVX1   g1679(.A(n2728), .Y(n2729));
  OAI21X1 g1680(.A0(n2045), .A1(n2038), .B0(n2727), .Y(n2730));
  INVX1   g1681(.A(n2730), .Y(n2731));
  INVX1   g1682(.A(n2720), .Y(n2732));
  OAI21X1 g1683(.A0(n2040), .A1(n2029), .B0(n2732), .Y(n2733));
  OAI21X1 g1684(.A0(n2720), .A1(n2192), .B0(n2733), .Y(n2734));
  NOR4X1  g1685(.A(n2731), .B(n2729), .C(n2721), .D(n2734), .Y(n2735));
  INVX1   g1686(.A(n2735), .Y(n2736));
  NOR2X1  g1687(.A(n2726), .B(n2049), .Y(n2737));
  NOR3X1  g1688(.A(n2665), .B(n2614), .C(n2691), .Y(n2738));
  NAND4X1 g1689(.A(n2671), .B(n2642), .C(n2641), .D(n2714), .Y(n2739));
  OAI21X1 g1690(.A0(n2714), .A1(n2738), .B0(n2739), .Y(n2740));
  INVX1   g1691(.A(n2714), .Y(n2741));
  INVX1   g1692(.A(P1_REG3_REG_15__SCAN_IN), .Y(n2742));
  NOR3X1  g1693(.A(n2644), .B(n2694), .C(n2695), .Y(n2743));
  XOR2X1  g1694(.A(n2743), .B(n2742), .Y(n2744));
  INVX1   g1695(.A(n2744), .Y(n2745));
  NAND3X1 g1696(.A(n2745), .B(n2017), .C(n2015), .Y(n2746));
  NAND3X1 g1697(.A(n2017), .B(n2021), .C(P1_REG1_REG_15__SCAN_IN), .Y(n2747));
  AOI22X1 g1698(.A0(n2094), .A1(P1_REG0_REG_15__SCAN_IN), .B0(P1_REG2_REG_15__SCAN_IN), .B1(n2095), .Y(n2748));
  NAND3X1 g1699(.A(n2748), .B(n2747), .C(n2746), .Y(n2749));
  AOI22X1 g1700(.A0(n2741), .A1(n2302), .B0(n2050), .B1(n2749), .Y(n2750));
  OAI21X1 g1701(.A0(n2740), .A1(n2064), .B0(n2750), .Y(n2751));
  NOR3X1  g1702(.A(n2751), .B(n2737), .C(n2736), .Y(n2752));
  NAND2X1 g1703(.A(n1998), .B(P1_REG0_REG_14__SCAN_IN), .Y(n2753));
  OAI21X1 g1704(.A0(n2752), .A1(n1998), .B0(n2753), .Y(P1_U3495));
  NOR2X1  g1705(.A(P1_IR_REG_31__SCAN_IN), .B(n1489), .Y(n2755));
  AOI21X1 g1706(.A0(n1490), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2755), .Y(n2756));
  INVX1   g1707(.A(n2756), .Y(n2757));
  NOR2X1  g1708(.A(n2003), .B(n1488), .Y(n2758));
  AOI21X1 g1709(.A0(n2757), .A1(n2003), .B0(n2758), .Y(n2759));
  XOR2X1  g1710(.A(n2759), .B(n2749), .Y(n2760));
  NOR2X1  g1711(.A(n2714), .B(n2709), .Y(n2761));
  INVX1   g1712(.A(n2761), .Y(n2762));
  NOR2X1  g1713(.A(n2741), .B(n2702), .Y(n2763));
  AOI21X1 g1714(.A0(n2719), .A1(n2762), .B0(n2763), .Y(n2764));
  XOR2X1  g1715(.A(n2764), .B(n2760), .Y(n2765));
  NOR2X1  g1716(.A(n2765), .B(n2177), .Y(n2766));
  NOR2X1  g1717(.A(n2714), .B(n2702), .Y(n2767));
  NOR2X1  g1718(.A(n2741), .B(n2709), .Y(n2768));
  INVX1   g1719(.A(n2768), .Y(n2769));
  AOI21X1 g1720(.A0(n2769), .A1(n2725), .B0(n2767), .Y(n2770));
  INVX1   g1721(.A(n2770), .Y(n2771));
  XOR2X1  g1722(.A(n2771), .B(n2760), .Y(n2772));
  INVX1   g1723(.A(n2772), .Y(n2773));
  AOI22X1 g1724(.A0(n2709), .A1(n2081), .B0(n2043), .B1(n2773), .Y(n2774));
  INVX1   g1725(.A(n2774), .Y(n2775));
  OAI21X1 g1726(.A0(n2045), .A1(n2038), .B0(n2773), .Y(n2776));
  INVX1   g1727(.A(n2776), .Y(n2777));
  INVX1   g1728(.A(n2765), .Y(n2778));
  OAI21X1 g1729(.A0(n2040), .A1(n2029), .B0(n2778), .Y(n2779));
  OAI21X1 g1730(.A0(n2765), .A1(n2192), .B0(n2779), .Y(n2780));
  NOR4X1  g1731(.A(n2777), .B(n2775), .C(n2766), .D(n2780), .Y(n2781));
  INVX1   g1732(.A(n2781), .Y(n2782));
  NOR2X1  g1733(.A(n2772), .B(n2049), .Y(n2783));
  XOR2X1  g1734(.A(n2759), .B(n2739), .Y(n2784));
  INVX1   g1735(.A(n2759), .Y(n2785));
  NOR4X1  g1736(.A(n2694), .B(n2695), .C(n2742), .D(n2644), .Y(n2786));
  XOR2X1  g1737(.A(n2786), .B(P1_REG3_REG_16__SCAN_IN), .Y(n2787));
  INVX1   g1738(.A(P1_REG1_REG_16__SCAN_IN), .Y(n2788));
  AOI22X1 g1739(.A0(n2094), .A1(P1_REG0_REG_16__SCAN_IN), .B0(P1_REG2_REG_16__SCAN_IN), .B1(n2095), .Y(n2789));
  OAI21X1 g1740(.A0(n2143), .A1(n2788), .B0(n2789), .Y(n2790));
  AOI21X1 g1741(.A0(n2787), .A1(n2100), .B0(n2790), .Y(n2791));
  INVX1   g1742(.A(n2791), .Y(n2792));
  AOI22X1 g1743(.A0(n2785), .A1(n2302), .B0(n2050), .B1(n2792), .Y(n2793));
  OAI21X1 g1744(.A0(n2784), .A1(n2064), .B0(n2793), .Y(n2794));
  NOR3X1  g1745(.A(n2794), .B(n2783), .C(n2782), .Y(n2795));
  NAND2X1 g1746(.A(n1998), .B(P1_REG0_REG_15__SCAN_IN), .Y(n2796));
  OAI21X1 g1747(.A0(n2795), .A1(n1998), .B0(n2796), .Y(P1_U3498));
  INVX1   g1748(.A(n2749), .Y(n2798));
  NOR2X1  g1749(.A(n2785), .B(n2798), .Y(n2799));
  NOR2X1  g1750(.A(n2759), .B(n2749), .Y(n2801));
  NOR2X1  g1751(.A(P1_IR_REG_31__SCAN_IN), .B(n1509), .Y(n2802));
  AOI21X1 g1752(.A0(n1522), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2802), .Y(n2803));
  INVX1   g1753(.A(n2803), .Y(n2804));
  NOR2X1  g1754(.A(n2003), .B(n1508), .Y(n2805));
  AOI21X1 g1755(.A0(n2804), .A1(n2003), .B0(n2805), .Y(n2806));
  XOR2X1  g1756(.A(n2806), .B(n2792), .Y(n2807));
  NOR2X1  g1757(.A(n2807), .B(n2801), .Y(n2808));
  OAI21X1 g1758(.A0(n4806), .A1(n2799), .B0(n2808), .Y(n2809));
  NOR2X1  g1759(.A(n2806), .B(n2792), .Y(n2810));
  INVX1   g1760(.A(n2806), .Y(n2811));
  OAI22X1 g1761(.A0(n2791), .A1(n2811), .B0(n2785), .B1(n2798), .Y(n2812));
  NOR2X1  g1762(.A(n2812), .B(n2810), .Y(n2813));
  OAI21X1 g1763(.A0(n2764), .A1(n2801), .B0(n2813), .Y(n2814));
  AOI21X1 g1764(.A0(n2814), .A1(n2809), .B0(n2177), .Y(n2815));
  NOR2X1  g1765(.A(n2759), .B(n2798), .Y(n2816));
  INVX1   g1766(.A(n2816), .Y(n2817));
  NOR2X1  g1767(.A(n2785), .B(n2749), .Y(n2818));
  OAI21X1 g1768(.A0(n2818), .A1(n2770), .B0(n2817), .Y(n2819));
  NOR2X1  g1769(.A(n2819), .B(n2807), .Y(n2820));
  AOI21X1 g1770(.A0(n2807), .A1(n2819), .B0(n2820), .Y(n2823));
  INVX1   g1771(.A(n2823), .Y(n2824));
  AOI22X1 g1772(.A0(n2749), .A1(n2081), .B0(n2043), .B1(n2824), .Y(n2825));
  OAI21X1 g1773(.A0(n2045), .A1(n2038), .B0(n2824), .Y(n2826));
  NAND2X1 g1774(.A(n2826), .B(n2825), .Y(n2827));
  AOI21X1 g1775(.A0(n2814), .A1(n2809), .B0(n2192), .Y(n2828));
  AOI22X1 g1776(.A0(n2809), .A1(n2814), .B0(n2176), .B1(n2030), .Y(n2829));
  NOR4X1  g1777(.A(n2828), .B(n2827), .C(n2815), .D(n2829), .Y(n2830));
  INVX1   g1778(.A(n2830), .Y(n2831));
  NOR2X1  g1779(.A(n2785), .B(n2739), .Y(n2832));
  XOR2X1  g1780(.A(n2806), .B(n2832), .Y(n2833));
  NAND2X1 g1781(.A(n2786), .B(P1_REG3_REG_16__SCAN_IN), .Y(n2834));
  XOR2X1  g1782(.A(n2834), .B(P1_REG3_REG_17__SCAN_IN), .Y(n2835));
  INVX1   g1783(.A(n2835), .Y(n2836));
  NAND3X1 g1784(.A(n2836), .B(n2017), .C(n2015), .Y(n2837));
  NAND3X1 g1785(.A(n2017), .B(n2021), .C(P1_REG1_REG_17__SCAN_IN), .Y(n2838));
  AOI22X1 g1786(.A0(n2094), .A1(P1_REG0_REG_17__SCAN_IN), .B0(P1_REG2_REG_17__SCAN_IN), .B1(n2095), .Y(n2839));
  NAND3X1 g1787(.A(n2839), .B(n2838), .C(n2837), .Y(n2840));
  INVX1   g1788(.A(n2840), .Y(n2841));
  OAI22X1 g1789(.A0(n2806), .A1(n2062), .B0(n2092), .B1(n2841), .Y(n2842));
  AOI21X1 g1790(.A0(n2833), .A1(n2063), .B0(n2842), .Y(n2843));
  OAI21X1 g1791(.A0(n2823), .A1(n2049), .B0(n2843), .Y(n2844));
  NOR2X1  g1792(.A(n2844), .B(n2831), .Y(n2845));
  NAND2X1 g1793(.A(n1998), .B(P1_REG0_REG_16__SCAN_IN), .Y(n2846));
  OAI21X1 g1794(.A0(n2845), .A1(n1998), .B0(n2846), .Y(P1_U3501));
  NOR2X1  g1795(.A(n2806), .B(n2791), .Y(n2848));
  NOR2X1  g1796(.A(P1_IR_REG_31__SCAN_IN), .B(n1539), .Y(n2849));
  AOI21X1 g1797(.A0(n1540), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2849), .Y(n2850));
  INVX1   g1798(.A(n2850), .Y(n2851));
  NOR2X1  g1799(.A(n2003), .B(n1538), .Y(n2852));
  AOI21X1 g1800(.A0(n2851), .A1(n2003), .B0(n2852), .Y(n2853));
  INVX1   g1801(.A(n2853), .Y(n2854));
  AOI22X1 g1802(.A0(n2841), .A1(n2853), .B0(n2806), .B1(n2791), .Y(n2855));
  INVX1   g1803(.A(n2855), .Y(n2856));
  AOI21X1 g1804(.A0(n2854), .A1(n2840), .B0(n2856), .Y(n2857));
  OAI21X1 g1805(.A0(n2848), .A1(n2819), .B0(n2857), .Y(n2858));
  INVX1   g1806(.A(n2819), .Y(n2859));
  AOI21X1 g1807(.A0(n2806), .A1(n2791), .B0(n2859), .Y(n2860));
  NOR2X1  g1808(.A(n2853), .B(n2840), .Y(n2861));
  NOR2X1  g1809(.A(n2854), .B(n2841), .Y(n2862));
  NOR3X1  g1810(.A(n2862), .B(n2861), .C(n2848), .Y(n2863));
  INVX1   g1811(.A(n2863), .Y(n2864));
  OAI21X1 g1812(.A0(n2864), .A1(n2860), .B0(n2858), .Y(n2865));
  INVX1   g1813(.A(n2865), .Y(n2866));
  OAI21X1 g1814(.A0(n2045), .A1(n2038), .B0(n2866), .Y(n2867));
  XOR2X1  g1815(.A(n2853), .B(n2840), .Y(n2868));
  INVX1   g1816(.A(n2810), .Y(n2869));
  NOR3X1  g1817(.A(n2801), .B(n2741), .C(n2702), .Y(n2870));
  OAI21X1 g1818(.A0(n2870), .A1(n2812), .B0(n2869), .Y(n2871));
  INVX1   g1819(.A(n2871), .Y(n2872));
  NOR3X1  g1820(.A(n2810), .B(n2801), .C(n2761), .Y(n2873));
  INVX1   g1821(.A(n2873), .Y(n2874));
  AOI21X1 g1822(.A0(n2718), .A1(n2717), .B0(n2874), .Y(n2875));
  NOR2X1  g1823(.A(n2875), .B(n2872), .Y(n2876));
  XOR2X1  g1824(.A(n2876), .B(n2868), .Y(n2877));
  INVX1   g1825(.A(n2877), .Y(n2878));
  AOI22X1 g1826(.A0(n2866), .A1(n2043), .B0(n2034), .B1(n2878), .Y(n2879));
  AOI22X1 g1827(.A0(n2792), .A1(n2081), .B0(n2041), .B1(n2878), .Y(n2880));
  OAI21X1 g1828(.A0(n2040), .A1(n2029), .B0(n2878), .Y(n2881));
  NAND4X1 g1829(.A(n2880), .B(n2879), .C(n2867), .D(n2881), .Y(n2882));
  NOR3X1  g1830(.A(n2811), .B(n2785), .C(n2739), .Y(n2883));
  XOR2X1  g1831(.A(n2853), .B(n2883), .Y(n2884));
  NAND3X1 g1832(.A(n2786), .B(P1_REG3_REG_16__SCAN_IN), .C(P1_REG3_REG_17__SCAN_IN), .Y(n2885));
  XOR2X1  g1833(.A(n2885), .B(P1_REG3_REG_18__SCAN_IN), .Y(n2886));
  INVX1   g1834(.A(n2886), .Y(n2887));
  INVX1   g1835(.A(P1_REG1_REG_18__SCAN_IN), .Y(n2888));
  AOI22X1 g1836(.A0(n2094), .A1(P1_REG0_REG_18__SCAN_IN), .B0(P1_REG2_REG_18__SCAN_IN), .B1(n2095), .Y(n2889));
  OAI21X1 g1837(.A0(n2143), .A1(n2888), .B0(n2889), .Y(n2890));
  AOI21X1 g1838(.A0(n2887), .A1(n2100), .B0(n2890), .Y(n2891));
  OAI22X1 g1839(.A0(n2853), .A1(n2062), .B0(n2092), .B1(n2891), .Y(n2892));
  AOI21X1 g1840(.A0(n2884), .A1(n2063), .B0(n2892), .Y(n2893));
  OAI21X1 g1841(.A0(n2865), .A1(n2049), .B0(n2893), .Y(n2894));
  NOR2X1  g1842(.A(n2894), .B(n2882), .Y(n2895));
  NAND2X1 g1843(.A(n1998), .B(P1_REG0_REG_17__SCAN_IN), .Y(n2896));
  OAI21X1 g1844(.A0(n2895), .A1(n1998), .B0(n2896), .Y(P1_U3504));
  NAND2X1 g1845(.A(n2854), .B(n2848), .Y(n2898));
  OAI21X1 g1846(.A0(n2854), .A1(n2848), .B0(n2840), .Y(n2899));
  NAND2X1 g1847(.A(n2899), .B(n2898), .Y(n2900));
  AOI21X1 g1848(.A0(n2855), .A1(n2819), .B0(n2900), .Y(n2901));
  INVX1   g1849(.A(n2891), .Y(n2902));
  NOR2X1  g1850(.A(P1_IR_REG_31__SCAN_IN), .B(n1562), .Y(n2903));
  AOI21X1 g1851(.A0(n1568), .A1(P1_IR_REG_31__SCAN_IN), .B0(n2903), .Y(n2904));
  INVX1   g1852(.A(n2904), .Y(n2905));
  NOR2X1  g1853(.A(n2003), .B(n1556), .Y(n2906));
  AOI21X1 g1854(.A0(n2905), .A1(n2003), .B0(n2906), .Y(n2907));
  XOR2X1  g1855(.A(n2907), .B(n2891), .Y(n2910));
  NOR2X1  g1856(.A(n2910), .B(n2901), .Y(n2911));
  AOI21X1 g1857(.A0(n2910), .A1(n2901), .B0(n2911), .Y(n2912));
  INVX1   g1858(.A(n2912), .Y(n2913));
  AOI22X1 g1859(.A0(n2840), .A1(n2081), .B0(n2043), .B1(n2913), .Y(n2914));
  OAI21X1 g1860(.A0(n2045), .A1(n2038), .B0(n2913), .Y(n2915));
  INVX1   g1861(.A(n2862), .Y(n2916));
  OAI22X1 g1862(.A0(n2872), .A1(n2875), .B0(n2853), .B1(n2840), .Y(n2917));
  NAND2X1 g1863(.A(n2917), .B(n2916), .Y(n2918));
  XOR2X1  g1864(.A(n2918), .B(n2910), .Y(n2919));
  INVX1   g1865(.A(n2919), .Y(n2920));
  OAI21X1 g1866(.A0(n2041), .A1(n2040), .B0(n2920), .Y(n2921));
  OAI21X1 g1867(.A0(n2034), .A1(n2029), .B0(n2920), .Y(n2922));
  NAND4X1 g1868(.A(n2921), .B(n2915), .C(n2914), .D(n2922), .Y(n2923));
  NAND2X1 g1869(.A(n2853), .B(n2883), .Y(n2924));
  INVX1   g1870(.A(n2907), .Y(n2925));
  XOR2X1  g1871(.A(n2925), .B(n2924), .Y(n2926));
  NAND4X1 g1872(.A(P1_REG3_REG_16__SCAN_IN), .B(P1_REG3_REG_17__SCAN_IN), .C(P1_REG3_REG_18__SCAN_IN), .D(n2786), .Y(n2927));
  XOR2X1  g1873(.A(n2927), .B(P1_REG3_REG_19__SCAN_IN), .Y(n2928));
  INVX1   g1874(.A(n2928), .Y(n2929));
  NAND3X1 g1875(.A(n2017), .B(n2021), .C(P1_REG1_REG_19__SCAN_IN), .Y(n2930));
  AOI22X1 g1876(.A0(n2094), .A1(P1_REG0_REG_19__SCAN_IN), .B0(P1_REG2_REG_19__SCAN_IN), .B1(n2095), .Y(n2931));
  NAND2X1 g1877(.A(n2931), .B(n2930), .Y(n2932));
  AOI21X1 g1878(.A0(n2929), .A1(n2100), .B0(n2932), .Y(n2933));
  OAI22X1 g1879(.A0(n2907), .A1(n2062), .B0(n2092), .B1(n2933), .Y(n2934));
  AOI21X1 g1880(.A0(n2926), .A1(n2063), .B0(n2934), .Y(n2935));
  OAI21X1 g1881(.A0(n2912), .A1(n2049), .B0(n2935), .Y(n2936));
  NOR2X1  g1882(.A(n2936), .B(n2923), .Y(n2937));
  NAND2X1 g1883(.A(n1998), .B(P1_REG0_REG_18__SCAN_IN), .Y(n2938));
  OAI21X1 g1884(.A0(n2937), .A1(n1998), .B0(n2938), .Y(P1_U3507));
  NAND2X1 g1885(.A(n2003), .B(n2037), .Y(n2940));
  OAI21X1 g1886(.A0(n2003), .A1(n1584), .B0(n2940), .Y(n2941));
  XOR2X1  g1887(.A(n2941), .B(n2933), .Y(n2942));
  AOI21X1 g1888(.A0(n2917), .A1(n2916), .B0(n2891), .Y(n2943));
  NAND3X1 g1889(.A(n2917), .B(n2891), .C(n2916), .Y(n2944));
  AOI21X1 g1890(.A0(n2944), .A1(n2907), .B0(n2943), .Y(n2945));
  XOR2X1  g1891(.A(n2945), .B(n2942), .Y(n2946));
  NOR2X1  g1892(.A(n2946), .B(n2177), .Y(n2947));
  INVX1   g1893(.A(n2901), .Y(n2948));
  NOR2X1  g1894(.A(n2925), .B(n2902), .Y(n2949));
  INVX1   g1895(.A(n2949), .Y(n2950));
  NOR2X1  g1896(.A(n2907), .B(n2891), .Y(n2951));
  AOI21X1 g1897(.A0(n2950), .A1(n2948), .B0(n2951), .Y(n2952));
  INVX1   g1898(.A(n2952), .Y(n2953));
  NOR2X1  g1899(.A(n2953), .B(n2942), .Y(n2954));
  AOI21X1 g1900(.A0(n2942), .A1(n2953), .B0(n2954), .Y(n2956));
  OAI22X1 g1901(.A0(n2891), .A1(n2212), .B0(n2211), .B1(n2956), .Y(n2957));
  AOI21X1 g1902(.A0(n2232), .A1(n2231), .B0(n2956), .Y(n2958));
  NOR3X1  g1903(.A(n2958), .B(n2957), .C(n2947), .Y(n2959));
  NOR2X1  g1904(.A(n2946), .B(n2192), .Y(n2960));
  AOI21X1 g1905(.A0(n2176), .A1(n2030), .B0(n2946), .Y(n2961));
  NOR2X1  g1906(.A(n2961), .B(n2960), .Y(n2962));
  NAND2X1 g1907(.A(n2962), .B(n2959), .Y(n2963));
  NOR2X1  g1908(.A(n2925), .B(n2924), .Y(n2964));
  NOR2X1  g1909(.A(n2003), .B(n1584), .Y(n2965));
  AOI21X1 g1910(.A0(n2003), .A1(n2037), .B0(n2965), .Y(n2966));
  XOR2X1  g1911(.A(n2966), .B(n2964), .Y(n2967));
  INVX1   g1912(.A(P1_REG3_REG_20__SCAN_IN), .Y(n2968));
  INVX1   g1913(.A(P1_REG3_REG_19__SCAN_IN), .Y(n2969));
  NOR2X1  g1914(.A(n2927), .B(n2969), .Y(n2970));
  XOR2X1  g1915(.A(n2970), .B(n2968), .Y(n2971));
  INVX1   g1916(.A(n2971), .Y(n2972));
  NAND3X1 g1917(.A(n2017), .B(n2021), .C(P1_REG1_REG_20__SCAN_IN), .Y(n2973));
  AOI22X1 g1918(.A0(n2094), .A1(P1_REG0_REG_20__SCAN_IN), .B0(P1_REG2_REG_20__SCAN_IN), .B1(n2095), .Y(n2974));
  NAND2X1 g1919(.A(n2974), .B(n2973), .Y(n2975));
  AOI21X1 g1920(.A0(n2972), .A1(n2100), .B0(n2975), .Y(n2976));
  OAI22X1 g1921(.A0(n2966), .A1(n2062), .B0(n2092), .B1(n2976), .Y(n2977));
  AOI21X1 g1922(.A0(n2967), .A1(n2063), .B0(n2977), .Y(n2978));
  OAI21X1 g1923(.A0(n2956), .A1(n2049), .B0(n2978), .Y(n2979));
  NOR2X1  g1924(.A(n2979), .B(n2963), .Y(n2980));
  NAND2X1 g1925(.A(n1998), .B(P1_REG0_REG_19__SCAN_IN), .Y(n2981));
  OAI21X1 g1926(.A0(n2980), .A1(n1998), .B0(n2981), .Y(P1_U3509));
  NOR2X1  g1927(.A(n2003), .B(n1607), .Y(n2983));
  XOR2X1  g1928(.A(n2983), .B(n2976), .Y(n2984));
  NAND2X1 g1929(.A(n2941), .B(n2933), .Y(n2985));
  NOR2X1  g1930(.A(n2941), .B(n2933), .Y(n2986));
  INVX1   g1931(.A(n2679), .Y(n2987));
  NAND2X1 g1932(.A(n2614), .B(n2602), .Y(n2988));
  OAI21X1 g1933(.A0(n2623), .A1(n2618), .B0(n2988), .Y(n2989));
  AOI21X1 g1934(.A0(n2989), .A1(n2987), .B0(n2672), .Y(n2990));
  OAI21X1 g1935(.A0(n2990), .A1(n2673), .B0(n2873), .Y(n2991));
  AOI21X1 g1936(.A0(n2991), .A1(n2871), .B0(n2861), .Y(n2992));
  OAI21X1 g1937(.A0(n2992), .A1(n2862), .B0(n2902), .Y(n2993));
  NOR3X1  g1938(.A(n2992), .B(n2902), .C(n2862), .Y(n2994));
  OAI21X1 g1939(.A0(n2994), .A1(n2925), .B0(n2993), .Y(n2995));
  AOI21X1 g1940(.A0(n2995), .A1(n2985), .B0(n2986), .Y(n2996));
  XOR2X1  g1941(.A(n2996), .B(n2984), .Y(n2997));
  NOR2X1  g1942(.A(n2997), .B(n2177), .Y(n2998));
  INVX1   g1943(.A(n2998), .Y(n2999));
  NOR2X1  g1944(.A(n2966), .B(n2933), .Y(n3000));
  INVX1   g1945(.A(n2976), .Y(n3001));
  INVX1   g1946(.A(n2933), .Y(n3002));
  OAI22X1 g1947(.A0(n3001), .A1(n2983), .B0(n2941), .B1(n3002), .Y(n3003));
  AOI21X1 g1948(.A0(n2983), .A1(n3001), .B0(n3003), .Y(n3004));
  OAI21X1 g1949(.A0(n3000), .A1(n2953), .B0(n3004), .Y(n3005));
  NOR2X1  g1950(.A(n2941), .B(n3002), .Y(n3006));
  NOR3X1  g1951(.A(n3001), .B(n2003), .C(n1607), .Y(n3007));
  NOR2X1  g1952(.A(n2983), .B(n2976), .Y(n3008));
  NOR3X1  g1953(.A(n3008), .B(n3007), .C(n3000), .Y(n3009));
  OAI21X1 g1954(.A0(n3006), .A1(n2952), .B0(n3009), .Y(n3010));
  NAND2X1 g1955(.A(n3010), .B(n3005), .Y(n3011));
  OAI22X1 g1956(.A0(n2933), .A1(n2212), .B0(n2211), .B1(n3011), .Y(n3012));
  AOI21X1 g1957(.A0(n2232), .A1(n2231), .B0(n3011), .Y(n3013));
  NOR2X1  g1958(.A(n3013), .B(n3012), .Y(n3014));
  NOR2X1  g1959(.A(n2997), .B(n2192), .Y(n3015));
  AOI21X1 g1960(.A0(n2176), .A1(n2030), .B0(n2997), .Y(n3016));
  NOR2X1  g1961(.A(n3016), .B(n3015), .Y(n3017));
  NAND3X1 g1962(.A(n3017), .B(n3014), .C(n2999), .Y(n3018));
  NAND4X1 g1963(.A(n2907), .B(n2853), .C(n2883), .D(n2966), .Y(n3019));
  XOR2X1  g1964(.A(n2983), .B(n3019), .Y(n3020));
  INVX1   g1965(.A(n2983), .Y(n3021));
  INVX1   g1966(.A(P1_REG3_REG_21__SCAN_IN), .Y(n3022));
  NOR3X1  g1967(.A(n2927), .B(n2969), .C(n2968), .Y(n3023));
  XOR2X1  g1968(.A(n3023), .B(n3022), .Y(n3024));
  AOI22X1 g1969(.A0(n2094), .A1(P1_REG0_REG_21__SCAN_IN), .B0(P1_REG2_REG_21__SCAN_IN), .B1(n2095), .Y(n3025));
  INVX1   g1970(.A(n3025), .Y(n3026));
  AOI21X1 g1971(.A0(n2099), .A1(P1_REG1_REG_21__SCAN_IN), .B0(n3026), .Y(n3027));
  OAI21X1 g1972(.A0(n3024), .A1(n2144), .B0(n3027), .Y(n3028));
  INVX1   g1973(.A(n3028), .Y(n3029));
  OAI22X1 g1974(.A0(n3021), .A1(n2062), .B0(n2092), .B1(n3029), .Y(n3030));
  AOI21X1 g1975(.A0(n3020), .A1(n2063), .B0(n3030), .Y(n3031));
  OAI21X1 g1976(.A0(n3011), .A1(n2049), .B0(n3031), .Y(n3032));
  NOR2X1  g1977(.A(n3032), .B(n3018), .Y(n3033));
  NAND2X1 g1978(.A(n1998), .B(P1_REG0_REG_20__SCAN_IN), .Y(n3034));
  OAI21X1 g1979(.A0(n3033), .A1(n1998), .B0(n3034), .Y(P1_U3510));
  NOR2X1  g1980(.A(n2003), .B(n1632), .Y(n3036));
  XOR2X1  g1981(.A(n3036), .B(n3029), .Y(n3037));
  INVX1   g1982(.A(n3007), .Y(n3038));
  INVX1   g1983(.A(n2985), .Y(n3039));
  INVX1   g1984(.A(n2986), .Y(n3040));
  OAI21X1 g1985(.A0(n2945), .A1(n3039), .B0(n3040), .Y(n3041));
  AOI21X1 g1986(.A0(n3041), .A1(n3038), .B0(n3008), .Y(n3042));
  XOR2X1  g1987(.A(n3042), .B(n3037), .Y(n3043));
  INVX1   g1988(.A(n3003), .Y(n3044));
  AOI21X1 g1989(.A0(n2941), .A1(n3002), .B0(n2983), .Y(n3045));
  NAND3X1 g1990(.A(n2983), .B(n2941), .C(n3002), .Y(n3046));
  AOI21X1 g1991(.A0(n3046), .A1(n2976), .B0(n3045), .Y(n3047));
  AOI21X1 g1992(.A0(n3044), .A1(n2953), .B0(n3047), .Y(n3048));
  NOR3X1  g1993(.A(n3028), .B(n2003), .C(n1632), .Y(n3049));
  OAI21X1 g1994(.A0(n2003), .A1(n1632), .B0(n3028), .Y(n3050));
  INVX1   g1995(.A(n3050), .Y(n3051));
  NOR3X1  g1996(.A(n3047), .B(n3051), .C(n3049), .Y(n3052));
  OAI21X1 g1997(.A0(n3003), .A1(n2952), .B0(n3052), .Y(n3053));
  OAI21X1 g1998(.A0(n3048), .A1(n3037), .B0(n3053), .Y(n3054));
  OAI22X1 g1999(.A0(n2976), .A1(n2212), .B0(n2211), .B1(n3054), .Y(n3055));
  AOI21X1 g2000(.A0(n2232), .A1(n2231), .B0(n3054), .Y(n3056));
  NOR2X1  g2001(.A(n3056), .B(n3055), .Y(n3057));
  OAI21X1 g2002(.A0(n3043), .A1(n2177), .B0(n3057), .Y(n3058));
  NOR2X1  g2003(.A(n3043), .B(n2192), .Y(n3059));
  AOI21X1 g2004(.A0(n2176), .A1(n2030), .B0(n3043), .Y(n3060));
  NAND3X1 g2005(.A(n3021), .B(n2966), .C(n2964), .Y(n3061));
  XOR2X1  g2006(.A(n3036), .B(n3061), .Y(n3062));
  INVX1   g2007(.A(n3036), .Y(n3063));
  NOR4X1  g2008(.A(n2969), .B(n3022), .C(n2968), .D(n2927), .Y(n3064));
  XOR2X1  g2009(.A(n3064), .B(P1_REG3_REG_22__SCAN_IN), .Y(n3065));
  INVX1   g2010(.A(n3065), .Y(n3066));
  AOI22X1 g2011(.A0(n2094), .A1(P1_REG0_REG_22__SCAN_IN), .B0(P1_REG2_REG_22__SCAN_IN), .B1(n2095), .Y(n3067));
  INVX1   g2012(.A(n3067), .Y(n3068));
  AOI21X1 g2013(.A0(n2099), .A1(P1_REG1_REG_22__SCAN_IN), .B0(n3068), .Y(n3069));
  OAI21X1 g2014(.A0(n3066), .A1(n2144), .B0(n3069), .Y(n3070));
  INVX1   g2015(.A(n3070), .Y(n3071));
  OAI22X1 g2016(.A0(n3063), .A1(n2062), .B0(n2092), .B1(n3071), .Y(n3072));
  AOI21X1 g2017(.A0(n3062), .A1(n2063), .B0(n3072), .Y(n3073));
  OAI21X1 g2018(.A0(n3054), .A1(n2049), .B0(n3073), .Y(n3074));
  NOR4X1  g2019(.A(n3060), .B(n3059), .C(n3058), .D(n3074), .Y(n3075));
  NAND2X1 g2020(.A(n1998), .B(P1_REG0_REG_21__SCAN_IN), .Y(n3076));
  OAI21X1 g2021(.A0(n3075), .A1(n1998), .B0(n3076), .Y(P1_U3511));
  NOR2X1  g2022(.A(n2003), .B(n1650), .Y(n3078));
  XOR2X1  g2023(.A(n3078), .B(n3071), .Y(n3079));
  INVX1   g2024(.A(n3049), .Y(n3080));
  INVX1   g2025(.A(n3008), .Y(n3081));
  OAI21X1 g2026(.A0(n2996), .A1(n3007), .B0(n3081), .Y(n3082));
  AOI21X1 g2027(.A0(n3082), .A1(n3080), .B0(n3051), .Y(n3083));
  XOR2X1  g2028(.A(n3083), .B(n3079), .Y(n3084));
  INVX1   g2029(.A(n3079), .Y(n3085));
  OAI21X1 g2030(.A0(n2003), .A1(n1632), .B0(n3029), .Y(n3086));
  NAND3X1 g2031(.A(n3086), .B(n3044), .C(n2950), .Y(n3087));
  NOR2X1  g2032(.A(n3087), .B(n2901), .Y(n3088));
  NOR3X1  g2033(.A(n3003), .B(n2907), .C(n2891), .Y(n3089));
  OAI21X1 g2034(.A0(n3089), .A1(n3047), .B0(n3086), .Y(n3090));
  NAND2X1 g2035(.A(n3036), .B(n3028), .Y(n3091));
  NAND2X1 g2036(.A(n3091), .B(n3090), .Y(n3092));
  NOR2X1  g2037(.A(n3092), .B(n3088), .Y(n3093));
  XOR2X1  g2038(.A(n3093), .B(n3085), .Y(n3094));
  OAI22X1 g2039(.A0(n3029), .A1(n2212), .B0(n2211), .B1(n3094), .Y(n3095));
  AOI21X1 g2040(.A0(n2232), .A1(n2231), .B0(n3094), .Y(n3096));
  NOR2X1  g2041(.A(n3096), .B(n3095), .Y(n3097));
  OAI21X1 g2042(.A0(n3084), .A1(n2177), .B0(n3097), .Y(n3098));
  NOR2X1  g2043(.A(n3084), .B(n2192), .Y(n3099));
  AOI21X1 g2044(.A0(n2176), .A1(n2030), .B0(n3084), .Y(n3100));
  NOR3X1  g2045(.A(n3036), .B(n2983), .C(n3019), .Y(n3101));
  INVX1   g2046(.A(n3078), .Y(n3102));
  XOR2X1  g2047(.A(n3102), .B(n3101), .Y(n3103));
  NAND2X1 g2048(.A(n3064), .B(P1_REG3_REG_22__SCAN_IN), .Y(n3104));
  XOR2X1  g2049(.A(n3104), .B(P1_REG3_REG_23__SCAN_IN), .Y(n3105));
  AOI22X1 g2050(.A0(n2094), .A1(P1_REG0_REG_23__SCAN_IN), .B0(P1_REG2_REG_23__SCAN_IN), .B1(n2095), .Y(n3106));
  INVX1   g2051(.A(n3106), .Y(n3107));
  AOI21X1 g2052(.A0(n2099), .A1(P1_REG1_REG_23__SCAN_IN), .B0(n3107), .Y(n3108));
  OAI21X1 g2053(.A0(n3105), .A1(n2144), .B0(n3108), .Y(n3109));
  INVX1   g2054(.A(n3109), .Y(n3110));
  OAI22X1 g2055(.A0(n3102), .A1(n2062), .B0(n2092), .B1(n3110), .Y(n3111));
  AOI21X1 g2056(.A0(n3103), .A1(n2063), .B0(n3111), .Y(n3112));
  OAI21X1 g2057(.A0(n3094), .A1(n2049), .B0(n3112), .Y(n3113));
  NOR4X1  g2058(.A(n3100), .B(n3099), .C(n3098), .D(n3113), .Y(n3114));
  NAND2X1 g2059(.A(n1998), .B(P1_REG0_REG_22__SCAN_IN), .Y(n3115));
  OAI21X1 g2060(.A0(n3114), .A1(n1998), .B0(n3115), .Y(P1_U3512));
  OAI21X1 g2061(.A0(n3078), .A1(n3071), .B0(n3083), .Y(n3117));
  NOR3X1  g2062(.A(n3070), .B(n2003), .C(n1650), .Y(n3118));
  INVX1   g2063(.A(n2003), .Y(n3119));
  OAI21X1 g2064(.A0(n1673), .A1(n1662), .B0(n3119), .Y(n3120));
  XOR2X1  g2065(.A(n3120), .B(n3109), .Y(n3121));
  NOR2X1  g2066(.A(n3121), .B(n3118), .Y(n3122));
  NAND2X1 g2067(.A(n3122), .B(n3117), .Y(n3123));
  NOR2X1  g2068(.A(n3120), .B(n3109), .Y(n3124));
  NOR2X1  g2069(.A(n3078), .B(n3071), .Y(n3125));
  AOI21X1 g2070(.A0(n3120), .A1(n3109), .B0(n3125), .Y(n3126));
  INVX1   g2071(.A(n3126), .Y(n3127));
  NOR2X1  g2072(.A(n3127), .B(n3124), .Y(n3128));
  OAI21X1 g2073(.A0(n3083), .A1(n3118), .B0(n3128), .Y(n3129));
  AOI21X1 g2074(.A0(n3129), .A1(n3123), .B0(n2177), .Y(n3130));
  OAI22X1 g2075(.A0(n3088), .A1(n3092), .B0(n3078), .B1(n3070), .Y(n3131));
  OAI21X1 g2076(.A0(n3102), .A1(n3071), .B0(n3131), .Y(n3132));
  XOR2X1  g2077(.A(n3132), .B(n3121), .Y(n3133));
  OAI22X1 g2078(.A0(n3071), .A1(n2212), .B0(n2211), .B1(n3133), .Y(n3134));
  AOI21X1 g2079(.A0(n2232), .A1(n2231), .B0(n3133), .Y(n3135));
  NOR3X1  g2080(.A(n3135), .B(n3134), .C(n3130), .Y(n3136));
  AOI21X1 g2081(.A0(n3129), .A1(n3123), .B0(n2192), .Y(n3137));
  AOI22X1 g2082(.A0(n3123), .A1(n3129), .B0(n2176), .B1(n2030), .Y(n3138));
  NOR2X1  g2083(.A(n3138), .B(n3137), .Y(n3139));
  NAND2X1 g2084(.A(n3139), .B(n3136), .Y(n3140));
  OAI21X1 g2085(.A0(n2003), .A1(n1650), .B0(n3101), .Y(n3141));
  INVX1   g2086(.A(n3120), .Y(n3142));
  XOR2X1  g2087(.A(n3142), .B(n3141), .Y(n3143));
  NAND3X1 g2088(.A(n3064), .B(P1_REG3_REG_23__SCAN_IN), .C(P1_REG3_REG_22__SCAN_IN), .Y(n3144));
  XOR2X1  g2089(.A(n3144), .B(P1_REG3_REG_24__SCAN_IN), .Y(n3145));
  AOI22X1 g2090(.A0(n2094), .A1(P1_REG0_REG_24__SCAN_IN), .B0(P1_REG2_REG_24__SCAN_IN), .B1(n2095), .Y(n3146));
  INVX1   g2091(.A(n3146), .Y(n3147));
  AOI21X1 g2092(.A0(n2099), .A1(P1_REG1_REG_24__SCAN_IN), .B0(n3147), .Y(n3148));
  OAI21X1 g2093(.A0(n3145), .A1(n2144), .B0(n3148), .Y(n3149));
  INVX1   g2094(.A(n3149), .Y(n3150));
  OAI22X1 g2095(.A0(n3120), .A1(n2062), .B0(n2092), .B1(n3150), .Y(n3151));
  AOI21X1 g2096(.A0(n3143), .A1(n2063), .B0(n3151), .Y(n3152));
  OAI21X1 g2097(.A0(n3133), .A1(n2049), .B0(n3152), .Y(n3153));
  NOR2X1  g2098(.A(n3153), .B(n3140), .Y(n3154));
  NAND2X1 g2099(.A(n1998), .B(P1_REG0_REG_23__SCAN_IN), .Y(n3155));
  OAI21X1 g2100(.A0(n3154), .A1(n1998), .B0(n3155), .Y(P1_U3513));
  NOR2X1  g2101(.A(n2003), .B(n1697), .Y(n3157));
  XOR2X1  g2102(.A(n3157), .B(n3150), .Y(n3158));
  INVX1   g2103(.A(n3124), .Y(n3159));
  OAI21X1 g2104(.A0(n3118), .A1(n3050), .B0(n3126), .Y(n3160));
  NOR3X1  g2105(.A(n3124), .B(n3118), .C(n3049), .Y(n3161));
  AOI22X1 g2106(.A0(n3160), .A1(n3159), .B0(n3082), .B1(n3161), .Y(n3162));
  XOR2X1  g2107(.A(n3162), .B(n3158), .Y(n3163));
  INVX1   g2108(.A(n3163), .Y(n3164));
  NAND2X1 g2109(.A(n3164), .B(n2041), .Y(n3165));
  NOR2X1  g2110(.A(n3120), .B(n3110), .Y(n3166));
  NAND2X1 g2111(.A(n3120), .B(n3110), .Y(n3167));
  AOI21X1 g2112(.A0(n3167), .A1(n3132), .B0(n3166), .Y(n3168));
  NOR3X1  g2113(.A(n3149), .B(n2003), .C(n1697), .Y(n3169));
  NOR2X1  g2114(.A(n3157), .B(n3150), .Y(n3170));
  OAI21X1 g2115(.A0(n3170), .A1(n3169), .B0(n3168), .Y(n3171));
  NAND2X1 g2116(.A(n1719), .B(n1713), .Y(n3172));
  XOR2X1  g2117(.A(n1695), .B(n3172), .Y(n3173));
  NOR2X1  g2118(.A(n3173), .B(n1152), .Y(n3174));
  OAI21X1 g2119(.A0(n3174), .A1(n1688), .B0(n3119), .Y(n3175));
  XOR2X1  g2120(.A(n3175), .B(n3150), .Y(n3176));
  OAI21X1 g2121(.A0(n3176), .A1(n3168), .B0(n3171), .Y(n3177));
  AOI22X1 g2122(.A0(n3109), .A1(n2081), .B0(n2043), .B1(n3177), .Y(n3178));
  OAI21X1 g2123(.A0(n2045), .A1(n2038), .B0(n3177), .Y(n3179));
  NAND3X1 g2124(.A(n3179), .B(n3178), .C(n3165), .Y(n3180));
  NOR2X1  g2125(.A(n3163), .B(n2192), .Y(n3181));
  AOI21X1 g2126(.A0(n2176), .A1(n2030), .B0(n3163), .Y(n3182));
  NAND2X1 g2127(.A(n3177), .B(n2048), .Y(n3183));
  NAND3X1 g2128(.A(n3120), .B(n3102), .C(n3101), .Y(n3184));
  XOR2X1  g2129(.A(n3157), .B(n3184), .Y(n3185));
  NAND4X1 g2130(.A(P1_REG3_REG_23__SCAN_IN), .B(P1_REG3_REG_24__SCAN_IN), .C(P1_REG3_REG_22__SCAN_IN), .D(n3064), .Y(n3186));
  XOR2X1  g2131(.A(n3186), .B(P1_REG3_REG_25__SCAN_IN), .Y(n3187));
  AOI22X1 g2132(.A0(n2094), .A1(P1_REG0_REG_25__SCAN_IN), .B0(P1_REG2_REG_25__SCAN_IN), .B1(n2095), .Y(n3188));
  INVX1   g2133(.A(n3188), .Y(n3189));
  AOI21X1 g2134(.A0(n2099), .A1(P1_REG1_REG_25__SCAN_IN), .B0(n3189), .Y(n3190));
  OAI21X1 g2135(.A0(n3187), .A1(n2144), .B0(n3190), .Y(n3191));
  INVX1   g2136(.A(n3191), .Y(n3192));
  OAI22X1 g2137(.A0(n3175), .A1(n2062), .B0(n2092), .B1(n3192), .Y(n3193));
  AOI21X1 g2138(.A0(n3185), .A1(n2063), .B0(n3193), .Y(n3194));
  NAND2X1 g2139(.A(n3194), .B(n3183), .Y(n3195));
  NOR4X1  g2140(.A(n3182), .B(n3181), .C(n3180), .D(n3195), .Y(n3196));
  NAND2X1 g2141(.A(n1998), .B(P1_REG0_REG_24__SCAN_IN), .Y(n3197));
  OAI21X1 g2142(.A0(n3196), .A1(n1998), .B0(n3197), .Y(P1_U3514));
  NOR2X1  g2143(.A(n2003), .B(n1726), .Y(n3199));
  XOR2X1  g2144(.A(n3199), .B(n3192), .Y(n3200));
  INVX1   g2145(.A(n3169), .Y(n3201));
  NAND2X1 g2146(.A(n3160), .B(n3159), .Y(n3202));
  INVX1   g2147(.A(n3161), .Y(n3203));
  OAI21X1 g2148(.A0(n3203), .A1(n3042), .B0(n3202), .Y(n3204));
  AOI21X1 g2149(.A0(n3204), .A1(n3201), .B0(n3170), .Y(n3205));
  XOR2X1  g2150(.A(n3205), .B(n3200), .Y(n3206));
  INVX1   g2151(.A(n3206), .Y(n3207));
  NAND2X1 g2152(.A(n3207), .B(n2041), .Y(n3208));
  NOR2X1  g2153(.A(n3157), .B(n3149), .Y(n3209));
  NAND2X1 g2154(.A(n3157), .B(n3149), .Y(n3210));
  OAI21X1 g2155(.A0(n3209), .A1(n3168), .B0(n3210), .Y(n3211));
  NAND2X1 g2156(.A(n1737), .B(n1735), .Y(n3212));
  XOR2X1  g2157(.A(n1724), .B(n3212), .Y(n3213));
  NOR2X1  g2158(.A(n3213), .B(n1152), .Y(n3214));
  OAI21X1 g2159(.A0(n3214), .A1(n1710), .B0(n3119), .Y(n3215));
  XOR2X1  g2160(.A(n3215), .B(n3192), .Y(n3216));
  NAND2X1 g2161(.A(n3200), .B(n3211), .Y(n3218));
  OAI21X1 g2162(.A0(n3211), .A1(n3200), .B0(n3218), .Y(n3219));
  AOI22X1 g2163(.A0(n3149), .A1(n2081), .B0(n2043), .B1(n3219), .Y(n3220));
  OAI21X1 g2164(.A0(n2045), .A1(n2038), .B0(n3219), .Y(n3221));
  NAND3X1 g2165(.A(n3221), .B(n3220), .C(n3208), .Y(n3222));
  NOR2X1  g2166(.A(n3206), .B(n2192), .Y(n3223));
  AOI21X1 g2167(.A0(n2176), .A1(n2030), .B0(n3206), .Y(n3224));
  NAND2X1 g2168(.A(n3219), .B(n2048), .Y(n3225));
  NAND4X1 g2169(.A(n3120), .B(n3102), .C(n3101), .D(n3175), .Y(n3226));
  XOR2X1  g2170(.A(n3199), .B(n3226), .Y(n3227));
  INVX1   g2171(.A(P1_REG3_REG_26__SCAN_IN), .Y(n3228));
  INVX1   g2172(.A(P1_REG3_REG_25__SCAN_IN), .Y(n3229));
  NOR2X1  g2173(.A(n3186), .B(n3229), .Y(n3230));
  XOR2X1  g2174(.A(n3230), .B(n3228), .Y(n3231));
  AOI22X1 g2175(.A0(n2094), .A1(P1_REG0_REG_26__SCAN_IN), .B0(P1_REG2_REG_26__SCAN_IN), .B1(n2095), .Y(n3232));
  INVX1   g2176(.A(n3232), .Y(n3233));
  AOI21X1 g2177(.A0(n2099), .A1(P1_REG1_REG_26__SCAN_IN), .B0(n3233), .Y(n3234));
  OAI21X1 g2178(.A0(n3231), .A1(n2144), .B0(n3234), .Y(n3235));
  INVX1   g2179(.A(n3235), .Y(n3236));
  OAI22X1 g2180(.A0(n3215), .A1(n2062), .B0(n2092), .B1(n3236), .Y(n3237));
  AOI21X1 g2181(.A0(n3227), .A1(n2063), .B0(n3237), .Y(n3238));
  NAND2X1 g2182(.A(n3238), .B(n3225), .Y(n3239));
  NOR4X1  g2183(.A(n3224), .B(n3223), .C(n3222), .D(n3239), .Y(n3240));
  NAND2X1 g2184(.A(n1998), .B(P1_REG0_REG_25__SCAN_IN), .Y(n3241));
  OAI21X1 g2185(.A0(n3240), .A1(n1998), .B0(n3241), .Y(P1_U3515));
  NOR2X1  g2186(.A(n2003), .B(n1744), .Y(n3243));
  XOR2X1  g2187(.A(n3243), .B(n3236), .Y(n3244));
  NOR3X1  g2188(.A(n3191), .B(n2003), .C(n1726), .Y(n3245));
  INVX1   g2189(.A(n3245), .Y(n3246));
  NOR2X1  g2190(.A(n3199), .B(n3192), .Y(n3247));
  OAI21X1 g2191(.A0(n3162), .A1(n3169), .B0(n4814), .Y(n3249));
  AOI21X1 g2192(.A0(n3249), .A1(n3246), .B0(n3247), .Y(n3250));
  XOR2X1  g2193(.A(n3250), .B(n3244), .Y(n3251));
  INVX1   g2194(.A(n3251), .Y(n3252));
  NAND2X1 g2195(.A(n3252), .B(n2041), .Y(n3253));
  NOR2X1  g2196(.A(n3209), .B(n3168), .Y(n3254));
  AOI21X1 g2197(.A0(n3157), .A1(n3149), .B0(n3254), .Y(n3255));
  OAI21X1 g2198(.A0(n3215), .A1(n3192), .B0(n3255), .Y(n3256));
  OAI21X1 g2199(.A0(n2003), .A1(n1726), .B0(n3192), .Y(n3257));
  OAI21X1 g2200(.A0(n3243), .A1(n3235), .B0(n3257), .Y(n3258));
  AOI21X1 g2201(.A0(n3243), .A1(n3235), .B0(n3258), .Y(n3259));
  OAI21X1 g2202(.A0(n3215), .A1(n3192), .B0(n3244), .Y(n3260));
  AOI21X1 g2203(.A0(n3257), .A1(n3211), .B0(n3260), .Y(n3261));
  AOI21X1 g2204(.A0(n3259), .A1(n3256), .B0(n3261), .Y(n3262));
  AOI22X1 g2205(.A0(n3191), .A1(n2081), .B0(n2043), .B1(n3262), .Y(n3263));
  OAI21X1 g2206(.A0(n2045), .A1(n2038), .B0(n3262), .Y(n3264));
  NAND3X1 g2207(.A(n3264), .B(n3263), .C(n3253), .Y(n3265));
  NOR2X1  g2208(.A(n3251), .B(n2192), .Y(n3266));
  AOI21X1 g2209(.A0(n2176), .A1(n2030), .B0(n3251), .Y(n3267));
  NAND2X1 g2210(.A(n3262), .B(n2048), .Y(n3268));
  NOR2X1  g2211(.A(n3199), .B(n3226), .Y(n3269));
  NAND2X1 g2212(.A(n1771), .B(n1769), .Y(n3270));
  XOR2X1  g2213(.A(n1742), .B(n3270), .Y(n3271));
  NOR2X1  g2214(.A(n3271), .B(n1152), .Y(n3272));
  OAI21X1 g2215(.A0(n3272), .A1(n1732), .B0(n3119), .Y(n3273));
  XOR2X1  g2216(.A(n3273), .B(n3269), .Y(n3274));
  INVX1   g2217(.A(P1_REG3_REG_27__SCAN_IN), .Y(n3275));
  NOR3X1  g2218(.A(n3186), .B(n3229), .C(n3228), .Y(n3276));
  XOR2X1  g2219(.A(n3276), .B(n3275), .Y(n3277));
  AOI22X1 g2220(.A0(n2094), .A1(P1_REG0_REG_27__SCAN_IN), .B0(P1_REG2_REG_27__SCAN_IN), .B1(n2095), .Y(n3278));
  INVX1   g2221(.A(n3278), .Y(n3279));
  AOI21X1 g2222(.A0(n2099), .A1(P1_REG1_REG_27__SCAN_IN), .B0(n3279), .Y(n3280));
  OAI21X1 g2223(.A0(n3277), .A1(n2144), .B0(n3280), .Y(n3281));
  INVX1   g2224(.A(n3281), .Y(n3282));
  OAI22X1 g2225(.A0(n3273), .A1(n2062), .B0(n2092), .B1(n3282), .Y(n3283));
  AOI21X1 g2226(.A0(n3274), .A1(n2063), .B0(n3283), .Y(n3284));
  NAND2X1 g2227(.A(n3284), .B(n3268), .Y(n3285));
  NOR4X1  g2228(.A(n3267), .B(n3266), .C(n3265), .D(n3285), .Y(n3286));
  NAND2X1 g2229(.A(n1998), .B(P1_REG0_REG_26__SCAN_IN), .Y(n3287));
  OAI21X1 g2230(.A0(n3286), .A1(n1998), .B0(n3287), .Y(P1_U3516));
  AOI22X1 g2231(.A0(n3236), .A1(n3273), .B0(n3215), .B1(n3192), .Y(n3289));
  OAI21X1 g2232(.A0(n3215), .A1(n3192), .B0(n3210), .Y(n3290));
  NAND2X1 g2233(.A(n3290), .B(n3289), .Y(n3291));
  AOI22X1 g2234(.A0(n3243), .A1(n3235), .B0(n3254), .B1(n3289), .Y(n3292));
  NAND2X1 g2235(.A(n3292), .B(n3291), .Y(n3293));
  OAI21X1 g2236(.A0(n1774), .A1(n1758), .B0(n3119), .Y(n3294));
  XOR2X1  g2237(.A(n3294), .B(n3282), .Y(n3295));
  XOR2X1  g2238(.A(n4834), .B(n3293), .Y(n3297));
  INVX1   g2239(.A(n3297), .Y(n3298));
  AOI22X1 g2240(.A0(n3235), .A1(n2081), .B0(n2043), .B1(n3298), .Y(n3299));
  OAI21X1 g2241(.A0(n2045), .A1(n2038), .B0(n3298), .Y(n3300));
  NAND2X1 g2242(.A(n3300), .B(n3299), .Y(n3301));
  NOR2X1  g2243(.A(n3243), .B(n3236), .Y(n3302));
  INVX1   g2244(.A(n3247), .Y(n3303));
  OAI21X1 g2245(.A0(n3205), .A1(n3245), .B0(n3303), .Y(n3304));
  NOR3X1  g2246(.A(n3235), .B(n2003), .C(n1744), .Y(n3305));
  NOR2X1  g2247(.A(n4834), .B(n3305), .Y(n3306));
  OAI21X1 g2248(.A0(n3304), .A1(n3302), .B0(n3306), .Y(n3307));
  NOR2X1  g2249(.A(n3295), .B(n3302), .Y(n3308));
  OAI21X1 g2250(.A0(n3250), .A1(n3305), .B0(n3308), .Y(n3309));
  AOI22X1 g2251(.A0(n3307), .A1(n3309), .B0(n2177), .B1(n2176), .Y(n3310));
  AOI22X1 g2252(.A0(n3307), .A1(n3309), .B0(n2192), .B1(n2030), .Y(n3311));
  NOR3X1  g2253(.A(n3243), .B(n3199), .C(n3226), .Y(n3312));
  XOR2X1  g2254(.A(n3294), .B(n3312), .Y(n3313));
  INVX1   g2255(.A(P1_REG3_REG_28__SCAN_IN), .Y(n3314));
  NOR4X1  g2256(.A(n3275), .B(n3229), .C(n3228), .D(n3186), .Y(n3315));
  XOR2X1  g2257(.A(n3315), .B(n3314), .Y(n3316));
  INVX1   g2258(.A(n3316), .Y(n3317));
  AOI22X1 g2259(.A0(n2094), .A1(P1_REG0_REG_28__SCAN_IN), .B0(P1_REG2_REG_28__SCAN_IN), .B1(n2095), .Y(n3318));
  INVX1   g2260(.A(n3318), .Y(n3319));
  AOI21X1 g2261(.A0(n2099), .A1(P1_REG1_REG_28__SCAN_IN), .B0(n3319), .Y(n3320));
  INVX1   g2262(.A(n3320), .Y(n3321));
  AOI21X1 g2263(.A0(n3317), .A1(n2100), .B0(n3321), .Y(n3322));
  OAI22X1 g2264(.A0(n3294), .A1(n2062), .B0(n2092), .B1(n3322), .Y(n3323));
  AOI21X1 g2265(.A0(n3313), .A1(n2063), .B0(n3323), .Y(n3324));
  OAI21X1 g2266(.A0(n3297), .A1(n2049), .B0(n3324), .Y(n3325));
  NOR4X1  g2267(.A(n3311), .B(n3310), .C(n3301), .D(n3325), .Y(n3326));
  NAND2X1 g2268(.A(n1998), .B(P1_REG0_REG_27__SCAN_IN), .Y(n3327));
  OAI21X1 g2269(.A0(n3326), .A1(n1998), .B0(n3327), .Y(P1_U3517));
  NOR2X1  g2270(.A(n2003), .B(n1790), .Y(n3329));
  XOR2X1  g2271(.A(n3329), .B(n3322), .Y(n3330));
  INVX1   g2272(.A(n3330), .Y(n3331));
  INVX1   g2273(.A(n3305), .Y(n3332));
  NOR2X1  g2274(.A(n2003), .B(n1775), .Y(n3333));
  NAND2X1 g2275(.A(n3333), .B(n3282), .Y(n3334));
  NAND3X1 g2276(.A(n3334), .B(n3304), .C(n3332), .Y(n3335));
  INVX1   g2277(.A(n3302), .Y(n3336));
  AOI21X1 g2278(.A0(n3282), .A1(n3336), .B0(n3333), .Y(n3337));
  NOR3X1  g2279(.A(n3282), .B(n3243), .C(n3236), .Y(n3338));
  NOR2X1  g2280(.A(n3338), .B(n3337), .Y(n3339));
  NAND2X1 g2281(.A(n3339), .B(n3335), .Y(n3340));
  XOR2X1  g2282(.A(n3340), .B(n3331), .Y(n3341));
  NOR2X1  g2283(.A(n3341), .B(n2177), .Y(n3342));
  NOR2X1  g2284(.A(n3333), .B(n3281), .Y(n3343));
  NAND2X1 g2285(.A(n3333), .B(n3281), .Y(n3344));
  OAI21X1 g2286(.A0(n3343), .A1(n3291), .B0(n3344), .Y(n3345));
  NOR3X1  g2287(.A(n3343), .B(n3273), .C(n3236), .Y(n3346));
  NOR4X1  g2288(.A(n3258), .B(n3209), .C(n3168), .D(n3343), .Y(n3347));
  NOR3X1  g2289(.A(n3347), .B(n3346), .C(n3345), .Y(n3348));
  XOR2X1  g2290(.A(n3348), .B(n3331), .Y(n3349));
  INVX1   g2291(.A(n3349), .Y(n3350));
  AOI22X1 g2292(.A0(n3281), .A1(n2081), .B0(n2043), .B1(n3350), .Y(n3351));
  OAI21X1 g2293(.A0(n2045), .A1(n2038), .B0(n3350), .Y(n3352));
  NAND2X1 g2294(.A(n3352), .B(n3351), .Y(n3353));
  XOR2X1  g2295(.A(n3340), .B(n3330), .Y(n3354));
  OAI21X1 g2296(.A0(n2040), .A1(n2029), .B0(n3354), .Y(n3355));
  OAI21X1 g2297(.A0(n3341), .A1(n2192), .B0(n3355), .Y(n3356));
  NOR4X1  g2298(.A(n3243), .B(n3199), .C(n3226), .D(n3333), .Y(n3357));
  INVX1   g2299(.A(n3329), .Y(n3358));
  XOR2X1  g2300(.A(n3358), .B(n3357), .Y(n3359));
  NAND4X1 g2301(.A(n2100), .B(P1_REG3_REG_27__SCAN_IN), .C(P1_REG3_REG_28__SCAN_IN), .D(n3276), .Y(n3360));
  NAND2X1 g2302(.A(n2094), .B(P1_REG0_REG_29__SCAN_IN), .Y(n3361));
  AOI22X1 g2303(.A0(n2095), .A1(P1_REG2_REG_29__SCAN_IN), .B0(P1_REG1_REG_29__SCAN_IN), .B1(n2099), .Y(n3362));
  NAND3X1 g2304(.A(n3362), .B(n3361), .C(n3360), .Y(n3363));
  INVX1   g2305(.A(n3363), .Y(n3364));
  OAI22X1 g2306(.A0(n3358), .A1(n2062), .B0(n2092), .B1(n3364), .Y(n3365));
  AOI21X1 g2307(.A0(n3359), .A1(n2063), .B0(n3365), .Y(n3366));
  OAI21X1 g2308(.A0(n3349), .A1(n2049), .B0(n3366), .Y(n3367));
  NOR4X1  g2309(.A(n3356), .B(n3353), .C(n3342), .D(n3367), .Y(n3368));
  NAND2X1 g2310(.A(n1998), .B(P1_REG0_REG_28__SCAN_IN), .Y(n3369));
  OAI21X1 g2311(.A0(n3368), .A1(n1998), .B0(n3369), .Y(P1_U3518));
  NOR2X1  g2312(.A(n2003), .B(n1820), .Y(n3371));
  XOR2X1  g2313(.A(n3371), .B(n3364), .Y(n3372));
  NOR2X1  g2314(.A(n3348), .B(n3358), .Y(n3373));
  AOI21X1 g2315(.A0(n3348), .A1(n3358), .B0(n3322), .Y(n3374));
  NOR2X1  g2316(.A(n3374), .B(n3373), .Y(n3375));
  XOR2X1  g2317(.A(n3375), .B(n3372), .Y(n3376));
  NAND2X1 g2318(.A(n3376), .B(n2045), .Y(n3377));
  NOR2X1  g2319(.A(n1987), .B(n1982), .Y(n3378));
  NOR3X1  g2320(.A(n2000), .B(n1999), .C(P1_B_REG_SCAN_IN), .Y(n3379));
  OAI21X1 g2321(.A0(n3379), .A1(n2003), .B0(n3378), .Y(n3380));
  NAND3X1 g2322(.A(n2017), .B(n2021), .C(P1_REG1_REG_30__SCAN_IN), .Y(n3381));
  AOI22X1 g2323(.A0(n2094), .A1(P1_REG0_REG_30__SCAN_IN), .B0(P1_REG2_REG_30__SCAN_IN), .B1(n2095), .Y(n3382));
  NAND2X1 g2324(.A(n3382), .B(n3381), .Y(n3383));
  INVX1   g2325(.A(n3383), .Y(n3384));
  OAI22X1 g2326(.A0(n3380), .A1(n3384), .B0(n3322), .B1(n2212), .Y(n3385));
  AOI21X1 g2327(.A0(n3376), .A1(n2038), .B0(n3385), .Y(n3386));
  NAND2X1 g2328(.A(n3386), .B(n3377), .Y(n3387));
  NAND2X1 g2329(.A(n3376), .B(n2048), .Y(n3388));
  INVX1   g2330(.A(n1781), .Y(n3389));
  NAND2X1 g2331(.A(n1813), .B(n1811), .Y(n3390));
  XOR2X1  g2332(.A(n1788), .B(n3390), .Y(n3391));
  OAI21X1 g2333(.A0(n3391), .A1(n1152), .B0(n3389), .Y(n3392));
  AOI21X1 g2334(.A0(n3119), .A1(n3392), .B0(n3322), .Y(n3393));
  INVX1   g2335(.A(n3334), .Y(n3394));
  NOR3X1  g2336(.A(n3394), .B(n3250), .C(n3305), .Y(n3395));
  NOR4X1  g2337(.A(n3337), .B(n3395), .C(n3393), .D(n3338), .Y(n3396));
  INVX1   g2338(.A(n3322), .Y(n3397));
  NAND2X1 g2339(.A(n1842), .B(n1840), .Y(n3398));
  XOR2X1  g2340(.A(n1818), .B(n3398), .Y(n3399));
  NOR2X1  g2341(.A(n3399), .B(n1152), .Y(n3400));
  OAI21X1 g2342(.A0(n3400), .A1(n1808), .B0(n3119), .Y(n3401));
  XOR2X1  g2343(.A(n3401), .B(n3364), .Y(n3402));
  OAI21X1 g2344(.A0(n3358), .A1(n3397), .B0(n3402), .Y(n3403));
  NOR3X1  g2345(.A(n3397), .B(n2003), .C(n1790), .Y(n3404));
  AOI21X1 g2346(.A0(n3339), .A1(n3335), .B0(n3404), .Y(n3405));
  OAI21X1 g2347(.A0(n2003), .A1(n1790), .B0(n3397), .Y(n3406));
  NAND2X1 g2348(.A(n3372), .B(n3406), .Y(n3407));
  OAI22X1 g2349(.A0(n3405), .A1(n3407), .B0(n3403), .B1(n3396), .Y(n3408));
  NAND2X1 g2350(.A(n3408), .B(n2034), .Y(n3409));
  OAI21X1 g2351(.A0(n2003), .A1(n1790), .B0(n3357), .Y(n3410));
  XOR2X1  g2352(.A(n3371), .B(n3410), .Y(n3411));
  AOI22X1 g2353(.A0(n3371), .A1(n2302), .B0(n2063), .B1(n3411), .Y(n3412));
  NAND3X1 g2354(.A(n3412), .B(n3409), .C(n3388), .Y(n3413));
  OAI21X1 g2355(.A0(n2040), .A1(n2029), .B0(n3408), .Y(n3414));
  AOI22X1 g2356(.A0(n3376), .A1(n2043), .B0(n2041), .B1(n3408), .Y(n3415));
  NAND2X1 g2357(.A(n3415), .B(n3414), .Y(n3416));
  NOR3X1  g2358(.A(n3416), .B(n3413), .C(n3387), .Y(n3417));
  NAND2X1 g2359(.A(n1998), .B(P1_REG0_REG_29__SCAN_IN), .Y(n3418));
  OAI21X1 g2360(.A0(n3417), .A1(n1998), .B0(n3418), .Y(P1_U3519));
  NAND3X1 g2361(.A(n3401), .B(n3358), .C(n3357), .Y(n3420));
  NOR2X1  g2362(.A(n2003), .B(n1846), .Y(n3421));
  XOR2X1  g2363(.A(n3421), .B(n3420), .Y(n3422));
  OAI21X1 g2364(.A0(n1845), .A1(n1829), .B0(n3119), .Y(n3423));
  NAND3X1 g2365(.A(n2017), .B(n2021), .C(P1_REG1_REG_31__SCAN_IN), .Y(n3424));
  AOI22X1 g2366(.A0(n2094), .A1(P1_REG0_REG_31__SCAN_IN), .B0(P1_REG2_REG_31__SCAN_IN), .B1(n2095), .Y(n3425));
  AOI21X1 g2367(.A0(n3425), .A1(n3424), .B0(n3380), .Y(n3426));
  INVX1   g2368(.A(n3426), .Y(n3427));
  OAI21X1 g2369(.A0(n3423), .A1(n2062), .B0(n3427), .Y(n3428));
  AOI21X1 g2370(.A0(n3422), .A1(n2063), .B0(n3428), .Y(n3429));
  NAND2X1 g2371(.A(n1998), .B(P1_REG0_REG_30__SCAN_IN), .Y(n3430));
  OAI21X1 g2372(.A0(n3429), .A1(n1998), .B0(n3430), .Y(P1_U3520));
  NOR2X1  g2373(.A(n3421), .B(n3420), .Y(n3432));
  OAI21X1 g2374(.A0(n1866), .A1(n1851), .B0(n3119), .Y(n3433));
  XOR2X1  g2375(.A(n3433), .B(n3432), .Y(n3434));
  OAI21X1 g2376(.A0(n3433), .A1(n2062), .B0(n3427), .Y(n3435));
  AOI21X1 g2377(.A0(n3434), .A1(n2063), .B0(n3435), .Y(n3436));
  NAND2X1 g2378(.A(n1998), .B(P1_REG0_REG_31__SCAN_IN), .Y(n3437));
  OAI21X1 g2379(.A0(n3436), .A1(n1998), .B0(n3437), .Y(P1_U3521));
  INVX1   g2380(.A(n1997), .Y(n3439));
  NAND3X1 g2381(.A(n3439), .B(n1995), .C(n1891), .Y(n3440));
  NAND2X1 g2382(.A(n3440), .B(P1_REG1_REG_0__SCAN_IN), .Y(n3441));
  OAI21X1 g2383(.A0(n3440), .A1(n2068), .B0(n3441), .Y(P1_U3522));
  NAND2X1 g2384(.A(n3440), .B(P1_REG1_REG_1__SCAN_IN), .Y(n3443));
  OAI21X1 g2385(.A0(n3440), .A1(n2107), .B0(n3443), .Y(P1_U3523));
  NAND2X1 g2386(.A(n3440), .B(P1_REG1_REG_2__SCAN_IN), .Y(n3445));
  OAI21X1 g2387(.A0(n3440), .A1(n2150), .B0(n3445), .Y(P1_U3524));
  NAND2X1 g2388(.A(n3440), .B(P1_REG1_REG_3__SCAN_IN), .Y(n3447));
  OAI21X1 g2389(.A0(n3440), .A1(n2208), .B0(n3447), .Y(P1_U3525));
  NAND2X1 g2390(.A(n3440), .B(P1_REG1_REG_4__SCAN_IN), .Y(n3449));
  OAI21X1 g2391(.A0(n3440), .A1(n2261), .B0(n3449), .Y(P1_U3526));
  NAND2X1 g2392(.A(n3440), .B(P1_REG1_REG_5__SCAN_IN), .Y(n3451));
  OAI21X1 g2393(.A0(n3440), .A1(n2316), .B0(n3451), .Y(P1_U3527));
  NAND2X1 g2394(.A(n3440), .B(P1_REG1_REG_6__SCAN_IN), .Y(n3453));
  OAI21X1 g2395(.A0(n3440), .A1(n2367), .B0(n3453), .Y(P1_U3528));
  NAND2X1 g2396(.A(n3440), .B(P1_REG1_REG_7__SCAN_IN), .Y(n3455));
  OAI21X1 g2397(.A0(n3440), .A1(n2413), .B0(n3455), .Y(P1_U3529));
  NAND2X1 g2398(.A(n3440), .B(P1_REG1_REG_8__SCAN_IN), .Y(n3457));
  OAI21X1 g2399(.A0(n3440), .A1(n2462), .B0(n3457), .Y(P1_U3530));
  NAND2X1 g2400(.A(n3440), .B(P1_REG1_REG_9__SCAN_IN), .Y(n3459));
  OAI21X1 g2401(.A0(n3440), .A1(n2508), .B0(n3459), .Y(P1_U3531));
  NAND2X1 g2402(.A(n3440), .B(P1_REG1_REG_10__SCAN_IN), .Y(n3461));
  OAI21X1 g2403(.A0(n3440), .A1(n2553), .B0(n3461), .Y(P1_U3532));
  NAND2X1 g2404(.A(n3440), .B(P1_REG1_REG_11__SCAN_IN), .Y(n3463));
  OAI21X1 g2405(.A0(n3440), .A1(n2606), .B0(n3463), .Y(P1_U3533));
  NAND2X1 g2406(.A(n3440), .B(P1_REG1_REG_12__SCAN_IN), .Y(n3465));
  OAI21X1 g2407(.A0(n3440), .A1(n2654), .B0(n3465), .Y(P1_U3534));
  NAND2X1 g2408(.A(n3440), .B(P1_REG1_REG_13__SCAN_IN), .Y(n3467));
  OAI21X1 g2409(.A0(n3440), .A1(n2706), .B0(n3467), .Y(P1_U3535));
  NAND2X1 g2410(.A(n3440), .B(P1_REG1_REG_14__SCAN_IN), .Y(n3469));
  OAI21X1 g2411(.A0(n3440), .A1(n2752), .B0(n3469), .Y(P1_U3536));
  NAND2X1 g2412(.A(n3440), .B(P1_REG1_REG_15__SCAN_IN), .Y(n3471));
  OAI21X1 g2413(.A0(n3440), .A1(n2795), .B0(n3471), .Y(P1_U3537));
  NAND2X1 g2414(.A(n3440), .B(P1_REG1_REG_16__SCAN_IN), .Y(n3473));
  OAI21X1 g2415(.A0(n3440), .A1(n2845), .B0(n3473), .Y(P1_U3538));
  NAND2X1 g2416(.A(n3440), .B(P1_REG1_REG_17__SCAN_IN), .Y(n3475));
  OAI21X1 g2417(.A0(n3440), .A1(n2895), .B0(n3475), .Y(P1_U3539));
  NAND2X1 g2418(.A(n3440), .B(P1_REG1_REG_18__SCAN_IN), .Y(n3477));
  OAI21X1 g2419(.A0(n3440), .A1(n2937), .B0(n3477), .Y(P1_U3540));
  NAND2X1 g2420(.A(n3440), .B(P1_REG1_REG_19__SCAN_IN), .Y(n3479));
  OAI21X1 g2421(.A0(n3440), .A1(n2980), .B0(n3479), .Y(P1_U3541));
  NAND2X1 g2422(.A(n3440), .B(P1_REG1_REG_20__SCAN_IN), .Y(n3481));
  OAI21X1 g2423(.A0(n3440), .A1(n3033), .B0(n3481), .Y(P1_U3542));
  NAND2X1 g2424(.A(n3440), .B(P1_REG1_REG_21__SCAN_IN), .Y(n3483));
  OAI21X1 g2425(.A0(n3440), .A1(n3075), .B0(n3483), .Y(P1_U3543));
  NAND2X1 g2426(.A(n3440), .B(P1_REG1_REG_22__SCAN_IN), .Y(n3485));
  OAI21X1 g2427(.A0(n3440), .A1(n3114), .B0(n3485), .Y(P1_U3544));
  NAND2X1 g2428(.A(n3440), .B(P1_REG1_REG_23__SCAN_IN), .Y(n3487));
  OAI21X1 g2429(.A0(n3440), .A1(n3154), .B0(n3487), .Y(P1_U3545));
  NAND2X1 g2430(.A(n3440), .B(P1_REG1_REG_24__SCAN_IN), .Y(n3489));
  OAI21X1 g2431(.A0(n3440), .A1(n3196), .B0(n3489), .Y(P1_U3546));
  NAND2X1 g2432(.A(n3440), .B(P1_REG1_REG_25__SCAN_IN), .Y(n3491));
  OAI21X1 g2433(.A0(n3440), .A1(n3240), .B0(n3491), .Y(P1_U3547));
  NAND2X1 g2434(.A(n3440), .B(P1_REG1_REG_26__SCAN_IN), .Y(n3493));
  OAI21X1 g2435(.A0(n3440), .A1(n3286), .B0(n3493), .Y(P1_U3548));
  NAND2X1 g2436(.A(n3440), .B(P1_REG1_REG_27__SCAN_IN), .Y(n3495));
  OAI21X1 g2437(.A0(n3440), .A1(n3326), .B0(n3495), .Y(P1_U3549));
  NAND2X1 g2438(.A(n3440), .B(P1_REG1_REG_28__SCAN_IN), .Y(n3497));
  OAI21X1 g2439(.A0(n3440), .A1(n3368), .B0(n3497), .Y(P1_U3550));
  NAND2X1 g2440(.A(n3440), .B(P1_REG1_REG_29__SCAN_IN), .Y(n3499));
  OAI21X1 g2441(.A0(n3440), .A1(n3417), .B0(n3499), .Y(P1_U3551));
  NAND2X1 g2442(.A(n3440), .B(P1_REG1_REG_30__SCAN_IN), .Y(n3501));
  OAI21X1 g2443(.A0(n3440), .A1(n3429), .B0(n3501), .Y(P1_U3552));
  NAND2X1 g2444(.A(n3440), .B(P1_REG1_REG_31__SCAN_IN), .Y(n3503));
  OAI21X1 g2445(.A0(n3440), .A1(n3436), .B0(n3503), .Y(P1_U3553));
  NOR4X1  g2446(.A(n1989), .B(n2028), .C(n1983), .D(n1991), .Y(n3505));
  INVX1   g2447(.A(n3505), .Y(n3506));
  INVX1   g2448(.A(n1980), .Y(n3507));
  INVX1   g2449(.A(n3378), .Y(n3508));
  AOI21X1 g2450(.A0(n1991), .A1(n1985), .B0(n3508), .Y(n3509));
  INVX1   g2451(.A(n3509), .Y(n3510));
  NAND4X1 g2452(.A(n1997), .B(n3507), .C(n1977), .D(n3510), .Y(n3511));
  NAND2X1 g2453(.A(n3511), .B(n3506), .Y(n3512));
  NAND4X1 g2454(.A(n2058), .B(n2050), .C(n1891), .D(n3512), .Y(n3513));
  NAND2X1 g2455(.A(n3512), .B(n1891), .Y(n3514));
  INVX1   g2456(.A(n3514), .Y(n3515));
  AOI21X1 g2457(.A0(n3512), .A1(n1891), .B0(n2019), .Y(n3516));
  AOI21X1 g2458(.A0(n3515), .A1(n2047), .B0(n3516), .Y(n3517));
  NAND3X1 g2459(.A(n1987), .B(n2028), .C(n1982), .Y(n3518));
  NOR2X1  g2460(.A(n3518), .B(n3514), .Y(n3519));
  NOR4X1  g2461(.A(n1991), .B(n1987), .C(n2028), .D(n3514), .Y(n3520));
  AOI22X1 g2462(.A0(n3519), .A1(n2010), .B0(n4841), .B1(n3520), .Y(n3521));
  NOR4X1  g2463(.A(n1989), .B(n2028), .C(n1983), .D(n2037), .Y(n3522));
  INVX1   g2464(.A(n3522), .Y(n3523));
  NOR2X1  g2465(.A(n3523), .B(n3514), .Y(n3524));
  NOR2X1  g2466(.A(n3514), .B(n3506), .Y(n3525));
  AOI22X1 g2467(.A0(n3524), .A1(n2010), .B0(P1_REG3_REG_0__SCAN_IN), .B1(n3525), .Y(n3526));
  NAND4X1 g2468(.A(n3521), .B(n3517), .C(n3513), .D(n3526), .Y(P1_U3293));
  NAND4X1 g2469(.A(n2102), .B(n2050), .C(n1891), .D(n3512), .Y(n3528));
  AOI21X1 g2470(.A0(n3512), .A1(n1891), .B0(n2051), .Y(n3529));
  AOI21X1 g2471(.A0(n3515), .A1(n2090), .B0(n3529), .Y(n3530));
  AOI22X1 g2472(.A0(n3519), .A1(n2075), .B0(n2079), .B1(n3520), .Y(n3531));
  AOI22X1 g2473(.A0(n3524), .A1(n2091), .B0(P1_REG3_REG_1__SCAN_IN), .B1(n3525), .Y(n3532));
  NAND4X1 g2474(.A(n3531), .B(n3530), .C(n3528), .D(n3532), .Y(P1_U3292));
  NAND4X1 g2475(.A(n2160), .B(n2050), .C(n1891), .D(n3512), .Y(n3534));
  AOI22X1 g2476(.A0(n3519), .A1(n2114), .B0(n2139), .B1(n3524), .Y(n3535));
  INVX1   g2477(.A(P1_REG2_REG_2__SCAN_IN), .Y(n3536));
  AOI21X1 g2478(.A0(n3512), .A1(n1891), .B0(n3536), .Y(n3537));
  AOI21X1 g2479(.A0(n3515), .A1(n2135), .B0(n3537), .Y(n3538));
  AOI22X1 g2480(.A0(n3520), .A1(n2124), .B0(P1_REG3_REG_2__SCAN_IN), .B1(n3525), .Y(n3539));
  NAND4X1 g2481(.A(n3538), .B(n3535), .C(n3534), .D(n3539), .Y(P1_U3291));
  AOI22X1 g2482(.A0(n3520), .A1(n2173), .B0(n2158), .B1(n3525), .Y(n3541));
  AOI22X1 g2483(.A0(n3519), .A1(n2169), .B0(n2197), .B1(n3524), .Y(n3542));
  INVX1   g2484(.A(P1_REG2_REG_3__SCAN_IN), .Y(n3543));
  NOR2X1  g2485(.A(n3514), .B(n2092), .Y(n3544));
  INVX1   g2486(.A(n3544), .Y(n3545));
  OAI22X1 g2487(.A0(n3515), .A1(n3543), .B0(n2204), .B1(n3545), .Y(n3546));
  AOI21X1 g2488(.A0(n3515), .A1(n2195), .B0(n3546), .Y(n3547));
  NAND3X1 g2489(.A(n3547), .B(n3542), .C(n3541), .Y(P1_U3290));
  NOR3X1  g2490(.A(n2244), .B(n2233), .C(n2230), .Y(n3549));
  INVX1   g2491(.A(P1_REG2_REG_4__SCAN_IN), .Y(n3550));
  INVX1   g2492(.A(n3519), .Y(n3551));
  OAI22X1 g2493(.A0(n3515), .A1(n3550), .B0(n2225), .B1(n3551), .Y(n3552));
  NAND4X1 g2494(.A(n3512), .B(n2246), .C(n1891), .D(n3522), .Y(n3553));
  OAI21X1 g2495(.A0(n3545), .A1(n2257), .B0(n3553), .Y(n3554));
  INVX1   g2496(.A(n3520), .Y(n3555));
  INVX1   g2497(.A(n3525), .Y(n3556));
  OAI22X1 g2498(.A0(n3555), .A1(n2229), .B0(n2202), .B1(n3556), .Y(n3557));
  NOR3X1  g2499(.A(n3557), .B(n3554), .C(n3552), .Y(n3558));
  OAI21X1 g2500(.A0(n3514), .A1(n3549), .B0(n3558), .Y(P1_U3289));
  OAI21X1 g2501(.A0(n2297), .A1(n2295), .B0(n3515), .Y(n3560));
  OAI22X1 g2502(.A0(n3515), .A1(n2247), .B0(n2283), .B1(n3551), .Y(n3561));
  INVX1   g2503(.A(n3524), .Y(n3562));
  OAI22X1 g2504(.A0(n3545), .A1(n2312), .B0(n2301), .B1(n3562), .Y(n3563));
  OAI22X1 g2505(.A0(n3555), .A1(n2298), .B0(n2253), .B1(n3556), .Y(n3564));
  NOR3X1  g2506(.A(n3564), .B(n3563), .C(n3561), .Y(n3565));
  NAND2X1 g2507(.A(n3565), .B(n3560), .Y(P1_U3288));
  NAND2X1 g2508(.A(n3515), .B(n2353), .Y(n3567));
  AOI22X1 g2509(.A0(n3514), .A1(P1_REG2_REG_6__SCAN_IN), .B0(n2324), .B1(n3519), .Y(n3568));
  AOI22X1 g2510(.A0(n3544), .A1(n2362), .B0(n2356), .B1(n3524), .Y(n3569));
  AOI22X1 g2511(.A0(n3520), .A1(n2346), .B0(n2309), .B1(n3525), .Y(n3570));
  NAND4X1 g2512(.A(n3569), .B(n3568), .C(n3567), .D(n3570), .Y(P1_U3287));
  NOR3X1  g2513(.A(n2396), .B(n2392), .C(n2384), .Y(n3572));
  AOI22X1 g2514(.A0(n3544), .A1(n2408), .B0(n2398), .B1(n3524), .Y(n3573));
  OAI21X1 g2515(.A0(n3556), .A1(n2359), .B0(n3573), .Y(n3574));
  AOI22X1 g2516(.A0(n3514), .A1(P1_REG2_REG_7__SCAN_IN), .B0(n2376), .B1(n3519), .Y(n3575));
  OAI21X1 g2517(.A0(n3555), .A1(n2383), .B0(n3575), .Y(n3576));
  NOR2X1  g2518(.A(n3576), .B(n3574), .Y(n3577));
  OAI21X1 g2519(.A0(n3514), .A1(n3572), .B0(n3577), .Y(P1_U3286));
  NOR3X1  g2520(.A(n2445), .B(n2441), .C(n2430), .Y(n3579));
  NOR2X1  g2521(.A(n3555), .B(n2429), .Y(n3580));
  AOI22X1 g2522(.A0(n3514), .A1(P1_REG2_REG_8__SCAN_IN), .B0(n2424), .B1(n3519), .Y(n3581));
  NAND4X1 g2523(.A(n3505), .B(n2406), .C(n1891), .D(n3512), .Y(n3582));
  AOI22X1 g2524(.A0(n3544), .A1(n2457), .B0(n2448), .B1(n3524), .Y(n3583));
  NAND3X1 g2525(.A(n3583), .B(n3582), .C(n3581), .Y(n3584));
  NOR2X1  g2526(.A(n3584), .B(n3580), .Y(n3585));
  OAI21X1 g2527(.A0(n3514), .A1(n3579), .B0(n3585), .Y(P1_U3285));
  NOR3X1  g2528(.A(n2493), .B(n2490), .C(n2481), .Y(n3587));
  AOI22X1 g2529(.A0(n3514), .A1(P1_REG2_REG_9__SCAN_IN), .B0(n2469), .B1(n3519), .Y(n3588));
  INVX1   g2530(.A(n2451), .Y(n3589));
  NAND4X1 g2531(.A(n3505), .B(n3589), .C(n1891), .D(n3512), .Y(n3590));
  AOI22X1 g2532(.A0(n3544), .A1(n2503), .B0(n2495), .B1(n3524), .Y(n3591));
  NAND3X1 g2533(.A(n3591), .B(n3590), .C(n3588), .Y(n3592));
  AOI21X1 g2534(.A0(n3520), .A1(n2491), .B0(n3592), .Y(n3593));
  OAI21X1 g2535(.A0(n3514), .A1(n3587), .B0(n3593), .Y(P1_U3284));
  NOR3X1  g2536(.A(n2537), .B(n2533), .C(n2527), .Y(n3595));
  NAND4X1 g2537(.A(n3512), .B(n2541), .C(n1891), .D(n3522), .Y(n3596));
  AOI22X1 g2538(.A0(n3514), .A1(P1_REG2_REG_10__SCAN_IN), .B0(n2516), .B1(n3519), .Y(n3597));
  AOI22X1 g2539(.A0(n3544), .A1(n2580), .B0(n2500), .B1(n3525), .Y(n3598));
  NAND3X1 g2540(.A(n3598), .B(n3597), .C(n3596), .Y(n3599));
  AOI21X1 g2541(.A0(n3520), .A1(n2525), .B0(n3599), .Y(n3600));
  OAI21X1 g2542(.A0(n3514), .A1(n3595), .B0(n3600), .Y(P1_U3283));
  NOR2X1  g2543(.A(n3555), .B(n2583), .Y(n3602));
  NAND4X1 g2544(.A(n3512), .B(n2594), .C(n1891), .D(n3522), .Y(n3603));
  AOI22X1 g2545(.A0(n3514), .A1(P1_REG2_REG_11__SCAN_IN), .B0(n2634), .B1(n3544), .Y(n3604));
  INVX1   g2546(.A(n2543), .Y(n3605));
  AOI22X1 g2547(.A0(n3519), .A1(n2562), .B0(n3605), .B1(n3525), .Y(n3606));
  NAND3X1 g2548(.A(n3606), .B(n3604), .C(n3603), .Y(n3607));
  NOR2X1  g2549(.A(n3607), .B(n3602), .Y(n3608));
  OAI21X1 g2550(.A0(n3514), .A1(n2591), .B0(n3608), .Y(P1_U3282));
  NOR3X1  g2551(.A(n2640), .B(n2639), .C(n2628), .Y(n3610));
  NOR2X1  g2552(.A(n3555), .B(n2637), .Y(n3611));
  NAND4X1 g2553(.A(n3512), .B(n2643), .C(n1891), .D(n3522), .Y(n3612));
  AOI22X1 g2554(.A0(n3514), .A1(P1_REG2_REG_12__SCAN_IN), .B0(n2649), .B1(n3544), .Y(n3613));
  INVX1   g2555(.A(n2596), .Y(n3614));
  AOI22X1 g2556(.A0(n3519), .A1(n2614), .B0(n3614), .B1(n3525), .Y(n3615));
  NAND3X1 g2557(.A(n3615), .B(n3613), .C(n3612), .Y(n3616));
  NOR2X1  g2558(.A(n3616), .B(n3611), .Y(n3617));
  OAI21X1 g2559(.A0(n3514), .A1(n3610), .B0(n3617), .Y(P1_U3281));
  NOR3X1  g2560(.A(n2690), .B(n2686), .C(n2677), .Y(n3619));
  NAND2X1 g2561(.A(n3524), .B(n2693), .Y(n3620));
  AOI22X1 g2562(.A0(n3514), .A1(P1_REG2_REG_13__SCAN_IN), .B0(n2709), .B1(n3544), .Y(n3621));
  AOI22X1 g2563(.A0(n3519), .A1(n2665), .B0(n2646), .B1(n3525), .Y(n3622));
  NAND3X1 g2564(.A(n3622), .B(n3621), .C(n3620), .Y(n3623));
  AOI21X1 g2565(.A0(n3520), .A1(n2675), .B0(n3623), .Y(n3624));
  OAI21X1 g2566(.A0(n3514), .A1(n3619), .B0(n3624), .Y(P1_U3280));
  NOR2X1  g2567(.A(n3555), .B(n2726), .Y(n3626));
  NOR2X1  g2568(.A(n3562), .B(n2740), .Y(n3627));
  INVX1   g2569(.A(P1_REG2_REG_14__SCAN_IN), .Y(n3628));
  OAI22X1 g2570(.A0(n3515), .A1(n3628), .B0(n2714), .B1(n3551), .Y(n3629));
  OAI22X1 g2571(.A0(n3545), .A1(n2798), .B0(n2697), .B1(n3556), .Y(n3630));
  NOR4X1  g2572(.A(n3629), .B(n3627), .C(n3626), .D(n3630), .Y(n3631));
  OAI21X1 g2573(.A0(n3514), .A1(n2735), .B0(n3631), .Y(P1_U3279));
  INVX1   g2574(.A(P1_REG2_REG_15__SCAN_IN), .Y(n3633));
  OAI22X1 g2575(.A0(n3515), .A1(n3633), .B0(n2759), .B1(n3551), .Y(n3634));
  OAI22X1 g2576(.A0(n3545), .A1(n2791), .B0(n2744), .B1(n3556), .Y(n3635));
  NOR2X1  g2577(.A(n3635), .B(n3634), .Y(n3636));
  OAI21X1 g2578(.A0(n3562), .A1(n2784), .B0(n3636), .Y(n3637));
  AOI21X1 g2579(.A0(n3520), .A1(n2773), .B0(n3637), .Y(n3638));
  OAI21X1 g2580(.A0(n3514), .A1(n2781), .B0(n3638), .Y(P1_U3278));
  NAND2X1 g2581(.A(n3524), .B(n2833), .Y(n3640));
  AOI22X1 g2582(.A0(n3514), .A1(P1_REG2_REG_16__SCAN_IN), .B0(n2811), .B1(n3519), .Y(n3641));
  AOI22X1 g2583(.A0(n3544), .A1(n2840), .B0(n2787), .B1(n3525), .Y(n3642));
  NAND3X1 g2584(.A(n3642), .B(n3641), .C(n3640), .Y(n3643));
  AOI21X1 g2585(.A0(n3520), .A1(n2824), .B0(n3643), .Y(n3644));
  OAI21X1 g2586(.A0(n3514), .A1(n2830), .B0(n3644), .Y(P1_U3277));
  NAND2X1 g2587(.A(n3515), .B(n2882), .Y(n3646));
  NAND2X1 g2588(.A(n3520), .B(n2866), .Y(n3647));
  NAND2X1 g2589(.A(n3524), .B(n2884), .Y(n3648));
  AOI22X1 g2590(.A0(n3514), .A1(P1_REG2_REG_17__SCAN_IN), .B0(n2836), .B1(n3525), .Y(n3649));
  OAI21X1 g2591(.A0(n3545), .A1(n2891), .B0(n3649), .Y(n3650));
  AOI21X1 g2592(.A0(n3519), .A1(n2854), .B0(n3650), .Y(n3651));
  NAND4X1 g2593(.A(n3648), .B(n3647), .C(n3646), .D(n3651), .Y(P1_U3276));
  NAND2X1 g2594(.A(n3515), .B(n2923), .Y(n3653));
  NAND2X1 g2595(.A(n3520), .B(n2913), .Y(n3654));
  NAND2X1 g2596(.A(n3524), .B(n2926), .Y(n3655));
  AOI22X1 g2597(.A0(n3514), .A1(P1_REG2_REG_18__SCAN_IN), .B0(n2887), .B1(n3525), .Y(n3656));
  OAI21X1 g2598(.A0(n3545), .A1(n2933), .B0(n3656), .Y(n3657));
  AOI21X1 g2599(.A0(n3519), .A1(n2925), .B0(n3657), .Y(n3658));
  NAND4X1 g2600(.A(n3655), .B(n3654), .C(n3653), .D(n3658), .Y(P1_U3275));
  NAND2X1 g2601(.A(n3515), .B(n2963), .Y(n3660));
  INVX1   g2602(.A(n2956), .Y(n3661));
  NAND2X1 g2603(.A(n3520), .B(n3661), .Y(n3662));
  NAND2X1 g2604(.A(n3524), .B(n2967), .Y(n3663));
  AOI22X1 g2605(.A0(n3514), .A1(P1_REG2_REG_19__SCAN_IN), .B0(n2929), .B1(n3525), .Y(n3664));
  OAI21X1 g2606(.A0(n3545), .A1(n2976), .B0(n3664), .Y(n3665));
  AOI21X1 g2607(.A0(n3519), .A1(n2941), .B0(n3665), .Y(n3666));
  NAND4X1 g2608(.A(n3663), .B(n3662), .C(n3660), .D(n3666), .Y(P1_U3274));
  NAND2X1 g2609(.A(n3515), .B(n3018), .Y(n3668));
  NAND3X1 g2610(.A(n3520), .B(n3010), .C(n3005), .Y(n3669));
  NAND2X1 g2611(.A(n3524), .B(n3020), .Y(n3670));
  AOI22X1 g2612(.A0(n3514), .A1(P1_REG2_REG_20__SCAN_IN), .B0(n3028), .B1(n3544), .Y(n3671));
  OAI21X1 g2613(.A0(n3556), .A1(n2971), .B0(n3671), .Y(n3672));
  AOI21X1 g2614(.A0(n3519), .A1(n2983), .B0(n3672), .Y(n3673));
  NAND4X1 g2615(.A(n3670), .B(n3669), .C(n3668), .D(n3673), .Y(P1_U3273));
  NOR3X1  g2616(.A(n3060), .B(n3059), .C(n3058), .Y(n3675));
  NOR2X1  g2617(.A(n3555), .B(n3054), .Y(n3676));
  NAND2X1 g2618(.A(n3524), .B(n3062), .Y(n3677));
  INVX1   g2619(.A(n3024), .Y(n3678));
  AOI22X1 g2620(.A0(n3514), .A1(P1_REG2_REG_21__SCAN_IN), .B0(n3678), .B1(n3525), .Y(n3679));
  OAI21X1 g2621(.A0(n3545), .A1(n3071), .B0(n3679), .Y(n3680));
  AOI21X1 g2622(.A0(n3519), .A1(n3036), .B0(n3680), .Y(n3681));
  NAND2X1 g2623(.A(n3681), .B(n3677), .Y(n3682));
  NOR2X1  g2624(.A(n3682), .B(n3676), .Y(n3683));
  OAI21X1 g2625(.A0(n3514), .A1(n3675), .B0(n3683), .Y(P1_U3272));
  NOR3X1  g2626(.A(n3100), .B(n3099), .C(n3098), .Y(n3685));
  NOR2X1  g2627(.A(n3555), .B(n3094), .Y(n3686));
  NAND2X1 g2628(.A(n3524), .B(n3103), .Y(n3687));
  AOI22X1 g2629(.A0(n3514), .A1(P1_REG2_REG_22__SCAN_IN), .B0(n3109), .B1(n3544), .Y(n3688));
  OAI21X1 g2630(.A0(n3556), .A1(n3066), .B0(n3688), .Y(n3689));
  AOI21X1 g2631(.A0(n3519), .A1(n3078), .B0(n3689), .Y(n3690));
  NAND2X1 g2632(.A(n3690), .B(n3687), .Y(n3691));
  NOR2X1  g2633(.A(n3691), .B(n3686), .Y(n3692));
  OAI21X1 g2634(.A0(n3514), .A1(n3685), .B0(n3692), .Y(P1_U3271));
  NAND2X1 g2635(.A(n3515), .B(n3140), .Y(n3694));
  INVX1   g2636(.A(n3133), .Y(n3695));
  NAND2X1 g2637(.A(n3520), .B(n3695), .Y(n3696));
  NAND2X1 g2638(.A(n3524), .B(n3143), .Y(n3697));
  AOI22X1 g2639(.A0(n3514), .A1(P1_REG2_REG_23__SCAN_IN), .B0(n3149), .B1(n3544), .Y(n3698));
  OAI21X1 g2640(.A0(n3556), .A1(n3105), .B0(n3698), .Y(n3699));
  AOI21X1 g2641(.A0(n3519), .A1(n3142), .B0(n3699), .Y(n3700));
  NAND4X1 g2642(.A(n3697), .B(n3696), .C(n3694), .D(n3700), .Y(P1_U3270));
  NOR3X1  g2643(.A(n3182), .B(n3181), .C(n3180), .Y(n3702));
  NAND2X1 g2644(.A(n3524), .B(n3185), .Y(n3703));
  INVX1   g2645(.A(n3145), .Y(n3704));
  AOI22X1 g2646(.A0(n3514), .A1(P1_REG2_REG_24__SCAN_IN), .B0(n3704), .B1(n3525), .Y(n3705));
  OAI21X1 g2647(.A0(n3545), .A1(n3192), .B0(n3705), .Y(n3706));
  AOI21X1 g2648(.A0(n3519), .A1(n3157), .B0(n3706), .Y(n3707));
  NAND2X1 g2649(.A(n3707), .B(n3703), .Y(n3708));
  AOI21X1 g2650(.A0(n3520), .A1(n3177), .B0(n3708), .Y(n3709));
  OAI21X1 g2651(.A0(n3514), .A1(n3702), .B0(n3709), .Y(P1_U3269));
  NOR3X1  g2652(.A(n3224), .B(n3223), .C(n3222), .Y(n3711));
  NAND2X1 g2653(.A(n3524), .B(n3227), .Y(n3712));
  INVX1   g2654(.A(n3187), .Y(n3713));
  AOI22X1 g2655(.A0(n3514), .A1(P1_REG2_REG_25__SCAN_IN), .B0(n3713), .B1(n3525), .Y(n3714));
  OAI21X1 g2656(.A0(n3545), .A1(n3236), .B0(n3714), .Y(n3715));
  AOI21X1 g2657(.A0(n3519), .A1(n3199), .B0(n3715), .Y(n3716));
  NAND2X1 g2658(.A(n3716), .B(n3712), .Y(n3717));
  AOI21X1 g2659(.A0(n3520), .A1(n3219), .B0(n3717), .Y(n3718));
  OAI21X1 g2660(.A0(n3514), .A1(n3711), .B0(n3718), .Y(P1_U3268));
  NOR3X1  g2661(.A(n3267), .B(n3266), .C(n3265), .Y(n3720));
  NAND2X1 g2662(.A(n3524), .B(n3274), .Y(n3721));
  INVX1   g2663(.A(n3231), .Y(n3722));
  AOI22X1 g2664(.A0(n3514), .A1(P1_REG2_REG_26__SCAN_IN), .B0(n3722), .B1(n3525), .Y(n3723));
  OAI21X1 g2665(.A0(n3545), .A1(n3282), .B0(n3723), .Y(n3724));
  AOI21X1 g2666(.A0(n3519), .A1(n3243), .B0(n3724), .Y(n3725));
  NAND2X1 g2667(.A(n3725), .B(n3721), .Y(n3726));
  AOI21X1 g2668(.A0(n3520), .A1(n3262), .B0(n3726), .Y(n3727));
  OAI21X1 g2669(.A0(n3514), .A1(n3720), .B0(n3727), .Y(P1_U3267));
  NOR3X1  g2670(.A(n3311), .B(n3310), .C(n3301), .Y(n3729));
  NAND2X1 g2671(.A(n3524), .B(n3313), .Y(n3730));
  INVX1   g2672(.A(n3277), .Y(n3731));
  AOI22X1 g2673(.A0(n3514), .A1(P1_REG2_REG_27__SCAN_IN), .B0(n3731), .B1(n3525), .Y(n3732));
  OAI21X1 g2674(.A0(n3545), .A1(n3322), .B0(n3732), .Y(n3733));
  AOI21X1 g2675(.A0(n3519), .A1(n3333), .B0(n3733), .Y(n3734));
  NAND2X1 g2676(.A(n3734), .B(n3730), .Y(n3735));
  AOI21X1 g2677(.A0(n3520), .A1(n3298), .B0(n3735), .Y(n3736));
  OAI21X1 g2678(.A0(n3514), .A1(n3729), .B0(n3736), .Y(P1_U3266));
  NOR3X1  g2679(.A(n3356), .B(n3353), .C(n3342), .Y(n3738));
  NAND2X1 g2680(.A(n3524), .B(n3359), .Y(n3739));
  AOI22X1 g2681(.A0(n3514), .A1(P1_REG2_REG_28__SCAN_IN), .B0(n3317), .B1(n3525), .Y(n3740));
  OAI21X1 g2682(.A0(n3545), .A1(n3364), .B0(n3740), .Y(n3741));
  AOI21X1 g2683(.A0(n3519), .A1(n3329), .B0(n3741), .Y(n3742));
  NAND2X1 g2684(.A(n3742), .B(n3739), .Y(n3743));
  AOI21X1 g2685(.A0(n3520), .A1(n3350), .B0(n3743), .Y(n3744));
  OAI21X1 g2686(.A0(n3514), .A1(n3738), .B0(n3744), .Y(P1_U3265));
  NAND3X1 g2687(.A(n3415), .B(n3414), .C(n3409), .Y(n3746));
  OAI21X1 g2688(.A0(n3746), .A1(n3387), .B0(n3515), .Y(n3747));
  NAND2X1 g2689(.A(n3520), .B(n3376), .Y(n3748));
  NAND3X1 g2690(.A(n3276), .B(P1_REG3_REG_27__SCAN_IN), .C(P1_REG3_REG_28__SCAN_IN), .Y(n3749));
  NOR3X1  g2691(.A(n3514), .B(n3506), .C(n3749), .Y(n3750));
  AOI21X1 g2692(.A0(n3514), .A1(P1_REG2_REG_29__SCAN_IN), .B0(n3750), .Y(n3751));
  OAI21X1 g2693(.A0(n3551), .A1(n3401), .B0(n3751), .Y(n3752));
  AOI21X1 g2694(.A0(n3524), .A1(n3411), .B0(n3752), .Y(n3753));
  NAND3X1 g2695(.A(n3753), .B(n3748), .C(n3747), .Y(P1_U3356));
  NAND2X1 g2696(.A(n3524), .B(n3422), .Y(n3755));
  INVX1   g2697(.A(n1829), .Y(n3756));
  NAND2X1 g2698(.A(n1834), .B(n1832), .Y(n3757));
  XOR2X1  g2699(.A(n1837), .B(n3757), .Y(n3758));
  OAI21X1 g2700(.A0(n3758), .A1(n1152), .B0(n3756), .Y(n3759));
  NAND3X1 g2701(.A(n3519), .B(n3119), .C(n3759), .Y(n3760));
  NAND3X1 g2702(.A(n3512), .B(n3426), .C(n1891), .Y(n3761));
  NAND2X1 g2703(.A(n3514), .B(P1_REG2_REG_30__SCAN_IN), .Y(n3762));
  NAND4X1 g2704(.A(n3761), .B(n3760), .C(n3755), .D(n3762), .Y(P1_U3264));
  NAND2X1 g2705(.A(n3524), .B(n3434), .Y(n3764));
  INVX1   g2706(.A(n1851), .Y(n3765));
  OAI21X1 g2707(.A0(n1843), .A1(n1831), .B0(n1856), .Y(n3766));
  NAND4X1 g2708(.A(n1855), .B(n1834), .C(n1832), .D(n1860), .Y(n3767));
  NAND4X1 g2709(.A(n3767), .B(n3766), .C(n1145), .D(n1864), .Y(n3768));
  AOI21X1 g2710(.A0(n3768), .A1(n3765), .B0(n2003), .Y(n3769));
  NAND2X1 g2711(.A(n3519), .B(n3769), .Y(n3770));
  NAND2X1 g2712(.A(n3514), .B(P1_REG2_REG_31__SCAN_IN), .Y(n3771));
  NAND4X1 g2713(.A(n3770), .B(n3764), .C(n3761), .D(n3771), .Y(P1_U3263));
  OAI21X1 g2714(.A0(n3378), .A1(n1882), .B0(n1872), .Y(n3773));
  NAND2X1 g2715(.A(n3773), .B(n3119), .Y(n3774));
  NOR4X1  g2716(.A(n1882), .B(n1873), .C(P1_U3086), .D(n3774), .Y(n3775));
  INVX1   g2717(.A(P1_REG2_REG_18__SCAN_IN), .Y(n3776));
  INVX1   g2718(.A(P1_REG2_REG_16__SCAN_IN), .Y(n3777));
  INVX1   g2719(.A(P1_REG2_REG_17__SCAN_IN), .Y(n3778));
  AOI22X1 g2720(.A0(n2803), .A1(n3777), .B0(n3778), .B1(n2850), .Y(n3779));
  INVX1   g2721(.A(P1_REG2_REG_13__SCAN_IN), .Y(n3780));
  NAND2X1 g2722(.A(n2662), .B(n3780), .Y(n3781));
  INVX1   g2723(.A(P1_REG2_REG_11__SCAN_IN), .Y(n3782));
  NOR2X1  g2724(.A(n2559), .B(n3782), .Y(n3783));
  INVX1   g2725(.A(n3783), .Y(n3784));
  INVX1   g2726(.A(P1_REG2_REG_12__SCAN_IN), .Y(n3785));
  AOI22X1 g2727(.A0(n2611), .A1(n3785), .B0(n3780), .B1(n2662), .Y(n3786));
  INVX1   g2728(.A(n3786), .Y(n3787));
  NOR2X1  g2729(.A(n2611), .B(n3785), .Y(n3788));
  AOI21X1 g2730(.A0(n2663), .A1(P1_REG2_REG_13__SCAN_IN), .B0(n3788), .Y(n3789));
  OAI21X1 g2731(.A0(n3787), .A1(n3784), .B0(n3789), .Y(n3790));
  INVX1   g2732(.A(P1_REG2_REG_10__SCAN_IN), .Y(n3791));
  INVX1   g2733(.A(P1_REG2_REG_8__SCAN_IN), .Y(n3792));
  NOR2X1  g2734(.A(n2421), .B(n3792), .Y(n3793));
  INVX1   g2735(.A(P1_REG2_REG_9__SCAN_IN), .Y(n3794));
  AOI22X1 g2736(.A0(n2466), .A1(n3794), .B0(n3791), .B1(n2513), .Y(n3795));
  OAI22X1 g2737(.A0(n2466), .A1(n3794), .B0(n3791), .B1(n2513), .Y(n3796));
  AOI21X1 g2738(.A0(n3795), .A1(n3793), .B0(n3796), .Y(n3797));
  AOI21X1 g2739(.A0(n2513), .A1(n3791), .B0(n3797), .Y(n3798));
  OAI22X1 g2740(.A0(n2322), .A1(P1_REG2_REG_6__SCAN_IN), .B0(P1_REG2_REG_7__SCAN_IN), .B1(n2374), .Y(n3799));
  AOI22X1 g2741(.A0(n2221), .A1(n3550), .B0(n2247), .B1(n2265), .Y(n3800));
  AOI22X1 g2742(.A0(n2111), .A1(n3536), .B0(n3543), .B1(n2162), .Y(n3801));
  NOR2X1  g2743(.A(n2004), .B(n2019), .Y(n3802));
  OAI21X1 g2744(.A0(n2073), .A1(P1_REG2_REG_1__SCAN_IN), .B0(n3802), .Y(n3803));
  INVX1   g2745(.A(n3803), .Y(n3804));
  NOR2X1  g2746(.A(n2072), .B(n2051), .Y(n3805));
  OAI21X1 g2747(.A0(n3805), .A1(n3804), .B0(n3801), .Y(n3806));
  NOR2X1  g2748(.A(n2162), .B(n3543), .Y(n3807));
  INVX1   g2749(.A(n3807), .Y(n3808));
  NOR2X1  g2750(.A(n2111), .B(n3536), .Y(n3809));
  OAI21X1 g2751(.A0(n2163), .A1(P1_REG2_REG_3__SCAN_IN), .B0(n3809), .Y(n3810));
  NAND3X1 g2752(.A(n3810), .B(n3808), .C(n3806), .Y(n3811));
  NAND2X1 g2753(.A(n3811), .B(n3800), .Y(n3812));
  NOR2X1  g2754(.A(n2221), .B(n3550), .Y(n3813));
  INVX1   g2755(.A(n3813), .Y(n3814));
  AOI21X1 g2756(.A0(n3814), .A1(n2247), .B0(n2265), .Y(n3815));
  AOI21X1 g2757(.A0(n3813), .A1(P1_REG2_REG_5__SCAN_IN), .B0(n3815), .Y(n3816));
  NAND2X1 g2758(.A(n3816), .B(n3812), .Y(n3817));
  INVX1   g2759(.A(n3817), .Y(n3818));
  NOR2X1  g2760(.A(n2321), .B(n2303), .Y(n3819));
  INVX1   g2761(.A(P1_REG2_REG_7__SCAN_IN), .Y(n3820));
  INVX1   g2762(.A(n3819), .Y(n3821));
  AOI21X1 g2763(.A0(n3821), .A1(n3820), .B0(n2373), .Y(n3822));
  AOI21X1 g2764(.A0(n3819), .A1(P1_REG2_REG_7__SCAN_IN), .B0(n3822), .Y(n3823));
  OAI21X1 g2765(.A0(n3818), .A1(n3799), .B0(n3823), .Y(n3824));
  NOR2X1  g2766(.A(n2422), .B(P1_REG2_REG_8__SCAN_IN), .Y(n3825));
  INVX1   g2767(.A(n3825), .Y(n3826));
  NAND3X1 g2768(.A(n3826), .B(n3824), .C(n3795), .Y(n3827));
  INVX1   g2769(.A(n3827), .Y(n3828));
  NOR2X1  g2770(.A(n3828), .B(n3798), .Y(n3829));
  NOR2X1  g2771(.A(n2560), .B(P1_REG2_REG_11__SCAN_IN), .Y(n3830));
  NOR3X1  g2772(.A(n3830), .B(n3829), .C(n3787), .Y(n3831));
  AOI21X1 g2773(.A0(n3790), .A1(n3781), .B0(n3831), .Y(n3832));
  AOI21X1 g2774(.A0(n2711), .A1(n3628), .B0(n3832), .Y(n3833));
  AOI21X1 g2775(.A0(n2712), .A1(P1_REG2_REG_14__SCAN_IN), .B0(n3833), .Y(n3834));
  AOI21X1 g2776(.A0(n2756), .A1(n3633), .B0(n3834), .Y(n3835));
  AOI21X1 g2777(.A0(n2757), .A1(P1_REG2_REG_15__SCAN_IN), .B0(n3835), .Y(n3836));
  INVX1   g2778(.A(n3836), .Y(n3837));
  NOR2X1  g2779(.A(n2803), .B(n3777), .Y(n3838));
  INVX1   g2780(.A(n3838), .Y(n3839));
  AOI21X1 g2781(.A0(n3839), .A1(n3778), .B0(n2850), .Y(n3840));
  AOI21X1 g2782(.A0(n3838), .A1(P1_REG2_REG_17__SCAN_IN), .B0(n3840), .Y(n3841));
  INVX1   g2783(.A(n3841), .Y(n3842));
  AOI21X1 g2784(.A0(n3837), .A1(n3779), .B0(n3842), .Y(n3843));
  OAI21X1 g2785(.A0(n2904), .A1(n3776), .B0(n3843), .Y(n3844));
  XOR2X1  g2786(.A(n1991), .B(P1_REG2_REG_19__SCAN_IN), .Y(n3845));
  AOI21X1 g2787(.A0(n2904), .A1(n3776), .B0(n3845), .Y(n3846));
  NAND2X1 g2788(.A(n3846), .B(n3844), .Y(n3847));
  AOI21X1 g2789(.A0(n2904), .A1(n3776), .B0(n3843), .Y(n3848));
  OAI21X1 g2790(.A0(n2904), .A1(n3776), .B0(n3845), .Y(n3849));
  OAI21X1 g2791(.A0(n3849), .A1(n3848), .B0(n3847), .Y(n3850));
  NOR4X1  g2792(.A(n2040), .B(n2038), .C(n2029), .D(n3522), .Y(n3851));
  NOR2X1  g2793(.A(n1992), .B(n1982), .Y(n3852));
  NOR4X1  g2794(.A(n3852), .B(n2041), .C(n2034), .D(n3505), .Y(n3853));
  NAND2X1 g2795(.A(n1989), .B(n1985), .Y(n3854));
  NAND4X1 g2796(.A(n3853), .B(n3851), .C(n3518), .D(n3854), .Y(n3855));
  INVX1   g2797(.A(n3855), .Y(n3856));
  INVX1   g2798(.A(n2002), .Y(n3857));
  NOR2X1  g2799(.A(n3857), .B(n2080), .Y(n3858));
  INVX1   g2800(.A(n3858), .Y(n3859));
  INVX1   g2801(.A(P1_REG1_REG_17__SCAN_IN), .Y(n3862));
  AOI22X1 g2802(.A0(n2803), .A1(n2788), .B0(n3862), .B1(n2850), .Y(n3863));
  INVX1   g2803(.A(P1_REG1_REG_15__SCAN_IN), .Y(n3864));
  NOR2X1  g2804(.A(n2663), .B(P1_REG1_REG_13__SCAN_IN), .Y(n3865));
  INVX1   g2805(.A(P1_REG1_REG_11__SCAN_IN), .Y(n3866));
  NOR2X1  g2806(.A(n2559), .B(n3866), .Y(n3867));
  INVX1   g2807(.A(P1_REG1_REG_12__SCAN_IN), .Y(n3868));
  INVX1   g2808(.A(P1_REG1_REG_13__SCAN_IN), .Y(n3869));
  AOI22X1 g2809(.A0(n2611), .A1(n3868), .B0(n3869), .B1(n2662), .Y(n3870));
  NAND2X1 g2810(.A(n3870), .B(n3867), .Y(n3871));
  NOR2X1  g2811(.A(n2611), .B(n3868), .Y(n3872));
  AOI21X1 g2812(.A0(n2663), .A1(P1_REG1_REG_13__SCAN_IN), .B0(n3872), .Y(n3873));
  AOI21X1 g2813(.A0(n3873), .A1(n3871), .B0(n3865), .Y(n3874));
  NOR2X1  g2814(.A(n2612), .B(P1_REG1_REG_12__SCAN_IN), .Y(n3875));
  INVX1   g2815(.A(P1_REG1_REG_10__SCAN_IN), .Y(n3876));
  NAND2X1 g2816(.A(n2513), .B(n3876), .Y(n3877));
  INVX1   g2817(.A(P1_REG1_REG_8__SCAN_IN), .Y(n3878));
  NOR2X1  g2818(.A(n2421), .B(n3878), .Y(n3879));
  INVX1   g2819(.A(P1_REG1_REG_9__SCAN_IN), .Y(n3880));
  AOI22X1 g2820(.A0(n2466), .A1(n3880), .B0(n3876), .B1(n2513), .Y(n3881));
  NAND2X1 g2821(.A(n3881), .B(n3879), .Y(n3882));
  AOI22X1 g2822(.A0(n2467), .A1(P1_REG1_REG_9__SCAN_IN), .B0(P1_REG1_REG_10__SCAN_IN), .B1(n2514), .Y(n3883));
  NAND2X1 g2823(.A(n3883), .B(n3882), .Y(n3884));
  INVX1   g2824(.A(P1_REG1_REG_6__SCAN_IN), .Y(n3885));
  INVX1   g2825(.A(P1_REG1_REG_7__SCAN_IN), .Y(n3886));
  AOI22X1 g2826(.A0(n2321), .A1(n3885), .B0(n3886), .B1(n2373), .Y(n3887));
  INVX1   g2827(.A(n3887), .Y(n3888));
  INVX1   g2828(.A(P1_REG1_REG_5__SCAN_IN), .Y(n3889));
  AOI22X1 g2829(.A0(n2221), .A1(n2200), .B0(n3889), .B1(n2265), .Y(n3890));
  AOI22X1 g2830(.A0(n2111), .A1(n2183), .B0(n2142), .B1(n2162), .Y(n3891));
  INVX1   g2831(.A(P1_REG1_REG_1__SCAN_IN), .Y(n3892));
  OAI21X1 g2832(.A0(n2006), .A1(n2005), .B0(P1_REG1_REG_0__SCAN_IN), .Y(n3893));
  AOI21X1 g2833(.A0(n2072), .A1(n3892), .B0(n3893), .Y(n3894));
  NOR2X1  g2834(.A(n2072), .B(n3892), .Y(n3895));
  OAI21X1 g2835(.A0(n3895), .A1(n3894), .B0(n3891), .Y(n3896));
  NOR2X1  g2836(.A(n2162), .B(n2142), .Y(n3897));
  INVX1   g2837(.A(n3897), .Y(n3898));
  NOR2X1  g2838(.A(n2111), .B(n2183), .Y(n3899));
  OAI21X1 g2839(.A0(n2163), .A1(P1_REG1_REG_3__SCAN_IN), .B0(n3899), .Y(n3900));
  NAND3X1 g2840(.A(n3900), .B(n3898), .C(n3896), .Y(n3901));
  NAND2X1 g2841(.A(n3901), .B(n3890), .Y(n3902));
  NOR2X1  g2842(.A(n2221), .B(n2200), .Y(n3903));
  INVX1   g2843(.A(n3903), .Y(n3904));
  AOI21X1 g2844(.A0(n3904), .A1(n3889), .B0(n2265), .Y(n3905));
  AOI21X1 g2845(.A0(n3903), .A1(P1_REG1_REG_5__SCAN_IN), .B0(n3905), .Y(n3906));
  NAND2X1 g2846(.A(n3906), .B(n3902), .Y(n3907));
  INVX1   g2847(.A(n3907), .Y(n3908));
  NOR3X1  g2848(.A(n2321), .B(n3886), .C(n3885), .Y(n3909));
  OAI21X1 g2849(.A0(n2321), .A1(n3885), .B0(n3886), .Y(n3910));
  AOI21X1 g2850(.A0(n3910), .A1(n2374), .B0(n3909), .Y(n3911));
  OAI21X1 g2851(.A0(n3908), .A1(n3888), .B0(n3911), .Y(n3912));
  INVX1   g2852(.A(n3881), .Y(n3913));
  NOR2X1  g2853(.A(n2422), .B(P1_REG1_REG_8__SCAN_IN), .Y(n3914));
  NOR2X1  g2854(.A(n3914), .B(n3913), .Y(n3915));
  AOI22X1 g2855(.A0(n3912), .A1(n3915), .B0(n3884), .B1(n3877), .Y(n3916));
  NOR2X1  g2856(.A(n2560), .B(P1_REG1_REG_11__SCAN_IN), .Y(n3917));
  NOR4X1  g2857(.A(n3916), .B(n3875), .C(n3865), .D(n3917), .Y(n3918));
  NOR2X1  g2858(.A(n3918), .B(n3874), .Y(n3919));
  AOI21X1 g2859(.A0(n2711), .A1(n2699), .B0(n3919), .Y(n3920));
  AOI21X1 g2860(.A0(n2712), .A1(P1_REG1_REG_14__SCAN_IN), .B0(n3920), .Y(n3921));
  AOI21X1 g2861(.A0(n2756), .A1(n3864), .B0(n3921), .Y(n3922));
  AOI21X1 g2862(.A0(n2757), .A1(P1_REG1_REG_15__SCAN_IN), .B0(n3922), .Y(n3923));
  INVX1   g2863(.A(n3923), .Y(n3924));
  NOR2X1  g2864(.A(n2803), .B(n2788), .Y(n3925));
  INVX1   g2865(.A(n3925), .Y(n3926));
  AOI21X1 g2866(.A0(n3926), .A1(n3862), .B0(n2850), .Y(n3927));
  AOI21X1 g2867(.A0(n3925), .A1(P1_REG1_REG_17__SCAN_IN), .B0(n3927), .Y(n3928));
  INVX1   g2868(.A(n3928), .Y(n3929));
  AOI21X1 g2869(.A0(n3924), .A1(n3863), .B0(n3929), .Y(n3930));
  INVX1   g2870(.A(n3930), .Y(n3931));
  NOR2X1  g2871(.A(n2904), .B(n2888), .Y(n3932));
  XOR2X1  g2872(.A(n1991), .B(P1_REG1_REG_19__SCAN_IN), .Y(n3933));
  AOI21X1 g2873(.A0(n2904), .A1(n2888), .B0(n3933), .Y(n3934));
  OAI21X1 g2874(.A0(n3932), .A1(n3931), .B0(n3934), .Y(n3935));
  AOI21X1 g2875(.A0(n2904), .A1(n2888), .B0(n3930), .Y(n3936));
  OAI21X1 g2876(.A0(n2904), .A1(n2888), .B0(n3933), .Y(n3937));
  OAI21X1 g2877(.A0(n3937), .A1(n3936), .B0(n3935), .Y(n3938));
  INVX1   g2878(.A(n3938), .Y(n3939));
  INVX1   g2879(.A(n2080), .Y(n3941));
  AOI22X1 g2880(.A0(n3857), .A1(n3939), .B0(n2037), .B1(n2080), .Y(n3943));
  OAI21X1 g2881(.A0(n3859), .A1(n3850), .B0(n3943), .Y(n3944));
  NAND2X1 g2882(.A(n3944), .B(n3775), .Y(n3945));
  NAND3X1 g2883(.A(n1884), .B(n1878), .C(n1875), .Y(n3946));
  NOR2X1  g2884(.A(n3946), .B(n1873), .Y(n3947));
  NAND2X1 g2885(.A(n3774), .B(P1_STATE_REG_SCAN_IN), .Y(P1_U3085));
  NOR2X1  g2886(.A(P1_U3085), .B(n3947), .Y(n3949));
  NOR4X1  g2887(.A(n2002), .B(n1872), .C(P1_U3086), .D(n3949), .Y(n3950));
  NOR4X1  g2888(.A(n3949), .B(n1872), .C(P1_U3086), .D(n3859), .Y(n3951));
  INVX1   g2889(.A(n3951), .Y(n3952));
  NOR4X1  g2890(.A(n3941), .B(n1872), .C(P1_U3086), .D(n3949), .Y(n3953));
  INVX1   g2891(.A(n3949), .Y(n3954));
  OAI22X1 g2892(.A0(P1_STATE_REG_SCAN_IN), .A1(n2969), .B0(n1086), .B1(n3954), .Y(n3955));
  AOI21X1 g2893(.A0(n3953), .A1(n2037), .B0(n3955), .Y(n3956));
  OAI21X1 g2894(.A0(n3952), .A1(n3850), .B0(n3956), .Y(n3957));
  AOI21X1 g2895(.A0(n3950), .A1(n3939), .B0(n3957), .Y(n3958));
  NAND2X1 g2896(.A(n3958), .B(n3945), .Y(P1_U3262));
  XOR2X1  g2897(.A(n2904), .B(P1_REG2_REG_18__SCAN_IN), .Y(n3960));
  INVX1   g2898(.A(n3960), .Y(n3961));
  XOR2X1  g2899(.A(n3961), .B(n3843), .Y(n3962));
  NOR2X1  g2900(.A(n3962), .B(n3859), .Y(n3963));
  XOR2X1  g2901(.A(n2904), .B(n2888), .Y(n3966));
  XOR2X1  g2902(.A(n3966), .B(n3930), .Y(n3967));
  OAI22X1 g2903(.A0(n3941), .A1(n2904), .B0(n2002), .B1(n3967), .Y(n3968));
  OAI21X1 g2904(.A0(n3968), .A1(n3963), .B0(n3775), .Y(n3969));
  INVX1   g2905(.A(n3950), .Y(n3970));
  NOR2X1  g2906(.A(n3967), .B(n3970), .Y(n3971));
  NOR2X1  g2907(.A(n3962), .B(n3952), .Y(n3972));
  INVX1   g2908(.A(n3953), .Y(n3973));
  AOI22X1 g2909(.A0(P1_U3086), .A1(P1_REG3_REG_18__SCAN_IN), .B0(P1_ADDR_REG_18__SCAN_IN), .B1(n3949), .Y(n3974));
  OAI21X1 g2910(.A0(n3973), .A1(n2904), .B0(n3974), .Y(n3975));
  NOR3X1  g2911(.A(n3975), .B(n3972), .C(n3971), .Y(n3976));
  NAND2X1 g2912(.A(n3976), .B(n3969), .Y(P1_U3261));
  INVX1   g2913(.A(n3775), .Y(n3978));
  OAI21X1 g2914(.A0(n2850), .A1(n3778), .B0(n3779), .Y(n3979));
  AOI21X1 g2915(.A0(n3839), .A1(n3836), .B0(n3979), .Y(n3980));
  NOR2X1  g2916(.A(n2804), .B(P1_REG2_REG_16__SCAN_IN), .Y(n3981));
  INVX1   g2917(.A(n3981), .Y(n3982));
  XOR2X1  g2918(.A(n2850), .B(P1_REG2_REG_17__SCAN_IN), .Y(n3983));
  OAI21X1 g2919(.A0(n2803), .A1(n3777), .B0(n3983), .Y(n3984));
  AOI21X1 g2920(.A0(n3837), .A1(n3982), .B0(n3984), .Y(n3985));
  NOR3X1  g2921(.A(n3985), .B(n3980), .C(n3859), .Y(n3986));
  OAI21X1 g2922(.A0(n2850), .A1(n3862), .B0(n3863), .Y(n3987));
  AOI21X1 g2923(.A0(n3926), .A1(n3923), .B0(n3987), .Y(n3988));
  AOI21X1 g2924(.A0(n2803), .A1(n2788), .B0(n3923), .Y(n3989));
  XOR2X1  g2925(.A(n2850), .B(n3862), .Y(n3990));
  NOR3X1  g2926(.A(n3990), .B(n3989), .C(n3925), .Y(n3991));
  NOR3X1  g2927(.A(n3991), .B(n3988), .C(n2002), .Y(n3992));
  NOR3X1  g2928(.A(n3856), .B(n2850), .C(n3941), .Y(n3993));
  NOR3X1  g2929(.A(n3993), .B(n3992), .C(n3986), .Y(n3994));
  NOR3X1  g2930(.A(n3991), .B(n3988), .C(n3970), .Y(n3995));
  NOR3X1  g2931(.A(n3985), .B(n3980), .C(n3952), .Y(n3996));
  AOI22X1 g2932(.A0(P1_U3086), .A1(P1_REG3_REG_17__SCAN_IN), .B0(P1_ADDR_REG_17__SCAN_IN), .B1(n3949), .Y(n3997));
  OAI21X1 g2933(.A0(n3973), .A1(n2850), .B0(n3997), .Y(n3998));
  NOR3X1  g2934(.A(n3998), .B(n3996), .C(n3995), .Y(n3999));
  OAI21X1 g2935(.A0(n3994), .A1(n3978), .B0(n3999), .Y(P1_U3260));
  XOR2X1  g2936(.A(n2803), .B(n3777), .Y(n4001));
  AOI21X1 g2937(.A0(n3839), .A1(n3982), .B0(n3836), .Y(n4002));
  AOI21X1 g2938(.A0(n4001), .A1(n3836), .B0(n4002), .Y(n4003));
  NOR2X1  g2939(.A(n4003), .B(n3859), .Y(n4004));
  XOR2X1  g2940(.A(n2803), .B(n2788), .Y(n4005));
  NOR2X1  g2941(.A(n4005), .B(n3923), .Y(n4007));
  AOI21X1 g2942(.A0(n4005), .A1(n3923), .B0(n4007), .Y(n4008));
  OAI22X1 g2943(.A0(n3941), .A1(n2803), .B0(n2002), .B1(n4008), .Y(n4009));
  OAI21X1 g2944(.A0(n4009), .A1(n4004), .B0(n3775), .Y(n4010));
  NOR2X1  g2945(.A(n4008), .B(n3970), .Y(n4011));
  NOR2X1  g2946(.A(n4003), .B(n3952), .Y(n4012));
  AOI22X1 g2947(.A0(P1_U3086), .A1(P1_REG3_REG_16__SCAN_IN), .B0(P1_ADDR_REG_16__SCAN_IN), .B1(n3949), .Y(n4013));
  OAI21X1 g2948(.A0(n3973), .A1(n2803), .B0(n4013), .Y(n4014));
  NOR3X1  g2949(.A(n4014), .B(n4012), .C(n4011), .Y(n4015));
  NAND2X1 g2950(.A(n4015), .B(n4010), .Y(P1_U3259));
  XOR2X1  g2951(.A(n2756), .B(P1_REG2_REG_15__SCAN_IN), .Y(n4017));
  XOR2X1  g2952(.A(n4017), .B(n3834), .Y(n4018));
  XOR2X1  g2953(.A(n2756), .B(n3864), .Y(n4019));
  XOR2X1  g2954(.A(n4019), .B(n3921), .Y(n4020));
  OAI22X1 g2955(.A0(n3941), .A1(n2756), .B0(n2002), .B1(n4020), .Y(n4021));
  AOI21X1 g2956(.A0(n4018), .A1(n3858), .B0(n4021), .Y(n4022));
  NOR2X1  g2957(.A(n4020), .B(n3970), .Y(n4023));
  NAND2X1 g2958(.A(n4018), .B(n3951), .Y(n4024));
  NAND2X1 g2959(.A(n3953), .B(n2757), .Y(n4025));
  AOI22X1 g2960(.A0(P1_U3086), .A1(P1_REG3_REG_15__SCAN_IN), .B0(P1_ADDR_REG_15__SCAN_IN), .B1(n3949), .Y(n4026));
  NAND3X1 g2961(.A(n4026), .B(n4025), .C(n4024), .Y(n4027));
  NOR2X1  g2962(.A(n4027), .B(n4023), .Y(n4028));
  OAI21X1 g2963(.A0(n4022), .A1(n3978), .B0(n4028), .Y(P1_U3258));
  XOR2X1  g2964(.A(n2711), .B(P1_REG2_REG_14__SCAN_IN), .Y(n4030));
  XOR2X1  g2965(.A(n4030), .B(n3832), .Y(n4031));
  NAND2X1 g2966(.A(n4031), .B(n3858), .Y(n4032));
  XOR2X1  g2967(.A(n2711), .B(P1_REG1_REG_14__SCAN_IN), .Y(n4033));
  XOR2X1  g2968(.A(n4033), .B(n3919), .Y(n4034));
  AOI22X1 g2969(.A0(n2080), .A1(n2712), .B0(n3857), .B1(n4034), .Y(n4035));
  NAND2X1 g2970(.A(n4035), .B(n4032), .Y(n4036));
  NAND2X1 g2971(.A(n4036), .B(n3775), .Y(n4037));
  NAND2X1 g2972(.A(n4031), .B(n3951), .Y(n4038));
  AOI22X1 g2973(.A0(P1_U3086), .A1(P1_REG3_REG_14__SCAN_IN), .B0(P1_ADDR_REG_14__SCAN_IN), .B1(n3949), .Y(n4039));
  AOI22X1 g2974(.A0(n3953), .A1(n2712), .B0(n3950), .B1(n4034), .Y(n4040));
  NAND4X1 g2975(.A(n4039), .B(n4038), .C(n4037), .D(n4040), .Y(P1_U3257));
  INVX1   g2976(.A(n3788), .Y(n4042));
  INVX1   g2977(.A(n3829), .Y(n4043));
  INVX1   g2978(.A(n3830), .Y(n4044));
  AOI21X1 g2979(.A0(n4044), .A1(n4043), .B0(n3783), .Y(n4045));
  OAI21X1 g2980(.A0(n2662), .A1(n3780), .B0(n3786), .Y(n4046));
  AOI21X1 g2981(.A0(n4045), .A1(n4042), .B0(n4046), .Y(n4047));
  NOR2X1  g2982(.A(n2612), .B(P1_REG2_REG_12__SCAN_IN), .Y(n4048));
  NOR2X1  g2983(.A(n4045), .B(n4048), .Y(n4049));
  XOR2X1  g2984(.A(n2662), .B(n3780), .Y(n4050));
  NOR3X1  g2985(.A(n4050), .B(n4049), .C(n3788), .Y(n4051));
  NOR3X1  g2986(.A(n4051), .B(n4047), .C(n3859), .Y(n4052));
  INVX1   g2987(.A(n3916), .Y(n4053));
  INVX1   g2988(.A(n3917), .Y(n4054));
  AOI21X1 g2989(.A0(n4054), .A1(n4053), .B0(n3867), .Y(n4055));
  INVX1   g2990(.A(n4055), .Y(n4056));
  NOR2X1  g2991(.A(n4056), .B(n3872), .Y(n4057));
  OAI21X1 g2992(.A0(n2662), .A1(n3869), .B0(n3870), .Y(n4058));
  XOR2X1  g2993(.A(n2662), .B(n3869), .Y(n4059));
  NOR2X1  g2994(.A(n4059), .B(n3872), .Y(n4060));
  OAI21X1 g2995(.A0(n4055), .A1(n3875), .B0(n4060), .Y(n4061));
  OAI21X1 g2996(.A0(n4058), .A1(n4057), .B0(n4061), .Y(n4062));
  OAI22X1 g2997(.A0(n3941), .A1(n2662), .B0(n2002), .B1(n4062), .Y(n4063));
  OAI21X1 g2998(.A0(n4063), .A1(n4052), .B0(n3775), .Y(n4064));
  NOR2X1  g2999(.A(n4062), .B(n3970), .Y(n4065));
  NOR3X1  g3000(.A(n4051), .B(n4047), .C(n3952), .Y(n4066));
  AOI22X1 g3001(.A0(P1_U3086), .A1(P1_REG3_REG_13__SCAN_IN), .B0(P1_ADDR_REG_13__SCAN_IN), .B1(n3949), .Y(n4067));
  OAI21X1 g3002(.A0(n3973), .A1(n2662), .B0(n4067), .Y(n4068));
  NOR3X1  g3003(.A(n4068), .B(n4066), .C(n4065), .Y(n4069));
  NAND2X1 g3004(.A(n4069), .B(n4064), .Y(P1_U3256));
  XOR2X1  g3005(.A(n2611), .B(n3785), .Y(n4073));
  NOR2X1  g3006(.A(n4073), .B(n4045), .Y(n4074));
  AOI21X1 g3007(.A0(n4073), .A1(n4045), .B0(n4074), .Y(n4075));
  NOR2X1  g3008(.A(n4075), .B(n3859), .Y(n4076));
  XOR2X1  g3009(.A(n2611), .B(n3868), .Y(n4077));
  NOR2X1  g3010(.A(n4077), .B(n4055), .Y(n4079));
  AOI21X1 g3011(.A0(n4077), .A1(n4055), .B0(n4079), .Y(n4080));
  OAI22X1 g3012(.A0(n3941), .A1(n2611), .B0(n2002), .B1(n4080), .Y(n4081));
  OAI21X1 g3013(.A0(n4081), .A1(n4076), .B0(n3775), .Y(n4082));
  AOI22X1 g3014(.A0(P1_U3086), .A1(P1_REG3_REG_12__SCAN_IN), .B0(P1_ADDR_REG_12__SCAN_IN), .B1(n3949), .Y(n4083));
  OAI21X1 g3015(.A0(n4075), .A1(n3952), .B0(n4083), .Y(n4084));
  OAI22X1 g3016(.A0(n3973), .A1(n2611), .B0(n3970), .B1(n4080), .Y(n4085));
  NOR2X1  g3017(.A(n4085), .B(n4084), .Y(n4086));
  NAND2X1 g3018(.A(n4086), .B(n4082), .Y(P1_U3255));
  XOR2X1  g3019(.A(n2559), .B(n3782), .Y(n4088));
  AOI21X1 g3020(.A0(n4044), .A1(n3784), .B0(n3829), .Y(n4089));
  AOI21X1 g3021(.A0(n4088), .A1(n3829), .B0(n4089), .Y(n4090));
  NOR2X1  g3022(.A(n4090), .B(n3859), .Y(n4091));
  XOR2X1  g3023(.A(n2559), .B(n3866), .Y(n4092));
  NOR2X1  g3024(.A(n4092), .B(n3916), .Y(n4094));
  AOI21X1 g3025(.A0(n4092), .A1(n3916), .B0(n4094), .Y(n4095));
  OAI22X1 g3026(.A0(n3941), .A1(n2559), .B0(n2002), .B1(n4095), .Y(n4096));
  OAI21X1 g3027(.A0(n4096), .A1(n4091), .B0(n3775), .Y(n4097));
  AOI22X1 g3028(.A0(P1_U3086), .A1(P1_REG3_REG_11__SCAN_IN), .B0(P1_ADDR_REG_11__SCAN_IN), .B1(n3949), .Y(n4098));
  OAI21X1 g3029(.A0(n4090), .A1(n3952), .B0(n4098), .Y(n4099));
  OAI22X1 g3030(.A0(n3973), .A1(n2559), .B0(n3970), .B1(n4095), .Y(n4100));
  NOR2X1  g3031(.A(n4100), .B(n4099), .Y(n4101));
  NAND2X1 g3032(.A(n4101), .B(n4097), .Y(P1_U3254));
  NAND2X1 g3033(.A(n2467), .B(P1_REG2_REG_9__SCAN_IN), .Y(n4103));
  AOI21X1 g3034(.A0(n3826), .A1(n3824), .B0(n3793), .Y(n4104));
  OAI21X1 g3035(.A0(n2513), .A1(n3791), .B0(n3795), .Y(n4105));
  AOI21X1 g3036(.A0(n4104), .A1(n4103), .B0(n4105), .Y(n4106));
  AOI21X1 g3037(.A0(n2466), .A1(n3794), .B0(n4104), .Y(n4107));
  AOI22X1 g3038(.A0(n2467), .A1(P1_REG2_REG_9__SCAN_IN), .B0(n3791), .B1(n2514), .Y(n4108));
  OAI21X1 g3039(.A0(n2514), .A1(n3791), .B0(n4108), .Y(n4109));
  NOR2X1  g3040(.A(n4109), .B(n4107), .Y(n4110));
  NOR3X1  g3041(.A(n4110), .B(n4106), .C(n3859), .Y(n4111));
  NAND2X1 g3042(.A(n2467), .B(P1_REG1_REG_9__SCAN_IN), .Y(n4112));
  INVX1   g3043(.A(n3914), .Y(n4113));
  AOI21X1 g3044(.A0(n4113), .A1(n3912), .B0(n3879), .Y(n4114));
  OAI21X1 g3045(.A0(n2513), .A1(n3876), .B0(n3881), .Y(n4115));
  AOI21X1 g3046(.A0(n4114), .A1(n4112), .B0(n4115), .Y(n4116));
  AOI21X1 g3047(.A0(n2466), .A1(n3880), .B0(n4114), .Y(n4117));
  AOI22X1 g3048(.A0(n2467), .A1(P1_REG1_REG_9__SCAN_IN), .B0(n3876), .B1(n2514), .Y(n4118));
  OAI21X1 g3049(.A0(n2514), .A1(n3876), .B0(n4118), .Y(n4119));
  NOR2X1  g3050(.A(n4119), .B(n4117), .Y(n4120));
  NOR3X1  g3051(.A(n4120), .B(n4116), .C(n2002), .Y(n4121));
  NOR3X1  g3052(.A(n3856), .B(n2513), .C(n3941), .Y(n4122));
  NOR3X1  g3053(.A(n4122), .B(n4121), .C(n4111), .Y(n4123));
  NOR3X1  g3054(.A(n4110), .B(n4106), .C(n3952), .Y(n4124));
  INVX1   g3055(.A(n3947), .Y(n4125));
  NAND4X1 g3056(.A(n4125), .B(P1_STATE_REG_SCAN_IN), .C(P1_ADDR_REG_10__SCAN_IN), .D(n3774), .Y(n4126));
  OAI21X1 g3057(.A0(P1_STATE_REG_SCAN_IN), .A1(n2497), .B0(n4126), .Y(n4127));
  NOR3X1  g3058(.A(n4120), .B(n4116), .C(n3970), .Y(n4128));
  NOR2X1  g3059(.A(n3973), .B(n2513), .Y(n4129));
  NOR4X1  g3060(.A(n4128), .B(n4127), .C(n4124), .D(n4129), .Y(n4130));
  OAI21X1 g3061(.A0(n4123), .A1(n3978), .B0(n4130), .Y(P1_U3253));
  XOR2X1  g3062(.A(n2466), .B(n3794), .Y(n4132));
  NOR2X1  g3063(.A(n4132), .B(n4104), .Y(n4134));
  AOI21X1 g3064(.A0(n4132), .A1(n4104), .B0(n4134), .Y(n4135));
  NOR2X1  g3065(.A(n4135), .B(n3859), .Y(n4136));
  XOR2X1  g3066(.A(n2466), .B(n3880), .Y(n4137));
  NOR2X1  g3067(.A(n4137), .B(n4114), .Y(n4139));
  AOI21X1 g3068(.A0(n4137), .A1(n4114), .B0(n4139), .Y(n4140));
  OAI22X1 g3069(.A0(n3941), .A1(n2466), .B0(n2002), .B1(n4140), .Y(n4141));
  OAI21X1 g3070(.A0(n4141), .A1(n4136), .B0(n3775), .Y(n4142));
  AOI22X1 g3071(.A0(P1_U3086), .A1(P1_REG3_REG_9__SCAN_IN), .B0(P1_ADDR_REG_9__SCAN_IN), .B1(n3949), .Y(n4143));
  OAI21X1 g3072(.A0(n4135), .A1(n3952), .B0(n4143), .Y(n4144));
  OAI22X1 g3073(.A0(n3973), .A1(n2466), .B0(n3970), .B1(n4140), .Y(n4145));
  NOR2X1  g3074(.A(n4145), .B(n4144), .Y(n4146));
  NAND2X1 g3075(.A(n4146), .B(n4142), .Y(P1_U3252));
  NOR3X1  g3076(.A(n3856), .B(n2421), .C(n3941), .Y(n4148));
  XOR2X1  g3077(.A(n2421), .B(P1_REG1_REG_8__SCAN_IN), .Y(n4149));
  NOR2X1  g3078(.A(n4149), .B(n3912), .Y(n4150));
  AOI21X1 g3079(.A0(n4149), .A1(n3912), .B0(n4150), .Y(n4152));
  XOR2X1  g3080(.A(n2421), .B(P1_REG2_REG_8__SCAN_IN), .Y(n4153));
  NOR2X1  g3081(.A(n4153), .B(n3824), .Y(n4154));
  AOI21X1 g3082(.A0(n4153), .A1(n3824), .B0(n4154), .Y(n4156));
  OAI22X1 g3083(.A0(n4152), .A1(n2002), .B0(n3859), .B1(n4156), .Y(n4157));
  OAI21X1 g3084(.A0(n4157), .A1(n4148), .B0(n3775), .Y(n4158));
  AOI22X1 g3085(.A0(P1_U3086), .A1(P1_REG3_REG_8__SCAN_IN), .B0(P1_ADDR_REG_8__SCAN_IN), .B1(n3949), .Y(n4159));
  NOR2X1  g3086(.A(n4156), .B(n3952), .Y(n4160));
  OAI22X1 g3087(.A0(n3973), .A1(n2421), .B0(n3970), .B1(n4152), .Y(n4161));
  NOR2X1  g3088(.A(n4161), .B(n4160), .Y(n4162));
  NAND3X1 g3089(.A(n4162), .B(n4159), .C(n4158), .Y(P1_U3251));
  NOR2X1  g3090(.A(n2321), .B(n3885), .Y(n4164));
  AOI21X1 g3091(.A0(n2374), .A1(P1_REG1_REG_7__SCAN_IN), .B0(n3888), .Y(n4165));
  OAI21X1 g3092(.A0(n4164), .A1(n3907), .B0(n4165), .Y(n4166));
  AOI22X1 g3093(.A0(n3902), .A1(n3906), .B0(n2321), .B1(n3885), .Y(n4167));
  AOI21X1 g3094(.A0(n2374), .A1(n3886), .B0(n4164), .Y(n4168));
  OAI21X1 g3095(.A0(n2374), .A1(n3886), .B0(n4168), .Y(n4169));
  OAI21X1 g3096(.A0(n4169), .A1(n4167), .B0(n4166), .Y(n4170));
  INVX1   g3097(.A(n4170), .Y(n4171));
  NAND3X1 g3098(.A(n3821), .B(n3816), .C(n3812), .Y(n4172));
  AOI21X1 g3099(.A0(n2374), .A1(P1_REG2_REG_7__SCAN_IN), .B0(n3799), .Y(n4173));
  AOI22X1 g3100(.A0(n3812), .A1(n3816), .B0(n2321), .B1(n2303), .Y(n4174));
  AOI21X1 g3101(.A0(n2374), .A1(n3820), .B0(n3819), .Y(n4175));
  OAI21X1 g3102(.A0(n2374), .A1(n3820), .B0(n4175), .Y(n4176));
  NOR2X1  g3103(.A(n4176), .B(n4174), .Y(n4177));
  AOI21X1 g3104(.A0(n4173), .A1(n4172), .B0(n4177), .Y(n4178));
  AOI22X1 g3105(.A0(n4171), .A1(n3857), .B0(n3858), .B1(n4178), .Y(n4179));
  OAI21X1 g3106(.A0(n3941), .A1(n2373), .B0(n4179), .Y(n4180));
  NAND2X1 g3107(.A(n4180), .B(n3775), .Y(n4181));
  AOI22X1 g3108(.A0(P1_U3086), .A1(P1_REG3_REG_7__SCAN_IN), .B0(P1_ADDR_REG_7__SCAN_IN), .B1(n3949), .Y(n4182));
  NAND2X1 g3109(.A(n4178), .B(n3951), .Y(n4183));
  AOI22X1 g3110(.A0(n3953), .A1(n2374), .B0(n3950), .B1(n4171), .Y(n4184));
  NAND4X1 g3111(.A(n4183), .B(n4182), .C(n4181), .D(n4184), .Y(P1_U3250));
  XOR2X1  g3112(.A(n2321), .B(n2303), .Y(n4186));
  NAND3X1 g3113(.A(n4186), .B(n3816), .C(n3812), .Y(n4187));
  OAI21X1 g3114(.A0(n4186), .A1(n3818), .B0(n4187), .Y(n4189));
  NAND2X1 g3115(.A(n4189), .B(n3951), .Y(n4190));
  AOI22X1 g3116(.A0(P1_U3086), .A1(P1_REG3_REG_6__SCAN_IN), .B0(P1_ADDR_REG_6__SCAN_IN), .B1(n3949), .Y(n4191));
  XOR2X1  g3117(.A(n2321), .B(n3885), .Y(n4192));
  NAND3X1 g3118(.A(n4192), .B(n3906), .C(n3902), .Y(n4193));
  OAI21X1 g3119(.A0(n4192), .A1(n3908), .B0(n4193), .Y(n4195));
  NAND2X1 g3120(.A(n4195), .B(n3950), .Y(n4196));
  AOI22X1 g3121(.A0(n4189), .A1(n3858), .B0(n3857), .B1(n4195), .Y(n4197));
  OAI21X1 g3122(.A0(n3941), .A1(n2321), .B0(n4197), .Y(n4198));
  AOI22X1 g3123(.A0(n3953), .A1(n2322), .B0(n3775), .B1(n4198), .Y(n4199));
  NAND4X1 g3124(.A(n4196), .B(n4191), .C(n4190), .D(n4199), .Y(P1_U3249));
  NOR2X1  g3125(.A(n2163), .B(P1_REG2_REG_3__SCAN_IN), .Y(n4201));
  NOR2X1  g3126(.A(n2112), .B(P1_REG2_REG_2__SCAN_IN), .Y(n4202));
  NOR3X1  g3127(.A(n3803), .B(n4202), .C(n4201), .Y(n4203));
  NOR3X1  g3128(.A(n4202), .B(n2072), .C(n2051), .Y(n4204));
  NOR2X1  g3129(.A(n4204), .B(n3809), .Y(n4205));
  OAI21X1 g3130(.A0(n4205), .A1(n4201), .B0(n3808), .Y(n4206));
  NOR2X1  g3131(.A(n4206), .B(n4203), .Y(n4207));
  OAI21X1 g3132(.A0(n2265), .A1(n2247), .B0(n3800), .Y(n4208));
  AOI21X1 g3133(.A0(n4207), .A1(n3814), .B0(n4208), .Y(n4209));
  OAI22X1 g3134(.A0(n4203), .A1(n4206), .B0(n2222), .B1(P1_REG2_REG_4__SCAN_IN), .Y(n4210));
  OAI22X1 g3135(.A0(n2221), .A1(n3550), .B0(P1_REG2_REG_5__SCAN_IN), .B1(n2265), .Y(n4211));
  AOI21X1 g3136(.A0(n2265), .A1(P1_REG2_REG_5__SCAN_IN), .B0(n4211), .Y(n4212));
  AOI21X1 g3137(.A0(n4212), .A1(n4210), .B0(n4209), .Y(n4213));
  NAND2X1 g3138(.A(n4213), .B(n3951), .Y(n4214));
  AOI22X1 g3139(.A0(P1_U3086), .A1(P1_REG3_REG_5__SCAN_IN), .B0(P1_ADDR_REG_5__SCAN_IN), .B1(n3949), .Y(n4215));
  NOR2X1  g3140(.A(n2163), .B(P1_REG1_REG_3__SCAN_IN), .Y(n4216));
  NOR2X1  g3141(.A(n2112), .B(P1_REG1_REG_2__SCAN_IN), .Y(n4217));
  INVX1   g3142(.A(n3894), .Y(n4218));
  NOR3X1  g3143(.A(n4218), .B(n4217), .C(n4216), .Y(n4219));
  NOR3X1  g3144(.A(n4217), .B(n2072), .C(n3892), .Y(n4220));
  NOR2X1  g3145(.A(n4220), .B(n3899), .Y(n4221));
  OAI21X1 g3146(.A0(n4221), .A1(n4216), .B0(n3898), .Y(n4222));
  NOR2X1  g3147(.A(n4222), .B(n4219), .Y(n4223));
  OAI21X1 g3148(.A0(n2265), .A1(n3889), .B0(n3890), .Y(n4224));
  AOI21X1 g3149(.A0(n4223), .A1(n3904), .B0(n4224), .Y(n4225));
  OAI22X1 g3150(.A0(n4219), .A1(n4222), .B0(n2222), .B1(P1_REG1_REG_4__SCAN_IN), .Y(n4226));
  OAI22X1 g3151(.A0(n2221), .A1(n2200), .B0(P1_REG1_REG_5__SCAN_IN), .B1(n2265), .Y(n4227));
  AOI21X1 g3152(.A0(n2265), .A1(P1_REG1_REG_5__SCAN_IN), .B0(n4227), .Y(n4228));
  AOI21X1 g3153(.A0(n4228), .A1(n4226), .B0(n4225), .Y(n4229));
  NAND2X1 g3154(.A(n4229), .B(n3950), .Y(n4230));
  AOI22X1 g3155(.A0(n4213), .A1(n3858), .B0(n3857), .B1(n4229), .Y(n4231));
  OAI21X1 g3156(.A0(n3941), .A1(n2265), .B0(n4231), .Y(n4232));
  AOI22X1 g3157(.A0(n3953), .A1(n2266), .B0(n3775), .B1(n4232), .Y(n4233));
  NAND4X1 g3158(.A(n4230), .B(n4215), .C(n4214), .D(n4233), .Y(P1_U3248));
  NOR3X1  g3159(.A(n3946), .B(n1873), .C(P1_U3086), .Y(P1_U3973));
  INVX1   g3160(.A(P1_U3973), .Y(n4236));
  NAND2X1 g3161(.A(n2037), .B(n1987), .Y(n4237));
  OAI21X1 g3162(.A0(n1987), .A1(n1985), .B0(n4237), .Y(n4238));
  OAI21X1 g3163(.A0(n4238), .A1(n2061), .B0(n3946), .Y(n4239));
  NOR3X1  g3164(.A(n3852), .B(n2059), .C(n2034), .Y(n4240));
  AOI21X1 g3165(.A0(n4240), .A1(n4237), .B0(n1882), .Y(n4241));
  NAND3X1 g3166(.A(n1989), .B(n1985), .C(n3946), .Y(n4242));
  OAI22X1 g3167(.A0(n2011), .A1(n4242), .B0(n2004), .B1(n3946), .Y(n4243));
  AOI21X1 g3168(.A0(n4241), .A1(n2026), .B0(n4243), .Y(n4244));
  XOR2X1  g3169(.A(n4244), .B(n4239), .Y(n4245));
  INVX1   g3170(.A(n4239), .Y(n4246));
  AOI21X1 g3171(.A0(n2061), .A1(n3946), .B0(n4241), .Y(n4247));
  INVX1   g3172(.A(n4242), .Y(n4248));
  AOI22X1 g3173(.A0(n2026), .A1(n4248), .B0(n1882), .B1(P1_REG1_REG_0__SCAN_IN), .Y(n4249));
  OAI21X1 g3174(.A0(n4247), .A1(n2011), .B0(n4249), .Y(n4250));
  XOR2X1  g3175(.A(n4250), .B(n4246), .Y(n4251));
  XOR2X1  g3176(.A(n4251), .B(n4245), .Y(n4252));
  NOR2X1  g3177(.A(n2002), .B(n2080), .Y(n4253));
  NAND3X1 g3178(.A(n3858), .B(n2004), .C(P1_REG2_REG_0__SCAN_IN), .Y(n4254));
  AOI21X1 g3179(.A0(n2002), .A1(n2019), .B0(n2080), .Y(n4255));
  OAI21X1 g3180(.A0(n4255), .A1(n2004), .B0(n4254), .Y(n4256));
  AOI21X1 g3181(.A0(n4253), .A1(n4252), .B0(n4256), .Y(n4257));
  XOR2X1  g3182(.A(n2221), .B(n3550), .Y(n4258));
  NOR2X1  g3183(.A(n4258), .B(n4207), .Y(n4260));
  AOI21X1 g3184(.A0(n4258), .A1(n4207), .B0(n4260), .Y(n4261));
  AOI22X1 g3185(.A0(P1_U3086), .A1(P1_REG3_REG_4__SCAN_IN), .B0(P1_ADDR_REG_4__SCAN_IN), .B1(n3949), .Y(n4262));
  OAI21X1 g3186(.A0(n4261), .A1(n3952), .B0(n4262), .Y(n4263));
  NOR2X1  g3187(.A(n3973), .B(n2221), .Y(n4264));
  XOR2X1  g3188(.A(n2221), .B(n2200), .Y(n4265));
  NOR2X1  g3189(.A(n4265), .B(n4223), .Y(n4267));
  AOI21X1 g3190(.A0(n4265), .A1(n4223), .B0(n4267), .Y(n4268));
  OAI22X1 g3191(.A0(n4261), .A1(n3859), .B0(n2002), .B1(n4268), .Y(n4269));
  AOI21X1 g3192(.A0(n2080), .A1(n2222), .B0(n4269), .Y(n4270));
  OAI22X1 g3193(.A0(n4268), .A1(n3970), .B0(n3978), .B1(n4270), .Y(n4271));
  NOR3X1  g3194(.A(n4271), .B(n4264), .C(n4263), .Y(n4272));
  OAI21X1 g3195(.A0(n4257), .A1(n4236), .B0(n4272), .Y(P1_U3247));
  OAI21X1 g3196(.A0(n3803), .A1(n4202), .B0(n4205), .Y(n4274));
  XOR2X1  g3197(.A(n2162), .B(P1_REG2_REG_3__SCAN_IN), .Y(n4275));
  OAI21X1 g3198(.A0(n3807), .A1(n4201), .B0(n4274), .Y(n4276));
  OAI21X1 g3199(.A0(n4275), .A1(n4274), .B0(n4276), .Y(n4277));
  NAND2X1 g3200(.A(n4277), .B(n3951), .Y(n4278));
  AOI22X1 g3201(.A0(P1_U3086), .A1(P1_REG3_REG_3__SCAN_IN), .B0(P1_ADDR_REG_3__SCAN_IN), .B1(n3949), .Y(n4279));
  OAI21X1 g3202(.A0(n4218), .A1(n4217), .B0(n4221), .Y(n4280));
  XOR2X1  g3203(.A(n2162), .B(P1_REG1_REG_3__SCAN_IN), .Y(n4281));
  OAI21X1 g3204(.A0(n3897), .A1(n4216), .B0(n4280), .Y(n4282));
  OAI21X1 g3205(.A0(n4281), .A1(n4280), .B0(n4282), .Y(n4283));
  NAND2X1 g3206(.A(n4283), .B(n3950), .Y(n4284));
  AOI22X1 g3207(.A0(n4277), .A1(n3858), .B0(n3857), .B1(n4283), .Y(n4285));
  OAI21X1 g3208(.A0(n3941), .A1(n2162), .B0(n4285), .Y(n4286));
  AOI22X1 g3209(.A0(n3953), .A1(n2163), .B0(n3775), .B1(n4286), .Y(n4287));
  NAND4X1 g3210(.A(n4284), .B(n4279), .C(n4278), .D(n4287), .Y(P1_U3246));
  NOR2X1  g3211(.A(n3805), .B(n3804), .Y(n4289));
  NOR3X1  g3212(.A(n3809), .B(n4289), .C(n4202), .Y(n4290));
  XOR2X1  g3213(.A(n2111), .B(P1_REG2_REG_2__SCAN_IN), .Y(n4291));
  AOI21X1 g3214(.A0(n4291), .A1(n4289), .B0(n4290), .Y(n4292));
  NAND2X1 g3215(.A(n4292), .B(n3951), .Y(n4293));
  AOI22X1 g3216(.A0(P1_U3086), .A1(P1_REG3_REG_2__SCAN_IN), .B0(P1_ADDR_REG_2__SCAN_IN), .B1(n3949), .Y(n4294));
  NAND2X1 g3217(.A(n4294), .B(n4293), .Y(n4295));
  NOR2X1  g3218(.A(n3895), .B(n3894), .Y(n4296));
  NOR3X1  g3219(.A(n3899), .B(n4296), .C(n4217), .Y(n4297));
  XOR2X1  g3220(.A(n2111), .B(P1_REG1_REG_2__SCAN_IN), .Y(n4298));
  AOI21X1 g3221(.A0(n4298), .A1(n4296), .B0(n4297), .Y(n4299));
  NAND3X1 g3222(.A(n3855), .B(n2112), .C(n2080), .Y(n4300));
  AOI22X1 g3223(.A0(n4292), .A1(n3858), .B0(n3857), .B1(n4299), .Y(n4301));
  AOI21X1 g3224(.A0(n4301), .A1(n4300), .B0(n3978), .Y(n4302));
  AOI21X1 g3225(.A0(n4299), .A1(n3950), .B0(n4302), .Y(n4303));
  OAI21X1 g3226(.A0(n3973), .A1(n2111), .B0(n4303), .Y(n4304));
  NOR2X1  g3227(.A(n4304), .B(n4295), .Y(n4305));
  OAI21X1 g3228(.A0(n4257), .A1(n4236), .B0(n4305), .Y(P1_U3245));
  XOR2X1  g3229(.A(n2072), .B(n2051), .Y(n4307));
  XOR2X1  g3230(.A(n4307), .B(n3802), .Y(n4308));
  INVX1   g3231(.A(P1_REG3_REG_1__SCAN_IN), .Y(n4309));
  OAI22X1 g3232(.A0(P1_STATE_REG_SCAN_IN), .A1(n4309), .B0(n1133), .B1(n3954), .Y(n4310));
  AOI21X1 g3233(.A0(n4308), .A1(n3951), .B0(n4310), .Y(n4311));
  XOR2X1  g3234(.A(n2072), .B(P1_REG1_REG_1__SCAN_IN), .Y(n4312));
  XOR2X1  g3235(.A(n4312), .B(n3893), .Y(n4313));
  NAND2X1 g3236(.A(n4313), .B(n3950), .Y(n4314));
  AOI22X1 g3237(.A0(n4308), .A1(n3858), .B0(n3857), .B1(n4313), .Y(n4315));
  OAI21X1 g3238(.A0(n3941), .A1(n2072), .B0(n4315), .Y(n4316));
  AOI22X1 g3239(.A0(n3953), .A1(n2073), .B0(n3775), .B1(n4316), .Y(n4317));
  NAND3X1 g3240(.A(n4317), .B(n4314), .C(n4311), .Y(P1_U3244));
  XOR2X1  g3241(.A(n2004), .B(n2019), .Y(n4319));
  NAND2X1 g3242(.A(n4319), .B(n3951), .Y(n4320));
  AOI22X1 g3243(.A0(P1_U3086), .A1(P1_REG3_REG_0__SCAN_IN), .B0(P1_ADDR_REG_0__SCAN_IN), .B1(n3949), .Y(n4321));
  XOR2X1  g3244(.A(n2008), .B(P1_REG1_REG_0__SCAN_IN), .Y(n4322));
  NAND2X1 g3245(.A(n4322), .B(n3950), .Y(n4323));
  AOI22X1 g3246(.A0(n4319), .A1(n3858), .B0(n3857), .B1(n4322), .Y(n4324));
  OAI21X1 g3247(.A0(n3941), .A1(n2004), .B0(n4324), .Y(n4325));
  AOI22X1 g3248(.A0(n3953), .A1(n2008), .B0(n3775), .B1(n4325), .Y(n4326));
  NAND4X1 g3249(.A(n4323), .B(n4321), .C(n4320), .D(n4326), .Y(P1_U3243));
  NAND2X1 g3250(.A(n4236), .B(P1_DATAO_REG_0__SCAN_IN), .Y(n4328));
  OAI21X1 g3251(.A0(n4236), .A1(n2128), .B0(n4328), .Y(P1_U3554));
  NAND2X1 g3252(.A(n4236), .B(P1_DATAO_REG_1__SCAN_IN), .Y(n4330));
  OAI21X1 g3253(.A0(n4236), .A1(n2117), .B0(n4330), .Y(P1_U3555));
  OAI21X1 g3254(.A0(n2185), .A1(n2182), .B0(P1_U3973), .Y(n4332));
  OAI21X1 g3255(.A0(P1_U3973), .A1(n1286), .B0(n4332), .Y(P1_U3556));
  NAND2X1 g3256(.A(n4236), .B(P1_DATAO_REG_3__SCAN_IN), .Y(n4334));
  OAI21X1 g3257(.A0(n4236), .A1(n2146), .B0(n4334), .Y(P1_U3557));
  NAND2X1 g3258(.A(n4236), .B(P1_DATAO_REG_4__SCAN_IN), .Y(n4336));
  OAI21X1 g3259(.A0(n4236), .A1(n2204), .B0(n4336), .Y(P1_U3558));
  NAND2X1 g3260(.A(n4236), .B(P1_DATAO_REG_5__SCAN_IN), .Y(n4338));
  OAI21X1 g3261(.A0(n4236), .A1(n2257), .B0(n4338), .Y(P1_U3559));
  NAND2X1 g3262(.A(n4236), .B(P1_DATAO_REG_6__SCAN_IN), .Y(n4340));
  OAI21X1 g3263(.A0(n4236), .A1(n2312), .B0(n4340), .Y(P1_U3560));
  NAND2X1 g3264(.A(n4236), .B(P1_DATAO_REG_7__SCAN_IN), .Y(n4342));
  OAI21X1 g3265(.A0(n4236), .A1(n2363), .B0(n4342), .Y(P1_U3561));
  NAND2X1 g3266(.A(n4236), .B(P1_DATAO_REG_8__SCAN_IN), .Y(n4344));
  OAI21X1 g3267(.A0(n4236), .A1(n2409), .B0(n4344), .Y(P1_U3562));
  NAND2X1 g3268(.A(n4236), .B(P1_DATAO_REG_9__SCAN_IN), .Y(n4346));
  OAI21X1 g3269(.A0(n4236), .A1(n2458), .B0(n4346), .Y(P1_U3563));
  NAND2X1 g3270(.A(n4236), .B(P1_DATAO_REG_10__SCAN_IN), .Y(n4348));
  OAI21X1 g3271(.A0(n4236), .A1(n2504), .B0(n4348), .Y(P1_U3564));
  NAND2X1 g3272(.A(n4236), .B(P1_DATAO_REG_11__SCAN_IN), .Y(n4350));
  OAI21X1 g3273(.A0(n4236), .A1(n2549), .B0(n4350), .Y(P1_U3565));
  NAND2X1 g3274(.A(n4236), .B(P1_DATAO_REG_12__SCAN_IN), .Y(n4352));
  OAI21X1 g3275(.A0(n4236), .A1(n2602), .B0(n4352), .Y(P1_U3566));
  NAND2X1 g3276(.A(n4236), .B(P1_DATAO_REG_13__SCAN_IN), .Y(n4354));
  OAI21X1 g3277(.A0(n4236), .A1(n2650), .B0(n4354), .Y(P1_U3567));
  NAND2X1 g3278(.A(n4236), .B(P1_DATAO_REG_14__SCAN_IN), .Y(n4356));
  OAI21X1 g3279(.A0(n4236), .A1(n2702), .B0(n4356), .Y(P1_U3568));
  NAND2X1 g3280(.A(n4236), .B(P1_DATAO_REG_15__SCAN_IN), .Y(n4358));
  OAI21X1 g3281(.A0(n4236), .A1(n2798), .B0(n4358), .Y(P1_U3569));
  NAND2X1 g3282(.A(n4236), .B(P1_DATAO_REG_16__SCAN_IN), .Y(n4360));
  OAI21X1 g3283(.A0(n4236), .A1(n2791), .B0(n4360), .Y(P1_U3570));
  NAND2X1 g3284(.A(n4236), .B(P1_DATAO_REG_17__SCAN_IN), .Y(n4362));
  OAI21X1 g3285(.A0(n4236), .A1(n2841), .B0(n4362), .Y(P1_U3571));
  NAND2X1 g3286(.A(n4236), .B(P1_DATAO_REG_18__SCAN_IN), .Y(n4364));
  OAI21X1 g3287(.A0(n4236), .A1(n2891), .B0(n4364), .Y(P1_U3572));
  NAND2X1 g3288(.A(n4236), .B(P1_DATAO_REG_19__SCAN_IN), .Y(n4366));
  OAI21X1 g3289(.A0(n4236), .A1(n2933), .B0(n4366), .Y(P1_U3573));
  NAND2X1 g3290(.A(n4236), .B(P1_DATAO_REG_20__SCAN_IN), .Y(n4368));
  OAI21X1 g3291(.A0(n4236), .A1(n2976), .B0(n4368), .Y(P1_U3574));
  NAND2X1 g3292(.A(n4236), .B(P1_DATAO_REG_21__SCAN_IN), .Y(n4370));
  OAI21X1 g3293(.A0(n4236), .A1(n3029), .B0(n4370), .Y(P1_U3575));
  NAND2X1 g3294(.A(n4236), .B(P1_DATAO_REG_22__SCAN_IN), .Y(n4372));
  OAI21X1 g3295(.A0(n4236), .A1(n3071), .B0(n4372), .Y(P1_U3576));
  NAND2X1 g3296(.A(n4236), .B(P1_DATAO_REG_23__SCAN_IN), .Y(n4374));
  OAI21X1 g3297(.A0(n4236), .A1(n3110), .B0(n4374), .Y(P1_U3577));
  NAND2X1 g3298(.A(n4236), .B(P1_DATAO_REG_24__SCAN_IN), .Y(n4376));
  OAI21X1 g3299(.A0(n4236), .A1(n3150), .B0(n4376), .Y(P1_U3578));
  NAND2X1 g3300(.A(n4236), .B(P1_DATAO_REG_25__SCAN_IN), .Y(n4378));
  OAI21X1 g3301(.A0(n4236), .A1(n3192), .B0(n4378), .Y(P1_U3579));
  NAND2X1 g3302(.A(n4236), .B(P1_DATAO_REG_26__SCAN_IN), .Y(n4380));
  OAI21X1 g3303(.A0(n4236), .A1(n3236), .B0(n4380), .Y(P1_U3580));
  NAND2X1 g3304(.A(n4236), .B(P1_DATAO_REG_27__SCAN_IN), .Y(n4382));
  OAI21X1 g3305(.A0(n4236), .A1(n3282), .B0(n4382), .Y(P1_U3581));
  NAND2X1 g3306(.A(n4236), .B(P1_DATAO_REG_28__SCAN_IN), .Y(n4384));
  OAI21X1 g3307(.A0(n4236), .A1(n3322), .B0(n4384), .Y(P1_U3582));
  NAND2X1 g3308(.A(n4236), .B(P1_DATAO_REG_29__SCAN_IN), .Y(n4386));
  OAI21X1 g3309(.A0(n4236), .A1(n3364), .B0(n4386), .Y(P1_U3583));
  NAND2X1 g3310(.A(n4236), .B(P1_DATAO_REG_30__SCAN_IN), .Y(n4388));
  OAI21X1 g3311(.A0(n4236), .A1(n3384), .B0(n4388), .Y(P1_U3584));
  NAND2X1 g3312(.A(n3425), .B(n3424), .Y(n4390));
  INVX1   g3313(.A(n4390), .Y(n4391));
  NAND2X1 g3314(.A(n4236), .B(P1_DATAO_REG_31__SCAN_IN), .Y(n4392));
  OAI21X1 g3315(.A0(n4236), .A1(n4391), .B0(n4392), .Y(P1_U3585));
  NAND2X1 g3316(.A(n3769), .B(n4391), .Y(n4394));
  NOR4X1  g3317(.A(n3295), .B(n3302), .C(n3246), .D(n3393), .Y(n4395));
  OAI21X1 g3318(.A0(n3433), .A1(n4390), .B0(n4395), .Y(n4396));
  NOR4X1  g3319(.A(n3124), .B(n3078), .C(n3071), .D(n3169), .Y(n4397));
  NOR3X1  g3320(.A(n3169), .B(n3142), .C(n3110), .Y(n4398));
  NOR4X1  g3321(.A(n4397), .B(n3247), .C(n3170), .D(n4398), .Y(n4399));
  NAND3X1 g3322(.A(n4399), .B(n3406), .C(n3308), .Y(n4400));
  NOR2X1  g3323(.A(n3393), .B(n3334), .Y(n4401));
  OAI21X1 g3324(.A0(n3433), .A1(n4390), .B0(n4401), .Y(n4402));
  NOR4X1  g3325(.A(n3295), .B(n3273), .C(n3235), .D(n3393), .Y(n4403));
  OAI22X1 g3326(.A0(n3433), .A1(n4390), .B0(n3404), .B1(n4403), .Y(n4404));
  NAND4X1 g3327(.A(n4402), .B(n4400), .C(n4396), .D(n4404), .Y(n4405));
  AOI22X1 g3328(.A0(n3383), .A1(n3423), .B0(n3401), .B1(n3363), .Y(n4406));
  NAND2X1 g3329(.A(n4406), .B(n4405), .Y(n4407));
  NOR3X1  g3330(.A(n3363), .B(n2003), .C(n1820), .Y(n4408));
  NAND2X1 g3331(.A(n3423), .B(n3383), .Y(n4409));
  NAND2X1 g3332(.A(n4409), .B(n4408), .Y(n4410));
  NOR2X1  g3333(.A(n3423), .B(n3383), .Y(n4411));
  NAND2X1 g3334(.A(n4411), .B(n4394), .Y(n4412));
  NAND2X1 g3335(.A(n3433), .B(n4390), .Y(n4413));
  NAND4X1 g3336(.A(n4412), .B(n4410), .C(n4407), .D(n4413), .Y(n4414));
  OAI21X1 g3337(.A0(n3433), .A1(n4390), .B0(n3404), .Y(n4415));
  AOI22X1 g3338(.A0(n4401), .A1(n4394), .B0(n4408), .B1(n4409), .Y(n4416));
  NAND3X1 g3339(.A(n3406), .B(n3308), .C(n3305), .Y(n4417));
  AOI21X1 g3340(.A0(n3769), .A1(n4391), .B0(n4417), .Y(n4418));
  NOR2X1  g3341(.A(n3769), .B(n4391), .Y(n4419));
  INVX1   g3342(.A(n2763), .Y(n4420));
  NOR3X1  g3343(.A(n2529), .B(n2432), .C(n2330), .Y(n4421));
  OAI21X1 g3344(.A0(n2424), .A1(n2409), .B0(n4421), .Y(n4422));
  INVX1   g3345(.A(n2290), .Y(n4423));
  NOR2X1  g3346(.A(n2128), .B(n2010), .Y(n4424));
  AOI21X1 g3347(.A0(n2084), .A1(n1987), .B0(n4424), .Y(n4425));
  AOI21X1 g3348(.A0(n4425), .A1(n2075), .B0(n2117), .Y(n4426));
  NOR2X1  g3349(.A(n4425), .B(n2075), .Y(n4427));
  OAI22X1 g3350(.A0(n2146), .A1(n2169), .B0(n2114), .B1(n2103), .Y(n4428));
  NOR4X1  g3351(.A(n4427), .B(n4426), .C(n2272), .D(n4428), .Y(n4429));
  OAI21X1 g3352(.A0(n2329), .A1(n4423), .B0(n4429), .Y(n4430));
  AOI22X1 g3353(.A0(n2504), .A1(n2516), .B0(n2469), .B1(n2458), .Y(n4431));
  OAI21X1 g3354(.A0(n4430), .A1(n4422), .B0(n4431), .Y(n4432));
  NAND2X1 g3355(.A(n2424), .B(n2409), .Y(n4433));
  OAI21X1 g3356(.A0(n2424), .A1(n2409), .B0(n2431), .Y(n4434));
  AOI21X1 g3357(.A0(n4434), .A1(n4433), .B0(n2529), .Y(n4435));
  AOI22X1 g3358(.A0(n2602), .A1(n2614), .B0(n2562), .B1(n2549), .Y(n4436));
  OAI21X1 g3359(.A0(n2169), .A1(n2146), .B0(n2186), .Y(n4437));
  AOI21X1 g3360(.A0(n4437), .A1(n2234), .B0(n2272), .Y(n4438));
  OAI22X1 g3361(.A0(n2388), .A1(n4438), .B0(n2329), .B1(n4423), .Y(n4439));
  OAI21X1 g3362(.A0(n4439), .A1(n4422), .B0(n4436), .Y(n4440));
  NOR3X1  g3363(.A(n4440), .B(n4435), .C(n4432), .Y(n4441));
  NAND2X1 g3364(.A(n4436), .B(n2556), .Y(n4442));
  NAND2X1 g3365(.A(n2988), .B(n2570), .Y(n4443));
  NAND4X1 g3366(.A(n4442), .B(n2717), .C(n2987), .D(n4443), .Y(n4444));
  OAI22X1 g3367(.A0(n4441), .A1(n4444), .B0(n2671), .B1(n2649), .Y(n4445));
  AOI21X1 g3368(.A0(n4445), .A1(n4420), .B0(n2761), .Y(n4446));
  NOR2X1  g3369(.A(n2907), .B(n2902), .Y(n4447));
  NOR4X1  g3370(.A(n2861), .B(n2810), .C(n2801), .D(n4447), .Y(n4448));
  OAI21X1 g3371(.A0(n4446), .A1(n2799), .B0(n4448), .Y(n4449));
  NOR2X1  g3372(.A(n2925), .B(n2891), .Y(n4450));
  NOR4X1  g3373(.A(n2861), .B(n2811), .C(n2791), .D(n4447), .Y(n4451));
  NOR3X1  g3374(.A(n4447), .B(n2854), .C(n2841), .Y(n4452));
  NOR4X1  g3375(.A(n4451), .B(n2986), .C(n4450), .D(n4452), .Y(n4453));
  AOI21X1 g3376(.A0(n4453), .A1(n4449), .B0(n3039), .Y(n4454));
  NOR3X1  g3377(.A(n4454), .B(n3051), .C(n3008), .Y(n4455));
  OAI21X1 g3378(.A0(n3051), .A1(n3038), .B0(n3080), .Y(n4456));
  NOR3X1  g3379(.A(n4456), .B(n4455), .C(n3118), .Y(n4457));
  NAND3X1 g3380(.A(n4457), .B(n3201), .C(n3159), .Y(n4458));
  NOR3X1  g3381(.A(n4458), .B(n4419), .C(n4418), .Y(n4459));
  OAI21X1 g3382(.A0(n4411), .A1(n4395), .B0(n4394), .Y(n4460));
  NAND4X1 g3383(.A(n4459), .B(n4416), .C(n4415), .D(n4460), .Y(n4461));
  NAND2X1 g3384(.A(n1991), .B(n1873), .Y(n4462));
  NOR2X1  g3385(.A(n4462), .B(n2028), .Y(n4463));
  NAND4X1 g3386(.A(n4461), .B(n4414), .C(n4394), .D(n4463), .Y(n4464));
  NAND3X1 g3387(.A(n4413), .B(n4412), .C(n4410), .Y(n4465));
  AOI21X1 g3388(.A0(n4406), .A1(n4405), .B0(n4465), .Y(n4466));
  NAND2X1 g3389(.A(n4461), .B(n4394), .Y(n4467));
  NOR3X1  g3390(.A(n1991), .B(n2028), .C(n1872), .Y(n4468));
  OAI21X1 g3391(.A0(n4467), .A1(n4466), .B0(n4468), .Y(n4469));
  NAND2X1 g3392(.A(n4469), .B(n4464), .Y(n4470));
  NOR3X1  g3393(.A(n1992), .B(n1987), .C(n1982), .Y(n4471));
  AOI21X1 g3394(.A0(n4471), .A1(n3858), .B0(n1873), .Y(n4472));
  NOR2X1  g3395(.A(n1982), .B(n1872), .Y(n4473));
  NOR2X1  g3396(.A(n4473), .B(P1_U3086), .Y(n4474));
  OAI21X1 g3397(.A0(n3946), .A1(n1873), .B0(n4474), .Y(n4475));
  OAI21X1 g3398(.A0(n4475), .A1(n4472), .B0(P1_B_REG_SCAN_IN), .Y(n4476));
  INVX1   g3399(.A(n2060), .Y(n4477));
  OAI21X1 g3400(.A0(n1991), .A1(n1983), .B0(n1873), .Y(n4478));
  OAI22X1 g3401(.A0(n4478), .A1(n4391), .B0(n3433), .B1(n4477), .Y(n4482));
  OAI22X1 g3402(.A0(n4478), .A1(n3433), .B0(n4477), .B1(n4391), .Y(n4483));
  XOR2X1  g3403(.A(n4483), .B(n4482), .Y(n4484));
  NAND3X1 g3404(.A(n4390), .B(n3383), .C(n2060), .Y(n4485));
  INVX1   g3405(.A(n4478), .Y(n4486));
  NAND3X1 g3406(.A(n4486), .B(n3119), .C(n3759), .Y(n4487));
  NAND2X1 g3407(.A(n4390), .B(n3383), .Y(n4488));
  OAI22X1 g3408(.A0(n4478), .A1(n4488), .B0(n3423), .B1(n4477), .Y(n4489));
  AOI21X1 g3409(.A0(n4487), .A1(n4485), .B0(n4489), .Y(n4490));
  NAND2X1 g3410(.A(n4486), .B(n3371), .Y(n4491));
  AOI22X1 g3411(.A0(n3397), .A1(n1872), .B0(n2060), .B1(n3363), .Y(n4492));
  AOI21X1 g3412(.A0(n4486), .A1(n3363), .B0(n1872), .Y(n4493));
  OAI21X1 g3413(.A0(n3401), .A1(n4477), .B0(n4493), .Y(n4494));
  AOI21X1 g3414(.A0(n4492), .A1(n4491), .B0(n4494), .Y(n4495));
  NOR3X1  g3415(.A(n4478), .B(n2003), .C(n1790), .Y(n4496));
  OAI22X1 g3416(.A0(n3282), .A1(n1873), .B0(n4477), .B1(n3322), .Y(n4497));
  OAI21X1 g3417(.A0(n4478), .A1(n3322), .B0(n1873), .Y(n4498));
  AOI21X1 g3418(.A0(n3329), .A1(n2060), .B0(n4498), .Y(n4499));
  OAI21X1 g3419(.A0(n4497), .A1(n4496), .B0(n4499), .Y(n4500));
  NOR3X1  g3420(.A(n4499), .B(n4497), .C(n4496), .Y(n4501));
  AOI22X1 g3421(.A0(n3235), .A1(n1872), .B0(n2060), .B1(n3281), .Y(n4502));
  OAI21X1 g3422(.A0(n4478), .A1(n3294), .B0(n4502), .Y(n4503));
  OAI21X1 g3423(.A0(n4478), .A1(n3282), .B0(n1873), .Y(n4504));
  AOI21X1 g3424(.A0(n3333), .A1(n2060), .B0(n4504), .Y(n4505));
  NOR2X1  g3425(.A(n4505), .B(n4503), .Y(n4506));
  OAI21X1 g3426(.A0(n4506), .A1(n4501), .B0(n4500), .Y(n4507));
  NOR4X1  g3427(.A(n4495), .B(n4490), .C(n4484), .D(n4507), .Y(n4508));
  AOI22X1 g3428(.A0(n4486), .A1(n4390), .B0(n3769), .B1(n2060), .Y(n4509));
  NOR4X1  g3429(.A(n4509), .B(n2060), .C(n1873), .D(n4483), .Y(n4510));
  AOI22X1 g3430(.A0(n4486), .A1(n3769), .B0(n2060), .B1(n4390), .Y(n4511));
  AOI21X1 g3431(.A0(n2037), .A1(n1982), .B0(n1873), .Y(n4512));
  NOR3X1  g3432(.A(n4512), .B(n4511), .C(n4482), .Y(n4513));
  NOR3X1  g3433(.A(n4513), .B(n4510), .C(n4508), .Y(n4514));
  NAND2X1 g3434(.A(n4505), .B(n4503), .Y(n4515));
  AOI21X1 g3435(.A0(n4486), .A1(n3191), .B0(n1872), .Y(n4516));
  OAI21X1 g3436(.A0(n3215), .A1(n4477), .B0(n4516), .Y(n4517));
  OAI22X1 g3437(.A0(n3150), .A1(n1873), .B0(n4477), .B1(n3192), .Y(n4518));
  AOI21X1 g3438(.A0(n4486), .A1(n3199), .B0(n4518), .Y(n4519));
  NAND2X1 g3439(.A(n4519), .B(n4517), .Y(n4520));
  AOI21X1 g3440(.A0(n4486), .A1(n3235), .B0(n1872), .Y(n4521));
  INVX1   g3441(.A(n4521), .Y(n4522));
  AOI21X1 g3442(.A0(n3243), .A1(n2060), .B0(n4522), .Y(n4523));
  AOI22X1 g3443(.A0(n3191), .A1(n1872), .B0(n2060), .B1(n3235), .Y(n4524));
  OAI21X1 g3444(.A0(n4478), .A1(n3273), .B0(n4524), .Y(n4525));
  OAI21X1 g3445(.A0(n4525), .A1(n4523), .B0(n4520), .Y(n4526));
  NAND2X1 g3446(.A(n4525), .B(n4523), .Y(n4527));
  NAND4X1 g3447(.A(n4526), .B(n4515), .C(n4500), .D(n4527), .Y(n4528));
  NOR4X1  g3448(.A(n4495), .B(n4490), .C(n4484), .D(n4528), .Y(n4529));
  OAI21X1 g3449(.A0(n4478), .A1(n3150), .B0(n1873), .Y(n4530));
  AOI21X1 g3450(.A0(n3157), .A1(n2060), .B0(n4530), .Y(n4531));
  AOI22X1 g3451(.A0(n3109), .A1(n1872), .B0(n2060), .B1(n3149), .Y(n4532));
  OAI21X1 g3452(.A0(n4478), .A1(n3175), .B0(n4532), .Y(n4533));
  OAI21X1 g3453(.A0(n4478), .A1(n3110), .B0(n1873), .Y(n4534));
  AOI21X1 g3454(.A0(n3142), .A1(n2060), .B0(n4534), .Y(n4535));
  AOI22X1 g3455(.A0(n3070), .A1(n1872), .B0(n2060), .B1(n3109), .Y(n4536));
  OAI21X1 g3456(.A0(n4478), .A1(n3120), .B0(n4536), .Y(n4537));
  OAI22X1 g3457(.A0(n4535), .A1(n4537), .B0(n4533), .B1(n4531), .Y(n4538));
  AOI21X1 g3458(.A0(n4486), .A1(n3001), .B0(n1872), .Y(n4539));
  OAI21X1 g3459(.A0(n3021), .A1(n4477), .B0(n4539), .Y(n4540));
  OAI22X1 g3460(.A0(n2933), .A1(n1873), .B0(n4477), .B1(n2976), .Y(n4541));
  AOI21X1 g3461(.A0(n4486), .A1(n2983), .B0(n4541), .Y(n4542));
  NAND2X1 g3462(.A(n4542), .B(n4540), .Y(n4543));
  OAI21X1 g3463(.A0(n4478), .A1(n2933), .B0(n1873), .Y(n4544));
  AOI21X1 g3464(.A0(n2941), .A1(n2060), .B0(n4544), .Y(n4545));
  AOI22X1 g3465(.A0(n2902), .A1(n1872), .B0(n2060), .B1(n3002), .Y(n4546));
  OAI21X1 g3466(.A0(n4478), .A1(n2966), .B0(n4546), .Y(n4547));
  NOR2X1  g3467(.A(n4547), .B(n4545), .Y(n4548));
  OAI21X1 g3468(.A0(n4478), .A1(n2702), .B0(n1873), .Y(n4549));
  AOI21X1 g3469(.A0(n2741), .A1(n2060), .B0(n4549), .Y(n4550));
  AOI22X1 g3470(.A0(n2649), .A1(n1872), .B0(n2060), .B1(n2709), .Y(n4551));
  OAI21X1 g3471(.A0(n4478), .A1(n2714), .B0(n4551), .Y(n4552));
  NOR2X1  g3472(.A(n4552), .B(n4550), .Y(n4553));
  OAI21X1 g3473(.A0(n4478), .A1(n2650), .B0(n1873), .Y(n4554));
  AOI21X1 g3474(.A0(n2665), .A1(n2060), .B0(n4554), .Y(n4555));
  AOI22X1 g3475(.A0(n2634), .A1(n1872), .B0(n2060), .B1(n2649), .Y(n4556));
  OAI21X1 g3476(.A0(n4478), .A1(n2671), .B0(n4556), .Y(n4557));
  NOR2X1  g3477(.A(n4557), .B(n4555), .Y(n4558));
  OAI21X1 g3478(.A0(n2203), .A1(n2199), .B0(n4486), .Y(n4559));
  AOI21X1 g3479(.A0(n2224), .A1(n2060), .B0(n1872), .Y(n4560));
  NAND2X1 g3480(.A(n4560), .B(n4559), .Y(n4561));
  OAI21X1 g3481(.A0(n2203), .A1(n2199), .B0(n2060), .Y(n4562));
  AOI22X1 g3482(.A0(n2224), .A1(n4486), .B0(n2160), .B1(n1872), .Y(n4563));
  NAND3X1 g3483(.A(n4563), .B(n4562), .C(n4561), .Y(n4564));
  OAI21X1 g3484(.A0(n2145), .A1(n2141), .B0(n4486), .Y(n4565));
  AOI21X1 g3485(.A0(n2169), .A1(n2060), .B0(n1872), .Y(n4566));
  OAI21X1 g3486(.A0(n2145), .A1(n2141), .B0(n2060), .Y(n4567));
  AOI22X1 g3487(.A0(n2169), .A1(n4486), .B0(n2102), .B1(n1872), .Y(n4568));
  NAND2X1 g3488(.A(n4568), .B(n4567), .Y(n4569));
  AOI21X1 g3489(.A0(n4566), .A1(n4565), .B0(n4569), .Y(n4570));
  OAI21X1 g3490(.A0(n2185), .A1(n2182), .B0(n4486), .Y(n4571));
  AOI21X1 g3491(.A0(n2114), .A1(n2060), .B0(n1872), .Y(n4572));
  NAND2X1 g3492(.A(n4572), .B(n4571), .Y(n4573));
  OAI21X1 g3493(.A0(n2185), .A1(n2182), .B0(n2060), .Y(n4574));
  AOI22X1 g3494(.A0(n2114), .A1(n4486), .B0(n2058), .B1(n1872), .Y(n4575));
  NAND3X1 g3495(.A(n4575), .B(n4574), .C(n4573), .Y(n4576));
  NAND2X1 g3496(.A(n4575), .B(n4574), .Y(n4577));
  NAND3X1 g3497(.A(n4577), .B(n4572), .C(n4571), .Y(n4578));
  AOI21X1 g3498(.A0(n2075), .A1(n2060), .B0(n1872), .Y(n4580));
  OAI21X1 g3499(.A0(n2117), .A1(n4478), .B0(n4580), .Y(n4581));
  OAI22X1 g3500(.A0(n2093), .A1(n4478), .B0(n2128), .B1(n1873), .Y(n4583));
  AOI21X1 g3501(.A0(n2058), .A1(n2060), .B0(n4583), .Y(n4584));
  NAND3X1 g3502(.A(n4584), .B(n4581), .C(n4578), .Y(n4585));
  NAND2X1 g3503(.A(n4566), .B(n4565), .Y(n4586));
  AOI21X1 g3504(.A0(n4568), .A1(n4567), .B0(n4586), .Y(n4587));
  AOI21X1 g3505(.A0(n4585), .A1(n4576), .B0(n4587), .Y(n4588));
  AOI21X1 g3506(.A0(n4563), .A1(n4562), .B0(n4561), .Y(n4589));
  INVX1   g3507(.A(n4589), .Y(n4590));
  OAI21X1 g3508(.A0(n4588), .A1(n4570), .B0(n4590), .Y(n4591));
  NAND2X1 g3509(.A(n4486), .B(n2268), .Y(n4592));
  NAND2X1 g3510(.A(n2095), .B(P1_REG2_REG_5__SCAN_IN), .Y(n4593));
  NAND4X1 g3511(.A(n2251), .B(n2249), .C(n4593), .D(n2255), .Y(n4594));
  AOI22X1 g3512(.A0(n2219), .A1(n1872), .B0(n2060), .B1(n4594), .Y(n4595));
  AOI21X1 g3513(.A0(n4594), .A1(n4486), .B0(n1872), .Y(n4596));
  OAI21X1 g3514(.A0(n2283), .A1(n4477), .B0(n4596), .Y(n4597));
  AOI21X1 g3515(.A0(n4595), .A1(n4592), .B0(n4597), .Y(n4598));
  AOI21X1 g3516(.A0(n4591), .A1(n4564), .B0(n4598), .Y(n4599));
  OAI21X1 g3517(.A0(n4584), .A1(n4581), .B0(n4578), .Y(n4600));
  OAI22X1 g3518(.A0(n4477), .A1(n2128), .B0(n2011), .B1(n4478), .Y(n4601));
  NOR2X1  g3519(.A(n4478), .B(n2128), .Y(n4602));
  OAI21X1 g3520(.A0(n4477), .A1(n2011), .B0(n1873), .Y(n4603));
  NOR2X1  g3521(.A(n4603), .B(n4602), .Y(n4604));
  NOR3X1  g3522(.A(n1991), .B(n1983), .C(n1872), .Y(n4605));
  OAI21X1 g3523(.A0(n4605), .A1(n4604), .B0(n4601), .Y(n4606));
  AOI21X1 g3524(.A0(n4605), .A1(n4604), .B0(n4587), .Y(n4607));
  NAND2X1 g3525(.A(n4607), .B(n4606), .Y(n4608));
  NOR4X1  g3526(.A(n4600), .B(n4598), .C(n4589), .D(n4608), .Y(n4609));
  AOI22X1 g3527(.A0(n4594), .A1(n1872), .B0(n2060), .B1(n2313), .Y(n4610));
  OAI21X1 g3528(.A0(n4478), .A1(n2355), .B0(n4610), .Y(n4611));
  OAI21X1 g3529(.A0(n4478), .A1(n2312), .B0(n1873), .Y(n4612));
  AOI21X1 g3530(.A0(n2324), .A1(n2060), .B0(n4612), .Y(n4613));
  NAND3X1 g3531(.A(n4597), .B(n4595), .C(n4592), .Y(n4614));
  OAI21X1 g3532(.A0(n4613), .A1(n4611), .B0(n4614), .Y(n4615));
  NOR3X1  g3533(.A(n4615), .B(n4609), .C(n4599), .Y(n4616));
  AOI22X1 g3534(.A0(n2408), .A1(n1872), .B0(n2060), .B1(n2457), .Y(n4617));
  OAI21X1 g3535(.A0(n4478), .A1(n2496), .B0(n4617), .Y(n4618));
  OAI21X1 g3536(.A0(n4478), .A1(n2458), .B0(n1873), .Y(n4619));
  AOI21X1 g3537(.A0(n2469), .A1(n2060), .B0(n4619), .Y(n4620));
  NAND2X1 g3538(.A(n4620), .B(n4618), .Y(n4621));
  AOI22X1 g3539(.A0(n2362), .A1(n1872), .B0(n2060), .B1(n2408), .Y(n4622));
  OAI21X1 g3540(.A0(n4478), .A1(n2447), .B0(n4622), .Y(n4623));
  AOI21X1 g3541(.A0(n4486), .A1(n2408), .B0(n1872), .Y(n4624));
  INVX1   g3542(.A(n4624), .Y(n4625));
  AOI21X1 g3543(.A0(n2424), .A1(n2060), .B0(n4625), .Y(n4626));
  NAND2X1 g3544(.A(n4626), .B(n4623), .Y(n4627));
  AOI22X1 g3545(.A0(n2313), .A1(n1872), .B0(n2060), .B1(n2362), .Y(n4628));
  OAI21X1 g3546(.A0(n4478), .A1(n2399), .B0(n4628), .Y(n4629));
  OAI21X1 g3547(.A0(n4478), .A1(n2363), .B0(n1873), .Y(n4630));
  AOI21X1 g3548(.A0(n2376), .A1(n2060), .B0(n4630), .Y(n4631));
  AOI22X1 g3549(.A0(n4629), .A1(n4631), .B0(n4613), .B1(n4611), .Y(n4632));
  NAND3X1 g3550(.A(n4632), .B(n4627), .C(n4621), .Y(n4633));
  OAI21X1 g3551(.A0(n4478), .A1(n2602), .B0(n1873), .Y(n4634));
  AOI21X1 g3552(.A0(n2614), .A1(n2060), .B0(n4634), .Y(n4635));
  AOI22X1 g3553(.A0(n2580), .A1(n1872), .B0(n2060), .B1(n2634), .Y(n4636));
  OAI21X1 g3554(.A0(n4478), .A1(n2642), .B0(n4636), .Y(n4637));
  OAI21X1 g3555(.A0(n4478), .A1(n2549), .B0(n1873), .Y(n4638));
  AOI21X1 g3556(.A0(n2562), .A1(n2060), .B0(n4638), .Y(n4639));
  AOI22X1 g3557(.A0(n2503), .A1(n1872), .B0(n2060), .B1(n2580), .Y(n4640));
  OAI21X1 g3558(.A0(n4478), .A1(n2593), .B0(n4640), .Y(n4641));
  OAI22X1 g3559(.A0(n4639), .A1(n4641), .B0(n4637), .B1(n4635), .Y(n4642));
  NOR2X1  g3560(.A(n4631), .B(n4629), .Y(n4643));
  NAND3X1 g3561(.A(n4643), .B(n4627), .C(n4621), .Y(n4644));
  NOR2X1  g3562(.A(n4626), .B(n4623), .Y(n4645));
  NAND2X1 g3563(.A(n4645), .B(n4621), .Y(n4646));
  OAI21X1 g3564(.A0(n4478), .A1(n2504), .B0(n1873), .Y(n4647));
  AOI21X1 g3565(.A0(n2516), .A1(n2060), .B0(n4647), .Y(n4648));
  INVX1   g3566(.A(n4648), .Y(n4649));
  AOI22X1 g3567(.A0(n2457), .A1(n1872), .B0(n2060), .B1(n2503), .Y(n4650));
  INVX1   g3568(.A(n4650), .Y(n4651));
  AOI21X1 g3569(.A0(n4486), .A1(n2516), .B0(n4651), .Y(n4652));
  NOR2X1  g3570(.A(n4620), .B(n4618), .Y(n4653));
  AOI21X1 g3571(.A0(n4652), .A1(n4649), .B0(n4653), .Y(n4654));
  NAND3X1 g3572(.A(n4654), .B(n4646), .C(n4644), .Y(n4655));
  NOR2X1  g3573(.A(n4655), .B(n4642), .Y(n4656));
  OAI21X1 g3574(.A0(n4633), .A1(n4616), .B0(n4656), .Y(n4657));
  NOR3X1  g3575(.A(n4652), .B(n4649), .C(n4642), .Y(n4658));
  NOR2X1  g3576(.A(n4637), .B(n4635), .Y(n4659));
  NAND2X1 g3577(.A(n4641), .B(n4639), .Y(n4660));
  AOI22X1 g3578(.A0(n4635), .A1(n4637), .B0(n4557), .B1(n4555), .Y(n4661));
  OAI21X1 g3579(.A0(n4660), .A1(n4659), .B0(n4661), .Y(n4662));
  NOR2X1  g3580(.A(n4662), .B(n4658), .Y(n4663));
  AOI21X1 g3581(.A0(n4663), .A1(n4657), .B0(n4558), .Y(n4664));
  AOI21X1 g3582(.A0(n4552), .A1(n4550), .B0(n4664), .Y(n4665));
  AOI22X1 g3583(.A0(n2709), .A1(n1872), .B0(n2060), .B1(n2749), .Y(n4666));
  OAI21X1 g3584(.A0(n4478), .A1(n2759), .B0(n4666), .Y(n4667));
  AOI21X1 g3585(.A0(n4486), .A1(n2749), .B0(n1872), .Y(n4668));
  OAI21X1 g3586(.A0(n2759), .A1(n4477), .B0(n4668), .Y(n4669));
  INVX1   g3587(.A(n4669), .Y(n4670));
  NAND2X1 g3588(.A(n4670), .B(n4667), .Y(n4671));
  OAI21X1 g3589(.A0(n4665), .A1(n4553), .B0(n4671), .Y(n4672));
  AOI21X1 g3590(.A0(n4486), .A1(n2902), .B0(n1872), .Y(n4673));
  OAI21X1 g3591(.A0(n2907), .A1(n4477), .B0(n4673), .Y(n4674));
  OAI22X1 g3592(.A0(n2841), .A1(n1873), .B0(n4477), .B1(n2891), .Y(n4675));
  AOI21X1 g3593(.A0(n4486), .A1(n2925), .B0(n4675), .Y(n4676));
  NAND2X1 g3594(.A(n4676), .B(n4674), .Y(n4677));
  AOI21X1 g3595(.A0(n4486), .A1(n2840), .B0(n1872), .Y(n4678));
  OAI21X1 g3596(.A0(n2853), .A1(n4477), .B0(n4678), .Y(n4679));
  AOI22X1 g3597(.A0(n2792), .A1(n1872), .B0(n2060), .B1(n2840), .Y(n4680));
  INVX1   g3598(.A(n4680), .Y(n4681));
  AOI21X1 g3599(.A0(n4486), .A1(n2854), .B0(n4681), .Y(n4682));
  NAND2X1 g3600(.A(n4682), .B(n4679), .Y(n4683));
  NAND2X1 g3601(.A(n4683), .B(n4677), .Y(n4684));
  OAI21X1 g3602(.A0(n4478), .A1(n2791), .B0(n1873), .Y(n4685));
  AOI21X1 g3603(.A0(n2811), .A1(n2060), .B0(n4685), .Y(n4686));
  AOI22X1 g3604(.A0(n2749), .A1(n1872), .B0(n2060), .B1(n2792), .Y(n4687));
  OAI21X1 g3605(.A0(n4478), .A1(n2806), .B0(n4687), .Y(n4688));
  OAI22X1 g3606(.A0(n4686), .A1(n4688), .B0(n4670), .B1(n4667), .Y(n4689));
  NOR2X1  g3607(.A(n4689), .B(n4684), .Y(n4690));
  NAND4X1 g3608(.A(n4686), .B(n4683), .C(n4677), .D(n4688), .Y(n4691));
  NAND2X1 g3609(.A(n4547), .B(n4545), .Y(n4692));
  NOR2X1  g3610(.A(n4676), .B(n4674), .Y(n4693));
  NOR2X1  g3611(.A(n4682), .B(n4679), .Y(n4694));
  AOI21X1 g3612(.A0(n4694), .A1(n4677), .B0(n4693), .Y(n4695));
  NAND3X1 g3613(.A(n4695), .B(n4692), .C(n4691), .Y(n4696));
  AOI21X1 g3614(.A0(n4690), .A1(n4672), .B0(n4696), .Y(n4697));
  OAI22X1 g3615(.A0(n4548), .A1(n4697), .B0(n4542), .B1(n4540), .Y(n4698));
  OAI21X1 g3616(.A0(n4478), .A1(n3029), .B0(n1873), .Y(n4699));
  AOI21X1 g3617(.A0(n3036), .A1(n2060), .B0(n4699), .Y(n4700));
  AOI22X1 g3618(.A0(n3001), .A1(n1872), .B0(n2060), .B1(n3028), .Y(n4701));
  OAI21X1 g3619(.A0(n4478), .A1(n3063), .B0(n4701), .Y(n4702));
  AOI22X1 g3620(.A0(n4700), .A1(n4702), .B0(n4698), .B1(n4543), .Y(n4703));
  AOI21X1 g3621(.A0(n4486), .A1(n3070), .B0(n1872), .Y(n4704));
  INVX1   g3622(.A(n4704), .Y(n4705));
  AOI21X1 g3623(.A0(n3078), .A1(n2060), .B0(n4705), .Y(n4706));
  AOI22X1 g3624(.A0(n3028), .A1(n1872), .B0(n2060), .B1(n3070), .Y(n4707));
  OAI21X1 g3625(.A0(n4478), .A1(n3102), .B0(n4707), .Y(n4708));
  OAI22X1 g3626(.A0(n4706), .A1(n4708), .B0(n4702), .B1(n4700), .Y(n4709));
  NOR3X1  g3627(.A(n4709), .B(n4703), .C(n4538), .Y(n4710));
  NOR2X1  g3628(.A(n4533), .B(n4531), .Y(n4711));
  NAND2X1 g3629(.A(n4533), .B(n4531), .Y(n4712));
  NAND2X1 g3630(.A(n4537), .B(n4535), .Y(n4713));
  OAI21X1 g3631(.A0(n4713), .A1(n4711), .B0(n4712), .Y(n4714));
  NAND2X1 g3632(.A(n4708), .B(n4706), .Y(n4715));
  OAI22X1 g3633(.A0(n4538), .A1(n4715), .B0(n4519), .B1(n4517), .Y(n4716));
  NOR3X1  g3634(.A(n4716), .B(n4714), .C(n4710), .Y(n4717));
  NAND4X1 g3635(.A(n4527), .B(n4515), .C(n4500), .D(n4717), .Y(n4718));
  NOR4X1  g3636(.A(n4495), .B(n4490), .C(n4484), .D(n4718), .Y(n4719));
  NAND3X1 g3637(.A(n4489), .B(n4487), .C(n4485), .Y(n4720));
  NOR2X1  g3638(.A(n4720), .B(n4484), .Y(n4721));
  NAND3X1 g3639(.A(n4494), .B(n4492), .C(n4491), .Y(n4722));
  NOR3X1  g3640(.A(n4722), .B(n4490), .C(n4484), .Y(n4723));
  NOR4X1  g3641(.A(n4721), .B(n4719), .C(n4529), .D(n4723), .Y(n4724));
  NAND2X1 g3642(.A(n4724), .B(n4514), .Y(n4725));
  NAND3X1 g3643(.A(n4471), .B(n3858), .C(n1891), .Y(n4726));
  OAI21X1 g3644(.A0(n4726), .A1(n4725), .B0(n4476), .Y(n4727));
  NOR3X1  g3645(.A(n4727), .B(n4470), .C(n2028), .Y(n4728));
  NOR2X1  g3646(.A(P1_STATE_REG_SCAN_IN), .B(P1_B_REG_SCAN_IN), .Y(n4729));
  NAND2X1 g3647(.A(n4473), .B(n2034), .Y(n4730));
  AOI21X1 g3648(.A0(n4724), .A1(n4514), .B0(n4730), .Y(n4731));
  NAND3X1 g3649(.A(n1989), .B(n1982), .C(n1873), .Y(n4732));
  NAND3X1 g3650(.A(n4488), .B(n3119), .C(n3759), .Y(n4733));
  NOR3X1  g3651(.A(n4419), .B(n4488), .C(n3421), .Y(n4735));
  OAI21X1 g3652(.A0(n2003), .A1(n1820), .B0(n3363), .Y(n4736));
  OAI21X1 g3653(.A0(n2003), .A1(n1650), .B0(n3070), .Y(n4740));
  NAND2X1 g3654(.A(n3050), .B(n4740), .Y(n4742));
  NOR2X1  g3655(.A(n3038), .B(n4742), .Y(n4744));
  AOI21X1 g3656(.A0(n3049), .A1(n4740), .B0(n3118), .Y(n4748));
  OAI21X1 g3657(.A0(n3109), .A1(n3120), .B0(n4748), .Y(n4749));
  AOI22X1 g3658(.A0(n2933), .A1(n2941), .B0(n2925), .B1(n2891), .Y(n4750));
  NAND2X1 g3659(.A(n2862), .B(n4750), .Y(n4752));
  OAI22X1 g3660(.A0(n2976), .A1(n2983), .B0(n2941), .B1(n2933), .Y(n4755));
  AOI21X1 g3661(.A0(n4450), .A1(n2985), .B0(n4755), .Y(n4756));
  NAND4X1 g3662(.A(n4752), .B(n3050), .C(n4740), .D(n4756), .Y(n4757));
  INVX1   g3663(.A(n4750), .Y(n4758));
  OAI22X1 g3664(.A0(n2840), .A1(n2853), .B0(n2806), .B1(n2792), .Y(n4759));
  NOR2X1  g3665(.A(n4759), .B(n4758), .Y(n4760));
  NAND2X1 g3666(.A(n2785), .B(n2798), .Y(n4761));
  NOR2X1  g3667(.A(n2496), .B(n2457), .Y(n4763));
  AOI22X1 g3668(.A0(n2363), .A1(n2376), .B0(n2324), .B1(n2312), .Y(n4766));
  NAND2X1 g3669(.A(n2225), .B(n2219), .Y(n4768));
  NOR2X1  g3670(.A(n2165), .B(n2160), .Y(n4769));
  AOI21X1 g3671(.A0(n4769), .A1(n4768), .B0(n2270), .Y(n4770));
  NAND2X1 g3672(.A(n4770), .B(n4766), .Y(n4771));
  NAND3X1 g3673(.A(n4766), .B(n4594), .C(n2283), .Y(n4772));
  AOI21X1 g3674(.A0(n4772), .A1(n4771), .B0(n2289), .Y(n4773));
  NAND2X1 g3675(.A(n2447), .B(n2408), .Y(n4774));
  NAND3X1 g3676(.A(n2376), .B(n2361), .C(n2357), .Y(n4776));
  NAND2X1 g3677(.A(n2330), .B(n4776), .Y(n4778));
  NAND3X1 g3678(.A(n4778), .B(n2474), .C(n4774), .Y(n4779));
  OAI21X1 g3679(.A0(n4779), .A1(n4773), .B0(n4433), .Y(n4780));
  NAND2X1 g3680(.A(n2496), .B(n2457), .Y(n4781));
  AOI21X1 g3681(.A0(n4781), .A1(n4780), .B0(n4763), .Y(n4782));
  AOI22X1 g3682(.A0(n2219), .A1(n2225), .B0(n2165), .B1(n2160), .Y(n4784));
  NAND4X1 g3683(.A(n4778), .B(n2474), .C(n4774), .D(n4784), .Y(n4785));
  NAND2X1 g3684(.A(n4781), .B(n4772), .Y(n4786));
  NAND3X1 g3685(.A(n2114), .B(n2101), .C(n2096), .Y(n4787));
  NOR4X1  g3686(.A(n4786), .B(n4785), .C(n2556), .D(n4787), .Y(n4788));
  OAI21X1 g3687(.A0(n2084), .A1(n2093), .B0(n2058), .Y(n4790));
  NAND2X1 g3688(.A(n2084), .B(n2093), .Y(n4791));
  OAI21X1 g3689(.A0(n2185), .A1(n2182), .B0(n2137), .Y(n4792));
  NAND3X1 g3690(.A(n4792), .B(n4791), .C(n4790), .Y(n4793));
  NOR4X1  g3691(.A(n4786), .B(n4785), .C(n2556), .D(n4793), .Y(n4794));
  OAI22X1 g3692(.A0(n2649), .A1(n2671), .B0(n2642), .B1(n2634), .Y(n4795));
  OAI22X1 g3693(.A0(n2580), .A1(n2593), .B0(n2517), .B1(n2503), .Y(n4796));
  NOR4X1  g3694(.A(n4795), .B(n4794), .C(n4788), .D(n4796), .Y(n4797));
  OAI21X1 g3695(.A0(n2556), .A1(n4782), .B0(n4797), .Y(n4798));
  NAND2X1 g3696(.A(n2593), .B(n2580), .Y(n4799));
  NOR2X1  g3697(.A(n4799), .B(n4795), .Y(n4800));
  AOI22X1 g3698(.A0(n2709), .A1(n2714), .B0(n2671), .B1(n2649), .Y(n4803));
  OAI21X1 g3699(.A0(n2987), .A1(n2672), .B0(n4803), .Y(n4804));
  NOR2X1  g3700(.A(n4804), .B(n4800), .Y(n4805));
  AOI21X1 g3701(.A0(n4805), .A1(n4798), .B0(n2761), .Y(n4806));
  OAI21X1 g3702(.A0(n2799), .A1(n4806), .B0(n4761), .Y(n4808));
  NAND2X1 g3703(.A(n2806), .B(n2792), .Y(n4809));
  NAND2X1 g3704(.A(n4809), .B(n4808), .Y(n4810));
  AOI21X1 g3705(.A0(n4810), .A1(n4760), .B0(n4757), .Y(n4811));
  NOR4X1  g3706(.A(n4749), .B(n4744), .C(n3169), .D(n4811), .Y(n4812));
  OAI21X1 g3707(.A0(n2003), .A1(n1697), .B0(n3149), .Y(n4814));
  NAND2X1 g3708(.A(n3109), .B(n3120), .Y(n4815));
  OAI21X1 g3709(.A0(n4815), .A1(n3169), .B0(n4814), .Y(n4816));
  NOR3X1  g3710(.A(n4816), .B(n3247), .C(n4812), .Y(n4817));
  OAI22X1 g3711(.A0(n3235), .A1(n3273), .B0(n3215), .B1(n3191), .Y(n4818));
  AOI22X1 g3712(.A0(n3281), .A1(n3294), .B0(n3273), .B1(n3235), .Y(n4819));
  OAI21X1 g3713(.A0(n4818), .A1(n4817), .B0(n4819), .Y(n4820));
  NAND2X1 g3714(.A(n4820), .B(n3334), .Y(n4821));
  OAI21X1 g3715(.A0(n4821), .A1(n3329), .B0(n3322), .Y(n4822));
  AOI21X1 g3716(.A0(n4821), .A1(n3329), .B0(n4408), .Y(n4824));
  NAND2X1 g3717(.A(n4824), .B(n4822), .Y(n4825));
  AOI21X1 g3718(.A0(n4825), .A1(n4736), .B0(n4419), .Y(n4826));
  OAI21X1 g3719(.A0(n4826), .A1(n4735), .B0(n4733), .Y(n4827));
  NAND3X1 g3720(.A(n3378), .B(n1991), .C(n1873), .Y(n4828));
  AOI21X1 g3721(.A0(n4391), .A1(n3769), .B0(n4828), .Y(n4829));
  XOR2X1  g3722(.A(n3423), .B(n3383), .Y(n4830));
  XOR2X1  g3723(.A(n3769), .B(n4390), .Y(n4831));
  XOR2X1  g3724(.A(n3294), .B(n3281), .Y(n4834));
  XOR2X1  g3725(.A(n3273), .B(n3236), .Y(n4835));
  XOR2X1  g3726(.A(n2853), .B(n2841), .Y(n4839));
  XOR2X1  g3727(.A(n2516), .B(n2503), .Y(n4840));
  XOR2X1  g3728(.A(n2026), .B(n2010), .Y(n4841));
  NOR4X1  g3729(.A(n2170), .B(n2115), .C(n2076), .D(n4841), .Y(n4842));
  NAND3X1 g3730(.A(n4842), .B(n2325), .C(n2226), .Y(n4843));
  XOR2X1  g3731(.A(n2268), .B(n4594), .Y(n4844));
  XOR2X1  g3732(.A(n2376), .B(n2362), .Y(n4845));
  NOR4X1  g3733(.A(n4844), .B(n4843), .C(n4840), .D(n4845), .Y(n4846));
  NOR3X1  g3734(.A(n2574), .B(n2486), .C(n2427), .Y(n4847));
  XOR2X1  g3735(.A(n2759), .B(n2798), .Y(n4848));
  XOR2X1  g3736(.A(n2665), .B(n2649), .Y(n4849));
  XOR2X1  g3737(.A(n2714), .B(n2702), .Y(n4850));
  NOR4X1  g3738(.A(n4849), .B(n4848), .C(n2635), .D(n4850), .Y(n4851));
  NAND4X1 g3739(.A(n4847), .B(n4846), .C(n2807), .D(n4851), .Y(n4852));
  NOR3X1  g3740(.A(n4852), .B(n4839), .C(n2910), .Y(n4853));
  NAND3X1 g3741(.A(n4853), .B(n2984), .C(n2942), .Y(n4854));
  AOI21X1 g3742(.A0(n3091), .A1(n3086), .B0(n4854), .Y(n4855));
  NAND3X1 g3743(.A(n4855), .B(n3079), .C(n3121), .Y(n4856));
  NOR4X1  g3744(.A(n4835), .B(n3216), .C(n3176), .D(n4856), .Y(n4857));
  NAND3X1 g3745(.A(n4857), .B(n4834), .C(n3330), .Y(n4858));
  NOR3X1  g3746(.A(n4858), .B(n3402), .C(n4831), .Y(n4859));
  NAND3X1 g3747(.A(n4859), .B(n4830), .C(n4462), .Y(n4860));
  AOI22X1 g3748(.A0(n4830), .A1(n4859), .B0(n2037), .B1(n1873), .Y(n4861));
  NOR2X1  g3749(.A(n4861), .B(n1989), .Y(n4862));
  AOI22X1 g3750(.A0(n4860), .A1(n4862), .B0(n4829), .B1(n4827), .Y(n4863));
  OAI21X1 g3751(.A0(n4732), .A1(n4725), .B0(n4863), .Y(n4864));
  NOR4X1  g3752(.A(n4731), .B(n4727), .C(n4470), .D(n4864), .Y(n4865));
  NOR3X1  g3753(.A(n4865), .B(n4729), .C(n4728), .Y(P1_U3242));
  AOI22X1 g3754(.A0(n4241), .A1(n2709), .B0(n2741), .B1(n4248), .Y(n4867));
  OAI22X1 g3755(.A0(n4242), .A1(n2702), .B0(n2714), .B1(n4247), .Y(n4868));
  XOR2X1  g3756(.A(n4868), .B(n4239), .Y(n4869));
  NOR2X1  g3757(.A(n4869), .B(n4867), .Y(n4870));
  NAND2X1 g3758(.A(n4869), .B(n4867), .Y(n4871));
  INVX1   g3759(.A(n2061), .Y(n4872));
  NOR2X1  g3760(.A(n2059), .B(n2034), .Y(n4873));
  AOI21X1 g3761(.A0(n4873), .A1(n2044), .B0(n1882), .Y(n4874));
  NOR2X1  g3762(.A(n4237), .B(n1882), .Y(n4875));
  NOR2X1  g3763(.A(n4875), .B(n4874), .Y(n4876));
  OAI21X1 g3764(.A0(n4872), .A1(n1882), .B0(n4876), .Y(n4877));
  AOI22X1 g3765(.A0(n4248), .A1(n2649), .B0(n2665), .B1(n4877), .Y(n4878));
  XOR2X1  g3766(.A(n4878), .B(n4246), .Y(n4879));
  AOI22X1 g3767(.A0(n4241), .A1(n2649), .B0(n2665), .B1(n4248), .Y(n4880));
  NAND2X1 g3768(.A(n4880), .B(n4879), .Y(n4881));
  INVX1   g3769(.A(n4881), .Y(n4882));
  AOI22X1 g3770(.A0(n4241), .A1(n2580), .B0(n2562), .B1(n4248), .Y(n4883));
  AOI22X1 g3771(.A0(n4248), .A1(n2580), .B0(n2562), .B1(n4877), .Y(n4884));
  XOR2X1  g3772(.A(n4884), .B(n4246), .Y(n4885));
  NOR2X1  g3773(.A(n4885), .B(n4883), .Y(n4886));
  AOI22X1 g3774(.A0(n4241), .A1(n2634), .B0(n2614), .B1(n4248), .Y(n4887));
  AOI22X1 g3775(.A0(n4248), .A1(n2634), .B0(n2614), .B1(n4877), .Y(n4888));
  XOR2X1  g3776(.A(n4888), .B(n4246), .Y(n4889));
  AOI22X1 g3777(.A0(n4887), .A1(n4889), .B0(n4880), .B1(n4879), .Y(n4890));
  OAI22X1 g3778(.A0(n4887), .A1(n4889), .B0(n4880), .B1(n4879), .Y(n4891));
  AOI21X1 g3779(.A0(n4890), .A1(n4886), .B0(n4891), .Y(n4892));
  AOI22X1 g3780(.A0(n4241), .A1(n2503), .B0(n2516), .B1(n4248), .Y(n4893));
  AOI22X1 g3781(.A0(n4248), .A1(n2503), .B0(n2516), .B1(n4877), .Y(n4894));
  XOR2X1  g3782(.A(n4894), .B(n4246), .Y(n4895));
  NOR2X1  g3783(.A(n4895), .B(n4893), .Y(n4896));
  NAND2X1 g3784(.A(n4895), .B(n4893), .Y(n4897));
  AOI22X1 g3785(.A0(n4248), .A1(n2457), .B0(n2469), .B1(n4877), .Y(n4898));
  XOR2X1  g3786(.A(n4898), .B(n4246), .Y(n4899));
  INVX1   g3787(.A(n4899), .Y(n4900));
  AOI22X1 g3788(.A0(n4241), .A1(n2457), .B0(n2469), .B1(n4248), .Y(n4901));
  INVX1   g3789(.A(n4901), .Y(n4902));
  NOR2X1  g3790(.A(n4902), .B(n4900), .Y(n4903));
  AOI22X1 g3791(.A0(n4241), .A1(n2408), .B0(n2424), .B1(n4248), .Y(n4904));
  AOI22X1 g3792(.A0(n4248), .A1(n2408), .B0(n2424), .B1(n4877), .Y(n4905));
  XOR2X1  g3793(.A(n4905), .B(n4246), .Y(n4906));
  NOR2X1  g3794(.A(n4906), .B(n4904), .Y(n4907));
  NAND2X1 g3795(.A(n4906), .B(n4904), .Y(n4908));
  AOI22X1 g3796(.A0(n4241), .A1(n2313), .B0(n2324), .B1(n4248), .Y(n4909));
  AOI22X1 g3797(.A0(n4248), .A1(n2313), .B0(n2324), .B1(n4877), .Y(n4910));
  XOR2X1  g3798(.A(n4910), .B(n4246), .Y(n4911));
  AOI22X1 g3799(.A0(n4241), .A1(n2362), .B0(n2376), .B1(n4248), .Y(n4912));
  AOI22X1 g3800(.A0(n4248), .A1(n2362), .B0(n2376), .B1(n4877), .Y(n4913));
  XOR2X1  g3801(.A(n4913), .B(n4246), .Y(n4914));
  AOI22X1 g3802(.A0(n4912), .A1(n4914), .B0(n4911), .B1(n4909), .Y(n4915));
  INVX1   g3803(.A(n4915), .Y(n4916));
  AOI22X1 g3804(.A0(n4241), .A1(n4594), .B0(n2268), .B1(n4248), .Y(n4917));
  AOI22X1 g3805(.A0(n4248), .A1(n4594), .B0(n2268), .B1(n4877), .Y(n4918));
  XOR2X1  g3806(.A(n4918), .B(n4246), .Y(n4919));
  NOR2X1  g3807(.A(n4919), .B(n4917), .Y(n4920));
  NAND2X1 g3808(.A(n4919), .B(n4917), .Y(n4921));
  AOI22X1 g3809(.A0(n4248), .A1(n2219), .B0(n2224), .B1(n4877), .Y(n4922));
  XOR2X1  g3810(.A(n4922), .B(n4246), .Y(n4923));
  AOI22X1 g3811(.A0(n4241), .A1(n2219), .B0(n2224), .B1(n4248), .Y(n4924));
  NAND2X1 g3812(.A(n4924), .B(n4923), .Y(n4925));
  INVX1   g3813(.A(n4925), .Y(n4926));
  AOI22X1 g3814(.A0(n4241), .A1(n2102), .B0(n2114), .B1(n4248), .Y(n4927));
  AOI22X1 g3815(.A0(n4248), .A1(n2102), .B0(n2114), .B1(n4877), .Y(n4928));
  XOR2X1  g3816(.A(n4928), .B(n4246), .Y(n4929));
  AOI22X1 g3817(.A0(n4241), .A1(n2160), .B0(n2169), .B1(n4248), .Y(n4930));
  AOI22X1 g3818(.A0(n4248), .A1(n2160), .B0(n2169), .B1(n4877), .Y(n4931));
  XOR2X1  g3819(.A(n4931), .B(n4246), .Y(n4932));
  AOI22X1 g3820(.A0(n4930), .A1(n4932), .B0(n4929), .B1(n4927), .Y(n4933));
  AOI22X1 g3821(.A0(n4241), .A1(n2058), .B0(n2075), .B1(n4248), .Y(n4934));
  INVX1   g3822(.A(n4934), .Y(n4935));
  AOI22X1 g3823(.A0(n4248), .A1(n2058), .B0(n2075), .B1(n4877), .Y(n4936));
  XOR2X1  g3824(.A(n4936), .B(n4239), .Y(n4937));
  NAND2X1 g3825(.A(n4937), .B(n4935), .Y(n4938));
  NOR2X1  g3826(.A(n4937), .B(n4935), .Y(n4939));
  NOR2X1  g3827(.A(n4244), .B(n4239), .Y(n4940));
  NAND2X1 g3828(.A(n4244), .B(n4239), .Y(n4941));
  AOI21X1 g3829(.A0(n4941), .A1(n4251), .B0(n4940), .Y(n4942));
  OAI21X1 g3830(.A0(n4942), .A1(n4939), .B0(n4938), .Y(n4943));
  INVX1   g3831(.A(n4927), .Y(n4944));
  XOR2X1  g3832(.A(n4928), .B(n4239), .Y(n4945));
  INVX1   g3833(.A(n4930), .Y(n4946));
  NAND3X1 g3834(.A(n4946), .B(n4945), .C(n4944), .Y(n4947));
  AOI21X1 g3835(.A0(n4945), .A1(n4944), .B0(n4946), .Y(n4948));
  OAI21X1 g3836(.A0(n4948), .A1(n4932), .B0(n4947), .Y(n4949));
  AOI21X1 g3837(.A0(n4943), .A1(n4933), .B0(n4949), .Y(n4950));
  NOR2X1  g3838(.A(n4924), .B(n4923), .Y(n4951));
  INVX1   g3839(.A(n4951), .Y(n4952));
  OAI21X1 g3840(.A0(n4950), .A1(n4926), .B0(n4952), .Y(n4953));
  AOI21X1 g3841(.A0(n4953), .A1(n4921), .B0(n4920), .Y(n4954));
  NOR2X1  g3842(.A(n4911), .B(n4909), .Y(n4955));
  INVX1   g3843(.A(n4955), .Y(n4956));
  INVX1   g3844(.A(n4912), .Y(n4957));
  INVX1   g3845(.A(n4914), .Y(n4958));
  OAI21X1 g3846(.A0(n4955), .A1(n4957), .B0(n4958), .Y(n4959));
  OAI21X1 g3847(.A0(n4956), .A1(n4912), .B0(n4959), .Y(n4960));
  INVX1   g3848(.A(n4960), .Y(n4961));
  OAI21X1 g3849(.A0(n4954), .A1(n4916), .B0(n4961), .Y(n4962));
  AOI21X1 g3850(.A0(n4962), .A1(n4908), .B0(n4907), .Y(n4963));
  NOR2X1  g3851(.A(n4901), .B(n4899), .Y(n4964));
  INVX1   g3852(.A(n4964), .Y(n4965));
  OAI21X1 g3853(.A0(n4963), .A1(n4903), .B0(n4965), .Y(n4966));
  AOI21X1 g3854(.A0(n4966), .A1(n4897), .B0(n4896), .Y(n4967));
  NAND2X1 g3855(.A(n4889), .B(n4887), .Y(n4968));
  INVX1   g3856(.A(n4968), .Y(n4969));
  NAND2X1 g3857(.A(n4885), .B(n4883), .Y(n4970));
  INVX1   g3858(.A(n4970), .Y(n4971));
  NOR3X1  g3859(.A(n4971), .B(n4969), .C(n4882), .Y(n4972));
  INVX1   g3860(.A(n4972), .Y(n4973));
  OAI22X1 g3861(.A0(n4967), .A1(n4973), .B0(n4892), .B1(n4882), .Y(n4974));
  AOI21X1 g3862(.A0(n4974), .A1(n4871), .B0(n4870), .Y(n4975));
  OAI22X1 g3863(.A0(n4242), .A1(n2798), .B0(n2759), .B1(n4247), .Y(n4976));
  XOR2X1  g3864(.A(n4976), .B(n4239), .Y(n4977));
  AOI22X1 g3865(.A0(n4241), .A1(n2749), .B0(n2785), .B1(n4248), .Y(n4978));
  XOR2X1  g3866(.A(n4978), .B(n4977), .Y(n4979));
  XOR2X1  g3867(.A(n4979), .B(n4975), .Y(n4980));
  NOR3X1  g3868(.A(n1997), .B(n1980), .C(n1978), .Y(n4981));
  OAI21X1 g3869(.A0(n2037), .A1(n2028), .B0(n1983), .Y(n4982));
  OAI21X1 g3870(.A0(n2037), .A1(n2028), .B0(n1989), .Y(n4983));
  NOR2X1  g3871(.A(n4983), .B(n1983), .Y(n4984));
  NOR4X1  g3872(.A(n3522), .B(n2045), .C(n2043), .D(n4984), .Y(n4985));
  OAI21X1 g3873(.A0(n4982), .A1(n1989), .B0(n4985), .Y(n4986));
  NAND3X1 g3874(.A(n4986), .B(n4981), .C(n1891), .Y(n4987));
  INVX1   g3875(.A(n4981), .Y(n4988));
  NOR4X1  g3876(.A(n1882), .B(n1873), .C(P1_U3086), .D(n3518), .Y(n4989));
  NAND3X1 g3877(.A(n3510), .B(n3946), .C(n1872), .Y(n4990));
  AOI21X1 g3878(.A0(n4986), .A1(n4988), .B0(n4990), .Y(n4991));
  NOR2X1  g3879(.A(n4991), .B(P1_U3086), .Y(n4992));
  AOI21X1 g3880(.A0(n4989), .A1(n4988), .B0(n4992), .Y(n4993));
  NOR4X1  g3881(.A(n1987), .B(n1982), .C(n1892), .D(n1992), .Y(n4995));
  INVX1   g3882(.A(n4995), .Y(n4996));
  NOR4X1  g3883(.A(n1997), .B(n1980), .C(n1978), .D(n2080), .Y(n4997));
  NOR4X1  g3884(.A(n1997), .B(n1980), .C(n1978), .D(n3941), .Y(n4998));
  INVX1   g3885(.A(n4998), .Y(n4999));
  OAI22X1 g3886(.A0(n4981), .A1(n2744), .B0(n2791), .B1(n4999), .Y(n5000));
  AOI21X1 g3887(.A0(n4997), .A1(n2709), .B0(n5000), .Y(n5001));
  AOI22X1 g3888(.A0(n4981), .A1(n4989), .B0(n3505), .B1(n1891), .Y(n5002));
  AOI22X1 g3889(.A0(n2785), .A1(n5150), .B0(P1_U3086), .B1(P1_REG3_REG_15__SCAN_IN), .Y(n5004));
  OAI21X1 g3890(.A0(n5001), .A1(n4996), .B0(n5004), .Y(n5005));
  AOI21X1 g3891(.A0(n5157), .A1(n2745), .B0(n5005), .Y(n5006));
  OAI21X1 g3892(.A0(n4987), .A1(n4980), .B0(n5006), .Y(P1_U3241));
  AOI22X1 g3893(.A0(n4241), .A1(n3149), .B0(n3157), .B1(n4248), .Y(n5008));
  INVX1   g3894(.A(n5008), .Y(n5009));
  OAI22X1 g3895(.A0(n4242), .A1(n3150), .B0(n3175), .B1(n4247), .Y(n5010));
  XOR2X1  g3896(.A(n5010), .B(n4246), .Y(n5011));
  NOR2X1  g3897(.A(n5011), .B(n5009), .Y(n5012));
  AOI22X1 g3898(.A0(n4241), .A1(n3109), .B0(n3142), .B1(n4248), .Y(n5013));
  OAI22X1 g3899(.A0(n4242), .A1(n3110), .B0(n3120), .B1(n4247), .Y(n5014));
  XOR2X1  g3900(.A(n5014), .B(n4239), .Y(n5015));
  NOR2X1  g3901(.A(n5015), .B(n5013), .Y(n5016));
  NAND2X1 g3902(.A(n5015), .B(n5013), .Y(n5017));
  AOI22X1 g3903(.A0(n4241), .A1(n3070), .B0(n3078), .B1(n4248), .Y(n5018));
  AOI22X1 g3904(.A0(n4248), .A1(n3070), .B0(n3078), .B1(n4877), .Y(n5019));
  XOR2X1  g3905(.A(n5019), .B(n4246), .Y(n5020));
  NOR2X1  g3906(.A(n5020), .B(n5018), .Y(n5021));
  INVX1   g3907(.A(n5021), .Y(n5022));
  NAND2X1 g3908(.A(n5020), .B(n5018), .Y(n5023));
  INVX1   g3909(.A(n5023), .Y(n5024));
  AOI22X1 g3910(.A0(n4248), .A1(n3028), .B0(n3036), .B1(n4877), .Y(n5025));
  XOR2X1  g3911(.A(n5025), .B(n4246), .Y(n5026));
  AOI22X1 g3912(.A0(n4241), .A1(n3028), .B0(n3036), .B1(n4248), .Y(n5027));
  NAND2X1 g3913(.A(n5027), .B(n5026), .Y(n5028));
  AOI22X1 g3914(.A0(n4241), .A1(n3002), .B0(n2941), .B1(n4248), .Y(n5029));
  AOI22X1 g3915(.A0(n4248), .A1(n3002), .B0(n2941), .B1(n4877), .Y(n5030));
  XOR2X1  g3916(.A(n5030), .B(n4246), .Y(n5031));
  NOR2X1  g3917(.A(n5031), .B(n5029), .Y(n5032));
  INVX1   g3918(.A(n5032), .Y(n5033));
  AOI22X1 g3919(.A0(n4241), .A1(n3001), .B0(n2983), .B1(n4248), .Y(n5034));
  AOI22X1 g3920(.A0(n4248), .A1(n3001), .B0(n2983), .B1(n4877), .Y(n5035));
  XOR2X1  g3921(.A(n5035), .B(n4246), .Y(n5036));
  NAND2X1 g3922(.A(n5036), .B(n5034), .Y(n5037));
  NAND2X1 g3923(.A(n5037), .B(n5028), .Y(n5038));
  INVX1   g3924(.A(n5026), .Y(n5039));
  INVX1   g3925(.A(n5027), .Y(n5040));
  NOR2X1  g3926(.A(n5036), .B(n5034), .Y(n5041));
  AOI21X1 g3927(.A0(n5040), .A1(n5039), .B0(n5041), .Y(n5042));
  OAI21X1 g3928(.A0(n5038), .A1(n5033), .B0(n5042), .Y(n5043));
  AOI22X1 g3929(.A0(n4241), .A1(n2902), .B0(n2925), .B1(n4248), .Y(n5044));
  OAI22X1 g3930(.A0(n4242), .A1(n2891), .B0(n2907), .B1(n4247), .Y(n5045));
  XOR2X1  g3931(.A(n5045), .B(n4239), .Y(n5046));
  NOR2X1  g3932(.A(n5046), .B(n5044), .Y(n5047));
  INVX1   g3933(.A(n5047), .Y(n5048));
  NAND2X1 g3934(.A(n5046), .B(n5044), .Y(n5049));
  INVX1   g3935(.A(n5049), .Y(n5050));
  AOI22X1 g3936(.A0(n4241), .A1(n2792), .B0(n2811), .B1(n4248), .Y(n5051));
  OAI22X1 g3937(.A0(n4242), .A1(n2791), .B0(n2806), .B1(n4247), .Y(n5052));
  XOR2X1  g3938(.A(n5052), .B(n4239), .Y(n5053));
  AOI22X1 g3939(.A0(n4241), .A1(n2840), .B0(n2854), .B1(n4248), .Y(n5054));
  AOI22X1 g3940(.A0(n4248), .A1(n2840), .B0(n2854), .B1(n4877), .Y(n5055));
  XOR2X1  g3941(.A(n5055), .B(n4246), .Y(n5056));
  AOI22X1 g3942(.A0(n5054), .A1(n5056), .B0(n5053), .B1(n5051), .Y(n5057));
  NOR2X1  g3943(.A(n4978), .B(n4977), .Y(n5058));
  INVX1   g3944(.A(n5058), .Y(n5059));
  NAND2X1 g3945(.A(n4978), .B(n4977), .Y(n5060));
  INVX1   g3946(.A(n5060), .Y(n5061));
  OAI21X1 g3947(.A0(n5061), .A1(n4975), .B0(n5059), .Y(n5062));
  NOR3X1  g3948(.A(n5054), .B(n5053), .C(n5051), .Y(n5063));
  NOR2X1  g3949(.A(n5053), .B(n5051), .Y(n5064));
  INVX1   g3950(.A(n5064), .Y(n5065));
  AOI21X1 g3951(.A0(n5065), .A1(n5054), .B0(n5056), .Y(n5066));
  NOR2X1  g3952(.A(n5066), .B(n5063), .Y(n5067));
  INVX1   g3953(.A(n5067), .Y(n5068));
  AOI21X1 g3954(.A0(n5062), .A1(n5057), .B0(n5068), .Y(n5069));
  OAI21X1 g3955(.A0(n5069), .A1(n5050), .B0(n5048), .Y(n5070));
  NAND2X1 g3956(.A(n5031), .B(n5029), .Y(n5071));
  INVX1   g3957(.A(n5071), .Y(n5072));
  NOR2X1  g3958(.A(n5072), .B(n5038), .Y(n5073));
  AOI22X1 g3959(.A0(n5070), .A1(n5073), .B0(n5043), .B1(n5028), .Y(n5074));
  OAI21X1 g3960(.A0(n5074), .A1(n5024), .B0(n5022), .Y(n5075));
  AOI21X1 g3961(.A0(n5075), .A1(n5017), .B0(n5016), .Y(n5076));
  AOI22X1 g3962(.A0(n4241), .A1(n3191), .B0(n3199), .B1(n4248), .Y(n5077));
  INVX1   g3963(.A(n5077), .Y(n5078));
  OAI22X1 g3964(.A0(n4242), .A1(n3192), .B0(n3215), .B1(n4247), .Y(n5079));
  XOR2X1  g3965(.A(n5079), .B(n4239), .Y(n5080));
  INVX1   g3966(.A(n5080), .Y(n5081));
  NAND2X1 g3967(.A(n5011), .B(n5009), .Y(n5082));
  INVX1   g3968(.A(n5082), .Y(n5083));
  AOI21X1 g3969(.A0(n5081), .A1(n5078), .B0(n5083), .Y(n5084));
  OAI21X1 g3970(.A0(n5076), .A1(n5012), .B0(n5084), .Y(n5085));
  OAI22X1 g3971(.A0(n4242), .A1(n3236), .B0(n3273), .B1(n4247), .Y(n5086));
  XOR2X1  g3972(.A(n5086), .B(n4239), .Y(n5087));
  OAI22X1 g3973(.A0(n4876), .A1(n3236), .B0(n3273), .B1(n4242), .Y(n5088));
  INVX1   g3974(.A(n5088), .Y(n5089));
  NOR2X1  g3975(.A(n5089), .B(n5087), .Y(n5090));
  INVX1   g3976(.A(n5090), .Y(n5091));
  AOI22X1 g3977(.A0(n5087), .A1(n5089), .B0(n5080), .B1(n5077), .Y(n5092));
  NAND3X1 g3978(.A(n5092), .B(n5091), .C(n5085), .Y(n5093));
  INVX1   g3979(.A(n5012), .Y(n5094));
  INVX1   g3980(.A(n5016), .Y(n5095));
  INVX1   g3981(.A(n5017), .Y(n5096));
  NAND2X1 g3982(.A(n5043), .B(n5028), .Y(n5097));
  INVX1   g3983(.A(n5057), .Y(n5098));
  INVX1   g3984(.A(n4870), .Y(n5099));
  INVX1   g3985(.A(n4871), .Y(n5100));
  NOR2X1  g3986(.A(n4892), .B(n4882), .Y(n5101));
  INVX1   g3987(.A(n4896), .Y(n5102));
  INVX1   g3988(.A(n4897), .Y(n5103));
  INVX1   g3989(.A(n4903), .Y(n5104));
  INVX1   g3990(.A(n4907), .Y(n5105));
  INVX1   g3991(.A(n4908), .Y(n5106));
  INVX1   g3992(.A(n4920), .Y(n5107));
  INVX1   g3993(.A(n4921), .Y(n5108));
  XOR2X1  g3994(.A(n4931), .B(n4239), .Y(n5109));
  OAI22X1 g3995(.A0(n4946), .A1(n5109), .B0(n4945), .B1(n4944), .Y(n5110));
  XOR2X1  g3996(.A(n4936), .B(n4246), .Y(n5111));
  NOR2X1  g3997(.A(n5111), .B(n4934), .Y(n5112));
  NAND2X1 g3998(.A(n5111), .B(n4934), .Y(n5113));
  XOR2X1  g3999(.A(n4250), .B(n4239), .Y(n5114));
  AOI22X1 g4000(.A0(n2010), .A1(n4248), .B0(n2008), .B1(n1882), .Y(n5115));
  OAI21X1 g4001(.A0(n4876), .A1(n2128), .B0(n5115), .Y(n5116));
  NAND2X1 g4002(.A(n5116), .B(n4246), .Y(n5117));
  NOR2X1  g4003(.A(n5116), .B(n4246), .Y(n5118));
  OAI21X1 g4004(.A0(n5118), .A1(n5114), .B0(n5117), .Y(n5119));
  AOI21X1 g4005(.A0(n5119), .A1(n5113), .B0(n5112), .Y(n5120));
  NOR3X1  g4006(.A(n4930), .B(n4929), .C(n4927), .Y(n5121));
  OAI21X1 g4007(.A0(n4929), .A1(n4927), .B0(n4930), .Y(n5122));
  AOI21X1 g4008(.A0(n5122), .A1(n5109), .B0(n5121), .Y(n5123));
  OAI21X1 g4009(.A0(n5120), .A1(n5110), .B0(n5123), .Y(n5124));
  AOI21X1 g4010(.A0(n5124), .A1(n4925), .B0(n4951), .Y(n5125));
  OAI21X1 g4011(.A0(n5125), .A1(n5108), .B0(n5107), .Y(n5126));
  AOI21X1 g4012(.A0(n5126), .A1(n4915), .B0(n4960), .Y(n5127));
  OAI21X1 g4013(.A0(n5127), .A1(n5106), .B0(n5105), .Y(n5128));
  AOI21X1 g4014(.A0(n5128), .A1(n5104), .B0(n4964), .Y(n5129));
  OAI21X1 g4015(.A0(n5129), .A1(n5103), .B0(n5102), .Y(n5130));
  AOI21X1 g4016(.A0(n4972), .A1(n5130), .B0(n5101), .Y(n5131));
  OAI21X1 g4017(.A0(n5131), .A1(n5100), .B0(n5099), .Y(n5132));
  AOI21X1 g4018(.A0(n5060), .A1(n5132), .B0(n5058), .Y(n5133));
  OAI21X1 g4019(.A0(n5133), .A1(n5098), .B0(n5067), .Y(n5134));
  AOI21X1 g4020(.A0(n5134), .A1(n5049), .B0(n5047), .Y(n5135));
  INVX1   g4021(.A(n5073), .Y(n5136));
  OAI21X1 g4022(.A0(n5136), .A1(n5135), .B0(n5097), .Y(n5137));
  AOI21X1 g4023(.A0(n5137), .A1(n5023), .B0(n5021), .Y(n5138));
  OAI21X1 g4024(.A0(n5138), .A1(n5096), .B0(n5095), .Y(n5139));
  AOI21X1 g4025(.A0(n5139), .A1(n5094), .B0(n5083), .Y(n5140));
  XOR2X1  g4026(.A(n5089), .B(n5087), .Y(n5141));
  AOI21X1 g4027(.A0(n5081), .A1(n5078), .B0(n5141), .Y(n5142));
  INVX1   g4028(.A(n4987), .Y(n5143));
  NAND2X1 g4029(.A(n5080), .B(n5077), .Y(n5144));
  OAI21X1 g4030(.A0(n5141), .A1(n5144), .B0(n5143), .Y(n5145));
  AOI21X1 g4031(.A0(n5142), .A1(n5140), .B0(n5145), .Y(n5146));
  NAND2X1 g4032(.A(n5146), .B(n5093), .Y(n5147));
  INVX1   g4033(.A(n3518), .Y(n5148));
  NAND4X1 g4034(.A(n3439), .B(n3507), .C(n1977), .D(n5148), .Y(n5149));
  AOI21X1 g4035(.A0(n5149), .A1(n3506), .B0(n1892), .Y(n5150));
  NAND2X1 g4036(.A(n5150), .B(n3243), .Y(n5151));
  NOR2X1  g4037(.A(n4999), .B(n3282), .Y(n5152));
  INVX1   g4038(.A(n4997), .Y(n5153));
  OAI22X1 g4039(.A0(n4981), .A1(n3231), .B0(n3192), .B1(n5153), .Y(n5154));
  OAI21X1 g4040(.A0(n5154), .A1(n5152), .B0(n4995), .Y(n5155));
  NAND2X1 g4041(.A(n4988), .B(n5148), .Y(n5156));
  AOI21X1 g4042(.A0(n5156), .A1(n4991), .B0(P1_U3086), .Y(n5157));
  AOI22X1 g4043(.A0(n3722), .A1(n5157), .B0(P1_U3086), .B1(P1_REG3_REG_26__SCAN_IN), .Y(n5158));
  NAND4X1 g4044(.A(n5155), .B(n5151), .C(n5147), .D(n5158), .Y(P1_U3240));
  INVX1   g4045(.A(n4909), .Y(n5160));
  XOR2X1  g4046(.A(n4911), .B(n5160), .Y(n5161));
  NOR2X1  g4047(.A(n5161), .B(n5126), .Y(n5162));
  XOR2X1  g4048(.A(n4911), .B(n4909), .Y(n5163));
  NOR2X1  g4049(.A(n5163), .B(n4954), .Y(n5164));
  OAI21X1 g4050(.A0(n5164), .A1(n5162), .B0(n5143), .Y(n5165));
  OAI22X1 g4051(.A0(n4981), .A1(n2308), .B0(n2257), .B1(n5153), .Y(n5166));
  AOI21X1 g4052(.A0(n4998), .A1(n2362), .B0(n5166), .Y(n5167));
  AOI22X1 g4053(.A0(n2324), .A1(n5150), .B0(P1_U3086), .B1(P1_REG3_REG_6__SCAN_IN), .Y(n5168));
  OAI21X1 g4054(.A0(n5167), .A1(n4996), .B0(n5168), .Y(n5169));
  AOI21X1 g4055(.A0(n5157), .A1(n2309), .B0(n5169), .Y(n5170));
  NAND2X1 g4056(.A(n5170), .B(n5165), .Y(P1_U3239));
  XOR2X1  g4057(.A(n5046), .B(n5044), .Y(n5172));
  XOR2X1  g4058(.A(n5172), .B(n5069), .Y(n5173));
  AOI22X1 g4059(.A0(n4988), .A1(n2887), .B0(n3002), .B1(n4998), .Y(n5174));
  OAI21X1 g4060(.A0(n5153), .A1(n2841), .B0(n5174), .Y(n5175));
  AOI22X1 g4061(.A0(n4995), .A1(n5175), .B0(P1_U3086), .B1(P1_REG3_REG_18__SCAN_IN), .Y(n5176));
  OAI21X1 g4062(.A0(n4993), .A1(n2886), .B0(n5176), .Y(n5177));
  AOI21X1 g4063(.A0(n5150), .A1(n2925), .B0(n5177), .Y(n5178));
  OAI21X1 g4064(.A0(n5173), .A1(n4987), .B0(n5178), .Y(P1_U3238));
  XOR2X1  g4065(.A(n4945), .B(n4927), .Y(n5180));
  NOR2X1  g4066(.A(n4945), .B(n4944), .Y(n5181));
  NOR2X1  g4067(.A(n4929), .B(n4927), .Y(n5182));
  OAI21X1 g4068(.A0(n5182), .A1(n5181), .B0(n4943), .Y(n5183));
  OAI21X1 g4069(.A0(n5180), .A1(n4943), .B0(n5183), .Y(n5184));
  NAND2X1 g4070(.A(n5184), .B(n5143), .Y(n5185));
  NAND2X1 g4071(.A(n4998), .B(n2160), .Y(n5186));
  AOI22X1 g4072(.A0(n4988), .A1(P1_REG3_REG_2__SCAN_IN), .B0(n2058), .B1(n4997), .Y(n5187));
  AOI21X1 g4073(.A0(n5187), .A1(n5186), .B0(n4996), .Y(n5188));
  AOI22X1 g4074(.A0(n2114), .A1(n5150), .B0(P1_U3086), .B1(P1_REG3_REG_2__SCAN_IN), .Y(n5189));
  OAI21X1 g4075(.A0(n4993), .A1(n2184), .B0(n5189), .Y(n5190));
  NOR2X1  g4076(.A(n5190), .B(n5188), .Y(n5191));
  NAND2X1 g4077(.A(n5191), .B(n5185), .Y(P1_U3237));
  INVX1   g4078(.A(n4883), .Y(n5193));
  XOR2X1  g4079(.A(n4885), .B(n5193), .Y(n5194));
  OAI21X1 g4080(.A0(n4971), .A1(n4886), .B0(n5130), .Y(n5195));
  OAI21X1 g4081(.A0(n5194), .A1(n5130), .B0(n5195), .Y(n5196));
  NAND2X1 g4082(.A(n5196), .B(n5143), .Y(n5197));
  OAI22X1 g4083(.A0(n4981), .A1(n2543), .B0(n2504), .B1(n5153), .Y(n5198));
  AOI21X1 g4084(.A0(n4998), .A1(n2634), .B0(n5198), .Y(n5199));
  AOI22X1 g4085(.A0(n2562), .A1(n5150), .B0(P1_U3086), .B1(P1_REG3_REG_11__SCAN_IN), .Y(n5200));
  OAI21X1 g4086(.A0(n5199), .A1(n4996), .B0(n5200), .Y(n5201));
  AOI21X1 g4087(.A0(n5157), .A1(n3605), .B0(n5201), .Y(n5202));
  NAND2X1 g4088(.A(n5202), .B(n5197), .Y(P1_U3236));
  XOR2X1  g4089(.A(n5020), .B(n5018), .Y(n5204));
  XOR2X1  g4090(.A(n5204), .B(n5074), .Y(n5205));
  AOI22X1 g4091(.A0(n4988), .A1(n3065), .B0(n3028), .B1(n4997), .Y(n5207));
  OAI21X1 g4092(.A0(n4999), .A1(n3110), .B0(n5207), .Y(n5208));
  AOI22X1 g4093(.A0(n4995), .A1(n5208), .B0(P1_U3086), .B1(P1_REG3_REG_22__SCAN_IN), .Y(n5209));
  OAI21X1 g4094(.A0(n4993), .A1(n3066), .B0(n5209), .Y(n5210));
  AOI21X1 g4095(.A0(n5150), .A1(n3078), .B0(n5210), .Y(n5211));
  OAI21X1 g4096(.A0(n5205), .A1(n4987), .B0(n5211), .Y(P1_U3235));
  NOR2X1  g4097(.A(n4889), .B(n4887), .Y(n5213));
  INVX1   g4098(.A(n5213), .Y(n5214));
  AOI21X1 g4099(.A0(n4970), .A1(n5130), .B0(n4886), .Y(n5215));
  OAI21X1 g4100(.A0(n4880), .A1(n4879), .B0(n4890), .Y(n5216));
  AOI21X1 g4101(.A0(n5215), .A1(n5214), .B0(n5216), .Y(n5217));
  INVX1   g4102(.A(n4880), .Y(n5218));
  OAI22X1 g4103(.A0(n4887), .A1(n4889), .B0(n5218), .B1(n4879), .Y(n5219));
  AOI21X1 g4104(.A0(n5218), .A1(n4879), .B0(n5219), .Y(n5220));
  OAI21X1 g4105(.A0(n5215), .A1(n4969), .B0(n5220), .Y(n5221));
  NAND2X1 g4106(.A(n5221), .B(n5143), .Y(n5222));
  OAI22X1 g4107(.A0(n4981), .A1(n2645), .B0(n2702), .B1(n4999), .Y(n5223));
  AOI21X1 g4108(.A0(n4997), .A1(n2634), .B0(n5223), .Y(n5224));
  AOI22X1 g4109(.A0(n2665), .A1(n5150), .B0(P1_U3086), .B1(P1_REG3_REG_13__SCAN_IN), .Y(n5225));
  OAI21X1 g4110(.A0(n5224), .A1(n4996), .B0(n5225), .Y(n5226));
  AOI21X1 g4111(.A0(n5157), .A1(n2646), .B0(n5226), .Y(n5227));
  OAI21X1 g4112(.A0(n5222), .A1(n5217), .B0(n5227), .Y(P1_U3234));
  AOI21X1 g4113(.A0(n5071), .A1(n5070), .B0(n5032), .Y(n5229));
  XOR2X1  g4114(.A(n5036), .B(n5034), .Y(n5230));
  NAND2X1 g4115(.A(n5229), .B(n5230), .Y(n5231));
  OAI21X1 g4116(.A0(n5230), .A1(n5229), .B0(n5231), .Y(n5233));
  NAND2X1 g4117(.A(n5233), .B(n5143), .Y(n5234));
  NAND2X1 g4118(.A(n5150), .B(n2983), .Y(n5235));
  OAI22X1 g4119(.A0(n4981), .A1(n2971), .B0(n3029), .B1(n4999), .Y(n5236));
  AOI21X1 g4120(.A0(n4997), .A1(n3002), .B0(n5236), .Y(n5237));
  OAI22X1 g4121(.A0(n4996), .A1(n5237), .B0(P1_STATE_REG_SCAN_IN), .B1(n2968), .Y(n5238));
  AOI21X1 g4122(.A0(n5157), .A1(n2972), .B0(n5238), .Y(n5239));
  NAND3X1 g4123(.A(n5239), .B(n5235), .C(n5234), .Y(P1_U3233));
  OAI21X1 g4124(.A0(n4995), .A1(n4989), .B0(n4988), .Y(n5241));
  OAI21X1 g4125(.A0(n4991), .A1(P1_U3086), .B0(n5241), .Y(n5242));
  NAND2X1 g4126(.A(n5242), .B(P1_REG3_REG_0__SCAN_IN), .Y(n5243));
  NOR2X1  g4127(.A(n4996), .B(n2117), .Y(n5244));
  AOI22X1 g4128(.A0(n4998), .A1(n5244), .B0(P1_U3086), .B1(P1_REG3_REG_0__SCAN_IN), .Y(n5245));
  OAI21X1 g4129(.A0(n5002), .A1(n2011), .B0(n5245), .Y(n5246));
  AOI21X1 g4130(.A0(n5143), .A1(n4252), .B0(n5246), .Y(n5247));
  NAND2X1 g4131(.A(n5247), .B(n5243), .Y(P1_U3232));
  XOR2X1  g4132(.A(n4901), .B(n4899), .Y(n5249));
  XOR2X1  g4133(.A(n5249), .B(n4963), .Y(n5250));
  OAI22X1 g4134(.A0(n4981), .A1(n2451), .B0(n2409), .B1(n5153), .Y(n5251));
  AOI21X1 g4135(.A0(n4998), .A1(n2503), .B0(n5251), .Y(n5252));
  AOI22X1 g4136(.A0(n2469), .A1(n5150), .B0(P1_U3086), .B1(P1_REG3_REG_9__SCAN_IN), .Y(n5253));
  OAI21X1 g4137(.A0(n5252), .A1(n4996), .B0(n5253), .Y(n5254));
  AOI21X1 g4138(.A0(n5157), .A1(n3589), .B0(n5254), .Y(n5255));
  OAI21X1 g4139(.A0(n5250), .A1(n4987), .B0(n5255), .Y(P1_U3231));
  XOR2X1  g4140(.A(n4924), .B(n4923), .Y(n5257));
  XOR2X1  g4141(.A(n5257), .B(n4950), .Y(n5258));
  NOR2X1  g4142(.A(n4993), .B(n2202), .Y(n5259));
  OAI22X1 g4143(.A0(n4981), .A1(n2202), .B0(n2146), .B1(n5153), .Y(n5260));
  AOI21X1 g4144(.A0(n4998), .A1(n4594), .B0(n5260), .Y(n5261));
  AOI22X1 g4145(.A0(n2224), .A1(n5150), .B0(P1_U3086), .B1(P1_REG3_REG_4__SCAN_IN), .Y(n5262));
  OAI21X1 g4146(.A0(n5261), .A1(n4996), .B0(n5262), .Y(n5263));
  NOR2X1  g4147(.A(n5263), .B(n5259), .Y(n5264));
  OAI21X1 g4148(.A0(n5258), .A1(n4987), .B0(n5264), .Y(P1_U3230));
  XOR2X1  g4149(.A(n5011), .B(n5008), .Y(n5266));
  NOR2X1  g4150(.A(n5266), .B(n5139), .Y(n5267));
  AOI21X1 g4151(.A0(n5082), .A1(n5094), .B0(n5076), .Y(n5268));
  OAI21X1 g4152(.A0(n5268), .A1(n5267), .B0(n5143), .Y(n5269));
  NAND2X1 g4153(.A(n5150), .B(n3157), .Y(n5270));
  NOR2X1  g4154(.A(n4999), .B(n3192), .Y(n5271));
  OAI22X1 g4155(.A0(n4981), .A1(n3145), .B0(n3110), .B1(n5153), .Y(n5272));
  OAI21X1 g4156(.A0(n5272), .A1(n5271), .B0(n4995), .Y(n5273));
  AOI22X1 g4157(.A0(n3704), .A1(n5157), .B0(P1_U3086), .B1(P1_REG3_REG_24__SCAN_IN), .Y(n5274));
  NAND4X1 g4158(.A(n5273), .B(n5270), .C(n5269), .D(n5274), .Y(P1_U3229));
  OAI21X1 g4159(.A0(n5056), .A1(n5054), .B0(n5057), .Y(n5276));
  AOI21X1 g4160(.A0(n5065), .A1(n5133), .B0(n5276), .Y(n5277));
  AOI21X1 g4161(.A0(n5053), .A1(n5051), .B0(n5133), .Y(n5278));
  INVX1   g4162(.A(n5056), .Y(n5279));
  AOI21X1 g4163(.A0(n5279), .A1(n5054), .B0(n5064), .Y(n5280));
  OAI21X1 g4164(.A0(n5279), .A1(n5054), .B0(n5280), .Y(n5281));
  OAI21X1 g4165(.A0(n5281), .A1(n5278), .B0(n5143), .Y(n5282));
  AOI22X1 g4166(.A0(n4988), .A1(n2836), .B0(n2902), .B1(n4998), .Y(n5283));
  OAI21X1 g4167(.A0(n5153), .A1(n2791), .B0(n5283), .Y(n5284));
  AOI22X1 g4168(.A0(n4995), .A1(n5284), .B0(P1_U3086), .B1(P1_REG3_REG_17__SCAN_IN), .Y(n5285));
  OAI21X1 g4169(.A0(n4993), .A1(n2835), .B0(n5285), .Y(n5286));
  AOI21X1 g4170(.A0(n5150), .A1(n2854), .B0(n5286), .Y(n5287));
  OAI21X1 g4171(.A0(n5282), .A1(n5277), .B0(n5287), .Y(P1_U3228));
  XOR2X1  g4172(.A(n4919), .B(n4917), .Y(n5289));
  XOR2X1  g4173(.A(n5289), .B(n5125), .Y(n5290));
  OAI22X1 g4174(.A0(n4981), .A1(n2253), .B0(n2204), .B1(n5153), .Y(n5291));
  AOI21X1 g4175(.A0(n4998), .A1(n2313), .B0(n5291), .Y(n5292));
  AOI22X1 g4176(.A0(n2268), .A1(n5150), .B0(P1_U3086), .B1(P1_REG3_REG_5__SCAN_IN), .Y(n5293));
  OAI21X1 g4177(.A0(n5292), .A1(n4996), .B0(n5293), .Y(n5294));
  AOI21X1 g4178(.A0(n5157), .A1(n2254), .B0(n5294), .Y(n5295));
  OAI21X1 g4179(.A0(n5290), .A1(n4987), .B0(n5295), .Y(P1_U3227));
  INVX1   g4180(.A(n5051), .Y(n5297));
  XOR2X1  g4181(.A(n5053), .B(n5297), .Y(n5298));
  NOR2X1  g4182(.A(n5298), .B(n5062), .Y(n5299));
  XOR2X1  g4183(.A(n5053), .B(n5051), .Y(n5300));
  NOR2X1  g4184(.A(n5300), .B(n5133), .Y(n5301));
  OAI21X1 g4185(.A0(n5301), .A1(n5299), .B0(n5143), .Y(n5302));
  NAND2X1 g4186(.A(n5157), .B(n2787), .Y(n5303));
  AOI22X1 g4187(.A0(n4988), .A1(n2787), .B0(n2840), .B1(n4998), .Y(n5304));
  OAI21X1 g4188(.A0(n5153), .A1(n2798), .B0(n5304), .Y(n5305));
  NAND2X1 g4189(.A(n5305), .B(n4995), .Y(n5306));
  AOI22X1 g4190(.A0(n2811), .A1(n5150), .B0(P1_U3086), .B1(P1_REG3_REG_16__SCAN_IN), .Y(n5307));
  NAND4X1 g4191(.A(n5306), .B(n5303), .C(n5302), .D(n5307), .Y(P1_U3226));
  OAI21X1 g4192(.A0(n5076), .A1(n5012), .B0(n5082), .Y(n5309));
  XOR2X1  g4193(.A(n5080), .B(n5078), .Y(n5310));
  NOR2X1  g4194(.A(n5310), .B(n5309), .Y(n5311));
  XOR2X1  g4195(.A(n5080), .B(n5077), .Y(n5312));
  NOR2X1  g4196(.A(n5312), .B(n5140), .Y(n5313));
  OAI21X1 g4197(.A0(n5313), .A1(n5311), .B0(n5143), .Y(n5314));
  NAND2X1 g4198(.A(n5150), .B(n3199), .Y(n5315));
  AOI22X1 g4199(.A0(n4988), .A1(n3713), .B0(n3149), .B1(n4997), .Y(n5316));
  OAI21X1 g4200(.A0(n4999), .A1(n3236), .B0(n5316), .Y(n5317));
  OAI22X1 g4201(.A0(n3187), .A1(n4993), .B0(P1_STATE_REG_SCAN_IN), .B1(n3229), .Y(n5318));
  AOI21X1 g4202(.A0(n5317), .A1(n4995), .B0(n5318), .Y(n5319));
  NAND3X1 g4203(.A(n5319), .B(n5315), .C(n5314), .Y(P1_U3225));
  NOR2X1  g4204(.A(n4971), .B(n4967), .Y(n5321));
  INVX1   g4205(.A(n4887), .Y(n5322));
  XOR2X1  g4206(.A(n4889), .B(n5322), .Y(n5323));
  NOR3X1  g4207(.A(n5323), .B(n5321), .C(n4886), .Y(n5324));
  AOI21X1 g4208(.A0(n5214), .A1(n4968), .B0(n5215), .Y(n5325));
  OAI21X1 g4209(.A0(n5325), .A1(n5324), .B0(n5143), .Y(n5326));
  OAI22X1 g4210(.A0(n4981), .A1(n2596), .B0(n2650), .B1(n4999), .Y(n5327));
  AOI21X1 g4211(.A0(n4997), .A1(n2580), .B0(n5327), .Y(n5328));
  AOI22X1 g4212(.A0(n2614), .A1(n5150), .B0(P1_U3086), .B1(P1_REG3_REG_12__SCAN_IN), .Y(n5329));
  OAI21X1 g4213(.A0(n5328), .A1(n4996), .B0(n5329), .Y(n5330));
  AOI21X1 g4214(.A0(n5157), .A1(n3614), .B0(n5330), .Y(n5331));
  NAND2X1 g4215(.A(n5331), .B(n5326), .Y(P1_U3224));
  INVX1   g4216(.A(n5229), .Y(n5333));
  AOI21X1 g4217(.A0(n5040), .A1(n5039), .B0(n5038), .Y(n5334));
  OAI21X1 g4218(.A0(n5333), .A1(n5041), .B0(n5334), .Y(n5335));
  AOI21X1 g4219(.A0(n5027), .A1(n5039), .B0(n5041), .Y(n5336));
  OAI21X1 g4220(.A0(n5027), .A1(n5039), .B0(n5336), .Y(n5337));
  AOI21X1 g4221(.A0(n5333), .A1(n5037), .B0(n5337), .Y(n5338));
  NOR2X1  g4222(.A(n5338), .B(n4987), .Y(n5339));
  NAND2X1 g4223(.A(n5339), .B(n5335), .Y(n5340));
  NAND2X1 g4224(.A(n5150), .B(n3036), .Y(n5341));
  OAI22X1 g4225(.A0(n4981), .A1(n3024), .B0(n3071), .B1(n4999), .Y(n5342));
  AOI21X1 g4226(.A0(n4997), .A1(n3001), .B0(n5342), .Y(n5343));
  OAI22X1 g4227(.A0(n4996), .A1(n5343), .B0(P1_STATE_REG_SCAN_IN), .B1(n3022), .Y(n5344));
  AOI21X1 g4228(.A0(n5157), .A1(n3678), .B0(n5344), .Y(n5345));
  NAND3X1 g4229(.A(n5345), .B(n5341), .C(n5340), .Y(P1_U3223));
  AOI22X1 g4230(.A0(n4988), .A1(P1_REG3_REG_1__SCAN_IN), .B0(n2026), .B1(n4997), .Y(n5347));
  OAI21X1 g4231(.A0(n4999), .A1(n2103), .B0(n5347), .Y(n5348));
  OAI22X1 g4232(.A0(n2093), .A1(n5002), .B0(P1_STATE_REG_SCAN_IN), .B1(n4309), .Y(n5349));
  AOI21X1 g4233(.A0(n5348), .A1(n4995), .B0(n5349), .Y(n5350));
  XOR2X1  g4234(.A(n5111), .B(n4934), .Y(n5351));
  XOR2X1  g4235(.A(n5351), .B(n5119), .Y(n5352));
  AOI22X1 g4236(.A0(n5157), .A1(P1_REG3_REG_1__SCAN_IN), .B0(n5143), .B1(n5352), .Y(n5353));
  NAND2X1 g4237(.A(n5353), .B(n5350), .Y(P1_U3222));
  XOR2X1  g4238(.A(n4906), .B(n4904), .Y(n5355));
  XOR2X1  g4239(.A(n5355), .B(n5127), .Y(n5356));
  OAI22X1 g4240(.A0(n4981), .A1(n2405), .B0(n2363), .B1(n5153), .Y(n5357));
  AOI21X1 g4241(.A0(n4998), .A1(n2457), .B0(n5357), .Y(n5358));
  AOI22X1 g4242(.A0(n2424), .A1(n5150), .B0(P1_U3086), .B1(P1_REG3_REG_8__SCAN_IN), .Y(n5359));
  OAI21X1 g4243(.A0(n5358), .A1(n4996), .B0(n5359), .Y(n5360));
  AOI21X1 g4244(.A0(n5157), .A1(n2406), .B0(n5360), .Y(n5361));
  OAI21X1 g4245(.A0(n5356), .A1(n4987), .B0(n5361), .Y(P1_U3221));
  INVX1   g4246(.A(n5092), .Y(n5363));
  OAI22X1 g4247(.A0(n4242), .A1(n3282), .B0(n3294), .B1(n4247), .Y(n5364));
  XOR2X1  g4248(.A(n5364), .B(n4239), .Y(n5365));
  AOI22X1 g4249(.A0(n4241), .A1(n3281), .B0(n3333), .B1(n4248), .Y(n5366));
  NAND2X1 g4250(.A(n5366), .B(n5365), .Y(n5367));
  INVX1   g4251(.A(n5367), .Y(n5368));
  NOR4X1  g4252(.A(n5363), .B(n5076), .C(n5012), .D(n5368), .Y(n5369));
  AOI22X1 g4253(.A0(n4241), .A1(n3397), .B0(n3329), .B1(n4248), .Y(n5370));
  XOR2X1  g4254(.A(n5370), .B(n4246), .Y(n5371));
  OAI22X1 g4255(.A0(n4242), .A1(n3322), .B0(n3358), .B1(n4247), .Y(n5372));
  XOR2X1  g4256(.A(n5372), .B(n5371), .Y(n5373));
  NOR2X1  g4257(.A(n5363), .B(n5084), .Y(n5374));
  NOR2X1  g4258(.A(n5366), .B(n5365), .Y(n5375));
  AOI21X1 g4259(.A0(n5374), .A1(n5367), .B0(n5375), .Y(n5376));
  OAI21X1 g4260(.A0(n5368), .A1(n5091), .B0(n5376), .Y(n5377));
  NOR3X1  g4261(.A(n5377), .B(n5373), .C(n5369), .Y(n5378));
  NAND3X1 g4262(.A(n5092), .B(n5139), .C(n5094), .Y(n5379));
  NOR3X1  g4263(.A(n5375), .B(n5374), .C(n5090), .Y(n5380));
  NAND2X1 g4264(.A(n5373), .B(n5367), .Y(n5381));
  AOI21X1 g4265(.A0(n5380), .A1(n5379), .B0(n5381), .Y(n5382));
  OAI21X1 g4266(.A0(n5382), .A1(n5378), .B0(n5143), .Y(n5383));
  NAND3X1 g4267(.A(n5150), .B(n3119), .C(n3392), .Y(n5384));
  AOI22X1 g4268(.A0(n4988), .A1(n3317), .B0(n3363), .B1(n4998), .Y(n5385));
  OAI21X1 g4269(.A0(n5153), .A1(n3282), .B0(n5385), .Y(n5386));
  OAI22X1 g4270(.A0(n3316), .A1(n4993), .B0(P1_STATE_REG_SCAN_IN), .B1(n3314), .Y(n5387));
  AOI21X1 g4271(.A0(n5386), .A1(n4995), .B0(n5387), .Y(n5388));
  NAND3X1 g4272(.A(n5388), .B(n5384), .C(n5383), .Y(P1_U3220));
  INVX1   g4273(.A(n5029), .Y(n5390));
  XOR2X1  g4274(.A(n5031), .B(n5390), .Y(n5391));
  NOR2X1  g4275(.A(n5391), .B(n5070), .Y(n5392));
  AOI21X1 g4276(.A0(n5071), .A1(n5033), .B0(n5135), .Y(n5393));
  OAI21X1 g4277(.A0(n5393), .A1(n5392), .B0(n5143), .Y(n5394));
  AOI22X1 g4278(.A0(n4988), .A1(n2929), .B0(n3001), .B1(n4998), .Y(n5395));
  OAI21X1 g4279(.A0(n5153), .A1(n2891), .B0(n5395), .Y(n5396));
  AOI22X1 g4280(.A0(n4995), .A1(n5396), .B0(P1_U3086), .B1(P1_REG3_REG_19__SCAN_IN), .Y(n5397));
  OAI21X1 g4281(.A0(n4993), .A1(n2928), .B0(n5397), .Y(n5398));
  AOI21X1 g4282(.A0(n5150), .A1(n2941), .B0(n5398), .Y(n5399));
  NAND2X1 g4283(.A(n5399), .B(n5394), .Y(P1_U3219));
  AOI21X1 g4284(.A0(n5109), .A1(n4946), .B0(n5110), .Y(n5401));
  OAI21X1 g4285(.A0(n5182), .A1(n4943), .B0(n5401), .Y(n5402));
  OAI22X1 g4286(.A0(n4946), .A1(n4932), .B0(n4929), .B1(n4927), .Y(n5403));
  AOI21X1 g4287(.A0(n4932), .A1(n4946), .B0(n5403), .Y(n5404));
  OAI21X1 g4288(.A0(n5120), .A1(n5181), .B0(n5404), .Y(n5405));
  NAND3X1 g4289(.A(n5405), .B(n5402), .C(n5143), .Y(n5406));
  OAI22X1 g4290(.A0(n4981), .A1(P1_REG3_REG_3__SCAN_IN), .B0(n2103), .B1(n5153), .Y(n5407));
  AOI21X1 g4291(.A0(n4998), .A1(n2219), .B0(n5407), .Y(n5408));
  AOI22X1 g4292(.A0(n2169), .A1(n5150), .B0(P1_U3086), .B1(P1_REG3_REG_3__SCAN_IN), .Y(n5409));
  OAI21X1 g4293(.A0(n5408), .A1(n4996), .B0(n5409), .Y(n5410));
  AOI21X1 g4294(.A0(n5157), .A1(n2158), .B0(n5410), .Y(n5411));
  NAND2X1 g4295(.A(n5411), .B(n5406), .Y(P1_U3218));
  XOR2X1  g4296(.A(n4895), .B(n4893), .Y(n5413));
  XOR2X1  g4297(.A(n5413), .B(n5129), .Y(n5414));
  OAI22X1 g4298(.A0(n4981), .A1(n2499), .B0(n2458), .B1(n5153), .Y(n5415));
  AOI21X1 g4299(.A0(n4998), .A1(n2580), .B0(n5415), .Y(n5416));
  AOI22X1 g4300(.A0(n2516), .A1(n5150), .B0(P1_U3086), .B1(P1_REG3_REG_10__SCAN_IN), .Y(n5417));
  OAI21X1 g4301(.A0(n5416), .A1(n4996), .B0(n5417), .Y(n5418));
  AOI21X1 g4302(.A0(n5157), .A1(n2500), .B0(n5418), .Y(n5419));
  OAI21X1 g4303(.A0(n5414), .A1(n4987), .B0(n5419), .Y(P1_U3217));
  XOR2X1  g4304(.A(n5015), .B(n5013), .Y(n5421));
  XOR2X1  g4305(.A(n5421), .B(n5138), .Y(n5422));
  NOR2X1  g4306(.A(n4999), .B(n3150), .Y(n5423));
  OAI22X1 g4307(.A0(n4981), .A1(n3105), .B0(n3071), .B1(n5153), .Y(n5424));
  OAI21X1 g4308(.A0(n5424), .A1(n5423), .B0(n4995), .Y(n5425));
  INVX1   g4309(.A(n3105), .Y(n5426));
  AOI22X1 g4310(.A0(n5426), .A1(n5157), .B0(P1_U3086), .B1(P1_REG3_REG_23__SCAN_IN), .Y(n5427));
  NAND2X1 g4311(.A(n5427), .B(n5425), .Y(n5428));
  AOI21X1 g4312(.A0(n5150), .A1(n3142), .B0(n5428), .Y(n5429));
  OAI21X1 g4313(.A0(n5422), .A1(n4987), .B0(n5429), .Y(P1_U3216));
  XOR2X1  g4314(.A(n4869), .B(n4867), .Y(n5431));
  XOR2X1  g4315(.A(n5431), .B(n5131), .Y(n5432));
  OAI22X1 g4316(.A0(n4981), .A1(n2697), .B0(n2798), .B1(n4999), .Y(n5433));
  AOI21X1 g4317(.A0(n4997), .A1(n2649), .B0(n5433), .Y(n5434));
  AOI22X1 g4318(.A0(n2741), .A1(n5150), .B0(P1_U3086), .B1(P1_REG3_REG_14__SCAN_IN), .Y(n5435));
  OAI21X1 g4319(.A0(n5434), .A1(n4996), .B0(n5435), .Y(n5436));
  AOI21X1 g4320(.A0(n5157), .A1(n2698), .B0(n5436), .Y(n5437));
  OAI21X1 g4321(.A0(n5432), .A1(n4987), .B0(n5437), .Y(P1_U3215));
  NOR3X1  g4322(.A(n5363), .B(n5076), .C(n5012), .Y(n5439));
  INVX1   g4323(.A(n5366), .Y(n5440));
  XOR2X1  g4324(.A(n5440), .B(n5365), .Y(n5441));
  NOR4X1  g4325(.A(n5439), .B(n5374), .C(n5090), .D(n5441), .Y(n5442));
  NOR2X1  g4326(.A(n5374), .B(n5090), .Y(n5443));
  INVX1   g4327(.A(n5441), .Y(n5444));
  AOI21X1 g4328(.A0(n5443), .A1(n5379), .B0(n5444), .Y(n5445));
  OAI21X1 g4329(.A0(n5445), .A1(n5442), .B0(n5143), .Y(n5446));
  NAND2X1 g4330(.A(n5150), .B(n3333), .Y(n5447));
  AOI22X1 g4331(.A0(n4988), .A1(n3731), .B0(n3235), .B1(n4997), .Y(n5448));
  OAI21X1 g4332(.A0(n4999), .A1(n3322), .B0(n5448), .Y(n5449));
  OAI22X1 g4333(.A0(n3277), .A1(n4993), .B0(P1_STATE_REG_SCAN_IN), .B1(n3275), .Y(n5450));
  AOI21X1 g4334(.A0(n5449), .A1(n4995), .B0(n5450), .Y(n5451));
  NAND3X1 g4335(.A(n5451), .B(n5447), .C(n5446), .Y(P1_U3214));
  OAI21X1 g4336(.A0(n4914), .A1(n4912), .B0(n4915), .Y(n5453));
  AOI21X1 g4337(.A0(n4956), .A1(n4954), .B0(n5453), .Y(n5454));
  AOI21X1 g4338(.A0(n4911), .A1(n4909), .B0(n4954), .Y(n5455));
  AOI21X1 g4339(.A0(n4958), .A1(n4912), .B0(n4955), .Y(n5456));
  OAI21X1 g4340(.A0(n4958), .A1(n4912), .B0(n5456), .Y(n5457));
  OAI21X1 g4341(.A0(n5457), .A1(n5455), .B0(n5143), .Y(n5458));
  OAI22X1 g4342(.A0(n4981), .A1(n2359), .B0(n2312), .B1(n5153), .Y(n5459));
  AOI21X1 g4343(.A0(n4998), .A1(n2408), .B0(n5459), .Y(n5460));
  AOI22X1 g4344(.A0(n2376), .A1(n5150), .B0(P1_U3086), .B1(P1_REG3_REG_7__SCAN_IN), .Y(n5461));
  OAI21X1 g4345(.A0(n5460), .A1(n4996), .B0(n5461), .Y(n5462));
  AOI21X1 g4346(.A0(n5157), .A1(n2360), .B0(n5462), .Y(n5463));
  OAI21X1 g4347(.A0(n5458), .A1(n5454), .B0(n5463), .Y(P1_U3213));
  AOI21X1 g4348(.A0(n1144), .A1(n1142), .B0(n1166), .Y(n5465));
  AOI21X1 g4349(.A0(n1155), .A1(n1152), .B0(n5465), .Y(n5466));
  NAND2X1 g4350(.A(P2_IR_REG_0__SCAN_IN), .B(P2_STATE_REG_SCAN_IN), .Y(n5467));
  OAI21X1 g4351(.A0(n5466), .A1(P2_STATE_REG_SCAN_IN), .B0(n5467), .Y(P2_U3295));
  AOI21X1 g4352(.A0(n1144), .A1(n1142), .B0(n1163), .Y(n5469));
  AOI21X1 g4353(.A0(n1179), .A1(n1152), .B0(n5469), .Y(n5470));
  INVX1   g4354(.A(P2_STATE_REG_SCAN_IN), .Y(P2_U3151));
  NOR2X1  g4355(.A(P2_IR_REG_31__SCAN_IN), .B(P2_U3151), .Y(n5472));
  INVX1   g4356(.A(P2_IR_REG_31__SCAN_IN), .Y(n5473));
  NOR2X1  g4357(.A(n5473), .B(P2_U3151), .Y(n5474));
  XOR2X1  g4358(.A(P2_IR_REG_1__SCAN_IN), .B(P2_IR_REG_0__SCAN_IN), .Y(n5475));
  AOI22X1 g4359(.A0(n5474), .A1(n5475), .B0(n5472), .B1(P2_IR_REG_1__SCAN_IN), .Y(n5476));
  OAI21X1 g4360(.A0(n5470), .A1(P2_STATE_REG_SCAN_IN), .B0(n5476), .Y(P2_U3294));
  AOI21X1 g4361(.A0(n1144), .A1(n1142), .B0(n1286), .Y(n5478));
  AOI21X1 g4362(.A0(n1195), .A1(n1152), .B0(n5478), .Y(n5479));
  INVX1   g4363(.A(P2_IR_REG_2__SCAN_IN), .Y(n5480));
  NOR2X1  g4364(.A(P2_IR_REG_1__SCAN_IN), .B(P2_IR_REG_0__SCAN_IN), .Y(n5481));
  XOR2X1  g4365(.A(n5481), .B(n5480), .Y(n5482));
  AOI22X1 g4366(.A0(n5474), .A1(n5482), .B0(n5472), .B1(P2_IR_REG_2__SCAN_IN), .Y(n5483));
  OAI21X1 g4367(.A0(n5479), .A1(P2_STATE_REG_SCAN_IN), .B0(n5483), .Y(P2_U3293));
  AOI21X1 g4368(.A0(n1144), .A1(n1142), .B0(n1289), .Y(n5485));
  AOI21X1 g4369(.A0(n1210), .A1(n1152), .B0(n5485), .Y(n5486));
  INVX1   g4370(.A(P2_IR_REG_3__SCAN_IN), .Y(n5487));
  NOR3X1  g4371(.A(P2_IR_REG_2__SCAN_IN), .B(P2_IR_REG_1__SCAN_IN), .C(P2_IR_REG_0__SCAN_IN), .Y(n5488));
  XOR2X1  g4372(.A(n5488), .B(n5487), .Y(n5489));
  AOI22X1 g4373(.A0(n5474), .A1(n5489), .B0(n5472), .B1(P2_IR_REG_3__SCAN_IN), .Y(n5490));
  OAI21X1 g4374(.A0(n5486), .A1(P2_STATE_REG_SCAN_IN), .B0(n5490), .Y(P2_U3292));
  AOI21X1 g4375(.A0(n1144), .A1(n1142), .B0(n1229), .Y(n5492));
  AOI21X1 g4376(.A0(n1234), .A1(n1152), .B0(n5492), .Y(n5493));
  INVX1   g4377(.A(P2_IR_REG_4__SCAN_IN), .Y(n5494));
  NOR4X1  g4378(.A(P2_IR_REG_2__SCAN_IN), .B(P2_IR_REG_1__SCAN_IN), .C(P2_IR_REG_0__SCAN_IN), .D(P2_IR_REG_3__SCAN_IN), .Y(n5495));
  XOR2X1  g4379(.A(n5495), .B(n5494), .Y(n5496));
  AOI22X1 g4380(.A0(n5474), .A1(n5496), .B0(n5472), .B1(P2_IR_REG_4__SCAN_IN), .Y(n5497));
  OAI21X1 g4381(.A0(n5493), .A1(P2_STATE_REG_SCAN_IN), .B0(n5497), .Y(P2_U3291));
  AOI21X1 g4382(.A0(n1144), .A1(n1142), .B0(n1250), .Y(n5499));
  AOI21X1 g4383(.A0(n1255), .A1(n1152), .B0(n5499), .Y(n5500));
  NAND2X1 g4384(.A(n5495), .B(n5494), .Y(n5501));
  XOR2X1  g4385(.A(n5501), .B(P2_IR_REG_5__SCAN_IN), .Y(n5502));
  AOI22X1 g4386(.A0(n5474), .A1(n5502), .B0(n5472), .B1(P2_IR_REG_5__SCAN_IN), .Y(n5503));
  OAI21X1 g4387(.A0(n5500), .A1(P2_STATE_REG_SCAN_IN), .B0(n5503), .Y(P2_U3290));
  AOI21X1 g4388(.A0(n1144), .A1(n1142), .B0(n1269), .Y(n5505));
  AOI21X1 g4389(.A0(n1274), .A1(n1152), .B0(n5505), .Y(n5506));
  INVX1   g4390(.A(P2_IR_REG_5__SCAN_IN), .Y(n5507));
  NAND3X1 g4391(.A(n5495), .B(n5507), .C(n5494), .Y(n5508));
  INVX1   g4392(.A(P2_IR_REG_6__SCAN_IN), .Y(n5509));
  NAND2X1 g4393(.A(n5509), .B(n5507), .Y(n5510));
  NOR2X1  g4394(.A(n5510), .B(n5501), .Y(n5511));
  AOI21X1 g4395(.A0(n5508), .A1(P2_IR_REG_6__SCAN_IN), .B0(n5511), .Y(n5512));
  AOI22X1 g4396(.A0(n5474), .A1(n5512), .B0(n5472), .B1(P2_IR_REG_6__SCAN_IN), .Y(n5513));
  OAI21X1 g4397(.A0(n5506), .A1(P2_STATE_REG_SCAN_IN), .B0(n5513), .Y(P2_U3289));
  AOI21X1 g4398(.A0(n1144), .A1(n1142), .B0(n1309), .Y(n5515));
  AOI21X1 g4399(.A0(n1314), .A1(n1152), .B0(n5515), .Y(n5516));
  INVX1   g4400(.A(P2_IR_REG_7__SCAN_IN), .Y(n5517));
  XOR2X1  g4401(.A(n5511), .B(n5517), .Y(n5518));
  AOI22X1 g4402(.A0(n5474), .A1(n5518), .B0(n5472), .B1(P2_IR_REG_7__SCAN_IN), .Y(n5519));
  OAI21X1 g4403(.A0(n5516), .A1(P2_STATE_REG_SCAN_IN), .B0(n5519), .Y(P2_U3288));
  INVX1   g4404(.A(P1_DATAO_REG_8__SCAN_IN), .Y(n5521));
  AOI21X1 g4405(.A0(n1144), .A1(n1142), .B0(n5521), .Y(n5522));
  AOI21X1 g4406(.A0(n1335), .A1(n1152), .B0(n5522), .Y(n5523));
  INVX1   g4407(.A(P2_IR_REG_8__SCAN_IN), .Y(n5524));
  AOI21X1 g4408(.A0(n5511), .A1(n5517), .B0(n5524), .Y(n5525));
  NOR4X1  g4409(.A(P2_IR_REG_7__SCAN_IN), .B(P2_IR_REG_6__SCAN_IN), .C(P2_IR_REG_5__SCAN_IN), .D(P2_IR_REG_8__SCAN_IN), .Y(n5526));
  NAND3X1 g4410(.A(n5526), .B(n5495), .C(n5494), .Y(n5527));
  INVX1   g4411(.A(n5527), .Y(n5528));
  NOR2X1  g4412(.A(n5528), .B(n5525), .Y(n5529));
  AOI22X1 g4413(.A0(n5474), .A1(n5529), .B0(n5472), .B1(P2_IR_REG_8__SCAN_IN), .Y(n5530));
  OAI21X1 g4414(.A0(n5523), .A1(P2_STATE_REG_SCAN_IN), .B0(n5530), .Y(P2_U3287));
  AOI21X1 g4415(.A0(n1144), .A1(n1142), .B0(n1367), .Y(n5532));
  AOI21X1 g4416(.A0(n1359), .A1(n1152), .B0(n5532), .Y(n5533));
  XOR2X1  g4417(.A(n5527), .B(P2_IR_REG_9__SCAN_IN), .Y(n5534));
  AOI22X1 g4418(.A0(n5474), .A1(n5534), .B0(n5472), .B1(P2_IR_REG_9__SCAN_IN), .Y(n5535));
  OAI21X1 g4419(.A0(n5533), .A1(P2_STATE_REG_SCAN_IN), .B0(n5535), .Y(P2_U3286));
  AOI21X1 g4420(.A0(n1144), .A1(n1142), .B0(n1389), .Y(n5537));
  AOI21X1 g4421(.A0(n1379), .A1(n1152), .B0(n5537), .Y(n5538));
  INVX1   g4422(.A(P2_IR_REG_9__SCAN_IN), .Y(n5539));
  NAND4X1 g4423(.A(n5495), .B(n5539), .C(n5494), .D(n5526), .Y(n5540));
  NOR3X1  g4424(.A(n5527), .B(P2_IR_REG_10__SCAN_IN), .C(P2_IR_REG_9__SCAN_IN), .Y(n5541));
  AOI21X1 g4425(.A0(n5540), .A1(P2_IR_REG_10__SCAN_IN), .B0(n5541), .Y(n5542));
  AOI22X1 g4426(.A0(n5474), .A1(n5542), .B0(n5472), .B1(P2_IR_REG_10__SCAN_IN), .Y(n5543));
  OAI21X1 g4427(.A0(n5538), .A1(P2_STATE_REG_SCAN_IN), .B0(n5543), .Y(P2_U3285));
  AOI21X1 g4428(.A0(n1144), .A1(n1142), .B0(n1414), .Y(n5545));
  AOI21X1 g4429(.A0(n1402), .A1(n1152), .B0(n5545), .Y(n5546));
  INVX1   g4430(.A(P2_IR_REG_11__SCAN_IN), .Y(n5547));
  XOR2X1  g4431(.A(n5541), .B(n5547), .Y(n5548));
  AOI22X1 g4432(.A0(n5474), .A1(n5548), .B0(n5472), .B1(P2_IR_REG_11__SCAN_IN), .Y(n5549));
  OAI21X1 g4433(.A0(n5546), .A1(P2_STATE_REG_SCAN_IN), .B0(n5549), .Y(P2_U3284));
  OAI21X1 g4434(.A0(n1149), .A1(n1148), .B0(P1_DATAO_REG_12__SCAN_IN), .Y(n5551));
  INVX1   g4435(.A(n5551), .Y(n5552));
  AOI21X1 g4436(.A0(n1423), .A1(n1152), .B0(n5552), .Y(n5553));
  INVX1   g4437(.A(P2_IR_REG_12__SCAN_IN), .Y(n5554));
  AOI21X1 g4438(.A0(n5541), .A1(n5547), .B0(n5554), .Y(n5555));
  NOR4X1  g4439(.A(P2_IR_REG_11__SCAN_IN), .B(P2_IR_REG_10__SCAN_IN), .C(P2_IR_REG_9__SCAN_IN), .D(P2_IR_REG_12__SCAN_IN), .Y(n5556));
  NAND4X1 g4440(.A(n5526), .B(n5495), .C(n5494), .D(n5556), .Y(n5557));
  INVX1   g4441(.A(n5557), .Y(n5558));
  NOR2X1  g4442(.A(n5558), .B(n5555), .Y(n5559));
  AOI22X1 g4443(.A0(n5474), .A1(n5559), .B0(n5472), .B1(P2_IR_REG_12__SCAN_IN), .Y(n5560));
  OAI21X1 g4444(.A0(n5553), .A1(P2_STATE_REG_SCAN_IN), .B0(n5560), .Y(P2_U3283));
  AOI21X1 g4445(.A0(n1144), .A1(n1142), .B0(n1438), .Y(n5562));
  AOI21X1 g4446(.A0(n1442), .A1(n1152), .B0(n5562), .Y(n5563));
  XOR2X1  g4447(.A(n5557), .B(P2_IR_REG_13__SCAN_IN), .Y(n5564));
  AOI22X1 g4448(.A0(n5474), .A1(n5564), .B0(n5472), .B1(P2_IR_REG_13__SCAN_IN), .Y(n5565));
  OAI21X1 g4449(.A0(n5563), .A1(P2_STATE_REG_SCAN_IN), .B0(n5565), .Y(P2_U3282));
  INVX1   g4450(.A(P1_DATAO_REG_14__SCAN_IN), .Y(n5567));
  AOI21X1 g4451(.A0(n1144), .A1(n1142), .B0(n5567), .Y(n5568));
  AOI21X1 g4452(.A0(n1460), .A1(n1152), .B0(n5568), .Y(n5569));
  INVX1   g4453(.A(P2_IR_REG_13__SCAN_IN), .Y(n5570));
  INVX1   g4454(.A(P2_IR_REG_14__SCAN_IN), .Y(n5571));
  AOI21X1 g4455(.A0(n5558), .A1(n5570), .B0(n5571), .Y(n5572));
  NOR3X1  g4456(.A(n5557), .B(P2_IR_REG_14__SCAN_IN), .C(P2_IR_REG_13__SCAN_IN), .Y(n5573));
  NOR2X1  g4457(.A(n5573), .B(n5572), .Y(n5574));
  AOI22X1 g4458(.A0(n5474), .A1(n5574), .B0(n5472), .B1(P2_IR_REG_14__SCAN_IN), .Y(n5575));
  OAI21X1 g4459(.A0(n5569), .A1(P2_STATE_REG_SCAN_IN), .B0(n5575), .Y(P2_U3281));
  OAI21X1 g4460(.A0(n1149), .A1(n1148), .B0(P1_DATAO_REG_15__SCAN_IN), .Y(n5577));
  INVX1   g4461(.A(n5577), .Y(n5578));
  AOI21X1 g4462(.A0(n1487), .A1(n1152), .B0(n5578), .Y(n5579));
  INVX1   g4463(.A(P2_IR_REG_15__SCAN_IN), .Y(n5580));
  XOR2X1  g4464(.A(n5573), .B(n5580), .Y(n5581));
  AOI22X1 g4465(.A0(n5474), .A1(n5581), .B0(n5472), .B1(P2_IR_REG_15__SCAN_IN), .Y(n5582));
  OAI21X1 g4466(.A0(n5579), .A1(P2_STATE_REG_SCAN_IN), .B0(n5582), .Y(P2_U3280));
  OAI21X1 g4467(.A0(n1149), .A1(n1148), .B0(P1_DATAO_REG_16__SCAN_IN), .Y(n5584));
  INVX1   g4468(.A(n5584), .Y(n5585));
  AOI21X1 g4469(.A0(n1507), .A1(n1152), .B0(n5585), .Y(n5586));
  INVX1   g4470(.A(P2_IR_REG_16__SCAN_IN), .Y(n5587));
  NOR4X1  g4471(.A(P2_IR_REG_15__SCAN_IN), .B(P2_IR_REG_14__SCAN_IN), .C(P2_IR_REG_13__SCAN_IN), .D(n5557), .Y(n5588));
  NOR4X1  g4472(.A(P2_IR_REG_15__SCAN_IN), .B(P2_IR_REG_14__SCAN_IN), .C(P2_IR_REG_13__SCAN_IN), .D(P2_IR_REG_16__SCAN_IN), .Y(n5589));
  NAND2X1 g4473(.A(n5589), .B(n5556), .Y(n5590));
  OAI22X1 g4474(.A0(n5588), .A1(n5587), .B0(n5527), .B1(n5590), .Y(n5591));
  INVX1   g4475(.A(n5591), .Y(n5592));
  AOI22X1 g4476(.A0(n5474), .A1(n5592), .B0(n5472), .B1(P2_IR_REG_16__SCAN_IN), .Y(n5593));
  OAI21X1 g4477(.A0(n5586), .A1(P2_STATE_REG_SCAN_IN), .B0(n5593), .Y(P2_U3279));
  OAI21X1 g4478(.A0(n1149), .A1(n1148), .B0(P1_DATAO_REG_17__SCAN_IN), .Y(n5595));
  INVX1   g4479(.A(n5595), .Y(n5596));
  AOI21X1 g4480(.A0(n1537), .A1(n1152), .B0(n5596), .Y(n5597));
  INVX1   g4481(.A(P2_IR_REG_17__SCAN_IN), .Y(n5598));
  NOR2X1  g4482(.A(n5590), .B(n5527), .Y(n5599));
  XOR2X1  g4483(.A(n5599), .B(n5598), .Y(n5600));
  AOI22X1 g4484(.A0(n5474), .A1(n5600), .B0(n5472), .B1(P2_IR_REG_17__SCAN_IN), .Y(n5601));
  OAI21X1 g4485(.A0(n5597), .A1(P2_STATE_REG_SCAN_IN), .B0(n5601), .Y(P2_U3278));
  OAI21X1 g4486(.A0(n1149), .A1(n1148), .B0(P1_DATAO_REG_18__SCAN_IN), .Y(n5603));
  INVX1   g4487(.A(n5603), .Y(n5604));
  AOI21X1 g4488(.A0(n1555), .A1(n1152), .B0(n5604), .Y(n5605));
  INVX1   g4489(.A(P2_IR_REG_18__SCAN_IN), .Y(n5606));
  NOR3X1  g4490(.A(n5590), .B(n5527), .C(P2_IR_REG_17__SCAN_IN), .Y(n5607));
  NOR4X1  g4491(.A(n5527), .B(P2_IR_REG_18__SCAN_IN), .C(P2_IR_REG_17__SCAN_IN), .D(n5590), .Y(n5608));
  INVX1   g4492(.A(n5608), .Y(n5609));
  OAI21X1 g4493(.A0(n5607), .A1(n5606), .B0(n5609), .Y(n5610));
  INVX1   g4494(.A(n5610), .Y(n5611));
  AOI22X1 g4495(.A0(n5474), .A1(n5611), .B0(n5472), .B1(P2_IR_REG_18__SCAN_IN), .Y(n5612));
  OAI21X1 g4496(.A0(n5605), .A1(P2_STATE_REG_SCAN_IN), .B0(n5612), .Y(P2_U3277));
  OAI21X1 g4497(.A0(n1149), .A1(n1148), .B0(P1_DATAO_REG_19__SCAN_IN), .Y(n5614));
  INVX1   g4498(.A(n5614), .Y(n5615));
  AOI21X1 g4499(.A0(n1583), .A1(n1152), .B0(n5615), .Y(n5616));
  INVX1   g4500(.A(P2_IR_REG_19__SCAN_IN), .Y(n5617));
  XOR2X1  g4501(.A(n5608), .B(n5617), .Y(n5618));
  AOI22X1 g4502(.A0(n5474), .A1(n5618), .B0(n5472), .B1(P2_IR_REG_19__SCAN_IN), .Y(n5619));
  OAI21X1 g4503(.A0(n5616), .A1(P2_STATE_REG_SCAN_IN), .B0(n5619), .Y(P2_U3276));
  OAI21X1 g4504(.A0(n1149), .A1(n1148), .B0(P1_DATAO_REG_20__SCAN_IN), .Y(n5621));
  INVX1   g4505(.A(n5621), .Y(n5622));
  AOI21X1 g4506(.A0(n1606), .A1(n1152), .B0(n5622), .Y(n5623));
  OAI21X1 g4507(.A0(n5609), .A1(P2_IR_REG_19__SCAN_IN), .B0(P2_IR_REG_20__SCAN_IN), .Y(n5624));
  NOR4X1  g4508(.A(P2_IR_REG_19__SCAN_IN), .B(P2_IR_REG_18__SCAN_IN), .C(P2_IR_REG_17__SCAN_IN), .D(P2_IR_REG_20__SCAN_IN), .Y(n5625));
  INVX1   g4509(.A(n5625), .Y(n5626));
  NOR3X1  g4510(.A(n5626), .B(n5590), .C(n5527), .Y(n5627));
  INVX1   g4511(.A(n5627), .Y(n5628));
  NAND2X1 g4512(.A(n5628), .B(n5624), .Y(n5629));
  NOR3X1  g4513(.A(n5629), .B(n5473), .C(P2_U3151), .Y(n5630));
  AOI21X1 g4514(.A0(n5472), .A1(P2_IR_REG_20__SCAN_IN), .B0(n5630), .Y(n5631));
  OAI21X1 g4515(.A0(n5623), .A1(P2_STATE_REG_SCAN_IN), .B0(n5631), .Y(P2_U3275));
  OAI21X1 g4516(.A0(n1149), .A1(n1148), .B0(P1_DATAO_REG_21__SCAN_IN), .Y(n5633));
  INVX1   g4517(.A(n5633), .Y(n5634));
  AOI21X1 g4518(.A0(n1631), .A1(n1152), .B0(n5634), .Y(n5635));
  INVX1   g4519(.A(P2_IR_REG_21__SCAN_IN), .Y(n5636));
  XOR2X1  g4520(.A(n5627), .B(n5636), .Y(n5637));
  AOI22X1 g4521(.A0(n5474), .A1(n5637), .B0(n5472), .B1(P2_IR_REG_21__SCAN_IN), .Y(n5638));
  OAI21X1 g4522(.A0(n5635), .A1(P2_STATE_REG_SCAN_IN), .B0(n5638), .Y(P2_U3274));
  OAI21X1 g4523(.A0(n1149), .A1(n1148), .B0(P1_DATAO_REG_22__SCAN_IN), .Y(n5640));
  INVX1   g4524(.A(n5640), .Y(n5641));
  AOI21X1 g4525(.A0(n1649), .A1(n1152), .B0(n5641), .Y(n5642));
  INVX1   g4526(.A(P2_IR_REG_22__SCAN_IN), .Y(n5643));
  AOI21X1 g4527(.A0(n5627), .A1(n5636), .B0(n5643), .Y(n5644));
  NOR2X1  g4528(.A(P2_IR_REG_22__SCAN_IN), .B(P2_IR_REG_21__SCAN_IN), .Y(n5645));
  AOI21X1 g4529(.A0(n5645), .A1(n5627), .B0(n5644), .Y(n5646));
  AOI22X1 g4530(.A0(n5474), .A1(n5646), .B0(n5472), .B1(P2_IR_REG_22__SCAN_IN), .Y(n5647));
  OAI21X1 g4531(.A0(n5642), .A1(P2_STATE_REG_SCAN_IN), .B0(n5647), .Y(P2_U3273));
  OAI21X1 g4532(.A0(n1149), .A1(n1148), .B0(P1_DATAO_REG_23__SCAN_IN), .Y(n5649));
  OAI21X1 g4533(.A0(n1672), .A1(n1145), .B0(n5649), .Y(n5650));
  INVX1   g4534(.A(n5650), .Y(n5651));
  INVX1   g4535(.A(P2_IR_REG_23__SCAN_IN), .Y(n5652));
  NOR3X1  g4536(.A(n5628), .B(P2_IR_REG_22__SCAN_IN), .C(P2_IR_REG_21__SCAN_IN), .Y(n5653));
  XOR2X1  g4537(.A(n5653), .B(n5652), .Y(n5654));
  AOI22X1 g4538(.A0(n5474), .A1(n5654), .B0(n5472), .B1(P2_IR_REG_23__SCAN_IN), .Y(n5655));
  OAI21X1 g4539(.A0(n5651), .A1(P2_STATE_REG_SCAN_IN), .B0(n5655), .Y(P2_U3272));
  OAI21X1 g4540(.A0(n1149), .A1(n1148), .B0(P1_DATAO_REG_24__SCAN_IN), .Y(n5657));
  OAI21X1 g4541(.A0(n3173), .A1(n1145), .B0(n5657), .Y(n5658));
  INVX1   g4542(.A(n5658), .Y(n5659));
  NAND3X1 g4543(.A(n5645), .B(n5627), .C(n5652), .Y(n5660));
  NOR4X1  g4544(.A(P2_IR_REG_23__SCAN_IN), .B(P2_IR_REG_22__SCAN_IN), .C(P2_IR_REG_21__SCAN_IN), .D(P2_IR_REG_24__SCAN_IN), .Y(n5661));
  NAND3X1 g4545(.A(n5661), .B(n5625), .C(n5599), .Y(n5662));
  INVX1   g4546(.A(n5662), .Y(n5663));
  AOI21X1 g4547(.A0(n5660), .A1(P2_IR_REG_24__SCAN_IN), .B0(n5663), .Y(n5664));
  AOI22X1 g4548(.A0(n5474), .A1(n5664), .B0(n5472), .B1(P2_IR_REG_24__SCAN_IN), .Y(n5665));
  OAI21X1 g4549(.A0(n5659), .A1(P2_STATE_REG_SCAN_IN), .B0(n5665), .Y(P2_U3271));
  OAI21X1 g4550(.A0(n1149), .A1(n1148), .B0(P1_DATAO_REG_25__SCAN_IN), .Y(n5667));
  INVX1   g4551(.A(n5667), .Y(n5668));
  AOI21X1 g4552(.A0(n1725), .A1(n1152), .B0(n5668), .Y(n5669));
  INVX1   g4553(.A(P2_IR_REG_25__SCAN_IN), .Y(n5670));
  XOR2X1  g4554(.A(n5662), .B(n5670), .Y(n5671));
  NOR3X1  g4555(.A(n5671), .B(n5473), .C(P2_U3151), .Y(n5672));
  AOI21X1 g4556(.A0(n5472), .A1(P2_IR_REG_25__SCAN_IN), .B0(n5672), .Y(n5673));
  OAI21X1 g4557(.A0(n5669), .A1(P2_STATE_REG_SCAN_IN), .B0(n5673), .Y(P2_U3270));
  OAI21X1 g4558(.A0(n1149), .A1(n1148), .B0(P1_DATAO_REG_26__SCAN_IN), .Y(n5675));
  INVX1   g4559(.A(n5675), .Y(n5676));
  AOI21X1 g4560(.A0(n1743), .A1(n1152), .B0(n5676), .Y(n5677));
  INVX1   g4561(.A(P2_IR_REG_26__SCAN_IN), .Y(n5678));
  AOI21X1 g4562(.A0(n5663), .A1(n5670), .B0(n5678), .Y(n5679));
  NAND2X1 g4563(.A(n5678), .B(n5670), .Y(n5680));
  NOR2X1  g4564(.A(n5680), .B(n5662), .Y(n5681));
  NOR2X1  g4565(.A(n5681), .B(n5679), .Y(n5682));
  AOI22X1 g4566(.A0(n5474), .A1(n5682), .B0(n5472), .B1(P2_IR_REG_26__SCAN_IN), .Y(n5683));
  OAI21X1 g4567(.A0(n5677), .A1(P2_STATE_REG_SCAN_IN), .B0(n5683), .Y(P2_U3269));
  AOI21X1 g4568(.A0(n1773), .A1(n1768), .B0(n1145), .Y(n5685));
  OAI21X1 g4569(.A0(n1149), .A1(n1148), .B0(P1_DATAO_REG_27__SCAN_IN), .Y(n5686));
  INVX1   g4570(.A(n5686), .Y(n5687));
  NOR2X1  g4571(.A(n5687), .B(n5685), .Y(n5688));
  XOR2X1  g4572(.A(n5681), .B(P2_IR_REG_27__SCAN_IN), .Y(n5689));
  INVX1   g4573(.A(n5689), .Y(n5690));
  AOI22X1 g4574(.A0(n5474), .A1(n5690), .B0(n5472), .B1(P2_IR_REG_27__SCAN_IN), .Y(n5691));
  OAI21X1 g4575(.A0(n5688), .A1(P2_STATE_REG_SCAN_IN), .B0(n5691), .Y(P2_U3268));
  OAI21X1 g4576(.A0(n1149), .A1(n1148), .B0(P1_DATAO_REG_28__SCAN_IN), .Y(n5693));
  INVX1   g4577(.A(n5693), .Y(n5694));
  AOI21X1 g4578(.A0(n1789), .A1(n1152), .B0(n5694), .Y(n5695));
  INVX1   g4579(.A(P2_IR_REG_28__SCAN_IN), .Y(n5696));
  NOR2X1  g4580(.A(n5681), .B(n5696), .Y(n5697));
  INVX1   g4581(.A(P2_IR_REG_27__SCAN_IN), .Y(n5698));
  NOR2X1  g4582(.A(n5696), .B(n5698), .Y(n5699));
  NOR4X1  g4583(.A(n5662), .B(P2_IR_REG_28__SCAN_IN), .C(P2_IR_REG_27__SCAN_IN), .D(n5680), .Y(n5700));
  NOR3X1  g4584(.A(n5700), .B(n5699), .C(n5697), .Y(n5701));
  AOI22X1 g4585(.A0(n5474), .A1(n5701), .B0(n5472), .B1(P2_IR_REG_28__SCAN_IN), .Y(n5702));
  OAI21X1 g4586(.A0(n5695), .A1(P2_STATE_REG_SCAN_IN), .B0(n5702), .Y(P2_U3267));
  OAI21X1 g4587(.A0(n1149), .A1(n1148), .B0(P1_DATAO_REG_29__SCAN_IN), .Y(n5704));
  INVX1   g4588(.A(n5704), .Y(n5705));
  AOI21X1 g4589(.A0(n1819), .A1(n1152), .B0(n5705), .Y(n5706));
  INVX1   g4590(.A(P2_IR_REG_29__SCAN_IN), .Y(n5707));
  XOR2X1  g4591(.A(n5700), .B(n5707), .Y(n5708));
  AOI22X1 g4592(.A0(n5474), .A1(n5708), .B0(n5472), .B1(P2_IR_REG_29__SCAN_IN), .Y(n5709));
  OAI21X1 g4593(.A0(n5706), .A1(P2_STATE_REG_SCAN_IN), .B0(n5709), .Y(P2_U3266));
  AOI21X1 g4594(.A0(n1844), .A1(n1839), .B0(n1145), .Y(n5711));
  OAI21X1 g4595(.A0(n1149), .A1(n1148), .B0(P1_DATAO_REG_30__SCAN_IN), .Y(n5712));
  INVX1   g4596(.A(n5712), .Y(n5713));
  NOR2X1  g4597(.A(n5713), .B(n5711), .Y(n5714));
  NAND2X1 g4598(.A(n5700), .B(n5707), .Y(n5715));
  XOR2X1  g4599(.A(n5715), .B(P2_IR_REG_30__SCAN_IN), .Y(n5716));
  AOI22X1 g4600(.A0(n5474), .A1(n5716), .B0(n5472), .B1(P2_IR_REG_30__SCAN_IN), .Y(n5717));
  OAI21X1 g4601(.A0(n5714), .A1(P2_STATE_REG_SCAN_IN), .B0(n5717), .Y(P2_U3265));
  NAND4X1 g4602(.A(n3767), .B(n3766), .C(n1152), .D(n1864), .Y(n5719));
  OAI21X1 g4603(.A0(n1149), .A1(n1148), .B0(P1_DATAO_REG_31__SCAN_IN), .Y(n5720));
  NAND2X1 g4604(.A(n5720), .B(n5719), .Y(n5721));
  NAND2X1 g4605(.A(n5721), .B(P2_U3151), .Y(n5722));
  NOR2X1  g4606(.A(n5715), .B(P2_IR_REG_30__SCAN_IN), .Y(n5723));
  NAND3X1 g4607(.A(n5723), .B(P2_IR_REG_31__SCAN_IN), .C(P2_STATE_REG_SCAN_IN), .Y(n5724));
  NAND2X1 g4608(.A(n5724), .B(n5722), .Y(P2_U3264));
  INVX1   g4609(.A(P2_D_REG_0__SCAN_IN), .Y(n5726));
  NOR2X1  g4610(.A(P2_IR_REG_31__SCAN_IN), .B(n5652), .Y(n5727));
  AOI21X1 g4611(.A0(n5654), .A1(P2_IR_REG_31__SCAN_IN), .B0(n5727), .Y(n5728));
  INVX1   g4612(.A(n5728), .Y(n5729));
  NAND2X1 g4613(.A(n5473), .B(P2_IR_REG_24__SCAN_IN), .Y(n5730));
  INVX1   g4614(.A(n5730), .Y(n5731));
  AOI21X1 g4615(.A0(n5664), .A1(P2_IR_REG_31__SCAN_IN), .B0(n5731), .Y(n5732));
  NOR2X1  g4616(.A(P2_IR_REG_31__SCAN_IN), .B(n5670), .Y(n5733));
  INVX1   g4617(.A(n5733), .Y(n5734));
  OAI21X1 g4618(.A0(n5671), .A1(n5473), .B0(n5734), .Y(n5735));
  INVX1   g4619(.A(n5735), .Y(n5736));
  NOR2X1  g4620(.A(P2_IR_REG_31__SCAN_IN), .B(n5678), .Y(n5737));
  AOI21X1 g4621(.A0(n5682), .A1(P2_IR_REG_31__SCAN_IN), .B0(n5737), .Y(n5738));
  NOR3X1  g4622(.A(n5738), .B(n5736), .C(n5732), .Y(n5739));
  XOR2X1  g4623(.A(n5732), .B(P2_B_REG_SCAN_IN), .Y(n5740));
  NOR3X1  g4624(.A(n5740), .B(n5738), .C(n5735), .Y(n5741));
  NOR2X1  g4625(.A(n5741), .B(n5738), .Y(n5742));
  NOR4X1  g4626(.A(n5739), .B(n5729), .C(P2_U3151), .D(n5742), .Y(n5743));
  NOR3X1  g4627(.A(n5739), .B(n5729), .C(P2_U3151), .Y(n5744));
  NOR3X1  g4628(.A(n5681), .B(n5679), .C(n5473), .Y(n5745));
  OAI22X1 g4629(.A0(n5737), .A1(n5745), .B0(n5735), .B1(n5740), .Y(n5746));
  OAI21X1 g4630(.A0(n5738), .A1(n5735), .B0(n5732), .Y(n5747));
  NAND3X1 g4631(.A(n5747), .B(n5746), .C(n5744), .Y(n5748));
  OAI21X1 g4632(.A0(n5743), .A1(n5726), .B0(n5748), .Y(P2_U3376));
  INVX1   g4633(.A(P2_D_REG_1__SCAN_IN), .Y(n5750));
  NAND2X1 g4634(.A(n5738), .B(n5736), .Y(n5751));
  NAND3X1 g4635(.A(n5751), .B(n5746), .C(n5744), .Y(n5752));
  OAI21X1 g4636(.A0(n5743), .A1(n5750), .B0(n5752), .Y(P2_U3377));
  INVX1   g4637(.A(P2_D_REG_2__SCAN_IN), .Y(n5754));
  AOI21X1 g4638(.A0(n5746), .A1(n5744), .B0(n5754), .Y(P2_U3263));
  INVX1   g4639(.A(P2_D_REG_3__SCAN_IN), .Y(n5756));
  AOI21X1 g4640(.A0(n5746), .A1(n5744), .B0(n5756), .Y(P2_U3262));
  INVX1   g4641(.A(P2_D_REG_4__SCAN_IN), .Y(n5758));
  AOI21X1 g4642(.A0(n5746), .A1(n5744), .B0(n5758), .Y(P2_U3261));
  INVX1   g4643(.A(P2_D_REG_5__SCAN_IN), .Y(n5760));
  AOI21X1 g4644(.A0(n5746), .A1(n5744), .B0(n5760), .Y(P2_U3260));
  INVX1   g4645(.A(P2_D_REG_6__SCAN_IN), .Y(n5762));
  AOI21X1 g4646(.A0(n5746), .A1(n5744), .B0(n5762), .Y(P2_U3259));
  INVX1   g4647(.A(P2_D_REG_7__SCAN_IN), .Y(n5764));
  AOI21X1 g4648(.A0(n5746), .A1(n5744), .B0(n5764), .Y(P2_U3258));
  INVX1   g4649(.A(P2_D_REG_8__SCAN_IN), .Y(n5766));
  AOI21X1 g4650(.A0(n5746), .A1(n5744), .B0(n5766), .Y(P2_U3257));
  INVX1   g4651(.A(P2_D_REG_9__SCAN_IN), .Y(n5768));
  AOI21X1 g4652(.A0(n5746), .A1(n5744), .B0(n5768), .Y(P2_U3256));
  INVX1   g4653(.A(P2_D_REG_10__SCAN_IN), .Y(n5770));
  AOI21X1 g4654(.A0(n5746), .A1(n5744), .B0(n5770), .Y(P2_U3255));
  INVX1   g4655(.A(P2_D_REG_11__SCAN_IN), .Y(n5772));
  AOI21X1 g4656(.A0(n5746), .A1(n5744), .B0(n5772), .Y(P2_U3254));
  INVX1   g4657(.A(P2_D_REG_12__SCAN_IN), .Y(n5774));
  AOI21X1 g4658(.A0(n5746), .A1(n5744), .B0(n5774), .Y(P2_U3253));
  INVX1   g4659(.A(P2_D_REG_13__SCAN_IN), .Y(n5776));
  AOI21X1 g4660(.A0(n5746), .A1(n5744), .B0(n5776), .Y(P2_U3252));
  INVX1   g4661(.A(P2_D_REG_14__SCAN_IN), .Y(n5778));
  AOI21X1 g4662(.A0(n5746), .A1(n5744), .B0(n5778), .Y(P2_U3251));
  INVX1   g4663(.A(P2_D_REG_15__SCAN_IN), .Y(n5780));
  AOI21X1 g4664(.A0(n5746), .A1(n5744), .B0(n5780), .Y(P2_U3250));
  INVX1   g4665(.A(P2_D_REG_16__SCAN_IN), .Y(n5782));
  AOI21X1 g4666(.A0(n5746), .A1(n5744), .B0(n5782), .Y(P2_U3249));
  INVX1   g4667(.A(P2_D_REG_17__SCAN_IN), .Y(n5784));
  AOI21X1 g4668(.A0(n5746), .A1(n5744), .B0(n5784), .Y(P2_U3248));
  INVX1   g4669(.A(P2_D_REG_18__SCAN_IN), .Y(n5786));
  AOI21X1 g4670(.A0(n5746), .A1(n5744), .B0(n5786), .Y(P2_U3247));
  INVX1   g4671(.A(P2_D_REG_19__SCAN_IN), .Y(n5788));
  AOI21X1 g4672(.A0(n5746), .A1(n5744), .B0(n5788), .Y(P2_U3246));
  INVX1   g4673(.A(P2_D_REG_20__SCAN_IN), .Y(n5790));
  AOI21X1 g4674(.A0(n5746), .A1(n5744), .B0(n5790), .Y(P2_U3245));
  INVX1   g4675(.A(P2_D_REG_21__SCAN_IN), .Y(n5792));
  AOI21X1 g4676(.A0(n5746), .A1(n5744), .B0(n5792), .Y(P2_U3244));
  INVX1   g4677(.A(P2_D_REG_22__SCAN_IN), .Y(n5794));
  AOI21X1 g4678(.A0(n5746), .A1(n5744), .B0(n5794), .Y(P2_U3243));
  INVX1   g4679(.A(P2_D_REG_23__SCAN_IN), .Y(n5796));
  AOI21X1 g4680(.A0(n5746), .A1(n5744), .B0(n5796), .Y(P2_U3242));
  INVX1   g4681(.A(P2_D_REG_24__SCAN_IN), .Y(n5798));
  AOI21X1 g4682(.A0(n5746), .A1(n5744), .B0(n5798), .Y(P2_U3241));
  INVX1   g4683(.A(P2_D_REG_25__SCAN_IN), .Y(n5800));
  AOI21X1 g4684(.A0(n5746), .A1(n5744), .B0(n5800), .Y(P2_U3240));
  INVX1   g4685(.A(P2_D_REG_26__SCAN_IN), .Y(n5802));
  AOI21X1 g4686(.A0(n5746), .A1(n5744), .B0(n5802), .Y(P2_U3239));
  INVX1   g4687(.A(P2_D_REG_27__SCAN_IN), .Y(n5804));
  AOI21X1 g4688(.A0(n5746), .A1(n5744), .B0(n5804), .Y(P2_U3238));
  INVX1   g4689(.A(P2_D_REG_28__SCAN_IN), .Y(n5806));
  AOI21X1 g4690(.A0(n5746), .A1(n5744), .B0(n5806), .Y(P2_U3237));
  INVX1   g4691(.A(P2_D_REG_29__SCAN_IN), .Y(n5808));
  AOI21X1 g4692(.A0(n5746), .A1(n5744), .B0(n5808), .Y(P2_U3236));
  INVX1   g4693(.A(P2_D_REG_30__SCAN_IN), .Y(n5810));
  AOI21X1 g4694(.A0(n5746), .A1(n5744), .B0(n5810), .Y(P2_U3235));
  INVX1   g4695(.A(P2_D_REG_31__SCAN_IN), .Y(n5812));
  AOI21X1 g4696(.A0(n5746), .A1(n5744), .B0(n5812), .Y(P2_U3234));
  INVX1   g4697(.A(P2_REG0_REG_0__SCAN_IN), .Y(n5814));
  INVX1   g4698(.A(n5744), .Y(n5815));
  OAI21X1 g4699(.A0(P2_D_REG_7__SCAN_IN), .A1(P2_D_REG_3__SCAN_IN), .B0(n5742), .Y(n5816));
  OAI21X1 g4700(.A0(P2_D_REG_9__SCAN_IN), .A1(P2_D_REG_8__SCAN_IN), .B0(n5742), .Y(n5817));
  OAI21X1 g4701(.A0(P2_D_REG_10__SCAN_IN), .A1(P2_D_REG_5__SCAN_IN), .B0(n5742), .Y(n5818));
  OAI21X1 g4702(.A0(P2_D_REG_6__SCAN_IN), .A1(P2_D_REG_4__SCAN_IN), .B0(n5742), .Y(n5819));
  NAND4X1 g4703(.A(n5818), .B(n5817), .C(n5816), .D(n5819), .Y(n5820));
  OAI21X1 g4704(.A0(P2_D_REG_28__SCAN_IN), .A1(P2_D_REG_27__SCAN_IN), .B0(n5742), .Y(n5821));
  OAI21X1 g4705(.A0(P2_D_REG_26__SCAN_IN), .A1(P2_D_REG_25__SCAN_IN), .B0(n5742), .Y(n5822));
  OAI21X1 g4706(.A0(P2_D_REG_31__SCAN_IN), .A1(P2_D_REG_30__SCAN_IN), .B0(n5742), .Y(n5823));
  OAI21X1 g4707(.A0(P2_D_REG_29__SCAN_IN), .A1(P2_D_REG_2__SCAN_IN), .B0(n5742), .Y(n5824));
  NAND4X1 g4708(.A(n5823), .B(n5822), .C(n5821), .D(n5824), .Y(n5825));
  OAI21X1 g4709(.A0(P2_D_REG_21__SCAN_IN), .A1(P2_D_REG_20__SCAN_IN), .B0(n5742), .Y(n5826));
  OAI21X1 g4710(.A0(P2_D_REG_19__SCAN_IN), .A1(P2_D_REG_18__SCAN_IN), .B0(n5742), .Y(n5827));
  OAI21X1 g4711(.A0(P2_D_REG_23__SCAN_IN), .A1(P2_D_REG_22__SCAN_IN), .B0(n5742), .Y(n5828));
  NAND3X1 g4712(.A(n5828), .B(n5827), .C(n5826), .Y(n5829));
  OAI21X1 g4713(.A0(P2_D_REG_14__SCAN_IN), .A1(P2_D_REG_12__SCAN_IN), .B0(n5742), .Y(n5830));
  OAI21X1 g4714(.A0(P2_D_REG_13__SCAN_IN), .A1(P2_D_REG_11__SCAN_IN), .B0(n5742), .Y(n5831));
  OAI21X1 g4715(.A0(P2_D_REG_24__SCAN_IN), .A1(P2_D_REG_16__SCAN_IN), .B0(n5742), .Y(n5832));
  OAI21X1 g4716(.A0(P2_D_REG_17__SCAN_IN), .A1(P2_D_REG_15__SCAN_IN), .B0(n5742), .Y(n5833));
  NAND4X1 g4717(.A(n5832), .B(n5831), .C(n5830), .D(n5833), .Y(n5834));
  NOR4X1  g4718(.A(n5829), .B(n5825), .C(n5820), .D(n5834), .Y(n5835));
  INVX1   g4719(.A(n5835), .Y(n5836));
  NOR2X1  g4720(.A(n5746), .B(n5750), .Y(n5837));
  AOI21X1 g4721(.A0(n5751), .A1(n5746), .B0(n5837), .Y(n5838));
  INVX1   g4722(.A(n5838), .Y(n5839));
  NAND2X1 g4723(.A(n5738), .B(n5732), .Y(n5840));
  NAND2X1 g4724(.A(n5840), .B(n5746), .Y(n5841));
  OAI21X1 g4725(.A0(n5746), .A1(n5726), .B0(n5841), .Y(n5842));
  NOR2X1  g4726(.A(P2_IR_REG_31__SCAN_IN), .B(n5636), .Y(n5843));
  AOI21X1 g4727(.A0(n5637), .A1(P2_IR_REG_31__SCAN_IN), .B0(n5843), .Y(n5844));
  NOR3X1  g4728(.A(n5653), .B(n5644), .C(n5473), .Y(n5845));
  AOI21X1 g4729(.A0(n5473), .A1(P2_IR_REG_22__SCAN_IN), .B0(n5845), .Y(n5846));
  INVX1   g4730(.A(n5844), .Y(n5847));
  NAND2X1 g4731(.A(n5473), .B(P2_IR_REG_20__SCAN_IN), .Y(n5848));
  OAI21X1 g4732(.A0(n5629), .A1(n5473), .B0(n5848), .Y(n5849));
  NOR2X1  g4733(.A(n5849), .B(n5847), .Y(n5850));
  XOR2X1  g4734(.A(n5850), .B(n5846), .Y(n5851));
  NOR2X1  g4735(.A(P2_IR_REG_31__SCAN_IN), .B(n5617), .Y(n5852));
  AOI21X1 g4736(.A0(n5618), .A1(P2_IR_REG_31__SCAN_IN), .B0(n5852), .Y(n5853));
  AOI21X1 g4737(.A0(n5853), .A1(n5844), .B0(n5851), .Y(n5854));
  NOR4X1  g4738(.A(n5842), .B(n5839), .C(n5836), .D(n5854), .Y(n5855));
  INVX1   g4739(.A(n5855), .Y(n5856));
  INVX1   g4740(.A(n5849), .Y(n5857));
  NOR3X1  g4741(.A(n5853), .B(n5847), .C(n5846), .Y(n5858));
  INVX1   g4742(.A(n5858), .Y(n5859));
  INVX1   g4743(.A(n5853), .Y(n5860));
  NOR4X1  g4744(.A(n5849), .B(n5844), .C(n5846), .D(n5860), .Y(n5861));
  INVX1   g4745(.A(n5861), .Y(n5862));
  OAI21X1 g4746(.A0(n5859), .A1(n5857), .B0(n5862), .Y(n5863));
  NAND4X1 g4747(.A(n5842), .B(n5839), .C(n5835), .D(n5863), .Y(n5864));
  AOI21X1 g4748(.A0(n5864), .A1(n5856), .B0(n5815), .Y(n5865));
  NAND2X1 g4749(.A(n5473), .B(P2_IR_REG_27__SCAN_IN), .Y(n5866));
  OAI21X1 g4750(.A0(n5689), .A1(n5473), .B0(n5866), .Y(n5867));
  NOR4X1  g4751(.A(n5699), .B(n5697), .C(n5473), .D(n5700), .Y(n5868));
  NOR2X1  g4752(.A(P2_IR_REG_31__SCAN_IN), .B(n5696), .Y(n5869));
  NOR3X1  g4753(.A(n5869), .B(n5868), .C(n5867), .Y(n5870));
  NAND2X1 g4754(.A(P2_IR_REG_31__SCAN_IN), .B(P2_IR_REG_0__SCAN_IN), .Y(n5871));
  INVX1   g4755(.A(n5871), .Y(n5872));
  INVX1   g4756(.A(P2_IR_REG_0__SCAN_IN), .Y(n5873));
  NOR2X1  g4757(.A(P2_IR_REG_31__SCAN_IN), .B(n5873), .Y(n5874));
  INVX1   g4758(.A(n5873), .Y(n5876));
  NAND2X1 g4759(.A(n5876), .B(n5870), .Y(n5877));
  OAI21X1 g4760(.A0(n5870), .A1(n5466), .B0(n5877), .Y(n5878));
  INVX1   g4761(.A(n5878), .Y(n5879));
  INVX1   g4762(.A(P2_IR_REG_30__SCAN_IN), .Y(n5880));
  NOR2X1  g4763(.A(P2_IR_REG_31__SCAN_IN), .B(n5880), .Y(n5881));
  AOI21X1 g4764(.A0(n5716), .A1(P2_IR_REG_31__SCAN_IN), .B0(n5881), .Y(n5882));
  NOR2X1  g4765(.A(P2_IR_REG_31__SCAN_IN), .B(n5707), .Y(n5883));
  AOI21X1 g4766(.A0(n5708), .A1(P2_IR_REG_31__SCAN_IN), .B0(n5883), .Y(n5884));
  NAND3X1 g4767(.A(n5884), .B(n5882), .C(P2_REG0_REG_0__SCAN_IN), .Y(n5885));
  XOR2X1  g4768(.A(n5715), .B(n5880), .Y(n5886));
  INVX1   g4769(.A(n5881), .Y(n5887));
  OAI21X1 g4770(.A0(n5886), .A1(n5473), .B0(n5887), .Y(n5888));
  NAND3X1 g4771(.A(n5884), .B(n5888), .C(P2_REG2_REG_0__SCAN_IN), .Y(n5889));
  NAND2X1 g4772(.A(n5708), .B(P2_IR_REG_31__SCAN_IN), .Y(n5890));
  OAI21X1 g4773(.A0(P2_IR_REG_31__SCAN_IN), .A1(n5707), .B0(n5890), .Y(n5891));
  NAND3X1 g4774(.A(n5891), .B(n5882), .C(P2_REG1_REG_0__SCAN_IN), .Y(n5892));
  NAND3X1 g4775(.A(n5891), .B(n5888), .C(P2_REG3_REG_0__SCAN_IN), .Y(n5893));
  NAND4X1 g4776(.A(n5892), .B(n5889), .C(n5885), .D(n5893), .Y(n5894));
  XOR2X1  g4777(.A(n5894), .B(n5879), .Y(n5895));
  NOR3X1  g4778(.A(n5853), .B(n5849), .C(n5846), .Y(n5896));
  INVX1   g4779(.A(n5896), .Y(n5897));
  NOR2X1  g4780(.A(n5897), .B(n5895), .Y(n5898));
  INVX1   g4781(.A(n5898), .Y(n5899));
  NOR3X1  g4782(.A(n5853), .B(n5857), .C(n5844), .Y(n5901));
  NOR3X1  g4783(.A(n5860), .B(n5857), .C(n5846), .Y(n5902));
  OAI21X1 g4784(.A0(n5902), .A1(n5901), .B0(n8531), .Y(n5903));
  NOR3X1  g4785(.A(n5853), .B(n5857), .C(n5846), .Y(n5904));
  NOR3X1  g4786(.A(n5860), .B(n5857), .C(n5844), .Y(n5905));
  OAI21X1 g4787(.A0(n5905), .A1(n5904), .B0(n8531), .Y(n5906));
  INVX1   g4788(.A(n5846), .Y(n5907));
  NOR4X1  g4789(.A(n5849), .B(n5844), .C(n5907), .D(n5860), .Y(n5908));
  NOR4X1  g4790(.A(n5849), .B(n5847), .C(n5846), .D(n5860), .Y(n5909));
  OAI21X1 g4791(.A0(n5909), .A1(n5908), .B0(n8531), .Y(n5910));
  NAND4X1 g4792(.A(n5906), .B(n5903), .C(n5899), .D(n5910), .Y(n5911));
  INVX1   g4793(.A(n5911), .Y(n5912));
  NOR3X1  g4794(.A(n5853), .B(n5849), .C(n5907), .Y(n5913));
  INVX1   g4795(.A(n5867), .Y(n5914));
  NOR2X1  g4796(.A(n5869), .B(n5868), .Y(n5915));
  XOR2X1  g4797(.A(n5915), .B(n5914), .Y(n5916));
  NOR3X1  g4798(.A(n5916), .B(n5844), .C(n5846), .Y(n5917));
  INVX1   g4799(.A(n5917), .Y(n5918));
  NAND3X1 g4800(.A(n5884), .B(n5882), .C(P2_REG0_REG_1__SCAN_IN), .Y(n5919));
  NAND3X1 g4801(.A(n5884), .B(n5888), .C(P2_REG2_REG_1__SCAN_IN), .Y(n5920));
  NAND2X1 g4802(.A(n5920), .B(n5919), .Y(n5921));
  NAND3X1 g4803(.A(n5891), .B(n5882), .C(P2_REG1_REG_1__SCAN_IN), .Y(n5922));
  NAND3X1 g4804(.A(n5891), .B(n5888), .C(P2_REG3_REG_1__SCAN_IN), .Y(n5923));
  NAND2X1 g4805(.A(n5923), .B(n5922), .Y(n5924));
  NOR2X1  g4806(.A(n5924), .B(n5921), .Y(n5925));
  NAND2X1 g4807(.A(n5844), .B(n5846), .Y(n5926));
  OAI22X1 g4808(.A0(n5925), .A1(n5918), .B0(n5879), .B1(n5926), .Y(n5927));
  AOI21X1 g4809(.A0(n5913), .A1(n8531), .B0(n5927), .Y(n5928));
  NAND2X1 g4810(.A(n5928), .B(n5912), .Y(n5929));
  NAND2X1 g4811(.A(n5929), .B(n5865), .Y(n5930));
  OAI21X1 g4812(.A0(n5865), .A1(n5814), .B0(n5930), .Y(P2_U3390));
  NOR2X1  g4813(.A(n5894), .B(n5879), .Y(n5932));
  NAND4X1 g4814(.A(n5922), .B(n5920), .C(n5919), .D(n5923), .Y(n5933));
  INVX1   g4815(.A(P2_IR_REG_1__SCAN_IN), .Y(n5934));
  NOR2X1  g4816(.A(P2_IR_REG_31__SCAN_IN), .B(n5934), .Y(n5935));
  AOI21X1 g4817(.A0(n5475), .A1(P2_IR_REG_31__SCAN_IN), .B0(n5935), .Y(n5936));
  INVX1   g4818(.A(n5936), .Y(n5937));
  NOR2X1  g4819(.A(n5870), .B(n5470), .Y(n5938));
  AOI21X1 g4820(.A0(n5937), .A1(n5870), .B0(n5938), .Y(n5939));
  XOR2X1  g4821(.A(n5939), .B(n5933), .Y(n5940));
  XOR2X1  g4822(.A(n5940), .B(n5932), .Y(n5941));
  INVX1   g4823(.A(n5941), .Y(n5942));
  OAI21X1 g4824(.A0(n5909), .A1(n5902), .B0(n5942), .Y(n5943));
  NAND2X1 g4825(.A(n5937), .B(n5870), .Y(n5944));
  OAI21X1 g4826(.A0(n5870), .A1(n5470), .B0(n5944), .Y(n5945));
  XOR2X1  g4827(.A(n5945), .B(n5933), .Y(n5946));
  NAND2X1 g4828(.A(n5894), .B(n5878), .Y(n5947));
  XOR2X1  g4829(.A(n5947), .B(n5946), .Y(n5948));
  INVX1   g4830(.A(n5948), .Y(n5949));
  AOI22X1 g4831(.A0(n5942), .A1(n5908), .B0(n5901), .B1(n5949), .Y(n5950));
  XOR2X1  g4832(.A(n5915), .B(n5867), .Y(n5951));
  NOR3X1  g4833(.A(n5951), .B(n5844), .C(n5846), .Y(n5952));
  AOI22X1 g4834(.A0(n5949), .A1(n5905), .B0(n5894), .B1(n5952), .Y(n5953));
  OAI21X1 g4835(.A0(n5904), .A1(n5896), .B0(n5949), .Y(n5954));
  NAND4X1 g4836(.A(n5953), .B(n5950), .C(n5943), .D(n5954), .Y(n5955));
  INVX1   g4837(.A(n5955), .Y(n5956));
  NOR2X1  g4838(.A(n5891), .B(n5888), .Y(n5957));
  NOR2X1  g4839(.A(n5891), .B(n5882), .Y(n5958));
  AOI22X1 g4840(.A0(n5957), .A1(P2_REG0_REG_2__SCAN_IN), .B0(P2_REG2_REG_2__SCAN_IN), .B1(n5958), .Y(n5959));
  INVX1   g4841(.A(n5959), .Y(n5960));
  NOR2X1  g4842(.A(n5884), .B(n5888), .Y(n5961));
  NOR2X1  g4843(.A(n5884), .B(n5882), .Y(n5962));
  AOI22X1 g4844(.A0(n5961), .A1(P2_REG1_REG_2__SCAN_IN), .B0(P2_REG3_REG_2__SCAN_IN), .B1(n5962), .Y(n5963));
  INVX1   g4845(.A(n5963), .Y(n5964));
  NOR2X1  g4846(.A(n5964), .B(n5960), .Y(n5965));
  OAI22X1 g4847(.A0(n5939), .A1(n5926), .B0(n5918), .B1(n5965), .Y(n5966));
  AOI21X1 g4848(.A0(n5942), .A1(n5913), .B0(n5966), .Y(n5967));
  NAND2X1 g4849(.A(n5967), .B(n5956), .Y(n5968));
  NAND2X1 g4850(.A(n5968), .B(n5865), .Y(n5969));
  INVX1   g4851(.A(n5865), .Y(n5970));
  NAND2X1 g4852(.A(n5970), .B(P2_REG0_REG_1__SCAN_IN), .Y(n5971));
  NAND2X1 g4853(.A(n5971), .B(n5969), .Y(P2_U3393));
  NOR2X1  g4854(.A(n5939), .B(n5925), .Y(n5973));
  NOR2X1  g4855(.A(n5945), .B(n5933), .Y(n5974));
  NOR2X1  g4856(.A(n5947), .B(n5974), .Y(n5975));
  NOR2X1  g4857(.A(n5975), .B(n5973), .Y(n5976));
  NOR2X1  g4858(.A(P2_IR_REG_31__SCAN_IN), .B(n5480), .Y(n5977));
  AOI21X1 g4859(.A0(n5482), .A1(P2_IR_REG_31__SCAN_IN), .B0(n5977), .Y(n5978));
  INVX1   g4860(.A(n5978), .Y(n5979));
  NOR2X1  g4861(.A(n5870), .B(n5479), .Y(n5980));
  AOI21X1 g4862(.A0(n5979), .A1(n5870), .B0(n5980), .Y(n5981));
  AOI21X1 g4863(.A0(n5963), .A1(n5959), .B0(n5981), .Y(n5982));
  NAND2X1 g4864(.A(n5979), .B(n5870), .Y(n5983));
  OAI21X1 g4865(.A0(n5870), .A1(n5479), .B0(n5983), .Y(n5984));
  NOR3X1  g4866(.A(n5984), .B(n5964), .C(n5960), .Y(n5985));
  NOR3X1  g4867(.A(n5976), .B(n5985), .C(n5982), .Y(n5986));
  XOR2X1  g4868(.A(n5984), .B(n5965), .Y(n5987));
  AOI21X1 g4869(.A0(n5987), .A1(n5976), .B0(n5986), .Y(n5988));
  NAND2X1 g4870(.A(n5988), .B(n5901), .Y(n5989));
  OAI21X1 g4871(.A0(n5904), .A1(n5896), .B0(n5988), .Y(n5990));
  INVX1   g4872(.A(n5902), .Y(n5991));
  NAND2X1 g4873(.A(n5889), .B(n5885), .Y(n5992));
  NAND2X1 g4874(.A(n5893), .B(n5892), .Y(n5993));
  NOR2X1  g4875(.A(n5993), .B(n5992), .Y(n5994));
  NAND2X1 g4876(.A(n5994), .B(n5878), .Y(n5995));
  OAI21X1 g4877(.A0(n5933), .A1(n5995), .B0(n5939), .Y(n5996));
  OAI21X1 g4878(.A0(n5925), .A1(n5932), .B0(n5996), .Y(n5997));
  INVX1   g4879(.A(n5997), .Y(n5998));
  XOR2X1  g4880(.A(n5998), .B(n5987), .Y(n5999));
  AOI22X1 g4881(.A0(n5952), .A1(n5933), .B0(n5905), .B1(n5988), .Y(n6000));
  OAI21X1 g4882(.A0(n5999), .A1(n5991), .B0(n6000), .Y(n6001));
  INVX1   g4883(.A(n5908), .Y(n6002));
  INVX1   g4884(.A(n5909), .Y(n6003));
  AOI21X1 g4885(.A0(n6003), .A1(n6002), .B0(n5999), .Y(n6004));
  NOR2X1  g4886(.A(n6004), .B(n6001), .Y(n6005));
  NAND3X1 g4887(.A(n6005), .B(n5990), .C(n5989), .Y(n6006));
  INVX1   g4888(.A(n5913), .Y(n6007));
  INVX1   g4889(.A(n5926), .Y(n6008));
  AOI22X1 g4890(.A0(n5957), .A1(P2_REG0_REG_3__SCAN_IN), .B0(P2_REG2_REG_3__SCAN_IN), .B1(n5958), .Y(n6009));
  INVX1   g4891(.A(P2_REG3_REG_3__SCAN_IN), .Y(n6010));
  AOI22X1 g4892(.A0(n5961), .A1(P2_REG1_REG_3__SCAN_IN), .B0(n6010), .B1(n5962), .Y(n6011));
  NAND2X1 g4893(.A(n6011), .B(n6009), .Y(n6012));
  AOI22X1 g4894(.A0(n5984), .A1(n6008), .B0(n5917), .B1(n6012), .Y(n6013));
  OAI21X1 g4895(.A0(n5999), .A1(n6007), .B0(n6013), .Y(n6014));
  NOR2X1  g4896(.A(n6014), .B(n6006), .Y(n6015));
  NAND2X1 g4897(.A(n5970), .B(P2_REG0_REG_2__SCAN_IN), .Y(n6016));
  OAI21X1 g4898(.A0(n6015), .A1(n5970), .B0(n6016), .Y(P2_U3396));
  INVX1   g4899(.A(n5901), .Y(n6018));
  NOR2X1  g4900(.A(P2_IR_REG_31__SCAN_IN), .B(n5487), .Y(n6019));
  AOI21X1 g4901(.A0(n5489), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6019), .Y(n6020));
  INVX1   g4902(.A(n6020), .Y(n6021));
  NAND2X1 g4903(.A(n6021), .B(n5870), .Y(n6022));
  OAI21X1 g4904(.A0(n5870), .A1(n5486), .B0(n6022), .Y(n6023));
  INVX1   g4905(.A(n6023), .Y(n6024));
  XOR2X1  g4906(.A(n6024), .B(n6012), .Y(n6025));
  INVX1   g4907(.A(n5985), .Y(n6027));
  AOI21X1 g4908(.A0(n6027), .A1(n5973), .B0(n5982), .Y(n6028));
  INVX1   g4909(.A(n6028), .Y(n6029));
  AOI21X1 g4910(.A0(n5975), .A1(n6027), .B0(n6029), .Y(n6030));
  XOR2X1  g4911(.A(n6023), .B(n6012), .Y(n6031));
  NOR2X1  g4912(.A(n6031), .B(n6030), .Y(n6032));
  AOI21X1 g4913(.A0(n6030), .A1(n6031), .B0(n6032), .Y(n6033));
  NOR2X1  g4914(.A(n6033), .B(n6018), .Y(n6034));
  INVX1   g4915(.A(n5904), .Y(n6035));
  AOI21X1 g4916(.A0(n6035), .A1(n5897), .B0(n6033), .Y(n6036));
  NOR2X1  g4917(.A(n6036), .B(n6034), .Y(n6037));
  AOI21X1 g4918(.A0(n5963), .A1(n5959), .B0(n5984), .Y(n6038));
  NOR3X1  g4919(.A(n5981), .B(n5964), .C(n5960), .Y(n6039));
  NOR2X1  g4920(.A(n6025), .B(n6039), .Y(n6040));
  OAI21X1 g4921(.A0(n5997), .A1(n6038), .B0(n6040), .Y(n6041));
  NOR2X1  g4922(.A(n6031), .B(n6038), .Y(n6042));
  OAI21X1 g4923(.A0(n5998), .A1(n6039), .B0(n6042), .Y(n6043));
  NAND2X1 g4924(.A(n6043), .B(n6041), .Y(n6044));
  INVX1   g4925(.A(n5905), .Y(n6045));
  INVX1   g4926(.A(n5952), .Y(n6046));
  OAI22X1 g4927(.A0(n5965), .A1(n6046), .B0(n6045), .B1(n6033), .Y(n6047));
  AOI21X1 g4928(.A0(n6044), .A1(n5902), .B0(n6047), .Y(n6048));
  OAI21X1 g4929(.A0(n5909), .A1(n5908), .B0(n6044), .Y(n6049));
  NAND3X1 g4930(.A(n6049), .B(n6048), .C(n6037), .Y(n6050));
  INVX1   g4931(.A(n6044), .Y(n6051));
  AOI22X1 g4932(.A0(n5957), .A1(P2_REG0_REG_4__SCAN_IN), .B0(P2_REG2_REG_4__SCAN_IN), .B1(n5958), .Y(n6052));
  XOR2X1  g4933(.A(P2_REG3_REG_4__SCAN_IN), .B(P2_REG3_REG_3__SCAN_IN), .Y(n6053));
  INVX1   g4934(.A(n6053), .Y(n6054));
  AOI22X1 g4935(.A0(n5962), .A1(n6054), .B0(n5961), .B1(P2_REG1_REG_4__SCAN_IN), .Y(n6055));
  NAND2X1 g4936(.A(n6055), .B(n6052), .Y(n6056));
  AOI22X1 g4937(.A0(n6023), .A1(n6008), .B0(n5917), .B1(n6056), .Y(n6057));
  OAI21X1 g4938(.A0(n6051), .A1(n6007), .B0(n6057), .Y(n6058));
  NOR2X1  g4939(.A(n6058), .B(n6050), .Y(n6059));
  NAND2X1 g4940(.A(n5970), .B(P2_REG0_REG_3__SCAN_IN), .Y(n6060));
  OAI21X1 g4941(.A0(n6059), .A1(n5970), .B0(n6060), .Y(P2_U3399));
  AOI21X1 g4942(.A0(n6011), .A1(n6009), .B0(n6024), .Y(n6062));
  NOR2X1  g4943(.A(P2_IR_REG_31__SCAN_IN), .B(n5494), .Y(n6063));
  AOI21X1 g4944(.A0(n5496), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6063), .Y(n6064));
  INVX1   g4945(.A(n6064), .Y(n6065));
  NAND2X1 g4946(.A(n6065), .B(n5870), .Y(n6066));
  OAI21X1 g4947(.A0(n5870), .A1(n5493), .B0(n6066), .Y(n6067));
  INVX1   g4948(.A(n6067), .Y(n6068));
  XOR2X1  g4949(.A(n6068), .B(n6056), .Y(n6069));
  NOR2X1  g4950(.A(n6023), .B(n6012), .Y(n6070));
  NOR2X1  g4951(.A(n6070), .B(n6028), .Y(n6071));
  NOR4X1  g4952(.A(n5985), .B(n5947), .C(n5974), .D(n6070), .Y(n6072));
  NOR4X1  g4953(.A(n6071), .B(n6069), .C(n6062), .D(n6072), .Y(n6073));
  NOR3X1  g4954(.A(n6072), .B(n6071), .C(n6062), .Y(n6074));
  XOR2X1  g4955(.A(n6067), .B(n6056), .Y(n6075));
  NOR2X1  g4956(.A(n6075), .B(n6074), .Y(n6076));
  OAI21X1 g4957(.A0(n6076), .A1(n6073), .B0(n5901), .Y(n6077));
  OAI22X1 g4958(.A0(n6073), .A1(n6076), .B0(n5904), .B1(n5896), .Y(n6078));
  INVX1   g4959(.A(n6012), .Y(n6079));
  AOI21X1 g4960(.A0(n6023), .A1(n6079), .B0(n6039), .Y(n6080));
  NAND2X1 g4961(.A(n6012), .B(n6038), .Y(n6081));
  OAI21X1 g4962(.A0(n6012), .A1(n6038), .B0(n6024), .Y(n6082));
  NAND2X1 g4963(.A(n6082), .B(n6081), .Y(n6083));
  AOI21X1 g4964(.A0(n6080), .A1(n5997), .B0(n6083), .Y(n6084));
  XOR2X1  g4965(.A(n6084), .B(n6069), .Y(n6085));
  INVX1   g4966(.A(n6085), .Y(n6086));
  NOR2X1  g4967(.A(n6076), .B(n6073), .Y(n6087));
  OAI22X1 g4968(.A0(n6079), .A1(n6046), .B0(n6045), .B1(n6087), .Y(n6088));
  AOI21X1 g4969(.A0(n6086), .A1(n5902), .B0(n6088), .Y(n6089));
  OAI21X1 g4970(.A0(n5909), .A1(n5908), .B0(n6086), .Y(n6090));
  NAND4X1 g4971(.A(n6089), .B(n6078), .C(n6077), .D(n6090), .Y(n6091));
  AOI22X1 g4972(.A0(n5957), .A1(P2_REG0_REG_5__SCAN_IN), .B0(P2_REG2_REG_5__SCAN_IN), .B1(n5958), .Y(n6092));
  INVX1   g4973(.A(P2_REG3_REG_5__SCAN_IN), .Y(n6093));
  NOR2X1  g4974(.A(P2_REG3_REG_4__SCAN_IN), .B(P2_REG3_REG_3__SCAN_IN), .Y(n6094));
  XOR2X1  g4975(.A(n6094), .B(n6093), .Y(n6095));
  INVX1   g4976(.A(n6095), .Y(n6096));
  AOI22X1 g4977(.A0(n5962), .A1(n6096), .B0(n5961), .B1(P2_REG1_REG_5__SCAN_IN), .Y(n6097));
  NAND2X1 g4978(.A(n6097), .B(n6092), .Y(n6098));
  AOI22X1 g4979(.A0(n6067), .A1(n6008), .B0(n5917), .B1(n6098), .Y(n6099));
  OAI21X1 g4980(.A0(n6085), .A1(n6007), .B0(n6099), .Y(n6100));
  NOR2X1  g4981(.A(n6100), .B(n6091), .Y(n6101));
  NAND2X1 g4982(.A(n5970), .B(P2_REG0_REG_4__SCAN_IN), .Y(n6102));
  OAI21X1 g4983(.A0(n6101), .A1(n5970), .B0(n6102), .Y(P2_U3402));
  INVX1   g4984(.A(n6056), .Y(n6104));
  AOI21X1 g4985(.A0(n6055), .A1(n6052), .B0(n6068), .Y(n6105));
  NOR4X1  g4986(.A(n6072), .B(n6071), .C(n6062), .D(n6105), .Y(n6106));
  INVX1   g4987(.A(P2_REG2_REG_5__SCAN_IN), .Y(n6107));
  NAND2X1 g4988(.A(n5884), .B(n5888), .Y(n6108));
  NAND3X1 g4989(.A(n5884), .B(n5882), .C(P2_REG0_REG_5__SCAN_IN), .Y(n6109));
  OAI21X1 g4990(.A0(n6108), .A1(n6107), .B0(n6109), .Y(n6110));
  INVX1   g4991(.A(P2_REG1_REG_5__SCAN_IN), .Y(n6111));
  NAND2X1 g4992(.A(n5891), .B(n5882), .Y(n6112));
  NAND2X1 g4993(.A(n5891), .B(n5888), .Y(n6113));
  OAI22X1 g4994(.A0(n6113), .A1(n6095), .B0(n6112), .B1(n6111), .Y(n6114));
  NOR2X1  g4995(.A(n6114), .B(n6110), .Y(n6115));
  NOR2X1  g4996(.A(P2_IR_REG_31__SCAN_IN), .B(n5507), .Y(n6116));
  AOI21X1 g4997(.A0(n5502), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6116), .Y(n6117));
  NOR4X1  g4998(.A(n5869), .B(n5868), .C(n5867), .D(n6117), .Y(n6118));
  NOR2X1  g4999(.A(n5870), .B(n5500), .Y(n6119));
  NOR2X1  g5000(.A(n6119), .B(n6118), .Y(n6120));
  NOR2X1  g5001(.A(n6067), .B(n6056), .Y(n6121));
  INVX1   g5002(.A(n6118), .Y(n6122));
  OAI21X1 g5003(.A0(n5870), .A1(n5500), .B0(n6122), .Y(n6123));
  NOR2X1  g5004(.A(n6123), .B(n6098), .Y(n6124));
  NOR2X1  g5005(.A(n6124), .B(n6121), .Y(n6125));
  OAI21X1 g5006(.A0(n6120), .A1(n6115), .B0(n6125), .Y(n6126));
  NOR2X1  g5007(.A(n6121), .B(n6074), .Y(n6127));
  XOR2X1  g5008(.A(n6123), .B(n6115), .Y(n6128));
  OAI21X1 g5009(.A0(n6068), .A1(n6104), .B0(n6128), .Y(n6129));
  OAI22X1 g5010(.A0(n6127), .A1(n6129), .B0(n6126), .B1(n6106), .Y(n6130));
  OAI22X1 g5011(.A0(n6104), .A1(n6046), .B0(n6045), .B1(n6130), .Y(n6131));
  NOR2X1  g5012(.A(n6130), .B(n6018), .Y(n6132));
  AOI21X1 g5013(.A0(n6035), .A1(n5897), .B0(n6130), .Y(n6133));
  NOR2X1  g5014(.A(n6068), .B(n6056), .Y(n6134));
  NOR2X1  g5015(.A(n6084), .B(n6134), .Y(n6135));
  AOI21X1 g5016(.A0(n6068), .A1(n6056), .B0(n6135), .Y(n6136));
  XOR2X1  g5017(.A(n6136), .B(n6128), .Y(n6137));
  INVX1   g5018(.A(n6137), .Y(n6138));
  OAI21X1 g5019(.A0(n5908), .A1(n5902), .B0(n6138), .Y(n6139));
  OAI21X1 g5020(.A0(n6137), .A1(n6003), .B0(n6139), .Y(n6140));
  NOR4X1  g5021(.A(n6133), .B(n6132), .C(n6131), .D(n6140), .Y(n6141));
  INVX1   g5022(.A(n6141), .Y(n6142));
  AOI22X1 g5023(.A0(n5957), .A1(P2_REG0_REG_6__SCAN_IN), .B0(P2_REG2_REG_6__SCAN_IN), .B1(n5958), .Y(n6143));
  NOR4X1  g5024(.A(P2_REG3_REG_4__SCAN_IN), .B(P2_REG3_REG_5__SCAN_IN), .C(P2_REG3_REG_3__SCAN_IN), .D(P2_REG3_REG_6__SCAN_IN), .Y(n6144));
  INVX1   g5025(.A(P2_REG3_REG_6__SCAN_IN), .Y(n6145));
  AOI21X1 g5026(.A0(n6094), .A1(n6093), .B0(n6145), .Y(n6146));
  NOR2X1  g5027(.A(n6146), .B(n6144), .Y(n6147));
  INVX1   g5028(.A(n6147), .Y(n6148));
  AOI22X1 g5029(.A0(n5962), .A1(n6148), .B0(n5961), .B1(P2_REG1_REG_6__SCAN_IN), .Y(n6149));
  NAND2X1 g5030(.A(n6149), .B(n6143), .Y(n6150));
  AOI22X1 g5031(.A0(n6123), .A1(n6008), .B0(n5917), .B1(n6150), .Y(n6151));
  OAI21X1 g5032(.A0(n6137), .A1(n6007), .B0(n6151), .Y(n6152));
  NOR2X1  g5033(.A(n6152), .B(n6142), .Y(n6153));
  NAND2X1 g5034(.A(n5970), .B(P2_REG0_REG_5__SCAN_IN), .Y(n6154));
  OAI21X1 g5035(.A0(n6153), .A1(n5970), .B0(n6154), .Y(P2_U3405));
  INVX1   g5036(.A(n6150), .Y(n6156));
  NOR2X1  g5037(.A(P2_IR_REG_31__SCAN_IN), .B(n5509), .Y(n6157));
  AOI21X1 g5038(.A0(n5512), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6157), .Y(n6158));
  INVX1   g5039(.A(n6158), .Y(n6159));
  NAND2X1 g5040(.A(n6159), .B(n5870), .Y(n6160));
  OAI21X1 g5041(.A0(n5870), .A1(n5506), .B0(n6160), .Y(n6161));
  XOR2X1  g5042(.A(n6161), .B(n6156), .Y(n6162));
  AOI21X1 g5043(.A0(n6023), .A1(n6012), .B0(n5982), .Y(n6163));
  OAI21X1 g5044(.A0(n5976), .A1(n5985), .B0(n6163), .Y(n6164));
  NOR3X1  g5045(.A(n6124), .B(n6121), .C(n6070), .Y(n6165));
  NAND3X1 g5046(.A(n6123), .B(n6067), .C(n6056), .Y(n6166));
  AOI21X1 g5047(.A0(n6067), .A1(n6056), .B0(n6123), .Y(n6167));
  OAI21X1 g5048(.A0(n6167), .A1(n6115), .B0(n6166), .Y(n6168));
  AOI21X1 g5049(.A0(n6165), .A1(n6164), .B0(n6168), .Y(n6169));
  INVX1   g5050(.A(n6169), .Y(n6170));
  NOR2X1  g5051(.A(n6170), .B(n6162), .Y(n6171));
  XOR2X1  g5052(.A(n6161), .B(n6150), .Y(n6172));
  NOR2X1  g5053(.A(n6172), .B(n6169), .Y(n6173));
  NOR2X1  g5054(.A(n6173), .B(n6171), .Y(n6174));
  OAI22X1 g5055(.A0(n6115), .A1(n6046), .B0(n6045), .B1(n6174), .Y(n6175));
  OAI22X1 g5056(.A0(n6171), .A1(n6173), .B0(n5904), .B1(n5896), .Y(n6176));
  OAI21X1 g5057(.A0(n6174), .A1(n6018), .B0(n6176), .Y(n6177));
  INVX1   g5058(.A(n6136), .Y(n6178));
  AOI21X1 g5059(.A0(n6120), .A1(n6098), .B0(n6178), .Y(n6179));
  NAND2X1 g5060(.A(n6123), .B(n6115), .Y(n6180));
  INVX1   g5061(.A(n6180), .Y(n6181));
  NOR2X1  g5062(.A(n6162), .B(n6181), .Y(n6182));
  INVX1   g5063(.A(n6182), .Y(n6183));
  NOR2X1  g5064(.A(n5870), .B(n5506), .Y(n6184));
  AOI21X1 g5065(.A0(n6159), .A1(n5870), .B0(n6184), .Y(n6185));
  NOR2X1  g5066(.A(n6185), .B(n6150), .Y(n6186));
  AOI22X1 g5067(.A0(n6150), .A1(n6185), .B0(n6120), .B1(n6098), .Y(n6187));
  INVX1   g5068(.A(n6187), .Y(n6188));
  NOR2X1  g5069(.A(n6188), .B(n6186), .Y(n6189));
  OAI21X1 g5070(.A0(n6136), .A1(n6181), .B0(n6189), .Y(n6190));
  OAI21X1 g5071(.A0(n6183), .A1(n6179), .B0(n6190), .Y(n6191));
  INVX1   g5072(.A(n6191), .Y(n6192));
  OAI21X1 g5073(.A0(n5908), .A1(n5902), .B0(n6191), .Y(n6193));
  OAI21X1 g5074(.A0(n6192), .A1(n6003), .B0(n6193), .Y(n6194));
  AOI22X1 g5075(.A0(n5957), .A1(P2_REG0_REG_7__SCAN_IN), .B0(P2_REG2_REG_7__SCAN_IN), .B1(n5958), .Y(n6195));
  INVX1   g5076(.A(P2_REG3_REG_7__SCAN_IN), .Y(n6196));
  XOR2X1  g5077(.A(n6144), .B(n6196), .Y(n6197));
  INVX1   g5078(.A(n6197), .Y(n6198));
  AOI22X1 g5079(.A0(n5962), .A1(n6198), .B0(n5961), .B1(P2_REG1_REG_7__SCAN_IN), .Y(n6199));
  NAND2X1 g5080(.A(n6199), .B(n6195), .Y(n6200));
  AOI22X1 g5081(.A0(n6161), .A1(n6008), .B0(n5917), .B1(n6200), .Y(n6201));
  OAI21X1 g5082(.A0(n6192), .A1(n6007), .B0(n6201), .Y(n6202));
  NOR4X1  g5083(.A(n6194), .B(n6177), .C(n6175), .D(n6202), .Y(n6203));
  NAND2X1 g5084(.A(n5970), .B(P2_REG0_REG_6__SCAN_IN), .Y(n6204));
  OAI21X1 g5085(.A0(n6203), .A1(n5970), .B0(n6204), .Y(P2_U3408));
  INVX1   g5086(.A(n6200), .Y(n6206));
  NOR2X1  g5087(.A(P2_IR_REG_31__SCAN_IN), .B(n5517), .Y(n6207));
  AOI21X1 g5088(.A0(n5518), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6207), .Y(n6208));
  INVX1   g5089(.A(n6208), .Y(n6209));
  NAND2X1 g5090(.A(n6209), .B(n5870), .Y(n6210));
  OAI21X1 g5091(.A0(n5870), .A1(n5516), .B0(n6210), .Y(n6211));
  XOR2X1  g5092(.A(n6211), .B(n6206), .Y(n6212));
  INVX1   g5093(.A(n6084), .Y(n6213));
  NAND3X1 g5094(.A(n6180), .B(n6068), .C(n6056), .Y(n6214));
  AOI21X1 g5095(.A0(n6214), .A1(n6187), .B0(n6186), .Y(n6215));
  NOR3X1  g5096(.A(n6186), .B(n6181), .C(n6134), .Y(n6216));
  AOI21X1 g5097(.A0(n6216), .A1(n6213), .B0(n6215), .Y(n6217));
  XOR2X1  g5098(.A(n6217), .B(n6212), .Y(n6218));
  INVX1   g5099(.A(n6218), .Y(n6219));
  OAI21X1 g5100(.A0(n5909), .A1(n5902), .B0(n6219), .Y(n6220));
  NAND2X1 g5101(.A(n6161), .B(n6150), .Y(n6221));
  INVX1   g5102(.A(n6211), .Y(n6222));
  OAI22X1 g5103(.A0(n6200), .A1(n6211), .B0(n6161), .B1(n6150), .Y(n6223));
  INVX1   g5104(.A(n6223), .Y(n6224));
  OAI21X1 g5105(.A0(n6222), .A1(n6206), .B0(n6224), .Y(n6225));
  AOI21X1 g5106(.A0(n6221), .A1(n6169), .B0(n6225), .Y(n6226));
  INVX1   g5107(.A(n6221), .Y(n6227));
  AOI21X1 g5108(.A0(n6199), .A1(n6195), .B0(n6211), .Y(n6228));
  NOR2X1  g5109(.A(n6222), .B(n6200), .Y(n6229));
  AOI21X1 g5110(.A0(n6185), .A1(n6156), .B0(n6169), .Y(n6230));
  NOR4X1  g5111(.A(n6229), .B(n6228), .C(n6227), .D(n6230), .Y(n6231));
  NOR2X1  g5112(.A(n6231), .B(n6226), .Y(n6232));
  AOI22X1 g5113(.A0(n6219), .A1(n5908), .B0(n5901), .B1(n6232), .Y(n6233));
  AOI22X1 g5114(.A0(n6150), .A1(n5952), .B0(n5905), .B1(n6232), .Y(n6234));
  OAI21X1 g5115(.A0(n5904), .A1(n5896), .B0(n6232), .Y(n6235));
  NAND4X1 g5116(.A(n6234), .B(n6233), .C(n6220), .D(n6235), .Y(n6236));
  AOI22X1 g5117(.A0(n5957), .A1(P2_REG0_REG_8__SCAN_IN), .B0(P2_REG2_REG_8__SCAN_IN), .B1(n5958), .Y(n6237));
  NAND2X1 g5118(.A(n6144), .B(n6196), .Y(n6238));
  XOR2X1  g5119(.A(n6238), .B(P2_REG3_REG_8__SCAN_IN), .Y(n6239));
  INVX1   g5120(.A(n6239), .Y(n6240));
  AOI22X1 g5121(.A0(n5962), .A1(n6240), .B0(n5961), .B1(P2_REG1_REG_8__SCAN_IN), .Y(n6241));
  NAND2X1 g5122(.A(n6241), .B(n6237), .Y(n6242));
  AOI22X1 g5123(.A0(n6211), .A1(n6008), .B0(n5917), .B1(n6242), .Y(n6243));
  OAI21X1 g5124(.A0(n6218), .A1(n6007), .B0(n6243), .Y(n6244));
  NOR2X1  g5125(.A(n6244), .B(n6236), .Y(n6245));
  NAND2X1 g5126(.A(n5970), .B(P2_REG0_REG_7__SCAN_IN), .Y(n6246));
  OAI21X1 g5127(.A0(n6245), .A1(n5970), .B0(n6246), .Y(P2_U3411));
  INVX1   g5128(.A(n6217), .Y(n6248));
  INVX1   g5129(.A(n6242), .Y(n6249));
  NOR2X1  g5130(.A(P2_IR_REG_31__SCAN_IN), .B(n5524), .Y(n6250));
  AOI21X1 g5131(.A0(n5529), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6250), .Y(n6251));
  INVX1   g5132(.A(n6251), .Y(n6252));
  NAND2X1 g5133(.A(n6252), .B(n5870), .Y(n6253));
  OAI21X1 g5134(.A0(n5870), .A1(n5523), .B0(n6253), .Y(n6254));
  XOR2X1  g5135(.A(n6254), .B(n6249), .Y(n6255));
  NOR2X1  g5136(.A(n6255), .B(n6229), .Y(n6256));
  OAI21X1 g5137(.A0(n6248), .A1(n6228), .B0(n6256), .Y(n6257));
  NOR2X1  g5138(.A(n6268), .B(n6228), .Y(n6259));
  OAI21X1 g5139(.A0(n6217), .A1(n6229), .B0(n6259), .Y(n6260));
  NAND2X1 g5140(.A(n6260), .B(n6257), .Y(n6261));
  OAI21X1 g5141(.A0(n5909), .A1(n5902), .B0(n6261), .Y(n6262));
  AOI21X1 g5142(.A0(n6222), .A1(n6221), .B0(n6206), .Y(n6263));
  AOI21X1 g5143(.A0(n6211), .A1(n6227), .B0(n6263), .Y(n6264));
  OAI21X1 g5144(.A0(n6223), .A1(n6169), .B0(n6264), .Y(n6265));
  NOR2X1  g5145(.A(n6265), .B(n6255), .Y(n6266));
  INVX1   g5146(.A(n6265), .Y(n6267));
  XOR2X1  g5147(.A(n6254), .B(n6242), .Y(n6268));
  NOR2X1  g5148(.A(n6268), .B(n6267), .Y(n6269));
  NOR2X1  g5149(.A(n6269), .B(n6266), .Y(n6270));
  NOR2X1  g5150(.A(n6270), .B(n6018), .Y(n6271));
  AOI21X1 g5151(.A0(n6261), .A1(n5908), .B0(n6271), .Y(n6272));
  NAND2X1 g5152(.A(n6272), .B(n6262), .Y(n6273));
  OAI22X1 g5153(.A0(n6206), .A1(n6046), .B0(n6045), .B1(n6270), .Y(n6274));
  AOI21X1 g5154(.A0(n6035), .A1(n5897), .B0(n6270), .Y(n6275));
  NAND2X1 g5155(.A(n6261), .B(n5913), .Y(n6276));
  AOI22X1 g5156(.A0(n5957), .A1(P2_REG0_REG_9__SCAN_IN), .B0(P2_REG2_REG_9__SCAN_IN), .B1(n5958), .Y(n6277));
  INVX1   g5157(.A(P2_REG3_REG_9__SCAN_IN), .Y(n6278));
  NOR2X1  g5158(.A(n6238), .B(P2_REG3_REG_8__SCAN_IN), .Y(n6279));
  NOR2X1  g5159(.A(P2_REG3_REG_9__SCAN_IN), .B(P2_REG3_REG_8__SCAN_IN), .Y(n6280));
  INVX1   g5160(.A(n6280), .Y(n6281));
  OAI22X1 g5161(.A0(n6279), .A1(n6278), .B0(n6238), .B1(n6281), .Y(n6282));
  AOI22X1 g5162(.A0(n5962), .A1(n6282), .B0(n5961), .B1(P2_REG1_REG_9__SCAN_IN), .Y(n6283));
  NAND2X1 g5163(.A(n6283), .B(n6277), .Y(n6284));
  AOI22X1 g5164(.A0(n6254), .A1(n6008), .B0(n5917), .B1(n6284), .Y(n6285));
  NAND2X1 g5165(.A(n6285), .B(n6276), .Y(n6286));
  NOR4X1  g5166(.A(n6275), .B(n6274), .C(n6273), .D(n6286), .Y(n6287));
  NAND2X1 g5167(.A(n5970), .B(P2_REG0_REG_8__SCAN_IN), .Y(n6288));
  OAI21X1 g5168(.A0(n6287), .A1(n5970), .B0(n6288), .Y(P2_U3414));
  NOR2X1  g5169(.A(n5870), .B(n5523), .Y(n6290));
  AOI21X1 g5170(.A0(n6252), .A1(n5870), .B0(n6290), .Y(n6291));
  NAND2X1 g5171(.A(n6291), .B(n6249), .Y(n6292));
  NOR2X1  g5172(.A(n6291), .B(n6249), .Y(n6293));
  AOI21X1 g5173(.A0(n6292), .A1(n6265), .B0(n6293), .Y(n6294));
  INVX1   g5174(.A(n6294), .Y(n6295));
  INVX1   g5175(.A(n6284), .Y(n6296));
  NOR2X1  g5176(.A(P2_IR_REG_31__SCAN_IN), .B(n5539), .Y(n6297));
  AOI21X1 g5177(.A0(n5534), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6297), .Y(n6298));
  INVX1   g5178(.A(n6298), .Y(n6299));
  NAND2X1 g5179(.A(n6299), .B(n5870), .Y(n6300));
  OAI21X1 g5180(.A0(n5870), .A1(n5533), .B0(n6300), .Y(n6301));
  XOR2X1  g5181(.A(n6301), .B(n6296), .Y(n6302));
  NOR2X1  g5182(.A(n6295), .B(n6302), .Y(n6303));
  AOI21X1 g5183(.A0(n6302), .A1(n6295), .B0(n6303), .Y(n6305));
  NOR2X1  g5184(.A(n6305), .B(n6045), .Y(n6306));
  AOI22X1 g5185(.A0(n6249), .A1(n6254), .B0(n6211), .B1(n6206), .Y(n6307));
  NAND2X1 g5186(.A(n6307), .B(n6216), .Y(n6308));
  NOR2X1  g5187(.A(n6308), .B(n6084), .Y(n6309));
  NAND2X1 g5188(.A(n6307), .B(n6215), .Y(n6310));
  OAI21X1 g5189(.A0(n6242), .A1(n6228), .B0(n6291), .Y(n6311));
  NAND2X1 g5190(.A(n6242), .B(n6228), .Y(n6312));
  NAND3X1 g5191(.A(n6312), .B(n6311), .C(n6310), .Y(n6313));
  NOR2X1  g5192(.A(n6313), .B(n6309), .Y(n6314));
  XOR2X1  g5193(.A(n6314), .B(n6302), .Y(n6315));
  INVX1   g5194(.A(n6315), .Y(n6316));
  AOI22X1 g5195(.A0(n6242), .A1(n5952), .B0(n5908), .B1(n6316), .Y(n6317));
  OAI21X1 g5196(.A0(n5909), .A1(n5902), .B0(n6316), .Y(n6318));
  NAND2X1 g5197(.A(n6318), .B(n6317), .Y(n6319));
  NOR2X1  g5198(.A(n6305), .B(n6018), .Y(n6320));
  AOI21X1 g5199(.A0(n6035), .A1(n5897), .B0(n6305), .Y(n6321));
  NOR4X1  g5200(.A(n6320), .B(n6319), .C(n6306), .D(n6321), .Y(n6322));
  INVX1   g5201(.A(n6322), .Y(n6323));
  AOI22X1 g5202(.A0(n5957), .A1(P2_REG0_REG_10__SCAN_IN), .B0(P2_REG2_REG_10__SCAN_IN), .B1(n5958), .Y(n6324));
  INVX1   g5203(.A(n6324), .Y(n6325));
  INVX1   g5204(.A(P2_REG3_REG_10__SCAN_IN), .Y(n6326));
  NOR2X1  g5205(.A(n6281), .B(n6238), .Y(n6327));
  NOR3X1  g5206(.A(n6281), .B(n6238), .C(P2_REG3_REG_10__SCAN_IN), .Y(n6328));
  INVX1   g5207(.A(n6328), .Y(n6329));
  OAI21X1 g5208(.A0(n6327), .A1(n6326), .B0(n6329), .Y(n6330));
  AOI22X1 g5209(.A0(n5962), .A1(n6330), .B0(n5961), .B1(P2_REG1_REG_10__SCAN_IN), .Y(n6331));
  INVX1   g5210(.A(n6331), .Y(n6332));
  NOR2X1  g5211(.A(n6332), .B(n6325), .Y(n6333));
  INVX1   g5212(.A(n6333), .Y(n6334));
  AOI22X1 g5213(.A0(n6301), .A1(n6008), .B0(n5917), .B1(n6334), .Y(n6335));
  OAI21X1 g5214(.A0(n6315), .A1(n6007), .B0(n6335), .Y(n6336));
  NOR2X1  g5215(.A(n6336), .B(n6323), .Y(n6337));
  NAND2X1 g5216(.A(n5970), .B(P2_REG0_REG_9__SCAN_IN), .Y(n6338));
  OAI21X1 g5217(.A0(n6337), .A1(n5970), .B0(n6338), .Y(P2_U3417));
  NAND2X1 g5218(.A(n6301), .B(n6284), .Y(n6340));
  INVX1   g5219(.A(P2_IR_REG_10__SCAN_IN), .Y(n6341));
  NOR2X1  g5220(.A(P2_IR_REG_31__SCAN_IN), .B(n6341), .Y(n6342));
  AOI21X1 g5221(.A0(n5542), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6342), .Y(n6343));
  INVX1   g5222(.A(n6343), .Y(n6344));
  NOR2X1  g5223(.A(n5870), .B(n5538), .Y(n6345));
  AOI21X1 g5224(.A0(n6344), .A1(n5870), .B0(n6345), .Y(n6346));
  NOR2X1  g5225(.A(n6301), .B(n6284), .Y(n6347));
  AOI21X1 g5226(.A0(n6346), .A1(n6333), .B0(n6347), .Y(n6348));
  OAI21X1 g5227(.A0(n6346), .A1(n6333), .B0(n6348), .Y(n6349));
  AOI21X1 g5228(.A0(n6340), .A1(n6294), .B0(n6349), .Y(n6350));
  NOR2X1  g5229(.A(n6347), .B(n6294), .Y(n6351));
  NAND2X1 g5230(.A(n6344), .B(n5870), .Y(n6352));
  OAI21X1 g5231(.A0(n5870), .A1(n5538), .B0(n6352), .Y(n6353));
  XOR2X1  g5232(.A(n6353), .B(n6333), .Y(n6354));
  NAND2X1 g5233(.A(n6354), .B(n6340), .Y(n6355));
  NOR2X1  g5234(.A(n6355), .B(n6351), .Y(n6356));
  NOR2X1  g5235(.A(n6356), .B(n6350), .Y(n6357));
  INVX1   g5236(.A(n6357), .Y(n6358));
  NOR2X1  g5237(.A(n6301), .B(n6296), .Y(n6359));
  INVX1   g5238(.A(n6301), .Y(n6360));
  NOR2X1  g5239(.A(n6360), .B(n6284), .Y(n6361));
  INVX1   g5240(.A(n6361), .Y(n6362));
  INVX1   g5241(.A(n6314), .Y(n6363));
  AOI21X1 g5242(.A0(n6363), .A1(n6362), .B0(n6359), .Y(n6364));
  XOR2X1  g5243(.A(n6364), .B(n6354), .Y(n6365));
  OAI22X1 g5244(.A0(n6296), .A1(n6046), .B0(n6002), .B1(n6365), .Y(n6366));
  AOI21X1 g5245(.A0(n6003), .A1(n5991), .B0(n6365), .Y(n6367));
  NOR2X1  g5246(.A(n6367), .B(n6366), .Y(n6368));
  OAI21X1 g5247(.A0(n6358), .A1(n6045), .B0(n6368), .Y(n6369));
  NOR3X1  g5248(.A(n6356), .B(n6350), .C(n6018), .Y(n6370));
  AOI21X1 g5249(.A0(n6035), .A1(n5897), .B0(n6358), .Y(n6371));
  NAND3X1 g5250(.A(n5884), .B(n5882), .C(P2_REG0_REG_11__SCAN_IN), .Y(n6372));
  NAND3X1 g5251(.A(n5884), .B(n5888), .C(P2_REG2_REG_11__SCAN_IN), .Y(n6373));
  NAND3X1 g5252(.A(n5891), .B(n5882), .C(P2_REG1_REG_11__SCAN_IN), .Y(n6374));
  NOR4X1  g5253(.A(n6238), .B(P2_REG3_REG_11__SCAN_IN), .C(P2_REG3_REG_10__SCAN_IN), .D(n6281), .Y(n6375));
  AOI21X1 g5254(.A0(n6329), .A1(P2_REG3_REG_11__SCAN_IN), .B0(n6375), .Y(n6376));
  INVX1   g5255(.A(n6376), .Y(n6377));
  NAND3X1 g5256(.A(n6377), .B(n5891), .C(n5888), .Y(n6378));
  NAND4X1 g5257(.A(n6374), .B(n6373), .C(n6372), .D(n6378), .Y(n6379));
  AOI22X1 g5258(.A0(n6353), .A1(n6008), .B0(n5917), .B1(n6379), .Y(n6380));
  OAI21X1 g5259(.A0(n6365), .A1(n6007), .B0(n6380), .Y(n6381));
  NOR4X1  g5260(.A(n6371), .B(n6370), .C(n6369), .D(n6381), .Y(n6382));
  NAND2X1 g5261(.A(n5970), .B(P2_REG0_REG_10__SCAN_IN), .Y(n6383));
  OAI21X1 g5262(.A0(n6382), .A1(n5970), .B0(n6383), .Y(P2_U3420));
  INVX1   g5263(.A(n6364), .Y(n6385));
  AOI21X1 g5264(.A0(n6346), .A1(n6334), .B0(n6385), .Y(n6386));
  NAND2X1 g5265(.A(n6353), .B(n6333), .Y(n6387));
  INVX1   g5266(.A(n6387), .Y(n6388));
  NOR2X1  g5267(.A(P2_IR_REG_31__SCAN_IN), .B(n5547), .Y(n6389));
  AOI21X1 g5268(.A0(n5548), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6389), .Y(n6390));
  INVX1   g5269(.A(n6390), .Y(n6391));
  NOR2X1  g5270(.A(n5870), .B(n5546), .Y(n6392));
  AOI21X1 g5271(.A0(n6391), .A1(n5870), .B0(n6392), .Y(n6393));
  XOR2X1  g5272(.A(n6393), .B(n6379), .Y(n6394));
  NOR2X1  g5273(.A(n6394), .B(n6388), .Y(n6395));
  INVX1   g5274(.A(n6395), .Y(n6396));
  NOR2X1  g5275(.A(n6393), .B(n6379), .Y(n6397));
  AOI22X1 g5276(.A0(n6379), .A1(n6393), .B0(n6346), .B1(n6334), .Y(n6398));
  INVX1   g5277(.A(n6398), .Y(n6399));
  NOR2X1  g5278(.A(n6399), .B(n6397), .Y(n6400));
  OAI21X1 g5279(.A0(n6364), .A1(n6388), .B0(n6400), .Y(n6401));
  OAI21X1 g5280(.A0(n6396), .A1(n6386), .B0(n6401), .Y(n6402));
  INVX1   g5281(.A(n6402), .Y(n6403));
  AOI21X1 g5282(.A0(n6003), .A1(n5991), .B0(n6403), .Y(n6404));
  NAND3X1 g5283(.A(n6348), .B(n6292), .C(n6265), .Y(n6406));
  AOI22X1 g5284(.A0(n6301), .A1(n6284), .B0(n6293), .B1(n6348), .Y(n6407));
  AOI21X1 g5285(.A0(n6346), .A1(n6333), .B0(n6407), .Y(n6408));
  AOI21X1 g5286(.A0(n6353), .A1(n6334), .B0(n6408), .Y(n6409));
  NAND2X1 g5287(.A(n6409), .B(n6406), .Y(n6410));
  INVX1   g5288(.A(n6410), .Y(n6411));
  INVX1   g5289(.A(n6379), .Y(n6412));
  XOR2X1  g5290(.A(n6393), .B(n6412), .Y(n6413));
  AOI21X1 g5291(.A0(n6409), .A1(n6406), .B0(n6413), .Y(n6414));
  AOI21X1 g5292(.A0(n6411), .A1(n6413), .B0(n6414), .Y(n6415));
  OAI22X1 g5293(.A0(n6403), .A1(n6002), .B0(n6018), .B1(n6415), .Y(n6416));
  OAI22X1 g5294(.A0(n6333), .A1(n6046), .B0(n6045), .B1(n6415), .Y(n6417));
  NOR2X1  g5295(.A(n6410), .B(n6394), .Y(n6418));
  OAI22X1 g5296(.A0(n6418), .A1(n6414), .B0(n5904), .B1(n5896), .Y(n6419));
  INVX1   g5297(.A(n6419), .Y(n6420));
  NOR4X1  g5298(.A(n6417), .B(n6416), .C(n6404), .D(n6420), .Y(n6421));
  INVX1   g5299(.A(n6421), .Y(n6422));
  INVX1   g5300(.A(n6393), .Y(n6423));
  AOI22X1 g5301(.A0(n5957), .A1(P2_REG0_REG_12__SCAN_IN), .B0(P2_REG2_REG_12__SCAN_IN), .B1(n5958), .Y(n6424));
  INVX1   g5302(.A(P2_REG3_REG_12__SCAN_IN), .Y(n6425));
  XOR2X1  g5303(.A(n6375), .B(n6425), .Y(n6426));
  INVX1   g5304(.A(n6426), .Y(n6427));
  AOI22X1 g5305(.A0(n5962), .A1(n6427), .B0(n5961), .B1(P2_REG1_REG_12__SCAN_IN), .Y(n6428));
  NAND2X1 g5306(.A(n6428), .B(n6424), .Y(n6429));
  AOI22X1 g5307(.A0(n6423), .A1(n6008), .B0(n5917), .B1(n6429), .Y(n6430));
  OAI21X1 g5308(.A0(n6403), .A1(n6007), .B0(n6430), .Y(n6431));
  NOR2X1  g5309(.A(n6431), .B(n6422), .Y(n6432));
  NAND2X1 g5310(.A(n5970), .B(P2_REG0_REG_11__SCAN_IN), .Y(n6433));
  OAI21X1 g5311(.A0(n6432), .A1(n5970), .B0(n6433), .Y(P2_U3423));
  NOR2X1  g5312(.A(n6393), .B(n6412), .Y(n6435));
  INVX1   g5313(.A(n6429), .Y(n6436));
  NOR2X1  g5314(.A(P2_IR_REG_31__SCAN_IN), .B(n5554), .Y(n6437));
  AOI21X1 g5315(.A0(n5559), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6437), .Y(n6438));
  INVX1   g5316(.A(n6438), .Y(n6439));
  NAND2X1 g5317(.A(n6439), .B(n5870), .Y(n6440));
  OAI21X1 g5318(.A0(n5870), .A1(n5553), .B0(n6440), .Y(n6441));
  XOR2X1  g5319(.A(n6441), .B(n6436), .Y(n6442));
  AOI22X1 g5320(.A0(n6406), .A1(n6409), .B0(n6393), .B1(n6412), .Y(n6443));
  NOR3X1  g5321(.A(n6443), .B(n6442), .C(n6435), .Y(n6444));
  NOR2X1  g5322(.A(n6443), .B(n6435), .Y(n6445));
  XOR2X1  g5323(.A(n6441), .B(n6429), .Y(n6446));
  NOR2X1  g5324(.A(n6446), .B(n6445), .Y(n6447));
  NOR2X1  g5325(.A(n6447), .B(n6444), .Y(n6448));
  NOR2X1  g5326(.A(n6448), .B(n6045), .Y(n6449));
  NOR4X1  g5327(.A(n6388), .B(n6314), .C(n6361), .D(n6397), .Y(n6450));
  NAND2X1 g5328(.A(n6387), .B(n6359), .Y(n6451));
  AOI21X1 g5329(.A0(n6451), .A1(n6398), .B0(n6397), .Y(n6452));
  NOR2X1  g5330(.A(n6452), .B(n6450), .Y(n6453));
  XOR2X1  g5331(.A(n6453), .B(n6442), .Y(n6454));
  INVX1   g5332(.A(n6454), .Y(n6455));
  AOI22X1 g5333(.A0(n6379), .A1(n5952), .B0(n5908), .B1(n6455), .Y(n6456));
  OAI21X1 g5334(.A0(n5909), .A1(n5902), .B0(n6455), .Y(n6457));
  NAND2X1 g5335(.A(n6457), .B(n6456), .Y(n6458));
  NOR2X1  g5336(.A(n6448), .B(n6018), .Y(n6459));
  AOI21X1 g5337(.A0(n6035), .A1(n5897), .B0(n6448), .Y(n6460));
  NOR4X1  g5338(.A(n6459), .B(n6458), .C(n6449), .D(n6460), .Y(n6461));
  INVX1   g5339(.A(n6461), .Y(n6462));
  AOI22X1 g5340(.A0(n5957), .A1(P2_REG0_REG_13__SCAN_IN), .B0(P2_REG2_REG_13__SCAN_IN), .B1(n5958), .Y(n6463));
  INVX1   g5341(.A(n6375), .Y(n6464));
  NOR2X1  g5342(.A(P2_REG3_REG_13__SCAN_IN), .B(P2_REG3_REG_12__SCAN_IN), .Y(n6465));
  INVX1   g5343(.A(n6465), .Y(n6466));
  OAI21X1 g5344(.A0(n6464), .A1(P2_REG3_REG_12__SCAN_IN), .B0(P2_REG3_REG_13__SCAN_IN), .Y(n6467));
  OAI21X1 g5345(.A0(n6466), .A1(n6464), .B0(n6467), .Y(n6468));
  AOI22X1 g5346(.A0(n5962), .A1(n6468), .B0(n5961), .B1(P2_REG1_REG_13__SCAN_IN), .Y(n6469));
  NAND2X1 g5347(.A(n6469), .B(n6463), .Y(n6470));
  AOI22X1 g5348(.A0(n6441), .A1(n6008), .B0(n5917), .B1(n6470), .Y(n6471));
  OAI21X1 g5349(.A0(n6454), .A1(n6007), .B0(n6471), .Y(n6472));
  NOR2X1  g5350(.A(n6472), .B(n6462), .Y(n6473));
  NAND2X1 g5351(.A(n5970), .B(P2_REG0_REG_12__SCAN_IN), .Y(n6474));
  OAI21X1 g5352(.A0(n6473), .A1(n5970), .B0(n6474), .Y(P2_U3426));
  NOR2X1  g5353(.A(n5870), .B(n5553), .Y(n6476));
  AOI21X1 g5354(.A0(n6439), .A1(n5870), .B0(n6476), .Y(n6477));
  NOR2X1  g5355(.A(n6477), .B(n6436), .Y(n6478));
  NOR3X1  g5356(.A(n6478), .B(n6443), .C(n6435), .Y(n6479));
  INVX1   g5357(.A(n6470), .Y(n6480));
  NOR2X1  g5358(.A(P2_IR_REG_31__SCAN_IN), .B(n5570), .Y(n6481));
  AOI21X1 g5359(.A0(n5564), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6481), .Y(n6482));
  INVX1   g5360(.A(n6482), .Y(n6483));
  NAND2X1 g5361(.A(n6483), .B(n5870), .Y(n6484));
  OAI21X1 g5362(.A0(n5870), .A1(n5563), .B0(n6484), .Y(n6485));
  INVX1   g5363(.A(n6485), .Y(n6486));
  OAI22X1 g5364(.A0(n6470), .A1(n6485), .B0(n6441), .B1(n6429), .Y(n6487));
  INVX1   g5365(.A(n6487), .Y(n6488));
  OAI21X1 g5366(.A0(n6486), .A1(n6480), .B0(n6488), .Y(n6489));
  AOI21X1 g5367(.A0(n6477), .A1(n6436), .B0(n6445), .Y(n6490));
  XOR2X1  g5368(.A(n6485), .B(n6480), .Y(n6491));
  OAI21X1 g5369(.A0(n6477), .A1(n6436), .B0(n6491), .Y(n6492));
  OAI22X1 g5370(.A0(n6490), .A1(n6492), .B0(n6489), .B1(n6479), .Y(n6493));
  NOR2X1  g5371(.A(n6477), .B(n6429), .Y(n6494));
  NOR4X1  g5372(.A(n6397), .B(n6388), .C(n6361), .D(n6494), .Y(n6495));
  OAI21X1 g5373(.A0(n6313), .A1(n6309), .B0(n6495), .Y(n6496));
  INVX1   g5374(.A(n6496), .Y(n6497));
  NOR2X1  g5375(.A(n6441), .B(n6436), .Y(n6498));
  NAND2X1 g5376(.A(n6441), .B(n6436), .Y(n6499));
  AOI21X1 g5377(.A0(n6452), .A1(n6499), .B0(n6498), .Y(n6500));
  INVX1   g5378(.A(n6500), .Y(n6501));
  NOR2X1  g5379(.A(n6501), .B(n6497), .Y(n6502));
  XOR2X1  g5380(.A(n6502), .B(n6491), .Y(n6503));
  OAI22X1 g5381(.A0(n6436), .A1(n6046), .B0(n6002), .B1(n6503), .Y(n6504));
  AOI21X1 g5382(.A0(n6003), .A1(n5991), .B0(n6503), .Y(n6505));
  NOR2X1  g5383(.A(n6505), .B(n6504), .Y(n6506));
  OAI21X1 g5384(.A0(n6493), .A1(n6045), .B0(n6506), .Y(n6507));
  NOR2X1  g5385(.A(n6493), .B(n6018), .Y(n6508));
  AOI21X1 g5386(.A0(n6035), .A1(n5897), .B0(n6493), .Y(n6509));
  AOI22X1 g5387(.A0(n5957), .A1(P2_REG0_REG_14__SCAN_IN), .B0(P2_REG2_REG_14__SCAN_IN), .B1(n5958), .Y(n6510));
  INVX1   g5388(.A(P2_REG3_REG_14__SCAN_IN), .Y(n6511));
  NOR2X1  g5389(.A(n6466), .B(n6464), .Y(n6512));
  XOR2X1  g5390(.A(n6512), .B(n6511), .Y(n6513));
  INVX1   g5391(.A(n6513), .Y(n6514));
  AOI22X1 g5392(.A0(n5962), .A1(n6514), .B0(n5961), .B1(P2_REG1_REG_14__SCAN_IN), .Y(n6515));
  NAND2X1 g5393(.A(n6515), .B(n6510), .Y(n6516));
  AOI22X1 g5394(.A0(n6485), .A1(n6008), .B0(n5917), .B1(n6516), .Y(n6517));
  OAI21X1 g5395(.A0(n6503), .A1(n6007), .B0(n6517), .Y(n6518));
  NOR4X1  g5396(.A(n6509), .B(n6508), .C(n6507), .D(n6518), .Y(n6519));
  NAND2X1 g5397(.A(n5970), .B(P2_REG0_REG_13__SCAN_IN), .Y(n6520));
  OAI21X1 g5398(.A0(n6519), .A1(n5970), .B0(n6520), .Y(P2_U3429));
  NOR2X1  g5399(.A(n6485), .B(n6480), .Y(n6522));
  INVX1   g5400(.A(n6522), .Y(n6523));
  AOI22X1 g5401(.A0(n6496), .A1(n6500), .B0(n6485), .B1(n6480), .Y(n6524));
  INVX1   g5402(.A(n6524), .Y(n6525));
  NAND2X1 g5403(.A(n6525), .B(n6523), .Y(n6526));
  INVX1   g5404(.A(n6516), .Y(n6527));
  NOR2X1  g5405(.A(P2_IR_REG_31__SCAN_IN), .B(n5571), .Y(n6528));
  AOI21X1 g5406(.A0(n5574), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6528), .Y(n6529));
  INVX1   g5407(.A(n6529), .Y(n6530));
  NAND2X1 g5408(.A(n6530), .B(n5870), .Y(n6531));
  OAI21X1 g5409(.A0(n5870), .A1(n5569), .B0(n6531), .Y(n6532));
  XOR2X1  g5410(.A(n6532), .B(n6527), .Y(n6533));
  INVX1   g5411(.A(n6533), .Y(n6534));
  XOR2X1  g5412(.A(n6534), .B(n6526), .Y(n6535));
  INVX1   g5413(.A(n6535), .Y(n6536));
  AOI22X1 g5414(.A0(n6470), .A1(n5952), .B0(n5908), .B1(n6536), .Y(n6537));
  OAI21X1 g5415(.A0(n5909), .A1(n5902), .B0(n6536), .Y(n6538));
  AOI21X1 g5416(.A0(n6393), .A1(n6412), .B0(n6487), .Y(n6539));
  NOR3X1  g5417(.A(n6487), .B(n6393), .C(n6412), .Y(n6540));
  OAI22X1 g5418(.A0(n6485), .A1(n6470), .B0(n6478), .B1(n6540), .Y(n6541));
  OAI21X1 g5419(.A0(n6486), .A1(n6480), .B0(n6541), .Y(n6542));
  AOI21X1 g5420(.A0(n6539), .A1(n6410), .B0(n6542), .Y(n6543));
  XOR2X1  g5421(.A(n6543), .B(n6534), .Y(n6544));
  INVX1   g5422(.A(n6544), .Y(n6545));
  OAI21X1 g5423(.A0(n5905), .A1(n5904), .B0(n6545), .Y(n6546));
  OAI21X1 g5424(.A0(n5901), .A1(n5896), .B0(n6545), .Y(n6547));
  NAND4X1 g5425(.A(n6546), .B(n6538), .C(n6537), .D(n6547), .Y(n6548));
  AOI22X1 g5426(.A0(n5957), .A1(P2_REG0_REG_15__SCAN_IN), .B0(P2_REG2_REG_15__SCAN_IN), .B1(n5958), .Y(n6549));
  INVX1   g5427(.A(n6549), .Y(n6550));
  INVX1   g5428(.A(P2_REG1_REG_15__SCAN_IN), .Y(n6551));
  NOR3X1  g5429(.A(n5884), .B(n5888), .C(n6551), .Y(n6552));
  NOR4X1  g5430(.A(n6464), .B(P2_REG3_REG_15__SCAN_IN), .C(P2_REG3_REG_14__SCAN_IN), .D(n6466), .Y(n6553));
  INVX1   g5431(.A(P2_REG3_REG_15__SCAN_IN), .Y(n6554));
  AOI21X1 g5432(.A0(n6512), .A1(n6511), .B0(n6554), .Y(n6555));
  NOR2X1  g5433(.A(n6555), .B(n6553), .Y(n6556));
  NOR3X1  g5434(.A(n6556), .B(n5884), .C(n5882), .Y(n6557));
  NOR3X1  g5435(.A(n6557), .B(n6552), .C(n6550), .Y(n6558));
  INVX1   g5436(.A(n6558), .Y(n6559));
  AOI22X1 g5437(.A0(n6532), .A1(n6008), .B0(n5917), .B1(n6559), .Y(n6560));
  OAI21X1 g5438(.A0(n6535), .A1(n6007), .B0(n6560), .Y(n6561));
  NOR2X1  g5439(.A(n6561), .B(n6548), .Y(n6562));
  NAND2X1 g5440(.A(n5970), .B(P2_REG0_REG_14__SCAN_IN), .Y(n6563));
  OAI21X1 g5441(.A0(n6562), .A1(n5970), .B0(n6563), .Y(P2_U3432));
  NOR2X1  g5442(.A(P2_IR_REG_31__SCAN_IN), .B(n5580), .Y(n6565));
  AOI21X1 g5443(.A0(n5581), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6565), .Y(n6566));
  INVX1   g5444(.A(n6566), .Y(n6567));
  NAND2X1 g5445(.A(n6567), .B(n5870), .Y(n6568));
  OAI21X1 g5446(.A0(n5870), .A1(n5579), .B0(n6568), .Y(n6569));
  XOR2X1  g5447(.A(n6569), .B(n6558), .Y(n6570));
  NOR2X1  g5448(.A(n6532), .B(n6527), .Y(n6571));
  INVX1   g5449(.A(n6532), .Y(n6572));
  NOR2X1  g5450(.A(n6572), .B(n6516), .Y(n6573));
  INVX1   g5451(.A(n6573), .Y(n6574));
  AOI21X1 g5452(.A0(n6574), .A1(n6526), .B0(n6571), .Y(n6575));
  XOR2X1  g5453(.A(n6575), .B(n6570), .Y(n6576));
  INVX1   g5454(.A(n6576), .Y(n6577));
  AOI22X1 g5455(.A0(n6516), .A1(n5952), .B0(n5908), .B1(n6577), .Y(n6578));
  OAI21X1 g5456(.A0(n5909), .A1(n5902), .B0(n6577), .Y(n6579));
  NAND2X1 g5457(.A(n6532), .B(n6516), .Y(n6580));
  NOR2X1  g5458(.A(n6532), .B(n6516), .Y(n6581));
  OAI21X1 g5459(.A0(n6581), .A1(n6543), .B0(n6580), .Y(n6582));
  XOR2X1  g5460(.A(n6582), .B(n6570), .Y(n6583));
  INVX1   g5461(.A(n6583), .Y(n6584));
  OAI21X1 g5462(.A0(n5905), .A1(n5904), .B0(n6584), .Y(n6585));
  OAI21X1 g5463(.A0(n5901), .A1(n5896), .B0(n6584), .Y(n6586));
  NAND4X1 g5464(.A(n6585), .B(n6579), .C(n6578), .D(n6586), .Y(n6587));
  AOI22X1 g5465(.A0(n5957), .A1(P2_REG0_REG_16__SCAN_IN), .B0(P2_REG2_REG_16__SCAN_IN), .B1(n5958), .Y(n6588));
  INVX1   g5466(.A(P2_REG3_REG_16__SCAN_IN), .Y(n6589));
  XOR2X1  g5467(.A(n6553), .B(n6589), .Y(n6590));
  INVX1   g5468(.A(n6590), .Y(n6591));
  AOI22X1 g5469(.A0(n5962), .A1(n6591), .B0(n5961), .B1(P2_REG1_REG_16__SCAN_IN), .Y(n6592));
  NAND2X1 g5470(.A(n6592), .B(n6588), .Y(n6593));
  AOI22X1 g5471(.A0(n6569), .A1(n6008), .B0(n5917), .B1(n6593), .Y(n6594));
  OAI21X1 g5472(.A0(n6576), .A1(n6007), .B0(n6594), .Y(n6595));
  NOR2X1  g5473(.A(n6595), .B(n6587), .Y(n6596));
  NAND2X1 g5474(.A(n5970), .B(P2_REG0_REG_15__SCAN_IN), .Y(n6597));
  OAI21X1 g5475(.A0(n6596), .A1(n5970), .B0(n6597), .Y(P2_U3435));
  INVX1   g5476(.A(n6593), .Y(n6599));
  NOR2X1  g5477(.A(P2_IR_REG_31__SCAN_IN), .B(n5587), .Y(n6600));
  AOI21X1 g5478(.A0(n5592), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6600), .Y(n6601));
  INVX1   g5479(.A(n6601), .Y(n6602));
  NAND2X1 g5480(.A(n6602), .B(n5870), .Y(n6603));
  OAI21X1 g5481(.A0(n5870), .A1(n5586), .B0(n6603), .Y(n6604));
  XOR2X1  g5482(.A(n6604), .B(n6599), .Y(n6605));
  INVX1   g5483(.A(n6569), .Y(n6607));
  NOR2X1  g5484(.A(n6607), .B(n6558), .Y(n6608));
  NAND2X1 g5485(.A(n6607), .B(n6558), .Y(n6609));
  AOI21X1 g5486(.A0(n6609), .A1(n6582), .B0(n6608), .Y(n6610));
  XOR2X1  g5487(.A(n6604), .B(n6593), .Y(n6611));
  NOR2X1  g5488(.A(n6611), .B(n6610), .Y(n6612));
  AOI21X1 g5489(.A0(n6610), .A1(n6611), .B0(n6612), .Y(n6613));
  NOR2X1  g5490(.A(n6613), .B(n6045), .Y(n6614));
  INVX1   g5491(.A(n6575), .Y(n6615));
  AOI21X1 g5492(.A0(n6607), .A1(n6559), .B0(n6615), .Y(n6616));
  NAND2X1 g5493(.A(n6569), .B(n6558), .Y(n6617));
  INVX1   g5494(.A(n6617), .Y(n6618));
  NOR2X1  g5495(.A(n6605), .B(n6618), .Y(n6619));
  INVX1   g5496(.A(n6619), .Y(n6620));
  NAND2X1 g5497(.A(n6604), .B(n6599), .Y(n6621));
  INVX1   g5498(.A(n6621), .Y(n6622));
  INVX1   g5499(.A(n6604), .Y(n6623));
  AOI22X1 g5500(.A0(n6593), .A1(n6623), .B0(n6607), .B1(n6559), .Y(n6624));
  INVX1   g5501(.A(n6624), .Y(n6625));
  NOR2X1  g5502(.A(n6625), .B(n6622), .Y(n6626));
  OAI21X1 g5503(.A0(n6575), .A1(n6618), .B0(n6626), .Y(n6627));
  OAI21X1 g5504(.A0(n6620), .A1(n6616), .B0(n6627), .Y(n6628));
  AOI22X1 g5505(.A0(n6559), .A1(n5952), .B0(n5908), .B1(n6628), .Y(n6629));
  OAI21X1 g5506(.A0(n5909), .A1(n5902), .B0(n6628), .Y(n6630));
  NAND2X1 g5507(.A(n6630), .B(n6629), .Y(n6631));
  INVX1   g5508(.A(n6610), .Y(n6632));
  NOR2X1  g5509(.A(n6632), .B(n6605), .Y(n6633));
  OAI22X1 g5510(.A0(n6633), .A1(n6612), .B0(n5904), .B1(n5896), .Y(n6634));
  OAI21X1 g5511(.A0(n6613), .A1(n6018), .B0(n6634), .Y(n6635));
  NAND2X1 g5512(.A(n6628), .B(n5913), .Y(n6636));
  AOI22X1 g5513(.A0(n5957), .A1(P2_REG0_REG_17__SCAN_IN), .B0(P2_REG2_REG_17__SCAN_IN), .B1(n5958), .Y(n6637));
  INVX1   g5514(.A(P2_REG3_REG_17__SCAN_IN), .Y(n6638));
  INVX1   g5515(.A(n6553), .Y(n6639));
  NOR2X1  g5516(.A(n6639), .B(P2_REG3_REG_16__SCAN_IN), .Y(n6640));
  NOR3X1  g5517(.A(n6639), .B(P2_REG3_REG_17__SCAN_IN), .C(P2_REG3_REG_16__SCAN_IN), .Y(n6641));
  INVX1   g5518(.A(n6641), .Y(n6642));
  OAI21X1 g5519(.A0(n6640), .A1(n6638), .B0(n6642), .Y(n6643));
  AOI22X1 g5520(.A0(n5962), .A1(n6643), .B0(n5961), .B1(P2_REG1_REG_17__SCAN_IN), .Y(n6644));
  NAND2X1 g5521(.A(n6644), .B(n6637), .Y(n6645));
  AOI22X1 g5522(.A0(n6604), .A1(n6008), .B0(n5917), .B1(n6645), .Y(n6646));
  NAND2X1 g5523(.A(n6646), .B(n6636), .Y(n6647));
  NOR4X1  g5524(.A(n6635), .B(n6631), .C(n6614), .D(n6647), .Y(n6648));
  NAND2X1 g5525(.A(n5970), .B(P2_REG0_REG_16__SCAN_IN), .Y(n6649));
  OAI21X1 g5526(.A0(n6648), .A1(n5970), .B0(n6649), .Y(P2_U3438));
  NAND2X1 g5527(.A(n6604), .B(n6593), .Y(n6651));
  INVX1   g5528(.A(n6651), .Y(n6652));
  NOR2X1  g5529(.A(P2_IR_REG_31__SCAN_IN), .B(n5598), .Y(n6653));
  AOI21X1 g5530(.A0(n5600), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6653), .Y(n6654));
  INVX1   g5531(.A(n6654), .Y(n6655));
  NOR2X1  g5532(.A(n5870), .B(n5597), .Y(n6656));
  AOI21X1 g5533(.A0(n6655), .A1(n5870), .B0(n6656), .Y(n6657));
  INVX1   g5534(.A(n6657), .Y(n6658));
  OAI22X1 g5535(.A0(n6645), .A1(n6658), .B0(n6604), .B1(n6593), .Y(n6659));
  AOI21X1 g5536(.A0(n6658), .A1(n6645), .B0(n6659), .Y(n6660));
  OAI21X1 g5537(.A0(n6652), .A1(n6632), .B0(n6660), .Y(n6661));
  AOI21X1 g5538(.A0(n6623), .A1(n6599), .B0(n6610), .Y(n6662));
  XOR2X1  g5539(.A(n6657), .B(n6645), .Y(n6663));
  NAND2X1 g5540(.A(n6663), .B(n6651), .Y(n6664));
  OAI21X1 g5541(.A0(n6664), .A1(n6662), .B0(n6661), .Y(n6665));
  NAND3X1 g5542(.A(n6621), .B(n6617), .C(n6571), .Y(n6666));
  AOI21X1 g5543(.A0(n6666), .A1(n6624), .B0(n6622), .Y(n6667));
  NOR3X1  g5544(.A(n6622), .B(n6618), .C(n6573), .Y(n6668));
  OAI21X1 g5545(.A0(n6524), .A1(n6522), .B0(n6668), .Y(n6669));
  INVX1   g5546(.A(n6669), .Y(n6670));
  NOR2X1  g5547(.A(n6670), .B(n6667), .Y(n6671));
  XOR2X1  g5548(.A(n6671), .B(n6663), .Y(n6672));
  OAI22X1 g5549(.A0(n6599), .A1(n6046), .B0(n6002), .B1(n6672), .Y(n6673));
  AOI21X1 g5550(.A0(n6003), .A1(n5991), .B0(n6672), .Y(n6674));
  NOR2X1  g5551(.A(n6674), .B(n6673), .Y(n6675));
  OAI21X1 g5552(.A0(n6665), .A1(n6045), .B0(n6675), .Y(n6676));
  NOR2X1  g5553(.A(n6665), .B(n6018), .Y(n6677));
  AOI21X1 g5554(.A0(n6035), .A1(n5897), .B0(n6665), .Y(n6678));
  AOI22X1 g5555(.A0(n5957), .A1(P2_REG0_REG_18__SCAN_IN), .B0(P2_REG2_REG_18__SCAN_IN), .B1(n5958), .Y(n6679));
  INVX1   g5556(.A(P2_REG3_REG_18__SCAN_IN), .Y(n6680));
  XOR2X1  g5557(.A(n6641), .B(n6680), .Y(n6681));
  INVX1   g5558(.A(n6681), .Y(n6682));
  AOI22X1 g5559(.A0(n5962), .A1(n6682), .B0(n5961), .B1(P2_REG1_REG_18__SCAN_IN), .Y(n6683));
  NAND2X1 g5560(.A(n6683), .B(n6679), .Y(n6684));
  AOI22X1 g5561(.A0(n6658), .A1(n6008), .B0(n5917), .B1(n6684), .Y(n6685));
  OAI21X1 g5562(.A0(n6672), .A1(n6007), .B0(n6685), .Y(n6686));
  NOR4X1  g5563(.A(n6678), .B(n6677), .C(n6676), .D(n6686), .Y(n6687));
  NAND2X1 g5564(.A(n5970), .B(P2_REG0_REG_17__SCAN_IN), .Y(n6688));
  OAI21X1 g5565(.A0(n6687), .A1(n5970), .B0(n6688), .Y(P2_U3441));
  NOR2X1  g5566(.A(n6657), .B(n6651), .Y(n6690));
  INVX1   g5567(.A(n6645), .Y(n6691));
  AOI21X1 g5568(.A0(n6657), .A1(n6651), .B0(n6691), .Y(n6692));
  NOR2X1  g5569(.A(n6692), .B(n6690), .Y(n6693));
  OAI21X1 g5570(.A0(n6659), .A1(n6610), .B0(n6693), .Y(n6694));
  NOR2X1  g5571(.A(P2_IR_REG_31__SCAN_IN), .B(n5606), .Y(n6695));
  AOI21X1 g5572(.A0(n5611), .A1(P2_IR_REG_31__SCAN_IN), .B0(n6695), .Y(n6696));
  INVX1   g5573(.A(n6696), .Y(n6697));
  NOR2X1  g5574(.A(n5870), .B(n5605), .Y(n6698));
  AOI21X1 g5575(.A0(n6697), .A1(n5870), .B0(n6698), .Y(n6699));
  XOR2X1  g5576(.A(n6699), .B(n6684), .Y(n6700));
  NOR2X1  g5577(.A(n6694), .B(n6700), .Y(n6701));
  INVX1   g5578(.A(n6684), .Y(n6702));
  XOR2X1  g5579(.A(n6699), .B(n6702), .Y(n6703));
  AOI21X1 g5580(.A0(n6700), .A1(n6694), .B0(n6701), .Y(n6705));
  NOR2X1  g5581(.A(n6705), .B(n6045), .Y(n6706));
  NOR2X1  g5582(.A(n6658), .B(n6691), .Y(n6708));
  INVX1   g5583(.A(n6667), .Y(n6709));
  AOI22X1 g5584(.A0(n6709), .A1(n6669), .B0(n6658), .B1(n6691), .Y(n6710));
  NOR2X1  g5585(.A(n6710), .B(n6708), .Y(n6711));
  XOR2X1  g5586(.A(n6711), .B(n6703), .Y(n6712));
  AOI22X1 g5587(.A0(n6645), .A1(n5952), .B0(n5908), .B1(n6712), .Y(n6713));
  OAI21X1 g5588(.A0(n5909), .A1(n5902), .B0(n6712), .Y(n6714));
  NAND2X1 g5589(.A(n6714), .B(n6713), .Y(n6715));
  NOR2X1  g5590(.A(n6705), .B(n6018), .Y(n6716));
  AOI21X1 g5591(.A0(n6035), .A1(n5897), .B0(n6705), .Y(n6717));
  NOR4X1  g5592(.A(n6716), .B(n6715), .C(n6706), .D(n6717), .Y(n6718));
  INVX1   g5593(.A(n6718), .Y(n6719));
  NAND2X1 g5594(.A(n6712), .B(n5913), .Y(n6720));
  INVX1   g5595(.A(n6699), .Y(n6721));
  AOI22X1 g5596(.A0(n5957), .A1(P2_REG0_REG_19__SCAN_IN), .B0(P2_REG2_REG_19__SCAN_IN), .B1(n5958), .Y(n6722));
  INVX1   g5597(.A(P2_REG3_REG_19__SCAN_IN), .Y(n6723));
  NOR4X1  g5598(.A(P2_REG3_REG_18__SCAN_IN), .B(P2_REG3_REG_17__SCAN_IN), .C(P2_REG3_REG_16__SCAN_IN), .D(n6639), .Y(n6724));
  NOR3X1  g5599(.A(n6642), .B(P2_REG3_REG_18__SCAN_IN), .C(P2_REG3_REG_19__SCAN_IN), .Y(n6725));
  INVX1   g5600(.A(n6725), .Y(n6726));
  OAI21X1 g5601(.A0(n6724), .A1(n6723), .B0(n6726), .Y(n6727));
  AOI22X1 g5602(.A0(n5962), .A1(n6727), .B0(n5961), .B1(P2_REG1_REG_19__SCAN_IN), .Y(n6728));
  NAND2X1 g5603(.A(n6728), .B(n6722), .Y(n6729));
  AOI22X1 g5604(.A0(n6721), .A1(n6008), .B0(n5917), .B1(n6729), .Y(n6730));
  NAND2X1 g5605(.A(n6730), .B(n6720), .Y(n6731));
  NOR2X1  g5606(.A(n6731), .B(n6719), .Y(n6732));
  NAND2X1 g5607(.A(n5970), .B(P2_REG0_REG_18__SCAN_IN), .Y(n6733));
  OAI21X1 g5608(.A0(n6732), .A1(n5970), .B0(n6733), .Y(P2_U3444));
  INVX1   g5609(.A(n6729), .Y(n6735));
  NAND2X1 g5610(.A(n5870), .B(n5860), .Y(n6736));
  OAI21X1 g5611(.A0(n5870), .A1(n5616), .B0(n6736), .Y(n6737));
  NOR2X1  g5612(.A(n6721), .B(n6684), .Y(n6740));
  INVX1   g5613(.A(n6740), .Y(n6741));
  NOR2X1  g5614(.A(n6699), .B(n6702), .Y(n6742));
  AOI21X1 g5615(.A0(n6741), .A1(n6694), .B0(n6742), .Y(n6743));
  XOR2X1  g5616(.A(n6737), .B(n6729), .Y(n6744));
  NOR2X1  g5617(.A(n6744), .B(n6743), .Y(n6745));
  AOI21X1 g5618(.A0(n6743), .A1(n6744), .B0(n6745), .Y(n6746));
  NOR2X1  g5619(.A(n6746), .B(n6045), .Y(n6747));
  NOR2X1  g5620(.A(n6721), .B(n6702), .Y(n6748));
  INVX1   g5621(.A(n6748), .Y(n6749));
  OAI21X1 g5622(.A0(n6710), .A1(n6708), .B0(n6684), .Y(n6750));
  OAI21X1 g5623(.A0(n6710), .A1(n6708), .B0(n6699), .Y(n6751));
  NAND3X1 g5624(.A(n6751), .B(n6750), .C(n6749), .Y(n6752));
  XOR2X1  g5625(.A(n6752), .B(n6744), .Y(n6753));
  INVX1   g5626(.A(n6753), .Y(n6754));
  AOI22X1 g5627(.A0(n6684), .A1(n5952), .B0(n5908), .B1(n6754), .Y(n6755));
  OAI21X1 g5628(.A0(n5909), .A1(n5902), .B0(n6754), .Y(n6756));
  NAND2X1 g5629(.A(n6756), .B(n6755), .Y(n6757));
  NOR2X1  g5630(.A(n6746), .B(n6018), .Y(n6758));
  AOI21X1 g5631(.A0(n6035), .A1(n5897), .B0(n6746), .Y(n6759));
  NOR4X1  g5632(.A(n6758), .B(n6757), .C(n6747), .D(n6759), .Y(n6760));
  INVX1   g5633(.A(n6760), .Y(n6761));
  AOI22X1 g5634(.A0(n5957), .A1(P2_REG0_REG_20__SCAN_IN), .B0(P2_REG2_REG_20__SCAN_IN), .B1(n5958), .Y(n6762));
  INVX1   g5635(.A(P2_REG3_REG_20__SCAN_IN), .Y(n6763));
  XOR2X1  g5636(.A(n6725), .B(n6763), .Y(n6764));
  INVX1   g5637(.A(n6764), .Y(n6765));
  AOI22X1 g5638(.A0(n5962), .A1(n6765), .B0(n5961), .B1(P2_REG1_REG_20__SCAN_IN), .Y(n6766));
  NAND2X1 g5639(.A(n6766), .B(n6762), .Y(n6767));
  AOI22X1 g5640(.A0(n6737), .A1(n6008), .B0(n5917), .B1(n6767), .Y(n6768));
  OAI21X1 g5641(.A0(n6753), .A1(n6007), .B0(n6768), .Y(n6769));
  NOR2X1  g5642(.A(n6769), .B(n6761), .Y(n6770));
  NAND2X1 g5643(.A(n5970), .B(P2_REG0_REG_19__SCAN_IN), .Y(n6771));
  OAI21X1 g5644(.A0(n6770), .A1(n5970), .B0(n6771), .Y(P2_U3446));
  INVX1   g5645(.A(n6767), .Y(n6773));
  NOR2X1  g5646(.A(n5870), .B(n5623), .Y(n6774));
  XOR2X1  g5647(.A(n6774), .B(n6773), .Y(n6775));
  NOR2X1  g5648(.A(n6737), .B(n6735), .Y(n6776));
  NAND2X1 g5649(.A(n6737), .B(n6735), .Y(n6777));
  AOI21X1 g5650(.A0(n6752), .A1(n6777), .B0(n6776), .Y(n6778));
  XOR2X1  g5651(.A(n6778), .B(n6775), .Y(n6779));
  INVX1   g5652(.A(n6779), .Y(n6780));
  AOI22X1 g5653(.A0(n6729), .A1(n5952), .B0(n5908), .B1(n6780), .Y(n6781));
  OAI21X1 g5654(.A0(n5909), .A1(n5902), .B0(n6780), .Y(n6782));
  INVX1   g5655(.A(n6743), .Y(n6783));
  NAND2X1 g5656(.A(n6737), .B(n6729), .Y(n6784));
  INVX1   g5657(.A(n6784), .Y(n6785));
  OAI22X1 g5658(.A0(n6767), .A1(n6774), .B0(n6737), .B1(n6729), .Y(n6786));
  AOI21X1 g5659(.A0(n6774), .A1(n6767), .B0(n6786), .Y(n6787));
  OAI21X1 g5660(.A0(n6785), .A1(n6783), .B0(n6787), .Y(n6788));
  NOR2X1  g5661(.A(n6737), .B(n6729), .Y(n6789));
  NOR2X1  g5662(.A(n6774), .B(n6773), .Y(n6790));
  NOR3X1  g5663(.A(n6767), .B(n5870), .C(n5623), .Y(n6791));
  NOR3X1  g5664(.A(n6791), .B(n6790), .C(n6785), .Y(n6792));
  OAI21X1 g5665(.A0(n6789), .A1(n6743), .B0(n6792), .Y(n6793));
  NAND2X1 g5666(.A(n6793), .B(n6788), .Y(n6794));
  INVX1   g5667(.A(n6794), .Y(n6795));
  OAI21X1 g5668(.A0(n5905), .A1(n5904), .B0(n6795), .Y(n6796));
  OAI21X1 g5669(.A0(n5901), .A1(n5896), .B0(n6795), .Y(n6797));
  NAND4X1 g5670(.A(n6796), .B(n6782), .C(n6781), .D(n6797), .Y(n6798));
  AOI22X1 g5671(.A0(n5957), .A1(P2_REG0_REG_21__SCAN_IN), .B0(P2_REG2_REG_21__SCAN_IN), .B1(n5958), .Y(n6799));
  NOR4X1  g5672(.A(P2_REG3_REG_18__SCAN_IN), .B(P2_REG3_REG_20__SCAN_IN), .C(P2_REG3_REG_19__SCAN_IN), .D(n6642), .Y(n6800));
  INVX1   g5673(.A(n6800), .Y(n6801));
  NOR3X1  g5674(.A(n6726), .B(P2_REG3_REG_20__SCAN_IN), .C(P2_REG3_REG_21__SCAN_IN), .Y(n6802));
  AOI21X1 g5675(.A0(n6801), .A1(P2_REG3_REG_21__SCAN_IN), .B0(n6802), .Y(n6803));
  INVX1   g5676(.A(n6803), .Y(n6804));
  AOI22X1 g5677(.A0(n5962), .A1(n6804), .B0(n5961), .B1(P2_REG1_REG_21__SCAN_IN), .Y(n6805));
  NAND2X1 g5678(.A(n6805), .B(n6799), .Y(n6806));
  AOI22X1 g5679(.A0(n6774), .A1(n6008), .B0(n5917), .B1(n6806), .Y(n6807));
  OAI21X1 g5680(.A0(n6779), .A1(n6007), .B0(n6807), .Y(n6808));
  NOR2X1  g5681(.A(n6808), .B(n6798), .Y(n6809));
  NAND2X1 g5682(.A(n5970), .B(P2_REG0_REG_20__SCAN_IN), .Y(n6810));
  OAI21X1 g5683(.A0(n6809), .A1(n5970), .B0(n6810), .Y(P2_U3447));
  INVX1   g5684(.A(n6790), .Y(n6812));
  OAI21X1 g5685(.A0(n6778), .A1(n6791), .B0(n6812), .Y(n6813));
  INVX1   g5686(.A(n6806), .Y(n6814));
  NOR2X1  g5687(.A(n5870), .B(n5635), .Y(n6815));
  XOR2X1  g5688(.A(n6815), .B(n6814), .Y(n6816));
  XOR2X1  g5689(.A(n8528), .B(n6813), .Y(n6818));
  AOI21X1 g5690(.A0(n6003), .A1(n5991), .B0(n6818), .Y(n6819));
  INVX1   g5691(.A(n6737), .Y(n6820));
  NAND2X1 g5692(.A(n1606), .B(n1152), .Y(n6821));
  NAND2X1 g5693(.A(n5621), .B(n6821), .Y(n6822));
  INVX1   g5694(.A(n5870), .Y(n6823));
  NAND2X1 g5695(.A(n6823), .B(n6822), .Y(n6824));
  AOI22X1 g5696(.A0(n6773), .A1(n6824), .B0(n6820), .B1(n6735), .Y(n6825));
  OAI21X1 g5697(.A0(n5870), .A1(n5623), .B0(n6784), .Y(n6826));
  OAI21X1 g5698(.A0(n6824), .A1(n6784), .B0(n6773), .Y(n6827));
  AOI22X1 g5699(.A0(n6826), .A1(n6827), .B0(n6825), .B1(n6783), .Y(n6828));
  AOI21X1 g5700(.A0(n6827), .A1(n6826), .B0(n8528), .Y(n6829));
  OAI21X1 g5701(.A0(n6786), .A1(n6743), .B0(n6829), .Y(n6830));
  OAI21X1 g5702(.A0(n6828), .A1(n6816), .B0(n6830), .Y(n6831));
  OAI22X1 g5703(.A0(n6818), .A1(n6002), .B0(n6018), .B1(n6831), .Y(n6832));
  OAI22X1 g5704(.A0(n6773), .A1(n6046), .B0(n6045), .B1(n6831), .Y(n6833));
  AOI21X1 g5705(.A0(n6035), .A1(n5897), .B0(n6831), .Y(n6834));
  NOR4X1  g5706(.A(n6833), .B(n6832), .C(n6819), .D(n6834), .Y(n6835));
  INVX1   g5707(.A(n6835), .Y(n6836));
  AOI22X1 g5708(.A0(n5957), .A1(P2_REG0_REG_22__SCAN_IN), .B0(P2_REG2_REG_22__SCAN_IN), .B1(n5958), .Y(n6837));
  INVX1   g5709(.A(P2_REG3_REG_22__SCAN_IN), .Y(n6838));
  XOR2X1  g5710(.A(n6802), .B(n6838), .Y(n6839));
  INVX1   g5711(.A(n6839), .Y(n6840));
  AOI22X1 g5712(.A0(n5962), .A1(n6840), .B0(n5961), .B1(P2_REG1_REG_22__SCAN_IN), .Y(n6841));
  NAND2X1 g5713(.A(n6841), .B(n6837), .Y(n6842));
  AOI22X1 g5714(.A0(n6815), .A1(n6008), .B0(n5917), .B1(n6842), .Y(n6843));
  OAI21X1 g5715(.A0(n6818), .A1(n6007), .B0(n6843), .Y(n6844));
  NOR2X1  g5716(.A(n6844), .B(n6836), .Y(n6845));
  NAND2X1 g5717(.A(n5970), .B(P2_REG0_REG_21__SCAN_IN), .Y(n6846));
  OAI21X1 g5718(.A0(n6845), .A1(n5970), .B0(n6846), .Y(P2_U3448));
  INVX1   g5719(.A(n6842), .Y(n6848));
  NOR2X1  g5720(.A(n5870), .B(n5642), .Y(n6849));
  XOR2X1  g5721(.A(n6849), .B(n6848), .Y(n6850));
  NOR2X1  g5722(.A(n6815), .B(n6814), .Y(n6851));
  NOR3X1  g5723(.A(n6806), .B(n5870), .C(n5635), .Y(n6852));
  INVX1   g5724(.A(n6852), .Y(n6853));
  AOI21X1 g5725(.A0(n6853), .A1(n6813), .B0(n6851), .Y(n6854));
  XOR2X1  g5726(.A(n6854), .B(n6850), .Y(n6855));
  NOR2X1  g5727(.A(n6855), .B(n5991), .Y(n6856));
  INVX1   g5728(.A(n6850), .Y(n6857));
  NOR2X1  g5729(.A(n6815), .B(n6806), .Y(n6858));
  NOR3X1  g5730(.A(n6858), .B(n6786), .C(n6740), .Y(n6859));
  AOI22X1 g5731(.A0(n6826), .A1(n6827), .B0(n6825), .B1(n6742), .Y(n6860));
  NAND2X1 g5732(.A(n6815), .B(n6806), .Y(n6861));
  OAI21X1 g5733(.A0(n6860), .A1(n6858), .B0(n6861), .Y(n6862));
  AOI21X1 g5734(.A0(n6859), .A1(n6694), .B0(n6862), .Y(n6863));
  XOR2X1  g5735(.A(n6863), .B(n6857), .Y(n6864));
  OAI22X1 g5736(.A0(n6814), .A1(n6046), .B0(n6045), .B1(n6864), .Y(n6865));
  NOR2X1  g5737(.A(n6864), .B(n6018), .Y(n6866));
  AOI21X1 g5738(.A0(n6035), .A1(n5897), .B0(n6864), .Y(n6867));
  NOR4X1  g5739(.A(n6866), .B(n6865), .C(n6856), .D(n6867), .Y(n6868));
  INVX1   g5740(.A(n6855), .Y(n6869));
  OAI21X1 g5741(.A0(n5909), .A1(n5908), .B0(n6869), .Y(n6870));
  NAND2X1 g5742(.A(n6870), .B(n6868), .Y(n6871));
  AOI22X1 g5743(.A0(n5957), .A1(P2_REG0_REG_23__SCAN_IN), .B0(P2_REG2_REG_23__SCAN_IN), .B1(n5958), .Y(n6872));
  INVX1   g5744(.A(P2_REG3_REG_23__SCAN_IN), .Y(n6873));
  NOR4X1  g5745(.A(P2_REG3_REG_22__SCAN_IN), .B(P2_REG3_REG_20__SCAN_IN), .C(P2_REG3_REG_21__SCAN_IN), .D(n6726), .Y(n6874));
  NAND3X1 g5746(.A(n6802), .B(n6838), .C(n6873), .Y(n6875));
  OAI21X1 g5747(.A0(n6874), .A1(n6873), .B0(n6875), .Y(n6876));
  AOI22X1 g5748(.A0(n5962), .A1(n6876), .B0(n5961), .B1(P2_REG1_REG_23__SCAN_IN), .Y(n6877));
  NAND2X1 g5749(.A(n6877), .B(n6872), .Y(n6878));
  AOI22X1 g5750(.A0(n6849), .A1(n6008), .B0(n5917), .B1(n6878), .Y(n6879));
  OAI21X1 g5751(.A0(n6855), .A1(n6007), .B0(n6879), .Y(n6880));
  NOR2X1  g5752(.A(n6880), .B(n6871), .Y(n6881));
  NAND2X1 g5753(.A(n5970), .B(P2_REG0_REG_22__SCAN_IN), .Y(n6882));
  OAI21X1 g5754(.A0(n6881), .A1(n5970), .B0(n6882), .Y(P2_U3449));
  OAI21X1 g5755(.A0(n6849), .A1(n6848), .B0(n6854), .Y(n6884));
  NOR3X1  g5756(.A(n6842), .B(n5870), .C(n5642), .Y(n6885));
  NAND2X1 g5757(.A(n6823), .B(n5650), .Y(n6886));
  XOR2X1  g5758(.A(n6886), .B(n6878), .Y(n6887));
  NOR2X1  g5759(.A(n6887), .B(n6885), .Y(n6888));
  NAND2X1 g5760(.A(n6888), .B(n6884), .Y(n6889));
  INVX1   g5761(.A(n6878), .Y(n6890));
  NAND3X1 g5762(.A(n6890), .B(n6823), .C(n5650), .Y(n6891));
  INVX1   g5763(.A(n6891), .Y(n6892));
  INVX1   g5764(.A(n6849), .Y(n6893));
  AOI22X1 g5765(.A0(n6878), .A1(n6886), .B0(n6893), .B1(n6842), .Y(n6894));
  INVX1   g5766(.A(n6894), .Y(n6895));
  NOR2X1  g5767(.A(n6895), .B(n6892), .Y(n6896));
  OAI21X1 g5768(.A0(n6854), .A1(n6885), .B0(n6896), .Y(n6897));
  AOI21X1 g5769(.A0(n6897), .A1(n6889), .B0(n5991), .Y(n6898));
  NAND2X1 g5770(.A(n6849), .B(n6842), .Y(n6899));
  NOR2X1  g5771(.A(n6849), .B(n6842), .Y(n6900));
  OAI21X1 g5772(.A0(n6900), .A1(n6863), .B0(n6899), .Y(n6901));
  XOR2X1  g5773(.A(n6901), .B(n6887), .Y(n6902));
  INVX1   g5774(.A(n6902), .Y(n6903));
  AOI22X1 g5775(.A0(n6842), .A1(n5952), .B0(n5905), .B1(n6903), .Y(n6904));
  AOI21X1 g5776(.A0(n6035), .A1(n5897), .B0(n6902), .Y(n6905));
  AOI21X1 g5777(.A0(n6903), .A1(n5901), .B0(n6905), .Y(n6906));
  NAND2X1 g5778(.A(n6906), .B(n6904), .Y(n6907));
  AOI22X1 g5779(.A0(n6889), .A1(n6897), .B0(n6003), .B1(n6002), .Y(n6908));
  INVX1   g5780(.A(n6897), .Y(n6909));
  AOI21X1 g5781(.A0(n6888), .A1(n6884), .B0(n6909), .Y(n6910));
  INVX1   g5782(.A(n6886), .Y(n6911));
  AOI22X1 g5783(.A0(n5957), .A1(P2_REG0_REG_24__SCAN_IN), .B0(P2_REG2_REG_24__SCAN_IN), .B1(n5958), .Y(n6912));
  XOR2X1  g5784(.A(n6875), .B(P2_REG3_REG_24__SCAN_IN), .Y(n6913));
  INVX1   g5785(.A(n6913), .Y(n6914));
  AOI22X1 g5786(.A0(n5962), .A1(n6914), .B0(n5961), .B1(P2_REG1_REG_24__SCAN_IN), .Y(n6915));
  NAND2X1 g5787(.A(n6915), .B(n6912), .Y(n6916));
  AOI22X1 g5788(.A0(n6911), .A1(n6008), .B0(n5917), .B1(n6916), .Y(n6917));
  OAI21X1 g5789(.A0(n6910), .A1(n6007), .B0(n6917), .Y(n6918));
  NOR4X1  g5790(.A(n6908), .B(n6907), .C(n6898), .D(n6918), .Y(n6919));
  NAND2X1 g5791(.A(n5970), .B(P2_REG0_REG_23__SCAN_IN), .Y(n6920));
  OAI21X1 g5792(.A0(n6919), .A1(n5970), .B0(n6920), .Y(P2_U3450));
  NOR2X1  g5793(.A(n6886), .B(n6890), .Y(n6922));
  NAND2X1 g5794(.A(n6886), .B(n6890), .Y(n6923));
  AOI21X1 g5795(.A0(n6923), .A1(n6901), .B0(n6922), .Y(n6924));
  NAND2X1 g5796(.A(n6823), .B(n5658), .Y(n6925));
  XOR2X1  g5797(.A(n6925), .B(n6916), .Y(n6926));
  NAND2X1 g5798(.A(n6924), .B(n6930), .Y(n6928));
  INVX1   g5799(.A(n6916), .Y(n6929));
  XOR2X1  g5800(.A(n6925), .B(n6929), .Y(n6930));
  OAI21X1 g5801(.A0(n6930), .A1(n6924), .B0(n6928), .Y(n6931));
  NAND2X1 g5802(.A(n6931), .B(n5901), .Y(n6932));
  OAI21X1 g5803(.A0(n5904), .A1(n5896), .B0(n6931), .Y(n6933));
  NAND2X1 g5804(.A(n6933), .B(n6932), .Y(n6934));
  INVX1   g5805(.A(n6885), .Y(n6935));
  NAND3X1 g5806(.A(n6891), .B(n6935), .C(n6851), .Y(n6936));
  AOI21X1 g5807(.A0(n6936), .A1(n6894), .B0(n6892), .Y(n6937));
  NOR3X1  g5808(.A(n6892), .B(n6885), .C(n6852), .Y(n6938));
  AOI21X1 g5809(.A0(n6938), .A1(n6813), .B0(n6937), .Y(n6939));
  XOR2X1  g5810(.A(n6939), .B(n6926), .Y(n6940));
  AOI22X1 g5811(.A0(n6878), .A1(n5952), .B0(n5905), .B1(n6931), .Y(n6941));
  OAI21X1 g5812(.A0(n6940), .A1(n5991), .B0(n6941), .Y(n6942));
  INVX1   g5813(.A(n6940), .Y(n6943));
  OAI21X1 g5814(.A0(n5909), .A1(n5908), .B0(n6943), .Y(n6944));
  INVX1   g5815(.A(n6944), .Y(n6945));
  INVX1   g5816(.A(n6925), .Y(n6946));
  AOI22X1 g5817(.A0(n5957), .A1(P2_REG0_REG_25__SCAN_IN), .B0(P2_REG2_REG_25__SCAN_IN), .B1(n5958), .Y(n6947));
  NOR3X1  g5818(.A(n6875), .B(P2_REG3_REG_24__SCAN_IN), .C(P2_REG3_REG_25__SCAN_IN), .Y(n6948));
  INVX1   g5819(.A(n6948), .Y(n6949));
  OAI21X1 g5820(.A0(n6875), .A1(P2_REG3_REG_24__SCAN_IN), .B0(P2_REG3_REG_25__SCAN_IN), .Y(n6950));
  NAND2X1 g5821(.A(n6950), .B(n6949), .Y(n6951));
  AOI22X1 g5822(.A0(n5962), .A1(n6951), .B0(n5961), .B1(P2_REG1_REG_25__SCAN_IN), .Y(n6952));
  NAND2X1 g5823(.A(n6952), .B(n6947), .Y(n6953));
  AOI22X1 g5824(.A0(n6946), .A1(n6008), .B0(n5917), .B1(n6953), .Y(n6954));
  OAI21X1 g5825(.A0(n6940), .A1(n6007), .B0(n6954), .Y(n6955));
  NOR4X1  g5826(.A(n6945), .B(n6942), .C(n6934), .D(n6955), .Y(n6956));
  NAND2X1 g5827(.A(n5970), .B(P2_REG0_REG_24__SCAN_IN), .Y(n6957));
  OAI21X1 g5828(.A0(n6956), .A1(n5970), .B0(n6957), .Y(P2_U3451));
  INVX1   g5829(.A(n6953), .Y(n6959));
  NOR2X1  g5830(.A(n5870), .B(n5669), .Y(n6960));
  XOR2X1  g5831(.A(n6960), .B(n6959), .Y(n6961));
  NOR2X1  g5832(.A(n6925), .B(n6929), .Y(n6962));
  AOI21X1 g5833(.A0(n6925), .A1(n6929), .B0(n6924), .Y(n6963));
  NOR2X1  g5834(.A(n6963), .B(n6962), .Y(n6964));
  INVX1   g5835(.A(n6964), .Y(n6965));
  NOR2X1  g5836(.A(n6960), .B(n6953), .Y(n6966));
  NOR3X1  g5837(.A(n6959), .B(n5870), .C(n5669), .Y(n6967));
  OAI22X1 g5838(.A0(n6966), .A1(n6967), .B0(n6963), .B1(n6962), .Y(n6968));
  OAI21X1 g5839(.A0(n6965), .A1(n6961), .B0(n6968), .Y(n6969));
  NAND2X1 g5840(.A(n6969), .B(n5901), .Y(n6970));
  OAI21X1 g5841(.A0(n5904), .A1(n5896), .B0(n6969), .Y(n6971));
  NAND2X1 g5842(.A(n6971), .B(n6970), .Y(n6972));
  NAND2X1 g5843(.A(n6925), .B(n6916), .Y(n6973));
  NOR2X1  g5844(.A(n6925), .B(n6916), .Y(n6974));
  OAI21X1 g5845(.A0(n6939), .A1(n6974), .B0(n6973), .Y(n6975));
  XOR2X1  g5846(.A(n6975), .B(n6961), .Y(n6976));
  INVX1   g5847(.A(n6976), .Y(n6977));
  AOI22X1 g5848(.A0(n6916), .A1(n5952), .B0(n5905), .B1(n6969), .Y(n6978));
  OAI21X1 g5849(.A0(n6977), .A1(n5991), .B0(n6978), .Y(n6979));
  OAI21X1 g5850(.A0(n5909), .A1(n5908), .B0(n6976), .Y(n6980));
  INVX1   g5851(.A(n6980), .Y(n6981));
  AOI22X1 g5852(.A0(n5957), .A1(P2_REG0_REG_26__SCAN_IN), .B0(P2_REG2_REG_26__SCAN_IN), .B1(n5958), .Y(n6982));
  INVX1   g5853(.A(P2_REG3_REG_26__SCAN_IN), .Y(n6983));
  XOR2X1  g5854(.A(n6948), .B(n6983), .Y(n6984));
  INVX1   g5855(.A(n6984), .Y(n6985));
  AOI22X1 g5856(.A0(n5962), .A1(n6985), .B0(n5961), .B1(P2_REG1_REG_26__SCAN_IN), .Y(n6986));
  NAND2X1 g5857(.A(n6986), .B(n6982), .Y(n6987));
  AOI22X1 g5858(.A0(n6960), .A1(n6008), .B0(n5917), .B1(n6987), .Y(n6988));
  OAI21X1 g5859(.A0(n6977), .A1(n6007), .B0(n6988), .Y(n6989));
  NOR4X1  g5860(.A(n6981), .B(n6979), .C(n6972), .D(n6989), .Y(n6990));
  NAND2X1 g5861(.A(n5970), .B(P2_REG0_REG_25__SCAN_IN), .Y(n6991));
  OAI21X1 g5862(.A0(n6990), .A1(n5970), .B0(n6991), .Y(P2_U3452));
  NOR3X1  g5863(.A(n6967), .B(n6963), .C(n6962), .Y(n6993));
  INVX1   g5864(.A(n6987), .Y(n6994));
  OAI21X1 g5865(.A0(n3271), .A1(n1145), .B0(n5675), .Y(n6995));
  NAND2X1 g5866(.A(n6823), .B(n6995), .Y(n6996));
  AOI21X1 g5867(.A0(n6996), .A1(n6994), .B0(n6966), .Y(n6997));
  INVX1   g5868(.A(n6997), .Y(n6998));
  NOR3X1  g5869(.A(n6994), .B(n5870), .C(n5677), .Y(n6999));
  NOR3X1  g5870(.A(n6999), .B(n6998), .C(n6993), .Y(n7000));
  OAI22X1 g5871(.A0(n6960), .A1(n6953), .B0(n6962), .B1(n6963), .Y(n7001));
  XOR2X1  g5872(.A(n6996), .B(n6994), .Y(n7002));
  NOR2X1  g5873(.A(n7002), .B(n6967), .Y(n7003));
  AOI21X1 g5874(.A0(n7003), .A1(n7001), .B0(n7000), .Y(n7004));
  NAND2X1 g5875(.A(n7004), .B(n5901), .Y(n7005));
  OAI21X1 g5876(.A0(n5904), .A1(n5896), .B0(n7004), .Y(n7006));
  NAND2X1 g5877(.A(n7006), .B(n7005), .Y(n7007));
  NAND2X1 g5878(.A(n6960), .B(n6959), .Y(n7008));
  XOR2X1  g5879(.A(n8505), .B(n7002), .Y(n7011));
  AOI22X1 g5880(.A0(n6953), .A1(n5952), .B0(n5905), .B1(n7004), .Y(n7012));
  OAI21X1 g5881(.A0(n7011), .A1(n5991), .B0(n7012), .Y(n7013));
  AOI21X1 g5882(.A0(n6003), .A1(n6002), .B0(n7011), .Y(n7014));
  INVX1   g5883(.A(n6996), .Y(n7015));
  AOI22X1 g5884(.A0(n5957), .A1(P2_REG0_REG_27__SCAN_IN), .B0(P2_REG2_REG_27__SCAN_IN), .B1(n5958), .Y(n7016));
  INVX1   g5885(.A(P2_REG3_REG_27__SCAN_IN), .Y(n7017));
  NOR4X1  g5886(.A(P2_REG3_REG_26__SCAN_IN), .B(P2_REG3_REG_24__SCAN_IN), .C(P2_REG3_REG_25__SCAN_IN), .D(n6875), .Y(n7018));
  NOR3X1  g5887(.A(n6949), .B(P2_REG3_REG_26__SCAN_IN), .C(P2_REG3_REG_27__SCAN_IN), .Y(n7019));
  INVX1   g5888(.A(n7019), .Y(n7020));
  OAI21X1 g5889(.A0(n7018), .A1(n7017), .B0(n7020), .Y(n7021));
  AOI22X1 g5890(.A0(n5962), .A1(n7021), .B0(n5961), .B1(P2_REG1_REG_27__SCAN_IN), .Y(n7022));
  NAND2X1 g5891(.A(n7022), .B(n7016), .Y(n7023));
  AOI22X1 g5892(.A0(n7015), .A1(n6008), .B0(n5917), .B1(n7023), .Y(n7024));
  OAI21X1 g5893(.A0(n7011), .A1(n6007), .B0(n7024), .Y(n7025));
  NOR4X1  g5894(.A(n7014), .B(n7013), .C(n7007), .D(n7025), .Y(n7026));
  NAND2X1 g5895(.A(n5970), .B(P2_REG0_REG_26__SCAN_IN), .Y(n7027));
  OAI21X1 g5896(.A0(n7026), .A1(n5970), .B0(n7027), .Y(P2_U3453));
  OAI21X1 g5897(.A0(n5870), .A1(n5677), .B0(n6987), .Y(n7029));
  NOR2X1  g5898(.A(n6960), .B(n6959), .Y(n7030));
  AOI21X1 g5899(.A0(n6975), .A1(n7008), .B0(n7030), .Y(n7031));
  NAND2X1 g5900(.A(n7031), .B(n7029), .Y(n7032));
  NOR3X1  g5901(.A(n6987), .B(n5870), .C(n5677), .Y(n7033));
  OAI21X1 g5902(.A0(n5687), .A1(n5685), .B0(n6823), .Y(n7034));
  XOR2X1  g5903(.A(n7034), .B(n7023), .Y(n7035));
  NOR2X1  g5904(.A(n7035), .B(n7033), .Y(n7036));
  NAND2X1 g5905(.A(n7036), .B(n7032), .Y(n7037));
  INVX1   g5906(.A(n7035), .Y(n7039));
  NOR2X1  g5907(.A(n7039), .B(n8426), .Y(n7040));
  OAI21X1 g5908(.A0(n7031), .A1(n7033), .B0(n7040), .Y(n7041));
  AOI22X1 g5909(.A0(n7037), .A1(n7041), .B0(n6003), .B1(n5991), .Y(n7042));
  NAND2X1 g5910(.A(n8505), .B(n8433), .Y(n7044));
  AOI22X1 g5911(.A0(n7044), .A1(n7040), .B0(n7036), .B1(n7032), .Y(n7045));
  INVX1   g5912(.A(n6960), .Y(n7046));
  OAI22X1 g5913(.A0(n6959), .A1(n7046), .B0(n6925), .B1(n6929), .Y(n7047));
  NAND2X1 g5914(.A(n7047), .B(n6997), .Y(n7048));
  AOI21X1 g5915(.A0(n6997), .A1(n6963), .B0(n6999), .Y(n7049));
  NAND2X1 g5916(.A(n7049), .B(n7048), .Y(n7050));
  XOR2X1  g5917(.A(n7050), .B(n7035), .Y(n7051));
  OAI22X1 g5918(.A0(n7045), .A1(n6002), .B0(n6018), .B1(n7051), .Y(n7052));
  NOR2X1  g5919(.A(n7052), .B(n7042), .Y(n7053));
  OAI22X1 g5920(.A0(n6994), .A1(n6046), .B0(n6045), .B1(n7051), .Y(n7054));
  AOI21X1 g5921(.A0(n6035), .A1(n5897), .B0(n7051), .Y(n7055));
  NOR2X1  g5922(.A(n7055), .B(n7054), .Y(n7056));
  NAND2X1 g5923(.A(n7056), .B(n7053), .Y(n7057));
  NOR2X1  g5924(.A(n5870), .B(n5688), .Y(n7058));
  AOI22X1 g5925(.A0(n5957), .A1(P2_REG0_REG_28__SCAN_IN), .B0(P2_REG2_REG_28__SCAN_IN), .B1(n5958), .Y(n7059));
  INVX1   g5926(.A(P2_REG3_REG_28__SCAN_IN), .Y(n7060));
  XOR2X1  g5927(.A(n7019), .B(n7060), .Y(n7061));
  INVX1   g5928(.A(n7061), .Y(n7062));
  AOI22X1 g5929(.A0(n5962), .A1(n7062), .B0(n5961), .B1(P2_REG1_REG_28__SCAN_IN), .Y(n7063));
  NAND2X1 g5930(.A(n7063), .B(n7059), .Y(n7064));
  AOI22X1 g5931(.A0(n7058), .A1(n6008), .B0(n5917), .B1(n7064), .Y(n7065));
  OAI21X1 g5932(.A0(n7045), .A1(n6007), .B0(n7065), .Y(n7066));
  NOR2X1  g5933(.A(n7066), .B(n7057), .Y(n7067));
  NAND2X1 g5934(.A(n5970), .B(P2_REG0_REG_27__SCAN_IN), .Y(n7068));
  OAI21X1 g5935(.A0(n7067), .A1(n5970), .B0(n7068), .Y(P2_U3454));
  OAI21X1 g5936(.A0(n3391), .A1(n1145), .B0(n5693), .Y(n7070));
  NAND2X1 g5937(.A(n6823), .B(n7070), .Y(n7071));
  XOR2X1  g5938(.A(n7071), .B(n7064), .Y(n7072));
  INVX1   g5939(.A(n7072), .Y(n7073));
  INVX1   g5940(.A(n7023), .Y(n7074));
  AOI21X1 g5941(.A0(n7074), .A1(n7029), .B0(n7058), .Y(n7075));
  AOI21X1 g5942(.A0(n7023), .A1(n8426), .B0(n7075), .Y(n7076));
  OAI22X1 g5943(.A0(n7023), .A1(n7034), .B0(n6996), .B1(n6987), .Y(n7077));
  OAI21X1 g5944(.A0(n7077), .A1(n7031), .B0(n7076), .Y(n7078));
  XOR2X1  g5945(.A(n7078), .B(n7073), .Y(n7079));
  AOI21X1 g5946(.A0(n6003), .A1(n5991), .B0(n7079), .Y(n7080));
  NAND2X1 g5947(.A(n7034), .B(n7074), .Y(n7081));
  NAND3X1 g5948(.A(n7081), .B(n7047), .C(n6997), .Y(n7082));
  NAND2X1 g5949(.A(n7058), .B(n7023), .Y(n7083));
  NAND2X1 g5950(.A(n7081), .B(n6999), .Y(n7084));
  NAND3X1 g5951(.A(n7081), .B(n6997), .C(n6963), .Y(n7085));
  NAND4X1 g5952(.A(n7084), .B(n7083), .C(n7082), .D(n7085), .Y(n7086));
  XOR2X1  g5953(.A(n7086), .B(n7072), .Y(n7087));
  OAI22X1 g5954(.A0(n7079), .A1(n6002), .B0(n6018), .B1(n7087), .Y(n7088));
  OAI22X1 g5955(.A0(n7074), .A1(n6046), .B0(n6045), .B1(n7087), .Y(n7089));
  AOI21X1 g5956(.A0(n6035), .A1(n5897), .B0(n7087), .Y(n7090));
  NOR4X1  g5957(.A(n7089), .B(n7088), .C(n7080), .D(n7090), .Y(n7091));
  INVX1   g5958(.A(n7091), .Y(n7092));
  NOR2X1  g5959(.A(n5870), .B(n5695), .Y(n7093));
  NOR4X1  g5960(.A(P2_REG3_REG_26__SCAN_IN), .B(P2_REG3_REG_28__SCAN_IN), .C(P2_REG3_REG_27__SCAN_IN), .D(n6949), .Y(n7094));
  INVX1   g5961(.A(n7094), .Y(n7095));
  NOR2X1  g5962(.A(n7095), .B(n6113), .Y(n7096));
  INVX1   g5963(.A(n7096), .Y(n7097));
  NAND3X1 g5964(.A(n5891), .B(n5882), .C(P2_REG1_REG_29__SCAN_IN), .Y(n7098));
  AOI22X1 g5965(.A0(n5957), .A1(P2_REG0_REG_29__SCAN_IN), .B0(P2_REG2_REG_29__SCAN_IN), .B1(n5958), .Y(n7099));
  NAND3X1 g5966(.A(n7099), .B(n7098), .C(n7097), .Y(n7100));
  AOI22X1 g5967(.A0(n7093), .A1(n6008), .B0(n5917), .B1(n7100), .Y(n7101));
  OAI21X1 g5968(.A0(n7079), .A1(n6007), .B0(n7101), .Y(n7102));
  NOR2X1  g5969(.A(n7102), .B(n7092), .Y(n7103));
  NAND2X1 g5970(.A(n5970), .B(P2_REG0_REG_28__SCAN_IN), .Y(n7104));
  OAI21X1 g5971(.A0(n7103), .A1(n5970), .B0(n7104), .Y(P2_U3455));
  INVX1   g5972(.A(n7100), .Y(n7106));
  NOR2X1  g5973(.A(n5870), .B(n5706), .Y(n7107));
  XOR2X1  g5974(.A(n7107), .B(n7106), .Y(n7108));
  AOI21X1 g5975(.A0(n7071), .A1(n7064), .B0(n7078), .Y(n7109));
  NAND2X1 g5976(.A(n7109), .B(n7108), .Y(n7110));
  INVX1   g5977(.A(n7064), .Y(n7111));
  NAND3X1 g5978(.A(n7111), .B(n6823), .C(n7070), .Y(n7112));
  OAI21X1 g5979(.A0(n3399), .A1(n1145), .B0(n5704), .Y(n7113));
  NAND2X1 g5980(.A(n6823), .B(n7113), .Y(n7114));
  XOR2X1  g5981(.A(n7114), .B(n7106), .Y(n7115));
  NAND3X1 g5982(.A(n7115), .B(n7078), .C(n7112), .Y(n7116));
  NOR2X1  g5983(.A(n7115), .B(n7112), .Y(n7117));
  NOR3X1  g5984(.A(n7108), .B(n7093), .C(n7111), .Y(n7118));
  NOR2X1  g5985(.A(n7118), .B(n7117), .Y(n7119));
  NAND3X1 g5986(.A(n7119), .B(n7116), .C(n7110), .Y(n7120));
  OAI21X1 g5987(.A0(n5909), .A1(n5908), .B0(n7120), .Y(n7121));
  NAND2X1 g5988(.A(n7086), .B(n7093), .Y(n7122));
  OAI21X1 g5989(.A0(n7086), .A1(n7093), .B0(n7064), .Y(n7123));
  NAND2X1 g5990(.A(n7123), .B(n7122), .Y(n7124));
  XOR2X1  g5991(.A(n7124), .B(n7115), .Y(n7125));
  OAI21X1 g5992(.A0(n5905), .A1(n5901), .B0(n7125), .Y(n7126));
  NAND2X1 g5993(.A(n7126), .B(n7121), .Y(n7127));
  NAND2X1 g5994(.A(n7125), .B(n5896), .Y(n7128));
  AOI22X1 g5995(.A0(n5957), .A1(P2_REG0_REG_30__SCAN_IN), .B0(P2_REG2_REG_30__SCAN_IN), .B1(n5958), .Y(n7129));
  NAND3X1 g5996(.A(n5891), .B(n5882), .C(P2_REG1_REG_30__SCAN_IN), .Y(n7130));
  NAND3X1 g5997(.A(n7130), .B(n7129), .C(n7097), .Y(n7131));
  NOR2X1  g5998(.A(n5844), .B(n5846), .Y(n7132));
  NOR3X1  g5999(.A(n5915), .B(n5914), .C(P2_B_REG_SCAN_IN), .Y(n7133));
  OAI21X1 g6000(.A0(n7133), .A1(n5870), .B0(n7132), .Y(n7134));
  INVX1   g6001(.A(n7134), .Y(n7135));
  AOI22X1 g6002(.A0(n7131), .A1(n7135), .B0(n7064), .B1(n5952), .Y(n7136));
  AOI22X1 g6003(.A0(n7120), .A1(n5902), .B0(n5904), .B1(n7125), .Y(n7137));
  NAND3X1 g6004(.A(n7137), .B(n7136), .C(n7128), .Y(n7138));
  NAND2X1 g6005(.A(n7120), .B(n5913), .Y(n7139));
  OAI21X1 g6006(.A0(n7114), .A1(n5926), .B0(n7139), .Y(n7140));
  NOR3X1  g6007(.A(n7140), .B(n7138), .C(n7127), .Y(n7141));
  NAND2X1 g6008(.A(n5970), .B(P2_REG0_REG_29__SCAN_IN), .Y(n7142));
  OAI21X1 g6009(.A0(n7141), .A1(n5970), .B0(n7142), .Y(P2_U3456));
  NAND3X1 g6010(.A(n5891), .B(n5882), .C(P2_REG1_REG_31__SCAN_IN), .Y(n7144));
  AOI22X1 g6011(.A0(n5957), .A1(P2_REG0_REG_31__SCAN_IN), .B0(P2_REG2_REG_31__SCAN_IN), .B1(n5958), .Y(n7145));
  NAND3X1 g6012(.A(n7145), .B(n7144), .C(n7097), .Y(n7146));
  INVX1   g6013(.A(n7146), .Y(n7147));
  NOR2X1  g6014(.A(n7147), .B(n7134), .Y(n7148));
  NOR2X1  g6015(.A(n5870), .B(n5714), .Y(n7149));
  AOI21X1 g6016(.A0(n7149), .A1(n6008), .B0(n7148), .Y(n7150));
  NAND2X1 g6017(.A(n5970), .B(P2_REG0_REG_30__SCAN_IN), .Y(n7151));
  OAI21X1 g6018(.A0(n7150), .A1(n5970), .B0(n7151), .Y(P2_U3457));
  AOI21X1 g6019(.A0(n5720), .A1(n5719), .B0(n5870), .Y(n7153));
  AOI21X1 g6020(.A0(n7153), .A1(n6008), .B0(n7148), .Y(n7154));
  NAND2X1 g6021(.A(n5970), .B(P2_REG0_REG_31__SCAN_IN), .Y(n7155));
  OAI21X1 g6022(.A0(n7154), .A1(n5970), .B0(n7155), .Y(P2_U3458));
  INVX1   g6023(.A(P2_REG1_REG_0__SCAN_IN), .Y(n7157));
  NAND2X1 g6024(.A(n5853), .B(n5850), .Y(n7158));
  OAI21X1 g6025(.A0(n5849), .A1(n5847), .B0(n5846), .Y(n7159));
  NAND3X1 g6026(.A(n7159), .B(n7158), .C(n5859), .Y(n7160));
  NAND4X1 g6027(.A(n5842), .B(n5838), .C(n5835), .D(n7160), .Y(n7161));
  NOR4X1  g6028(.A(n5857), .B(n5847), .C(n5846), .D(n5860), .Y(n7162));
  NOR2X1  g6029(.A(n7162), .B(n5861), .Y(n7163));
  NOR4X1  g6030(.A(n5842), .B(n5838), .C(n5836), .D(n7163), .Y(n7164));
  INVX1   g6031(.A(n7164), .Y(n7165));
  AOI21X1 g6032(.A0(n7165), .A1(n7161), .B0(n5815), .Y(n7166));
  NAND2X1 g6033(.A(n7166), .B(n5929), .Y(n7167));
  OAI21X1 g6034(.A0(n7166), .A1(n7157), .B0(n7167), .Y(P2_U3459));
  INVX1   g6035(.A(P2_REG1_REG_1__SCAN_IN), .Y(n7169));
  NAND2X1 g6036(.A(n7166), .B(n5968), .Y(n7170));
  OAI21X1 g6037(.A0(n7166), .A1(n7169), .B0(n7170), .Y(P2_U3460));
  INVX1   g6038(.A(n7166), .Y(n7172));
  NAND2X1 g6039(.A(n7172), .B(P2_REG1_REG_2__SCAN_IN), .Y(n7173));
  OAI21X1 g6040(.A0(n7172), .A1(n6015), .B0(n7173), .Y(P2_U3461));
  NAND2X1 g6041(.A(n7172), .B(P2_REG1_REG_3__SCAN_IN), .Y(n7175));
  OAI21X1 g6042(.A0(n7172), .A1(n6059), .B0(n7175), .Y(P2_U3462));
  NAND2X1 g6043(.A(n7172), .B(P2_REG1_REG_4__SCAN_IN), .Y(n7177));
  OAI21X1 g6044(.A0(n7172), .A1(n6101), .B0(n7177), .Y(P2_U3463));
  NAND2X1 g6045(.A(n7172), .B(P2_REG1_REG_5__SCAN_IN), .Y(n7179));
  OAI21X1 g6046(.A0(n7172), .A1(n6153), .B0(n7179), .Y(P2_U3464));
  NAND2X1 g6047(.A(n7172), .B(P2_REG1_REG_6__SCAN_IN), .Y(n7181));
  OAI21X1 g6048(.A0(n7172), .A1(n6203), .B0(n7181), .Y(P2_U3465));
  NAND2X1 g6049(.A(n7172), .B(P2_REG1_REG_7__SCAN_IN), .Y(n7183));
  OAI21X1 g6050(.A0(n7172), .A1(n6245), .B0(n7183), .Y(P2_U3466));
  NAND2X1 g6051(.A(n7172), .B(P2_REG1_REG_8__SCAN_IN), .Y(n7185));
  OAI21X1 g6052(.A0(n7172), .A1(n6287), .B0(n7185), .Y(P2_U3467));
  NAND2X1 g6053(.A(n7172), .B(P2_REG1_REG_9__SCAN_IN), .Y(n7187));
  OAI21X1 g6054(.A0(n7172), .A1(n6337), .B0(n7187), .Y(P2_U3468));
  NAND2X1 g6055(.A(n7172), .B(P2_REG1_REG_10__SCAN_IN), .Y(n7189));
  OAI21X1 g6056(.A0(n7172), .A1(n6382), .B0(n7189), .Y(P2_U3469));
  NAND2X1 g6057(.A(n7172), .B(P2_REG1_REG_11__SCAN_IN), .Y(n7191));
  OAI21X1 g6058(.A0(n7172), .A1(n6432), .B0(n7191), .Y(P2_U3470));
  NAND2X1 g6059(.A(n7172), .B(P2_REG1_REG_12__SCAN_IN), .Y(n7193));
  OAI21X1 g6060(.A0(n7172), .A1(n6473), .B0(n7193), .Y(P2_U3471));
  NAND2X1 g6061(.A(n7172), .B(P2_REG1_REG_13__SCAN_IN), .Y(n7195));
  OAI21X1 g6062(.A0(n7172), .A1(n6519), .B0(n7195), .Y(P2_U3472));
  NAND2X1 g6063(.A(n7172), .B(P2_REG1_REG_14__SCAN_IN), .Y(n7197));
  OAI21X1 g6064(.A0(n7172), .A1(n6562), .B0(n7197), .Y(P2_U3473));
  NAND2X1 g6065(.A(n7172), .B(P2_REG1_REG_15__SCAN_IN), .Y(n7199));
  OAI21X1 g6066(.A0(n7172), .A1(n6596), .B0(n7199), .Y(P2_U3474));
  NAND2X1 g6067(.A(n7172), .B(P2_REG1_REG_16__SCAN_IN), .Y(n7201));
  OAI21X1 g6068(.A0(n7172), .A1(n6648), .B0(n7201), .Y(P2_U3475));
  NAND2X1 g6069(.A(n7172), .B(P2_REG1_REG_17__SCAN_IN), .Y(n7203));
  OAI21X1 g6070(.A0(n7172), .A1(n6687), .B0(n7203), .Y(P2_U3476));
  NAND2X1 g6071(.A(n7172), .B(P2_REG1_REG_18__SCAN_IN), .Y(n7205));
  OAI21X1 g6072(.A0(n7172), .A1(n6732), .B0(n7205), .Y(P2_U3477));
  NAND2X1 g6073(.A(n7172), .B(P2_REG1_REG_19__SCAN_IN), .Y(n7207));
  OAI21X1 g6074(.A0(n7172), .A1(n6770), .B0(n7207), .Y(P2_U3478));
  NAND2X1 g6075(.A(n7172), .B(P2_REG1_REG_20__SCAN_IN), .Y(n7209));
  OAI21X1 g6076(.A0(n7172), .A1(n6809), .B0(n7209), .Y(P2_U3479));
  NAND2X1 g6077(.A(n7172), .B(P2_REG1_REG_21__SCAN_IN), .Y(n7211));
  OAI21X1 g6078(.A0(n7172), .A1(n6845), .B0(n7211), .Y(P2_U3480));
  NAND2X1 g6079(.A(n7172), .B(P2_REG1_REG_22__SCAN_IN), .Y(n7213));
  OAI21X1 g6080(.A0(n7172), .A1(n6881), .B0(n7213), .Y(P2_U3481));
  NAND2X1 g6081(.A(n7172), .B(P2_REG1_REG_23__SCAN_IN), .Y(n7215));
  OAI21X1 g6082(.A0(n7172), .A1(n6919), .B0(n7215), .Y(P2_U3482));
  NAND2X1 g6083(.A(n7172), .B(P2_REG1_REG_24__SCAN_IN), .Y(n7217));
  OAI21X1 g6084(.A0(n7172), .A1(n6956), .B0(n7217), .Y(P2_U3483));
  NAND2X1 g6085(.A(n7172), .B(P2_REG1_REG_25__SCAN_IN), .Y(n7219));
  OAI21X1 g6086(.A0(n7172), .A1(n6990), .B0(n7219), .Y(P2_U3484));
  NAND2X1 g6087(.A(n7172), .B(P2_REG1_REG_26__SCAN_IN), .Y(n7221));
  OAI21X1 g6088(.A0(n7172), .A1(n7026), .B0(n7221), .Y(P2_U3485));
  NAND2X1 g6089(.A(n7172), .B(P2_REG1_REG_27__SCAN_IN), .Y(n7223));
  OAI21X1 g6090(.A0(n7172), .A1(n7067), .B0(n7223), .Y(P2_U3486));
  NAND2X1 g6091(.A(n7172), .B(P2_REG1_REG_28__SCAN_IN), .Y(n7225));
  OAI21X1 g6092(.A0(n7172), .A1(n7103), .B0(n7225), .Y(P2_U3487));
  NAND2X1 g6093(.A(n7172), .B(P2_REG1_REG_29__SCAN_IN), .Y(n7227));
  OAI21X1 g6094(.A0(n7172), .A1(n7141), .B0(n7227), .Y(P2_U3488));
  NAND2X1 g6095(.A(n7172), .B(P2_REG1_REG_30__SCAN_IN), .Y(n7229));
  OAI21X1 g6096(.A0(n7172), .A1(n7150), .B0(n7229), .Y(P2_U3489));
  NAND2X1 g6097(.A(n7172), .B(P2_REG1_REG_31__SCAN_IN), .Y(n7231));
  OAI21X1 g6098(.A0(n7172), .A1(n7154), .B0(n7231), .Y(P2_U3490));
  NOR4X1  g6099(.A(n5849), .B(n5847), .C(n5907), .D(n5853), .Y(n7233));
  NOR2X1  g6100(.A(n5746), .B(n5726), .Y(n7234));
  AOI21X1 g6101(.A0(n5840), .A1(n5746), .B0(n7234), .Y(n7235));
  AOI21X1 g6102(.A0(n5860), .A1(n5844), .B0(n5846), .Y(n7236));
  OAI21X1 g6103(.A0(n5849), .A1(n5847), .B0(n7236), .Y(n7237));
  NAND4X1 g6104(.A(n7235), .B(n5839), .C(n5835), .D(n7237), .Y(n7238));
  INVX1   g6105(.A(n7238), .Y(n7239));
  NOR4X1  g6106(.A(n7235), .B(n5839), .C(n5836), .D(n7163), .Y(n7240));
  NAND3X1 g6107(.A(n7233), .B(n5744), .C(P2_REG3_REG_0__SCAN_IN), .Y(n7241));
  NOR3X1  g6108(.A(n7240), .B(n7239), .C(n7233), .Y(n7242));
  NOR2X1  g6109(.A(n7242), .B(n5815), .Y(n7243));
  INVX1   g6110(.A(P2_REG2_REG_0__SCAN_IN), .Y(n7244));
  NOR2X1  g6111(.A(n7243), .B(n7244), .Y(n7245));
  AOI21X1 g6112(.A0(n7243), .A1(n5911), .B0(n7245), .Y(n7246));
  NOR3X1  g6113(.A(n7242), .B(n5918), .C(n5815), .Y(n7247));
  NAND2X1 g6114(.A(n7247), .B(n5933), .Y(n7248));
  NOR3X1  g6115(.A(n5860), .B(n5847), .C(n5907), .Y(n7249));
  NOR4X1  g6116(.A(n5857), .B(n5847), .C(n5907), .D(n5853), .Y(n7250));
  NOR2X1  g6117(.A(n7250), .B(n7249), .Y(n7251));
  NOR3X1  g6118(.A(n7251), .B(n7242), .C(n5815), .Y(n7252));
  NOR2X1  g6119(.A(n5849), .B(n5844), .Y(n7253));
  INVX1   g6120(.A(n7253), .Y(n7254));
  NOR4X1  g6121(.A(n7242), .B(n5853), .C(n5815), .D(n7254), .Y(n7255));
  AOI22X1 g6122(.A0(n7252), .A1(n5878), .B0(n8531), .B1(n7255), .Y(n7256));
  NAND4X1 g6123(.A(n7248), .B(n7246), .C(n7241), .D(n7256), .Y(P2_U3233));
  NAND3X1 g6124(.A(n7233), .B(n5744), .C(P2_REG3_REG_1__SCAN_IN), .Y(n7258));
  INVX1   g6125(.A(P2_REG2_REG_1__SCAN_IN), .Y(n7259));
  NOR2X1  g6126(.A(n7243), .B(n7259), .Y(n7260));
  AOI21X1 g6127(.A0(n7243), .A1(n5955), .B0(n7260), .Y(n7261));
  INVX1   g6128(.A(n5965), .Y(n7262));
  NAND2X1 g6129(.A(n7247), .B(n7262), .Y(n7263));
  AOI22X1 g6130(.A0(n7252), .A1(n5945), .B0(n5942), .B1(n7255), .Y(n7264));
  NAND4X1 g6131(.A(n7263), .B(n7261), .C(n7258), .D(n7264), .Y(P2_U3232));
  NAND3X1 g6132(.A(n7233), .B(n5744), .C(P2_REG3_REG_2__SCAN_IN), .Y(n7266));
  INVX1   g6133(.A(P2_REG2_REG_2__SCAN_IN), .Y(n7267));
  NOR2X1  g6134(.A(n7243), .B(n7267), .Y(n7268));
  AOI21X1 g6135(.A0(n7243), .A1(n6006), .B0(n7268), .Y(n7269));
  INVX1   g6136(.A(n7252), .Y(n7270));
  INVX1   g6137(.A(n7255), .Y(n7271));
  OAI22X1 g6138(.A0(n7270), .A1(n5981), .B0(n5999), .B1(n7271), .Y(n7272));
  AOI21X1 g6139(.A0(n7247), .A1(n6012), .B0(n7272), .Y(n7273));
  NAND3X1 g6140(.A(n7273), .B(n7269), .C(n7266), .Y(P2_U3231));
  NAND3X1 g6141(.A(n7233), .B(n5744), .C(n6010), .Y(n7275));
  INVX1   g6142(.A(P2_REG2_REG_3__SCAN_IN), .Y(n7276));
  NOR2X1  g6143(.A(n7243), .B(n7276), .Y(n7277));
  AOI21X1 g6144(.A0(n7243), .A1(n6050), .B0(n7277), .Y(n7278));
  OAI22X1 g6145(.A0(n7270), .A1(n6024), .B0(n6051), .B1(n7271), .Y(n7279));
  AOI21X1 g6146(.A0(n7247), .A1(n6056), .B0(n7279), .Y(n7280));
  NAND3X1 g6147(.A(n7280), .B(n7278), .C(n7275), .Y(P2_U3230));
  INVX1   g6148(.A(n7243), .Y(n7282));
  INVX1   g6149(.A(n7233), .Y(n7283));
  NOR2X1  g6150(.A(n7283), .B(n5815), .Y(n7284));
  AOI22X1 g6151(.A0(n7282), .A1(P2_REG2_REG_4__SCAN_IN), .B0(n6054), .B1(n7284), .Y(n7285));
  AOI22X1 g6152(.A0(n7252), .A1(n6067), .B0(n6086), .B1(n7255), .Y(n7286));
  AOI22X1 g6153(.A0(n7243), .A1(n6091), .B0(n6098), .B1(n7247), .Y(n7287));
  NAND3X1 g6154(.A(n7287), .B(n7286), .C(n7285), .Y(P2_U3229));
  INVX1   g6155(.A(n7284), .Y(n7289));
  OAI22X1 g6156(.A0(n7243), .A1(n6107), .B0(n6095), .B1(n7289), .Y(n7290));
  NOR4X1  g6157(.A(n6156), .B(n5918), .C(n5815), .D(n7242), .Y(n7291));
  OAI22X1 g6158(.A0(n7270), .A1(n6120), .B0(n6137), .B1(n7271), .Y(n7292));
  NOR3X1  g6159(.A(n7292), .B(n7291), .C(n7290), .Y(n7293));
  OAI21X1 g6160(.A0(n7282), .A1(n6141), .B0(n7293), .Y(P2_U3228));
  NOR3X1  g6161(.A(n6194), .B(n6177), .C(n6175), .Y(n7295));
  INVX1   g6162(.A(P2_REG2_REG_6__SCAN_IN), .Y(n7296));
  OAI22X1 g6163(.A0(n7243), .A1(n7296), .B0(n6147), .B1(n7289), .Y(n7297));
  INVX1   g6164(.A(n7247), .Y(n7298));
  AOI22X1 g6165(.A0(n7252), .A1(n6161), .B0(n6191), .B1(n7255), .Y(n7299));
  OAI21X1 g6166(.A0(n7298), .A1(n6206), .B0(n7299), .Y(n7300));
  NOR2X1  g6167(.A(n7300), .B(n7297), .Y(n7301));
  OAI21X1 g6168(.A0(n7282), .A1(n7295), .B0(n7301), .Y(P2_U3227));
  NAND2X1 g6169(.A(n7243), .B(n6236), .Y(n7303));
  AOI22X1 g6170(.A0(n7282), .A1(P2_REG2_REG_7__SCAN_IN), .B0(n6211), .B1(n7252), .Y(n7304));
  OAI22X1 g6171(.A0(n7289), .A1(n6197), .B0(n6218), .B1(n7271), .Y(n7305));
  AOI21X1 g6172(.A0(n7247), .A1(n6242), .B0(n7305), .Y(n7306));
  NAND3X1 g6173(.A(n7306), .B(n7304), .C(n7303), .Y(P2_U3226));
  NOR3X1  g6174(.A(n6275), .B(n6274), .C(n6273), .Y(n7308));
  INVX1   g6175(.A(P2_REG2_REG_8__SCAN_IN), .Y(n7309));
  OAI22X1 g6176(.A0(n7243), .A1(n7309), .B0(n6291), .B1(n7270), .Y(n7310));
  AOI22X1 g6177(.A0(n7284), .A1(n6240), .B0(n6261), .B1(n7255), .Y(n7311));
  OAI21X1 g6178(.A0(n7298), .A1(n6296), .B0(n7311), .Y(n7312));
  NOR2X1  g6179(.A(n7312), .B(n7310), .Y(n7313));
  OAI21X1 g6180(.A0(n7282), .A1(n7308), .B0(n7313), .Y(P2_U3225));
  NAND2X1 g6181(.A(n7243), .B(n6323), .Y(n7315));
  AOI22X1 g6182(.A0(n7282), .A1(P2_REG2_REG_9__SCAN_IN), .B0(n6334), .B1(n7247), .Y(n7316));
  INVX1   g6183(.A(n6282), .Y(n7317));
  OAI22X1 g6184(.A0(n7289), .A1(n7317), .B0(n6360), .B1(n7270), .Y(n7318));
  AOI21X1 g6185(.A0(n7255), .A1(n6316), .B0(n7318), .Y(n7319));
  NAND3X1 g6186(.A(n7319), .B(n7316), .C(n7315), .Y(P2_U3224));
  NOR3X1  g6187(.A(n6371), .B(n6370), .C(n6369), .Y(n7321));
  INVX1   g6188(.A(P2_REG2_REG_10__SCAN_IN), .Y(n7322));
  OAI22X1 g6189(.A0(n7243), .A1(n7322), .B0(n6412), .B1(n7298), .Y(n7323));
  AOI22X1 g6190(.A0(n7284), .A1(n6330), .B0(n6353), .B1(n7252), .Y(n7324));
  OAI21X1 g6191(.A0(n7271), .A1(n6365), .B0(n7324), .Y(n7325));
  NOR2X1  g6192(.A(n7325), .B(n7323), .Y(n7326));
  OAI21X1 g6193(.A0(n7282), .A1(n7321), .B0(n7326), .Y(P2_U3223));
  AOI22X1 g6194(.A0(n7282), .A1(P2_REG2_REG_11__SCAN_IN), .B0(n6429), .B1(n7247), .Y(n7328));
  AOI22X1 g6195(.A0(n7284), .A1(n6377), .B0(n6423), .B1(n7252), .Y(n7329));
  NAND2X1 g6196(.A(n7329), .B(n7328), .Y(n7330));
  AOI21X1 g6197(.A0(n7255), .A1(n6402), .B0(n7330), .Y(n7331));
  OAI21X1 g6198(.A0(n7282), .A1(n6421), .B0(n7331), .Y(P2_U3222));
  INVX1   g6199(.A(P2_REG2_REG_12__SCAN_IN), .Y(n7333));
  OAI22X1 g6200(.A0(n7243), .A1(n7333), .B0(n6480), .B1(n7298), .Y(n7334));
  AOI22X1 g6201(.A0(n7284), .A1(n6427), .B0(n6441), .B1(n7252), .Y(n7335));
  OAI21X1 g6202(.A0(n7271), .A1(n6454), .B0(n7335), .Y(n7336));
  NOR2X1  g6203(.A(n7336), .B(n7334), .Y(n7337));
  OAI21X1 g6204(.A0(n7282), .A1(n6461), .B0(n7337), .Y(P2_U3221));
  NOR3X1  g6205(.A(n6509), .B(n6508), .C(n6507), .Y(n7339));
  OAI21X1 g6206(.A0(n7242), .A1(n5815), .B0(P2_REG2_REG_13__SCAN_IN), .Y(n7340));
  OAI21X1 g6207(.A0(n7298), .A1(n6527), .B0(n7340), .Y(n7341));
  AOI22X1 g6208(.A0(n7284), .A1(n6468), .B0(n6485), .B1(n7252), .Y(n7342));
  OAI21X1 g6209(.A0(n7271), .A1(n6503), .B0(n7342), .Y(n7343));
  NOR2X1  g6210(.A(n7343), .B(n7341), .Y(n7344));
  OAI21X1 g6211(.A0(n7282), .A1(n7339), .B0(n7344), .Y(P2_U3220));
  NAND2X1 g6212(.A(n7243), .B(n6548), .Y(n7346));
  NAND2X1 g6213(.A(n7255), .B(n6536), .Y(n7347));
  AOI22X1 g6214(.A0(n7282), .A1(P2_REG2_REG_14__SCAN_IN), .B0(n6559), .B1(n7247), .Y(n7348));
  AOI22X1 g6215(.A0(n7284), .A1(n6514), .B0(n6532), .B1(n7252), .Y(n7349));
  NAND4X1 g6216(.A(n7348), .B(n7347), .C(n7346), .D(n7349), .Y(P2_U3219));
  NAND2X1 g6217(.A(n7243), .B(n6587), .Y(n7351));
  NAND2X1 g6218(.A(n7255), .B(n6577), .Y(n7352));
  AOI22X1 g6219(.A0(n7282), .A1(P2_REG2_REG_15__SCAN_IN), .B0(n6593), .B1(n7247), .Y(n7353));
  INVX1   g6220(.A(n6556), .Y(n7354));
  AOI22X1 g6221(.A0(n7284), .A1(n7354), .B0(n6569), .B1(n7252), .Y(n7355));
  NAND4X1 g6222(.A(n7353), .B(n7352), .C(n7351), .D(n7355), .Y(P2_U3218));
  NOR3X1  g6223(.A(n6635), .B(n6631), .C(n6614), .Y(n7357));
  AOI22X1 g6224(.A0(n7282), .A1(P2_REG2_REG_16__SCAN_IN), .B0(n6645), .B1(n7247), .Y(n7358));
  AOI22X1 g6225(.A0(n7284), .A1(n6591), .B0(n6604), .B1(n7252), .Y(n7359));
  NAND2X1 g6226(.A(n7359), .B(n7358), .Y(n7360));
  AOI21X1 g6227(.A0(n7255), .A1(n6628), .B0(n7360), .Y(n7361));
  OAI21X1 g6228(.A0(n7282), .A1(n7357), .B0(n7361), .Y(P2_U3217));
  NOR3X1  g6229(.A(n6678), .B(n6677), .C(n6676), .Y(n7363));
  NOR2X1  g6230(.A(n7271), .B(n6672), .Y(n7364));
  INVX1   g6231(.A(P2_REG2_REG_17__SCAN_IN), .Y(n7365));
  OAI22X1 g6232(.A0(n7243), .A1(n7365), .B0(n6702), .B1(n7298), .Y(n7366));
  INVX1   g6233(.A(n6643), .Y(n7367));
  OAI22X1 g6234(.A0(n7289), .A1(n7367), .B0(n6657), .B1(n7270), .Y(n7368));
  NOR3X1  g6235(.A(n7368), .B(n7366), .C(n7364), .Y(n7369));
  OAI21X1 g6236(.A0(n7282), .A1(n7363), .B0(n7369), .Y(P2_U3216));
  AOI22X1 g6237(.A0(n7282), .A1(P2_REG2_REG_18__SCAN_IN), .B0(n6729), .B1(n7247), .Y(n7371));
  AOI22X1 g6238(.A0(n7284), .A1(n6682), .B0(n6721), .B1(n7252), .Y(n7372));
  NAND2X1 g6239(.A(n7372), .B(n7371), .Y(n7373));
  AOI21X1 g6240(.A0(n7255), .A1(n6712), .B0(n7373), .Y(n7374));
  OAI21X1 g6241(.A0(n7282), .A1(n6718), .B0(n7374), .Y(P2_U3215));
  INVX1   g6242(.A(P2_REG2_REG_19__SCAN_IN), .Y(n7376));
  OAI22X1 g6243(.A0(n7243), .A1(n7376), .B0(n6773), .B1(n7298), .Y(n7377));
  AOI21X1 g6244(.A0(n7284), .A1(n6727), .B0(n7377), .Y(n7378));
  OAI21X1 g6245(.A0(n7270), .A1(n6820), .B0(n7378), .Y(n7379));
  AOI21X1 g6246(.A0(n7255), .A1(n6754), .B0(n7379), .Y(n7380));
  OAI21X1 g6247(.A0(n7282), .A1(n6760), .B0(n7380), .Y(P2_U3214));
  NAND2X1 g6248(.A(n7243), .B(n6798), .Y(n7382));
  NAND2X1 g6249(.A(n7255), .B(n6780), .Y(n7383));
  AOI22X1 g6250(.A0(n7282), .A1(P2_REG2_REG_20__SCAN_IN), .B0(n6806), .B1(n7247), .Y(n7384));
  OAI21X1 g6251(.A0(n7289), .A1(n6764), .B0(n7384), .Y(n7385));
  AOI21X1 g6252(.A0(n7252), .A1(n6774), .B0(n7385), .Y(n7386));
  NAND3X1 g6253(.A(n7386), .B(n7383), .C(n7382), .Y(P2_U3213));
  NOR2X1  g6254(.A(n7271), .B(n6818), .Y(n7388));
  NOR3X1  g6255(.A(n7270), .B(n5870), .C(n5635), .Y(n7389));
  AOI22X1 g6256(.A0(n7282), .A1(P2_REG2_REG_21__SCAN_IN), .B0(n6842), .B1(n7247), .Y(n7390));
  OAI21X1 g6257(.A0(n7289), .A1(n6803), .B0(n7390), .Y(n7391));
  NOR3X1  g6258(.A(n7391), .B(n7389), .C(n7388), .Y(n7392));
  OAI21X1 g6259(.A0(n7282), .A1(n6835), .B0(n7392), .Y(P2_U3212));
  NAND2X1 g6260(.A(n7243), .B(n6871), .Y(n7394));
  NAND2X1 g6261(.A(n7255), .B(n6869), .Y(n7395));
  AOI22X1 g6262(.A0(n7282), .A1(P2_REG2_REG_22__SCAN_IN), .B0(n6878), .B1(n7247), .Y(n7396));
  OAI21X1 g6263(.A0(n7289), .A1(n6839), .B0(n7396), .Y(n7397));
  AOI21X1 g6264(.A0(n7252), .A1(n6849), .B0(n7397), .Y(n7398));
  NAND3X1 g6265(.A(n7398), .B(n7395), .C(n7394), .Y(P2_U3211));
  NOR3X1  g6266(.A(n6908), .B(n6907), .C(n6898), .Y(n7400));
  AOI21X1 g6267(.A0(n6897), .A1(n6889), .B0(n7271), .Y(n7401));
  NOR2X1  g6268(.A(n7270), .B(n6886), .Y(n7402));
  INVX1   g6269(.A(n6876), .Y(n7403));
  AOI22X1 g6270(.A0(n7282), .A1(P2_REG2_REG_23__SCAN_IN), .B0(n6916), .B1(n7247), .Y(n7404));
  OAI21X1 g6271(.A0(n7289), .A1(n7403), .B0(n7404), .Y(n7405));
  NOR3X1  g6272(.A(n7405), .B(n7402), .C(n7401), .Y(n7406));
  OAI21X1 g6273(.A0(n7282), .A1(n7400), .B0(n7406), .Y(P2_U3210));
  NOR3X1  g6274(.A(n6945), .B(n6942), .C(n6934), .Y(n7408));
  OAI21X1 g6275(.A0(n7242), .A1(n5815), .B0(P2_REG2_REG_24__SCAN_IN), .Y(n7409));
  OAI21X1 g6276(.A0(n7298), .A1(n6959), .B0(n7409), .Y(n7410));
  AOI21X1 g6277(.A0(n7284), .A1(n6914), .B0(n7410), .Y(n7411));
  OAI21X1 g6278(.A0(n7270), .A1(n6925), .B0(n7411), .Y(n7412));
  AOI21X1 g6279(.A0(n7255), .A1(n6943), .B0(n7412), .Y(n7413));
  OAI21X1 g6280(.A0(n7282), .A1(n7408), .B0(n7413), .Y(P2_U3209));
  NOR3X1  g6281(.A(n6981), .B(n6979), .C(n6972), .Y(n7415));
  OAI21X1 g6282(.A0(n7242), .A1(n5815), .B0(P2_REG2_REG_25__SCAN_IN), .Y(n7416));
  OAI21X1 g6283(.A0(n7298), .A1(n6994), .B0(n7416), .Y(n7417));
  AOI21X1 g6284(.A0(n7284), .A1(n6951), .B0(n7417), .Y(n7418));
  OAI21X1 g6285(.A0(n7270), .A1(n7046), .B0(n7418), .Y(n7419));
  AOI21X1 g6286(.A0(n7255), .A1(n6976), .B0(n7419), .Y(n7420));
  OAI21X1 g6287(.A0(n7282), .A1(n7415), .B0(n7420), .Y(P2_U3208));
  NOR3X1  g6288(.A(n7014), .B(n7013), .C(n7007), .Y(n7422));
  NOR2X1  g6289(.A(n7271), .B(n7011), .Y(n7423));
  NOR3X1  g6290(.A(n7270), .B(n5870), .C(n5677), .Y(n7424));
  AOI22X1 g6291(.A0(n7282), .A1(P2_REG2_REG_26__SCAN_IN), .B0(n7023), .B1(n7247), .Y(n7425));
  OAI21X1 g6292(.A0(n7289), .A1(n6984), .B0(n7425), .Y(n7426));
  NOR3X1  g6293(.A(n7426), .B(n7424), .C(n7423), .Y(n7427));
  OAI21X1 g6294(.A0(n7282), .A1(n7422), .B0(n7427), .Y(P2_U3207));
  NOR4X1  g6295(.A(n7054), .B(n7052), .C(n7042), .D(n7055), .Y(n7429));
  AOI21X1 g6296(.A0(n7041), .A1(n7037), .B0(n7271), .Y(n7430));
  NOR2X1  g6297(.A(n7270), .B(n7034), .Y(n7431));
  INVX1   g6298(.A(n7021), .Y(n7432));
  AOI22X1 g6299(.A0(n7282), .A1(P2_REG2_REG_27__SCAN_IN), .B0(n7064), .B1(n7247), .Y(n7433));
  OAI21X1 g6300(.A0(n7289), .A1(n7432), .B0(n7433), .Y(n7434));
  NOR3X1  g6301(.A(n7434), .B(n7431), .C(n7430), .Y(n7435));
  OAI21X1 g6302(.A0(n7282), .A1(n7429), .B0(n7435), .Y(P2_U3206));
  NOR2X1  g6303(.A(n7271), .B(n7079), .Y(n7437));
  NOR3X1  g6304(.A(n7270), .B(n5870), .C(n5695), .Y(n7438));
  AOI22X1 g6305(.A0(n7282), .A1(P2_REG2_REG_28__SCAN_IN), .B0(n7100), .B1(n7247), .Y(n7439));
  OAI21X1 g6306(.A0(n7289), .A1(n7061), .B0(n7439), .Y(n7440));
  NOR3X1  g6307(.A(n7440), .B(n7438), .C(n7437), .Y(n7441));
  OAI21X1 g6308(.A0(n7282), .A1(n7091), .B0(n7441), .Y(P2_U3205));
  OAI21X1 g6309(.A0(n7138), .A1(n7127), .B0(n7243), .Y(n7443));
  AOI22X1 g6310(.A0(n7282), .A1(P2_REG2_REG_29__SCAN_IN), .B0(n7094), .B1(n7284), .Y(n7444));
  OAI21X1 g6311(.A0(n7270), .A1(n7114), .B0(n7444), .Y(n7445));
  AOI21X1 g6312(.A0(n7255), .A1(n7120), .B0(n7445), .Y(n7446));
  NAND2X1 g6313(.A(n7446), .B(n7443), .Y(P2_U3204));
  OAI21X1 g6314(.A0(n5713), .A1(n5711), .B0(n6823), .Y(n7448));
  NAND3X1 g6315(.A(n7243), .B(n7146), .C(n7135), .Y(n7449));
  OAI21X1 g6316(.A0(n7289), .A1(n7095), .B0(n7449), .Y(n7450));
  AOI21X1 g6317(.A0(n7282), .A1(P2_REG2_REG_30__SCAN_IN), .B0(n7450), .Y(n7451));
  OAI21X1 g6318(.A0(n7270), .A1(n7448), .B0(n7451), .Y(P2_U3203));
  NAND2X1 g6319(.A(n6823), .B(n5721), .Y(n7453));
  AOI21X1 g6320(.A0(n7282), .A1(P2_REG2_REG_31__SCAN_IN), .B0(n7450), .Y(n7454));
  OAI21X1 g6321(.A0(n7270), .A1(n7453), .B0(n7454), .Y(P2_U3202));
  AOI21X1 g6322(.A0(n5739), .A1(n5728), .B0(P2_U3151), .Y(n7456));
  NAND2X1 g6323(.A(n6823), .B(n5729), .Y(n7457));
  OAI21X1 g6324(.A0(n5844), .A1(n5846), .B0(n6823), .Y(n7458));
  NAND3X1 g6325(.A(n7458), .B(n7457), .C(n7456), .Y(n7459));
  INVX1   g6326(.A(n7459), .Y(n7460));
  NOR2X1  g6327(.A(n7460), .B(n5815), .Y(n7461));
  NOR2X1  g6328(.A(n6601), .B(P2_REG2_REG_16__SCAN_IN), .Y(n7462));
  INVX1   g6329(.A(P2_REG2_REG_15__SCAN_IN), .Y(n7463));
  INVX1   g6330(.A(P2_REG2_REG_14__SCAN_IN), .Y(n7464));
  NAND2X1 g6331(.A(n6530), .B(n7464), .Y(n7465));
  NOR2X1  g6332(.A(n6530), .B(n7464), .Y(n7466));
  NOR2X1  g6333(.A(n6482), .B(P2_REG2_REG_13__SCAN_IN), .Y(n7467));
  NAND2X1 g6334(.A(n6482), .B(P2_REG2_REG_13__SCAN_IN), .Y(n7468));
  NAND2X1 g6335(.A(n6439), .B(n7333), .Y(n7469));
  NOR2X1  g6336(.A(n6439), .B(n7333), .Y(n7470));
  NOR2X1  g6337(.A(n6390), .B(P2_REG2_REG_11__SCAN_IN), .Y(n7471));
  NAND2X1 g6338(.A(n6390), .B(P2_REG2_REG_11__SCAN_IN), .Y(n7472));
  NAND2X1 g6339(.A(n6344), .B(n7322), .Y(n7473));
  NOR2X1  g6340(.A(n6344), .B(n7322), .Y(n7474));
  NOR2X1  g6341(.A(n6298), .B(P2_REG2_REG_9__SCAN_IN), .Y(n7475));
  NAND2X1 g6342(.A(n6298), .B(P2_REG2_REG_9__SCAN_IN), .Y(n7476));
  NAND2X1 g6343(.A(n6252), .B(n7309), .Y(n7477));
  NOR2X1  g6344(.A(n6252), .B(n7309), .Y(n7478));
  NOR2X1  g6345(.A(n6208), .B(P2_REG2_REG_7__SCAN_IN), .Y(n7479));
  NAND2X1 g6346(.A(n6208), .B(P2_REG2_REG_7__SCAN_IN), .Y(n7480));
  NAND2X1 g6347(.A(n6159), .B(n7296), .Y(n7481));
  NOR2X1  g6348(.A(n6159), .B(n7296), .Y(n7482));
  NOR2X1  g6349(.A(n6117), .B(P2_REG2_REG_5__SCAN_IN), .Y(n7483));
  NAND2X1 g6350(.A(n6117), .B(P2_REG2_REG_5__SCAN_IN), .Y(n7484));
  INVX1   g6351(.A(P2_REG2_REG_4__SCAN_IN), .Y(n7485));
  NAND2X1 g6352(.A(n6065), .B(n7485), .Y(n7486));
  NOR2X1  g6353(.A(n6065), .B(n7485), .Y(n7487));
  NOR3X1  g6354(.A(n5874), .B(n5872), .C(n7244), .Y(n7488));
  NOR2X1  g6355(.A(n7488), .B(P2_REG2_REG_1__SCAN_IN), .Y(n7489));
  AOI21X1 g6356(.A0(n7488), .A1(P2_REG2_REG_1__SCAN_IN), .B0(n5936), .Y(n7490));
  NOR2X1  g6357(.A(n7490), .B(n7489), .Y(n7491));
  AOI21X1 g6358(.A0(n5978), .A1(P2_REG2_REG_2__SCAN_IN), .B0(n7491), .Y(n7492));
  AOI21X1 g6359(.A0(n5979), .A1(n7267), .B0(n7492), .Y(n7493));
  AOI21X1 g6360(.A0(n6020), .A1(P2_REG2_REG_3__SCAN_IN), .B0(n7493), .Y(n7494));
  AOI21X1 g6361(.A0(n6021), .A1(n7276), .B0(n7494), .Y(n7495));
  OAI21X1 g6362(.A0(n7495), .A1(n7487), .B0(n7486), .Y(n7496));
  AOI21X1 g6363(.A0(n7496), .A1(n7484), .B0(n7483), .Y(n7497));
  OAI21X1 g6364(.A0(n7497), .A1(n7482), .B0(n7481), .Y(n7498));
  AOI21X1 g6365(.A0(n7498), .A1(n7480), .B0(n7479), .Y(n7499));
  OAI21X1 g6366(.A0(n7499), .A1(n7478), .B0(n7477), .Y(n7500));
  AOI21X1 g6367(.A0(n7500), .A1(n7476), .B0(n7475), .Y(n7501));
  OAI21X1 g6368(.A0(n7501), .A1(n7474), .B0(n7473), .Y(n7502));
  AOI21X1 g6369(.A0(n7502), .A1(n7472), .B0(n7471), .Y(n7503));
  OAI21X1 g6370(.A0(n7503), .A1(n7470), .B0(n7469), .Y(n7504));
  AOI21X1 g6371(.A0(n7504), .A1(n7468), .B0(n7467), .Y(n7505));
  OAI21X1 g6372(.A0(n7505), .A1(n7466), .B0(n7465), .Y(n7506));
  NAND2X1 g6373(.A(n7506), .B(n7463), .Y(n7507));
  OAI21X1 g6374(.A0(n7506), .A1(n7463), .B0(n6567), .Y(n7508));
  AOI22X1 g6375(.A0(n7507), .A1(n7508), .B0(n6601), .B1(P2_REG2_REG_16__SCAN_IN), .Y(n7509));
  OAI22X1 g6376(.A0(n7462), .A1(n7509), .B0(n6655), .B1(n7365), .Y(n7510));
  OAI21X1 g6377(.A0(n6654), .A1(P2_REG2_REG_17__SCAN_IN), .B0(n7510), .Y(n7511));
  NOR2X1  g6378(.A(n6696), .B(P2_REG2_REG_18__SCAN_IN), .Y(n7512));
  XOR2X1  g6379(.A(n5853), .B(P2_REG2_REG_19__SCAN_IN), .Y(n7513));
  AOI21X1 g6380(.A0(n6696), .A1(P2_REG2_REG_18__SCAN_IN), .B0(n7513), .Y(n7514));
  OAI21X1 g6381(.A0(n7512), .A1(n7511), .B0(n7514), .Y(n7515));
  INVX1   g6382(.A(n7512), .Y(n7516));
  INVX1   g6383(.A(P2_REG2_REG_18__SCAN_IN), .Y(n7517));
  OAI21X1 g6384(.A0(n6697), .A1(n7517), .B0(n7511), .Y(n7518));
  NAND3X1 g6385(.A(n7518), .B(n7513), .C(n7516), .Y(n7519));
  NOR2X1  g6386(.A(n5915), .B(n5914), .Y(n7520));
  INVX1   g6387(.A(n7520), .Y(n7521));
  NAND4X1 g6388(.A(n5846), .B(n7251), .C(n7283), .D(n5844), .Y(n7524));
  INVX1   g6389(.A(n7524), .Y(n7525));
  AOI21X1 g6390(.A0(n7519), .A1(n7515), .B0(n7521), .Y(n7528));
  NOR2X1  g6391(.A(n6654), .B(P2_REG1_REG_17__SCAN_IN), .Y(n7529));
  INVX1   g6392(.A(P2_REG1_REG_17__SCAN_IN), .Y(n7530));
  NOR2X1  g6393(.A(n6655), .B(n7530), .Y(n7531));
  INVX1   g6394(.A(n7531), .Y(n7532));
  INVX1   g6395(.A(P2_REG1_REG_16__SCAN_IN), .Y(n7533));
  INVX1   g6396(.A(P2_REG1_REG_14__SCAN_IN), .Y(n7534));
  NOR2X1  g6397(.A(n6530), .B(n7534), .Y(n7535));
  NOR2X1  g6398(.A(n6482), .B(P2_REG1_REG_13__SCAN_IN), .Y(n7536));
  NAND2X1 g6399(.A(n6482), .B(P2_REG1_REG_13__SCAN_IN), .Y(n7537));
  INVX1   g6400(.A(P2_REG1_REG_12__SCAN_IN), .Y(n7538));
  NAND2X1 g6401(.A(n6439), .B(n7538), .Y(n7539));
  NOR2X1  g6402(.A(n6439), .B(n7538), .Y(n7540));
  NOR2X1  g6403(.A(n6390), .B(P2_REG1_REG_11__SCAN_IN), .Y(n7541));
  NAND2X1 g6404(.A(n6390), .B(P2_REG1_REG_11__SCAN_IN), .Y(n7542));
  INVX1   g6405(.A(P2_REG1_REG_10__SCAN_IN), .Y(n7543));
  NAND2X1 g6406(.A(n6344), .B(n7543), .Y(n7544));
  NOR2X1  g6407(.A(n6344), .B(n7543), .Y(n7545));
  INVX1   g6408(.A(P2_REG1_REG_9__SCAN_IN), .Y(n7546));
  INVX1   g6409(.A(P2_REG1_REG_8__SCAN_IN), .Y(n7547));
  NOR2X1  g6410(.A(n6208), .B(P2_REG1_REG_7__SCAN_IN), .Y(n7548));
  NAND2X1 g6411(.A(n6208), .B(P2_REG1_REG_7__SCAN_IN), .Y(n7549));
  INVX1   g6412(.A(P2_REG1_REG_6__SCAN_IN), .Y(n7550));
  NAND2X1 g6413(.A(n6159), .B(n7550), .Y(n7551));
  NOR2X1  g6414(.A(n6159), .B(n7550), .Y(n7552));
  NOR2X1  g6415(.A(n6117), .B(P2_REG1_REG_5__SCAN_IN), .Y(n7553));
  NAND2X1 g6416(.A(n6117), .B(P2_REG1_REG_5__SCAN_IN), .Y(n7554));
  INVX1   g6417(.A(P2_REG1_REG_4__SCAN_IN), .Y(n7555));
  NAND2X1 g6418(.A(n6065), .B(n7555), .Y(n7556));
  NOR2X1  g6419(.A(n6065), .B(n7555), .Y(n7557));
  INVX1   g6420(.A(P2_REG1_REG_3__SCAN_IN), .Y(n7558));
  NOR2X1  g6421(.A(n5978), .B(P2_REG1_REG_2__SCAN_IN), .Y(n7559));
  INVX1   g6422(.A(n7559), .Y(n7560));
  INVX1   g6423(.A(P2_REG1_REG_2__SCAN_IN), .Y(n7561));
  NOR3X1  g6424(.A(n5874), .B(n5872), .C(n7157), .Y(n7562));
  NOR2X1  g6425(.A(n7562), .B(P2_REG1_REG_1__SCAN_IN), .Y(n7563));
  AOI21X1 g6426(.A0(n7562), .A1(P2_REG1_REG_1__SCAN_IN), .B0(n5936), .Y(n7564));
  OAI22X1 g6427(.A0(n7563), .A1(n7564), .B0(n5979), .B1(n7561), .Y(n7565));
  AOI22X1 g6428(.A0(n7560), .A1(n7565), .B0(n6020), .B1(P2_REG1_REG_3__SCAN_IN), .Y(n7566));
  AOI21X1 g6429(.A0(n6021), .A1(n7558), .B0(n7566), .Y(n7567));
  OAI21X1 g6430(.A0(n7567), .A1(n7557), .B0(n7556), .Y(n7568));
  AOI21X1 g6431(.A0(n7568), .A1(n7554), .B0(n7553), .Y(n7569));
  OAI21X1 g6432(.A0(n7569), .A1(n7552), .B0(n7551), .Y(n7570));
  AOI21X1 g6433(.A0(n7570), .A1(n7549), .B0(n7548), .Y(n7571));
  AOI21X1 g6434(.A0(n6251), .A1(P2_REG1_REG_8__SCAN_IN), .B0(n7571), .Y(n7572));
  AOI21X1 g6435(.A0(n6252), .A1(n7547), .B0(n7572), .Y(n7573));
  AOI21X1 g6436(.A0(n6298), .A1(P2_REG1_REG_9__SCAN_IN), .B0(n7573), .Y(n7574));
  AOI21X1 g6437(.A0(n6299), .A1(n7546), .B0(n7574), .Y(n7575));
  OAI21X1 g6438(.A0(n7575), .A1(n7545), .B0(n7544), .Y(n7576));
  AOI21X1 g6439(.A0(n7576), .A1(n7542), .B0(n7541), .Y(n7577));
  OAI21X1 g6440(.A0(n7577), .A1(n7540), .B0(n7539), .Y(n7578));
  AOI21X1 g6441(.A0(n7578), .A1(n7537), .B0(n7536), .Y(n7579));
  NOR2X1  g6442(.A(n7579), .B(n7535), .Y(n7580));
  AOI21X1 g6443(.A0(n6530), .A1(n7534), .B0(n7580), .Y(n7581));
  NOR2X1  g6444(.A(n7581), .B(P2_REG1_REG_15__SCAN_IN), .Y(n7582));
  AOI21X1 g6445(.A0(n7581), .A1(P2_REG1_REG_15__SCAN_IN), .B0(n6566), .Y(n7583));
  OAI22X1 g6446(.A0(n7582), .A1(n7583), .B0(n6602), .B1(n7533), .Y(n7584));
  OAI21X1 g6447(.A0(n6601), .A1(P2_REG1_REG_16__SCAN_IN), .B0(n7584), .Y(n7585));
  AOI21X1 g6448(.A0(n7585), .A1(n7532), .B0(n7529), .Y(n7586));
  OAI21X1 g6449(.A0(n6696), .A1(P2_REG1_REG_18__SCAN_IN), .B0(n7586), .Y(n7587));
  XOR2X1  g6450(.A(n5853), .B(P2_REG1_REG_19__SCAN_IN), .Y(n7588));
  AOI21X1 g6451(.A0(n6696), .A1(P2_REG1_REG_18__SCAN_IN), .B0(n7588), .Y(n7589));
  AOI21X1 g6452(.A0(n6696), .A1(P2_REG1_REG_18__SCAN_IN), .B0(n7586), .Y(n7590));
  OAI21X1 g6453(.A0(n6696), .A1(P2_REG1_REG_18__SCAN_IN), .B0(n7588), .Y(n7591));
  NOR2X1  g6454(.A(n7591), .B(n7590), .Y(n7592));
  AOI21X1 g6455(.A0(n7589), .A1(n7587), .B0(n7592), .Y(n7593));
  INVX1   g6456(.A(n5915), .Y(n7596));
  OAI22X1 g6457(.A0(n5867), .A1(n7593), .B0(n5853), .B1(n7596), .Y(n7599));
  OAI21X1 g6458(.A0(n7599), .A1(n7528), .B0(n7461), .Y(n7600));
  NOR4X1  g6459(.A(n5867), .B(n5728), .C(P2_U3151), .D(n7460), .Y(n7601));
  INVX1   g6460(.A(n7601), .Y(n7602));
  NOR2X1  g6461(.A(n7602), .B(n7593), .Y(n7603));
  NOR4X1  g6462(.A(n7521), .B(n5728), .C(P2_U3151), .D(n7460), .Y(n7604));
  INVX1   g6463(.A(n7604), .Y(n7605));
  AOI21X1 g6464(.A0(n7519), .A1(n7515), .B0(n7605), .Y(n7606));
  NOR2X1  g6465(.A(n5914), .B(n7376), .Y(n7607));
  AOI21X1 g6466(.A0(n5914), .A1(P2_REG1_REG_19__SCAN_IN), .B0(n7607), .Y(n7608));
  XOR2X1  g6467(.A(n7608), .B(n5853), .Y(n7609));
  NAND2X1 g6468(.A(n5914), .B(P2_REG1_REG_18__SCAN_IN), .Y(n7610));
  OAI21X1 g6469(.A0(n5914), .A1(n7517), .B0(n7610), .Y(n7611));
  NOR2X1  g6470(.A(n5867), .B(n7530), .Y(n7612));
  AOI21X1 g6471(.A0(n5867), .A1(P2_REG2_REG_17__SCAN_IN), .B0(n7612), .Y(n7613));
  INVX1   g6472(.A(n7613), .Y(n7614));
  NAND2X1 g6473(.A(n7614), .B(n6654), .Y(n7615));
  NOR2X1  g6474(.A(n7614), .B(n6654), .Y(n7616));
  NOR2X1  g6475(.A(n5867), .B(n7533), .Y(n7617));
  AOI21X1 g6476(.A0(n5867), .A1(P2_REG2_REG_16__SCAN_IN), .B0(n7617), .Y(n7618));
  INVX1   g6477(.A(n7618), .Y(n7619));
  NOR2X1  g6478(.A(n7619), .B(n6601), .Y(n7620));
  NOR2X1  g6479(.A(n5867), .B(n6551), .Y(n7621));
  AOI21X1 g6480(.A0(n5867), .A1(P2_REG2_REG_15__SCAN_IN), .B0(n7621), .Y(n7622));
  NOR2X1  g6481(.A(n7622), .B(n6567), .Y(n7623));
  AOI21X1 g6482(.A0(n7619), .A1(n6601), .B0(n7623), .Y(n7624));
  INVX1   g6483(.A(n7620), .Y(n7625));
  NOR2X1  g6484(.A(n5867), .B(n7534), .Y(n7626));
  AOI21X1 g6485(.A0(n5867), .A1(P2_REG2_REG_14__SCAN_IN), .B0(n7626), .Y(n7627));
  NOR2X1  g6486(.A(n7627), .B(n6530), .Y(n7628));
  NAND2X1 g6487(.A(n7622), .B(n6567), .Y(n7629));
  NAND3X1 g6488(.A(n7629), .B(n7628), .C(n7625), .Y(n7630));
  AOI21X1 g6489(.A0(n7630), .A1(n7624), .B0(n7620), .Y(n7631));
  INVX1   g6490(.A(P2_REG1_REG_13__SCAN_IN), .Y(n7632));
  NOR2X1  g6491(.A(n5867), .B(n7632), .Y(n7633));
  AOI21X1 g6492(.A0(n5867), .A1(P2_REG2_REG_13__SCAN_IN), .B0(n7633), .Y(n7634));
  NAND2X1 g6493(.A(n7634), .B(n6483), .Y(n7635));
  NOR2X1  g6494(.A(n5867), .B(n7538), .Y(n7636));
  AOI21X1 g6495(.A0(n5867), .A1(P2_REG2_REG_12__SCAN_IN), .B0(n7636), .Y(n7637));
  NAND2X1 g6496(.A(n7637), .B(n6439), .Y(n7638));
  INVX1   g6497(.A(P2_REG1_REG_11__SCAN_IN), .Y(n7639));
  NOR2X1  g6498(.A(n5867), .B(n7639), .Y(n7640));
  AOI21X1 g6499(.A0(n5867), .A1(P2_REG2_REG_11__SCAN_IN), .B0(n7640), .Y(n7641));
  INVX1   g6500(.A(n7641), .Y(n7642));
  NOR2X1  g6501(.A(n7642), .B(n6390), .Y(n7643));
  NOR2X1  g6502(.A(n5867), .B(n7543), .Y(n7644));
  AOI21X1 g6503(.A0(n5867), .A1(P2_REG2_REG_10__SCAN_IN), .B0(n7644), .Y(n7645));
  NOR2X1  g6504(.A(n7645), .B(n6344), .Y(n7646));
  NOR2X1  g6505(.A(n7641), .B(n6391), .Y(n7647));
  NOR2X1  g6506(.A(n7647), .B(n7646), .Y(n7648));
  INVX1   g6507(.A(n7648), .Y(n7649));
  NOR2X1  g6508(.A(n5867), .B(n7546), .Y(n7650));
  AOI21X1 g6509(.A0(n5867), .A1(P2_REG2_REG_9__SCAN_IN), .B0(n7650), .Y(n7651));
  INVX1   g6510(.A(n7645), .Y(n7652));
  NOR2X1  g6511(.A(n7652), .B(n6343), .Y(n7653));
  NOR4X1  g6512(.A(n7651), .B(n7643), .C(n6299), .D(n7653), .Y(n7654));
  NOR2X1  g6513(.A(n7654), .B(n7649), .Y(n7655));
  AOI22X1 g6514(.A0(n7641), .A1(n6391), .B0(n6344), .B1(n7645), .Y(n7656));
  NOR2X1  g6515(.A(n5867), .B(n7550), .Y(n7657));
  AOI21X1 g6516(.A0(n5867), .A1(P2_REG2_REG_6__SCAN_IN), .B0(n7657), .Y(n7658));
  INVX1   g6517(.A(n7658), .Y(n7659));
  NOR2X1  g6518(.A(n7659), .B(n6158), .Y(n7660));
  INVX1   g6519(.A(n7660), .Y(n7661));
  INVX1   g6520(.A(n6117), .Y(n7662));
  NOR2X1  g6521(.A(n5867), .B(n6111), .Y(n7663));
  AOI21X1 g6522(.A0(n5867), .A1(P2_REG2_REG_5__SCAN_IN), .B0(n7663), .Y(n7664));
  NOR2X1  g6523(.A(n7664), .B(n7662), .Y(n7665));
  AOI21X1 g6524(.A0(n7659), .A1(n6158), .B0(n7665), .Y(n7666));
  INVX1   g6525(.A(n7666), .Y(n7667));
  NOR2X1  g6526(.A(n5867), .B(n7555), .Y(n7668));
  AOI21X1 g6527(.A0(n5867), .A1(P2_REG2_REG_4__SCAN_IN), .B0(n7668), .Y(n7669));
  NAND2X1 g6528(.A(n7664), .B(n7662), .Y(n7670));
  INVX1   g6529(.A(n7670), .Y(n7671));
  NOR4X1  g6530(.A(n7669), .B(n7660), .C(n6065), .D(n7671), .Y(n7672));
  OAI21X1 g6531(.A0(n7672), .A1(n7667), .B0(n7661), .Y(n7673));
  NOR2X1  g6532(.A(n5867), .B(n7169), .Y(n7674));
  AOI21X1 g6533(.A0(n5867), .A1(P2_REG2_REG_1__SCAN_IN), .B0(n7674), .Y(n7675));
  NOR2X1  g6534(.A(n5867), .B(n7157), .Y(n7676));
  AOI21X1 g6535(.A0(n5867), .A1(P2_REG2_REG_0__SCAN_IN), .B0(n7676), .Y(n7677));
  NAND2X1 g6536(.A(n7677), .B(n5876), .Y(n7678));
  INVX1   g6537(.A(n7678), .Y(n7679));
  NAND3X1 g6538(.A(n7677), .B(n7675), .C(n5876), .Y(n7680));
  NAND2X1 g6539(.A(n7680), .B(n5936), .Y(n7681));
  OAI21X1 g6540(.A0(n7679), .A1(n7675), .B0(n7681), .Y(n7682));
  NOR2X1  g6541(.A(n5867), .B(n7558), .Y(n7683));
  AOI21X1 g6542(.A0(n5867), .A1(P2_REG2_REG_3__SCAN_IN), .B0(n7683), .Y(n7684));
  NOR2X1  g6543(.A(n5867), .B(n7561), .Y(n7685));
  AOI21X1 g6544(.A0(n5867), .A1(P2_REG2_REG_2__SCAN_IN), .B0(n7685), .Y(n7686));
  AOI22X1 g6545(.A0(n7684), .A1(n6021), .B0(n5979), .B1(n7686), .Y(n7687));
  NAND2X1 g6546(.A(n7687), .B(n7682), .Y(n7688));
  OAI21X1 g6547(.A0(n7686), .A1(n5979), .B0(n7684), .Y(n7689));
  NOR3X1  g6548(.A(n7686), .B(n7684), .C(n5979), .Y(n7690));
  AOI21X1 g6549(.A0(n7689), .A1(n6020), .B0(n7690), .Y(n7691));
  NAND2X1 g6550(.A(n7691), .B(n7688), .Y(n7692));
  NAND2X1 g6551(.A(n7669), .B(n6065), .Y(n7693));
  NAND4X1 g6552(.A(n7692), .B(n7670), .C(n7661), .D(n7693), .Y(n7694));
  NAND2X1 g6553(.A(n7694), .B(n7673), .Y(n7695));
  INVX1   g6554(.A(n7695), .Y(n7696));
  NOR2X1  g6555(.A(n5867), .B(n7547), .Y(n7697));
  AOI21X1 g6556(.A0(n5867), .A1(P2_REG2_REG_8__SCAN_IN), .B0(n7697), .Y(n7698));
  INVX1   g6557(.A(n7698), .Y(n7699));
  INVX1   g6558(.A(P2_REG1_REG_7__SCAN_IN), .Y(n7700));
  NOR2X1  g6559(.A(n5867), .B(n7700), .Y(n7701));
  AOI21X1 g6560(.A0(n5867), .A1(P2_REG2_REG_7__SCAN_IN), .B0(n7701), .Y(n7702));
  INVX1   g6561(.A(n7702), .Y(n7703));
  OAI22X1 g6562(.A0(n7699), .A1(n6251), .B0(n6208), .B1(n7703), .Y(n7704));
  OAI21X1 g6563(.A0(n7702), .A1(n6209), .B0(n7698), .Y(n7705));
  NOR3X1  g6564(.A(n7702), .B(n7698), .C(n6209), .Y(n7706));
  AOI21X1 g6565(.A0(n7705), .A1(n6251), .B0(n7706), .Y(n7707));
  OAI21X1 g6566(.A0(n7704), .A1(n7696), .B0(n7707), .Y(n7708));
  NAND2X1 g6567(.A(n7651), .B(n6299), .Y(n7709));
  NAND3X1 g6568(.A(n7709), .B(n7708), .C(n7656), .Y(n7710));
  OAI21X1 g6569(.A0(n7655), .A1(n7643), .B0(n7710), .Y(n7711));
  NAND2X1 g6570(.A(n7711), .B(n7638), .Y(n7712));
  OAI21X1 g6571(.A0(n7637), .A1(n6439), .B0(n7712), .Y(n7713));
  NAND2X1 g6572(.A(n7713), .B(n7635), .Y(n7714));
  OAI21X1 g6573(.A0(n7634), .A1(n6483), .B0(n7714), .Y(n7715));
  OAI21X1 g6574(.A0(n7619), .A1(n6601), .B0(n7629), .Y(n7716));
  AOI21X1 g6575(.A0(n7627), .A1(n6530), .B0(n7716), .Y(n7717));
  AOI21X1 g6576(.A0(n7717), .A1(n7715), .B0(n7631), .Y(n7718));
  OAI21X1 g6577(.A0(n7718), .A1(n7616), .B0(n7615), .Y(n7719));
  NAND2X1 g6578(.A(n7719), .B(n7611), .Y(n7720));
  OAI21X1 g6579(.A0(n7719), .A1(n7611), .B0(n6696), .Y(n7721));
  NAND2X1 g6580(.A(n7721), .B(n7720), .Y(n7722));
  XOR2X1  g6581(.A(n7722), .B(n7609), .Y(n7723));
  NOR3X1  g6582(.A(n5869), .B(n5868), .C(n5914), .Y(n7724));
  NAND3X1 g6583(.A(n5739), .B(n5728), .C(P2_STATE_REG_SCAN_IN), .Y(n7725));
  INVX1   g6584(.A(n7725), .Y(P2_U3893));
  OAI21X1 g6585(.A0(n7724), .A1(n5870), .B0(P2_U3893), .Y(n7727));
  NOR4X1  g6586(.A(n7596), .B(n5728), .C(P2_U3151), .D(n7460), .Y(n7728));
  AOI21X1 g6587(.A0(P2_U3893), .A1(n7596), .B0(n7728), .Y(n7729));
  INVX1   g6588(.A(n7729), .Y(n7730));
  OAI22X1 g6589(.A0(n1147), .A1(n7459), .B0(n6723), .B1(P2_STATE_REG_SCAN_IN), .Y(n7731));
  AOI21X1 g6590(.A0(n7730), .A1(n5860), .B0(n7731), .Y(n7732));
  OAI21X1 g6591(.A0(n7727), .A1(n7723), .B0(n7732), .Y(n7733));
  NOR3X1  g6592(.A(n7733), .B(n7606), .C(n7603), .Y(n7734));
  NAND2X1 g6593(.A(n7734), .B(n7600), .Y(P2_U3201));
  INVX1   g6594(.A(n7461), .Y(n7736));
  XOR2X1  g6595(.A(n6696), .B(P2_REG2_REG_18__SCAN_IN), .Y(n7737));
  XOR2X1  g6596(.A(n7737), .B(n7511), .Y(n7738));
  XOR2X1  g6597(.A(n6696), .B(P2_REG1_REG_18__SCAN_IN), .Y(n7739));
  XOR2X1  g6598(.A(n7739), .B(n7586), .Y(n7740));
  OAI22X1 g6599(.A0(n7596), .A1(n6696), .B0(n5867), .B1(n7740), .Y(n7741));
  AOI21X1 g6600(.A0(n7738), .A1(n7520), .B0(n7741), .Y(n7742));
  NOR2X1  g6601(.A(n7740), .B(n7602), .Y(n7743));
  INVX1   g6602(.A(n7738), .Y(n7744));
  NOR2X1  g6603(.A(n7744), .B(n7605), .Y(n7745));
  XOR2X1  g6604(.A(n7611), .B(n6697), .Y(n7746));
  XOR2X1  g6605(.A(n7746), .B(n7719), .Y(n7747));
  NOR2X1  g6606(.A(n7747), .B(n7727), .Y(n7748));
  AOI22X1 g6607(.A0(P2_ADDR_REG_18__SCAN_IN), .A1(n7460), .B0(P2_REG3_REG_18__SCAN_IN), .B1(P2_U3151), .Y(n7749));
  OAI21X1 g6608(.A0(n7729), .A1(n6696), .B0(n7749), .Y(n7750));
  NOR4X1  g6609(.A(n7748), .B(n7745), .C(n7743), .D(n7750), .Y(n7751));
  OAI21X1 g6610(.A0(n7742), .A1(n7736), .B0(n7751), .Y(P2_U3200));
  NOR2X1  g6611(.A(n7509), .B(n7462), .Y(n7753));
  XOR2X1  g6612(.A(n6654), .B(P2_REG2_REG_17__SCAN_IN), .Y(n7754));
  XOR2X1  g6613(.A(n7754), .B(n7753), .Y(n7755));
  XOR2X1  g6614(.A(n6654), .B(P2_REG1_REG_17__SCAN_IN), .Y(n7756));
  XOR2X1  g6615(.A(n7756), .B(n7585), .Y(n7757));
  AOI22X1 g6616(.A0(n5915), .A1(n6655), .B0(n5914), .B1(n7757), .Y(n7758));
  OAI21X1 g6617(.A0(n7755), .A1(n7521), .B0(n7758), .Y(n7759));
  NAND2X1 g6618(.A(n7759), .B(n7461), .Y(n7760));
  INVX1   g6619(.A(n7727), .Y(n7761));
  XOR2X1  g6620(.A(n7613), .B(n6654), .Y(n7762));
  XOR2X1  g6621(.A(n7762), .B(n7718), .Y(n7763));
  AOI22X1 g6622(.A0(P2_ADDR_REG_17__SCAN_IN), .A1(n7460), .B0(P2_REG3_REG_17__SCAN_IN), .B1(P2_U3151), .Y(n7764));
  OAI21X1 g6623(.A0(n7729), .A1(n6654), .B0(n7764), .Y(n7765));
  AOI21X1 g6624(.A0(n7763), .A1(n7761), .B0(n7765), .Y(n7766));
  OAI21X1 g6625(.A0(n7755), .A1(n7605), .B0(n7766), .Y(n7767));
  AOI21X1 g6626(.A0(n7757), .A1(n7601), .B0(n7767), .Y(n7768));
  NAND2X1 g6627(.A(n7768), .B(n7760), .Y(P2_U3199));
  NAND2X1 g6628(.A(n7508), .B(n7507), .Y(n7770));
  XOR2X1  g6629(.A(n6601), .B(P2_REG2_REG_16__SCAN_IN), .Y(n7771));
  XOR2X1  g6630(.A(n7771), .B(n7770), .Y(n7772));
  INVX1   g6631(.A(n7581), .Y(n7773));
  AOI21X1 g6632(.A0(n7773), .A1(n6551), .B0(n7583), .Y(n7774));
  XOR2X1  g6633(.A(n6601), .B(P2_REG1_REG_16__SCAN_IN), .Y(n7775));
  XOR2X1  g6634(.A(n7775), .B(n7774), .Y(n7776));
  OAI22X1 g6635(.A0(n7596), .A1(n6601), .B0(n5867), .B1(n7776), .Y(n7777));
  AOI21X1 g6636(.A0(n7772), .A1(n7520), .B0(n7777), .Y(n7778));
  NOR2X1  g6637(.A(n7776), .B(n7602), .Y(n7779));
  INVX1   g6638(.A(n7772), .Y(n7780));
  NOR2X1  g6639(.A(n7780), .B(n7605), .Y(n7781));
  NAND2X1 g6640(.A(n7627), .B(n6530), .Y(n7782));
  AOI21X1 g6641(.A0(n7782), .A1(n7715), .B0(n7628), .Y(n7783));
  INVX1   g6642(.A(n7783), .Y(n7784));
  XOR2X1  g6643(.A(n7618), .B(n6602), .Y(n7785));
  AOI21X1 g6644(.A0(n7622), .A1(n6567), .B0(n7785), .Y(n7786));
  OAI21X1 g6645(.A0(n7784), .A1(n7623), .B0(n7786), .Y(n7787));
  NAND2X1 g6646(.A(n7784), .B(n7629), .Y(n7788));
  NAND3X1 g6647(.A(n7788), .B(n7624), .C(n7625), .Y(n7789));
  AOI21X1 g6648(.A0(n7789), .A1(n7787), .B0(n7727), .Y(n7790));
  AOI22X1 g6649(.A0(P2_ADDR_REG_16__SCAN_IN), .A1(n7460), .B0(P2_REG3_REG_16__SCAN_IN), .B1(P2_U3151), .Y(n7791));
  OAI21X1 g6650(.A0(n7729), .A1(n6601), .B0(n7791), .Y(n7792));
  NOR4X1  g6651(.A(n7790), .B(n7781), .C(n7779), .D(n7792), .Y(n7793));
  OAI21X1 g6652(.A0(n7778), .A1(n7736), .B0(n7793), .Y(P2_U3198));
  XOR2X1  g6653(.A(n6566), .B(P2_REG2_REG_15__SCAN_IN), .Y(n7795));
  XOR2X1  g6654(.A(n7795), .B(n7506), .Y(n7796));
  XOR2X1  g6655(.A(n6566), .B(P2_REG1_REG_15__SCAN_IN), .Y(n7797));
  XOR2X1  g6656(.A(n7797), .B(n7581), .Y(n7798));
  OAI22X1 g6657(.A0(n7596), .A1(n6566), .B0(n5867), .B1(n7798), .Y(n7799));
  AOI21X1 g6658(.A0(n7796), .A1(n7520), .B0(n7799), .Y(n7800));
  NAND2X1 g6659(.A(n7796), .B(n7604), .Y(n7801));
  NAND2X1 g6660(.A(n7730), .B(n6567), .Y(n7802));
  AOI22X1 g6661(.A0(P2_ADDR_REG_15__SCAN_IN), .A1(n7460), .B0(P2_REG3_REG_15__SCAN_IN), .B1(P2_U3151), .Y(n7803));
  NAND3X1 g6662(.A(n7803), .B(n7802), .C(n7801), .Y(n7804));
  XOR2X1  g6663(.A(n7622), .B(n6567), .Y(n7805));
  XOR2X1  g6664(.A(n7805), .B(n7783), .Y(n7806));
  OAI22X1 g6665(.A0(n7798), .A1(n7602), .B0(n7727), .B1(n7806), .Y(n7807));
  NOR2X1  g6666(.A(n7807), .B(n7804), .Y(n7808));
  OAI21X1 g6667(.A0(n7800), .A1(n7736), .B0(n7808), .Y(P2_U3197));
  XOR2X1  g6668(.A(n6529), .B(P2_REG2_REG_14__SCAN_IN), .Y(n7810));
  XOR2X1  g6669(.A(n7810), .B(n7505), .Y(n7811));
  NOR2X1  g6670(.A(n7811), .B(n7521), .Y(n7812));
  XOR2X1  g6671(.A(n6529), .B(P2_REG1_REG_14__SCAN_IN), .Y(n7813));
  XOR2X1  g6672(.A(n7813), .B(n7579), .Y(n7814));
  OAI22X1 g6673(.A0(n7596), .A1(n6529), .B0(n5867), .B1(n7814), .Y(n7815));
  OAI21X1 g6674(.A0(n7815), .A1(n7812), .B0(n7461), .Y(n7816));
  NOR2X1  g6675(.A(n7811), .B(n7605), .Y(n7817));
  AOI22X1 g6676(.A0(P2_ADDR_REG_14__SCAN_IN), .A1(n7460), .B0(P2_REG3_REG_14__SCAN_IN), .B1(P2_U3151), .Y(n7818));
  OAI21X1 g6677(.A0(n7729), .A1(n6529), .B0(n7818), .Y(n7819));
  XOR2X1  g6678(.A(n7627), .B(n6529), .Y(n7820));
  XOR2X1  g6679(.A(n7820), .B(n7715), .Y(n7821));
  OAI22X1 g6680(.A0(n7814), .A1(n7602), .B0(n7727), .B1(n7821), .Y(n7822));
  NOR3X1  g6681(.A(n7822), .B(n7819), .C(n7817), .Y(n7823));
  NAND2X1 g6682(.A(n7823), .B(n7816), .Y(P2_U3196));
  XOR2X1  g6683(.A(n6482), .B(P2_REG2_REG_13__SCAN_IN), .Y(n7825));
  XOR2X1  g6684(.A(n7825), .B(n7504), .Y(n7826));
  XOR2X1  g6685(.A(n6482), .B(n7632), .Y(n7827));
  XOR2X1  g6686(.A(n7827), .B(n7578), .Y(n7828));
  OAI22X1 g6687(.A0(n7596), .A1(n6482), .B0(n5867), .B1(n7828), .Y(n7829));
  AOI21X1 g6688(.A0(n7826), .A1(n7520), .B0(n7829), .Y(n7830));
  NAND2X1 g6689(.A(n7826), .B(n7604), .Y(n7831));
  NAND2X1 g6690(.A(n7730), .B(n6483), .Y(n7832));
  AOI22X1 g6691(.A0(P2_ADDR_REG_13__SCAN_IN), .A1(n7460), .B0(P2_REG3_REG_13__SCAN_IN), .B1(P2_U3151), .Y(n7833));
  NAND3X1 g6692(.A(n7833), .B(n7832), .C(n7831), .Y(n7834));
  XOR2X1  g6693(.A(n7634), .B(n6482), .Y(n7835));
  XOR2X1  g6694(.A(n7835), .B(n7713), .Y(n7836));
  OAI22X1 g6695(.A0(n7828), .A1(n7602), .B0(n7727), .B1(n7836), .Y(n7837));
  NOR2X1  g6696(.A(n7837), .B(n7834), .Y(n7838));
  OAI21X1 g6697(.A0(n7830), .A1(n7736), .B0(n7838), .Y(P2_U3195));
  XOR2X1  g6698(.A(n6438), .B(P2_REG2_REG_12__SCAN_IN), .Y(n7840));
  XOR2X1  g6699(.A(n7840), .B(n7503), .Y(n7841));
  NOR2X1  g6700(.A(n7841), .B(n7521), .Y(n7842));
  XOR2X1  g6701(.A(n6438), .B(P2_REG1_REG_12__SCAN_IN), .Y(n7843));
  XOR2X1  g6702(.A(n7843), .B(n7577), .Y(n7844));
  OAI22X1 g6703(.A0(n7596), .A1(n6438), .B0(n5867), .B1(n7844), .Y(n7845));
  OAI21X1 g6704(.A0(n7845), .A1(n7842), .B0(n7461), .Y(n7846));
  NOR2X1  g6705(.A(n7841), .B(n7605), .Y(n7847));
  AOI22X1 g6706(.A0(P2_ADDR_REG_12__SCAN_IN), .A1(n7460), .B0(P2_REG3_REG_12__SCAN_IN), .B1(P2_U3151), .Y(n7848));
  OAI21X1 g6707(.A0(n7729), .A1(n6438), .B0(n7848), .Y(n7849));
  XOR2X1  g6708(.A(n7637), .B(n6438), .Y(n7850));
  XOR2X1  g6709(.A(n7850), .B(n7711), .Y(n7851));
  OAI22X1 g6710(.A0(n7844), .A1(n7602), .B0(n7727), .B1(n7851), .Y(n7852));
  NOR3X1  g6711(.A(n7852), .B(n7849), .C(n7847), .Y(n7853));
  NAND2X1 g6712(.A(n7853), .B(n7846), .Y(P2_U3194));
  INVX1   g6713(.A(n7646), .Y(n7855));
  NOR2X1  g6714(.A(n7651), .B(n6299), .Y(n7856));
  AOI21X1 g6715(.A0(n7709), .A1(n7708), .B0(n7856), .Y(n7857));
  OAI22X1 g6716(.A0(n7652), .A1(n6343), .B0(n7643), .B1(n7647), .Y(n7858));
  AOI21X1 g6717(.A0(n7857), .A1(n7855), .B0(n7858), .Y(n7859));
  NOR2X1  g6718(.A(n7857), .B(n7653), .Y(n7860));
  NOR3X1  g6719(.A(n7860), .B(n7649), .C(n7643), .Y(n7861));
  OAI21X1 g6720(.A0(n7861), .A1(n7859), .B0(n7761), .Y(n7862));
  XOR2X1  g6721(.A(n6390), .B(P2_REG2_REG_11__SCAN_IN), .Y(n7863));
  XOR2X1  g6722(.A(n7863), .B(n7502), .Y(n7864));
  NAND2X1 g6723(.A(n7864), .B(n7520), .Y(n7865));
  XOR2X1  g6724(.A(n6390), .B(P2_REG1_REG_11__SCAN_IN), .Y(n7866));
  XOR2X1  g6725(.A(n7866), .B(n7576), .Y(n7867));
  AOI22X1 g6726(.A0(n5915), .A1(n6391), .B0(n5914), .B1(n7867), .Y(n7868));
  NAND2X1 g6727(.A(n7868), .B(n7865), .Y(n7869));
  NAND2X1 g6728(.A(n7869), .B(n7461), .Y(n7870));
  NAND2X1 g6729(.A(n7867), .B(n7601), .Y(n7871));
  AOI22X1 g6730(.A0(P2_ADDR_REG_11__SCAN_IN), .A1(n7460), .B0(P2_REG3_REG_11__SCAN_IN), .B1(P2_U3151), .Y(n7872));
  OAI21X1 g6731(.A0(n7729), .A1(n6390), .B0(n7872), .Y(n7873));
  AOI21X1 g6732(.A0(n7864), .A1(n7604), .B0(n7873), .Y(n7874));
  NAND4X1 g6733(.A(n7871), .B(n7870), .C(n7862), .D(n7874), .Y(P2_U3193));
  XOR2X1  g6734(.A(n7645), .B(n6344), .Y(n7876));
  XOR2X1  g6735(.A(n7876), .B(n7857), .Y(n7877));
  XOR2X1  g6736(.A(n6343), .B(P2_REG2_REG_10__SCAN_IN), .Y(n7878));
  XOR2X1  g6737(.A(n7878), .B(n7501), .Y(n7879));
  NOR2X1  g6738(.A(n7879), .B(n7521), .Y(n7880));
  XOR2X1  g6739(.A(n6343), .B(P2_REG1_REG_10__SCAN_IN), .Y(n7881));
  XOR2X1  g6740(.A(n7881), .B(n7575), .Y(n7882));
  OAI22X1 g6741(.A0(n7596), .A1(n6343), .B0(n5867), .B1(n7882), .Y(n7883));
  NOR2X1  g6742(.A(n7883), .B(n7880), .Y(n7884));
  NOR2X1  g6743(.A(n7884), .B(n7736), .Y(n7885));
  NOR2X1  g6744(.A(n7882), .B(n7602), .Y(n7886));
  NOR2X1  g6745(.A(n7879), .B(n7605), .Y(n7887));
  AOI22X1 g6746(.A0(P2_ADDR_REG_10__SCAN_IN), .A1(n7460), .B0(P2_REG3_REG_10__SCAN_IN), .B1(P2_U3151), .Y(n7888));
  OAI21X1 g6747(.A0(n7729), .A1(n6343), .B0(n7888), .Y(n7889));
  NOR4X1  g6748(.A(n7887), .B(n7886), .C(n7885), .D(n7889), .Y(n7890));
  OAI21X1 g6749(.A0(n7877), .A1(n7727), .B0(n7890), .Y(P2_U3192));
  XOR2X1  g6750(.A(n7651), .B(n6298), .Y(n7892));
  XOR2X1  g6751(.A(n7892), .B(n7708), .Y(n7893));
  XOR2X1  g6752(.A(n6298), .B(P2_REG2_REG_9__SCAN_IN), .Y(n7894));
  XOR2X1  g6753(.A(n7894), .B(n7500), .Y(n7895));
  XOR2X1  g6754(.A(n6298), .B(P2_REG1_REG_9__SCAN_IN), .Y(n7896));
  XOR2X1  g6755(.A(n7896), .B(n7573), .Y(n7897));
  OAI22X1 g6756(.A0(n7596), .A1(n6298), .B0(n5867), .B1(n7897), .Y(n7898));
  AOI21X1 g6757(.A0(n7895), .A1(n7520), .B0(n7898), .Y(n7899));
  NOR2X1  g6758(.A(n7899), .B(n7736), .Y(n7900));
  NOR2X1  g6759(.A(n7897), .B(n7602), .Y(n7901));
  INVX1   g6760(.A(n7895), .Y(n7902));
  NOR2X1  g6761(.A(n7902), .B(n7605), .Y(n7903));
  AOI22X1 g6762(.A0(P2_ADDR_REG_9__SCAN_IN), .A1(n7460), .B0(P2_REG3_REG_9__SCAN_IN), .B1(P2_U3151), .Y(n7904));
  OAI21X1 g6763(.A0(n7729), .A1(n6298), .B0(n7904), .Y(n7905));
  NOR4X1  g6764(.A(n7903), .B(n7901), .C(n7900), .D(n7905), .Y(n7906));
  OAI21X1 g6765(.A0(n7893), .A1(n7727), .B0(n7906), .Y(P2_U3191));
  NOR2X1  g6766(.A(n7703), .B(n6208), .Y(n7908));
  AOI21X1 g6767(.A0(n7703), .A1(n6208), .B0(n7695), .Y(n7909));
  XOR2X1  g6768(.A(n7698), .B(n6252), .Y(n7910));
  NOR3X1  g6769(.A(n7910), .B(n7909), .C(n7908), .Y(n7911));
  AOI21X1 g6770(.A0(n7694), .A1(n7673), .B0(n7908), .Y(n7912));
  OAI21X1 g6771(.A0(n7702), .A1(n6209), .B0(n7910), .Y(n7913));
  NOR2X1  g6772(.A(n7913), .B(n7912), .Y(n7914));
  OAI21X1 g6773(.A0(n7914), .A1(n7911), .B0(n7761), .Y(n7915));
  XOR2X1  g6774(.A(n6251), .B(P2_REG2_REG_8__SCAN_IN), .Y(n7916));
  XOR2X1  g6775(.A(n7916), .B(n7499), .Y(n7917));
  NOR2X1  g6776(.A(n7917), .B(n7521), .Y(n7918));
  XOR2X1  g6777(.A(n6251), .B(P2_REG1_REG_8__SCAN_IN), .Y(n7919));
  XOR2X1  g6778(.A(n7919), .B(n7571), .Y(n7920));
  OAI22X1 g6779(.A0(n7596), .A1(n6251), .B0(n5867), .B1(n7920), .Y(n7921));
  OAI21X1 g6780(.A0(n7921), .A1(n7918), .B0(n7461), .Y(n7922));
  AOI22X1 g6781(.A0(P2_ADDR_REG_8__SCAN_IN), .A1(n7460), .B0(P2_REG3_REG_8__SCAN_IN), .B1(P2_U3151), .Y(n7923));
  OAI21X1 g6782(.A0(n7729), .A1(n6251), .B0(n7923), .Y(n7924));
  OAI22X1 g6783(.A0(n7917), .A1(n7605), .B0(n7602), .B1(n7920), .Y(n7925));
  NOR2X1  g6784(.A(n7925), .B(n7924), .Y(n7926));
  NAND3X1 g6785(.A(n7926), .B(n7922), .C(n7915), .Y(P2_U3190));
  XOR2X1  g6786(.A(n7702), .B(n6209), .Y(n7928));
  XOR2X1  g6787(.A(n7928), .B(n7695), .Y(n7929));
  NAND2X1 g6788(.A(n7929), .B(n7761), .Y(n7930));
  NOR3X1  g6789(.A(n7525), .B(n6208), .C(n7596), .Y(n7931));
  XOR2X1  g6790(.A(n6208), .B(n7700), .Y(n7932));
  XOR2X1  g6791(.A(n7932), .B(n7570), .Y(n7933));
  XOR2X1  g6792(.A(n6209), .B(P2_REG2_REG_7__SCAN_IN), .Y(n7934));
  XOR2X1  g6793(.A(n7934), .B(n7498), .Y(n7935));
  OAI22X1 g6794(.A0(n7933), .A1(n5867), .B0(n7521), .B1(n7935), .Y(n7936));
  OAI21X1 g6795(.A0(n7936), .A1(n7931), .B0(n7461), .Y(n7937));
  NOR2X1  g6796(.A(n7729), .B(n6208), .Y(n7938));
  NOR2X1  g6797(.A(n7933), .B(n7602), .Y(n7939));
  AOI22X1 g6798(.A0(P2_ADDR_REG_7__SCAN_IN), .A1(n7460), .B0(P2_REG3_REG_7__SCAN_IN), .B1(P2_U3151), .Y(n7940));
  OAI21X1 g6799(.A0(n7935), .A1(n7605), .B0(n7940), .Y(n7941));
  NOR3X1  g6800(.A(n7941), .B(n7939), .C(n7938), .Y(n7942));
  NAND3X1 g6801(.A(n7942), .B(n7937), .C(n7930), .Y(P2_U3189));
  NOR2X1  g6802(.A(n7669), .B(n6065), .Y(n7944));
  AOI21X1 g6803(.A0(n7693), .A1(n7692), .B0(n7944), .Y(n7945));
  OAI21X1 g6804(.A0(n7664), .A1(n7662), .B0(n7945), .Y(n7946));
  XOR2X1  g6805(.A(n7658), .B(n6159), .Y(n7947));
  AOI21X1 g6806(.A0(n7664), .A1(n7662), .B0(n7947), .Y(n7948));
  NOR2X1  g6807(.A(n7945), .B(n7671), .Y(n7949));
  NOR3X1  g6808(.A(n7949), .B(n7667), .C(n7660), .Y(n7950));
  AOI21X1 g6809(.A0(n7948), .A1(n7946), .B0(n7950), .Y(n7951));
  XOR2X1  g6810(.A(n6158), .B(n7550), .Y(n7952));
  XOR2X1  g6811(.A(n7952), .B(n7569), .Y(n7953));
  XOR2X1  g6812(.A(n6158), .B(n7296), .Y(n7954));
  XOR2X1  g6813(.A(n7954), .B(n7497), .Y(n7955));
  AOI22X1 g6814(.A0(n7953), .A1(n5914), .B0(n7520), .B1(n7955), .Y(n7956));
  OAI21X1 g6815(.A0(n7596), .A1(n6158), .B0(n7956), .Y(n7957));
  NAND2X1 g6816(.A(n7955), .B(n7604), .Y(n7958));
  AOI22X1 g6817(.A0(P2_ADDR_REG_6__SCAN_IN), .A1(n7460), .B0(P2_REG3_REG_6__SCAN_IN), .B1(P2_U3151), .Y(n7959));
  NAND2X1 g6818(.A(n7959), .B(n7958), .Y(n7960));
  AOI21X1 g6819(.A0(n7953), .A1(n7601), .B0(n7960), .Y(n7961));
  OAI21X1 g6820(.A0(n7729), .A1(n6158), .B0(n7961), .Y(n7962));
  AOI21X1 g6821(.A0(n7957), .A1(n7461), .B0(n7962), .Y(n7963));
  OAI21X1 g6822(.A0(n7951), .A1(n7727), .B0(n7963), .Y(P2_U3188));
  XOR2X1  g6823(.A(n7664), .B(n7662), .Y(n7965));
  XOR2X1  g6824(.A(n7965), .B(n7945), .Y(n7966));
  NAND3X1 g6825(.A(n7524), .B(n7662), .C(n5915), .Y(n7967));
  XOR2X1  g6826(.A(n6117), .B(P2_REG1_REG_5__SCAN_IN), .Y(n7968));
  XOR2X1  g6827(.A(n7968), .B(n7568), .Y(n7969));
  XOR2X1  g6828(.A(n6117), .B(P2_REG2_REG_5__SCAN_IN), .Y(n7970));
  XOR2X1  g6829(.A(n7970), .B(n7496), .Y(n7971));
  AOI22X1 g6830(.A0(n7969), .A1(n5914), .B0(n7520), .B1(n7971), .Y(n7972));
  AOI21X1 g6831(.A0(n7972), .A1(n7967), .B0(n7736), .Y(n7973));
  NOR2X1  g6832(.A(n7729), .B(n6117), .Y(n7974));
  NAND2X1 g6833(.A(n7969), .B(n7601), .Y(n7975));
  NAND2X1 g6834(.A(n7971), .B(n7604), .Y(n7976));
  AOI22X1 g6835(.A0(P2_ADDR_REG_5__SCAN_IN), .A1(n7460), .B0(P2_REG3_REG_5__SCAN_IN), .B1(P2_U3151), .Y(n7977));
  NAND3X1 g6836(.A(n7977), .B(n7976), .C(n7975), .Y(n7978));
  NOR3X1  g6837(.A(n7978), .B(n7974), .C(n7973), .Y(n7979));
  OAI21X1 g6838(.A0(n7966), .A1(n7727), .B0(n7979), .Y(P2_U3187));
  NOR3X1  g6839(.A(n7525), .B(n6064), .C(n7596), .Y(n7981));
  XOR2X1  g6840(.A(n6064), .B(P2_REG1_REG_4__SCAN_IN), .Y(n7982));
  XOR2X1  g6841(.A(n7982), .B(n7567), .Y(n7983));
  XOR2X1  g6842(.A(n6064), .B(P2_REG2_REG_4__SCAN_IN), .Y(n7984));
  XOR2X1  g6843(.A(n7984), .B(n7495), .Y(n7985));
  OAI22X1 g6844(.A0(n7983), .A1(n5867), .B0(n7521), .B1(n7985), .Y(n7986));
  OAI21X1 g6845(.A0(n7986), .A1(n7981), .B0(n7461), .Y(n7987));
  XOR2X1  g6846(.A(n7669), .B(n6065), .Y(n7988));
  XOR2X1  g6847(.A(n7988), .B(n7692), .Y(n7989));
  NAND2X1 g6848(.A(n7989), .B(n7761), .Y(n7990));
  NOR2X1  g6849(.A(n7729), .B(n6064), .Y(n7991));
  NOR2X1  g6850(.A(n7983), .B(n7602), .Y(n7992));
  AOI22X1 g6851(.A0(P2_ADDR_REG_4__SCAN_IN), .A1(n7460), .B0(P2_REG3_REG_4__SCAN_IN), .B1(P2_U3151), .Y(n7993));
  OAI21X1 g6852(.A0(n7985), .A1(n7605), .B0(n7993), .Y(n7994));
  NOR3X1  g6853(.A(n7994), .B(n7992), .C(n7991), .Y(n7995));
  NAND3X1 g6854(.A(n7995), .B(n7990), .C(n7987), .Y(P2_U3186));
  NOR3X1  g6855(.A(n7525), .B(n6020), .C(n7596), .Y(n7997));
  NOR2X1  g6856(.A(n5979), .B(n7561), .Y(n7998));
  NOR2X1  g6857(.A(n7564), .B(n7563), .Y(n7999));
  OAI21X1 g6858(.A0(n7999), .A1(n7998), .B0(n7560), .Y(n8000));
  XOR2X1  g6859(.A(n6020), .B(n7558), .Y(n8001));
  XOR2X1  g6860(.A(n8001), .B(n8000), .Y(n8002));
  XOR2X1  g6861(.A(n6020), .B(P2_REG2_REG_3__SCAN_IN), .Y(n8003));
  XOR2X1  g6862(.A(n8003), .B(n7493), .Y(n8004));
  OAI22X1 g6863(.A0(n8002), .A1(n5867), .B0(n7521), .B1(n8004), .Y(n8005));
  OAI21X1 g6864(.A0(n8005), .A1(n7997), .B0(n7461), .Y(n8006));
  INVX1   g6865(.A(n7686), .Y(n8007));
  NOR2X1  g6866(.A(n8007), .B(n5978), .Y(n8008));
  AOI21X1 g6867(.A0(n8007), .A1(n5978), .B0(n7682), .Y(n8009));
  XOR2X1  g6868(.A(n7684), .B(n6021), .Y(n8010));
  NOR3X1  g6869(.A(n8010), .B(n8009), .C(n8008), .Y(n8011));
  INVX1   g6870(.A(n8008), .Y(n8012));
  OAI21X1 g6871(.A0(n7686), .A1(n5979), .B0(n8010), .Y(n8013));
  AOI21X1 g6872(.A0(n8012), .A1(n7682), .B0(n8013), .Y(n8014));
  OAI21X1 g6873(.A0(n8014), .A1(n8011), .B0(n7761), .Y(n8015));
  NOR2X1  g6874(.A(n7729), .B(n6020), .Y(n8016));
  NOR2X1  g6875(.A(n8002), .B(n7602), .Y(n8017));
  AOI22X1 g6876(.A0(P2_ADDR_REG_3__SCAN_IN), .A1(n7460), .B0(P2_REG3_REG_3__SCAN_IN), .B1(P2_U3151), .Y(n8018));
  OAI21X1 g6877(.A0(n8004), .A1(n7605), .B0(n8018), .Y(n8019));
  NOR3X1  g6878(.A(n8019), .B(n8017), .C(n8016), .Y(n8020));
  NAND3X1 g6879(.A(n8020), .B(n8015), .C(n8006), .Y(P2_U3185));
  NOR3X1  g6880(.A(n7525), .B(n5978), .C(n7596), .Y(n8022));
  XOR2X1  g6881(.A(n5978), .B(P2_REG1_REG_2__SCAN_IN), .Y(n8023));
  XOR2X1  g6882(.A(n8023), .B(n7999), .Y(n8024));
  XOR2X1  g6883(.A(n5978), .B(P2_REG2_REG_2__SCAN_IN), .Y(n8025));
  XOR2X1  g6884(.A(n8025), .B(n7491), .Y(n8026));
  OAI22X1 g6885(.A0(n8024), .A1(n5867), .B0(n7521), .B1(n8026), .Y(n8027));
  OAI21X1 g6886(.A0(n8027), .A1(n8022), .B0(n7461), .Y(n8028));
  NOR2X1  g6887(.A(n8024), .B(n7602), .Y(n8029));
  AOI22X1 g6888(.A0(P2_ADDR_REG_2__SCAN_IN), .A1(n7460), .B0(P2_REG3_REG_2__SCAN_IN), .B1(P2_U3151), .Y(n8030));
  OAI21X1 g6889(.A0(n8026), .A1(n7605), .B0(n8030), .Y(n8031));
  NOR2X1  g6890(.A(n8031), .B(n8029), .Y(n8032));
  XOR2X1  g6891(.A(n7686), .B(n5979), .Y(n8033));
  XOR2X1  g6892(.A(n8033), .B(n7682), .Y(n8034));
  AOI22X1 g6893(.A0(n7730), .A1(n5979), .B0(n7761), .B1(n8034), .Y(n8035));
  NAND3X1 g6894(.A(n8035), .B(n8032), .C(n8028), .Y(P2_U3184));
  NOR3X1  g6895(.A(n7525), .B(n5936), .C(n7596), .Y(n8037));
  XOR2X1  g6896(.A(n7562), .B(n7169), .Y(n8038));
  XOR2X1  g6897(.A(n8038), .B(n5937), .Y(n8039));
  XOR2X1  g6898(.A(n7488), .B(n7259), .Y(n8040));
  XOR2X1  g6899(.A(n8040), .B(n5937), .Y(n8041));
  OAI22X1 g6900(.A0(n8039), .A1(n5867), .B0(n7521), .B1(n8041), .Y(n8042));
  OAI21X1 g6901(.A0(n8042), .A1(n8037), .B0(n7461), .Y(n8043));
  NOR2X1  g6902(.A(n7729), .B(n5936), .Y(n8044));
  NOR2X1  g6903(.A(n8039), .B(n7602), .Y(n8045));
  NOR2X1  g6904(.A(n8041), .B(n7605), .Y(n8046));
  XOR2X1  g6905(.A(n7675), .B(n5936), .Y(n8047));
  XOR2X1  g6906(.A(n8047), .B(n7678), .Y(n8048));
  AOI22X1 g6907(.A0(P2_ADDR_REG_1__SCAN_IN), .A1(n7460), .B0(P2_REG3_REG_1__SCAN_IN), .B1(P2_U3151), .Y(n8049));
  OAI21X1 g6908(.A0(n8048), .A1(n7727), .B0(n8049), .Y(n8050));
  NOR4X1  g6909(.A(n8046), .B(n8045), .C(n8044), .D(n8050), .Y(n8051));
  NAND2X1 g6910(.A(n8051), .B(n8043), .Y(P2_U3183));
  NOR3X1  g6911(.A(n7525), .B(n5873), .C(n7596), .Y(n8053));
  XOR2X1  g6912(.A(n5873), .B(P2_REG1_REG_0__SCAN_IN), .Y(n8054));
  XOR2X1  g6913(.A(n5873), .B(P2_REG2_REG_0__SCAN_IN), .Y(n8055));
  OAI22X1 g6914(.A0(n8054), .A1(n5867), .B0(n7521), .B1(n8055), .Y(n8056));
  OAI21X1 g6915(.A0(n8056), .A1(n8053), .B0(n7461), .Y(n8057));
  NAND2X1 g6916(.A(n7730), .B(n5876), .Y(n8058));
  NOR2X1  g6917(.A(n8054), .B(n7602), .Y(n8059));
  NOR2X1  g6918(.A(n8055), .B(n7605), .Y(n8060));
  INVX1   g6919(.A(P2_ADDR_REG_0__SCAN_IN), .Y(n8061));
  NOR2X1  g6920(.A(n7459), .B(n8061), .Y(n8062));
  INVX1   g6921(.A(P2_REG3_REG_0__SCAN_IN), .Y(n8063));
  XOR2X1  g6922(.A(n7677), .B(n5876), .Y(n8064));
  OAI22X1 g6923(.A0(n7727), .A1(n8064), .B0(n8063), .B1(P2_STATE_REG_SCAN_IN), .Y(n8065));
  NOR4X1  g6924(.A(n8062), .B(n8060), .C(n8059), .D(n8065), .Y(n8066));
  NAND3X1 g6925(.A(n8066), .B(n8058), .C(n8057), .Y(P2_U3182));
  NAND2X1 g6926(.A(n7725), .B(P2_DATAO_REG_0__SCAN_IN), .Y(n8068));
  OAI21X1 g6927(.A0(n7725), .A1(n5994), .B0(n8068), .Y(P2_U3491));
  NAND2X1 g6928(.A(n7725), .B(P2_DATAO_REG_1__SCAN_IN), .Y(n8070));
  OAI21X1 g6929(.A0(n7725), .A1(n5925), .B0(n8070), .Y(P2_U3492));
  NAND2X1 g6930(.A(n7725), .B(P2_DATAO_REG_2__SCAN_IN), .Y(n8072));
  OAI21X1 g6931(.A0(n7725), .A1(n5965), .B0(n8072), .Y(P2_U3493));
  NAND2X1 g6932(.A(n7725), .B(P2_DATAO_REG_3__SCAN_IN), .Y(n8074));
  OAI21X1 g6933(.A0(n7725), .A1(n6079), .B0(n8074), .Y(P2_U3494));
  NAND2X1 g6934(.A(n7725), .B(P2_DATAO_REG_4__SCAN_IN), .Y(n8076));
  OAI21X1 g6935(.A0(n7725), .A1(n6104), .B0(n8076), .Y(P2_U3495));
  NAND2X1 g6936(.A(n7725), .B(P2_DATAO_REG_5__SCAN_IN), .Y(n8078));
  OAI21X1 g6937(.A0(n7725), .A1(n6115), .B0(n8078), .Y(P2_U3496));
  NAND2X1 g6938(.A(n7725), .B(P2_DATAO_REG_6__SCAN_IN), .Y(n8080));
  OAI21X1 g6939(.A0(n7725), .A1(n6156), .B0(n8080), .Y(P2_U3497));
  NAND2X1 g6940(.A(n7725), .B(P2_DATAO_REG_7__SCAN_IN), .Y(n8082));
  OAI21X1 g6941(.A0(n7725), .A1(n6206), .B0(n8082), .Y(P2_U3498));
  NAND2X1 g6942(.A(n7725), .B(P2_DATAO_REG_8__SCAN_IN), .Y(n8084));
  OAI21X1 g6943(.A0(n7725), .A1(n6249), .B0(n8084), .Y(P2_U3499));
  NAND2X1 g6944(.A(n7725), .B(P2_DATAO_REG_9__SCAN_IN), .Y(n8086));
  OAI21X1 g6945(.A0(n7725), .A1(n6296), .B0(n8086), .Y(P2_U3500));
  NAND2X1 g6946(.A(n7725), .B(P2_DATAO_REG_10__SCAN_IN), .Y(n8088));
  OAI21X1 g6947(.A0(n7725), .A1(n6333), .B0(n8088), .Y(P2_U3501));
  NAND2X1 g6948(.A(n7725), .B(P2_DATAO_REG_11__SCAN_IN), .Y(n8090));
  OAI21X1 g6949(.A0(n7725), .A1(n6412), .B0(n8090), .Y(P2_U3502));
  NAND2X1 g6950(.A(n7725), .B(P2_DATAO_REG_12__SCAN_IN), .Y(n8092));
  OAI21X1 g6951(.A0(n7725), .A1(n6436), .B0(n8092), .Y(P2_U3503));
  NAND2X1 g6952(.A(n7725), .B(P2_DATAO_REG_13__SCAN_IN), .Y(n8094));
  OAI21X1 g6953(.A0(n7725), .A1(n6480), .B0(n8094), .Y(P2_U3504));
  NAND2X1 g6954(.A(n7725), .B(P2_DATAO_REG_14__SCAN_IN), .Y(n8096));
  OAI21X1 g6955(.A0(n7725), .A1(n6527), .B0(n8096), .Y(P2_U3505));
  NAND2X1 g6956(.A(n7725), .B(P2_DATAO_REG_15__SCAN_IN), .Y(n8098));
  OAI21X1 g6957(.A0(n7725), .A1(n6558), .B0(n8098), .Y(P2_U3506));
  NAND2X1 g6958(.A(n7725), .B(P2_DATAO_REG_16__SCAN_IN), .Y(n8100));
  OAI21X1 g6959(.A0(n7725), .A1(n6599), .B0(n8100), .Y(P2_U3507));
  NAND2X1 g6960(.A(n7725), .B(P2_DATAO_REG_17__SCAN_IN), .Y(n8102));
  OAI21X1 g6961(.A0(n7725), .A1(n6691), .B0(n8102), .Y(P2_U3508));
  NAND2X1 g6962(.A(n7725), .B(P2_DATAO_REG_18__SCAN_IN), .Y(n8104));
  OAI21X1 g6963(.A0(n7725), .A1(n6702), .B0(n8104), .Y(P2_U3509));
  NAND2X1 g6964(.A(n7725), .B(P2_DATAO_REG_19__SCAN_IN), .Y(n8106));
  OAI21X1 g6965(.A0(n7725), .A1(n6735), .B0(n8106), .Y(P2_U3510));
  NAND2X1 g6966(.A(n7725), .B(P2_DATAO_REG_20__SCAN_IN), .Y(n8108));
  OAI21X1 g6967(.A0(n7725), .A1(n6773), .B0(n8108), .Y(P2_U3511));
  NAND2X1 g6968(.A(n7725), .B(P2_DATAO_REG_21__SCAN_IN), .Y(n8110));
  OAI21X1 g6969(.A0(n7725), .A1(n6814), .B0(n8110), .Y(P2_U3512));
  NAND2X1 g6970(.A(n7725), .B(P2_DATAO_REG_22__SCAN_IN), .Y(n8112));
  OAI21X1 g6971(.A0(n7725), .A1(n6848), .B0(n8112), .Y(P2_U3513));
  NAND2X1 g6972(.A(n7725), .B(P2_DATAO_REG_23__SCAN_IN), .Y(n8114));
  OAI21X1 g6973(.A0(n7725), .A1(n6890), .B0(n8114), .Y(P2_U3514));
  NAND2X1 g6974(.A(n7725), .B(P2_DATAO_REG_24__SCAN_IN), .Y(n8116));
  OAI21X1 g6975(.A0(n7725), .A1(n6929), .B0(n8116), .Y(P2_U3515));
  NAND2X1 g6976(.A(n7725), .B(P2_DATAO_REG_25__SCAN_IN), .Y(n8118));
  OAI21X1 g6977(.A0(n7725), .A1(n6959), .B0(n8118), .Y(P2_U3516));
  NAND2X1 g6978(.A(n7725), .B(P2_DATAO_REG_26__SCAN_IN), .Y(n8120));
  OAI21X1 g6979(.A0(n7725), .A1(n6994), .B0(n8120), .Y(P2_U3517));
  NAND2X1 g6980(.A(n7725), .B(P2_DATAO_REG_27__SCAN_IN), .Y(n8122));
  OAI21X1 g6981(.A0(n7725), .A1(n7074), .B0(n8122), .Y(P2_U3518));
  NAND2X1 g6982(.A(n7725), .B(P2_DATAO_REG_28__SCAN_IN), .Y(n8124));
  OAI21X1 g6983(.A0(n7725), .A1(n7111), .B0(n8124), .Y(P2_U3519));
  NAND2X1 g6984(.A(n7725), .B(P2_DATAO_REG_29__SCAN_IN), .Y(n8126));
  OAI21X1 g6985(.A0(n7725), .A1(n7106), .B0(n8126), .Y(P2_U3520));
  INVX1   g6986(.A(n7131), .Y(n8128));
  NAND2X1 g6987(.A(n7725), .B(P2_DATAO_REG_30__SCAN_IN), .Y(n8129));
  OAI21X1 g6988(.A0(n7725), .A1(n8128), .B0(n8129), .Y(P2_U3521));
  NAND2X1 g6989(.A(n7725), .B(P2_DATAO_REG_31__SCAN_IN), .Y(n8131));
  OAI21X1 g6990(.A0(n7725), .A1(n7147), .B0(n8131), .Y(P2_U3522));
  INVX1   g6991(.A(n7132), .Y(n8134));
  NOR2X1  g6992(.A(n5853), .B(n5846), .Y(n8135));
  NOR2X1  g6993(.A(n5860), .B(n5846), .Y(n8136));
  NOR2X1  g6994(.A(n5844), .B(n5728), .Y(n8137));
  AOI22X1 g6995(.A0(n8136), .A1(n8137), .B0(n8135), .B1(n5847), .Y(n8138));
  INVX1   g6996(.A(n8138), .Y(n8139));
  AOI22X1 g6997(.A0(n8134), .A1(n7146), .B0(n7153), .B1(n8139), .Y(n8140));
  OAI22X1 g6998(.A0(n7132), .A1(n7453), .B0(n7147), .B1(n8138), .Y(n8141));
  XOR2X1  g6999(.A(n8141), .B(n8140), .Y(n8142));
  OAI22X1 g7000(.A0(n7132), .A1(n7448), .B0(n8128), .B1(n8138), .Y(n8143));
  AOI22X1 g7001(.A0(n7100), .A1(n8139), .B0(n7064), .B1(n5728), .Y(n8144));
  OAI21X1 g7002(.A0(n7132), .A1(n7114), .B0(n8144), .Y(n8145));
  AOI21X1 g7003(.A0(n8134), .A1(n7100), .B0(n5728), .Y(n8146));
  INVX1   g7004(.A(n8146), .Y(n8147));
  AOI21X1 g7005(.A0(n8139), .A1(n7107), .B0(n8147), .Y(n8148));
  AOI22X1 g7006(.A0(n8134), .A1(n7131), .B0(n7149), .B1(n8139), .Y(n8149));
  AOI22X1 g7007(.A0(n8148), .A1(n8145), .B0(n8143), .B1(n8149), .Y(n8150));
  AOI22X1 g7008(.A0(n7064), .A1(n8139), .B0(n7023), .B1(n5728), .Y(n8151));
  OAI21X1 g7009(.A0(n7132), .A1(n7071), .B0(n8151), .Y(n8152));
  AOI21X1 g7010(.A0(n8134), .A1(n7064), .B0(n5728), .Y(n8153));
  INVX1   g7011(.A(n8153), .Y(n8154));
  AOI21X1 g7012(.A0(n8139), .A1(n7093), .B0(n8154), .Y(n8155));
  AOI22X1 g7013(.A0(n6987), .A1(n8139), .B0(n6953), .B1(n5728), .Y(n8156));
  OAI21X1 g7014(.A0(n7132), .A1(n6996), .B0(n8156), .Y(n8157));
  INVX1   g7015(.A(n8157), .Y(n8158));
  AOI21X1 g7016(.A0(n8134), .A1(n6987), .B0(n5728), .Y(n8159));
  OAI21X1 g7017(.A0(n8138), .A1(n6996), .B0(n8159), .Y(n8160));
  AOI22X1 g7018(.A0(n7023), .A1(n8139), .B0(n6987), .B1(n5728), .Y(n8161));
  OAI21X1 g7019(.A0(n7132), .A1(n7034), .B0(n8161), .Y(n8162));
  INVX1   g7020(.A(n8162), .Y(n8163));
  AOI21X1 g7021(.A0(n8134), .A1(n7023), .B0(n5728), .Y(n8164));
  OAI21X1 g7022(.A0(n8138), .A1(n7034), .B0(n8164), .Y(n8165));
  OAI22X1 g7023(.A0(n8163), .A1(n8165), .B0(n8160), .B1(n8158), .Y(n8166));
  AOI21X1 g7024(.A0(n8155), .A1(n8152), .B0(n8166), .Y(n8167));
  NAND2X1 g7025(.A(n8134), .B(n6960), .Y(n8168));
  AOI22X1 g7026(.A0(n6953), .A1(n8139), .B0(n6916), .B1(n5728), .Y(n8169));
  NAND2X1 g7027(.A(n8169), .B(n8168), .Y(n8170));
  NAND2X1 g7028(.A(n8139), .B(n6960), .Y(n8171));
  AOI21X1 g7029(.A0(n8134), .A1(n6953), .B0(n5728), .Y(n8172));
  AOI21X1 g7030(.A0(n8172), .A1(n8171), .B0(n8170), .Y(n8173));
  NAND4X1 g7031(.A(n8167), .B(n8150), .C(n8142), .D(n8173), .Y(n8174));
  AOI22X1 g7032(.A0(n8134), .A1(n7153), .B0(n7146), .B1(n8139), .Y(n8175));
  XOR2X1  g7033(.A(n8175), .B(n8140), .Y(n8176));
  AOI22X1 g7034(.A0(n8134), .A1(n7149), .B0(n7131), .B1(n8139), .Y(n8177));
  INVX1   g7035(.A(n8144), .Y(n8178));
  AOI21X1 g7036(.A0(n8134), .A1(n7107), .B0(n8178), .Y(n8179));
  OAI21X1 g7037(.A0(n8138), .A1(n7114), .B0(n8146), .Y(n8180));
  OAI22X1 g7038(.A0(n7132), .A1(n8128), .B0(n7448), .B1(n8138), .Y(n8181));
  OAI22X1 g7039(.A0(n8180), .A1(n8179), .B0(n8177), .B1(n8181), .Y(n8182));
  NOR4X1  g7040(.A(n8152), .B(n8182), .C(n8176), .D(n8155), .Y(n8183));
  INVX1   g7041(.A(n8151), .Y(n8184));
  AOI21X1 g7042(.A0(n8134), .A1(n7093), .B0(n8184), .Y(n8185));
  OAI21X1 g7043(.A0(n8138), .A1(n7071), .B0(n8153), .Y(n8186));
  INVX1   g7044(.A(n8165), .Y(n8187));
  NOR2X1  g7045(.A(n8187), .B(n8162), .Y(n8188));
  OAI21X1 g7046(.A0(n8186), .A1(n8185), .B0(n8188), .Y(n8189));
  NOR3X1  g7047(.A(n8189), .B(n8182), .C(n8176), .Y(n8190));
  NOR2X1  g7048(.A(n8190), .B(n8183), .Y(n8191));
  NOR4X1  g7049(.A(n5844), .B(n5846), .C(n5729), .D(n5860), .Y(n8192));
  NOR2X1  g7050(.A(n8192), .B(n8141), .Y(n8193));
  NAND2X1 g7051(.A(n8192), .B(n8140), .Y(n8194));
  OAI21X1 g7052(.A0(n8175), .A1(n8140), .B0(n8194), .Y(n8195));
  NOR2X1  g7053(.A(n8195), .B(n8193), .Y(n8196));
  NAND2X1 g7054(.A(n8181), .B(n8177), .Y(n8197));
  NOR2X1  g7055(.A(n8148), .B(n8145), .Y(n8198));
  OAI21X1 g7056(.A0(n8181), .A1(n8177), .B0(n8198), .Y(n8199));
  AOI21X1 g7057(.A0(n8199), .A1(n8197), .B0(n8176), .Y(n8200));
  INVX1   g7058(.A(n8160), .Y(n8201));
  AOI22X1 g7059(.A0(n8162), .A1(n8187), .B0(n8201), .B1(n8157), .Y(n8202));
  OAI21X1 g7060(.A0(n8186), .A1(n8185), .B0(n8202), .Y(n8203));
  NAND2X1 g7061(.A(n8160), .B(n8158), .Y(n8204));
  NOR4X1  g7062(.A(n8203), .B(n8182), .C(n8176), .D(n8204), .Y(n8205));
  OAI21X1 g7063(.A0(n8138), .A1(n7046), .B0(n8172), .Y(n8206));
  AOI21X1 g7064(.A0(n8169), .A1(n8168), .B0(n8206), .Y(n8207));
  AOI21X1 g7065(.A0(n8134), .A1(n6916), .B0(n5728), .Y(n8208));
  INVX1   g7066(.A(n8208), .Y(n8209));
  AOI21X1 g7067(.A0(n8139), .A1(n6946), .B0(n8209), .Y(n8210));
  AOI22X1 g7068(.A0(n6916), .A1(n8139), .B0(n6878), .B1(n5728), .Y(n8211));
  OAI21X1 g7069(.A0(n7132), .A1(n6925), .B0(n8211), .Y(n8212));
  NOR2X1  g7070(.A(n8212), .B(n8210), .Y(n8213));
  AOI22X1 g7071(.A0(n6878), .A1(n8139), .B0(n6842), .B1(n5728), .Y(n8214));
  OAI21X1 g7072(.A0(n7132), .A1(n6886), .B0(n8214), .Y(n8215));
  AOI21X1 g7073(.A0(n8134), .A1(n6878), .B0(n5728), .Y(n8216));
  INVX1   g7074(.A(n8216), .Y(n8217));
  AOI21X1 g7075(.A0(n8139), .A1(n6911), .B0(n8217), .Y(n8218));
  NOR2X1  g7076(.A(n8218), .B(n8215), .Y(n8219));
  AOI22X1 g7077(.A0(n6842), .A1(n8139), .B0(n6806), .B1(n5728), .Y(n8220));
  INVX1   g7078(.A(n8220), .Y(n8221));
  AOI21X1 g7079(.A0(n8134), .A1(n6849), .B0(n8221), .Y(n8222));
  AOI21X1 g7080(.A0(n8134), .A1(n6842), .B0(n5728), .Y(n8223));
  OAI21X1 g7081(.A0(n8138), .A1(n6893), .B0(n8223), .Y(n8224));
  NAND2X1 g7082(.A(n8224), .B(n8222), .Y(n8225));
  INVX1   g7083(.A(n6815), .Y(n8226));
  AOI22X1 g7084(.A0(n6806), .A1(n8139), .B0(n6767), .B1(n5728), .Y(n8227));
  OAI21X1 g7085(.A0(n7132), .A1(n8226), .B0(n8227), .Y(n8228));
  AOI21X1 g7086(.A0(n8134), .A1(n6806), .B0(n5728), .Y(n8229));
  INVX1   g7087(.A(n8229), .Y(n8230));
  AOI21X1 g7088(.A0(n8139), .A1(n6815), .B0(n8230), .Y(n8231));
  AOI22X1 g7089(.A0(n6767), .A1(n8139), .B0(n6729), .B1(n5728), .Y(n8232));
  OAI21X1 g7090(.A0(n7132), .A1(n6824), .B0(n8232), .Y(n8233));
  OAI21X1 g7091(.A0(n7132), .A1(n6773), .B0(n5729), .Y(n8234));
  AOI21X1 g7092(.A0(n8139), .A1(n6774), .B0(n8234), .Y(n8235));
  AOI22X1 g7093(.A0(n8233), .A1(n8235), .B0(n8231), .B1(n8228), .Y(n8236));
  AOI22X1 g7094(.A0(n6729), .A1(n8139), .B0(n6684), .B1(n5728), .Y(n8237));
  OAI21X1 g7095(.A0(n7132), .A1(n6820), .B0(n8237), .Y(n8238));
  AOI21X1 g7096(.A0(n8134), .A1(n6729), .B0(n5728), .Y(n8239));
  OAI21X1 g7097(.A0(n8138), .A1(n6820), .B0(n8239), .Y(n8240));
  INVX1   g7098(.A(n8240), .Y(n8241));
  NOR2X1  g7099(.A(n8241), .B(n8238), .Y(n8242));
  NAND2X1 g7100(.A(n8242), .B(n8236), .Y(n8243));
  NAND2X1 g7101(.A(n8231), .B(n8228), .Y(n8244));
  NOR2X1  g7102(.A(n8235), .B(n8233), .Y(n8245));
  NOR2X1  g7103(.A(n8231), .B(n8228), .Y(n8246));
  AOI21X1 g7104(.A0(n8245), .A1(n8244), .B0(n8246), .Y(n8247));
  NAND3X1 g7105(.A(n8247), .B(n8243), .C(n8225), .Y(n8248));
  AOI22X1 g7106(.A0(n6684), .A1(n8139), .B0(n6645), .B1(n5728), .Y(n8249));
  OAI21X1 g7107(.A0(n7132), .A1(n6699), .B0(n8249), .Y(n8250));
  OAI21X1 g7108(.A0(n7132), .A1(n6702), .B0(n5729), .Y(n8251));
  AOI21X1 g7109(.A0(n8139), .A1(n6721), .B0(n8251), .Y(n8252));
  AOI22X1 g7110(.A0(n6645), .A1(n8139), .B0(n6593), .B1(n5728), .Y(n8253));
  OAI21X1 g7111(.A0(n7132), .A1(n6657), .B0(n8253), .Y(n8254));
  AOI21X1 g7112(.A0(n8134), .A1(n6645), .B0(n5728), .Y(n8255));
  OAI21X1 g7113(.A0(n8138), .A1(n6657), .B0(n8255), .Y(n8256));
  INVX1   g7114(.A(n8256), .Y(n8257));
  OAI22X1 g7115(.A0(n8254), .A1(n8257), .B0(n8252), .B1(n8250), .Y(n8258));
  INVX1   g7116(.A(n8258), .Y(n8259));
  AOI22X1 g7117(.A0(n6593), .A1(n8139), .B0(n6559), .B1(n5728), .Y(n8260));
  OAI21X1 g7118(.A0(n7132), .A1(n6623), .B0(n8260), .Y(n8261));
  OAI21X1 g7119(.A0(n7132), .A1(n6599), .B0(n5729), .Y(n8262));
  AOI21X1 g7120(.A0(n8139), .A1(n6604), .B0(n8262), .Y(n8263));
  NAND3X1 g7121(.A(n8263), .B(n8261), .C(n8259), .Y(n8264));
  NOR2X1  g7122(.A(n8252), .B(n8250), .Y(n8265));
  NAND2X1 g7123(.A(n8252), .B(n8250), .Y(n8266));
  NAND2X1 g7124(.A(n8257), .B(n8254), .Y(n8267));
  OAI21X1 g7125(.A0(n8267), .A1(n8265), .B0(n8266), .Y(n8268));
  AOI21X1 g7126(.A0(n8241), .A1(n8238), .B0(n8268), .Y(n8269));
  NAND3X1 g7127(.A(n8269), .B(n8264), .C(n8236), .Y(n8270));
  OAI21X1 g7128(.A0(n7132), .A1(n6527), .B0(n5729), .Y(n8271));
  AOI21X1 g7129(.A0(n8139), .A1(n6532), .B0(n8271), .Y(n8272));
  AOI22X1 g7130(.A0(n6516), .A1(n8139), .B0(n6470), .B1(n5728), .Y(n8273));
  OAI21X1 g7131(.A0(n7132), .A1(n6572), .B0(n8273), .Y(n8274));
  NOR2X1  g7132(.A(n8274), .B(n8272), .Y(n8275));
  AOI21X1 g7133(.A0(n8134), .A1(n6470), .B0(n5728), .Y(n8276));
  OAI21X1 g7134(.A0(n8138), .A1(n6486), .B0(n8276), .Y(n8277));
  AOI22X1 g7135(.A0(n6470), .A1(n8139), .B0(n6429), .B1(n5728), .Y(n8278));
  OAI21X1 g7136(.A0(n7132), .A1(n6486), .B0(n8278), .Y(n8279));
  INVX1   g7137(.A(n8279), .Y(n8280));
  OAI21X1 g7138(.A0(n7132), .A1(n6436), .B0(n5729), .Y(n8281));
  AOI21X1 g7139(.A0(n8139), .A1(n6441), .B0(n8281), .Y(n8282));
  AOI22X1 g7140(.A0(n6429), .A1(n8139), .B0(n6379), .B1(n5728), .Y(n8283));
  OAI21X1 g7141(.A0(n7132), .A1(n6477), .B0(n8283), .Y(n8284));
  AOI21X1 g7142(.A0(n8134), .A1(n6379), .B0(n5728), .Y(n8285));
  OAI21X1 g7143(.A0(n8138), .A1(n6393), .B0(n8285), .Y(n8286));
  INVX1   g7144(.A(n8286), .Y(n8287));
  AOI22X1 g7145(.A0(n6379), .A1(n8139), .B0(n6334), .B1(n5728), .Y(n8288));
  OAI21X1 g7146(.A0(n7132), .A1(n6393), .B0(n8288), .Y(n8289));
  OAI22X1 g7147(.A0(n8287), .A1(n8289), .B0(n8284), .B1(n8282), .Y(n8290));
  OAI22X1 g7148(.A0(n6296), .A1(n8138), .B0(n6249), .B1(n5729), .Y(n8291));
  AOI21X1 g7149(.A0(n8134), .A1(n6301), .B0(n8291), .Y(n8292));
  AOI21X1 g7150(.A0(n8134), .A1(n6284), .B0(n5728), .Y(n8293));
  OAI21X1 g7151(.A0(n8138), .A1(n6360), .B0(n8293), .Y(n8294));
  AOI22X1 g7152(.A0(n6242), .A1(n8139), .B0(n6200), .B1(n5728), .Y(n8295));
  OAI21X1 g7153(.A0(n7132), .A1(n6291), .B0(n8295), .Y(n8296));
  AOI21X1 g7154(.A0(n8134), .A1(n6242), .B0(n5728), .Y(n8297));
  INVX1   g7155(.A(n8297), .Y(n8298));
  AOI21X1 g7156(.A0(n8139), .A1(n6254), .B0(n8298), .Y(n8299));
  NAND2X1 g7157(.A(n8299), .B(n8296), .Y(n8300));
  OAI21X1 g7158(.A0(n8294), .A1(n8292), .B0(n8300), .Y(n8301));
  AOI22X1 g7159(.A0(n6150), .A1(n8139), .B0(n6098), .B1(n5728), .Y(n8302));
  OAI21X1 g7160(.A0(n7132), .A1(n6185), .B0(n8302), .Y(n8303));
  OAI21X1 g7161(.A0(n7132), .A1(n6156), .B0(n5729), .Y(n8304));
  AOI21X1 g7162(.A0(n8139), .A1(n6161), .B0(n8304), .Y(n8305));
  AOI22X1 g7163(.A0(n6098), .A1(n8139), .B0(n6056), .B1(n5728), .Y(n8306));
  OAI21X1 g7164(.A0(n7132), .A1(n6120), .B0(n8306), .Y(n8307));
  OAI21X1 g7165(.A0(n7132), .A1(n6115), .B0(n5729), .Y(n8308));
  AOI21X1 g7166(.A0(n8139), .A1(n6123), .B0(n8308), .Y(n8309));
  OAI22X1 g7167(.A0(n8307), .A1(n8309), .B0(n8305), .B1(n8303), .Y(n8310));
  OAI22X1 g7168(.A0(n6068), .A1(n7132), .B0(n6079), .B1(n5729), .Y(n8311));
  AOI21X1 g7169(.A0(n8139), .A1(n6056), .B0(n8311), .Y(n8312));
  AOI21X1 g7170(.A0(n8139), .A1(n6067), .B0(n5728), .Y(n8313));
  OAI21X1 g7171(.A0(n7132), .A1(n6104), .B0(n8313), .Y(n8314));
  NOR3X1  g7172(.A(n8314), .B(n8312), .C(n8310), .Y(n8315));
  NOR2X1  g7173(.A(n8305), .B(n8303), .Y(n8316));
  NAND2X1 g7174(.A(n8309), .B(n8307), .Y(n8317));
  AOI22X1 g7175(.A0(n6200), .A1(n8139), .B0(n6150), .B1(n5728), .Y(n8318));
  OAI21X1 g7176(.A0(n7132), .A1(n6222), .B0(n8318), .Y(n8319));
  OAI21X1 g7177(.A0(n7132), .A1(n6206), .B0(n5729), .Y(n8320));
  AOI21X1 g7178(.A0(n8139), .A1(n6211), .B0(n8320), .Y(n8321));
  AOI22X1 g7179(.A0(n8319), .A1(n8321), .B0(n8305), .B1(n8303), .Y(n8322));
  OAI21X1 g7180(.A0(n8317), .A1(n8316), .B0(n8322), .Y(n8323));
  OAI22X1 g7181(.A0(n6024), .A1(n7132), .B0(n5965), .B1(n5729), .Y(n8324));
  AOI21X1 g7182(.A0(n8139), .A1(n6012), .B0(n8324), .Y(n8325));
  AOI21X1 g7183(.A0(n8139), .A1(n6023), .B0(n5728), .Y(n8326));
  OAI21X1 g7184(.A0(n7132), .A1(n6079), .B0(n8326), .Y(n8327));
  NOR2X1  g7185(.A(n8327), .B(n8325), .Y(n8328));
  AOI22X1 g7186(.A0(n5984), .A1(n8134), .B0(n5933), .B1(n5728), .Y(n8329));
  OAI21X1 g7187(.A0(n8138), .A1(n5965), .B0(n8329), .Y(n8330));
  INVX1   g7188(.A(n8330), .Y(n8331));
  AOI21X1 g7189(.A0(n8139), .A1(n5984), .B0(n5728), .Y(n8332));
  OAI21X1 g7190(.A0(n7132), .A1(n5965), .B0(n8332), .Y(n8333));
  NAND2X1 g7191(.A(n8333), .B(n8331), .Y(n8334));
  AOI22X1 g7192(.A0(n8325), .A1(n8327), .B0(n8314), .B1(n8312), .Y(n8335));
  OAI21X1 g7193(.A0(n8334), .A1(n8328), .B0(n8335), .Y(n8336));
  NOR2X1  g7194(.A(n8336), .B(n8310), .Y(n8337));
  NOR4X1  g7195(.A(n8323), .B(n8315), .C(n8301), .D(n8337), .Y(n8338));
  NOR3X1  g7196(.A(n8321), .B(n8319), .C(n8301), .Y(n8339));
  NOR2X1  g7197(.A(n8299), .B(n8296), .Y(n8340));
  OAI21X1 g7198(.A0(n8294), .A1(n8292), .B0(n8340), .Y(n8341));
  AOI21X1 g7199(.A0(n8134), .A1(n6334), .B0(n5728), .Y(n8342));
  OAI21X1 g7200(.A0(n8138), .A1(n6346), .B0(n8342), .Y(n8343));
  AOI22X1 g7201(.A0(n6334), .A1(n8139), .B0(n6284), .B1(n5728), .Y(n8344));
  OAI21X1 g7202(.A0(n7132), .A1(n6346), .B0(n8344), .Y(n8345));
  INVX1   g7203(.A(n8345), .Y(n8346));
  AOI22X1 g7204(.A0(n8343), .A1(n8346), .B0(n8294), .B1(n8292), .Y(n8347));
  NAND2X1 g7205(.A(n8347), .B(n8341), .Y(n8348));
  NOR4X1  g7206(.A(n8339), .B(n8338), .C(n8290), .D(n8348), .Y(n8349));
  OAI22X1 g7207(.A0(n8331), .A1(n8333), .B0(n8327), .B1(n8325), .Y(n8350));
  NOR4X1  g7208(.A(n8323), .B(n8315), .C(n8301), .D(n8350), .Y(n8351));
  AOI21X1 g7209(.A0(n8139), .A1(n5945), .B0(n5728), .Y(n8352));
  OAI21X1 g7210(.A0(n7132), .A1(n5925), .B0(n8352), .Y(n8353));
  INVX1   g7211(.A(n8353), .Y(n8354));
  AOI22X1 g7212(.A0(n5945), .A1(n8134), .B0(n5894), .B1(n5728), .Y(n8355));
  OAI21X1 g7213(.A0(n8138), .A1(n5925), .B0(n8355), .Y(n8356));
  AOI22X1 g7214(.A0(n8134), .A1(n5878), .B0(n5894), .B1(n8139), .Y(n8357));
  NAND2X1 g7215(.A(n8134), .B(n5894), .Y(n8358));
  AOI21X1 g7216(.A0(n8139), .A1(n5878), .B0(n5728), .Y(n8359));
  AOI22X1 g7217(.A0(n8358), .A1(n8359), .B0(n8137), .B1(n5846), .Y(n8360));
  NAND4X1 g7218(.A(n8358), .B(n8137), .C(n5846), .D(n8359), .Y(n8361));
  OAI21X1 g7219(.A0(n8360), .A1(n8357), .B0(n8361), .Y(n8362));
  AOI21X1 g7220(.A0(n8356), .A1(n8354), .B0(n8362), .Y(n8363));
  NOR2X1  g7221(.A(n8356), .B(n8354), .Y(n8364));
  OAI21X1 g7222(.A0(n8364), .A1(n8363), .B0(n8351), .Y(n8365));
  NAND2X1 g7223(.A(n8365), .B(n8349), .Y(n8366));
  NOR3X1  g7224(.A(n8346), .B(n8343), .C(n8290), .Y(n8367));
  NOR2X1  g7225(.A(n8284), .B(n8282), .Y(n8368));
  NAND2X1 g7226(.A(n8289), .B(n8287), .Y(n8369));
  NOR2X1  g7227(.A(n8369), .B(n8368), .Y(n8370));
  NAND2X1 g7228(.A(n8284), .B(n8282), .Y(n8371));
  OAI21X1 g7229(.A0(n8280), .A1(n8277), .B0(n8371), .Y(n8372));
  NOR3X1  g7230(.A(n8372), .B(n8370), .C(n8367), .Y(n8373));
  AOI22X1 g7231(.A0(n8366), .A1(n8373), .B0(n8280), .B1(n8277), .Y(n8374));
  AOI21X1 g7232(.A0(n8274), .A1(n8272), .B0(n8374), .Y(n8375));
  AOI22X1 g7233(.A0(n6559), .A1(n8139), .B0(n6516), .B1(n5728), .Y(n8376));
  OAI21X1 g7234(.A0(n7132), .A1(n6607), .B0(n8376), .Y(n8377));
  AOI21X1 g7235(.A0(n8134), .A1(n6559), .B0(n5728), .Y(n8378));
  OAI21X1 g7236(.A0(n8138), .A1(n6607), .B0(n8378), .Y(n8379));
  INVX1   g7237(.A(n8379), .Y(n8380));
  NAND2X1 g7238(.A(n8380), .B(n8377), .Y(n8381));
  OAI21X1 g7239(.A0(n8375), .A1(n8275), .B0(n8381), .Y(n8382));
  OAI22X1 g7240(.A0(n8377), .A1(n8380), .B0(n8263), .B1(n8261), .Y(n8383));
  NOR2X1  g7241(.A(n8383), .B(n8258), .Y(n8384));
  AOI21X1 g7242(.A0(n8384), .A1(n8382), .B0(n8270), .Y(n8385));
  NOR4X1  g7243(.A(n8248), .B(n8219), .C(n8213), .D(n8385), .Y(n8386));
  NAND2X1 g7244(.A(n8212), .B(n8210), .Y(n8387));
  NOR3X1  g7245(.A(n8224), .B(n8222), .C(n8219), .Y(n8388));
  AOI21X1 g7246(.A0(n8218), .A1(n8215), .B0(n8388), .Y(n8389));
  OAI21X1 g7247(.A0(n8389), .A1(n8213), .B0(n8387), .Y(n8390));
  NOR3X1  g7248(.A(n8390), .B(n8386), .C(n8207), .Y(n8391));
  NAND2X1 g7249(.A(n8391), .B(n8167), .Y(n8392));
  NOR3X1  g7250(.A(n8392), .B(n8182), .C(n8176), .Y(n8393));
  NOR4X1  g7251(.A(n8205), .B(n8200), .C(n8196), .D(n8393), .Y(n8394));
  XOR2X1  g7252(.A(n7132), .B(n5853), .Y(n8395));
  INVX1   g7253(.A(n8395), .Y(n8396));
  NAND4X1 g7254(.A(n8394), .B(n8191), .C(n8174), .D(n8396), .Y(n8397));
  NAND4X1 g7255(.A(n8185), .B(n8150), .C(n8142), .D(n8186), .Y(n8398));
  NAND2X1 g7256(.A(n8155), .B(n8152), .Y(n8399));
  NAND4X1 g7257(.A(n8399), .B(n8150), .C(n8142), .D(n8188), .Y(n8400));
  NAND3X1 g7258(.A(n8400), .B(n8398), .C(n8174), .Y(n8401));
  NOR2X1  g7259(.A(n8175), .B(n8140), .Y(n8402));
  AOI21X1 g7260(.A0(n8192), .A1(n8140), .B0(n8402), .Y(n8403));
  OAI21X1 g7261(.A0(n8192), .A1(n8141), .B0(n8403), .Y(n8404));
  NOR2X1  g7262(.A(n8149), .B(n8143), .Y(n8405));
  NAND2X1 g7263(.A(n8180), .B(n8179), .Y(n8406));
  AOI21X1 g7264(.A0(n8149), .A1(n8143), .B0(n8406), .Y(n8407));
  OAI21X1 g7265(.A0(n8407), .A1(n8405), .B0(n8142), .Y(n8408));
  NOR2X1  g7266(.A(n8204), .B(n8203), .Y(n8409));
  NAND3X1 g7267(.A(n8409), .B(n8150), .C(n8142), .Y(n8410));
  NAND4X1 g7268(.A(n8167), .B(n8150), .C(n8142), .D(n8391), .Y(n8411));
  NAND4X1 g7269(.A(n8410), .B(n8408), .C(n8404), .D(n8411), .Y(n8412));
  OAI21X1 g7270(.A0(n8412), .A1(n8401), .B0(n8395), .Y(n8413));
  NAND3X1 g7271(.A(n8413), .B(n8397), .C(n5857), .Y(n8414));
  NOR3X1  g7272(.A(n5915), .B(n5867), .C(n5862), .Y(n8415));
  INVX1   g7273(.A(n8415), .Y(n8416));
  NOR4X1  g7274(.A(n8412), .B(n8401), .C(n5815), .D(n8416), .Y(n8417));
  NAND2X1 g7275(.A(n7146), .B(n7131), .Y(n8421));
  INVX1   g7276(.A(n8421), .Y(n8422));
  OAI22X1 g7277(.A0(n7147), .A1(n7153), .B0(n7448), .B1(n8422), .Y(n8423));
  NAND3X1 g7278(.A(n7106), .B(n6823), .C(n7113), .Y(n8424));
  AOI22X1 g7279(.A0(n7111), .A1(n7093), .B0(n7058), .B1(n7074), .Y(n8425));
  AOI21X1 g7280(.A0(n6823), .A1(n6995), .B0(n6994), .Y(n8426));
  NAND3X1 g7281(.A(n8426), .B(n8425), .C(n8424), .Y(n8427));
  NOR2X1  g7282(.A(n8427), .B(n8423), .Y(n8428));
  NAND4X1 g7283(.A(n7448), .B(n7146), .C(n7131), .D(n7153), .Y(n8429));
  OAI21X1 g7284(.A0(n7146), .A1(n7453), .B0(n8429), .Y(n8430));
  NOR2X1  g7285(.A(n8430), .B(n8428), .Y(n8431));
  OAI21X1 g7286(.A0(n5870), .A1(n5706), .B0(n7100), .Y(n8432));
  NAND3X1 g7287(.A(n6994), .B(n6823), .C(n6995), .Y(n8433));
  OAI21X1 g7288(.A0(n5870), .A1(n5669), .B0(n6953), .Y(n8434));
  AOI21X1 g7289(.A0(n6823), .A1(n5658), .B0(n6929), .Y(n8435));
  NAND2X1 g7290(.A(n6886), .B(n6878), .Y(n8436));
  NOR2X1  g7291(.A(n6852), .B(n6885), .Y(n8439));
  NAND2X1 g7292(.A(n6790), .B(n8439), .Y(n8441));
  NOR2X1  g7293(.A(n6849), .B(n6848), .Y(n8444));
  AOI21X1 g7294(.A0(n6851), .A1(n6935), .B0(n8444), .Y(n8445));
  NAND3X1 g7295(.A(n8445), .B(n8441), .C(n8436), .Y(n8446));
  AOI22X1 g7296(.A0(n6729), .A1(n6820), .B0(n6699), .B1(n6684), .Y(n8447));
  NOR2X1  g7297(.A(n6657), .B(n6645), .Y(n8448));
  NAND2X1 g7298(.A(n8448), .B(n8447), .Y(n8449));
  NAND2X1 g7299(.A(n6820), .B(n6729), .Y(n8450));
  NOR2X1  g7300(.A(n6699), .B(n6684), .Y(n8451));
  OAI22X1 g7301(.A0(n6767), .A1(n6824), .B0(n6820), .B1(n6729), .Y(n8452));
  AOI21X1 g7302(.A0(n8451), .A1(n8450), .B0(n8452), .Y(n8453));
  NAND3X1 g7303(.A(n8453), .B(n8449), .C(n8439), .Y(n8454));
  NOR2X1  g7304(.A(n6569), .B(n6558), .Y(n8455));
  NAND2X1 g7305(.A(n6572), .B(n6516), .Y(n8456));
  AOI22X1 g7306(.A0(n6333), .A1(n6353), .B0(n6211), .B1(n6206), .Y(n8457));
  AOI22X1 g7307(.A0(n6296), .A1(n6301), .B0(n6254), .B1(n6249), .Y(n8458));
  NAND2X1 g7308(.A(n8458), .B(n8457), .Y(n8459));
  OAI22X1 g7309(.A0(n6150), .A1(n6185), .B0(n6120), .B1(n6098), .Y(n8460));
  NOR3X1  g7310(.A(n6134), .B(n8460), .C(n8459), .Y(n8462));
  AOI21X1 g7311(.A0(n6011), .A1(n6009), .B0(n6023), .Y(n8463));
  NAND2X1 g7312(.A(n8463), .B(n8462), .Y(n8464));
  AOI22X1 g7313(.A0(n6098), .A1(n6120), .B0(n6068), .B1(n6056), .Y(n8465));
  AOI22X1 g7314(.A0(n6200), .A1(n6222), .B0(n6185), .B1(n6150), .Y(n8466));
  OAI21X1 g7315(.A0(n8465), .A1(n8460), .B0(n8466), .Y(n8467));
  NAND3X1 g7316(.A(n8467), .B(n8458), .C(n8457), .Y(n8468));
  OAI22X1 g7317(.A0(n6480), .A1(n6485), .B0(n6441), .B1(n6436), .Y(n8469));
  INVX1   g7318(.A(n8469), .Y(n8470));
  OAI22X1 g7319(.A0(n6296), .A1(n6301), .B0(n6254), .B1(n6249), .Y(n8471));
  AOI22X1 g7320(.A0(n6333), .A1(n6353), .B0(n6301), .B1(n6296), .Y(n8472));
  AOI21X1 g7321(.A0(n8472), .A1(n8471), .B0(n6399), .Y(n8474));
  NAND4X1 g7322(.A(n8470), .B(n8468), .C(n8464), .D(n8474), .Y(n8475));
  NAND3X1 g7323(.A(n6023), .B(n6011), .C(n6009), .Y(n8476));
  NAND2X1 g7324(.A(n8476), .B(n8462), .Y(n8477));
  NOR2X1  g7325(.A(n5945), .B(n5925), .Y(n8478));
  AOI22X1 g7326(.A0(n5965), .A1(n5984), .B0(n5945), .B1(n5925), .Y(n8480));
  OAI21X1 g7327(.A0(n5995), .A1(n8478), .B0(n8480), .Y(n8481));
  OAI21X1 g7328(.A0(n5964), .A1(n5960), .B0(n5981), .Y(n8482));
  AOI21X1 g7329(.A0(n8482), .A1(n8481), .B0(n8477), .Y(n8483));
  AOI22X1 g7330(.A0(n6527), .A1(n6532), .B0(n6485), .B1(n6480), .Y(n8487));
  OAI21X1 g7331(.A0(n6499), .A1(n6522), .B0(n8487), .Y(n8488));
  AOI21X1 g7332(.A0(n6397), .A1(n8470), .B0(n8488), .Y(n8489));
  OAI21X1 g7333(.A0(n8483), .A1(n8475), .B0(n8489), .Y(n8490));
  AOI21X1 g7334(.A0(n8490), .A1(n8456), .B0(n6618), .Y(n8492));
  OAI21X1 g7335(.A0(n8492), .A1(n8455), .B0(n6621), .Y(n8494));
  INVX1   g7336(.A(n8447), .Y(n8495));
  OAI22X1 g7337(.A0(n6691), .A1(n6658), .B0(n6604), .B1(n6599), .Y(n8496));
  NOR2X1  g7338(.A(n8496), .B(n8495), .Y(n8497));
  AOI21X1 g7339(.A0(n8497), .A1(n8494), .B0(n8454), .Y(n8498));
  NOR3X1  g7340(.A(n8498), .B(n8446), .C(n8435), .Y(n8499));
  OAI22X1 g7341(.A0(n6916), .A1(n6925), .B0(n6886), .B1(n6878), .Y(n8502));
  NAND3X1 g7342(.A(n8502), .B(n6973), .C(n8434), .Y(n8503));
  NAND2X1 g7343(.A(n8503), .B(n7008), .Y(n8504));
  AOI21X1 g7344(.A0(n8499), .A1(n8434), .B0(n8504), .Y(n8505));
  NAND4X1 g7345(.A(n8433), .B(n8425), .C(n8424), .D(n8505), .Y(n8506));
  AOI21X1 g7346(.A0(n8506), .A1(n8432), .B0(n8423), .Y(n8507));
  NOR2X1  g7347(.A(n7058), .B(n7074), .Y(n8508));
  NAND3X1 g7348(.A(n8508), .B(n8425), .C(n8424), .Y(n8509));
  AOI21X1 g7349(.A0(n6823), .A1(n7070), .B0(n7111), .Y(n8510));
  NAND2X1 g7350(.A(n8510), .B(n8424), .Y(n8511));
  AOI21X1 g7351(.A0(n8511), .A1(n8509), .B0(n8423), .Y(n8512));
  NOR2X1  g7352(.A(n8512), .B(n8507), .Y(n8513));
  AOI21X1 g7353(.A0(n8513), .A1(n8431), .B0(n6018), .Y(n8514));
  NAND3X1 g7354(.A(n8513), .B(n8431), .C(n5905), .Y(n8515));
  NOR2X1  g7355(.A(n8415), .B(n5729), .Y(n8516));
  OAI21X1 g7356(.A0(n5846), .A1(n5728), .B0(n7456), .Y(n8517));
  OAI21X1 g7357(.A0(n8517), .A1(n8516), .B0(P2_B_REG_SCAN_IN), .Y(n8518));
  XOR2X1  g7358(.A(n7448), .B(n8128), .Y(n8519));
  XOR2X1  g7359(.A(n7153), .B(n7146), .Y(n8520));
  XOR2X1  g7360(.A(n6960), .B(n6953), .Y(n8524));
  XOR2X1  g7361(.A(n6815), .B(n6806), .Y(n8528));
  XOR2X1  g7362(.A(n6774), .B(n6767), .Y(n8529));
  XOR2X1  g7363(.A(n6657), .B(n6691), .Y(n8530));
  XOR2X1  g7364(.A(n5894), .B(n5878), .Y(n8531));
  OAI22X1 g7365(.A0(n6062), .A1(n6070), .B0(n5985), .B1(n5982), .Y(n8532));
  NOR2X1  g7366(.A(n8532), .B(n6172), .Y(n8533));
  NAND3X1 g7367(.A(n6128), .B(n6212), .C(n8533), .Y(n8536));
  NOR4X1  g7368(.A(n8531), .B(n6075), .C(n5946), .D(n8536), .Y(n8537));
  NOR2X1  g7369(.A(n6413), .B(n6268), .Y(n8538));
  NAND4X1 g7370(.A(n8538), .B(n8537), .C(n6302), .D(n6354), .Y(n8540));
  XOR2X1  g7371(.A(n6569), .B(n6559), .Y(n8541));
  NOR2X1  g7372(.A(n8541), .B(n6446), .Y(n8542));
  NAND3X1 g7373(.A(n6491), .B(n6533), .C(n8542), .Y(n8545));
  NOR4X1  g7374(.A(n8540), .B(n8530), .C(n6611), .D(n8545), .Y(n8546));
  NAND2X1 g7375(.A(n8546), .B(n6700), .Y(n8547));
  NOR4X1  g7376(.A(n8529), .B(n8528), .C(n6744), .D(n8547), .Y(n8548));
  NAND3X1 g7377(.A(n8548), .B(n6850), .C(n6887), .Y(n8549));
  NOR4X1  g7378(.A(n7002), .B(n8524), .C(n6930), .D(n8549), .Y(n8550));
  NAND3X1 g7379(.A(n8550), .B(n7035), .C(n7072), .Y(n8551));
  NOR4X1  g7380(.A(n7115), .B(n8520), .C(n8519), .D(n8551), .Y(n8552));
  XOR2X1  g7381(.A(n8552), .B(n5860), .Y(n8553));
  NOR2X1  g7382(.A(n5857), .B(n5847), .Y(n8554));
  NAND2X1 g7383(.A(n8554), .B(n8553), .Y(n8555));
  NAND3X1 g7384(.A(n8555), .B(n8518), .C(n8515), .Y(n8556));
  NOR3X1  g7385(.A(n8556), .B(n8514), .C(n8417), .Y(n8557));
  NAND2X1 g7386(.A(n8518), .B(n5728), .Y(n8558));
  NAND2X1 g7387(.A(n8518), .B(P2_U3151), .Y(n8559));
  OAI21X1 g7388(.A0(n8558), .A1(n8417), .B0(n8559), .Y(n8560));
  AOI21X1 g7389(.A0(n8557), .A1(n8414), .B0(n8560), .Y(P2_U3296));
  OAI21X1 g7390(.A0(n5853), .A1(n5847), .B0(n5857), .Y(n8562));
  INVX1   g7391(.A(n8562), .Y(n8563));
  AOI21X1 g7392(.A0(n8554), .A1(n5842), .B0(n8563), .Y(n8564));
  XOR2X1  g7393(.A(n8564), .B(n6353), .Y(n8565));
  INVX1   g7394(.A(n8565), .Y(n8566));
  NAND2X1 g7395(.A(n8566), .B(n6334), .Y(n8567));
  XOR2X1  g7396(.A(n8564), .B(n6485), .Y(n8568));
  INVX1   g7397(.A(n8568), .Y(n8569));
  NOR2X1  g7398(.A(n8569), .B(n6470), .Y(n8570));
  XOR2X1  g7399(.A(n8564), .B(n6441), .Y(n8571));
  AOI22X1 g7400(.A0(n8571), .A1(n6436), .B0(n6480), .B1(n8568), .Y(n8572));
  INVX1   g7401(.A(n8554), .Y(n8573));
  OAI21X1 g7402(.A0(n8573), .A1(n7235), .B0(n8562), .Y(n8574));
  XOR2X1  g7403(.A(n8574), .B(n6393), .Y(n8575));
  NAND2X1 g7404(.A(n8575), .B(n6412), .Y(n8576));
  NAND2X1 g7405(.A(n8576), .B(n8572), .Y(n8577));
  NOR2X1  g7406(.A(n8575), .B(n6412), .Y(n8578));
  OAI22X1 g7407(.A0(n8571), .A1(n6436), .B0(n6480), .B1(n8568), .Y(n8579));
  AOI21X1 g7408(.A0(n8578), .A1(n8572), .B0(n8579), .Y(n8580));
  OAI22X1 g7409(.A0(n8577), .A1(n8567), .B0(n8570), .B1(n8580), .Y(n8581));
  XOR2X1  g7410(.A(n8564), .B(n6532), .Y(n8582));
  NAND2X1 g7411(.A(n8582), .B(n6527), .Y(n8583));
  NOR2X1  g7412(.A(n8582), .B(n6527), .Y(n8584));
  AOI21X1 g7413(.A0(n8583), .A1(n8581), .B0(n8584), .Y(n8585));
  NAND2X1 g7414(.A(n8565), .B(n6333), .Y(n8586));
  NAND4X1 g7415(.A(n8583), .B(n8576), .C(n8572), .D(n8586), .Y(n8587));
  XOR2X1  g7416(.A(n8564), .B(n5984), .Y(n8588));
  XOR2X1  g7417(.A(n8574), .B(n6024), .Y(n8589));
  AOI22X1 g7418(.A0(n8588), .A1(n5965), .B0(n6079), .B1(n8589), .Y(n8590));
  XOR2X1  g7419(.A(n8564), .B(n5945), .Y(n8591));
  OAI21X1 g7420(.A0(n8574), .A1(n5878), .B0(n5894), .Y(n8592));
  AOI21X1 g7421(.A0(n8591), .A1(n5925), .B0(n8592), .Y(n8593));
  NAND2X1 g7422(.A(n8574), .B(n5879), .Y(n8594));
  AOI21X1 g7423(.A0(n8591), .A1(n5925), .B0(n8594), .Y(n8595));
  NOR2X1  g7424(.A(n8591), .B(n5925), .Y(n8596));
  NOR3X1  g7425(.A(n8596), .B(n8595), .C(n8593), .Y(n8597));
  INVX1   g7426(.A(n8597), .Y(n8598));
  NOR2X1  g7427(.A(n8588), .B(n5965), .Y(n8599));
  NAND2X1 g7428(.A(n8599), .B(n6012), .Y(n8600));
  INVX1   g7429(.A(n8589), .Y(n8601));
  OAI21X1 g7430(.A0(n8599), .A1(n6012), .B0(n8601), .Y(n8602));
  NAND2X1 g7431(.A(n8602), .B(n8600), .Y(n8603));
  AOI21X1 g7432(.A0(n8598), .A1(n8590), .B0(n8603), .Y(n8604));
  XOR2X1  g7433(.A(n8564), .B(n6067), .Y(n8605));
  NOR2X1  g7434(.A(n8605), .B(n6104), .Y(n8606));
  NOR2X1  g7435(.A(n8605), .B(n8604), .Y(n8607));
  NOR2X1  g7436(.A(n8607), .B(n8606), .Y(n8608));
  OAI21X1 g7437(.A0(n8604), .A1(n6104), .B0(n8608), .Y(n8609));
  XOR2X1  g7438(.A(n8564), .B(n6254), .Y(n8610));
  NAND2X1 g7439(.A(n8610), .B(n6249), .Y(n8611));
  XOR2X1  g7440(.A(n8564), .B(n6161), .Y(n8612));
  XOR2X1  g7441(.A(n8564), .B(n6211), .Y(n8613));
  AOI22X1 g7442(.A0(n8612), .A1(n6156), .B0(n6206), .B1(n8613), .Y(n8614));
  INVX1   g7443(.A(n8614), .Y(n8615));
  XOR2X1  g7444(.A(n8564), .B(n6123), .Y(n8616));
  INVX1   g7445(.A(n8616), .Y(n8617));
  NOR2X1  g7446(.A(n8617), .B(n6098), .Y(n8618));
  NOR2X1  g7447(.A(n8618), .B(n8615), .Y(n8619));
  NAND2X1 g7448(.A(n8619), .B(n8611), .Y(n8620));
  INVX1   g7449(.A(n8620), .Y(n8621));
  NOR2X1  g7450(.A(n8612), .B(n6156), .Y(n8622));
  NOR2X1  g7451(.A(n8622), .B(n6200), .Y(n8623));
  NOR2X1  g7452(.A(n8616), .B(n6115), .Y(n8624));
  AOI22X1 g7453(.A0(n8622), .A1(n6200), .B0(n8614), .B1(n8624), .Y(n8625));
  OAI21X1 g7454(.A0(n8623), .A1(n8613), .B0(n8625), .Y(n8626));
  NOR2X1  g7455(.A(n8610), .B(n6249), .Y(n8627));
  AOI21X1 g7456(.A0(n8626), .A1(n8611), .B0(n8627), .Y(n8628));
  INVX1   g7457(.A(n8628), .Y(n8629));
  AOI21X1 g7458(.A0(n8621), .A1(n8609), .B0(n8629), .Y(n8630));
  NOR2X1  g7459(.A(n8630), .B(n6296), .Y(n8631));
  XOR2X1  g7460(.A(n8564), .B(n6301), .Y(n8632));
  AOI21X1 g7461(.A0(n8630), .A1(n6296), .B0(n8632), .Y(n8633));
  NOR2X1  g7462(.A(n8633), .B(n8631), .Y(n8634));
  OAI21X1 g7463(.A0(n8634), .A1(n8587), .B0(n8585), .Y(n8635));
  XOR2X1  g7464(.A(n8564), .B(n6569), .Y(n8636));
  XOR2X1  g7465(.A(n8636), .B(n6559), .Y(n8637));
  XOR2X1  g7466(.A(n8637), .B(n8635), .Y(n8638));
  NOR3X1  g7467(.A(n5842), .B(n5839), .C(n5836), .Y(n8639));
  INVX1   g7468(.A(n8639), .Y(n8640));
  NOR3X1  g7469(.A(n5859), .B(n5857), .C(n8640), .Y(n8641));
  NAND2X1 g7470(.A(n5847), .B(n5846), .Y(n8642));
  INVX1   g7471(.A(n8642), .Y(n8643));
  NOR4X1  g7472(.A(n5849), .B(n5847), .C(n5846), .D(n5853), .Y(n8644));
  NOR4X1  g7473(.A(n8643), .B(n7162), .C(n5909), .D(n8644), .Y(n8645));
  NOR4X1  g7474(.A(n7235), .B(n5838), .C(n5836), .D(n8645), .Y(n8646));
  OAI21X1 g7475(.A0(n8646), .A1(n8641), .B0(n5744), .Y(n8647));
  NOR3X1  g7476(.A(n7235), .B(n5838), .C(n5836), .Y(n8648));
  INVX1   g7477(.A(n8648), .Y(n8649));
  NOR4X1  g7478(.A(n5739), .B(n5729), .C(P2_U3151), .D(n7251), .Y(n8650));
  NOR2X1  g7479(.A(n8645), .B(n8648), .Y(n8651));
  NOR3X1  g7480(.A(n5859), .B(n5857), .C(n8639), .Y(n8652));
  NOR2X1  g7481(.A(n5739), .B(n5729), .Y(n8653));
  AOI22X1 g7482(.A0(n8135), .A1(n5847), .B0(n5849), .B1(n7132), .Y(n8654));
  NAND2X1 g7483(.A(n8654), .B(n8653), .Y(n8655));
  NOR3X1  g7484(.A(n8655), .B(n8652), .C(n8651), .Y(n8656));
  INVX1   g7485(.A(n8656), .Y(n8657));
  AOI22X1 g7486(.A0(n8650), .A1(n8649), .B0(P2_STATE_REG_SCAN_IN), .B1(n8657), .Y(n8658));
  INVX1   g7487(.A(n8658), .Y(n8659));
  NOR4X1  g7488(.A(n5739), .B(n5729), .C(P2_U3151), .D(n5862), .Y(n8660));
  NOR4X1  g7489(.A(n5842), .B(n5839), .C(n5836), .D(n5916), .Y(n8661));
  INVX1   g7490(.A(n8661), .Y(n8662));
  NOR2X1  g7491(.A(n8662), .B(n6599), .Y(n8663));
  NOR4X1  g7492(.A(n5842), .B(n5839), .C(n5836), .D(n5951), .Y(n8664));
  INVX1   g7493(.A(n8664), .Y(n8665));
  OAI22X1 g7494(.A0(n6556), .A1(n8639), .B0(n6527), .B1(n8665), .Y(n8666));
  OAI21X1 g7495(.A0(n8666), .A1(n8663), .B0(n8660), .Y(n8667));
  AOI22X1 g7496(.A0(n7233), .A1(n5744), .B0(n8648), .B1(n8650), .Y(n8668));
  INVX1   g7497(.A(n8668), .Y(n8669));
  AOI22X1 g7498(.A0(n6569), .A1(n8669), .B0(P2_REG3_REG_15__SCAN_IN), .B1(P2_U3151), .Y(n8670));
  NAND2X1 g7499(.A(n8670), .B(n8667), .Y(n8671));
  AOI21X1 g7500(.A0(n8659), .A1(n7354), .B0(n8671), .Y(n8672));
  OAI21X1 g7501(.A0(n8647), .A1(n8638), .B0(n8672), .Y(P2_U3181));
  XOR2X1  g7502(.A(n8564), .B(n6925), .Y(n8674));
  NOR2X1  g7503(.A(n8674), .B(n6916), .Y(n8675));
  XOR2X1  g7504(.A(n8574), .B(n6886), .Y(n8676));
  NOR2X1  g7505(.A(n8676), .B(n6890), .Y(n8677));
  NAND2X1 g7506(.A(n8676), .B(n6890), .Y(n8678));
  XOR2X1  g7507(.A(n8574), .B(n6849), .Y(n8679));
  NAND2X1 g7508(.A(n8679), .B(n6842), .Y(n8680));
  NOR2X1  g7509(.A(n8679), .B(n6842), .Y(n8681));
  XOR2X1  g7510(.A(n8564), .B(n6815), .Y(n8682));
  XOR2X1  g7511(.A(n8564), .B(n6737), .Y(n8683));
  NOR2X1  g7512(.A(n8683), .B(n6735), .Y(n8684));
  XOR2X1  g7513(.A(n8574), .B(n6774), .Y(n8685));
  NOR2X1  g7514(.A(n8685), .B(n6767), .Y(n8686));
  AOI21X1 g7515(.A0(n8682), .A1(n6814), .B0(n8686), .Y(n8687));
  NAND2X1 g7516(.A(n8687), .B(n8684), .Y(n8688));
  NOR2X1  g7517(.A(n8682), .B(n6814), .Y(n8689));
  AOI21X1 g7518(.A0(n8685), .A1(n6767), .B0(n8689), .Y(n8690));
  AOI22X1 g7519(.A0(n8688), .A1(n8690), .B0(n8682), .B1(n6814), .Y(n8691));
  XOR2X1  g7520(.A(n8574), .B(n6699), .Y(n8692));
  INVX1   g7521(.A(n8692), .Y(n8693));
  NAND2X1 g7522(.A(n8693), .B(n6684), .Y(n8694));
  NOR2X1  g7523(.A(n8693), .B(n6684), .Y(n8695));
  XOR2X1  g7524(.A(n8564), .B(n6604), .Y(n8696));
  XOR2X1  g7525(.A(n8574), .B(n6657), .Y(n8697));
  AOI22X1 g7526(.A0(n8696), .A1(n6599), .B0(n6691), .B1(n8697), .Y(n8698));
  INVX1   g7527(.A(n8636), .Y(n8699));
  NOR2X1  g7528(.A(n8699), .B(n6559), .Y(n8700));
  NOR2X1  g7529(.A(n8700), .B(n8587), .Y(n8701));
  OAI21X1 g7530(.A0(n8633), .A1(n8631), .B0(n8701), .Y(n8702));
  NOR2X1  g7531(.A(n8700), .B(n8585), .Y(n8703));
  AOI21X1 g7532(.A0(n8699), .A1(n6559), .B0(n8703), .Y(n8704));
  NAND2X1 g7533(.A(n8704), .B(n8702), .Y(n8705));
  NOR2X1  g7534(.A(n8696), .B(n6599), .Y(n8706));
  INVX1   g7535(.A(n8706), .Y(n8707));
  AOI21X1 g7536(.A0(n8707), .A1(n6691), .B0(n8697), .Y(n8708));
  AOI21X1 g7537(.A0(n8706), .A1(n6645), .B0(n8708), .Y(n8709));
  INVX1   g7538(.A(n8709), .Y(n8710));
  AOI21X1 g7539(.A0(n8705), .A1(n8698), .B0(n8710), .Y(n8711));
  OAI21X1 g7540(.A0(n8711), .A1(n8695), .B0(n8694), .Y(n8712));
  NAND2X1 g7541(.A(n8683), .B(n6735), .Y(n8713));
  NAND2X1 g7542(.A(n8713), .B(n8687), .Y(n8714));
  INVX1   g7543(.A(n8714), .Y(n8715));
  AOI21X1 g7544(.A0(n8715), .A1(n8712), .B0(n8691), .Y(n8716));
  OAI21X1 g7545(.A0(n8716), .A1(n8681), .B0(n8680), .Y(n8717));
  AOI21X1 g7546(.A0(n8717), .A1(n8678), .B0(n8677), .Y(n8718));
  NOR2X1  g7547(.A(n8718), .B(n8675), .Y(n8719));
  XOR2X1  g7548(.A(n8574), .B(n6996), .Y(n8720));
  XOR2X1  g7549(.A(n8720), .B(n6987), .Y(n8721));
  NAND2X1 g7550(.A(n8674), .B(n6916), .Y(n8722));
  INVX1   g7551(.A(n8722), .Y(n8723));
  XOR2X1  g7552(.A(n8564), .B(n6960), .Y(n8724));
  NOR2X1  g7553(.A(n8724), .B(n6959), .Y(n8725));
  NOR2X1  g7554(.A(n8725), .B(n8723), .Y(n8726));
  NAND2X1 g7555(.A(n8726), .B(n8721), .Y(n8727));
  NOR2X1  g7556(.A(n8727), .B(n8719), .Y(n8728));
  NOR2X1  g7557(.A(n8720), .B(n6994), .Y(n8729));
  INVX1   g7558(.A(n8729), .Y(n8730));
  INVX1   g7559(.A(n8720), .Y(n8731));
  INVX1   g7560(.A(n8724), .Y(n8732));
  OAI22X1 g7561(.A0(n8731), .A1(n6987), .B0(n6953), .B1(n8732), .Y(n8733));
  INVX1   g7562(.A(n8733), .Y(n8734));
  NAND3X1 g7563(.A(n8734), .B(n8730), .C(n8719), .Y(n8735));
  NAND3X1 g7564(.A(n8734), .B(n8730), .C(n8723), .Y(n8736));
  NAND3X1 g7565(.A(n8734), .B(n8730), .C(n8725), .Y(n8737));
  NOR2X1  g7566(.A(n8732), .B(n6953), .Y(n8738));
  AOI21X1 g7567(.A0(n8738), .A1(n8721), .B0(n8647), .Y(n8739));
  NAND4X1 g7568(.A(n8737), .B(n8736), .C(n8735), .D(n8739), .Y(n8740));
  AOI22X1 g7569(.A0(n6985), .A1(n8640), .B0(n6953), .B1(n8664), .Y(n8745));
  OAI21X1 g7570(.A0(n8662), .A1(n7074), .B0(n8745), .Y(n8746));
  AOI22X1 g7571(.A0(n8660), .A1(n8746), .B0(P2_REG3_REG_26__SCAN_IN), .B1(P2_U3151), .Y(n8747));
  OAI21X1 g7572(.A0(n8658), .A1(n6984), .B0(n8747), .Y(n8748));
  AOI21X1 g7573(.A0(n8669), .A1(n7015), .B0(n8748), .Y(n8749));
  OAI21X1 g7574(.A0(n8740), .A1(n8728), .B0(n8749), .Y(P2_U3180));
  XOR2X1  g7575(.A(n8612), .B(n6156), .Y(n8751));
  INVX1   g7576(.A(n8618), .Y(n8752));
  AOI21X1 g7577(.A0(n8752), .A1(n8609), .B0(n8624), .Y(n8753));
  NOR2X1  g7578(.A(n8751), .B(n8753), .Y(n8755));
  AOI21X1 g7579(.A0(n8753), .A1(n8751), .B0(n8755), .Y(n8756));
  NOR2X1  g7580(.A(n8662), .B(n6206), .Y(n8757));
  OAI22X1 g7581(.A0(n6147), .A1(n8639), .B0(n6115), .B1(n8665), .Y(n8758));
  OAI21X1 g7582(.A0(n8758), .A1(n8757), .B0(n8660), .Y(n8759));
  AOI22X1 g7583(.A0(n6161), .A1(n8669), .B0(P2_REG3_REG_6__SCAN_IN), .B1(P2_U3151), .Y(n8760));
  NAND2X1 g7584(.A(n8760), .B(n8759), .Y(n8761));
  AOI21X1 g7585(.A0(n8659), .A1(n6148), .B0(n8761), .Y(n8762));
  OAI21X1 g7586(.A0(n8756), .A1(n8647), .B0(n8762), .Y(P2_U3179));
  XOR2X1  g7587(.A(n8692), .B(n6702), .Y(n8764));
  XOR2X1  g7588(.A(n8764), .B(n8711), .Y(n8765));
  NOR2X1  g7589(.A(n8658), .B(n6681), .Y(n8766));
  INVX1   g7590(.A(n8660), .Y(n8767));
  NAND2X1 g7591(.A(n8661), .B(n6729), .Y(n8768));
  AOI22X1 g7592(.A0(n6682), .A1(n8640), .B0(n6645), .B1(n8664), .Y(n8769));
  AOI21X1 g7593(.A0(n8769), .A1(n8768), .B0(n8767), .Y(n8770));
  OAI22X1 g7594(.A0(n6699), .A1(n8668), .B0(n6680), .B1(P2_STATE_REG_SCAN_IN), .Y(n8771));
  NOR3X1  g7595(.A(n8771), .B(n8770), .C(n8766), .Y(n8772));
  OAI21X1 g7596(.A0(n8765), .A1(n8647), .B0(n8772), .Y(P2_U3178));
  INVX1   g7597(.A(n8647), .Y(n8774));
  XOR2X1  g7598(.A(n8588), .B(n7262), .Y(n8775));
  INVX1   g7599(.A(n8588), .Y(n8776));
  NOR2X1  g7600(.A(n8776), .B(n7262), .Y(n8777));
  OAI21X1 g7601(.A0(n8599), .A1(n8777), .B0(n8598), .Y(n8778));
  OAI21X1 g7602(.A0(n8775), .A1(n8598), .B0(n8778), .Y(n8779));
  NAND2X1 g7603(.A(n8779), .B(n8774), .Y(n8780));
  NAND2X1 g7604(.A(n8659), .B(P2_REG3_REG_2__SCAN_IN), .Y(n8781));
  AOI22X1 g7605(.A0(n5933), .A1(n8664), .B0(n8640), .B1(P2_REG3_REG_2__SCAN_IN), .Y(n8782));
  OAI21X1 g7606(.A0(n8662), .A1(n6079), .B0(n8782), .Y(n8783));
  NAND2X1 g7607(.A(n8783), .B(n8660), .Y(n8784));
  AOI22X1 g7608(.A0(n5984), .A1(n8669), .B0(P2_REG3_REG_2__SCAN_IN), .B1(P2_U3151), .Y(n8785));
  NAND4X1 g7609(.A(n8784), .B(n8781), .C(n8780), .D(n8785), .Y(P2_U3177));
  NOR2X1  g7610(.A(n8566), .B(n6334), .Y(n8787));
  OAI21X1 g7611(.A0(n8634), .A1(n8787), .B0(n8567), .Y(n8788));
  XOR2X1  g7612(.A(n8575), .B(n6379), .Y(n8789));
  NOR2X1  g7613(.A(n8789), .B(n8788), .Y(n8790));
  AOI21X1 g7614(.A0(n8789), .A1(n8788), .B0(n8790), .Y(n8792));
  NOR2X1  g7615(.A(n8662), .B(n6436), .Y(n8793));
  OAI22X1 g7616(.A0(n6376), .A1(n8639), .B0(n6333), .B1(n8665), .Y(n8794));
  OAI21X1 g7617(.A0(n8794), .A1(n8793), .B0(n8660), .Y(n8795));
  AOI22X1 g7618(.A0(n6423), .A1(n8669), .B0(P2_REG3_REG_11__SCAN_IN), .B1(P2_U3151), .Y(n8796));
  NAND2X1 g7619(.A(n8796), .B(n8795), .Y(n8797));
  AOI21X1 g7620(.A0(n8659), .A1(n6377), .B0(n8797), .Y(n8798));
  OAI21X1 g7621(.A0(n8792), .A1(n8647), .B0(n8798), .Y(P2_U3176));
  XOR2X1  g7622(.A(n8679), .B(n6842), .Y(n8800));
  XOR2X1  g7623(.A(n8800), .B(n8716), .Y(n8801));
  AOI22X1 g7624(.A0(n6840), .A1(n8640), .B0(n6806), .B1(n8664), .Y(n8802));
  OAI21X1 g7625(.A0(n8662), .A1(n6890), .B0(n8802), .Y(n8803));
  AOI22X1 g7626(.A0(n8660), .A1(n8803), .B0(P2_REG3_REG_22__SCAN_IN), .B1(P2_U3151), .Y(n8804));
  OAI21X1 g7627(.A0(n8658), .A1(n6839), .B0(n8804), .Y(n8805));
  AOI21X1 g7628(.A0(n8669), .A1(n6849), .B0(n8805), .Y(n8806));
  OAI21X1 g7629(.A0(n8801), .A1(n8647), .B0(n8806), .Y(P2_U3175));
  INVX1   g7630(.A(n8571), .Y(n8808));
  NAND2X1 g7631(.A(n8808), .B(n6429), .Y(n8809));
  AOI21X1 g7632(.A0(n8788), .A1(n8576), .B0(n8578), .Y(n8810));
  OAI21X1 g7633(.A0(n8568), .A1(n6480), .B0(n8572), .Y(n8811));
  AOI21X1 g7634(.A0(n8810), .A1(n8809), .B0(n8811), .Y(n8812));
  AOI21X1 g7635(.A0(n8571), .A1(n6436), .B0(n8810), .Y(n8813));
  AOI22X1 g7636(.A0(n8808), .A1(n6429), .B0(n6480), .B1(n8569), .Y(n8814));
  OAI21X1 g7637(.A0(n8569), .A1(n6480), .B0(n8814), .Y(n8815));
  OAI21X1 g7638(.A0(n8815), .A1(n8813), .B0(n8774), .Y(n8816));
  INVX1   g7639(.A(n6468), .Y(n8817));
  OAI22X1 g7640(.A0(n8817), .A1(n8639), .B0(n6436), .B1(n8665), .Y(n8818));
  AOI21X1 g7641(.A0(n8661), .A1(n6516), .B0(n8818), .Y(n8819));
  AOI22X1 g7642(.A0(n6485), .A1(n8669), .B0(P2_REG3_REG_13__SCAN_IN), .B1(P2_U3151), .Y(n8820));
  OAI21X1 g7643(.A0(n8819), .A1(n8767), .B0(n8820), .Y(n8821));
  AOI21X1 g7644(.A0(n8659), .A1(n6468), .B0(n8821), .Y(n8822));
  OAI21X1 g7645(.A0(n8816), .A1(n8812), .B0(n8822), .Y(P2_U3174));
  XOR2X1  g7646(.A(n8685), .B(n6767), .Y(n8824));
  AOI21X1 g7647(.A0(n8713), .A1(n8712), .B0(n8684), .Y(n8825));
  NOR2X1  g7648(.A(n8824), .B(n8825), .Y(n8827));
  AOI21X1 g7649(.A0(n8825), .A1(n8824), .B0(n8827), .Y(n8828));
  AOI22X1 g7650(.A0(n6765), .A1(n8640), .B0(n6729), .B1(n8664), .Y(n8829));
  OAI21X1 g7651(.A0(n8662), .A1(n6814), .B0(n8829), .Y(n8830));
  AOI22X1 g7652(.A0(n8660), .A1(n8830), .B0(P2_REG3_REG_20__SCAN_IN), .B1(P2_U3151), .Y(n8831));
  OAI21X1 g7653(.A0(n8658), .A1(n6764), .B0(n8831), .Y(n8832));
  AOI21X1 g7654(.A0(n8669), .A1(n6774), .B0(n8832), .Y(n8833));
  OAI21X1 g7655(.A0(n8828), .A1(n8647), .B0(n8833), .Y(P2_U3173));
  AOI21X1 g7656(.A0(n8660), .A1(n8640), .B0(n8659), .Y(n8835));
  NOR2X1  g7657(.A(n8767), .B(n5925), .Y(n8837));
  AOI22X1 g7658(.A0(n8661), .A1(n8837), .B0(P2_REG3_REG_0__SCAN_IN), .B1(P2_U3151), .Y(n8838));
  OAI21X1 g7659(.A0(n8668), .A1(n5879), .B0(n8838), .Y(n8839));
  AOI21X1 g7660(.A0(n8531), .A1(n8774), .B0(n8839), .Y(n8840));
  OAI21X1 g7661(.A0(n8835), .A1(n8063), .B0(n8840), .Y(P2_U3172));
  XOR2X1  g7662(.A(n8632), .B(n6296), .Y(n8842));
  XOR2X1  g7663(.A(n8842), .B(n8630), .Y(n8843));
  NOR2X1  g7664(.A(n8662), .B(n6333), .Y(n8844));
  OAI22X1 g7665(.A0(n7317), .A1(n8639), .B0(n6249), .B1(n8665), .Y(n8845));
  OAI21X1 g7666(.A0(n8845), .A1(n8844), .B0(n8660), .Y(n8846));
  AOI22X1 g7667(.A0(n6301), .A1(n8669), .B0(P2_REG3_REG_9__SCAN_IN), .B1(P2_U3151), .Y(n8847));
  NAND2X1 g7668(.A(n8847), .B(n8846), .Y(n8848));
  AOI21X1 g7669(.A0(n8659), .A1(n6282), .B0(n8848), .Y(n8849));
  OAI21X1 g7670(.A0(n8843), .A1(n8647), .B0(n8849), .Y(P2_U3171));
  XOR2X1  g7671(.A(n8605), .B(n6104), .Y(n8851));
  XOR2X1  g7672(.A(n8851), .B(n8604), .Y(n8852));
  OAI22X1 g7673(.A0(n6053), .A1(n8639), .B0(n6079), .B1(n8665), .Y(n8853));
  AOI21X1 g7674(.A0(n8661), .A1(n6098), .B0(n8853), .Y(n8854));
  AOI22X1 g7675(.A0(n6067), .A1(n8669), .B0(P2_REG3_REG_4__SCAN_IN), .B1(P2_U3151), .Y(n8855));
  OAI21X1 g7676(.A0(n8854), .A1(n8767), .B0(n8855), .Y(n8856));
  AOI21X1 g7677(.A0(n8659), .A1(n6054), .B0(n8856), .Y(n8857));
  OAI21X1 g7678(.A0(n8852), .A1(n8647), .B0(n8857), .Y(P2_U3170));
  XOR2X1  g7679(.A(n8674), .B(n6916), .Y(n8859));
  INVX1   g7680(.A(n8675), .Y(n8860));
  AOI21X1 g7681(.A0(n8722), .A1(n8860), .B0(n8718), .Y(n8861));
  AOI21X1 g7682(.A0(n8859), .A1(n8718), .B0(n8861), .Y(n8862));
  AOI22X1 g7683(.A0(n6914), .A1(n8640), .B0(n6878), .B1(n8664), .Y(n8863));
  OAI21X1 g7684(.A0(n8662), .A1(n6959), .B0(n8863), .Y(n8864));
  AOI22X1 g7685(.A0(n8660), .A1(n8864), .B0(P2_REG3_REG_24__SCAN_IN), .B1(P2_U3151), .Y(n8865));
  OAI21X1 g7686(.A0(n8658), .A1(n6913), .B0(n8865), .Y(n8866));
  AOI21X1 g7687(.A0(n8669), .A1(n6946), .B0(n8866), .Y(n8867));
  OAI21X1 g7688(.A0(n8862), .A1(n8647), .B0(n8867), .Y(P2_U3169));
  INVX1   g7689(.A(n8705), .Y(n8869));
  OAI21X1 g7690(.A0(n8697), .A1(n6691), .B0(n8698), .Y(n8870));
  AOI21X1 g7691(.A0(n8707), .A1(n8869), .B0(n8870), .Y(n8871));
  AOI22X1 g7692(.A0(n8702), .A1(n8704), .B0(n8696), .B1(n6599), .Y(n8872));
  INVX1   g7693(.A(n8697), .Y(n8873));
  AOI21X1 g7694(.A0(n8873), .A1(n6691), .B0(n8706), .Y(n8874));
  OAI21X1 g7695(.A0(n8873), .A1(n6691), .B0(n8874), .Y(n8875));
  OAI21X1 g7696(.A0(n8875), .A1(n8872), .B0(n8774), .Y(n8876));
  OAI22X1 g7697(.A0(n7367), .A1(n8639), .B0(n6599), .B1(n8665), .Y(n8877));
  AOI21X1 g7698(.A0(n8661), .A1(n6684), .B0(n8877), .Y(n8878));
  AOI22X1 g7699(.A0(n6658), .A1(n8669), .B0(P2_REG3_REG_17__SCAN_IN), .B1(P2_U3151), .Y(n8879));
  OAI21X1 g7700(.A0(n8878), .A1(n8767), .B0(n8879), .Y(n8880));
  AOI21X1 g7701(.A0(n8659), .A1(n6643), .B0(n8880), .Y(n8881));
  OAI21X1 g7702(.A0(n8876), .A1(n8871), .B0(n8881), .Y(P2_U3168));
  XOR2X1  g7703(.A(n8616), .B(n6098), .Y(n8883));
  XOR2X1  g7704(.A(n8883), .B(n8609), .Y(n8884));
  NOR2X1  g7705(.A(n8662), .B(n6156), .Y(n8885));
  OAI22X1 g7706(.A0(n6095), .A1(n8639), .B0(n6104), .B1(n8665), .Y(n8886));
  OAI21X1 g7707(.A0(n8886), .A1(n8885), .B0(n8660), .Y(n8887));
  AOI22X1 g7708(.A0(n6123), .A1(n8669), .B0(P2_REG3_REG_5__SCAN_IN), .B1(P2_U3151), .Y(n8888));
  NAND2X1 g7709(.A(n8888), .B(n8887), .Y(n8889));
  AOI21X1 g7710(.A0(n8659), .A1(n6096), .B0(n8889), .Y(n8890));
  OAI21X1 g7711(.A0(n8884), .A1(n8647), .B0(n8890), .Y(P2_U3167));
  XOR2X1  g7712(.A(n8696), .B(n6599), .Y(n8892));
  AOI21X1 g7713(.A0(n8704), .A1(n8702), .B0(n8892), .Y(n8894));
  AOI21X1 g7714(.A0(n8892), .A1(n8869), .B0(n8894), .Y(n8895));
  OAI22X1 g7715(.A0(n6590), .A1(n8639), .B0(n6558), .B1(n8665), .Y(n8896));
  AOI21X1 g7716(.A0(n8661), .A1(n6645), .B0(n8896), .Y(n8897));
  AOI22X1 g7717(.A0(n6604), .A1(n8669), .B0(P2_REG3_REG_16__SCAN_IN), .B1(P2_U3151), .Y(n8898));
  OAI21X1 g7718(.A0(n8897), .A1(n8767), .B0(n8898), .Y(n8899));
  AOI21X1 g7719(.A0(n8659), .A1(n6591), .B0(n8899), .Y(n8900));
  OAI21X1 g7720(.A0(n8895), .A1(n8647), .B0(n8900), .Y(P2_U3166));
  OAI21X1 g7721(.A0(n8718), .A1(n8675), .B0(n8722), .Y(n8902));
  XOR2X1  g7722(.A(n8724), .B(n6953), .Y(n8903));
  NOR2X1  g7723(.A(n8903), .B(n8902), .Y(n8904));
  AOI21X1 g7724(.A0(n8903), .A1(n8902), .B0(n8904), .Y(n8906));
  INVX1   g7725(.A(n6951), .Y(n8907));
  AOI22X1 g7726(.A0(n6951), .A1(n8640), .B0(n6916), .B1(n8664), .Y(n8908));
  OAI21X1 g7727(.A0(n8662), .A1(n6994), .B0(n8908), .Y(n8909));
  AOI22X1 g7728(.A0(n8660), .A1(n8909), .B0(P2_REG3_REG_25__SCAN_IN), .B1(P2_U3151), .Y(n8910));
  OAI21X1 g7729(.A0(n8658), .A1(n8907), .B0(n8910), .Y(n8911));
  AOI21X1 g7730(.A0(n8669), .A1(n6960), .B0(n8911), .Y(n8912));
  OAI21X1 g7731(.A0(n8906), .A1(n8647), .B0(n8912), .Y(P2_U3165));
  XOR2X1  g7732(.A(n8571), .B(n6436), .Y(n8914));
  NOR2X1  g7733(.A(n8914), .B(n8810), .Y(n8916));
  AOI21X1 g7734(.A0(n8914), .A1(n8810), .B0(n8916), .Y(n8917));
  NOR2X1  g7735(.A(n8662), .B(n6480), .Y(n8918));
  OAI22X1 g7736(.A0(n6426), .A1(n8639), .B0(n6412), .B1(n8665), .Y(n8919));
  OAI21X1 g7737(.A0(n8919), .A1(n8918), .B0(n8660), .Y(n8920));
  AOI22X1 g7738(.A0(n6441), .A1(n8669), .B0(P2_REG3_REG_12__SCAN_IN), .B1(P2_U3151), .Y(n8921));
  NAND2X1 g7739(.A(n8921), .B(n8920), .Y(n8922));
  AOI21X1 g7740(.A0(n8659), .A1(n6427), .B0(n8922), .Y(n8923));
  OAI21X1 g7741(.A0(n8917), .A1(n8647), .B0(n8923), .Y(P2_U3164));
  NAND2X1 g7742(.A(n8685), .B(n6767), .Y(n8925));
  OAI21X1 g7743(.A0(n8682), .A1(n6814), .B0(n8687), .Y(n8926));
  AOI21X1 g7744(.A0(n8825), .A1(n8925), .B0(n8926), .Y(n8927));
  OAI21X1 g7745(.A0(n8682), .A1(n6806), .B0(n8925), .Y(n8928));
  AOI21X1 g7746(.A0(n8682), .A1(n6806), .B0(n8928), .Y(n8929));
  OAI21X1 g7747(.A0(n8825), .A1(n8686), .B0(n8929), .Y(n8930));
  NAND2X1 g7748(.A(n8930), .B(n8774), .Y(n8931));
  AOI22X1 g7749(.A0(n6804), .A1(n8640), .B0(n6767), .B1(n8664), .Y(n8932));
  OAI21X1 g7750(.A0(n8662), .A1(n6848), .B0(n8932), .Y(n8933));
  AOI22X1 g7751(.A0(n8660), .A1(n8933), .B0(P2_REG3_REG_21__SCAN_IN), .B1(P2_U3151), .Y(n8934));
  OAI21X1 g7752(.A0(n8658), .A1(n6803), .B0(n8934), .Y(n8935));
  AOI21X1 g7753(.A0(n8669), .A1(n6815), .B0(n8935), .Y(n8936));
  OAI21X1 g7754(.A0(n8931), .A1(n8927), .B0(n8936), .Y(P2_U3163));
  NAND2X1 g7755(.A(n8659), .B(P2_REG3_REG_1__SCAN_IN), .Y(n8938));
  NAND2X1 g7756(.A(n8594), .B(n8592), .Y(n8939));
  XOR2X1  g7757(.A(n8591), .B(n5925), .Y(n8940));
  XOR2X1  g7758(.A(n8940), .B(n8939), .Y(n8941));
  NAND2X1 g7759(.A(n8941), .B(n8774), .Y(n8942));
  AOI22X1 g7760(.A0(n5894), .A1(n8664), .B0(n8640), .B1(P2_REG3_REG_1__SCAN_IN), .Y(n8943));
  OAI21X1 g7761(.A0(n8662), .A1(n5965), .B0(n8943), .Y(n8944));
  NAND2X1 g7762(.A(n8944), .B(n8660), .Y(n8945));
  AOI22X1 g7763(.A0(n5945), .A1(n8669), .B0(P2_REG3_REG_1__SCAN_IN), .B1(P2_U3151), .Y(n8946));
  NAND4X1 g7764(.A(n8945), .B(n8942), .C(n8938), .D(n8946), .Y(P2_U3162));
  AOI21X1 g7765(.A0(n8619), .A1(n8609), .B0(n8626), .Y(n8948));
  XOR2X1  g7766(.A(n8610), .B(n6249), .Y(n8949));
  XOR2X1  g7767(.A(n8949), .B(n8948), .Y(n8950));
  NOR2X1  g7768(.A(n8662), .B(n6296), .Y(n8951));
  OAI22X1 g7769(.A0(n6239), .A1(n8639), .B0(n6206), .B1(n8665), .Y(n8952));
  OAI21X1 g7770(.A0(n8952), .A1(n8951), .B0(n8660), .Y(n8953));
  AOI22X1 g7771(.A0(n6254), .A1(n8669), .B0(P2_REG3_REG_8__SCAN_IN), .B1(P2_U3151), .Y(n8954));
  NAND2X1 g7772(.A(n8954), .B(n8953), .Y(n8955));
  AOI21X1 g7773(.A0(n8659), .A1(n6240), .B0(n8955), .Y(n8956));
  OAI21X1 g7774(.A0(n8950), .A1(n8647), .B0(n8956), .Y(P2_U3161));
  XOR2X1  g7775(.A(n8574), .B(n7034), .Y(n8958));
  INVX1   g7776(.A(n8958), .Y(n8959));
  OAI21X1 g7777(.A0(n8720), .A1(n6994), .B0(n8726), .Y(n8960));
  OAI21X1 g7778(.A0(n8959), .A1(n7023), .B0(n8960), .Y(n8961));
  AOI21X1 g7779(.A0(n8733), .A1(n8730), .B0(n8961), .Y(n8962));
  AOI21X1 g7780(.A0(n8724), .A1(n6959), .B0(n6994), .Y(n8963));
  AOI21X1 g7781(.A0(n8724), .A1(n6959), .B0(n8675), .Y(n8964));
  AOI22X1 g7782(.A0(n8963), .A1(n8860), .B0(n8731), .B1(n8964), .Y(n8965));
  INVX1   g7783(.A(n8965), .Y(n8966));
  OAI21X1 g7784(.A0(n8959), .A1(n7023), .B0(n8966), .Y(n8967));
  XOR2X1  g7785(.A(n8564), .B(n7064), .Y(n8968));
  XOR2X1  g7786(.A(n8968), .B(n7093), .Y(n8969));
  NOR2X1  g7787(.A(n8958), .B(n7074), .Y(n8970));
  NOR2X1  g7788(.A(n8970), .B(n8969), .Y(n8971));
  OAI21X1 g7789(.A0(n8967), .A1(n8718), .B0(n8971), .Y(n8972));
  NOR2X1  g7790(.A(n8965), .B(n8718), .Y(n8973));
  OAI21X1 g7791(.A0(n8733), .A1(n8726), .B0(n8730), .Y(n8974));
  NOR3X1  g7792(.A(n8974), .B(n8973), .C(n8970), .Y(n8975));
  OAI21X1 g7793(.A0(n8959), .A1(n7023), .B0(n8969), .Y(n8976));
  OAI22X1 g7794(.A0(n8975), .A1(n8976), .B0(n8972), .B1(n8962), .Y(n8977));
  NAND2X1 g7795(.A(n8977), .B(n8774), .Y(n8978));
  NAND3X1 g7796(.A(n8669), .B(n6823), .C(n7070), .Y(n8979));
  NOR2X1  g7797(.A(n8658), .B(n7061), .Y(n8980));
  OAI22X1 g7798(.A0(n7061), .A1(n8639), .B0(n7074), .B1(n8665), .Y(n8981));
  AOI21X1 g7799(.A0(n8661), .A1(n7100), .B0(n8981), .Y(n8982));
  OAI22X1 g7800(.A0(n8767), .A1(n8982), .B0(n7060), .B1(P2_STATE_REG_SCAN_IN), .Y(n8983));
  NOR2X1  g7801(.A(n8983), .B(n8980), .Y(n8984));
  NAND3X1 g7802(.A(n8984), .B(n8979), .C(n8978), .Y(P2_U3160));
  XOR2X1  g7803(.A(n8683), .B(n6729), .Y(n8986));
  NOR2X1  g7804(.A(n8986), .B(n8712), .Y(n8987));
  AOI21X1 g7805(.A0(n8986), .A1(n8712), .B0(n8987), .Y(n8989));
  INVX1   g7806(.A(n6727), .Y(n8990));
  AOI22X1 g7807(.A0(n6727), .A1(n8640), .B0(n6684), .B1(n8664), .Y(n8991));
  OAI21X1 g7808(.A0(n8662), .A1(n6773), .B0(n8991), .Y(n8992));
  AOI22X1 g7809(.A0(n8660), .A1(n8992), .B0(P2_REG3_REG_19__SCAN_IN), .B1(P2_U3151), .Y(n8993));
  OAI21X1 g7810(.A0(n8658), .A1(n8990), .B0(n8993), .Y(n8994));
  AOI21X1 g7811(.A0(n8669), .A1(n6737), .B0(n8994), .Y(n8995));
  OAI21X1 g7812(.A0(n8989), .A1(n8647), .B0(n8995), .Y(P2_U3159));
  OAI21X1 g7813(.A0(n8588), .A1(n5965), .B0(n8597), .Y(n8997));
  NAND2X1 g7814(.A(n8601), .B(n6012), .Y(n8998));
  NAND3X1 g7815(.A(n8998), .B(n8997), .C(n8590), .Y(n8999));
  OAI22X1 g7816(.A0(n8588), .A1(n5965), .B0(n6012), .B1(n8589), .Y(n9000));
  AOI21X1 g7817(.A0(n8589), .A1(n6012), .B0(n9000), .Y(n9001));
  OAI21X1 g7818(.A0(n8597), .A1(n8777), .B0(n9001), .Y(n9002));
  NAND3X1 g7819(.A(n9002), .B(n8999), .C(n8774), .Y(n9003));
  NAND2X1 g7820(.A(n8659), .B(n6010), .Y(n9004));
  AOI22X1 g7821(.A0(n7262), .A1(n8664), .B0(n8640), .B1(n6010), .Y(n9005));
  OAI21X1 g7822(.A0(n8662), .A1(n6104), .B0(n9005), .Y(n9006));
  OAI22X1 g7823(.A0(n6024), .A1(n8668), .B0(n6010), .B1(P2_STATE_REG_SCAN_IN), .Y(n9007));
  AOI21X1 g7824(.A0(n9006), .A1(n8660), .B0(n9007), .Y(n9008));
  NAND3X1 g7825(.A(n9008), .B(n9004), .C(n9003), .Y(P2_U3158));
  XOR2X1  g7826(.A(n8565), .B(n6333), .Y(n9010));
  XOR2X1  g7827(.A(n9010), .B(n8634), .Y(n9011));
  AOI22X1 g7828(.A0(n6330), .A1(n8640), .B0(n6284), .B1(n8664), .Y(n9012));
  OAI21X1 g7829(.A0(n8662), .A1(n6412), .B0(n9012), .Y(n9013));
  NAND2X1 g7830(.A(n9013), .B(n8660), .Y(n9014));
  AOI22X1 g7831(.A0(n6353), .A1(n8669), .B0(P2_REG3_REG_10__SCAN_IN), .B1(P2_U3151), .Y(n9015));
  NAND2X1 g7832(.A(n9015), .B(n9014), .Y(n9016));
  AOI21X1 g7833(.A0(n8659), .A1(n6330), .B0(n9016), .Y(n9017));
  OAI21X1 g7834(.A0(n9011), .A1(n8647), .B0(n9017), .Y(P2_U3157));
  XOR2X1  g7835(.A(n8676), .B(n6878), .Y(n9019));
  XOR2X1  g7836(.A(n9019), .B(n8717), .Y(n9020));
  AOI22X1 g7837(.A0(n6876), .A1(n8640), .B0(n6842), .B1(n8664), .Y(n9021));
  OAI21X1 g7838(.A0(n8662), .A1(n6929), .B0(n9021), .Y(n9022));
  AOI22X1 g7839(.A0(n8660), .A1(n9022), .B0(P2_REG3_REG_23__SCAN_IN), .B1(P2_U3151), .Y(n9023));
  OAI21X1 g7840(.A0(n8658), .A1(n7403), .B0(n9023), .Y(n9024));
  AOI21X1 g7841(.A0(n8669), .A1(n6911), .B0(n9024), .Y(n9025));
  OAI21X1 g7842(.A0(n9020), .A1(n8647), .B0(n9025), .Y(P2_U3156));
  NOR3X1  g7843(.A(n8634), .B(n8787), .C(n8577), .Y(n9027));
  NOR2X1  g7844(.A(n9027), .B(n8581), .Y(n9028));
  XOR2X1  g7845(.A(n8582), .B(n6527), .Y(n9029));
  XOR2X1  g7846(.A(n9029), .B(n9028), .Y(n9030));
  NOR2X1  g7847(.A(n8662), .B(n6558), .Y(n9031));
  OAI22X1 g7848(.A0(n6513), .A1(n8639), .B0(n6480), .B1(n8665), .Y(n9032));
  OAI21X1 g7849(.A0(n9032), .A1(n9031), .B0(n8660), .Y(n9033));
  AOI22X1 g7850(.A0(n6532), .A1(n8669), .B0(P2_REG3_REG_14__SCAN_IN), .B1(P2_U3151), .Y(n9034));
  NAND2X1 g7851(.A(n9034), .B(n9033), .Y(n9035));
  AOI21X1 g7852(.A0(n8659), .A1(n6514), .B0(n9035), .Y(n9036));
  OAI21X1 g7853(.A0(n9030), .A1(n8647), .B0(n9036), .Y(P2_U3155));
  NOR2X1  g7854(.A(n8974), .B(n8973), .Y(n9038));
  XOR2X1  g7855(.A(n8958), .B(n7074), .Y(n9039));
  XOR2X1  g7856(.A(n9039), .B(n9038), .Y(n9040));
  AOI22X1 g7857(.A0(n7021), .A1(n8640), .B0(n6987), .B1(n8664), .Y(n9041));
  OAI21X1 g7858(.A0(n8662), .A1(n7111), .B0(n9041), .Y(n9042));
  AOI22X1 g7859(.A0(n8660), .A1(n9042), .B0(P2_REG3_REG_27__SCAN_IN), .B1(P2_U3151), .Y(n9043));
  OAI21X1 g7860(.A0(n8658), .A1(n7432), .B0(n9043), .Y(n9044));
  AOI21X1 g7861(.A0(n8669), .A1(n7058), .B0(n9044), .Y(n9045));
  OAI21X1 g7862(.A0(n9040), .A1(n8647), .B0(n9045), .Y(P2_U3154));
  INVX1   g7863(.A(n8753), .Y(n9047));
  NOR2X1  g7864(.A(n9047), .B(n8622), .Y(n9048));
  OAI21X1 g7865(.A0(n8613), .A1(n6206), .B0(n8614), .Y(n9049));
  INVX1   g7866(.A(n8612), .Y(n9050));
  OAI21X1 g7867(.A0(n9050), .A1(n6150), .B0(n9047), .Y(n9051));
  OAI22X1 g7868(.A0(n8612), .A1(n6156), .B0(n6200), .B1(n8613), .Y(n9052));
  AOI21X1 g7869(.A0(n8613), .A1(n6200), .B0(n9052), .Y(n9053));
  AOI21X1 g7870(.A0(n9053), .A1(n9051), .B0(n8647), .Y(n9054));
  OAI21X1 g7871(.A0(n9049), .A1(n9048), .B0(n9054), .Y(n9055));
  NAND2X1 g7872(.A(n8659), .B(n6198), .Y(n9056));
  AOI22X1 g7873(.A0(n6198), .A1(n8640), .B0(n6150), .B1(n8664), .Y(n9057));
  OAI21X1 g7874(.A0(n8662), .A1(n6249), .B0(n9057), .Y(n9058));
  OAI22X1 g7875(.A0(n6222), .A1(n8668), .B0(n6196), .B1(P2_STATE_REG_SCAN_IN), .Y(n9059));
  AOI21X1 g7876(.A0(n9058), .A1(n8660), .B0(n9059), .Y(n9060));
  NAND3X1 g7877(.A(n9060), .B(n9056), .C(n9055), .Y(P2_U3153));
  INVX1   g7878(.A(n8653), .Y(n9062));
  AOI21X1 g7879(.A0(n6823), .A1(n5729), .B0(P2_U3151), .Y(n9063));
  OAI21X1 g7880(.A0(n7458), .A1(n9062), .B0(n9063), .Y(P2_U3150));
endmodule


