//Converted to Combinational (Partial output: n460) , Module name: s15850_n460
module s15850_n460 ( g1822, g1882, g1834, g1814, g1828, g1840, g1936, g1945, g1864, g1868, g1861, g1872, g1887, g1845, g1857, g1900, g1891, g1927, g1918, g1909, n460 );
input g1822, g1882, g1834, g1814, g1828, g1840, g1936, g1945, g1864, g1868, g1861, g1872, g1887, g1845, g1857, g1900, g1891, g1927, g1918, g1909;
output n460;
wire n2348, n2330, n2342, n2347, n2345, n2346_1, n2341_1, n2320, n2329, n2306_1, n2331_1, n2313, n2343, n2344, n2314, n2337, n2340, n2319, n2328, n2312, n2308, n2311_1, n2336_1, n2326_1, n2339, n2318, n2327, n2321_1, n2307, n2309, n2310, n2335, n2332, n2333, n2334, n2325, n2324, n2338, n2317, n2322, n2323, n2315, n2316_1;
OAI21X1  g0512(.A0(n2342), .A1(n2330), .B0(n2348), .Y(n460));
NAND4X1  g0511(.A(n2341_1), .B(n2346_1), .C(n2345), .D(n2347), .Y(n2348));
MX2X1    g0493(.A(n2306_1), .B(n2329), .S0(n2320), .Y(n2330));
OR2X1    g0505(.A(n2341_1), .B(n2331_1), .Y(n2342));
AOI21X1  g0510(.A0(n2343), .A1(g1822), .B0(n2313), .Y(n2347));
INVX1    g0508(.A(n2344), .Y(n2345));
INVX1    g0509(.A(n2331_1), .Y(n2346_1));
AOI21X1  g0504(.A0(n2340), .A1(n2337), .B0(n2314), .Y(n2341_1));
NAND2X1  g0483(.A(n2319), .B(n2314), .Y(n2320));
XOR2X1   g0492(.A(n2328), .B(g1882), .Y(n2329));
INVX1    g0469(.A(g1882), .Y(n2306_1));
NOR4X1   g0494(.A(g1828), .B(g1822), .C(g1814), .D(g1834), .Y(n2331_1));
NOR2X1   g0476(.A(n2312), .B(g1840), .Y(n2313));
INVX1    g0506(.A(g1828), .Y(n2343));
NOR3X1   g0507(.A(n2343), .B(g1822), .C(g1814), .Y(n2344));
OAI21X1  g0477(.A0(n2313), .A1(n2311_1), .B0(n2308), .Y(n2314));
OR4X1    g0500(.A(n2326_1), .B(g1945), .C(g1936), .D(n2336_1), .Y(n2337));
NAND4X1  g0503(.A(n2326_1), .B(g1945), .C(g1936), .D(n2339), .Y(n2340));
OAI21X1  g0482(.A0(n2318), .A1(g1840), .B0(n2308), .Y(n2319));
MX2X1    g0491(.A(n2321_1), .B(n2327), .S0(n2319), .Y(n2328));
NAND2X1  g0475(.A(g1834), .B(g1814), .Y(n2312));
NOR4X1   g0471(.A(g1861), .B(g1868), .C(g1864), .D(n2307), .Y(n2308));
NOR2X1   g0474(.A(n2310), .B(n2309), .Y(n2311_1));
NAND4X1  g0499(.A(n2334), .B(n2333), .C(n2332), .D(n2335), .Y(n2336_1));
OAI21X1  g0489(.A0(n2324), .A1(g1828), .B0(n2325), .Y(n2326_1));
NOR4X1   g0502(.A(n2334), .B(n2333), .C(n2332), .D(n2338), .Y(n2339));
INVX1    g0481(.A(n2317), .Y(n2318));
XOR2X1   g0490(.A(n2326_1), .B(g1872), .Y(n2327));
INVX1    g0484(.A(g1887), .Y(n2321_1));
INVX1    g0470(.A(g1845), .Y(n2307));
INVX1    g0472(.A(g1857), .Y(n2309));
NOR2X1   g0473(.A(g1828), .B(g1822), .Y(n2310));
NOR4X1   g0498(.A(g1891), .B(g1900), .C(g1882), .D(g1872), .Y(n2335));
INVX1    g0495(.A(g1927), .Y(n2332));
INVX1    g0496(.A(g1918), .Y(n2333));
INVX1    g0497(.A(g1909), .Y(n2334));
OAI21X1  g0488(.A0(g1828), .A1(g1814), .B0(n2322), .Y(n2325));
INVX1    g0487(.A(n2323), .Y(n2324));
NAND4X1  g0501(.A(g1891), .B(g1900), .C(g1882), .D(g1872), .Y(n2338));
NAND4X1  g0480(.A(n2316_1), .B(g1814), .C(n2315), .D(n2310), .Y(n2317));
INVX1    g0485(.A(g1822), .Y(n2322));
NOR2X1   g0486(.A(n2322), .B(g1814), .Y(n2323));
INVX1    g0478(.A(g1840), .Y(n2315));
INVX1    g0479(.A(g1834), .Y(n2316_1));

endmodule
