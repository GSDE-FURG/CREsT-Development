//Converted to Combinational , Module name: s35932 , Timestamp: 2018-12-03T15:51:08.347404 
module s35932 ( DATA_0_31, DATA_0_30, DATA_0_29, DATA_0_28, DATA_0_27, DATA_0_26, DATA_0_25, DATA_0_24, DATA_0_23, DATA_0_22, DATA_0_21, DATA_0_20, DATA_0_19, DATA_0_18, DATA_0_17, DATA_0_16, DATA_0_15, DATA_0_14, DATA_0_13, DATA_0_12, DATA_0_11, DATA_0_10, DATA_0_9, DATA_0_8, DATA_0_7, DATA_0_6, DATA_0_5, DATA_0_4, DATA_0_0, RESET, TM1, TM0, WX485, WX487, WX489, WX491, WX493, WX495, WX497, WX499, WX501, WX503, WX505, WX507, WX509, WX511, WX513, WX515, WX517, WX519, WX521, WX523, WX525, WX527, WX529, WX531, WX533, WX535, WX537, WX539, WX541, WX543, WX545, WX547, WX645, WX647, WX649, WX651, WX653, WX655, WX657, WX659, WX661, WX663, WX665, WX667, WX669, WX671, WX673, WX675, WX677, WX679, WX681, WX683, WX685, WX687, WX689, WX691, WX693, WX695, WX697, WX699, WX701, WX703, WX705, WX707, WX709, WX711, WX713, WX715, WX717, WX719, WX721, WX723, WX725, WX727, WX729, WX731, WX733, WX735, WX737, WX739, WX741, WX743, WX745, WX747, WX749, WX751, WX753, WX755, WX757, WX759, WX761, WX763, WX765, WX767, WX769, WX771, WX773, WX775, WX777, WX779, WX781, WX783, WX785, WX787, WX789, WX791, WX793, WX795, WX797, WX799, WX801, WX803, WX805, WX807, WX809, WX811, WX813, WX815, WX817, WX819, WX821, WX823, WX825, WX827, WX829, WX831, WX833, WX835, WX837, WX839, WX841, WX843, WX845, WX847, WX849, WX851, WX853, WX855, WX857, WX859, WX861, WX863, WX865, WX867, WX869, WX871, WX873, WX875, WX877, WX879, WX881, WX883, WX885, WX887, WX889, WX891, WX893, WX895, WX897, WX899, WX1778, WX1780, WX1782, WX1784, WX1786, WX1788, WX1790, WX1792, WX1794, WX1796, WX1798, WX1800, WX1802, WX1804, WX1806, WX1808, WX1810, WX1812, WX1814, WX1816, WX1818, WX1820, WX1822, WX1824, WX1826, WX1828, WX1830, WX1832, WX1834, WX1836, WX1838, WX1840, WX1938, WX1940, WX1942, WX1944, WX1946, WX1948, WX1950, WX1952, WX1954, WX1956, WX1958, WX1960, WX1962, WX1964, WX1966, WX1968, WX1970, WX1972, WX1974, WX1976, WX1978, WX1980, WX1982, WX1984, WX1986, WX1988, WX1990, WX1992, WX1994, WX1996, WX1998, WX2000, WX2002, WX2004, WX2006, WX2008, WX2010, WX2012, WX2014, WX2016, WX2018, WX2020, WX2022, WX2024, WX2026, WX2028, WX2030, WX2032, WX2034, WX2036, WX2038, WX2040, WX2042, WX2044, WX2046, WX2048, WX2050, WX2052, WX2054, WX2056, WX2058, WX2060, WX2062, WX2064, WX2066, WX2068, WX2070, WX2072, WX2074, WX2076, WX2078, WX2080, WX2082, WX2084, WX2086, WX2088, WX2090, WX2092, WX2094, WX2096, WX2098, WX2100, WX2102, WX2104, WX2106, WX2108, WX2110, WX2112, WX2114, WX2116, WX2118, WX2120, WX2122, WX2124, WX2126, WX2128, WX2130, WX2132, WX2134, WX2136, WX2138, WX2140, WX2142, WX2144, WX2146, WX2148, WX2150, WX2152, WX2154, WX2156, WX2158, WX2160, WX2162, WX2164, WX2166, WX2168, WX2170, WX2172, WX2174, WX2176, WX2178, WX2180, WX2182, WX2184, WX2186, WX2188, WX2190, WX2192, WX3071, WX3073, WX3075, WX3077, WX3079, WX3081, WX3083, WX3085, WX3087, WX3089, WX3091, WX3093, WX3095, WX3097, WX3099, WX3101, WX3103, WX3105, WX3107, WX3109, WX3111, WX3113, WX3115, WX3117, WX3119, WX3121, WX3123, WX3125, WX3127, WX3129, WX3131, WX3133, WX3231, WX3233, WX3235, WX3237, WX3239, WX3241, WX3243, WX3245, WX3247, WX3249, WX3251, WX3253, WX3255, WX3257, WX3259, WX3261, WX3263, WX3265, WX3267, WX3269, WX3271, WX3273, WX3275, WX3277, WX3279, WX3281, WX3283, WX3285, WX3287, WX3289, WX3291, WX3293, WX3295, WX3297, WX3299, WX3301, WX3303, WX3305, WX3307, WX3309, WX3311, WX3313, WX3315, WX3317, WX3319, WX3321, WX3323, WX3325, WX3327, WX3329, WX3331, WX3333, WX3335, WX3337, WX3339, WX3341, WX3343, WX3345, WX3347, WX3349, WX3351, WX3353, WX3355, WX3357, WX3359, WX3361, WX3363, WX3365, WX3367, WX3369, WX3371, WX3373, WX3375, WX3377, WX3379, WX3381, WX3383, WX3385, WX3387, WX3389, WX3391, WX3393, WX3395, WX3397, WX3399, WX3401, WX3403, WX3405, WX3407, WX3409, WX3411, WX3413, WX3415, WX3417, WX3419, WX3421, WX3423, WX3425, WX3427, WX3429, WX3431, WX3433, WX3435, WX3437, WX3439, WX3441, WX3443, WX3445, WX3447, WX3449, WX3451, WX3453, WX3455, WX3457, WX3459, WX3461, WX3463, WX3465, WX3467, WX3469, WX3471, WX3473, WX3475, WX3477, WX3479, WX3481, WX3483, WX3485, WX4364, WX4366, WX4368, WX4370, WX4372, WX4374, WX4376, WX4378, WX4380, WX4382, WX4384, WX4386, WX4388, WX4390, WX4392, WX4394, WX4396, WX4398, WX4400, WX4402, WX4404, WX4406, WX4408, WX4410, WX4412, WX4414, WX4416, WX4418, WX4420, WX4422, WX4424, WX4426, WX4524, WX4526, WX4528, WX4530, WX4532, WX4534, WX4536, WX4538, WX4540, WX4542, WX4544, WX4546, WX4548, WX4550, WX4552, WX4554, WX4556, WX4558, WX4560, WX4562, WX4564, WX4566, WX4568, WX4570, WX4572, WX4574, WX4576, WX4578, WX4580, WX4582, WX4584, WX4586, WX4588, WX4590, WX4592, WX4594, WX4596, WX4598, WX4600, WX4602, WX4604, WX4606, WX4608, WX4610, WX4612, WX4614, WX4616, WX4618, WX4620, WX4622, WX4624, WX4626, WX4628, WX4630, WX4632, WX4634, WX4636, WX4638, WX4640, WX4642, WX4644, WX4646, WX4648, WX4650, WX4652, WX4654, WX4656, WX4658, WX4660, WX4662, WX4664, WX4666, WX4668, WX4670, WX4672, WX4674, WX4676, WX4678, WX4680, WX4682, WX4684, WX4686, WX4688, WX4690, WX4692, WX4694, WX4696, WX4698, WX4700, WX4702, WX4704, WX4706, WX4708, WX4710, WX4712, WX4714, WX4716, WX4718, WX4720, WX4722, WX4724, WX4726, WX4728, WX4730, WX4732, WX4734, WX4736, WX4738, WX4740, WX4742, WX4744, WX4746, WX4748, WX4750, WX4752, WX4754, WX4756, WX4758, WX4760, WX4762, WX4764, WX4766, WX4768, WX4770, WX4772, WX4774, WX4776, WX4778, WX5657, WX5659, WX5661, WX5663, WX5665, WX5667, WX5669, WX5671, WX5673, WX5675, WX5677, WX5679, WX5681, WX5683, WX5685, WX5687, WX5689, WX5691, WX5693, WX5695, WX5697, WX5699, WX5701, WX5703, WX5705, WX5707, WX5709, WX5711, WX5713, WX5715, WX5717, WX5719, WX5817, WX5819, WX5821, WX5823, WX5825, WX5827, WX5829, WX5831, WX5833, WX5835, WX5837, WX5839, WX5841, WX5843, WX5845, WX5847, WX5849, WX5851, WX5853, WX5855, WX5857, WX5859, WX5861, WX5863, WX5865, WX5867, WX5869, WX5871, WX5873, WX5875, WX5877, WX5879, WX5881, WX5883, WX5885, WX5887, WX5889, WX5891, WX5893, WX5895, WX5897, WX5899, WX5901, WX5903, WX5905, WX5907, WX5909, WX5911, WX5913, WX5915, WX5917, WX5919, WX5921, WX5923, WX5925, WX5927, WX5929, WX5931, WX5933, WX5935, WX5937, WX5939, WX5941, WX5943, WX5945, WX5947, WX5949, WX5951, WX5953, WX5955, WX5957, WX5959, WX5961, WX5963, WX5965, WX5967, WX5969, WX5971, WX5973, WX5975, WX5977, WX5979, WX5981, WX5983, WX5985, WX5987, WX5989, WX5991, WX5993, WX5995, WX5997, WX5999, WX6001, WX6003, WX6005, WX6007, WX6009, WX6011, WX6013, WX6015, WX6017, WX6019, WX6021, WX6023, WX6025, WX6027, WX6029, WX6031, WX6033, WX6035, WX6037, WX6039, WX6041, WX6043, WX6045, WX6047, WX6049, WX6051, WX6053, WX6055, WX6057, WX6059, WX6061, WX6063, WX6065, WX6067, WX6069, WX6071, WX6950, WX6952, WX6954, WX6956, WX6958, WX6960, WX6962, WX6964, WX6966, WX6968, WX6970, WX6972, WX6974, WX6976, WX6978, WX6980, WX6982, WX6984, WX6986, WX6988, WX6990, WX6992, WX6994, WX6996, WX6998, WX7000, WX7002, WX7004, WX7006, WX7008, WX7010, WX7012, WX7110, WX7112, WX7114, WX7116, WX7118, WX7120, WX7122, WX7124, WX7126, WX7128, WX7130, WX7132, WX7134, WX7136, WX7138, WX7140, WX7142, WX7144, WX7146, WX7148, WX7150, WX7152, WX7154, WX7156, WX7158, WX7160, WX7162, WX7164, WX7166, WX7168, WX7170, WX7172, WX7174, WX7176, WX7178, WX7180, WX7182, WX7184, WX7186, WX7188, WX7190, WX7192, WX7194, WX7196, WX7198, WX7200, WX7202, WX7204, WX7206, WX7208, WX7210, WX7212, WX7214, WX7216, WX7218, WX7220, WX7222, WX7224, WX7226, WX7228, WX7230, WX7232, WX7234, WX7236, WX7238, WX7240, WX7242, WX7244, WX7246, WX7248, WX7250, WX7252, WX7254, WX7256, WX7258, WX7260, WX7262, WX7264, WX7266, WX7268, WX7270, WX7272, WX7274, WX7276, WX7278, WX7280, WX7282, WX7284, WX7286, WX7288, WX7290, WX7292, WX7294, WX7296, WX7298, WX7300, WX7302, WX7304, WX7306, WX7308, WX7310, WX7312, WX7314, WX7316, WX7318, WX7320, WX7322, WX7324, WX7326, WX7328, WX7330, WX7332, WX7334, WX7336, WX7338, WX7340, WX7342, WX7344, WX7346, WX7348, WX7350, WX7352, WX7354, WX7356, WX7358, WX7360, WX7362, WX7364, WX8243, WX8245, WX8247, WX8249, WX8251, WX8253, WX8255, WX8257, WX8259, WX8261, WX8263, WX8265, WX8267, WX8269, WX8271, WX8273, WX8275, WX8277, WX8279, WX8281, WX8283, WX8285, WX8287, WX8289, WX8291, WX8293, WX8295, WX8297, WX8299, WX8301, WX8303, WX8305, WX8403, WX8405, WX8407, WX8409, WX8411, WX8413, WX8415, WX8417, WX8419, WX8421, WX8423, WX8425, WX8427, WX8429, WX8431, WX8433, WX8435, WX8437, WX8439, WX8441, WX8443, WX8445, WX8447, WX8449, WX8451, WX8453, WX8455, WX8457, WX8459, WX8461, WX8463, WX8465, WX8467, WX8469, WX8471, WX8473, WX8475, WX8477, WX8479, WX8481, WX8483, WX8485, WX8487, WX8489, WX8491, WX8493, WX8495, WX8497, WX8499, WX8501, WX8503, WX8505, WX8507, WX8509, WX8511, WX8513, WX8515, WX8517, WX8519, WX8521, WX8523, WX8525, WX8527, WX8529, WX8531, WX8533, WX8535, WX8537, WX8539, WX8541, WX8543, WX8545, WX8547, WX8549, WX8551, WX8553, WX8555, WX8557, WX8559, WX8561, WX8563, WX8565, WX8567, WX8569, WX8571, WX8573, WX8575, WX8577, WX8579, WX8581, WX8583, WX8585, WX8587, WX8589, WX8591, WX8593, WX8595, WX8597, WX8599, WX8601, WX8603, WX8605, WX8607, WX8609, WX8611, WX8613, WX8615, WX8617, WX8619, WX8621, WX8623, WX8625, WX8627, WX8629, WX8631, WX8633, WX8635, WX8637, WX8639, WX8641, WX8643, WX8645, WX8647, WX8649, WX8651, WX8653, WX8655, WX8657, WX9536, WX9538, WX9540, WX9542, WX9544, WX9546, WX9548, WX9550, WX9552, WX9554, WX9556, WX9558, WX9560, WX9562, WX9564, WX9566, WX9568, WX9570, WX9572, WX9574, WX9576, WX9578, WX9580, WX9582, WX9584, WX9586, WX9588, WX9590, WX9592, WX9594, WX9596, WX9598, WX9696, WX9698, WX9700, WX9702, WX9704, WX9706, WX9708, WX9710, WX9712, WX9714, WX9716, WX9718, WX9720, WX9722, WX9724, WX9726, WX9728, WX9730, WX9732, WX9734, WX9736, WX9738, WX9740, WX9742, WX9744, WX9746, WX9748, WX9750, WX9752, WX9754, WX9756, WX9758, WX9760, WX9762, WX9764, WX9766, WX9768, WX9770, WX9772, WX9774, WX9776, WX9778, WX9780, WX9782, WX9784, WX9786, WX9788, WX9790, WX9792, WX9794, WX9796, WX9798, WX9800, WX9802, WX9804, WX9806, WX9808, WX9810, WX9812, WX9814, WX9816, WX9818, WX9820, WX9822, WX9824, WX9826, WX9828, WX9830, WX9832, WX9834, WX9836, WX9838, WX9840, WX9842, WX9844, WX9846, WX9848, WX9850, WX9852, WX9854, WX9856, WX9858, WX9860, WX9862, WX9864, WX9866, WX9868, WX9870, WX9872, WX9874, WX9876, WX9878, WX9880, WX9882, WX9884, WX9886, WX9888, WX9890, WX9892, WX9894, WX9896, WX9898, WX9900, WX9902, WX9904, WX9906, WX9908, WX9910, WX9912, WX9914, WX9916, WX9918, WX9920, WX9922, WX9924, WX9926, WX9928, WX9930, WX9932, WX9934, WX9936, WX9938, WX9940, WX9942, WX9944, WX9946, WX9948, WX9950, WX10829, WX10831, WX10833, WX10835, WX10837, WX10839, WX10841, WX10843, WX10845, WX10847, WX10849, WX10851, WX10853, WX10855, WX10857, WX10859, WX10861, WX10863, WX10865, WX10867, WX10869, WX10871, WX10873, WX10875, WX10877, WX10879, WX10881, WX10883, WX10885, WX10887, WX10889, WX10891, WX10989, WX10991, WX10993, WX10995, WX10997, WX10999, WX11001, WX11003, WX11005, WX11007, WX11009, WX11011, WX11013, WX11015, WX11017, WX11019, WX11021, WX11023, WX11025, WX11027, WX11029, WX11031, WX11033, WX11035, WX11037, WX11039, WX11041, WX11043, WX11045, WX11047, WX11049, WX11051, WX11053, WX11055, WX11057, WX11059, WX11061, WX11063, WX11065, WX11067, WX11069, WX11071, WX11073, WX11075, WX11077, WX11079, WX11081, WX11083, WX11085, WX11087, WX11089, WX11091, WX11093, WX11095, WX11097, WX11099, WX11101, WX11103, WX11105, WX11107, WX11109, WX11111, WX11113, WX11115, WX11117, WX11119, WX11121, WX11123, WX11125, WX11127, WX11129, WX11131, WX11133, WX11135, WX11137, WX11139, WX11141, WX11143, WX11145, WX11147, WX11149, WX11151, WX11153, WX11155, WX11157, WX11159, WX11161, WX11163, WX11165, WX11167, WX11169, WX11171, WX11173, WX11175, WX11177, WX11179, WX11181, WX11183, WX11185, WX11187, WX11189, WX11191, WX11193, WX11195, WX11197, WX11199, WX11201, WX11203, WX11205, WX11207, WX11209, WX11211, WX11213, WX11215, WX11217, WX11219, WX11221, WX11223, WX11225, WX11227, WX11229, WX11231, WX11233, WX11235, WX11237, WX11239, WX11241, WX11243, DATA_9_31, DATA_9_30, DATA_9_29, DATA_9_28, DATA_9_27, DATA_9_26, DATA_9_25, DATA_9_24, DATA_9_23, DATA_9_22, DATA_9_21, DATA_9_20, DATA_9_19, DATA_9_18, DATA_9_17, DATA_9_16, DATA_9_15, DATA_9_14, DATA_9_13, DATA_9_12, DATA_9_11, DATA_9_10, DATA_9_9, DATA_9_8, DATA_9_7, DATA_9_6, DATA_9_5, DATA_9_4, DATA_9_0, CRC_OUT_9_0, CRC_OUT_9_1, CRC_OUT_9_2, CRC_OUT_9_3, CRC_OUT_9_4, CRC_OUT_9_5, CRC_OUT_9_6, CRC_OUT_9_7, CRC_OUT_9_8, CRC_OUT_9_9, CRC_OUT_9_10, CRC_OUT_9_11, CRC_OUT_9_12, CRC_OUT_9_13, CRC_OUT_9_14, CRC_OUT_9_15, CRC_OUT_9_16, CRC_OUT_9_17, CRC_OUT_9_18, CRC_OUT_9_19, CRC_OUT_9_20, CRC_OUT_9_21, CRC_OUT_9_22, CRC_OUT_9_23, CRC_OUT_9_24, CRC_OUT_9_25, CRC_OUT_9_26, CRC_OUT_9_27, CRC_OUT_9_28, CRC_OUT_9_29, CRC_OUT_9_30, CRC_OUT_9_31, CRC_OUT_8_0, CRC_OUT_8_1, CRC_OUT_8_2, CRC_OUT_8_3, CRC_OUT_8_4, CRC_OUT_8_5, CRC_OUT_8_6, CRC_OUT_8_7, CRC_OUT_8_8, CRC_OUT_8_9, CRC_OUT_8_10, CRC_OUT_8_11, CRC_OUT_8_12, CRC_OUT_8_13, CRC_OUT_8_14, CRC_OUT_8_15, CRC_OUT_8_16, CRC_OUT_8_17, CRC_OUT_8_18, CRC_OUT_8_19, CRC_OUT_8_20, CRC_OUT_8_21, CRC_OUT_8_22, CRC_OUT_8_23, CRC_OUT_8_24, CRC_OUT_8_25, CRC_OUT_8_26, CRC_OUT_8_27, CRC_OUT_8_28, CRC_OUT_8_29, CRC_OUT_8_30, CRC_OUT_8_31, CRC_OUT_7_0, CRC_OUT_7_1, CRC_OUT_7_2, CRC_OUT_7_3, CRC_OUT_7_4, CRC_OUT_7_5, CRC_OUT_7_6, CRC_OUT_7_7, CRC_OUT_7_8, CRC_OUT_7_9, CRC_OUT_7_10, CRC_OUT_7_11, CRC_OUT_7_12, CRC_OUT_7_13, CRC_OUT_7_14, CRC_OUT_7_15, CRC_OUT_7_16, CRC_OUT_7_17, CRC_OUT_7_18, CRC_OUT_7_19, CRC_OUT_7_20, CRC_OUT_7_21, CRC_OUT_7_22, CRC_OUT_7_23, CRC_OUT_7_24, CRC_OUT_7_25, CRC_OUT_7_26, CRC_OUT_7_27, CRC_OUT_7_28, CRC_OUT_7_29, CRC_OUT_7_30, CRC_OUT_7_31, CRC_OUT_6_0, CRC_OUT_6_1, CRC_OUT_6_2, CRC_OUT_6_3, CRC_OUT_6_4, CRC_OUT_6_5, CRC_OUT_6_6, CRC_OUT_6_7, CRC_OUT_6_8, CRC_OUT_6_9, CRC_OUT_6_10, CRC_OUT_6_11, CRC_OUT_6_12, CRC_OUT_6_13, CRC_OUT_6_14, CRC_OUT_6_15, CRC_OUT_6_16, CRC_OUT_6_17, CRC_OUT_6_18, CRC_OUT_6_19, CRC_OUT_6_20, CRC_OUT_6_21, CRC_OUT_6_22, CRC_OUT_6_23, CRC_OUT_6_24, CRC_OUT_6_25, CRC_OUT_6_26, CRC_OUT_6_27, CRC_OUT_6_28, CRC_OUT_6_29, CRC_OUT_6_30, CRC_OUT_6_31, CRC_OUT_5_0, CRC_OUT_5_1, CRC_OUT_5_2, CRC_OUT_5_3, CRC_OUT_5_4, CRC_OUT_5_5, CRC_OUT_5_6, CRC_OUT_5_7, CRC_OUT_5_8, CRC_OUT_5_9, CRC_OUT_5_10, CRC_OUT_5_11, CRC_OUT_5_12, CRC_OUT_5_13, CRC_OUT_5_14, CRC_OUT_5_15, CRC_OUT_5_16, CRC_OUT_5_17, CRC_OUT_5_18, CRC_OUT_5_19, CRC_OUT_5_20, CRC_OUT_5_21, CRC_OUT_5_22, CRC_OUT_5_23, CRC_OUT_5_24, CRC_OUT_5_25, CRC_OUT_5_26, CRC_OUT_5_27, CRC_OUT_5_28, CRC_OUT_5_29, CRC_OUT_5_30, CRC_OUT_5_31, CRC_OUT_4_0, CRC_OUT_4_1, CRC_OUT_4_2, CRC_OUT_4_3, CRC_OUT_4_4, CRC_OUT_4_5, CRC_OUT_4_6, CRC_OUT_4_7, CRC_OUT_4_8, CRC_OUT_4_9, CRC_OUT_4_10, CRC_OUT_4_11, CRC_OUT_4_12, CRC_OUT_4_13, CRC_OUT_4_14, CRC_OUT_4_15, CRC_OUT_4_16, CRC_OUT_4_17, CRC_OUT_4_18, CRC_OUT_4_19, CRC_OUT_4_20, CRC_OUT_4_21, CRC_OUT_4_22, CRC_OUT_4_23, CRC_OUT_4_24, CRC_OUT_4_25, CRC_OUT_4_26, CRC_OUT_4_27, CRC_OUT_4_28, CRC_OUT_4_29, CRC_OUT_4_30, CRC_OUT_4_31, CRC_OUT_3_0, CRC_OUT_3_1, CRC_OUT_3_2, CRC_OUT_3_3, CRC_OUT_3_4, CRC_OUT_3_5, CRC_OUT_3_6, CRC_OUT_3_7, CRC_OUT_3_8, CRC_OUT_3_9, CRC_OUT_3_10, CRC_OUT_3_11, CRC_OUT_3_12, CRC_OUT_3_13, CRC_OUT_3_14, CRC_OUT_3_15, CRC_OUT_3_16, CRC_OUT_3_17, CRC_OUT_3_18, CRC_OUT_3_19, CRC_OUT_3_20, CRC_OUT_3_21, CRC_OUT_3_22, CRC_OUT_3_23, CRC_OUT_3_24, CRC_OUT_3_25, CRC_OUT_3_26, CRC_OUT_3_27, CRC_OUT_3_28, CRC_OUT_3_29, CRC_OUT_3_30, CRC_OUT_3_31, CRC_OUT_2_0, CRC_OUT_2_1, CRC_OUT_2_2, CRC_OUT_2_3, CRC_OUT_2_4, CRC_OUT_2_5, CRC_OUT_2_6, CRC_OUT_2_7, CRC_OUT_2_8, CRC_OUT_2_9, CRC_OUT_2_10, CRC_OUT_2_11, CRC_OUT_2_12, CRC_OUT_2_13, CRC_OUT_2_14, CRC_OUT_2_15, CRC_OUT_2_16, CRC_OUT_2_17, CRC_OUT_2_18, CRC_OUT_2_19, CRC_OUT_2_20, CRC_OUT_2_21, CRC_OUT_2_22, CRC_OUT_2_23, CRC_OUT_2_24, CRC_OUT_2_25, CRC_OUT_2_26, CRC_OUT_2_27, CRC_OUT_2_28, CRC_OUT_2_29, CRC_OUT_2_30, CRC_OUT_2_31, CRC_OUT_1_0, CRC_OUT_1_1, CRC_OUT_1_2, CRC_OUT_1_3, CRC_OUT_1_4, CRC_OUT_1_5, CRC_OUT_1_6, CRC_OUT_1_7, CRC_OUT_1_8, CRC_OUT_1_9, CRC_OUT_1_10, CRC_OUT_1_11, CRC_OUT_1_12, CRC_OUT_1_13, CRC_OUT_1_14, CRC_OUT_1_15, CRC_OUT_1_16, CRC_OUT_1_17, CRC_OUT_1_18, CRC_OUT_1_19, CRC_OUT_1_20, CRC_OUT_1_21, CRC_OUT_1_22, CRC_OUT_1_23, CRC_OUT_1_24, CRC_OUT_1_25, CRC_OUT_1_26, CRC_OUT_1_27, CRC_OUT_1_28, CRC_OUT_1_29, CRC_OUT_1_30, CRC_OUT_1_31, n711, n716, n721, n726, n731, n736, n741, n746, n751, n756, n761, n766, n771, n776, n781, n786, n791, n796, n801, n806, n811, n816, n821, n826, n831, n836, n841, n846, n851, n856, n861, n866, n871, n876, n881, n886, n891, n896, n901, n906, n911, n916, n921, n926, n931, n936, n941, n946, n951, n956, n961, n966, n971, n976, n981, n986, n991, n996, n1001, n1006, n1011, n1016, n1021, n1026, n1031, n1036, n1041, n1046, n1051, n1056, n1061, n1066, n1071, n1076, n1081, n1086, n1091, n1096, n1101, n1106, n1111, n1116, n1121, n1126, n1131, n1136, n1141, n1146, n1151, n1156, n1161, n1166, n1171, n1176, n1181, n1186, n1191, n1196, n1201, n1206, n1211, n1216, n1221, n1226, n1231, n1236, n1241, n1246, n1251, n1256, n1261, n1266, n1271, n1276, n1281, n1286, n1291, n1296, n1301, n1306, n1311, n1316, n1321, n1326, n1331, n1336, n1341, n1346, n1351, n1356, n1361, n1366, n1371, n1376, n1381, n1386, n1391, n1396, n1401, n1406, n1411, n1416, n1421, n1426, n1431, n1436, n1441, n1446, n1451, n1456, n1461, n1466, n1471, n1476, n1481, n1486, n1491, n1496, n1501, n1506, n1639, n1644, n1649, n1654, n1659, n1664, n1669, n1674, n1679, n1684, n1689, n1694, n1699, n1704, n1709, n1714, n1719, n1724, n1729, n1734, n1739, n1744, n1749, n1754, n1759, n1764, n1769, n1774, n1779, n1784, n1789, n1794, n1799, n1804, n1809, n1814, n1819, n1824, n1829, n1834, n1839, n1844, n1849, n1854, n1859, n1864, n1869, n1874, n1879, n1884, n1889, n1894, n1899, n1904, n1909, n1914, n1919, n1924, n1929, n1934, n1939, n1944, n1949, n1954, n1959, n1964, n1969, n1974, n1979, n1984, n1989, n1994, n1999, n2004, n2009, n2014, n2019, n2024, n2029, n2034, n2039, n2044, n2049, n2054, n2059, n2064, n2069, n2074, n2079, n2084, n2089, n2094, n2099, n2104, n2109, n2114, n2119, n2124, n2129, n2134, n2139, n2144, n2149, n2154, n2159, n2164, n2169, n2174, n2179, n2184, n2189, n2194, n2199, n2204, n2209, n2214, n2219, n2224, n2229, n2234, n2239, n2244, n2249, n2254, n2259, n2264, n2269, n2274, n2279, n2284, n2289, n2294, n2299, n2304, n2309, n2314, n2319, n2324, n2329, n2334, n2339, n2344, n2349, n2354, n2359, n2364, n2369, n2374, n2379, n2384, n2389, n2394, n2399, n2404, n2409, n2414, n2419, n2424, n2429, n2434, n2567, n2572, n2577, n2582, n2587, n2592, n2597, n2602, n2607, n2612, n2617, n2622, n2627, n2632, n2637, n2642, n2647, n2652, n2657, n2662, n2667, n2672, n2677, n2682, n2687, n2692, n2697, n2702, n2707, n2712, n2717, n2722, n2727, n2732, n2737, n2742, n2747, n2752, n2757, n2762, n2767, n2772, n2777, n2782, n2787, n2792, n2797, n2802, n2807, n2812, n2817, n2822, n2827, n2832, n2837, n2842, n2847, n2852, n2857, n2862, n2867, n2872, n2877, n2882, n2887, n2892, n2897, n2902, n2907, n2912, n2917, n2922, n2927, n2932, n2937, n2942, n2947, n2952, n2957, n2962, n2967, n2972, n2977, n2982, n2987, n2992, n2997, n3002, n3007, n3012, n3017, n3022, n3027, n3032, n3037, n3042, n3047, n3052, n3057, n3062, n3067, n3072, n3077, n3082, n3087, n3092, n3097, n3102, n3107, n3112, n3117, n3122, n3127, n3132, n3137, n3142, n3147, n3152, n3157, n3162, n3167, n3172, n3177, n3182, n3187, n3192, n3197, n3202, n3207, n3212, n3217, n3222, n3227, n3232, n3237, n3242, n3247, n3252, n3257, n3262, n3267, n3272, n3277, n3282, n3287, n3292, n3297, n3302, n3307, n3312, n3317, n3322, n3327, n3332, n3337, n3342, n3347, n3352, n3357, n3362, n3495, n3500, n3505, n3510, n3515, n3520, n3525, n3530, n3535, n3540, n3545, n3550, n3555, n3560, n3565, n3570, n3575, n3580, n3585, n3590, n3595, n3600, n3605, n3610, n3615, n3620, n3625, n3630, n3635, n3640, n3645, n3650, n3655, n3660, n3665, n3670, n3675, n3680, n3685, n3690, n3695, n3700, n3705, n3710, n3715, n3720, n3725, n3730, n3735, n3740, n3745, n3750, n3755, n3760, n3765, n3770, n3775, n3780, n3785, n3790, n3795, n3800, n3805, n3810, n3815, n3820, n3825, n3830, n3835, n3840, n3845, n3850, n3855, n3860, n3865, n3870, n3875, n3880, n3885, n3890, n3895, n3900, n3905, n3910, n3915, n3920, n3925, n3930, n3935, n3940, n3945, n3950, n3955, n3960, n3965, n3970, n3975, n3980, n3985, n3990, n3995, n4000, n4005, n4010, n4015, n4020, n4025, n4030, n4035, n4040, n4045, n4050, n4055, n4060, n4065, n4070, n4075, n4080, n4085, n4090, n4095, n4100, n4105, n4110, n4115, n4120, n4125, n4130, n4135, n4140, n4145, n4150, n4155, n4160, n4165, n4170, n4175, n4180, n4185, n4190, n4195, n4200, n4205, n4210, n4215, n4220, n4225, n4230, n4235, n4240, n4245, n4250, n4255, n4260, n4265, n4270, n4275, n4280, n4285, n4290, n4423, n4428, n4433, n4438, n4443, n4448, n4453, n4458, n4463, n4468, n4473, n4478, n4483, n4488, n4493, n4498, n4503, n4508, n4513, n4518, n4523, n4528, n4533, n4538, n4543, n4548, n4553, n4558, n4563, n4568, n4573, n4578, n4583, n4588, n4593, n4598, n4603, n4608, n4613, n4618, n4623, n4628, n4633, n4638, n4643, n4648, n4653, n4658, n4663, n4668, n4673, n4678, n4683, n4688, n4693, n4698, n4703, n4708, n4713, n4718, n4723, n4728, n4733, n4738, n4743, n4748, n4753, n4758, n4763, n4768, n4773, n4778, n4783, n4788, n4793, n4798, n4803, n4808, n4813, n4818, n4823, n4828, n4833, n4838, n4843, n4848, n4853, n4858, n4863, n4868, n4873, n4878, n4883, n4888, n4893, n4898, n4903, n4908, n4913, n4918, n4923, n4928, n4933, n4938, n4943, n4948, n4953, n4958, n4963, n4968, n4973, n4978, n4983, n4988, n4993, n4998, n5003, n5008, n5013, n5018, n5023, n5028, n5033, n5038, n5043, n5048, n5053, n5058, n5063, n5068, n5073, n5078, n5083, n5088, n5093, n5098, n5103, n5108, n5113, n5118, n5123, n5128, n5133, n5138, n5143, n5148, n5153, n5158, n5163, n5168, n5173, n5178, n5183, n5188, n5193, n5198, n5203, n5208, n5213, n5218, n5351, n5356, n5361, n5366, n5371, n5376, n5381, n5386, n5391, n5396, n5401, n5406, n5411, n5416, n5421, n5426, n5431, n5436, n5441, n5446, n5451, n5456, n5461, n5466, n5471, n5476, n5481, n5486, n5491, n5496, n5501, n5506, n5511, n5516, n5521, n5526, n5531, n5536, n5541, n5546, n5551, n5556, n5561, n5566, n5571, n5576, n5581, n5586, n5591, n5596, n5601, n5606, n5611, n5616, n5621, n5626, n5631, n5636, n5641, n5646, n5651, n5656, n5661, n5666, n5671, n5676, n5681, n5686, n5691, n5696, n5701, n5706, n5711, n5716, n5721, n5726, n5731, n5736, n5741, n5746, n5751, n5756, n5761, n5766, n5771, n5776, n5781, n5786, n5791, n5796, n5801, n5806, n5811, n5816, n5821, n5826, n5831, n5836, n5841, n5846, n5851, n5856, n5861, n5866, n5871, n5876, n5881, n5886, n5891, n5896, n5901, n5906, n5911, n5916, n5921, n5926, n5931, n5936, n5941, n5946, n5951, n5956, n5961, n5966, n5971, n5976, n5981, n5986, n5991, n5996, n6001, n6006, n6011, n6016, n6021, n6026, n6031, n6036, n6041, n6046, n6051, n6056, n6061, n6066, n6071, n6076, n6081, n6086, n6091, n6096, n6101, n6106, n6111, n6116, n6121, n6126, n6131, n6136, n6141, n6146, n6279, n6284, n6289, n6294, n6299, n6304, n6309, n6314, n6319, n6324, n6329, n6334, n6339, n6344, n6349, n6354, n6359, n6364, n6369, n6374, n6379, n6384, n6389, n6394, n6399, n6404, n6409, n6414, n6419, n6424, n6429, n6434, n6439, n6444, n6449, n6454, n6459, n6464, n6469, n6474, n6479, n6484, n6489, n6494, n6499, n6504, n6509, n6514, n6519, n6524, n6529, n6534, n6539, n6544, n6549, n6554, n6559, n6564, n6569, n6574, n6579, n6584, n6589, n6594, n6599, n6604, n6609, n6614, n6619, n6624, n6629, n6634, n6639, n6644, n6649, n6654, n6659, n6664, n6669, n6674, n6679, n6684, n6689, n6694, n6699, n6704, n6709, n6714, n6719, n6724, n6729, n6734, n6739, n6744, n6749, n6754, n6759, n6764, n6769, n6774, n6779, n6784, n6789, n6794, n6799, n6804, n6809, n6814, n6819, n6824, n6829, n6834, n6839, n6844, n6849, n6854, n6859, n6864, n6869, n6874, n6879, n6884, n6889, n6894, n6899, n6904, n6909, n6914, n6919, n6924, n6929, n6934, n6939, n6944, n6949, n6954, n6959, n6964, n6969, n6974, n6979, n6984, n6989, n6994, n6999, n7004, n7009, n7014, n7019, n7024, n7029, n7034, n7039, n7044, n7049, n7054, n7059, n7064, n7069, n7074, n7207, n7212, n7217, n7222, n7227, n7232, n7237, n7242, n7247, n7252, n7257, n7262, n7267, n7272, n7277, n7282, n7287, n7292, n7297, n7302, n7307, n7312, n7317, n7322, n7327, n7332, n7337, n7342, n7347, n7352, n7357, n7362, n7367, n7372, n7377, n7382, n7387, n7392, n7397, n7402, n7407, n7412, n7417, n7422, n7427, n7432, n7437, n7442, n7447, n7452, n7457, n7462, n7467, n7472, n7477, n7482, n7487, n7492, n7497, n7502, n7507, n7512, n7517, n7522, n7527, n7532, n7537, n7542, n7547, n7552, n7557, n7562, n7567, n7572, n7577, n7582, n7587, n7592, n7597, n7602, n7607, n7612, n7617, n7622, n7627, n7632, n7637, n7642, n7647, n7652, n7657, n7662, n7667, n7672, n7677, n7682, n7687, n7692, n7697, n7702, n7707, n7712, n7717, n7722, n7727, n7732, n7737, n7742, n7747, n7752, n7757, n7762, n7767, n7772, n7777, n7782, n7787, n7792, n7797, n7802, n7807, n7812, n7817, n7822, n7827, n7832, n7837, n7842, n7847, n7852, n7857, n7862, n7867, n7872, n7877, n7882, n7887, n7892, n7897, n7902, n7907, n7912, n7917, n7922, n7927, n7932, n7937, n7942, n7947, n7952, n7957, n7962, n7967, n7972, n7977, n7982, n7987, n7992, n7997, n8002, n8135, n8140, n8145, n8150, n8155, n8160, n8165, n8170, n8175, n8180, n8185, n8190, n8195, n8200, n8205, n8210, n8215, n8220, n8225, n8230, n8235, n8240, n8245, n8250, n8255, n8260, n8265, n8270, n8275, n8280, n8285, n8290, n8295, n8300, n8305, n8310, n8315, n8320, n8325, n8330, n8335, n8340, n8345, n8350, n8355, n8360, n8365, n8370, n8375, n8380, n8385, n8390, n8395, n8400, n8405, n8410, n8415, n8420, n8425, n8430, n8435, n8440, n8445, n8450, n8455, n8460, n8465, n8470, n8475, n8480, n8485, n8490, n8495, n8500, n8505, n8510, n8515, n8520, n8525, n8530, n8535, n8540, n8545, n8550, n8555, n8560, n8565, n8570, n8575, n8580, n8585, n8590, n8595, n8600, n8605, n8610, n8615, n8620, n8625, n8630, n8635, n8640, n8645, n8650, n8655, n8660, n8665, n8670, n8675, n8680, n8685, n8690, n8695, n8700, n8705, n8710, n8715, n8720, n8725, n8730, n8735, n8740, n8745, n8750, n8755, n8760, n8765, n8770, n8775, n8780, n8785, n8790, n8795, n8800, n8805, n8810, n8815, n8820, n8825, n8830, n8835, n8840, n8845, n8850, n8855, n8860, n8865, n8870, n8875, n8880, n8885, n8890, n8895, n8900, n8905, n8910, n8915, n8920, n8925, n8930 );
input DATA_0_1, DATA_0_2, DATA_0_3, DATA_0_31, DATA_0_30, DATA_0_29, DATA_0_28, DATA_0_27, DATA_0_26, DATA_0_25, DATA_0_24, DATA_0_23, DATA_0_22, DATA_0_21, DATA_0_20, DATA_0_19, DATA_0_18, DATA_0_17, DATA_0_16, DATA_0_15, DATA_0_14, DATA_0_13, DATA_0_12, DATA_0_11, DATA_0_10, DATA_0_9, DATA_0_8, DATA_0_7, DATA_0_6, DATA_0_5, DATA_0_4, DATA_0_0, RESET, TM1, TM0, WX485, WX487, WX489, WX491, WX493, WX495, WX497, WX499, WX501, WX503, WX505, WX507, WX509, WX511, WX513, WX515, WX517, WX519, WX521, WX523, WX525, WX527, WX529, WX531, WX533, WX535, WX537, WX539, WX541, WX543, WX545, WX547, WX645, WX647, WX649, WX651, WX653, WX655, WX657, WX659, WX661, WX663, WX665, WX667, WX669, WX671, WX673, WX675, WX677, WX679, WX681, WX683, WX685, WX687, WX689, WX691, WX693, WX695, WX697, WX699, WX701, WX703, WX705, WX707, WX709, WX711, WX713, WX715, WX717, WX719, WX721, WX723, WX725, WX727, WX729, WX731, WX733, WX735, WX737, WX739, WX741, WX743, WX745, WX747, WX749, WX751, WX753, WX755, WX757, WX759, WX761, WX763, WX765, WX767, WX769, WX771, WX773, WX775, WX777, WX779, WX781, WX783, WX785, WX787, WX789, WX791, WX793, WX795, WX797, WX799, WX801, WX803, WX805, WX807, WX809, WX811, WX813, WX815, WX817, WX819, WX821, WX823, WX825, WX827, WX829, WX831, WX833, WX835, WX837, WX839, WX841, WX843, WX845, WX847, WX849, WX851, WX853, WX855, WX857, WX859, WX861, WX863, WX865, WX867, WX869, WX871, WX873, WX875, WX877, WX879, WX881, WX883, WX885, WX887, WX889, WX891, WX893, WX895, WX897, WX899, WX1778, WX1780, WX1782, WX1784, WX1786, WX1788, WX1790, WX1792, WX1794, WX1796, WX1798, WX1800, WX1802, WX1804, WX1806, WX1808, WX1810, WX1812, WX1814, WX1816, WX1818, WX1820, WX1822, WX1824, WX1826, WX1828, WX1830, WX1832, WX1834, WX1836, WX1838, WX1840, WX1938, WX1940, WX1942, WX1944, WX1946, WX1948, WX1950, WX1952, WX1954, WX1956, WX1958, WX1960, WX1962, WX1964, WX1966, WX1968, WX1970, WX1972, WX1974, WX1976, WX1978, WX1980, WX1982, WX1984, WX1986, WX1988, WX1990, WX1992, WX1994, WX1996, WX1998, WX2000, WX2002, WX2004, WX2006, WX2008, WX2010, WX2012, WX2014, WX2016, WX2018, WX2020, WX2022, WX2024, WX2026, WX2028, WX2030, WX2032, WX2034, WX2036, WX2038, WX2040, WX2042, WX2044, WX2046, WX2048, WX2050, WX2052, WX2054, WX2056, WX2058, WX2060, WX2062, WX2064, WX2066, WX2068, WX2070, WX2072, WX2074, WX2076, WX2078, WX2080, WX2082, WX2084, WX2086, WX2088, WX2090, WX2092, WX2094, WX2096, WX2098, WX2100, WX2102, WX2104, WX2106, WX2108, WX2110, WX2112, WX2114, WX2116, WX2118, WX2120, WX2122, WX2124, WX2126, WX2128, WX2130, WX2132, WX2134, WX2136, WX2138, WX2140, WX2142, WX2144, WX2146, WX2148, WX2150, WX2152, WX2154, WX2156, WX2158, WX2160, WX2162, WX2164, WX2166, WX2168, WX2170, WX2172, WX2174, WX2176, WX2178, WX2180, WX2182, WX2184, WX2186, WX2188, WX2190, WX2192, WX3071, WX3073, WX3075, WX3077, WX3079, WX3081, WX3083, WX3085, WX3087, WX3089, WX3091, WX3093, WX3095, WX3097, WX3099, WX3101, WX3103, WX3105, WX3107, WX3109, WX3111, WX3113, WX3115, WX3117, WX3119, WX3121, WX3123, WX3125, WX3127, WX3129, WX3131, WX3133, WX3231, WX3233, WX3235, WX3237, WX3239, WX3241, WX3243, WX3245, WX3247, WX3249, WX3251, WX3253, WX3255, WX3257, WX3259, WX3261, WX3263, WX3265, WX3267, WX3269, WX3271, WX3273, WX3275, WX3277, WX3279, WX3281, WX3283, WX3285, WX3287, WX3289, WX3291, WX3293, WX3295, WX3297, WX3299, WX3301, WX3303, WX3305, WX3307, WX3309, WX3311, WX3313, WX3315, WX3317, WX3319, WX3321, WX3323, WX3325, WX3327, WX3329, WX3331, WX3333, WX3335, WX3337, WX3339, WX3341, WX3343, WX3345, WX3347, WX3349, WX3351, WX3353, WX3355, WX3357, WX3359, WX3361, WX3363, WX3365, WX3367, WX3369, WX3371, WX3373, WX3375, WX3377, WX3379, WX3381, WX3383, WX3385, WX3387, WX3389, WX3391, WX3393, WX3395, WX3397, WX3399, WX3401, WX3403, WX3405, WX3407, WX3409, WX3411, WX3413, WX3415, WX3417, WX3419, WX3421, WX3423, WX3425, WX3427, WX3429, WX3431, WX3433, WX3435, WX3437, WX3439, WX3441, WX3443, WX3445, WX3447, WX3449, WX3451, WX3453, WX3455, WX3457, WX3459, WX3461, WX3463, WX3465, WX3467, WX3469, WX3471, WX3473, WX3475, WX3477, WX3479, WX3481, WX3483, WX3485, WX4364, WX4366, WX4368, WX4370, WX4372, WX4374, WX4376, WX4378, WX4380, WX4382, WX4384, WX4386, WX4388, WX4390, WX4392, WX4394, WX4396, WX4398, WX4400, WX4402, WX4404, WX4406, WX4408, WX4410, WX4412, WX4414, WX4416, WX4418, WX4420, WX4422, WX4424, WX4426, WX4524, WX4526, WX4528, WX4530, WX4532, WX4534, WX4536, WX4538, WX4540, WX4542, WX4544, WX4546, WX4548, WX4550, WX4552, WX4554, WX4556, WX4558, WX4560, WX4562, WX4564, WX4566, WX4568, WX4570, WX4572, WX4574, WX4576, WX4578, WX4580, WX4582, WX4584, WX4586, WX4588, WX4590, WX4592, WX4594, WX4596, WX4598, WX4600, WX4602, WX4604, WX4606, WX4608, WX4610, WX4612, WX4614, WX4616, WX4618, WX4620, WX4622, WX4624, WX4626, WX4628, WX4630, WX4632, WX4634, WX4636, WX4638, WX4640, WX4642, WX4644, WX4646, WX4648, WX4650, WX4652, WX4654, WX4656, WX4658, WX4660, WX4662, WX4664, WX4666, WX4668, WX4670, WX4672, WX4674, WX4676, WX4678, WX4680, WX4682, WX4684, WX4686, WX4688, WX4690, WX4692, WX4694, WX4696, WX4698, WX4700, WX4702, WX4704, WX4706, WX4708, WX4710, WX4712, WX4714, WX4716, WX4718, WX4720, WX4722, WX4724, WX4726, WX4728, WX4730, WX4732, WX4734, WX4736, WX4738, WX4740, WX4742, WX4744, WX4746, WX4748, WX4750, WX4752, WX4754, WX4756, WX4758, WX4760, WX4762, WX4764, WX4766, WX4768, WX4770, WX4772, WX4774, WX4776, WX4778, WX5657, WX5659, WX5661, WX5663, WX5665, WX5667, WX5669, WX5671, WX5673, WX5675, WX5677, WX5679, WX5681, WX5683, WX5685, WX5687, WX5689, WX5691, WX5693, WX5695, WX5697, WX5699, WX5701, WX5703, WX5705, WX5707, WX5709, WX5711, WX5713, WX5715, WX5717, WX5719, WX5817, WX5819, WX5821, WX5823, WX5825, WX5827, WX5829, WX5831, WX5833, WX5835, WX5837, WX5839, WX5841, WX5843, WX5845, WX5847, WX5849, WX5851, WX5853, WX5855, WX5857, WX5859, WX5861, WX5863, WX5865, WX5867, WX5869, WX5871, WX5873, WX5875, WX5877, WX5879, WX5881, WX5883, WX5885, WX5887, WX5889, WX5891, WX5893, WX5895, WX5897, WX5899, WX5901, WX5903, WX5905, WX5907, WX5909, WX5911, WX5913, WX5915, WX5917, WX5919, WX5921, WX5923, WX5925, WX5927, WX5929, WX5931, WX5933, WX5935, WX5937, WX5939, WX5941, WX5943, WX5945, WX5947, WX5949, WX5951, WX5953, WX5955, WX5957, WX5959, WX5961, WX5963, WX5965, WX5967, WX5969, WX5971, WX5973, WX5975, WX5977, WX5979, WX5981, WX5983, WX5985, WX5987, WX5989, WX5991, WX5993, WX5995, WX5997, WX5999, WX6001, WX6003, WX6005, WX6007, WX6009, WX6011, WX6013, WX6015, WX6017, WX6019, WX6021, WX6023, WX6025, WX6027, WX6029, WX6031, WX6033, WX6035, WX6037, WX6039, WX6041, WX6043, WX6045, WX6047, WX6049, WX6051, WX6053, WX6055, WX6057, WX6059, WX6061, WX6063, WX6065, WX6067, WX6069, WX6071, WX6950, WX6952, WX6954, WX6956, WX6958, WX6960, WX6962, WX6964, WX6966, WX6968, WX6970, WX6972, WX6974, WX6976, WX6978, WX6980, WX6982, WX6984, WX6986, WX6988, WX6990, WX6992, WX6994, WX6996, WX6998, WX7000, WX7002, WX7004, WX7006, WX7008, WX7010, WX7012, WX7110, WX7112, WX7114, WX7116, WX7118, WX7120, WX7122, WX7124, WX7126, WX7128, WX7130, WX7132, WX7134, WX7136, WX7138, WX7140, WX7142, WX7144, WX7146, WX7148, WX7150, WX7152, WX7154, WX7156, WX7158, WX7160, WX7162, WX7164, WX7166, WX7168, WX7170, WX7172, WX7174, WX7176, WX7178, WX7180, WX7182, WX7184, WX7186, WX7188, WX7190, WX7192, WX7194, WX7196, WX7198, WX7200, WX7202, WX7204, WX7206, WX7208, WX7210, WX7212, WX7214, WX7216, WX7218, WX7220, WX7222, WX7224, WX7226, WX7228, WX7230, WX7232, WX7234, WX7236, WX7238, WX7240, WX7242, WX7244, WX7246, WX7248, WX7250, WX7252, WX7254, WX7256, WX7258, WX7260, WX7262, WX7264, WX7266, WX7268, WX7270, WX7272, WX7274, WX7276, WX7278, WX7280, WX7282, WX7284, WX7286, WX7288, WX7290, WX7292, WX7294, WX7296, WX7298, WX7300, WX7302, WX7304, WX7306, WX7308, WX7310, WX7312, WX7314, WX7316, WX7318, WX7320, WX7322, WX7324, WX7326, WX7328, WX7330, WX7332, WX7334, WX7336, WX7338, WX7340, WX7342, WX7344, WX7346, WX7348, WX7350, WX7352, WX7354, WX7356, WX7358, WX7360, WX7362, WX7364, WX8243, WX8245, WX8247, WX8249, WX8251, WX8253, WX8255, WX8257, WX8259, WX8261, WX8263, WX8265, WX8267, WX8269, WX8271, WX8273, WX8275, WX8277, WX8279, WX8281, WX8283, WX8285, WX8287, WX8289, WX8291, WX8293, WX8295, WX8297, WX8299, WX8301, WX8303, WX8305, WX8403, WX8405, WX8407, WX8409, WX8411, WX8413, WX8415, WX8417, WX8419, WX8421, WX8423, WX8425, WX8427, WX8429, WX8431, WX8433, WX8435, WX8437, WX8439, WX8441, WX8443, WX8445, WX8447, WX8449, WX8451, WX8453, WX8455, WX8457, WX8459, WX8461, WX8463, WX8465, WX8467, WX8469, WX8471, WX8473, WX8475, WX8477, WX8479, WX8481, WX8483, WX8485, WX8487, WX8489, WX8491, WX8493, WX8495, WX8497, WX8499, WX8501, WX8503, WX8505, WX8507, WX8509, WX8511, WX8513, WX8515, WX8517, WX8519, WX8521, WX8523, WX8525, WX8527, WX8529, WX8531, WX8533, WX8535, WX8537, WX8539, WX8541, WX8543, WX8545, WX8547, WX8549, WX8551, WX8553, WX8555, WX8557, WX8559, WX8561, WX8563, WX8565, WX8567, WX8569, WX8571, WX8573, WX8575, WX8577, WX8579, WX8581, WX8583, WX8585, WX8587, WX8589, WX8591, WX8593, WX8595, WX8597, WX8599, WX8601, WX8603, WX8605, WX8607, WX8609, WX8611, WX8613, WX8615, WX8617, WX8619, WX8621, WX8623, WX8625, WX8627, WX8629, WX8631, WX8633, WX8635, WX8637, WX8639, WX8641, WX8643, WX8645, WX8647, WX8649, WX8651, WX8653, WX8655, WX8657, WX9536, WX9538, WX9540, WX9542, WX9544, WX9546, WX9548, WX9550, WX9552, WX9554, WX9556, WX9558, WX9560, WX9562, WX9564, WX9566, WX9568, WX9570, WX9572, WX9574, WX9576, WX9578, WX9580, WX9582, WX9584, WX9586, WX9588, WX9590, WX9592, WX9594, WX9596, WX9598, WX9696, WX9698, WX9700, WX9702, WX9704, WX9706, WX9708, WX9710, WX9712, WX9714, WX9716, WX9718, WX9720, WX9722, WX9724, WX9726, WX9728, WX9730, WX9732, WX9734, WX9736, WX9738, WX9740, WX9742, WX9744, WX9746, WX9748, WX9750, WX9752, WX9754, WX9756, WX9758, WX9760, WX9762, WX9764, WX9766, WX9768, WX9770, WX9772, WX9774, WX9776, WX9778, WX9780, WX9782, WX9784, WX9786, WX9788, WX9790, WX9792, WX9794, WX9796, WX9798, WX9800, WX9802, WX9804, WX9806, WX9808, WX9810, WX9812, WX9814, WX9816, WX9818, WX9820, WX9822, WX9824, WX9826, WX9828, WX9830, WX9832, WX9834, WX9836, WX9838, WX9840, WX9842, WX9844, WX9846, WX9848, WX9850, WX9852, WX9854, WX9856, WX9858, WX9860, WX9862, WX9864, WX9866, WX9868, WX9870, WX9872, WX9874, WX9876, WX9878, WX9880, WX9882, WX9884, WX9886, WX9888, WX9890, WX9892, WX9894, WX9896, WX9898, WX9900, WX9902, WX9904, WX9906, WX9908, WX9910, WX9912, WX9914, WX9916, WX9918, WX9920, WX9922, WX9924, WX9926, WX9928, WX9930, WX9932, WX9934, WX9936, WX9938, WX9940, WX9942, WX9944, WX9946, WX9948, WX9950, WX10829, WX10831, WX10833, WX10835, WX10837, WX10839, WX10841, WX10843, WX10845, WX10847, WX10849, WX10851, WX10853, WX10855, WX10857, WX10859, WX10861, WX10863, WX10865, WX10867, WX10869, WX10871, WX10873, WX10875, WX10877, WX10879, WX10881, WX10883, WX10885, WX10887, WX10889, WX10891, WX10989, WX10991, WX10993, WX10995, WX10997, WX10999, WX11001, WX11003, WX11005, WX11007, WX11009, WX11011, WX11013, WX11015, WX11017, WX11019, WX11021, WX11023, WX11025, WX11027, WX11029, WX11031, WX11033, WX11035, WX11037, WX11039, WX11041, WX11043, WX11045, WX11047, WX11049, WX11051, WX11053, WX11055, WX11057, WX11059, WX11061, WX11063, WX11065, WX11067, WX11069, WX11071, WX11073, WX11075, WX11077, WX11079, WX11081, WX11083, WX11085, WX11087, WX11089, WX11091, WX11093, WX11095, WX11097, WX11099, WX11101, WX11103, WX11105, WX11107, WX11109, WX11111, WX11113, WX11115, WX11117, WX11119, WX11121, WX11123, WX11125, WX11127, WX11129, WX11131, WX11133, WX11135, WX11137, WX11139, WX11141, WX11143, WX11145, WX11147, WX11149, WX11151, WX11153, WX11155, WX11157, WX11159, WX11161, WX11163, WX11165, WX11167, WX11169, WX11171, WX11173, WX11175, WX11177, WX11179, WX11181, WX11183, WX11185, WX11187, WX11189, WX11191, WX11193, WX11195, WX11197, WX11199, WX11201, WX11203, WX11205, WX11207, WX11209, WX11211, WX11213, WX11215, WX11217, WX11219, WX11221, WX11223, WX11225, WX11227, WX11229, WX11231, WX11233, WX11235, WX11237, WX11239, WX11241, WX11243;
output DATA_9_1, DATA_9_2, DATA_9_3, DATA_9_31, DATA_9_30, DATA_9_29, DATA_9_28, DATA_9_27, DATA_9_26, DATA_9_25, DATA_9_24, DATA_9_23, DATA_9_22, DATA_9_21, DATA_9_20, DATA_9_19, DATA_9_18, DATA_9_17, DATA_9_16, DATA_9_15, DATA_9_14, DATA_9_13, DATA_9_12, DATA_9_11, DATA_9_10, DATA_9_9, DATA_9_8, DATA_9_7, DATA_9_6, DATA_9_5, DATA_9_4, DATA_9_0, CRC_OUT_9_0, CRC_OUT_9_1, CRC_OUT_9_2, CRC_OUT_9_3, CRC_OUT_9_4, CRC_OUT_9_5, CRC_OUT_9_6, CRC_OUT_9_7, CRC_OUT_9_8, CRC_OUT_9_9, CRC_OUT_9_10, CRC_OUT_9_11, CRC_OUT_9_12, CRC_OUT_9_13, CRC_OUT_9_14, CRC_OUT_9_15, CRC_OUT_9_16, CRC_OUT_9_17, CRC_OUT_9_18, CRC_OUT_9_19, CRC_OUT_9_20, CRC_OUT_9_21, CRC_OUT_9_22, CRC_OUT_9_23, CRC_OUT_9_24, CRC_OUT_9_25, CRC_OUT_9_26, CRC_OUT_9_27, CRC_OUT_9_28, CRC_OUT_9_29, CRC_OUT_9_30, CRC_OUT_9_31, CRC_OUT_8_0, CRC_OUT_8_1, CRC_OUT_8_2, CRC_OUT_8_3, CRC_OUT_8_4, CRC_OUT_8_5, CRC_OUT_8_6, CRC_OUT_8_7, CRC_OUT_8_8, CRC_OUT_8_9, CRC_OUT_8_10, CRC_OUT_8_11, CRC_OUT_8_12, CRC_OUT_8_13, CRC_OUT_8_14, CRC_OUT_8_15, CRC_OUT_8_16, CRC_OUT_8_17, CRC_OUT_8_18, CRC_OUT_8_19, CRC_OUT_8_20, CRC_OUT_8_21, CRC_OUT_8_22, CRC_OUT_8_23, CRC_OUT_8_24, CRC_OUT_8_25, CRC_OUT_8_26, CRC_OUT_8_27, CRC_OUT_8_28, CRC_OUT_8_29, CRC_OUT_8_30, CRC_OUT_8_31, CRC_OUT_7_0, CRC_OUT_7_1, CRC_OUT_7_2, CRC_OUT_7_3, CRC_OUT_7_4, CRC_OUT_7_5, CRC_OUT_7_6, CRC_OUT_7_7, CRC_OUT_7_8, CRC_OUT_7_9, CRC_OUT_7_10, CRC_OUT_7_11, CRC_OUT_7_12, CRC_OUT_7_13, CRC_OUT_7_14, CRC_OUT_7_15, CRC_OUT_7_16, CRC_OUT_7_17, CRC_OUT_7_18, CRC_OUT_7_19, CRC_OUT_7_20, CRC_OUT_7_21, CRC_OUT_7_22, CRC_OUT_7_23, CRC_OUT_7_24, CRC_OUT_7_25, CRC_OUT_7_26, CRC_OUT_7_27, CRC_OUT_7_28, CRC_OUT_7_29, CRC_OUT_7_30, CRC_OUT_7_31, CRC_OUT_6_0, CRC_OUT_6_1, CRC_OUT_6_2, CRC_OUT_6_3, CRC_OUT_6_4, CRC_OUT_6_5, CRC_OUT_6_6, CRC_OUT_6_7, CRC_OUT_6_8, CRC_OUT_6_9, CRC_OUT_6_10, CRC_OUT_6_11, CRC_OUT_6_12, CRC_OUT_6_13, CRC_OUT_6_14, CRC_OUT_6_15, CRC_OUT_6_16, CRC_OUT_6_17, CRC_OUT_6_18, CRC_OUT_6_19, CRC_OUT_6_20, CRC_OUT_6_21, CRC_OUT_6_22, CRC_OUT_6_23, CRC_OUT_6_24, CRC_OUT_6_25, CRC_OUT_6_26, CRC_OUT_6_27, CRC_OUT_6_28, CRC_OUT_6_29, CRC_OUT_6_30, CRC_OUT_6_31, CRC_OUT_5_0, CRC_OUT_5_1, CRC_OUT_5_2, CRC_OUT_5_3, CRC_OUT_5_4, CRC_OUT_5_5, CRC_OUT_5_6, CRC_OUT_5_7, CRC_OUT_5_8, CRC_OUT_5_9, CRC_OUT_5_10, CRC_OUT_5_11, CRC_OUT_5_12, CRC_OUT_5_13, CRC_OUT_5_14, CRC_OUT_5_15, CRC_OUT_5_16, CRC_OUT_5_17, CRC_OUT_5_18, CRC_OUT_5_19, CRC_OUT_5_20, CRC_OUT_5_21, CRC_OUT_5_22, CRC_OUT_5_23, CRC_OUT_5_24, CRC_OUT_5_25, CRC_OUT_5_26, CRC_OUT_5_27, CRC_OUT_5_28, CRC_OUT_5_29, CRC_OUT_5_30, CRC_OUT_5_31, CRC_OUT_4_0, CRC_OUT_4_1, CRC_OUT_4_2, CRC_OUT_4_3, CRC_OUT_4_4, CRC_OUT_4_5, CRC_OUT_4_6, CRC_OUT_4_7, CRC_OUT_4_8, CRC_OUT_4_9, CRC_OUT_4_10, CRC_OUT_4_11, CRC_OUT_4_12, CRC_OUT_4_13, CRC_OUT_4_14, CRC_OUT_4_15, CRC_OUT_4_16, CRC_OUT_4_17, CRC_OUT_4_18, CRC_OUT_4_19, CRC_OUT_4_20, CRC_OUT_4_21, CRC_OUT_4_22, CRC_OUT_4_23, CRC_OUT_4_24, CRC_OUT_4_25, CRC_OUT_4_26, CRC_OUT_4_27, CRC_OUT_4_28, CRC_OUT_4_29, CRC_OUT_4_30, CRC_OUT_4_31, CRC_OUT_3_0, CRC_OUT_3_1, CRC_OUT_3_2, CRC_OUT_3_3, CRC_OUT_3_4, CRC_OUT_3_5, CRC_OUT_3_6, CRC_OUT_3_7, CRC_OUT_3_8, CRC_OUT_3_9, CRC_OUT_3_10, CRC_OUT_3_11, CRC_OUT_3_12, CRC_OUT_3_13, CRC_OUT_3_14, CRC_OUT_3_15, CRC_OUT_3_16, CRC_OUT_3_17, CRC_OUT_3_18, CRC_OUT_3_19, CRC_OUT_3_20, CRC_OUT_3_21, CRC_OUT_3_22, CRC_OUT_3_23, CRC_OUT_3_24, CRC_OUT_3_25, CRC_OUT_3_26, CRC_OUT_3_27, CRC_OUT_3_28, CRC_OUT_3_29, CRC_OUT_3_30, CRC_OUT_3_31, CRC_OUT_2_0, CRC_OUT_2_1, CRC_OUT_2_2, CRC_OUT_2_3, CRC_OUT_2_4, CRC_OUT_2_5, CRC_OUT_2_6, CRC_OUT_2_7, CRC_OUT_2_8, CRC_OUT_2_9, CRC_OUT_2_10, CRC_OUT_2_11, CRC_OUT_2_12, CRC_OUT_2_13, CRC_OUT_2_14, CRC_OUT_2_15, CRC_OUT_2_16, CRC_OUT_2_17, CRC_OUT_2_18, CRC_OUT_2_19, CRC_OUT_2_20, CRC_OUT_2_21, CRC_OUT_2_22, CRC_OUT_2_23, CRC_OUT_2_24, CRC_OUT_2_25, CRC_OUT_2_26, CRC_OUT_2_27, CRC_OUT_2_28, CRC_OUT_2_29, CRC_OUT_2_30, CRC_OUT_2_31, CRC_OUT_1_0, CRC_OUT_1_1, CRC_OUT_1_2, CRC_OUT_1_3, CRC_OUT_1_4, CRC_OUT_1_5, CRC_OUT_1_6, CRC_OUT_1_7, CRC_OUT_1_8, CRC_OUT_1_9, CRC_OUT_1_10, CRC_OUT_1_11, CRC_OUT_1_12, CRC_OUT_1_13, CRC_OUT_1_14, CRC_OUT_1_15, CRC_OUT_1_16, CRC_OUT_1_17, CRC_OUT_1_18, CRC_OUT_1_19, CRC_OUT_1_20, CRC_OUT_1_21, CRC_OUT_1_22, CRC_OUT_1_23, CRC_OUT_1_24, CRC_OUT_1_25, CRC_OUT_1_26, CRC_OUT_1_27, CRC_OUT_1_28, CRC_OUT_1_29, CRC_OUT_1_30, CRC_OUT_1_31, n711, n716, n721, n726, n731, n736, n741, n746, n751, n756, n761, n766, n771, n776, n781, n786, n791, n796, n801, n806, n811, n816, n821, n826, n831, n836, n841, n846, n851, n856, n861, n866, n871, n876, n881, n886, n891, n896, n901, n906, n911, n916, n921, n926, n931, n936, n941, n946, n951, n956, n961, n966, n971, n976, n981, n986, n991, n996, n1001, n1006, n1011, n1016, n1021, n1026, n1031, n1036, n1041, n1046, n1051, n1056, n1061, n1066, n1071, n1076, n1081, n1086, n1091, n1096, n1101, n1106, n1111, n1116, n1121, n1126, n1131, n1136, n1141, n1146, n1151, n1156, n1161, n1166, n1171, n1176, n1181, n1186, n1191, n1196, n1201, n1206, n1211, n1216, n1221, n1226, n1231, n1236, n1241, n1246, n1251, n1256, n1261, n1266, n1271, n1276, n1281, n1286, n1291, n1296, n1301, n1306, n1311, n1316, n1321, n1326, n1331, n1336, n1341, n1346, n1351, n1356, n1361, n1366, n1371, n1376, n1381, n1386, n1391, n1396, n1401, n1406, n1411, n1416, n1421, n1426, n1431, n1436, n1441, n1446, n1451, n1456, n1461, n1466, n1471, n1476, n1481, n1486, n1491, n1496, n1501, n1506, n1639, n1644, n1649, n1654, n1659, n1664, n1669, n1674, n1679, n1684, n1689, n1694, n1699, n1704, n1709, n1714, n1719, n1724, n1729, n1734, n1739, n1744, n1749, n1754, n1759, n1764, n1769, n1774, n1779, n1784, n1789, n1794, n1799, n1804, n1809, n1814, n1819, n1824, n1829, n1834, n1839, n1844, n1849, n1854, n1859, n1864, n1869, n1874, n1879, n1884, n1889, n1894, n1899, n1904, n1909, n1914, n1919, n1924, n1929, n1934, n1939, n1944, n1949, n1954, n1959, n1964, n1969, n1974, n1979, n1984, n1989, n1994, n1999, n2004, n2009, n2014, n2019, n2024, n2029, n2034, n2039, n2044, n2049, n2054, n2059, n2064, n2069, n2074, n2079, n2084, n2089, n2094, n2099, n2104, n2109, n2114, n2119, n2124, n2129, n2134, n2139, n2144, n2149, n2154, n2159, n2164, n2169, n2174, n2179, n2184, n2189, n2194, n2199, n2204, n2209, n2214, n2219, n2224, n2229, n2234, n2239, n2244, n2249, n2254, n2259, n2264, n2269, n2274, n2279, n2284, n2289, n2294, n2299, n2304, n2309, n2314, n2319, n2324, n2329, n2334, n2339, n2344, n2349, n2354, n2359, n2364, n2369, n2374, n2379, n2384, n2389, n2394, n2399, n2404, n2409, n2414, n2419, n2424, n2429, n2434, n2567, n2572, n2577, n2582, n2587, n2592, n2597, n2602, n2607, n2612, n2617, n2622, n2627, n2632, n2637, n2642, n2647, n2652, n2657, n2662, n2667, n2672, n2677, n2682, n2687, n2692, n2697, n2702, n2707, n2712, n2717, n2722, n2727, n2732, n2737, n2742, n2747, n2752, n2757, n2762, n2767, n2772, n2777, n2782, n2787, n2792, n2797, n2802, n2807, n2812, n2817, n2822, n2827, n2832, n2837, n2842, n2847, n2852, n2857, n2862, n2867, n2872, n2877, n2882, n2887, n2892, n2897, n2902, n2907, n2912, n2917, n2922, n2927, n2932, n2937, n2942, n2947, n2952, n2957, n2962, n2967, n2972, n2977, n2982, n2987, n2992, n2997, n3002, n3007, n3012, n3017, n3022, n3027, n3032, n3037, n3042, n3047, n3052, n3057, n3062, n3067, n3072, n3077, n3082, n3087, n3092, n3097, n3102, n3107, n3112, n3117, n3122, n3127, n3132, n3137, n3142, n3147, n3152, n3157, n3162, n3167, n3172, n3177, n3182, n3187, n3192, n3197, n3202, n3207, n3212, n3217, n3222, n3227, n3232, n3237, n3242, n3247, n3252, n3257, n3262, n3267, n3272, n3277, n3282, n3287, n3292, n3297, n3302, n3307, n3312, n3317, n3322, n3327, n3332, n3337, n3342, n3347, n3352, n3357, n3362, n3495, n3500, n3505, n3510, n3515, n3520, n3525, n3530, n3535, n3540, n3545, n3550, n3555, n3560, n3565, n3570, n3575, n3580, n3585, n3590, n3595, n3600, n3605, n3610, n3615, n3620, n3625, n3630, n3635, n3640, n3645, n3650, n3655, n3660, n3665, n3670, n3675, n3680, n3685, n3690, n3695, n3700, n3705, n3710, n3715, n3720, n3725, n3730, n3735, n3740, n3745, n3750, n3755, n3760, n3765, n3770, n3775, n3780, n3785, n3790, n3795, n3800, n3805, n3810, n3815, n3820, n3825, n3830, n3835, n3840, n3845, n3850, n3855, n3860, n3865, n3870, n3875, n3880, n3885, n3890, n3895, n3900, n3905, n3910, n3915, n3920, n3925, n3930, n3935, n3940, n3945, n3950, n3955, n3960, n3965, n3970, n3975, n3980, n3985, n3990, n3995, n4000, n4005, n4010, n4015, n4020, n4025, n4030, n4035, n4040, n4045, n4050, n4055, n4060, n4065, n4070, n4075, n4080, n4085, n4090, n4095, n4100, n4105, n4110, n4115, n4120, n4125, n4130, n4135, n4140, n4145, n4150, n4155, n4160, n4165, n4170, n4175, n4180, n4185, n4190, n4195, n4200, n4205, n4210, n4215, n4220, n4225, n4230, n4235, n4240, n4245, n4250, n4255, n4260, n4265, n4270, n4275, n4280, n4285, n4290, n4423, n4428, n4433, n4438, n4443, n4448, n4453, n4458, n4463, n4468, n4473, n4478, n4483, n4488, n4493, n4498, n4503, n4508, n4513, n4518, n4523, n4528, n4533, n4538, n4543, n4548, n4553, n4558, n4563, n4568, n4573, n4578, n4583, n4588, n4593, n4598, n4603, n4608, n4613, n4618, n4623, n4628, n4633, n4638, n4643, n4648, n4653, n4658, n4663, n4668, n4673, n4678, n4683, n4688, n4693, n4698, n4703, n4708, n4713, n4718, n4723, n4728, n4733, n4738, n4743, n4748, n4753, n4758, n4763, n4768, n4773, n4778, n4783, n4788, n4793, n4798, n4803, n4808, n4813, n4818, n4823, n4828, n4833, n4838, n4843, n4848, n4853, n4858, n4863, n4868, n4873, n4878, n4883, n4888, n4893, n4898, n4903, n4908, n4913, n4918, n4923, n4928, n4933, n4938, n4943, n4948, n4953, n4958, n4963, n4968, n4973, n4978, n4983, n4988, n4993, n4998, n5003, n5008, n5013, n5018, n5023, n5028, n5033, n5038, n5043, n5048, n5053, n5058, n5063, n5068, n5073, n5078, n5083, n5088, n5093, n5098, n5103, n5108, n5113, n5118, n5123, n5128, n5133, n5138, n5143, n5148, n5153, n5158, n5163, n5168, n5173, n5178, n5183, n5188, n5193, n5198, n5203, n5208, n5213, n5218, n5351, n5356, n5361, n5366, n5371, n5376, n5381, n5386, n5391, n5396, n5401, n5406, n5411, n5416, n5421, n5426, n5431, n5436, n5441, n5446, n5451, n5456, n5461, n5466, n5471, n5476, n5481, n5486, n5491, n5496, n5501, n5506, n5511, n5516, n5521, n5526, n5531, n5536, n5541, n5546, n5551, n5556, n5561, n5566, n5571, n5576, n5581, n5586, n5591, n5596, n5601, n5606, n5611, n5616, n5621, n5626, n5631, n5636, n5641, n5646, n5651, n5656, n5661, n5666, n5671, n5676, n5681, n5686, n5691, n5696, n5701, n5706, n5711, n5716, n5721, n5726, n5731, n5736, n5741, n5746, n5751, n5756, n5761, n5766, n5771, n5776, n5781, n5786, n5791, n5796, n5801, n5806, n5811, n5816, n5821, n5826, n5831, n5836, n5841, n5846, n5851, n5856, n5861, n5866, n5871, n5876, n5881, n5886, n5891, n5896, n5901, n5906, n5911, n5916, n5921, n5926, n5931, n5936, n5941, n5946, n5951, n5956, n5961, n5966, n5971, n5976, n5981, n5986, n5991, n5996, n6001, n6006, n6011, n6016, n6021, n6026, n6031, n6036, n6041, n6046, n6051, n6056, n6061, n6066, n6071, n6076, n6081, n6086, n6091, n6096, n6101, n6106, n6111, n6116, n6121, n6126, n6131, n6136, n6141, n6146, n6279, n6284, n6289, n6294, n6299, n6304, n6309, n6314, n6319, n6324, n6329, n6334, n6339, n6344, n6349, n6354, n6359, n6364, n6369, n6374, n6379, n6384, n6389, n6394, n6399, n6404, n6409, n6414, n6419, n6424, n6429, n6434, n6439, n6444, n6449, n6454, n6459, n6464, n6469, n6474, n6479, n6484, n6489, n6494, n6499, n6504, n6509, n6514, n6519, n6524, n6529, n6534, n6539, n6544, n6549, n6554, n6559, n6564, n6569, n6574, n6579, n6584, n6589, n6594, n6599, n6604, n6609, n6614, n6619, n6624, n6629, n6634, n6639, n6644, n6649, n6654, n6659, n6664, n6669, n6674, n6679, n6684, n6689, n6694, n6699, n6704, n6709, n6714, n6719, n6724, n6729, n6734, n6739, n6744, n6749, n6754, n6759, n6764, n6769, n6774, n6779, n6784, n6789, n6794, n6799, n6804, n6809, n6814, n6819, n6824, n6829, n6834, n6839, n6844, n6849, n6854, n6859, n6864, n6869, n6874, n6879, n6884, n6889, n6894, n6899, n6904, n6909, n6914, n6919, n6924, n6929, n6934, n6939, n6944, n6949, n6954, n6959, n6964, n6969, n6974, n6979, n6984, n6989, n6994, n6999, n7004, n7009, n7014, n7019, n7024, n7029, n7034, n7039, n7044, n7049, n7054, n7059, n7064, n7069, n7074, n7207, n7212, n7217, n7222, n7227, n7232, n7237, n7242, n7247, n7252, n7257, n7262, n7267, n7272, n7277, n7282, n7287, n7292, n7297, n7302, n7307, n7312, n7317, n7322, n7327, n7332, n7337, n7342, n7347, n7352, n7357, n7362, n7367, n7372, n7377, n7382, n7387, n7392, n7397, n7402, n7407, n7412, n7417, n7422, n7427, n7432, n7437, n7442, n7447, n7452, n7457, n7462, n7467, n7472, n7477, n7482, n7487, n7492, n7497, n7502, n7507, n7512, n7517, n7522, n7527, n7532, n7537, n7542, n7547, n7552, n7557, n7562, n7567, n7572, n7577, n7582, n7587, n7592, n7597, n7602, n7607, n7612, n7617, n7622, n7627, n7632, n7637, n7642, n7647, n7652, n7657, n7662, n7667, n7672, n7677, n7682, n7687, n7692, n7697, n7702, n7707, n7712, n7717, n7722, n7727, n7732, n7737, n7742, n7747, n7752, n7757, n7762, n7767, n7772, n7777, n7782, n7787, n7792, n7797, n7802, n7807, n7812, n7817, n7822, n7827, n7832, n7837, n7842, n7847, n7852, n7857, n7862, n7867, n7872, n7877, n7882, n7887, n7892, n7897, n7902, n7907, n7912, n7917, n7922, n7927, n7932, n7937, n7942, n7947, n7952, n7957, n7962, n7967, n7972, n7977, n7982, n7987, n7992, n7997, n8002, n8135, n8140, n8145, n8150, n8155, n8160, n8165, n8170, n8175, n8180, n8185, n8190, n8195, n8200, n8205, n8210, n8215, n8220, n8225, n8230, n8235, n8240, n8245, n8250, n8255, n8260, n8265, n8270, n8275, n8280, n8285, n8290, n8295, n8300, n8305, n8310, n8315, n8320, n8325, n8330, n8335, n8340, n8345, n8350, n8355, n8360, n8365, n8370, n8375, n8380, n8385, n8390, n8395, n8400, n8405, n8410, n8415, n8420, n8425, n8430, n8435, n8440, n8445, n8450, n8455, n8460, n8465, n8470, n8475, n8480, n8485, n8490, n8495, n8500, n8505, n8510, n8515, n8520, n8525, n8530, n8535, n8540, n8545, n8550, n8555, n8560, n8565, n8570, n8575, n8580, n8585, n8590, n8595, n8600, n8605, n8610, n8615, n8620, n8625, n8630, n8635, n8640, n8645, n8650, n8655, n8660, n8665, n8670, n8675, n8680, n8685, n8690, n8695, n8700, n8705, n8710, n8715, n8720, n8725, n8730, n8735, n8740, n8745, n8750, n8755, n8760, n8765, n8770, n8775, n8780, n8785, n8790, n8795, n8800, n8805, n8810, n8815, n8820, n8825, n8830, n8835, n8840, n8845, n8850, n8855, n8860, n8865, n8870, n8875, n8880, n8885, n8890, n8895, n8900, n8905, n8910, n8915, n8920, n8925, n8930;
wire n5539, n5540, n5541_1, n5542, n5543, n5544, n5545, n5546_1, n5548, n5549, n5550, n5551_1, n5552, n5553, n5554, n5556_1, n5557, n5558, n5559, n5560, n5561_1, n5562, n5564, n5565, n5566_1, n5567, n5568, n5569, n5570, n5572, n5573, n5574, n5575, n5576_1, n5577, n5578, n5580, n5581_1, n5582, n5583, n5584, n5585, n5586_1, n5588, n5589, n5590, n5591_1, n5592, n5593, n5594, n5596_1, n5597, n5598, n5599, n5600, n5601_1, n5602, n5604, n5605, n5606_1, n5607, n5608, n5609, n5610, n5612, n5613, n5614, n5615, n5616_1, n5617, n5618, n5620, n5621_1, n5622, n5623, n5624, n5625, n5626_1, n5628, n5629, n5630, n5631_1, n5632, n5633, n5634, n5636_1, n5637, n5638, n5639, n5640, n5641_1, n5642, n5644, n5645, n5646_1, n5647, n5648, n5649, n5650, n5652, n5653, n5654, n5655, n5656_1, n5657, n5658, n5660, n5661_1, n5662, n5663, n5664, n5665, n5666_1, n5668, n5669, n5670, n5671_1, n5672, n5673, n5674, n5676_1, n5677, n5678, n5679, n5680, n5681_1, n5682, n5684, n5685, n5686_1, n5687, n5688, n5689, n5690, n5692, n5693, n5694, n5695, n5696_1, n5697, n5698, n5700, n5701_1, n5702, n5703, n5704, n5705, n5706_1, n5708, n5709, n5710, n5711_1, n5712, n5713, n5714, n5716_1, n5717, n5718, n5719, n5720, n5721_1, n5722, n5724, n5725, n5726_1, n5727, n5728, n5729, n5730, n5732, n5733, n5734, n5735, n5736_1, n5737, n5738, n5740, n5741_1, n5742, n5743, n5744, n5745, n5746_1, n5748, n5749, n5750, n5751_1, n5752, n5753, n5754, n5756_1, n5757, n5758, n5759, n5760, n5761_1, n5762, n5764, n5765, n5766_1, n5767, n5768, n5769, n5770, n5772, n5773, n5774, n5775, n5776_1, n5777, n5778, n5780, n5781_1, n5782, n5783, n5784, n5785, n5786_1, n5788, n5789, n5790, n5791_1, n5792, n5793, n5794, n5827, n5829, n5830, n5831_1, n5832, n5833, n5834, n5836_1, n5837, n5838, n5839, n5841_1, n5842, n5843, n5844, n5845, n5846_1, n5848, n5849, n5850, n5851_1, n5853, n5854, n5855, n5856_1, n5857, n5858, n5860, n5861_1, n5862, n5863, n5865, n5866_1, n5867, n5868, n5869, n5870, n5872, n5873, n5874, n5875, n5877, n5878, n5879, n5880, n5881_1, n5882, n5884, n5885, n5886_1, n5887, n5889, n5890, n5891_1, n5892, n5893, n5894, n5896_1, n5897, n5898, n5899, n5901_1, n5902, n5903, n5904, n5905, n5906_1, n5908, n5909, n5910, n5911_1, n5913, n5914, n5915, n5916_1, n5917, n5918, n5920, n5921_1, n5922, n5923, n5925, n5926_1, n5927, n5928, n5929, n5930, n5932, n5933, n5934, n5935, n5937, n5938, n5939, n5940, n5941_1, n5942, n5944, n5945, n5946_1, n5947, n5949, n5950, n5951_1, n5952, n5953, n5954, n5956_1, n5957, n5958, n5959, n5961_1, n5962, n5963, n5964, n5965, n5966_1, n5968, n5969, n5970, n5971_1, n5973, n5974, n5975, n5976_1, n5977, n5978, n5980, n5981_1, n5982, n5983, n5985, n5986_1, n5987, n5988, n5989, n5990, n5992, n5993, n5994, n5995, n5997, n5998, n5999, n6000, n6001_1, n6002, n6004, n6005, n6006_1, n6007, n6009, n6010, n6011_1, n6012, n6013, n6014, n6016_1, n6017, n6018, n6019, n6021_1, n6022, n6023, n6024, n6025, n6026_1, n6028, n6029, n6030, n6031_1, n6033, n6034, n6035, n6036_1, n6037, n6038, n6040, n6041_1, n6042, n6043, n6045, n6046_1, n6047, n6048, n6049, n6050, n6052, n6053, n6054, n6055, n6057, n6058, n6059, n6060, n6061_1, n6062, n6064, n6065, n6066_1, n6067, n6069, n6070, n6071_1, n6072, n6073, n6074, n6076_1, n6077, n6078, n6079, n6081_1, n6082, n6083, n6084, n6085, n6086_1, n6088, n6089, n6090, n6091_1, n6093, n6094, n6095, n6096_1, n6097, n6098, n6100, n6101_1, n6102, n6103, n6105, n6106_1, n6107, n6108, n6109, n6110, n6112, n6113, n6114, n6115, n6117, n6118, n6119, n6120, n6121_1, n6122, n6124, n6125, n6126_1, n6127, n6129, n6130, n6131_1, n6132, n6133, n6134, n6136_1, n6137, n6138, n6139, n6141_1, n6142, n6143, n6144, n6145, n6146_1, n6148, n6149, n6150, n6151_1, n6153, n6154, n6155_1, n6156, n6157, n6158, n6160, n6161, n6162, n6163_1, n6165, n6166, n6167_1, n6168, n6169, n6170, n6172, n6173, n6174, n6175_1, n6177, n6178, n6179_1, n6180, n6181, n6182, n6184, n6185, n6186, n6187_1, n6189, n6190, n6191_1, n6192, n6193, n6194, n6196, n6197, n6198, n6199_1, n6201, n6202, n6203_1, n6204, n6205, n6206, n6208, n6209, n6210, n6211_1, n6309_1, n6311, n6313, n6315, n6317, n6318, n6320, n6322, n6324_1, n6326, n6328, n6330, n6332, n6333, n6335, n6337, n6339_1, n6341, n6343, n6344_1, n6346, n6348, n6350, n6352, n6354_1, n6356, n6358, n6360, n6362, n6364_1, n6366, n6368, n6370, n6372, n6374_1, n6408, n6409_1, n6410, n6411, n6412, n6413, n6415, n6416, n6417, n6418, n6420, n6421, n6422, n6423, n6424_1, n6425, n6427, n6428, n6429_1, n6430, n6432, n6433, n6434_1, n6435, n6436, n6437, n6439_1, n6440, n6441, n6442, n6444_1, n6445, n6446, n6447, n6448, n6449_1, n6451, n6452, n6453, n6454_1, n6456, n6457, n6458, n6459_1, n6460, n6461, n6463, n6464_1, n6465, n6466, n6468, n6469_1, n6470, n6471, n6472, n6473, n6475, n6476, n6477, n6478, n6480, n6481, n6482, n6483, n6484_1, n6485, n6487, n6488, n6489_1, n6490, n6492, n6493, n6494_1, n6495, n6496, n6497, n6499_1, n6500, n6501, n6502, n6504_1, n6505, n6506, n6507, n6508, n6509_1, n6511, n6512, n6513, n6514_1, n6516, n6517, n6518, n6519_1, n6520, n6521, n6523, n6524_1, n6525, n6526, n6528, n6529_1, n6530, n6531, n6532, n6533, n6535, n6536, n6537, n6538, n6540, n6541, n6542, n6543, n6544_1, n6545, n6547, n6548, n6549_1, n6550, n6552, n6553, n6554_1, n6555, n6556, n6557, n6559_1, n6560, n6561, n6562, n6564_1, n6565, n6566, n6567, n6568, n6569_1, n6571, n6572, n6573, n6574_1, n6576, n6577, n6578, n6579_1, n6580, n6581, n6583, n6584_1, n6585, n6586, n6588, n6589_1, n6590, n6591, n6592, n6593, n6595, n6596, n6597, n6598, n6600, n6601, n6602, n6603, n6604_1, n6605, n6607, n6608, n6609_1, n6610, n6612, n6613, n6614_1, n6615, n6616, n6617, n6619_1, n6620, n6621, n6622, n6624_1, n6625, n6626, n6627, n6628, n6629_1, n6631, n6632, n6633, n6634_1, n6636, n6637, n6638, n6639_1, n6640, n6641, n6643, n6644_1, n6645, n6646, n6648, n6649_1, n6650, n6651, n6652, n6653, n6655, n6656, n6657, n6658, n6660, n6661, n6662, n6663, n6664_1, n6665, n6667, n6668, n6669_1, n6670, n6672, n6673, n6674_1, n6675, n6676, n6677, n6679_1, n6680, n6681, n6682, n6684_1, n6685, n6686, n6687, n6688, n6689_1, n6691, n6692, n6693, n6694_1, n6696, n6697, n6698, n6699_1, n6700, n6701, n6703, n6704_1, n6705, n6706, n6708, n6709_1, n6710, n6711, n6712, n6713, n6715, n6716, n6717, n6718, n6720, n6721, n6722, n6723, n6724_1, n6725, n6727, n6728, n6729_1, n6730, n6732, n6733, n6734_1, n6735, n6736, n6737, n6739_1, n6740, n6741, n6742, n6744_1, n6745, n6746, n6747, n6748, n6749_1, n6751, n6752, n6753, n6754_1, n6756, n6757, n6758, n6759_1, n6760, n6761, n6763, n6764_1, n6765, n6766, n6768, n6769_1, n6770, n6771, n6772, n6773, n6775, n6776, n6777, n6778, n6780, n6781, n6782, n6783, n6784_1, n6785, n6787, n6788, n6789_1, n6790, n6888, n6890, n6892, n6894_1, n6896, n6897, n6899_1, n6901, n6903, n6905, n6907, n6909_1, n6911, n6912, n6914_1, n6916, n6918, n6920, n6922, n6923, n6925, n6927, n6929_1, n6931, n6933, n6935, n6937, n6939_1, n6941, n6943, n6945, n6947, n6949_1, n6951, n6953, n6987, n6988, n6989_1, n6990, n6991, n6992, n6994_1, n6995, n6996, n6997, n6999_1, n7000, n7001, n7002, n7003, n7004_1, n7006, n7007, n7008, n7009_1, n7011, n7012, n7013, n7014_1, n7015, n7016, n7018, n7019_1, n7020, n7021, n7023, n7024_1, n7025, n7026, n7027, n7028, n7030, n7031, n7032, n7033, n7035, n7036, n7037, n7038, n7039_1, n7040, n7042, n7043, n7044_1, n7045, n7047, n7048, n7049_1, n7050, n7051, n7052, n7054_1, n7055, n7056, n7057, n7059_1, n7060, n7061, n7062, n7063, n7064_1, n7066, n7067, n7068, n7069_1, n7071, n7072, n7073, n7074_1, n7075, n7076, n7078, n7079_1, n7080, n7081, n7083_1, n7084, n7085, n7086, n7087_1, n7088, n7090, n7091_1, n7092, n7093, n7095_1, n7096, n7097, n7098, n7099_1, n7100, n7102, n7103_1, n7104, n7105, n7107_1, n7108, n7109, n7110, n7111_1, n7112, n7114, n7115_1, n7116, n7117, n7119_1, n7120, n7121, n7122, n7123_1, n7124, n7126, n7127_1, n7128, n7129, n7131_1, n7132, n7133, n7134, n7135_1, n7136, n7138, n7139_1, n7140, n7141, n7143_1, n7144, n7145, n7146, n7147_1, n7148, n7150, n7151_1, n7152, n7153, n7155_1, n7156, n7157, n7158, n7159_1, n7160, n7162, n7163_1, n7164, n7165, n7167_1, n7168, n7169, n7170, n7171_1, n7172, n7174, n7175_1, n7176, n7177, n7179_1, n7180, n7181, n7182, n7183_1, n7184, n7186, n7187_1, n7188, n7189, n7191_1, n7192, n7193, n7194, n7195_1, n7196, n7198, n7199_1, n7200, n7201, n7203_1, n7204, n7205, n7206, n7207_1, n7208, n7210, n7211, n7212_1, n7213, n7215, n7216, n7217_1, n7218, n7219, n7220, n7222_1, n7223, n7224, n7225, n7227_1, n7228, n7229, n7230, n7231, n7232_1, n7234, n7235, n7236, n7237_1, n7239, n7240, n7241, n7242_1, n7243, n7244, n7246, n7247_1, n7248, n7249, n7251, n7252_1, n7253, n7254, n7255, n7256, n7258, n7259, n7260, n7261, n7263, n7264, n7265, n7266, n7267_1, n7268, n7270, n7271, n7272_1, n7273, n7275, n7276, n7277_1, n7278, n7279, n7280, n7282_1, n7283, n7284, n7285, n7287_1, n7288, n7289, n7290, n7291, n7292_1, n7294, n7295, n7296, n7297_1, n7299, n7300, n7301, n7302_1, n7303, n7304, n7306, n7307_1, n7308, n7309, n7311, n7312_1, n7313, n7314, n7315, n7316, n7318, n7319, n7320, n7321, n7323, n7324, n7325, n7326, n7327_1, n7328, n7330, n7331, n7332_1, n7333, n7335, n7336, n7337_1, n7338, n7339, n7340, n7342_1, n7343, n7344, n7345, n7347_1, n7348, n7349, n7350, n7351, n7352_1, n7354, n7355, n7356, n7357_1, n7359, n7360, n7361, n7362_1, n7363, n7364, n7366, n7367_1, n7368, n7369, n7467_1, n7469, n7471, n7473, n7475, n7476, n7478, n7480, n7482_1, n7484, n7486, n7488, n7490, n7491, n7493, n7495, n7497_1, n7499, n7501, n7502_1, n7504, n7506, n7508, n7510, n7512_1, n7514, n7516, n7518, n7520, n7522_1, n7524, n7526, n7528, n7530, n7532_1, n7566, n7567_1, n7568, n7569, n7570, n7571, n7573, n7574, n7575, n7576, n7578, n7579, n7580, n7581, n7582_1, n7583, n7585, n7586, n7587_1, n7588, n7590, n7591, n7592_1, n7593, n7594, n7595, n7597_1, n7598, n7599, n7600, n7602_1, n7603, n7604, n7605, n7606, n7607_1, n7609, n7610, n7611, n7612_1, n7614, n7615, n7616, n7617_1, n7618, n7619, n7621, n7622_1, n7623, n7624, n7626, n7627_1, n7628, n7629, n7630, n7631, n7633, n7634, n7635, n7636, n7638, n7639, n7640, n7641, n7642_1, n7643, n7645, n7646, n7647_1, n7648, n7650, n7651, n7652_1, n7653, n7654, n7655, n7657_1, n7658, n7659, n7660, n7662_1, n7663, n7664, n7665, n7666, n7667_1, n7669, n7670, n7671, n7672_1, n7674, n7675, n7676, n7677_1, n7678, n7679, n7681, n7682_1, n7683, n7684, n7686, n7687_1, n7688, n7689, n7690, n7691, n7693, n7694, n7695, n7696, n7698, n7699, n7700, n7701, n7702_1, n7703, n7705, n7706, n7707_1, n7708, n7710, n7711, n7712_1, n7713, n7714, n7715, n7717_1, n7718, n7719, n7720, n7722_1, n7723, n7724, n7725, n7726, n7727_1, n7729, n7730, n7731, n7732_1, n7734, n7735, n7736, n7737_1, n7738, n7739, n7741, n7742_1, n7743, n7744, n7746, n7747_1, n7748, n7749, n7750, n7751, n7753, n7754, n7755, n7756, n7758, n7759, n7760, n7761, n7762_1, n7763, n7765, n7766, n7767_1, n7768, n7770, n7771, n7772_1, n7773, n7774, n7775, n7777_1, n7778, n7779, n7780, n7782_1, n7783, n7784, n7785, n7786, n7787_1, n7789, n7790, n7791, n7792_1, n7794, n7795, n7796, n7797_1, n7798, n7799, n7801, n7802_1, n7803, n7804, n7806, n7807_1, n7808, n7809, n7810, n7811, n7813, n7814, n7815, n7816, n7818, n7819, n7820, n7821, n7822_1, n7823, n7825, n7826, n7827_1, n7828, n7830, n7831, n7832_1, n7833, n7834, n7835, n7837_1, n7838, n7839, n7840, n7842_1, n7843, n7844, n7845, n7846, n7847_1, n7849, n7850, n7851, n7852_1, n7854, n7855, n7856, n7857_1, n7858, n7859, n7861, n7862_1, n7863, n7864, n7866, n7867_1, n7868, n7869, n7870, n7871, n7873, n7874, n7875, n7876, n7878, n7879, n7880, n7881, n7882_1, n7883, n7885, n7886, n7887_1, n7888, n7890, n7891, n7892_1, n7893, n7894, n7895, n7897_1, n7898, n7899, n7900, n7902_1, n7903, n7904, n7905, n7906, n7907_1, n7909, n7910, n7911, n7912_1, n7914, n7915, n7916, n7917_1, n7918, n7919, n7921, n7922_1, n7923, n7924, n7926, n7927_1, n7928, n7929, n7930, n7931, n7933, n7934, n7935, n7936, n7938, n7939, n7940, n7941, n7942_1, n7943, n7945, n7946, n7947_1, n7948, n8046, n8048, n8050, n8052, n8054, n8055_1, n8057, n8059_1, n8061, n8063_1, n8065, n8067_1, n8069, n8070, n8072, n8074, n8076, n8078, n8080, n8081, n8083_1, n8085, n8087_1, n8089, n8091_1, n8093, n8095_1, n8097, n8099_1, n8101, n8103_1, n8105, n8107_1, n8109, n8111_1, n8145_1, n8146, n8147, n8148, n8149, n8150_1, n8152, n8153, n8154, n8155_1, n8157, n8158, n8159, n8160_1, n8161, n8162, n8164, n8165_1, n8166, n8167, n8169, n8170_1, n8171, n8172, n8173, n8174, n8176, n8177, n8178, n8179, n8181, n8182, n8183, n8184, n8185_1, n8186, n8188, n8189, n8190_1, n8191, n8193, n8194, n8195_1, n8196, n8197, n8198, n8200_1, n8201, n8202, n8203, n8205_1, n8206, n8207, n8208, n8209, n8210_1, n8212, n8213, n8214, n8215_1, n8217, n8218, n8219, n8220_1, n8221, n8222, n8224, n8225_1, n8226, n8227, n8229, n8230_1, n8231, n8232, n8233, n8234, n8236, n8237, n8238, n8239, n8241, n8242, n8243, n8244, n8245_1, n8246, n8248, n8249, n8250_1, n8251, n8253, n8254, n8255_1, n8256, n8257, n8258, n8260_1, n8261, n8262, n8263, n8265_1, n8266, n8267, n8268, n8269, n8270_1, n8272, n8273, n8274, n8275_1, n8277, n8278, n8279, n8280_1, n8281, n8282, n8284, n8285_1, n8286, n8287, n8289, n8290_1, n8291, n8292, n8293, n8294, n8296, n8297, n8298, n8299, n8301, n8302, n8303, n8304, n8305_1, n8306, n8308, n8309, n8310_1, n8311, n8313, n8314, n8315_1, n8316, n8317, n8318, n8320_1, n8321, n8322, n8323, n8325_1, n8326, n8327, n8328, n8329, n8330_1, n8332, n8333, n8334, n8335_1, n8337, n8338, n8339, n8340_1, n8341, n8342, n8344, n8345_1, n8346, n8347, n8349, n8350_1, n8351, n8352, n8353, n8354, n8356, n8357, n8358, n8359, n8361, n8362, n8363, n8364, n8365_1, n8366, n8368, n8369, n8370_1, n8371, n8373, n8374, n8375_1, n8376, n8377, n8378, n8380_1, n8381, n8382, n8383, n8385_1, n8386, n8387, n8388, n8389, n8390_1, n8392, n8393, n8394, n8395_1, n8397, n8398, n8399, n8400_1, n8401, n8402, n8404, n8405_1, n8406, n8407, n8409, n8410_1, n8411, n8412, n8413, n8414, n8416, n8417, n8418, n8419, n8421, n8422, n8423, n8424, n8425_1, n8426, n8428, n8429, n8430_1, n8431, n8433, n8434, n8435_1, n8436, n8437, n8438, n8440_1, n8441, n8442, n8443, n8445_1, n8446, n8447, n8448, n8449, n8450_1, n8452, n8453, n8454, n8455_1, n8457, n8458, n8459, n8460_1, n8461, n8462, n8464, n8465_1, n8466, n8467, n8469, n8470_1, n8471, n8472, n8473, n8474, n8476, n8477, n8478, n8479, n8481, n8482, n8483, n8484, n8485_1, n8486, n8488, n8489, n8490_1, n8491, n8493, n8494, n8495_1, n8496, n8497, n8498, n8500_1, n8501, n8502, n8503, n8505_1, n8506, n8507, n8508, n8509, n8510_1, n8512, n8513, n8514, n8515_1, n8517, n8518, n8519, n8520_1, n8521, n8522, n8524, n8525_1, n8526, n8527, n8625_1, n8627, n8629, n8631, n8633, n8634, n8636, n8638, n8640_1, n8642, n8644, n8646, n8648, n8649, n8651, n8653, n8655_1, n8657, n8659, n8660_1, n8662, n8664, n8666, n8668, n8670_1, n8672, n8674, n8676, n8678, n8680_1, n8682, n8684, n8686, n8688, n8690_1, n8724, n8725_1, n8726, n8727, n8728, n8729, n8731, n8732, n8733, n8734, n8736, n8737, n8738, n8739, n8740_1, n8741, n8743, n8744, n8745_1, n8746, n8748, n8749, n8750_1, n8751, n8752, n8753, n8755_1, n8756, n8757, n8758, n8760_1, n8761, n8762, n8763, n8764, n8765_1, n8767, n8768, n8769, n8770_1, n8772, n8773, n8774, n8775_1, n8776, n8777, n8779, n8780_1, n8781, n8782, n8784, n8785_1, n8786, n8787, n8788, n8789, n8791, n8792, n8793, n8794, n8796, n8797, n8798, n8799, n8800_1, n8801, n8803, n8804, n8805_1, n8806, n8808, n8809, n8810_1, n8811, n8812, n8813, n8815_1, n8816, n8817, n8818, n8820_1, n8821, n8822, n8823, n8824, n8825_1, n8827, n8828, n8829, n8830_1, n8832, n8833, n8834, n8835_1, n8836, n8837, n8839, n8840_1, n8841, n8842, n8844, n8845_1, n8846, n8847, n8848, n8849, n8851, n8852, n8853, n8854, n8856, n8857, n8858, n8859, n8860_1, n8861, n8863, n8864, n8865_1, n8866, n8868, n8869, n8870_1, n8871, n8872, n8873, n8875_1, n8876, n8877, n8878, n8880_1, n8881, n8882, n8883, n8884, n8885_1, n8887, n8888, n8889, n8890_1, n8892, n8893, n8894, n8895_1, n8896, n8897, n8899, n8900_1, n8901, n8902, n8904, n8905_1, n8906, n8907, n8908, n8909, n8911, n8912, n8913, n8914, n8916, n8917, n8918, n8919, n8920_1, n8921, n8923, n8924, n8925_1, n8926, n8928, n8929, n8930_1, n8931, n8932, n8933, n8935_1, n8936, n8937, n8938, n8940, n8941, n8942, n8943_1, n8944, n8945, n8947_1, n8948, n8949, n8950, n8952, n8953, n8954, n8955_1, n8956, n8957, n8959_1, n8960, n8961, n8962, n8964, n8965, n8966, n8967_1, n8968, n8969, n8971_1, n8972, n8973, n8974, n8976, n8977, n8978, n8979_1, n8980, n8981, n8983_1, n8984, n8985, n8986, n8988, n8989, n8990, n8991_1, n8992, n8993, n8995_1, n8996, n8997, n8998, n9000, n9001, n9002, n9003_1, n9004, n9005, n9007_1, n9008, n9009, n9010, n9012, n9013, n9014, n9015_1, n9016, n9017, n9019_1, n9020, n9021, n9022, n9024, n9025, n9026, n9027_1, n9028, n9029, n9031_1, n9032, n9033, n9034, n9036, n9037, n9038, n9039_1, n9040, n9041, n9043_1, n9044, n9045, n9046, n9048, n9049, n9050, n9051_1, n9052, n9053, n9055_1, n9056, n9057, n9058, n9060, n9061, n9062, n9063, n9064, n9065, n9067, n9068, n9069, n9070, n9072, n9073, n9074, n9075, n9076, n9077, n9079, n9080, n9081, n9082, n9084, n9085, n9086, n9087, n9088, n9089, n9091, n9092, n9093, n9094, n9096, n9097, n9098, n9099, n9100, n9101, n9103, n9104, n9105, n9106, n9204, n9206, n9208, n9210, n9212, n9213, n9215, n9217, n9219, n9221, n9223, n9225, n9227, n9228, n9230, n9232, n9234, n9236, n9238, n9239, n9241, n9243, n9245, n9247, n9249, n9251, n9253, n9255, n9257, n9259, n9261, n9263, n9265, n9267, n9269, n9303, n9304, n9305, n9306, n9307, n9308, n9310, n9311, n9312, n9313, n9315, n9316, n9317, n9318, n9319, n9320, n9322, n9323, n9324, n9325, n9327, n9328, n9329, n9330, n9331, n9332, n9334, n9335, n9336, n9337, n9339, n9340, n9341, n9342, n9343, n9344, n9346, n9347, n9348, n9349, n9351, n9352, n9353, n9354, n9355, n9356, n9358, n9359, n9360, n9361, n9363, n9364, n9365, n9366, n9367, n9368, n9370, n9371, n9372, n9373, n9375, n9376, n9377, n9378, n9379, n9380, n9382, n9383, n9384, n9385, n9387, n9388, n9389, n9390, n9391, n9392, n9394, n9395, n9396, n9397, n9399, n9400, n9401, n9402, n9403, n9404, n9406, n9407, n9408, n9409, n9411, n9412, n9413, n9414, n9415, n9416, n9418, n9419, n9420, n9421, n9423, n9424, n9425, n9426, n9427, n9428, n9430, n9431, n9432, n9433, n9435, n9436, n9437, n9438, n9439, n9440, n9442, n9443, n9444, n9445, n9447, n9448, n9449, n9450, n9451, n9452, n9454, n9455, n9456, n9457, n9459, n9460, n9461, n9462, n9463, n9464, n9466, n9467, n9468, n9469, n9471, n9472, n9473, n9474, n9475, n9476, n9478, n9479, n9480, n9481, n9483, n9484, n9485, n9486, n9487, n9488, n9490, n9491, n9492, n9493, n9495, n9496, n9497, n9498, n9499, n9500, n9502, n9503, n9504, n9505, n9507, n9508, n9509, n9510, n9511, n9512, n9514, n9515, n9516, n9517, n9519, n9520, n9521, n9522, n9523, n9524, n9526, n9527, n9528, n9529, n9531, n9532, n9533, n9534, n9535, n9536, n9538, n9539, n9540, n9541, n9543, n9544, n9545, n9546, n9547, n9548, n9550, n9551, n9552, n9553, n9555, n9556, n9557, n9558, n9559, n9560, n9562, n9563, n9564, n9565, n9567, n9568, n9569, n9570, n9571, n9572, n9574, n9575, n9576, n9577, n9579, n9580, n9581, n9582, n9583, n9584, n9586, n9587, n9588, n9589, n9591, n9592, n9593, n9594, n9595, n9596, n9598, n9599, n9600, n9601, n9603, n9604, n9605, n9606, n9607, n9608, n9610, n9611, n9612, n9613, n9615, n9616, n9617, n9618, n9619, n9620, n9622, n9623, n9624, n9625, n9627, n9628, n9629, n9630, n9631, n9632, n9634, n9635, n9636, n9637, n9639, n9640, n9641, n9642, n9643, n9644, n9646, n9647, n9648, n9649, n9651, n9652, n9653, n9654, n9655, n9656, n9658, n9659, n9660, n9661, n9663, n9664, n9665, n9666, n9667, n9668, n9670, n9671, n9672, n9673, n9675, n9676, n9677, n9678, n9679, n9680, n9682, n9683, n9684, n9685, n9783, n9785, n9787, n9789, n9791, n9792, n9794, n9796, n9798, n9800, n9802, n9804, n9806, n9807, n9809, n9811, n9813, n9815, n9817, n9818, n9820, n9822, n9824, n9826, n9828, n9830, n9832, n9834, n9836, n9838, n9840, n9842, n9844, n9846, n9848, n9882, n9883, n9884, n9885, n9886, n9887, n9889, n9890, n9891, n9892, n9894, n9895, n9896, n9897, n9898, n9899, n9901, n9902, n9903, n9904, n9906, n9907, n9908, n9909, n9910, n9911, n9913, n9914, n9915, n9916, n9918, n9919, n9920, n9921, n9922, n9923, n9925, n9926, n9927, n9928, n9930, n9931, n9932, n9933, n9934, n9935, n9937, n9938, n9939, n9940, n9942, n9943, n9944, n9945, n9946, n9947, n9949, n9950, n9951, n9952, n9954, n9955, n9956, n9957, n9958, n9959, n9961, n9962, n9963, n9964, n9966, n9967, n9968, n9969, n9970, n9971, n9973, n9974, n9975, n9976, n9978, n9979, n9980, n9981, n9982, n9983, n9985, n9986, n9987, n9988, n9990, n9991, n9992, n9993, n9994, n9995, n9997, n9998, n9999, n10000, n10002, n10003, n10004, n10005, n10006, n10007, n10009, n10010, n10011, n10012, n10014, n10015, n10016, n10017, n10018, n10019, n10021, n10022, n10023, n10024, n10026, n10027, n10028, n10029, n10030, n10031, n10033, n10034, n10035, n10036, n10038, n10039, n10040, n10041, n10042, n10043, n10045, n10046, n10047, n10048, n10050, n10051, n10052, n10053, n10054, n10055, n10057, n10058, n10059, n10060, n10062, n10063, n10064, n10065, n10066, n10067, n10069, n10070, n10071, n10072, n10074, n10075, n10076, n10077, n10078, n10079, n10081, n10082, n10083, n10084, n10086, n10087, n10088, n10089, n10090, n10091, n10093, n10094, n10095, n10096, n10098, n10099, n10100, n10101, n10102, n10103, n10105, n10106, n10107, n10108, n10110, n10111, n10112, n10113, n10114, n10115, n10117, n10118, n10119, n10120, n10122, n10123, n10124, n10125, n10126, n10127, n10129, n10130, n10131, n10132, n10134, n10135, n10136, n10137, n10138, n10139, n10141, n10142, n10143, n10144, n10146, n10147, n10148, n10149, n10150, n10151, n10153, n10154, n10155, n10156, n10158, n10159, n10160, n10161, n10162, n10163, n10165, n10166, n10167, n10168, n10170, n10171, n10172, n10173, n10174, n10175, n10177, n10178, n10179, n10180, n10182, n10183, n10184, n10185, n10186, n10187, n10189, n10190, n10191, n10192, n10194, n10195, n10196, n10197, n10198, n10199, n10201, n10202, n10203, n10204, n10206, n10207, n10208, n10209, n10210, n10211, n10213, n10214, n10215, n10216, n10218, n10219, n10220, n10221, n10222, n10223, n10225, n10226, n10227, n10228, n10230, n10231, n10232, n10233, n10234, n10235, n10237, n10238, n10239, n10240, n10242, n10243, n10244, n10245, n10246, n10247, n10249, n10250, n10251, n10252, n10254, n10255, n10256, n10257, n10258, n10259, n10261, n10262, n10263, n10264, n10362, n10364, n10366, n10368, n10370, n10371, n10373, n10375, n10377, n10379, n10381, n10383, n10385, n10386, n10388, n10390, n10392, n10394, n10396, n10397, n10399, n10401, n10403, n10405, n10407, n10409, n10411, n10413, n10415, n10417, n10419, n10421, n10423, n10425, n10427, n10461, n10462, n10463, n10464, n10465, n10467, n10468, n10469, n10470, n10471, n10473, n10474, n10475, n10476, n10477, n10479, n10480, n10481, n10482, n10483, n10485, n10486, n10487, n10488, n10489, n10491, n10492, n10493, n10494, n10495, n10497, n10498, n10499, n10500, n10501, n10503, n10504, n10505, n10506, n10507, n10509, n10510, n10511, n10512, n10513, n10515, n10516, n10517, n10518, n10519, n10521, n10522, n10523, n10524, n10525, n10527, n10528, n10529, n10530, n10531, n10533, n10534, n10535, n10536, n10537, n10539, n10540, n10541, n10542, n10543, n10545, n10546, n10547, n10548, n10549, n10551, n10552, n10553, n10554, n10555, n10557, n10558, n10559, n10560, n10561, n10563, n10564, n10565, n10566, n10567, n10569, n10570, n10571, n10572, n10573, n10575, n10576, n10577, n10578, n10579, n10581, n10582, n10583, n10584, n10585, n10587, n10588, n10589, n10590, n10591, n10593, n10594, n10595, n10596, n10597, n10599, n10600, n10601, n10602, n10603, n10605, n10606, n10607, n10608, n10609, n10611, n10612, n10613, n10614, n10615, n10617, n10618, n10619, n10620, n10621, n10623, n10624, n10625, n10626, n10627, n10629, n10630, n10631, n10632, n10633, n10635, n10636, n10637, n10638, n10639, n10641, n10642, n10643, n10644, n10645, n10647, n10648, n10649, n10650, n10651, n10749, n10751, n10753, n10755, n10757, n10758, n10760, n10762, n10764, n10766, n10768, n10770, n10772, n10773, n10775, n10777, n10779, n10781, n10783, n10784, n10786, n10788, n10790, n10792, n10794, n10796, n10798, n10800, n10802, n10804, n10806, n10808, n10810, n10812, n10814;
INVX1    g0000(.A(TM0), .Y(n5539));
XOR2X1   g0001(.A(WX645), .B(TM1), .Y(n5540));
XOR2X1   g0002(.A(n5540), .B(WX709), .Y(n5541_1));
INVX1    g0003(.A(WX773), .Y(n5542));
XOR2X1   g0004(.A(WX837), .B(n5542), .Y(n5543));
XOR2X1   g0005(.A(n5543), .B(n5541_1), .Y(n5544));
OR2X1    g0006(.A(n5544), .B(TM0), .Y(n5545));
XOR2X1   g0007(.A(n5544), .B(WX485), .Y(n5546_1));
OAI21X1  g0008(.A0(n5546_1), .A1(n5539), .B0(n5545), .Y(DATA_9_31));
XOR2X1   g0009(.A(WX647), .B(TM1), .Y(n5548));
XOR2X1   g0010(.A(n5548), .B(WX711), .Y(n5549));
INVX1    g0011(.A(WX775), .Y(n5550));
XOR2X1   g0012(.A(WX839), .B(n5550), .Y(n5551_1));
XOR2X1   g0013(.A(n5551_1), .B(n5549), .Y(n5552));
OR2X1    g0014(.A(n5552), .B(TM0), .Y(n5553));
XOR2X1   g0015(.A(n5552), .B(WX487), .Y(n5554));
OAI21X1  g0016(.A0(n5554), .A1(n5539), .B0(n5553), .Y(DATA_9_30));
XOR2X1   g0017(.A(WX649), .B(TM1), .Y(n5556_1));
XOR2X1   g0018(.A(n5556_1), .B(WX713), .Y(n5557));
INVX1    g0019(.A(WX777), .Y(n5558));
XOR2X1   g0020(.A(WX841), .B(n5558), .Y(n5559));
XOR2X1   g0021(.A(n5559), .B(n5557), .Y(n5560));
OR2X1    g0022(.A(n5560), .B(TM0), .Y(n5561_1));
XOR2X1   g0023(.A(n5560), .B(WX489), .Y(n5562));
OAI21X1  g0024(.A0(n5562), .A1(n5539), .B0(n5561_1), .Y(DATA_9_29));
XOR2X1   g0025(.A(WX651), .B(TM1), .Y(n5564));
XOR2X1   g0026(.A(n5564), .B(WX715), .Y(n5565));
INVX1    g0027(.A(WX779), .Y(n5566_1));
XOR2X1   g0028(.A(WX843), .B(n5566_1), .Y(n5567));
XOR2X1   g0029(.A(n5567), .B(n5565), .Y(n5568));
OR2X1    g0030(.A(n5568), .B(TM0), .Y(n5569));
XOR2X1   g0031(.A(n5568), .B(WX491), .Y(n5570));
OAI21X1  g0032(.A0(n5570), .A1(n5539), .B0(n5569), .Y(DATA_9_28));
XOR2X1   g0033(.A(WX653), .B(TM1), .Y(n5572));
XOR2X1   g0034(.A(n5572), .B(WX717), .Y(n5573));
INVX1    g0035(.A(WX781), .Y(n5574));
XOR2X1   g0036(.A(WX845), .B(n5574), .Y(n5575));
XOR2X1   g0037(.A(n5575), .B(n5573), .Y(n5576_1));
OR2X1    g0038(.A(n5576_1), .B(TM0), .Y(n5577));
XOR2X1   g0039(.A(n5576_1), .B(WX493), .Y(n5578));
OAI21X1  g0040(.A0(n5578), .A1(n5539), .B0(n5577), .Y(DATA_9_27));
XOR2X1   g0041(.A(WX655), .B(TM1), .Y(n5580));
XOR2X1   g0042(.A(n5580), .B(WX719), .Y(n5581_1));
INVX1    g0043(.A(WX783), .Y(n5582));
XOR2X1   g0044(.A(WX847), .B(n5582), .Y(n5583));
XOR2X1   g0045(.A(n5583), .B(n5581_1), .Y(n5584));
OR2X1    g0046(.A(n5584), .B(TM0), .Y(n5585));
XOR2X1   g0047(.A(n5584), .B(WX495), .Y(n5586_1));
OAI21X1  g0048(.A0(n5586_1), .A1(n5539), .B0(n5585), .Y(DATA_9_26));
XOR2X1   g0049(.A(WX657), .B(TM1), .Y(n5588));
XOR2X1   g0050(.A(n5588), .B(WX721), .Y(n5589));
INVX1    g0051(.A(WX785), .Y(n5590));
XOR2X1   g0052(.A(WX849), .B(n5590), .Y(n5591_1));
XOR2X1   g0053(.A(n5591_1), .B(n5589), .Y(n5592));
OR2X1    g0054(.A(n5592), .B(TM0), .Y(n5593));
XOR2X1   g0055(.A(n5592), .B(WX497), .Y(n5594));
OAI21X1  g0056(.A0(n5594), .A1(n5539), .B0(n5593), .Y(DATA_9_25));
XOR2X1   g0057(.A(WX659), .B(TM1), .Y(n5596_1));
XOR2X1   g0058(.A(n5596_1), .B(WX723), .Y(n5597));
INVX1    g0059(.A(WX787), .Y(n5598));
XOR2X1   g0060(.A(WX851), .B(n5598), .Y(n5599));
XOR2X1   g0061(.A(n5599), .B(n5597), .Y(n5600));
OR2X1    g0062(.A(n5600), .B(TM0), .Y(n5601_1));
XOR2X1   g0063(.A(n5600), .B(WX499), .Y(n5602));
OAI21X1  g0064(.A0(n5602), .A1(n5539), .B0(n5601_1), .Y(DATA_9_24));
XOR2X1   g0065(.A(WX661), .B(TM1), .Y(n5604));
XOR2X1   g0066(.A(n5604), .B(WX725), .Y(n5605));
INVX1    g0067(.A(WX789), .Y(n5606_1));
XOR2X1   g0068(.A(WX853), .B(n5606_1), .Y(n5607));
XOR2X1   g0069(.A(n5607), .B(n5605), .Y(n5608));
OR2X1    g0070(.A(n5608), .B(TM0), .Y(n5609));
XOR2X1   g0071(.A(n5608), .B(WX501), .Y(n5610));
OAI21X1  g0072(.A0(n5610), .A1(n5539), .B0(n5609), .Y(DATA_9_23));
XOR2X1   g0073(.A(WX663), .B(TM1), .Y(n5612));
XOR2X1   g0074(.A(n5612), .B(WX727), .Y(n5613));
INVX1    g0075(.A(WX791), .Y(n5614));
XOR2X1   g0076(.A(WX855), .B(n5614), .Y(n5615));
XOR2X1   g0077(.A(n5615), .B(n5613), .Y(n5616_1));
OR2X1    g0078(.A(n5616_1), .B(TM0), .Y(n5617));
XOR2X1   g0079(.A(n5616_1), .B(WX503), .Y(n5618));
OAI21X1  g0080(.A0(n5618), .A1(n5539), .B0(n5617), .Y(DATA_9_22));
XOR2X1   g0081(.A(WX665), .B(TM1), .Y(n5620));
XOR2X1   g0082(.A(n5620), .B(WX729), .Y(n5621_1));
INVX1    g0083(.A(WX793), .Y(n5622));
XOR2X1   g0084(.A(WX857), .B(n5622), .Y(n5623));
XOR2X1   g0085(.A(n5623), .B(n5621_1), .Y(n5624));
OR2X1    g0086(.A(n5624), .B(TM0), .Y(n5625));
XOR2X1   g0087(.A(n5624), .B(WX505), .Y(n5626_1));
OAI21X1  g0088(.A0(n5626_1), .A1(n5539), .B0(n5625), .Y(DATA_9_21));
XOR2X1   g0089(.A(WX667), .B(TM1), .Y(n5628));
XOR2X1   g0090(.A(n5628), .B(WX731), .Y(n5629));
INVX1    g0091(.A(WX795), .Y(n5630));
XOR2X1   g0092(.A(WX859), .B(n5630), .Y(n5631_1));
XOR2X1   g0093(.A(n5631_1), .B(n5629), .Y(n5632));
OR2X1    g0094(.A(n5632), .B(TM0), .Y(n5633));
XOR2X1   g0095(.A(n5632), .B(WX507), .Y(n5634));
OAI21X1  g0096(.A0(n5634), .A1(n5539), .B0(n5633), .Y(DATA_9_20));
XOR2X1   g0097(.A(WX669), .B(TM1), .Y(n5636_1));
XOR2X1   g0098(.A(n5636_1), .B(WX733), .Y(n5637));
INVX1    g0099(.A(WX797), .Y(n5638));
XOR2X1   g0100(.A(WX861), .B(n5638), .Y(n5639));
XOR2X1   g0101(.A(n5639), .B(n5637), .Y(n5640));
OR2X1    g0102(.A(n5640), .B(TM0), .Y(n5641_1));
XOR2X1   g0103(.A(n5640), .B(WX509), .Y(n5642));
OAI21X1  g0104(.A0(n5642), .A1(n5539), .B0(n5641_1), .Y(DATA_9_19));
XOR2X1   g0105(.A(WX671), .B(TM1), .Y(n5644));
XOR2X1   g0106(.A(n5644), .B(WX735), .Y(n5645));
INVX1    g0107(.A(WX799), .Y(n5646_1));
XOR2X1   g0108(.A(WX863), .B(n5646_1), .Y(n5647));
XOR2X1   g0109(.A(n5647), .B(n5645), .Y(n5648));
OR2X1    g0110(.A(n5648), .B(TM0), .Y(n5649));
XOR2X1   g0111(.A(n5648), .B(WX511), .Y(n5650));
OAI21X1  g0112(.A0(n5650), .A1(n5539), .B0(n5649), .Y(DATA_9_18));
XOR2X1   g0113(.A(WX673), .B(TM1), .Y(n5652));
XOR2X1   g0114(.A(n5652), .B(WX737), .Y(n5653));
INVX1    g0115(.A(WX801), .Y(n5654));
XOR2X1   g0116(.A(WX865), .B(n5654), .Y(n5655));
XOR2X1   g0117(.A(n5655), .B(n5653), .Y(n5656_1));
OR2X1    g0118(.A(n5656_1), .B(TM0), .Y(n5657));
XOR2X1   g0119(.A(n5656_1), .B(WX513), .Y(n5658));
OAI21X1  g0120(.A0(n5658), .A1(n5539), .B0(n5657), .Y(DATA_9_17));
XOR2X1   g0121(.A(WX675), .B(TM1), .Y(n5660));
XOR2X1   g0122(.A(n5660), .B(WX739), .Y(n5661_1));
INVX1    g0123(.A(WX803), .Y(n5662));
XOR2X1   g0124(.A(WX867), .B(n5662), .Y(n5663));
XOR2X1   g0125(.A(n5663), .B(n5661_1), .Y(n5664));
OR2X1    g0126(.A(n5664), .B(TM0), .Y(n5665));
XOR2X1   g0127(.A(n5664), .B(WX515), .Y(n5666_1));
OAI21X1  g0128(.A0(n5666_1), .A1(n5539), .B0(n5665), .Y(DATA_9_16));
XOR2X1   g0129(.A(WX677), .B(TM0), .Y(n5668));
XOR2X1   g0130(.A(n5668), .B(WX741), .Y(n5669));
INVX1    g0131(.A(WX805), .Y(n5670));
XOR2X1   g0132(.A(WX869), .B(n5670), .Y(n5671_1));
XOR2X1   g0133(.A(n5671_1), .B(n5669), .Y(n5672));
OR2X1    g0134(.A(n5672), .B(TM0), .Y(n5673));
XOR2X1   g0135(.A(n5672), .B(WX517), .Y(n5674));
OAI21X1  g0136(.A0(n5674), .A1(n5539), .B0(n5673), .Y(DATA_9_15));
XOR2X1   g0137(.A(WX679), .B(TM0), .Y(n5676_1));
XOR2X1   g0138(.A(n5676_1), .B(WX743), .Y(n5677));
INVX1    g0139(.A(WX807), .Y(n5678));
XOR2X1   g0140(.A(WX871), .B(n5678), .Y(n5679));
XOR2X1   g0141(.A(n5679), .B(n5677), .Y(n5680));
OR2X1    g0142(.A(n5680), .B(TM0), .Y(n5681_1));
XOR2X1   g0143(.A(n5680), .B(WX519), .Y(n5682));
OAI21X1  g0144(.A0(n5682), .A1(n5539), .B0(n5681_1), .Y(DATA_9_14));
XOR2X1   g0145(.A(WX681), .B(TM0), .Y(n5684));
XOR2X1   g0146(.A(n5684), .B(WX745), .Y(n5685));
INVX1    g0147(.A(WX809), .Y(n5686_1));
XOR2X1   g0148(.A(WX873), .B(n5686_1), .Y(n5687));
XOR2X1   g0149(.A(n5687), .B(n5685), .Y(n5688));
OR2X1    g0150(.A(n5688), .B(TM0), .Y(n5689));
XOR2X1   g0151(.A(n5688), .B(WX521), .Y(n5690));
OAI21X1  g0152(.A0(n5690), .A1(n5539), .B0(n5689), .Y(DATA_9_13));
XOR2X1   g0153(.A(WX683), .B(TM0), .Y(n5692));
XOR2X1   g0154(.A(n5692), .B(WX747), .Y(n5693));
INVX1    g0155(.A(WX811), .Y(n5694));
XOR2X1   g0156(.A(WX875), .B(n5694), .Y(n5695));
XOR2X1   g0157(.A(n5695), .B(n5693), .Y(n5696_1));
OR2X1    g0158(.A(n5696_1), .B(TM0), .Y(n5697));
XOR2X1   g0159(.A(n5696_1), .B(WX523), .Y(n5698));
OAI21X1  g0160(.A0(n5698), .A1(n5539), .B0(n5697), .Y(DATA_9_12));
XOR2X1   g0161(.A(WX685), .B(TM0), .Y(n5700));
XOR2X1   g0162(.A(n5700), .B(WX749), .Y(n5701_1));
INVX1    g0163(.A(WX813), .Y(n5702));
XOR2X1   g0164(.A(WX877), .B(n5702), .Y(n5703));
XOR2X1   g0165(.A(n5703), .B(n5701_1), .Y(n5704));
OR2X1    g0166(.A(n5704), .B(TM0), .Y(n5705));
XOR2X1   g0167(.A(n5704), .B(WX525), .Y(n5706_1));
OAI21X1  g0168(.A0(n5706_1), .A1(n5539), .B0(n5705), .Y(DATA_9_11));
XOR2X1   g0169(.A(WX687), .B(TM0), .Y(n5708));
XOR2X1   g0170(.A(n5708), .B(WX751), .Y(n5709));
INVX1    g0171(.A(WX815), .Y(n5710));
XOR2X1   g0172(.A(WX879), .B(n5710), .Y(n5711_1));
XOR2X1   g0173(.A(n5711_1), .B(n5709), .Y(n5712));
OR2X1    g0174(.A(n5712), .B(TM0), .Y(n5713));
XOR2X1   g0175(.A(n5712), .B(WX527), .Y(n5714));
OAI21X1  g0176(.A0(n5714), .A1(n5539), .B0(n5713), .Y(DATA_9_10));
XOR2X1   g0177(.A(WX689), .B(TM0), .Y(n5716_1));
XOR2X1   g0178(.A(n5716_1), .B(WX753), .Y(n5717));
INVX1    g0179(.A(WX817), .Y(n5718));
XOR2X1   g0180(.A(WX881), .B(n5718), .Y(n5719));
XOR2X1   g0181(.A(n5719), .B(n5717), .Y(n5720));
OR2X1    g0182(.A(n5720), .B(TM0), .Y(n5721_1));
XOR2X1   g0183(.A(n5720), .B(WX529), .Y(n5722));
OAI21X1  g0184(.A0(n5722), .A1(n5539), .B0(n5721_1), .Y(DATA_9_9));
XOR2X1   g0185(.A(WX691), .B(TM0), .Y(n5724));
XOR2X1   g0186(.A(n5724), .B(WX755), .Y(n5725));
INVX1    g0187(.A(WX819), .Y(n5726_1));
XOR2X1   g0188(.A(WX883), .B(n5726_1), .Y(n5727));
XOR2X1   g0189(.A(n5727), .B(n5725), .Y(n5728));
OR2X1    g0190(.A(n5728), .B(TM0), .Y(n5729));
XOR2X1   g0191(.A(n5728), .B(WX531), .Y(n5730));
OAI21X1  g0192(.A0(n5730), .A1(n5539), .B0(n5729), .Y(DATA_9_8));
XOR2X1   g0193(.A(WX693), .B(TM0), .Y(n5732));
XOR2X1   g0194(.A(n5732), .B(WX757), .Y(n5733));
INVX1    g0195(.A(WX821), .Y(n5734));
XOR2X1   g0196(.A(WX885), .B(n5734), .Y(n5735));
XOR2X1   g0197(.A(n5735), .B(n5733), .Y(n5736_1));
OR2X1    g0198(.A(n5736_1), .B(TM0), .Y(n5737));
XOR2X1   g0199(.A(n5736_1), .B(WX533), .Y(n5738));
OAI21X1  g0200(.A0(n5738), .A1(n5539), .B0(n5737), .Y(DATA_9_7));
XOR2X1   g0201(.A(WX695), .B(TM0), .Y(n5740));
XOR2X1   g0202(.A(n5740), .B(WX759), .Y(n5741_1));
INVX1    g0203(.A(WX823), .Y(n5742));
XOR2X1   g0204(.A(WX887), .B(n5742), .Y(n5743));
XOR2X1   g0205(.A(n5743), .B(n5741_1), .Y(n5744));
OR2X1    g0206(.A(n5744), .B(TM0), .Y(n5745));
XOR2X1   g0207(.A(n5744), .B(WX535), .Y(n5746_1));
OAI21X1  g0208(.A0(n5746_1), .A1(n5539), .B0(n5745), .Y(DATA_9_6));
XOR2X1   g0209(.A(WX697), .B(TM0), .Y(n5748));
XOR2X1   g0210(.A(n5748), .B(WX761), .Y(n5749));
INVX1    g0211(.A(WX825), .Y(n5750));
XOR2X1   g0212(.A(WX889), .B(n5750), .Y(n5751_1));
XOR2X1   g0213(.A(n5751_1), .B(n5749), .Y(n5752));
OR2X1    g0214(.A(n5752), .B(TM0), .Y(n5753));
XOR2X1   g0215(.A(n5752), .B(WX537), .Y(n5754));
OAI21X1  g0216(.A0(n5754), .A1(n5539), .B0(n5753), .Y(DATA_9_5));
XOR2X1   g0217(.A(WX699), .B(TM0), .Y(n5756_1));
XOR2X1   g0218(.A(n5756_1), .B(WX763), .Y(n5757));
INVX1    g0219(.A(WX827), .Y(n5758));
XOR2X1   g0220(.A(WX891), .B(n5758), .Y(n5759));
XOR2X1   g0221(.A(n5759), .B(n5757), .Y(n5760));
OR2X1    g0222(.A(n5760), .B(TM0), .Y(n5761_1));
XOR2X1   g0223(.A(n5760), .B(WX539), .Y(n5762));
OAI21X1  g0224(.A0(n5762), .A1(n5539), .B0(n5761_1), .Y(DATA_9_4));
XOR2X1   g0225(.A(WX701), .B(TM0), .Y(n5764));
XOR2X1   g0226(.A(n5764), .B(WX765), .Y(n5765));
INVX1    g0227(.A(WX829), .Y(n5766_1));
XOR2X1   g0228(.A(WX893), .B(n5766_1), .Y(n5767));
XOR2X1   g0229(.A(n5767), .B(n5765), .Y(n5768));
OR2X1    g0230(.A(n5768), .B(TM0), .Y(n5769));
XOR2X1   g0231(.A(n5768), .B(WX541), .Y(n5770));
OAI21X1  g0232(.A0(n5770), .A1(n5539), .B0(n5769), .Y(DATA_9_3));
XOR2X1   g0233(.A(WX703), .B(TM0), .Y(n5772));
XOR2X1   g0234(.A(n5772), .B(WX767), .Y(n5773));
INVX1    g0235(.A(WX831), .Y(n5774));
XOR2X1   g0236(.A(WX895), .B(n5774), .Y(n5775));
XOR2X1   g0237(.A(n5775), .B(n5773), .Y(n5776_1));
OR2X1    g0238(.A(n5776_1), .B(TM0), .Y(n5777));
XOR2X1   g0239(.A(n5776_1), .B(WX543), .Y(n5778));
OAI21X1  g0240(.A0(n5778), .A1(n5539), .B0(n5777), .Y(DATA_9_2));
XOR2X1   g0241(.A(WX705), .B(TM0), .Y(n5780));
XOR2X1   g0242(.A(n5780), .B(WX769), .Y(n5781_1));
INVX1    g0243(.A(WX833), .Y(n5782));
XOR2X1   g0244(.A(WX897), .B(n5782), .Y(n5783));
XOR2X1   g0245(.A(n5783), .B(n5781_1), .Y(n5784));
OR2X1    g0246(.A(n5784), .B(TM0), .Y(n5785));
XOR2X1   g0247(.A(n5784), .B(WX545), .Y(n5786_1));
OAI21X1  g0248(.A0(n5786_1), .A1(n5539), .B0(n5785), .Y(DATA_9_1));
XOR2X1   g0249(.A(WX707), .B(TM0), .Y(n5788));
XOR2X1   g0250(.A(n5788), .B(WX771), .Y(n5789));
INVX1    g0251(.A(WX835), .Y(n5790));
XOR2X1   g0252(.A(WX899), .B(n5790), .Y(n5791_1));
XOR2X1   g0253(.A(n5791_1), .B(n5789), .Y(n5792));
OR2X1    g0254(.A(n5792), .B(TM0), .Y(n5793));
XOR2X1   g0255(.A(n5792), .B(WX547), .Y(n5794));
OAI21X1  g0256(.A0(n5794), .A1(n5539), .B0(n5793), .Y(DATA_9_0));
AND2X1   g0257(.A(WX487), .B(RESET), .Y(n711));
AND2X1   g0258(.A(WX489), .B(RESET), .Y(n716));
AND2X1   g0259(.A(WX491), .B(RESET), .Y(n721));
AND2X1   g0260(.A(WX493), .B(RESET), .Y(n726));
AND2X1   g0261(.A(WX495), .B(RESET), .Y(n731));
AND2X1   g0262(.A(WX497), .B(RESET), .Y(n736));
AND2X1   g0263(.A(WX499), .B(RESET), .Y(n741));
AND2X1   g0264(.A(WX501), .B(RESET), .Y(n746));
AND2X1   g0265(.A(WX503), .B(RESET), .Y(n751));
AND2X1   g0266(.A(WX505), .B(RESET), .Y(n756));
AND2X1   g0267(.A(WX507), .B(RESET), .Y(n761));
AND2X1   g0268(.A(WX509), .B(RESET), .Y(n766));
AND2X1   g0269(.A(WX511), .B(RESET), .Y(n771));
AND2X1   g0270(.A(WX513), .B(RESET), .Y(n776));
AND2X1   g0271(.A(WX515), .B(RESET), .Y(n781));
AND2X1   g0272(.A(WX517), .B(RESET), .Y(n786));
AND2X1   g0273(.A(WX519), .B(RESET), .Y(n791));
AND2X1   g0274(.A(WX521), .B(RESET), .Y(n796));
AND2X1   g0275(.A(WX523), .B(RESET), .Y(n801));
AND2X1   g0276(.A(WX525), .B(RESET), .Y(n806));
AND2X1   g0277(.A(WX527), .B(RESET), .Y(n811));
AND2X1   g0278(.A(WX529), .B(RESET), .Y(n816));
AND2X1   g0279(.A(WX531), .B(RESET), .Y(n821));
AND2X1   g0280(.A(WX533), .B(RESET), .Y(n826));
AND2X1   g0281(.A(WX535), .B(RESET), .Y(n831));
AND2X1   g0282(.A(WX537), .B(RESET), .Y(n836));
AND2X1   g0283(.A(WX539), .B(RESET), .Y(n841));
AND2X1   g0284(.A(WX541), .B(RESET), .Y(n846));
AND2X1   g0285(.A(WX543), .B(RESET), .Y(n851));
AND2X1   g0286(.A(WX545), .B(RESET), .Y(n856));
AND2X1   g0287(.A(WX547), .B(RESET), .Y(n861));
INVX1    g0288(.A(RESET), .Y(n5827));
NOR2X1   g0289(.A(WX485), .B(n5827), .Y(n866));
INVX1    g0290(.A(CRC_OUT_9_31), .Y(n5829));
XOR2X1   g0291(.A(WX1938), .B(TM1), .Y(n5830));
XOR2X1   g0292(.A(n5830), .B(WX2002), .Y(n5831_1));
INVX1    g0293(.A(WX2066), .Y(n5832));
XOR2X1   g0294(.A(WX2130), .B(n5832), .Y(n5833));
XOR2X1   g0295(.A(n5833), .B(n5831_1), .Y(n5834));
MX2X1    g0296(.A(n5829), .B(n5834), .S0(n5539), .Y(n5836_1));
INVX1    g0297(.A(WX485), .Y(n5837));
MX2X1    g0298(.A(n5837), .B(n5544), .S0(n5539), .Y(n5838));
MX2X1    g0299(.A(n5836_1), .B(n5838), .S0(TM1), .Y(n5839));
NOR2X1   g0300(.A(n5839), .B(n5827), .Y(n871));
INVX1    g0301(.A(CRC_OUT_9_30), .Y(n5841_1));
XOR2X1   g0302(.A(WX1940), .B(TM1), .Y(n5842));
XOR2X1   g0303(.A(n5842), .B(WX2004), .Y(n5843));
INVX1    g0304(.A(WX2068), .Y(n5844));
XOR2X1   g0305(.A(WX2132), .B(n5844), .Y(n5845));
XOR2X1   g0306(.A(n5845), .B(n5843), .Y(n5846_1));
MX2X1    g0307(.A(n5841_1), .B(n5846_1), .S0(n5539), .Y(n5848));
INVX1    g0308(.A(WX487), .Y(n5849));
MX2X1    g0309(.A(n5849), .B(n5552), .S0(n5539), .Y(n5850));
MX2X1    g0310(.A(n5848), .B(n5850), .S0(TM1), .Y(n5851_1));
NOR2X1   g0311(.A(n5851_1), .B(n5827), .Y(n876));
INVX1    g0312(.A(CRC_OUT_9_29), .Y(n5853));
XOR2X1   g0313(.A(WX1942), .B(TM1), .Y(n5854));
XOR2X1   g0314(.A(n5854), .B(WX2006), .Y(n5855));
INVX1    g0315(.A(WX2070), .Y(n5856_1));
XOR2X1   g0316(.A(WX2134), .B(n5856_1), .Y(n5857));
XOR2X1   g0317(.A(n5857), .B(n5855), .Y(n5858));
MX2X1    g0318(.A(n5853), .B(n5858), .S0(n5539), .Y(n5860));
INVX1    g0319(.A(WX489), .Y(n5861_1));
MX2X1    g0320(.A(n5861_1), .B(n5560), .S0(n5539), .Y(n5862));
MX2X1    g0321(.A(n5860), .B(n5862), .S0(TM1), .Y(n5863));
NOR2X1   g0322(.A(n5863), .B(n5827), .Y(n881));
INVX1    g0323(.A(CRC_OUT_9_28), .Y(n5865));
XOR2X1   g0324(.A(WX1944), .B(TM1), .Y(n5866_1));
XOR2X1   g0325(.A(n5866_1), .B(WX2008), .Y(n5867));
INVX1    g0326(.A(WX2072), .Y(n5868));
XOR2X1   g0327(.A(WX2136), .B(n5868), .Y(n5869));
XOR2X1   g0328(.A(n5869), .B(n5867), .Y(n5870));
MX2X1    g0329(.A(n5865), .B(n5870), .S0(n5539), .Y(n5872));
INVX1    g0330(.A(WX491), .Y(n5873));
MX2X1    g0331(.A(n5873), .B(n5568), .S0(n5539), .Y(n5874));
MX2X1    g0332(.A(n5872), .B(n5874), .S0(TM1), .Y(n5875));
NOR2X1   g0333(.A(n5875), .B(n5827), .Y(n886));
INVX1    g0334(.A(CRC_OUT_9_27), .Y(n5877));
XOR2X1   g0335(.A(WX1946), .B(TM1), .Y(n5878));
XOR2X1   g0336(.A(n5878), .B(WX2010), .Y(n5879));
INVX1    g0337(.A(WX2074), .Y(n5880));
XOR2X1   g0338(.A(WX2138), .B(n5880), .Y(n5881_1));
XOR2X1   g0339(.A(n5881_1), .B(n5879), .Y(n5882));
MX2X1    g0340(.A(n5877), .B(n5882), .S0(n5539), .Y(n5884));
INVX1    g0341(.A(WX493), .Y(n5885));
MX2X1    g0342(.A(n5885), .B(n5576_1), .S0(n5539), .Y(n5886_1));
MX2X1    g0343(.A(n5884), .B(n5886_1), .S0(TM1), .Y(n5887));
NOR2X1   g0344(.A(n5887), .B(n5827), .Y(n891));
INVX1    g0345(.A(CRC_OUT_9_26), .Y(n5889));
XOR2X1   g0346(.A(WX1948), .B(TM1), .Y(n5890));
XOR2X1   g0347(.A(n5890), .B(WX2012), .Y(n5891_1));
INVX1    g0348(.A(WX2076), .Y(n5892));
XOR2X1   g0349(.A(WX2140), .B(n5892), .Y(n5893));
XOR2X1   g0350(.A(n5893), .B(n5891_1), .Y(n5894));
MX2X1    g0351(.A(n5889), .B(n5894), .S0(n5539), .Y(n5896_1));
INVX1    g0352(.A(WX495), .Y(n5897));
MX2X1    g0353(.A(n5897), .B(n5584), .S0(n5539), .Y(n5898));
MX2X1    g0354(.A(n5896_1), .B(n5898), .S0(TM1), .Y(n5899));
NOR2X1   g0355(.A(n5899), .B(n5827), .Y(n896));
INVX1    g0356(.A(CRC_OUT_9_25), .Y(n5901_1));
XOR2X1   g0357(.A(WX1950), .B(TM1), .Y(n5902));
XOR2X1   g0358(.A(n5902), .B(WX2014), .Y(n5903));
INVX1    g0359(.A(WX2078), .Y(n5904));
XOR2X1   g0360(.A(WX2142), .B(n5904), .Y(n5905));
XOR2X1   g0361(.A(n5905), .B(n5903), .Y(n5906_1));
MX2X1    g0362(.A(n5901_1), .B(n5906_1), .S0(n5539), .Y(n5908));
INVX1    g0363(.A(WX497), .Y(n5909));
MX2X1    g0364(.A(n5909), .B(n5592), .S0(n5539), .Y(n5910));
MX2X1    g0365(.A(n5908), .B(n5910), .S0(TM1), .Y(n5911_1));
NOR2X1   g0366(.A(n5911_1), .B(n5827), .Y(n901));
INVX1    g0367(.A(CRC_OUT_9_24), .Y(n5913));
XOR2X1   g0368(.A(WX1952), .B(TM1), .Y(n5914));
XOR2X1   g0369(.A(n5914), .B(WX2016), .Y(n5915));
INVX1    g0370(.A(WX2080), .Y(n5916_1));
XOR2X1   g0371(.A(WX2144), .B(n5916_1), .Y(n5917));
XOR2X1   g0372(.A(n5917), .B(n5915), .Y(n5918));
MX2X1    g0373(.A(n5913), .B(n5918), .S0(n5539), .Y(n5920));
INVX1    g0374(.A(WX499), .Y(n5921_1));
MX2X1    g0375(.A(n5921_1), .B(n5600), .S0(n5539), .Y(n5922));
MX2X1    g0376(.A(n5920), .B(n5922), .S0(TM1), .Y(n5923));
NOR2X1   g0377(.A(n5923), .B(n5827), .Y(n906));
INVX1    g0378(.A(CRC_OUT_9_23), .Y(n5925));
XOR2X1   g0379(.A(WX1954), .B(TM1), .Y(n5926_1));
XOR2X1   g0380(.A(n5926_1), .B(WX2018), .Y(n5927));
INVX1    g0381(.A(WX2082), .Y(n5928));
XOR2X1   g0382(.A(WX2146), .B(n5928), .Y(n5929));
XOR2X1   g0383(.A(n5929), .B(n5927), .Y(n5930));
MX2X1    g0384(.A(n5925), .B(n5930), .S0(n5539), .Y(n5932));
INVX1    g0385(.A(WX501), .Y(n5933));
MX2X1    g0386(.A(n5933), .B(n5608), .S0(n5539), .Y(n5934));
MX2X1    g0387(.A(n5932), .B(n5934), .S0(TM1), .Y(n5935));
NOR2X1   g0388(.A(n5935), .B(n5827), .Y(n911));
INVX1    g0389(.A(CRC_OUT_9_22), .Y(n5937));
XOR2X1   g0390(.A(WX1956), .B(TM1), .Y(n5938));
XOR2X1   g0391(.A(n5938), .B(WX2020), .Y(n5939));
INVX1    g0392(.A(WX2084), .Y(n5940));
XOR2X1   g0393(.A(WX2148), .B(n5940), .Y(n5941_1));
XOR2X1   g0394(.A(n5941_1), .B(n5939), .Y(n5942));
MX2X1    g0395(.A(n5937), .B(n5942), .S0(n5539), .Y(n5944));
INVX1    g0396(.A(WX503), .Y(n5945));
MX2X1    g0397(.A(n5945), .B(n5616_1), .S0(n5539), .Y(n5946_1));
MX2X1    g0398(.A(n5944), .B(n5946_1), .S0(TM1), .Y(n5947));
NOR2X1   g0399(.A(n5947), .B(n5827), .Y(n916));
INVX1    g0400(.A(CRC_OUT_9_21), .Y(n5949));
XOR2X1   g0401(.A(WX1958), .B(TM1), .Y(n5950));
XOR2X1   g0402(.A(n5950), .B(WX2022), .Y(n5951_1));
INVX1    g0403(.A(WX2086), .Y(n5952));
XOR2X1   g0404(.A(WX2150), .B(n5952), .Y(n5953));
XOR2X1   g0405(.A(n5953), .B(n5951_1), .Y(n5954));
MX2X1    g0406(.A(n5949), .B(n5954), .S0(n5539), .Y(n5956_1));
INVX1    g0407(.A(WX505), .Y(n5957));
MX2X1    g0408(.A(n5957), .B(n5624), .S0(n5539), .Y(n5958));
MX2X1    g0409(.A(n5956_1), .B(n5958), .S0(TM1), .Y(n5959));
NOR2X1   g0410(.A(n5959), .B(n5827), .Y(n921));
INVX1    g0411(.A(CRC_OUT_9_20), .Y(n5961_1));
XOR2X1   g0412(.A(WX1960), .B(TM1), .Y(n5962));
XOR2X1   g0413(.A(n5962), .B(WX2024), .Y(n5963));
INVX1    g0414(.A(WX2088), .Y(n5964));
XOR2X1   g0415(.A(WX2152), .B(n5964), .Y(n5965));
XOR2X1   g0416(.A(n5965), .B(n5963), .Y(n5966_1));
MX2X1    g0417(.A(n5961_1), .B(n5966_1), .S0(n5539), .Y(n5968));
INVX1    g0418(.A(WX507), .Y(n5969));
MX2X1    g0419(.A(n5969), .B(n5632), .S0(n5539), .Y(n5970));
MX2X1    g0420(.A(n5968), .B(n5970), .S0(TM1), .Y(n5971_1));
NOR2X1   g0421(.A(n5971_1), .B(n5827), .Y(n926));
INVX1    g0422(.A(CRC_OUT_9_19), .Y(n5973));
XOR2X1   g0423(.A(WX1962), .B(TM1), .Y(n5974));
XOR2X1   g0424(.A(n5974), .B(WX2026), .Y(n5975));
INVX1    g0425(.A(WX2090), .Y(n5976_1));
XOR2X1   g0426(.A(WX2154), .B(n5976_1), .Y(n5977));
XOR2X1   g0427(.A(n5977), .B(n5975), .Y(n5978));
MX2X1    g0428(.A(n5973), .B(n5978), .S0(n5539), .Y(n5980));
INVX1    g0429(.A(WX509), .Y(n5981_1));
MX2X1    g0430(.A(n5981_1), .B(n5640), .S0(n5539), .Y(n5982));
MX2X1    g0431(.A(n5980), .B(n5982), .S0(TM1), .Y(n5983));
NOR2X1   g0432(.A(n5983), .B(n5827), .Y(n931));
INVX1    g0433(.A(CRC_OUT_9_18), .Y(n5985));
XOR2X1   g0434(.A(WX1964), .B(TM1), .Y(n5986_1));
XOR2X1   g0435(.A(n5986_1), .B(WX2028), .Y(n5987));
INVX1    g0436(.A(WX2092), .Y(n5988));
XOR2X1   g0437(.A(WX2156), .B(n5988), .Y(n5989));
XOR2X1   g0438(.A(n5989), .B(n5987), .Y(n5990));
MX2X1    g0439(.A(n5985), .B(n5990), .S0(n5539), .Y(n5992));
INVX1    g0440(.A(WX511), .Y(n5993));
MX2X1    g0441(.A(n5993), .B(n5648), .S0(n5539), .Y(n5994));
MX2X1    g0442(.A(n5992), .B(n5994), .S0(TM1), .Y(n5995));
NOR2X1   g0443(.A(n5995), .B(n5827), .Y(n936));
INVX1    g0444(.A(CRC_OUT_9_17), .Y(n5997));
XOR2X1   g0445(.A(WX1966), .B(TM1), .Y(n5998));
XOR2X1   g0446(.A(n5998), .B(WX2030), .Y(n5999));
INVX1    g0447(.A(WX2094), .Y(n6000));
XOR2X1   g0448(.A(WX2158), .B(n6000), .Y(n6001_1));
XOR2X1   g0449(.A(n6001_1), .B(n5999), .Y(n6002));
MX2X1    g0450(.A(n5997), .B(n6002), .S0(n5539), .Y(n6004));
INVX1    g0451(.A(WX513), .Y(n6005));
MX2X1    g0452(.A(n6005), .B(n5656_1), .S0(n5539), .Y(n6006_1));
MX2X1    g0453(.A(n6004), .B(n6006_1), .S0(TM1), .Y(n6007));
NOR2X1   g0454(.A(n6007), .B(n5827), .Y(n941));
INVX1    g0455(.A(CRC_OUT_9_16), .Y(n6009));
XOR2X1   g0456(.A(WX1968), .B(TM1), .Y(n6010));
XOR2X1   g0457(.A(n6010), .B(WX2032), .Y(n6011_1));
INVX1    g0458(.A(WX2096), .Y(n6012));
XOR2X1   g0459(.A(WX2160), .B(n6012), .Y(n6013));
XOR2X1   g0460(.A(n6013), .B(n6011_1), .Y(n6014));
MX2X1    g0461(.A(n6009), .B(n6014), .S0(n5539), .Y(n6016_1));
INVX1    g0462(.A(WX515), .Y(n6017));
MX2X1    g0463(.A(n6017), .B(n5664), .S0(n5539), .Y(n6018));
MX2X1    g0464(.A(n6016_1), .B(n6018), .S0(TM1), .Y(n6019));
NOR2X1   g0465(.A(n6019), .B(n5827), .Y(n946));
INVX1    g0466(.A(CRC_OUT_9_15), .Y(n6021_1));
XOR2X1   g0467(.A(WX1970), .B(TM0), .Y(n6022));
XOR2X1   g0468(.A(n6022), .B(WX2034), .Y(n6023));
INVX1    g0469(.A(WX2098), .Y(n6024));
XOR2X1   g0470(.A(WX2162), .B(n6024), .Y(n6025));
XOR2X1   g0471(.A(n6025), .B(n6023), .Y(n6026_1));
MX2X1    g0472(.A(n6021_1), .B(n6026_1), .S0(n5539), .Y(n6028));
INVX1    g0473(.A(WX517), .Y(n6029));
MX2X1    g0474(.A(n6029), .B(n5672), .S0(n5539), .Y(n6030));
MX2X1    g0475(.A(n6028), .B(n6030), .S0(TM1), .Y(n6031_1));
NOR2X1   g0476(.A(n6031_1), .B(n5827), .Y(n951));
INVX1    g0477(.A(CRC_OUT_9_14), .Y(n6033));
XOR2X1   g0478(.A(WX1972), .B(TM0), .Y(n6034));
XOR2X1   g0479(.A(n6034), .B(WX2036), .Y(n6035));
INVX1    g0480(.A(WX2100), .Y(n6036_1));
XOR2X1   g0481(.A(WX2164), .B(n6036_1), .Y(n6037));
XOR2X1   g0482(.A(n6037), .B(n6035), .Y(n6038));
MX2X1    g0483(.A(n6033), .B(n6038), .S0(n5539), .Y(n6040));
INVX1    g0484(.A(WX519), .Y(n6041_1));
MX2X1    g0485(.A(n6041_1), .B(n5680), .S0(n5539), .Y(n6042));
MX2X1    g0486(.A(n6040), .B(n6042), .S0(TM1), .Y(n6043));
NOR2X1   g0487(.A(n6043), .B(n5827), .Y(n956));
INVX1    g0488(.A(CRC_OUT_9_13), .Y(n6045));
XOR2X1   g0489(.A(WX1974), .B(TM0), .Y(n6046_1));
XOR2X1   g0490(.A(n6046_1), .B(WX2038), .Y(n6047));
INVX1    g0491(.A(WX2102), .Y(n6048));
XOR2X1   g0492(.A(WX2166), .B(n6048), .Y(n6049));
XOR2X1   g0493(.A(n6049), .B(n6047), .Y(n6050));
MX2X1    g0494(.A(n6045), .B(n6050), .S0(n5539), .Y(n6052));
INVX1    g0495(.A(WX521), .Y(n6053));
MX2X1    g0496(.A(n6053), .B(n5688), .S0(n5539), .Y(n6054));
MX2X1    g0497(.A(n6052), .B(n6054), .S0(TM1), .Y(n6055));
NOR2X1   g0498(.A(n6055), .B(n5827), .Y(n961));
INVX1    g0499(.A(CRC_OUT_9_12), .Y(n6057));
XOR2X1   g0500(.A(WX1976), .B(TM0), .Y(n6058));
XOR2X1   g0501(.A(n6058), .B(WX2040), .Y(n6059));
INVX1    g0502(.A(WX2104), .Y(n6060));
XOR2X1   g0503(.A(WX2168), .B(n6060), .Y(n6061_1));
XOR2X1   g0504(.A(n6061_1), .B(n6059), .Y(n6062));
MX2X1    g0505(.A(n6057), .B(n6062), .S0(n5539), .Y(n6064));
INVX1    g0506(.A(WX523), .Y(n6065));
MX2X1    g0507(.A(n6065), .B(n5696_1), .S0(n5539), .Y(n6066_1));
MX2X1    g0508(.A(n6064), .B(n6066_1), .S0(TM1), .Y(n6067));
NOR2X1   g0509(.A(n6067), .B(n5827), .Y(n966));
INVX1    g0510(.A(CRC_OUT_9_11), .Y(n6069));
XOR2X1   g0511(.A(WX1978), .B(TM0), .Y(n6070));
XOR2X1   g0512(.A(n6070), .B(WX2042), .Y(n6071_1));
INVX1    g0513(.A(WX2106), .Y(n6072));
XOR2X1   g0514(.A(WX2170), .B(n6072), .Y(n6073));
XOR2X1   g0515(.A(n6073), .B(n6071_1), .Y(n6074));
MX2X1    g0516(.A(n6069), .B(n6074), .S0(n5539), .Y(n6076_1));
INVX1    g0517(.A(WX525), .Y(n6077));
MX2X1    g0518(.A(n6077), .B(n5704), .S0(n5539), .Y(n6078));
MX2X1    g0519(.A(n6076_1), .B(n6078), .S0(TM1), .Y(n6079));
NOR2X1   g0520(.A(n6079), .B(n5827), .Y(n971));
INVX1    g0521(.A(CRC_OUT_9_10), .Y(n6081_1));
XOR2X1   g0522(.A(WX1980), .B(TM0), .Y(n6082));
XOR2X1   g0523(.A(n6082), .B(WX2044), .Y(n6083));
INVX1    g0524(.A(WX2108), .Y(n6084));
XOR2X1   g0525(.A(WX2172), .B(n6084), .Y(n6085));
XOR2X1   g0526(.A(n6085), .B(n6083), .Y(n6086_1));
MX2X1    g0527(.A(n6081_1), .B(n6086_1), .S0(n5539), .Y(n6088));
INVX1    g0528(.A(WX527), .Y(n6089));
MX2X1    g0529(.A(n6089), .B(n5712), .S0(n5539), .Y(n6090));
MX2X1    g0530(.A(n6088), .B(n6090), .S0(TM1), .Y(n6091_1));
NOR2X1   g0531(.A(n6091_1), .B(n5827), .Y(n976));
INVX1    g0532(.A(CRC_OUT_9_9), .Y(n6093));
XOR2X1   g0533(.A(WX1982), .B(TM0), .Y(n6094));
XOR2X1   g0534(.A(n6094), .B(WX2046), .Y(n6095));
INVX1    g0535(.A(WX2110), .Y(n6096_1));
XOR2X1   g0536(.A(WX2174), .B(n6096_1), .Y(n6097));
XOR2X1   g0537(.A(n6097), .B(n6095), .Y(n6098));
MX2X1    g0538(.A(n6093), .B(n6098), .S0(n5539), .Y(n6100));
INVX1    g0539(.A(WX529), .Y(n6101_1));
MX2X1    g0540(.A(n6101_1), .B(n5720), .S0(n5539), .Y(n6102));
MX2X1    g0541(.A(n6100), .B(n6102), .S0(TM1), .Y(n6103));
NOR2X1   g0542(.A(n6103), .B(n5827), .Y(n981));
INVX1    g0543(.A(CRC_OUT_9_8), .Y(n6105));
XOR2X1   g0544(.A(WX1984), .B(TM0), .Y(n6106_1));
XOR2X1   g0545(.A(n6106_1), .B(WX2048), .Y(n6107));
INVX1    g0546(.A(WX2112), .Y(n6108));
XOR2X1   g0547(.A(WX2176), .B(n6108), .Y(n6109));
XOR2X1   g0548(.A(n6109), .B(n6107), .Y(n6110));
MX2X1    g0549(.A(n6105), .B(n6110), .S0(n5539), .Y(n6112));
INVX1    g0550(.A(WX531), .Y(n6113));
MX2X1    g0551(.A(n6113), .B(n5728), .S0(n5539), .Y(n6114));
MX2X1    g0552(.A(n6112), .B(n6114), .S0(TM1), .Y(n6115));
NOR2X1   g0553(.A(n6115), .B(n5827), .Y(n986));
INVX1    g0554(.A(CRC_OUT_9_7), .Y(n6117));
XOR2X1   g0555(.A(WX1986), .B(TM0), .Y(n6118));
XOR2X1   g0556(.A(n6118), .B(WX2050), .Y(n6119));
INVX1    g0557(.A(WX2114), .Y(n6120));
XOR2X1   g0558(.A(WX2178), .B(n6120), .Y(n6121_1));
XOR2X1   g0559(.A(n6121_1), .B(n6119), .Y(n6122));
MX2X1    g0560(.A(n6117), .B(n6122), .S0(n5539), .Y(n6124));
INVX1    g0561(.A(WX533), .Y(n6125));
MX2X1    g0562(.A(n6125), .B(n5736_1), .S0(n5539), .Y(n6126_1));
MX2X1    g0563(.A(n6124), .B(n6126_1), .S0(TM1), .Y(n6127));
NOR2X1   g0564(.A(n6127), .B(n5827), .Y(n991));
INVX1    g0565(.A(CRC_OUT_9_6), .Y(n6129));
XOR2X1   g0566(.A(WX1988), .B(TM0), .Y(n6130));
XOR2X1   g0567(.A(n6130), .B(WX2052), .Y(n6131_1));
INVX1    g0568(.A(WX2116), .Y(n6132));
XOR2X1   g0569(.A(WX2180), .B(n6132), .Y(n6133));
XOR2X1   g0570(.A(n6133), .B(n6131_1), .Y(n6134));
MX2X1    g0571(.A(n6129), .B(n6134), .S0(n5539), .Y(n6136_1));
INVX1    g0572(.A(WX535), .Y(n6137));
MX2X1    g0573(.A(n6137), .B(n5744), .S0(n5539), .Y(n6138));
MX2X1    g0574(.A(n6136_1), .B(n6138), .S0(TM1), .Y(n6139));
NOR2X1   g0575(.A(n6139), .B(n5827), .Y(n996));
INVX1    g0576(.A(CRC_OUT_9_5), .Y(n6141_1));
XOR2X1   g0577(.A(WX1990), .B(TM0), .Y(n6142));
XOR2X1   g0578(.A(n6142), .B(WX2054), .Y(n6143));
INVX1    g0579(.A(WX2118), .Y(n6144));
XOR2X1   g0580(.A(WX2182), .B(n6144), .Y(n6145));
XOR2X1   g0581(.A(n6145), .B(n6143), .Y(n6146_1));
MX2X1    g0582(.A(n6141_1), .B(n6146_1), .S0(n5539), .Y(n6148));
INVX1    g0583(.A(WX537), .Y(n6149));
MX2X1    g0584(.A(n6149), .B(n5752), .S0(n5539), .Y(n6150));
MX2X1    g0585(.A(n6148), .B(n6150), .S0(TM1), .Y(n6151_1));
NOR2X1   g0586(.A(n6151_1), .B(n5827), .Y(n1001));
INVX1    g0587(.A(CRC_OUT_9_4), .Y(n6153));
XOR2X1   g0588(.A(WX1992), .B(TM0), .Y(n6154));
XOR2X1   g0589(.A(n6154), .B(WX2056), .Y(n6155_1));
INVX1    g0590(.A(WX2120), .Y(n6156));
XOR2X1   g0591(.A(WX2184), .B(n6156), .Y(n6157));
XOR2X1   g0592(.A(n6157), .B(n6155_1), .Y(n6158));
MX2X1    g0593(.A(n6153), .B(n6158), .S0(n5539), .Y(n6160));
INVX1    g0594(.A(WX539), .Y(n6161));
MX2X1    g0595(.A(n6161), .B(n5760), .S0(n5539), .Y(n6162));
MX2X1    g0596(.A(n6160), .B(n6162), .S0(TM1), .Y(n6163_1));
NOR2X1   g0597(.A(n6163_1), .B(n5827), .Y(n1006));
INVX1    g0598(.A(CRC_OUT_9_3), .Y(n6165));
XOR2X1   g0599(.A(WX1994), .B(TM0), .Y(n6166));
XOR2X1   g0600(.A(n6166), .B(WX2058), .Y(n6167_1));
INVX1    g0601(.A(WX2122), .Y(n6168));
XOR2X1   g0602(.A(WX2186), .B(n6168), .Y(n6169));
XOR2X1   g0603(.A(n6169), .B(n6167_1), .Y(n6170));
MX2X1    g0604(.A(n6165), .B(n6170), .S0(n5539), .Y(n6172));
INVX1    g0605(.A(WX541), .Y(n6173));
MX2X1    g0606(.A(n6173), .B(n5768), .S0(n5539), .Y(n6174));
MX2X1    g0607(.A(n6172), .B(n6174), .S0(TM1), .Y(n6175_1));
NOR2X1   g0608(.A(n6175_1), .B(n5827), .Y(n1011));
INVX1    g0609(.A(CRC_OUT_9_2), .Y(n6177));
XOR2X1   g0610(.A(WX1996), .B(TM0), .Y(n6178));
XOR2X1   g0611(.A(n6178), .B(WX2060), .Y(n6179_1));
INVX1    g0612(.A(WX2124), .Y(n6180));
XOR2X1   g0613(.A(WX2188), .B(n6180), .Y(n6181));
XOR2X1   g0614(.A(n6181), .B(n6179_1), .Y(n6182));
MX2X1    g0615(.A(n6177), .B(n6182), .S0(n5539), .Y(n6184));
INVX1    g0616(.A(WX543), .Y(n6185));
MX2X1    g0617(.A(n6185), .B(n5776_1), .S0(n5539), .Y(n6186));
MX2X1    g0618(.A(n6184), .B(n6186), .S0(TM1), .Y(n6187_1));
NOR2X1   g0619(.A(n6187_1), .B(n5827), .Y(n1016));
INVX1    g0620(.A(CRC_OUT_9_1), .Y(n6189));
XOR2X1   g0621(.A(WX1998), .B(TM0), .Y(n6190));
XOR2X1   g0622(.A(n6190), .B(WX2062), .Y(n6191_1));
INVX1    g0623(.A(WX2126), .Y(n6192));
XOR2X1   g0624(.A(WX2190), .B(n6192), .Y(n6193));
XOR2X1   g0625(.A(n6193), .B(n6191_1), .Y(n6194));
MX2X1    g0626(.A(n6189), .B(n6194), .S0(n5539), .Y(n6196));
INVX1    g0627(.A(WX545), .Y(n6197));
MX2X1    g0628(.A(n6197), .B(n5784), .S0(n5539), .Y(n6198));
MX2X1    g0629(.A(n6196), .B(n6198), .S0(TM1), .Y(n6199_1));
NOR2X1   g0630(.A(n6199_1), .B(n5827), .Y(n1021));
INVX1    g0631(.A(CRC_OUT_9_0), .Y(n6201));
XOR2X1   g0632(.A(WX2000), .B(TM0), .Y(n6202));
XOR2X1   g0633(.A(n6202), .B(WX2064), .Y(n6203_1));
INVX1    g0634(.A(WX2128), .Y(n6204));
XOR2X1   g0635(.A(WX2192), .B(n6204), .Y(n6205));
XOR2X1   g0636(.A(n6205), .B(n6203_1), .Y(n6206));
MX2X1    g0637(.A(n6201), .B(n6206), .S0(n5539), .Y(n6208));
INVX1    g0638(.A(WX547), .Y(n6209));
MX2X1    g0639(.A(n6209), .B(n5792), .S0(n5539), .Y(n6210));
MX2X1    g0640(.A(n6208), .B(n6210), .S0(TM1), .Y(n6211_1));
NOR2X1   g0641(.A(n6211_1), .B(n5827), .Y(n1026));
AND2X1   g0642(.A(WX645), .B(RESET), .Y(n1031));
AND2X1   g0643(.A(WX647), .B(RESET), .Y(n1036));
AND2X1   g0644(.A(WX649), .B(RESET), .Y(n1041));
AND2X1   g0645(.A(WX651), .B(RESET), .Y(n1046));
AND2X1   g0646(.A(WX653), .B(RESET), .Y(n1051));
AND2X1   g0647(.A(WX655), .B(RESET), .Y(n1056));
AND2X1   g0648(.A(WX657), .B(RESET), .Y(n1061));
AND2X1   g0649(.A(WX659), .B(RESET), .Y(n1066));
AND2X1   g0650(.A(WX661), .B(RESET), .Y(n1071));
AND2X1   g0651(.A(WX663), .B(RESET), .Y(n1076));
AND2X1   g0652(.A(WX665), .B(RESET), .Y(n1081));
AND2X1   g0653(.A(WX667), .B(RESET), .Y(n1086));
AND2X1   g0654(.A(WX669), .B(RESET), .Y(n1091));
AND2X1   g0655(.A(WX671), .B(RESET), .Y(n1096));
AND2X1   g0656(.A(WX673), .B(RESET), .Y(n1101));
AND2X1   g0657(.A(WX675), .B(RESET), .Y(n1106));
AND2X1   g0658(.A(WX677), .B(RESET), .Y(n1111));
AND2X1   g0659(.A(WX679), .B(RESET), .Y(n1116));
AND2X1   g0660(.A(WX681), .B(RESET), .Y(n1121));
AND2X1   g0661(.A(WX683), .B(RESET), .Y(n1126));
AND2X1   g0662(.A(WX685), .B(RESET), .Y(n1131));
AND2X1   g0663(.A(WX687), .B(RESET), .Y(n1136));
AND2X1   g0664(.A(WX689), .B(RESET), .Y(n1141));
AND2X1   g0665(.A(WX691), .B(RESET), .Y(n1146));
AND2X1   g0666(.A(WX693), .B(RESET), .Y(n1151));
AND2X1   g0667(.A(WX695), .B(RESET), .Y(n1156));
AND2X1   g0668(.A(WX697), .B(RESET), .Y(n1161));
AND2X1   g0669(.A(WX699), .B(RESET), .Y(n1166));
AND2X1   g0670(.A(WX701), .B(RESET), .Y(n1171));
AND2X1   g0671(.A(WX703), .B(RESET), .Y(n1176));
AND2X1   g0672(.A(WX705), .B(RESET), .Y(n1181));
AND2X1   g0673(.A(WX707), .B(RESET), .Y(n1186));
AND2X1   g0674(.A(WX709), .B(RESET), .Y(n1191));
AND2X1   g0675(.A(WX711), .B(RESET), .Y(n1196));
AND2X1   g0676(.A(WX713), .B(RESET), .Y(n1201));
AND2X1   g0677(.A(WX715), .B(RESET), .Y(n1206));
AND2X1   g0678(.A(WX717), .B(RESET), .Y(n1211));
AND2X1   g0679(.A(WX719), .B(RESET), .Y(n1216));
AND2X1   g0680(.A(WX721), .B(RESET), .Y(n1221));
AND2X1   g0681(.A(WX723), .B(RESET), .Y(n1226));
AND2X1   g0682(.A(WX725), .B(RESET), .Y(n1231));
AND2X1   g0683(.A(WX727), .B(RESET), .Y(n1236));
AND2X1   g0684(.A(WX729), .B(RESET), .Y(n1241));
AND2X1   g0685(.A(WX731), .B(RESET), .Y(n1246));
AND2X1   g0686(.A(WX733), .B(RESET), .Y(n1251));
AND2X1   g0687(.A(WX735), .B(RESET), .Y(n1256));
AND2X1   g0688(.A(WX737), .B(RESET), .Y(n1261));
AND2X1   g0689(.A(WX739), .B(RESET), .Y(n1266));
AND2X1   g0690(.A(WX741), .B(RESET), .Y(n1271));
AND2X1   g0691(.A(WX743), .B(RESET), .Y(n1276));
AND2X1   g0692(.A(WX745), .B(RESET), .Y(n1281));
AND2X1   g0693(.A(WX747), .B(RESET), .Y(n1286));
AND2X1   g0694(.A(WX749), .B(RESET), .Y(n1291));
AND2X1   g0695(.A(WX751), .B(RESET), .Y(n1296));
AND2X1   g0696(.A(WX753), .B(RESET), .Y(n1301));
AND2X1   g0697(.A(WX755), .B(RESET), .Y(n1306));
AND2X1   g0698(.A(WX757), .B(RESET), .Y(n1311));
AND2X1   g0699(.A(WX759), .B(RESET), .Y(n1316));
AND2X1   g0700(.A(WX761), .B(RESET), .Y(n1321));
AND2X1   g0701(.A(WX763), .B(RESET), .Y(n1326));
AND2X1   g0702(.A(WX765), .B(RESET), .Y(n1331));
AND2X1   g0703(.A(WX767), .B(RESET), .Y(n1336));
AND2X1   g0704(.A(WX769), .B(RESET), .Y(n1341));
AND2X1   g0705(.A(WX771), .B(RESET), .Y(n1346));
AND2X1   g0706(.A(WX773), .B(RESET), .Y(n1351));
AND2X1   g0707(.A(WX775), .B(RESET), .Y(n1356));
AND2X1   g0708(.A(WX777), .B(RESET), .Y(n1361));
AND2X1   g0709(.A(WX779), .B(RESET), .Y(n1366));
AND2X1   g0710(.A(WX781), .B(RESET), .Y(n1371));
AND2X1   g0711(.A(WX783), .B(RESET), .Y(n1376));
AND2X1   g0712(.A(WX785), .B(RESET), .Y(n1381));
AND2X1   g0713(.A(WX787), .B(RESET), .Y(n1386));
AND2X1   g0714(.A(WX789), .B(RESET), .Y(n1391));
AND2X1   g0715(.A(WX791), .B(RESET), .Y(n1396));
AND2X1   g0716(.A(WX793), .B(RESET), .Y(n1401));
AND2X1   g0717(.A(WX795), .B(RESET), .Y(n1406));
AND2X1   g0718(.A(WX797), .B(RESET), .Y(n1411));
AND2X1   g0719(.A(WX799), .B(RESET), .Y(n1416));
AND2X1   g0720(.A(WX801), .B(RESET), .Y(n1421));
AND2X1   g0721(.A(WX803), .B(RESET), .Y(n1426));
AND2X1   g0722(.A(WX805), .B(RESET), .Y(n1431));
AND2X1   g0723(.A(WX807), .B(RESET), .Y(n1436));
AND2X1   g0724(.A(WX809), .B(RESET), .Y(n1441));
AND2X1   g0725(.A(WX811), .B(RESET), .Y(n1446));
AND2X1   g0726(.A(WX813), .B(RESET), .Y(n1451));
AND2X1   g0727(.A(WX815), .B(RESET), .Y(n1456));
AND2X1   g0728(.A(WX817), .B(RESET), .Y(n1461));
AND2X1   g0729(.A(WX819), .B(RESET), .Y(n1466));
AND2X1   g0730(.A(WX821), .B(RESET), .Y(n1471));
AND2X1   g0731(.A(WX823), .B(RESET), .Y(n1476));
AND2X1   g0732(.A(WX825), .B(RESET), .Y(n1481));
AND2X1   g0733(.A(WX827), .B(RESET), .Y(n1486));
AND2X1   g0734(.A(WX829), .B(RESET), .Y(n1491));
AND2X1   g0735(.A(WX831), .B(RESET), .Y(n1496));
AND2X1   g0736(.A(WX833), .B(RESET), .Y(n1501));
AND2X1   g0737(.A(WX835), .B(RESET), .Y(n1506));
XOR2X1   g0738(.A(CRC_OUT_9_31), .B(WX899), .Y(n6309_1));
NOR2X1   g0739(.A(n6309_1), .B(n5827), .Y(CRC_OUT_9_0));
XOR2X1   g0740(.A(CRC_OUT_9_0), .B(WX897), .Y(n6311));
NOR2X1   g0741(.A(n6311), .B(n5827), .Y(CRC_OUT_9_1));
XOR2X1   g0742(.A(CRC_OUT_9_1), .B(WX895), .Y(n6313));
NOR2X1   g0743(.A(n6313), .B(n5827), .Y(CRC_OUT_9_2));
XOR2X1   g0744(.A(CRC_OUT_9_2), .B(WX893), .Y(n6315));
NOR2X1   g0745(.A(n6315), .B(n5827), .Y(CRC_OUT_9_3));
XOR2X1   g0746(.A(CRC_OUT_9_31), .B(WX891), .Y(n6317));
XOR2X1   g0747(.A(n6317), .B(CRC_OUT_9_3), .Y(n6318));
NOR2X1   g0748(.A(n6318), .B(n5827), .Y(CRC_OUT_9_4));
XOR2X1   g0749(.A(CRC_OUT_9_4), .B(WX889), .Y(n6320));
NOR2X1   g0750(.A(n6320), .B(n5827), .Y(CRC_OUT_9_5));
XOR2X1   g0751(.A(CRC_OUT_9_5), .B(WX887), .Y(n6322));
NOR2X1   g0752(.A(n6322), .B(n5827), .Y(CRC_OUT_9_6));
XOR2X1   g0753(.A(CRC_OUT_9_6), .B(WX885), .Y(n6324_1));
NOR2X1   g0754(.A(n6324_1), .B(n5827), .Y(CRC_OUT_9_7));
XOR2X1   g0755(.A(CRC_OUT_9_7), .B(WX883), .Y(n6326));
NOR2X1   g0756(.A(n6326), .B(n5827), .Y(CRC_OUT_9_8));
XOR2X1   g0757(.A(CRC_OUT_9_8), .B(WX881), .Y(n6328));
NOR2X1   g0758(.A(n6328), .B(n5827), .Y(CRC_OUT_9_9));
XOR2X1   g0759(.A(CRC_OUT_9_9), .B(WX879), .Y(n6330));
NOR2X1   g0760(.A(n6330), .B(n5827), .Y(CRC_OUT_9_10));
XOR2X1   g0761(.A(CRC_OUT_9_31), .B(WX877), .Y(n6332));
XOR2X1   g0762(.A(n6332), .B(CRC_OUT_9_10), .Y(n6333));
NOR2X1   g0763(.A(n6333), .B(n5827), .Y(CRC_OUT_9_11));
XOR2X1   g0764(.A(CRC_OUT_9_11), .B(WX875), .Y(n6335));
NOR2X1   g0765(.A(n6335), .B(n5827), .Y(CRC_OUT_9_12));
XOR2X1   g0766(.A(CRC_OUT_9_12), .B(WX873), .Y(n6337));
NOR2X1   g0767(.A(n6337), .B(n5827), .Y(CRC_OUT_9_13));
XOR2X1   g0768(.A(CRC_OUT_9_13), .B(WX871), .Y(n6339_1));
NOR2X1   g0769(.A(n6339_1), .B(n5827), .Y(CRC_OUT_9_14));
XOR2X1   g0770(.A(CRC_OUT_9_14), .B(WX869), .Y(n6341));
NOR2X1   g0771(.A(n6341), .B(n5827), .Y(CRC_OUT_9_15));
XOR2X1   g0772(.A(CRC_OUT_9_31), .B(WX867), .Y(n6343));
XOR2X1   g0773(.A(n6343), .B(CRC_OUT_9_15), .Y(n6344_1));
NOR2X1   g0774(.A(n6344_1), .B(n5827), .Y(CRC_OUT_9_16));
XOR2X1   g0775(.A(CRC_OUT_9_16), .B(WX865), .Y(n6346));
NOR2X1   g0776(.A(n6346), .B(n5827), .Y(CRC_OUT_9_17));
XOR2X1   g0777(.A(CRC_OUT_9_17), .B(WX863), .Y(n6348));
NOR2X1   g0778(.A(n6348), .B(n5827), .Y(CRC_OUT_9_18));
XOR2X1   g0779(.A(CRC_OUT_9_18), .B(WX861), .Y(n6350));
NOR2X1   g0780(.A(n6350), .B(n5827), .Y(CRC_OUT_9_19));
XOR2X1   g0781(.A(CRC_OUT_9_19), .B(WX859), .Y(n6352));
NOR2X1   g0782(.A(n6352), .B(n5827), .Y(CRC_OUT_9_20));
XOR2X1   g0783(.A(CRC_OUT_9_20), .B(WX857), .Y(n6354_1));
NOR2X1   g0784(.A(n6354_1), .B(n5827), .Y(CRC_OUT_9_21));
XOR2X1   g0785(.A(CRC_OUT_9_21), .B(WX855), .Y(n6356));
NOR2X1   g0786(.A(n6356), .B(n5827), .Y(CRC_OUT_9_22));
XOR2X1   g0787(.A(CRC_OUT_9_22), .B(WX853), .Y(n6358));
NOR2X1   g0788(.A(n6358), .B(n5827), .Y(CRC_OUT_9_23));
XOR2X1   g0789(.A(CRC_OUT_9_23), .B(WX851), .Y(n6360));
NOR2X1   g0790(.A(n6360), .B(n5827), .Y(CRC_OUT_9_24));
XOR2X1   g0791(.A(CRC_OUT_9_24), .B(WX849), .Y(n6362));
NOR2X1   g0792(.A(n6362), .B(n5827), .Y(CRC_OUT_9_25));
XOR2X1   g0793(.A(CRC_OUT_9_25), .B(WX847), .Y(n6364_1));
NOR2X1   g0794(.A(n6364_1), .B(n5827), .Y(CRC_OUT_9_26));
XOR2X1   g0795(.A(CRC_OUT_9_26), .B(WX845), .Y(n6366));
NOR2X1   g0796(.A(n6366), .B(n5827), .Y(CRC_OUT_9_27));
XOR2X1   g0797(.A(CRC_OUT_9_27), .B(WX843), .Y(n6368));
NOR2X1   g0798(.A(n6368), .B(n5827), .Y(CRC_OUT_9_28));
XOR2X1   g0799(.A(CRC_OUT_9_28), .B(WX841), .Y(n6370));
NOR2X1   g0800(.A(n6370), .B(n5827), .Y(CRC_OUT_9_29));
XOR2X1   g0801(.A(CRC_OUT_9_29), .B(WX839), .Y(n6372));
NOR2X1   g0802(.A(n6372), .B(n5827), .Y(CRC_OUT_9_30));
XOR2X1   g0803(.A(CRC_OUT_9_30), .B(WX837), .Y(n6374_1));
NOR2X1   g0804(.A(n6374_1), .B(n5827), .Y(CRC_OUT_9_31));
AND2X1   g0805(.A(WX1780), .B(RESET), .Y(n1639));
AND2X1   g0806(.A(WX1782), .B(RESET), .Y(n1644));
AND2X1   g0807(.A(WX1784), .B(RESET), .Y(n1649));
AND2X1   g0808(.A(WX1786), .B(RESET), .Y(n1654));
AND2X1   g0809(.A(WX1788), .B(RESET), .Y(n1659));
AND2X1   g0810(.A(WX1790), .B(RESET), .Y(n1664));
AND2X1   g0811(.A(WX1792), .B(RESET), .Y(n1669));
AND2X1   g0812(.A(WX1794), .B(RESET), .Y(n1674));
AND2X1   g0813(.A(WX1796), .B(RESET), .Y(n1679));
AND2X1   g0814(.A(WX1798), .B(RESET), .Y(n1684));
AND2X1   g0815(.A(WX1800), .B(RESET), .Y(n1689));
AND2X1   g0816(.A(WX1802), .B(RESET), .Y(n1694));
AND2X1   g0817(.A(WX1804), .B(RESET), .Y(n1699));
AND2X1   g0818(.A(WX1806), .B(RESET), .Y(n1704));
AND2X1   g0819(.A(WX1808), .B(RESET), .Y(n1709));
AND2X1   g0820(.A(WX1810), .B(RESET), .Y(n1714));
AND2X1   g0821(.A(WX1812), .B(RESET), .Y(n1719));
AND2X1   g0822(.A(WX1814), .B(RESET), .Y(n1724));
AND2X1   g0823(.A(WX1816), .B(RESET), .Y(n1729));
AND2X1   g0824(.A(WX1818), .B(RESET), .Y(n1734));
AND2X1   g0825(.A(WX1820), .B(RESET), .Y(n1739));
AND2X1   g0826(.A(WX1822), .B(RESET), .Y(n1744));
AND2X1   g0827(.A(WX1824), .B(RESET), .Y(n1749));
AND2X1   g0828(.A(WX1826), .B(RESET), .Y(n1754));
AND2X1   g0829(.A(WX1828), .B(RESET), .Y(n1759));
AND2X1   g0830(.A(WX1830), .B(RESET), .Y(n1764));
AND2X1   g0831(.A(WX1832), .B(RESET), .Y(n1769));
AND2X1   g0832(.A(WX1834), .B(RESET), .Y(n1774));
AND2X1   g0833(.A(WX1836), .B(RESET), .Y(n1779));
AND2X1   g0834(.A(WX1838), .B(RESET), .Y(n1784));
AND2X1   g0835(.A(WX1840), .B(RESET), .Y(n1789));
NOR2X1   g0836(.A(WX1778), .B(n5827), .Y(n1794));
INVX1    g0837(.A(CRC_OUT_8_31), .Y(n6408));
XOR2X1   g0838(.A(WX3231), .B(TM1), .Y(n6409_1));
XOR2X1   g0839(.A(n6409_1), .B(WX3295), .Y(n6410));
INVX1    g0840(.A(WX3359), .Y(n6411));
XOR2X1   g0841(.A(WX3423), .B(n6411), .Y(n6412));
XOR2X1   g0842(.A(n6412), .B(n6410), .Y(n6413));
MX2X1    g0843(.A(n6408), .B(n6413), .S0(n5539), .Y(n6415));
INVX1    g0844(.A(WX1778), .Y(n6416));
MX2X1    g0845(.A(n6416), .B(n5834), .S0(n5539), .Y(n6417));
MX2X1    g0846(.A(n6415), .B(n6417), .S0(TM1), .Y(n6418));
NOR2X1   g0847(.A(n6418), .B(n5827), .Y(n1799));
INVX1    g0848(.A(CRC_OUT_8_30), .Y(n6420));
XOR2X1   g0849(.A(WX3233), .B(TM1), .Y(n6421));
XOR2X1   g0850(.A(n6421), .B(WX3297), .Y(n6422));
INVX1    g0851(.A(WX3361), .Y(n6423));
XOR2X1   g0852(.A(WX3425), .B(n6423), .Y(n6424_1));
XOR2X1   g0853(.A(n6424_1), .B(n6422), .Y(n6425));
MX2X1    g0854(.A(n6420), .B(n6425), .S0(n5539), .Y(n6427));
INVX1    g0855(.A(WX1780), .Y(n6428));
MX2X1    g0856(.A(n6428), .B(n5846_1), .S0(n5539), .Y(n6429_1));
MX2X1    g0857(.A(n6427), .B(n6429_1), .S0(TM1), .Y(n6430));
NOR2X1   g0858(.A(n6430), .B(n5827), .Y(n1804));
INVX1    g0859(.A(CRC_OUT_8_29), .Y(n6432));
XOR2X1   g0860(.A(WX3235), .B(TM1), .Y(n6433));
XOR2X1   g0861(.A(n6433), .B(WX3299), .Y(n6434_1));
INVX1    g0862(.A(WX3363), .Y(n6435));
XOR2X1   g0863(.A(WX3427), .B(n6435), .Y(n6436));
XOR2X1   g0864(.A(n6436), .B(n6434_1), .Y(n6437));
MX2X1    g0865(.A(n6432), .B(n6437), .S0(n5539), .Y(n6439_1));
INVX1    g0866(.A(WX1782), .Y(n6440));
MX2X1    g0867(.A(n6440), .B(n5858), .S0(n5539), .Y(n6441));
MX2X1    g0868(.A(n6439_1), .B(n6441), .S0(TM1), .Y(n6442));
NOR2X1   g0869(.A(n6442), .B(n5827), .Y(n1809));
INVX1    g0870(.A(CRC_OUT_8_28), .Y(n6444_1));
XOR2X1   g0871(.A(WX3237), .B(TM1), .Y(n6445));
XOR2X1   g0872(.A(n6445), .B(WX3301), .Y(n6446));
INVX1    g0873(.A(WX3365), .Y(n6447));
XOR2X1   g0874(.A(WX3429), .B(n6447), .Y(n6448));
XOR2X1   g0875(.A(n6448), .B(n6446), .Y(n6449_1));
MX2X1    g0876(.A(n6444_1), .B(n6449_1), .S0(n5539), .Y(n6451));
INVX1    g0877(.A(WX1784), .Y(n6452));
MX2X1    g0878(.A(n6452), .B(n5870), .S0(n5539), .Y(n6453));
MX2X1    g0879(.A(n6451), .B(n6453), .S0(TM1), .Y(n6454_1));
NOR2X1   g0880(.A(n6454_1), .B(n5827), .Y(n1814));
INVX1    g0881(.A(CRC_OUT_8_27), .Y(n6456));
XOR2X1   g0882(.A(WX3239), .B(TM1), .Y(n6457));
XOR2X1   g0883(.A(n6457), .B(WX3303), .Y(n6458));
INVX1    g0884(.A(WX3367), .Y(n6459_1));
XOR2X1   g0885(.A(WX3431), .B(n6459_1), .Y(n6460));
XOR2X1   g0886(.A(n6460), .B(n6458), .Y(n6461));
MX2X1    g0887(.A(n6456), .B(n6461), .S0(n5539), .Y(n6463));
INVX1    g0888(.A(WX1786), .Y(n6464_1));
MX2X1    g0889(.A(n6464_1), .B(n5882), .S0(n5539), .Y(n6465));
MX2X1    g0890(.A(n6463), .B(n6465), .S0(TM1), .Y(n6466));
NOR2X1   g0891(.A(n6466), .B(n5827), .Y(n1819));
INVX1    g0892(.A(CRC_OUT_8_26), .Y(n6468));
XOR2X1   g0893(.A(WX3241), .B(TM1), .Y(n6469_1));
XOR2X1   g0894(.A(n6469_1), .B(WX3305), .Y(n6470));
INVX1    g0895(.A(WX3369), .Y(n6471));
XOR2X1   g0896(.A(WX3433), .B(n6471), .Y(n6472));
XOR2X1   g0897(.A(n6472), .B(n6470), .Y(n6473));
MX2X1    g0898(.A(n6468), .B(n6473), .S0(n5539), .Y(n6475));
INVX1    g0899(.A(WX1788), .Y(n6476));
MX2X1    g0900(.A(n6476), .B(n5894), .S0(n5539), .Y(n6477));
MX2X1    g0901(.A(n6475), .B(n6477), .S0(TM1), .Y(n6478));
NOR2X1   g0902(.A(n6478), .B(n5827), .Y(n1824));
INVX1    g0903(.A(CRC_OUT_8_25), .Y(n6480));
XOR2X1   g0904(.A(WX3243), .B(TM1), .Y(n6481));
XOR2X1   g0905(.A(n6481), .B(WX3307), .Y(n6482));
INVX1    g0906(.A(WX3371), .Y(n6483));
XOR2X1   g0907(.A(WX3435), .B(n6483), .Y(n6484_1));
XOR2X1   g0908(.A(n6484_1), .B(n6482), .Y(n6485));
MX2X1    g0909(.A(n6480), .B(n6485), .S0(n5539), .Y(n6487));
INVX1    g0910(.A(WX1790), .Y(n6488));
MX2X1    g0911(.A(n6488), .B(n5906_1), .S0(n5539), .Y(n6489_1));
MX2X1    g0912(.A(n6487), .B(n6489_1), .S0(TM1), .Y(n6490));
NOR2X1   g0913(.A(n6490), .B(n5827), .Y(n1829));
INVX1    g0914(.A(CRC_OUT_8_24), .Y(n6492));
XOR2X1   g0915(.A(WX3245), .B(TM1), .Y(n6493));
XOR2X1   g0916(.A(n6493), .B(WX3309), .Y(n6494_1));
INVX1    g0917(.A(WX3373), .Y(n6495));
XOR2X1   g0918(.A(WX3437), .B(n6495), .Y(n6496));
XOR2X1   g0919(.A(n6496), .B(n6494_1), .Y(n6497));
MX2X1    g0920(.A(n6492), .B(n6497), .S0(n5539), .Y(n6499_1));
INVX1    g0921(.A(WX1792), .Y(n6500));
MX2X1    g0922(.A(n6500), .B(n5918), .S0(n5539), .Y(n6501));
MX2X1    g0923(.A(n6499_1), .B(n6501), .S0(TM1), .Y(n6502));
NOR2X1   g0924(.A(n6502), .B(n5827), .Y(n1834));
INVX1    g0925(.A(CRC_OUT_8_23), .Y(n6504_1));
XOR2X1   g0926(.A(WX3247), .B(TM1), .Y(n6505));
XOR2X1   g0927(.A(n6505), .B(WX3311), .Y(n6506));
INVX1    g0928(.A(WX3375), .Y(n6507));
XOR2X1   g0929(.A(WX3439), .B(n6507), .Y(n6508));
XOR2X1   g0930(.A(n6508), .B(n6506), .Y(n6509_1));
MX2X1    g0931(.A(n6504_1), .B(n6509_1), .S0(n5539), .Y(n6511));
INVX1    g0932(.A(WX1794), .Y(n6512));
MX2X1    g0933(.A(n6512), .B(n5930), .S0(n5539), .Y(n6513));
MX2X1    g0934(.A(n6511), .B(n6513), .S0(TM1), .Y(n6514_1));
NOR2X1   g0935(.A(n6514_1), .B(n5827), .Y(n1839));
INVX1    g0936(.A(CRC_OUT_8_22), .Y(n6516));
XOR2X1   g0937(.A(WX3249), .B(TM1), .Y(n6517));
XOR2X1   g0938(.A(n6517), .B(WX3313), .Y(n6518));
INVX1    g0939(.A(WX3377), .Y(n6519_1));
XOR2X1   g0940(.A(WX3441), .B(n6519_1), .Y(n6520));
XOR2X1   g0941(.A(n6520), .B(n6518), .Y(n6521));
MX2X1    g0942(.A(n6516), .B(n6521), .S0(n5539), .Y(n6523));
INVX1    g0943(.A(WX1796), .Y(n6524_1));
MX2X1    g0944(.A(n6524_1), .B(n5942), .S0(n5539), .Y(n6525));
MX2X1    g0945(.A(n6523), .B(n6525), .S0(TM1), .Y(n6526));
NOR2X1   g0946(.A(n6526), .B(n5827), .Y(n1844));
INVX1    g0947(.A(CRC_OUT_8_21), .Y(n6528));
XOR2X1   g0948(.A(WX3251), .B(TM1), .Y(n6529_1));
XOR2X1   g0949(.A(n6529_1), .B(WX3315), .Y(n6530));
INVX1    g0950(.A(WX3379), .Y(n6531));
XOR2X1   g0951(.A(WX3443), .B(n6531), .Y(n6532));
XOR2X1   g0952(.A(n6532), .B(n6530), .Y(n6533));
MX2X1    g0953(.A(n6528), .B(n6533), .S0(n5539), .Y(n6535));
INVX1    g0954(.A(WX1798), .Y(n6536));
MX2X1    g0955(.A(n6536), .B(n5954), .S0(n5539), .Y(n6537));
MX2X1    g0956(.A(n6535), .B(n6537), .S0(TM1), .Y(n6538));
NOR2X1   g0957(.A(n6538), .B(n5827), .Y(n1849));
INVX1    g0958(.A(CRC_OUT_8_20), .Y(n6540));
XOR2X1   g0959(.A(WX3253), .B(TM1), .Y(n6541));
XOR2X1   g0960(.A(n6541), .B(WX3317), .Y(n6542));
INVX1    g0961(.A(WX3381), .Y(n6543));
XOR2X1   g0962(.A(WX3445), .B(n6543), .Y(n6544_1));
XOR2X1   g0963(.A(n6544_1), .B(n6542), .Y(n6545));
MX2X1    g0964(.A(n6540), .B(n6545), .S0(n5539), .Y(n6547));
INVX1    g0965(.A(WX1800), .Y(n6548));
MX2X1    g0966(.A(n6548), .B(n5966_1), .S0(n5539), .Y(n6549_1));
MX2X1    g0967(.A(n6547), .B(n6549_1), .S0(TM1), .Y(n6550));
NOR2X1   g0968(.A(n6550), .B(n5827), .Y(n1854));
INVX1    g0969(.A(CRC_OUT_8_19), .Y(n6552));
XOR2X1   g0970(.A(WX3255), .B(TM1), .Y(n6553));
XOR2X1   g0971(.A(n6553), .B(WX3319), .Y(n6554_1));
INVX1    g0972(.A(WX3383), .Y(n6555));
XOR2X1   g0973(.A(WX3447), .B(n6555), .Y(n6556));
XOR2X1   g0974(.A(n6556), .B(n6554_1), .Y(n6557));
MX2X1    g0975(.A(n6552), .B(n6557), .S0(n5539), .Y(n6559_1));
INVX1    g0976(.A(WX1802), .Y(n6560));
MX2X1    g0977(.A(n6560), .B(n5978), .S0(n5539), .Y(n6561));
MX2X1    g0978(.A(n6559_1), .B(n6561), .S0(TM1), .Y(n6562));
NOR2X1   g0979(.A(n6562), .B(n5827), .Y(n1859));
INVX1    g0980(.A(CRC_OUT_8_18), .Y(n6564_1));
XOR2X1   g0981(.A(WX3257), .B(TM1), .Y(n6565));
XOR2X1   g0982(.A(n6565), .B(WX3321), .Y(n6566));
INVX1    g0983(.A(WX3385), .Y(n6567));
XOR2X1   g0984(.A(WX3449), .B(n6567), .Y(n6568));
XOR2X1   g0985(.A(n6568), .B(n6566), .Y(n6569_1));
MX2X1    g0986(.A(n6564_1), .B(n6569_1), .S0(n5539), .Y(n6571));
INVX1    g0987(.A(WX1804), .Y(n6572));
MX2X1    g0988(.A(n6572), .B(n5990), .S0(n5539), .Y(n6573));
MX2X1    g0989(.A(n6571), .B(n6573), .S0(TM1), .Y(n6574_1));
NOR2X1   g0990(.A(n6574_1), .B(n5827), .Y(n1864));
INVX1    g0991(.A(CRC_OUT_8_17), .Y(n6576));
XOR2X1   g0992(.A(WX3259), .B(TM1), .Y(n6577));
XOR2X1   g0993(.A(n6577), .B(WX3323), .Y(n6578));
INVX1    g0994(.A(WX3387), .Y(n6579_1));
XOR2X1   g0995(.A(WX3451), .B(n6579_1), .Y(n6580));
XOR2X1   g0996(.A(n6580), .B(n6578), .Y(n6581));
MX2X1    g0997(.A(n6576), .B(n6581), .S0(n5539), .Y(n6583));
INVX1    g0998(.A(WX1806), .Y(n6584_1));
MX2X1    g0999(.A(n6584_1), .B(n6002), .S0(n5539), .Y(n6585));
MX2X1    g1000(.A(n6583), .B(n6585), .S0(TM1), .Y(n6586));
NOR2X1   g1001(.A(n6586), .B(n5827), .Y(n1869));
INVX1    g1002(.A(CRC_OUT_8_16), .Y(n6588));
XOR2X1   g1003(.A(WX3261), .B(TM1), .Y(n6589_1));
XOR2X1   g1004(.A(n6589_1), .B(WX3325), .Y(n6590));
INVX1    g1005(.A(WX3389), .Y(n6591));
XOR2X1   g1006(.A(WX3453), .B(n6591), .Y(n6592));
XOR2X1   g1007(.A(n6592), .B(n6590), .Y(n6593));
MX2X1    g1008(.A(n6588), .B(n6593), .S0(n5539), .Y(n6595));
INVX1    g1009(.A(WX1808), .Y(n6596));
MX2X1    g1010(.A(n6596), .B(n6014), .S0(n5539), .Y(n6597));
MX2X1    g1011(.A(n6595), .B(n6597), .S0(TM1), .Y(n6598));
NOR2X1   g1012(.A(n6598), .B(n5827), .Y(n1874));
INVX1    g1013(.A(CRC_OUT_8_15), .Y(n6600));
XOR2X1   g1014(.A(WX3263), .B(TM0), .Y(n6601));
XOR2X1   g1015(.A(n6601), .B(WX3327), .Y(n6602));
INVX1    g1016(.A(WX3391), .Y(n6603));
XOR2X1   g1017(.A(WX3455), .B(n6603), .Y(n6604_1));
XOR2X1   g1018(.A(n6604_1), .B(n6602), .Y(n6605));
MX2X1    g1019(.A(n6600), .B(n6605), .S0(n5539), .Y(n6607));
INVX1    g1020(.A(WX1810), .Y(n6608));
MX2X1    g1021(.A(n6608), .B(n6026_1), .S0(n5539), .Y(n6609_1));
MX2X1    g1022(.A(n6607), .B(n6609_1), .S0(TM1), .Y(n6610));
NOR2X1   g1023(.A(n6610), .B(n5827), .Y(n1879));
INVX1    g1024(.A(CRC_OUT_8_14), .Y(n6612));
XOR2X1   g1025(.A(WX3265), .B(TM0), .Y(n6613));
XOR2X1   g1026(.A(n6613), .B(WX3329), .Y(n6614_1));
INVX1    g1027(.A(WX3393), .Y(n6615));
XOR2X1   g1028(.A(WX3457), .B(n6615), .Y(n6616));
XOR2X1   g1029(.A(n6616), .B(n6614_1), .Y(n6617));
MX2X1    g1030(.A(n6612), .B(n6617), .S0(n5539), .Y(n6619_1));
INVX1    g1031(.A(WX1812), .Y(n6620));
MX2X1    g1032(.A(n6620), .B(n6038), .S0(n5539), .Y(n6621));
MX2X1    g1033(.A(n6619_1), .B(n6621), .S0(TM1), .Y(n6622));
NOR2X1   g1034(.A(n6622), .B(n5827), .Y(n1884));
INVX1    g1035(.A(CRC_OUT_8_13), .Y(n6624_1));
XOR2X1   g1036(.A(WX3267), .B(TM0), .Y(n6625));
XOR2X1   g1037(.A(n6625), .B(WX3331), .Y(n6626));
INVX1    g1038(.A(WX3395), .Y(n6627));
XOR2X1   g1039(.A(WX3459), .B(n6627), .Y(n6628));
XOR2X1   g1040(.A(n6628), .B(n6626), .Y(n6629_1));
MX2X1    g1041(.A(n6624_1), .B(n6629_1), .S0(n5539), .Y(n6631));
INVX1    g1042(.A(WX1814), .Y(n6632));
MX2X1    g1043(.A(n6632), .B(n6050), .S0(n5539), .Y(n6633));
MX2X1    g1044(.A(n6631), .B(n6633), .S0(TM1), .Y(n6634_1));
NOR2X1   g1045(.A(n6634_1), .B(n5827), .Y(n1889));
INVX1    g1046(.A(CRC_OUT_8_12), .Y(n6636));
XOR2X1   g1047(.A(WX3269), .B(TM0), .Y(n6637));
XOR2X1   g1048(.A(n6637), .B(WX3333), .Y(n6638));
INVX1    g1049(.A(WX3397), .Y(n6639_1));
XOR2X1   g1050(.A(WX3461), .B(n6639_1), .Y(n6640));
XOR2X1   g1051(.A(n6640), .B(n6638), .Y(n6641));
MX2X1    g1052(.A(n6636), .B(n6641), .S0(n5539), .Y(n6643));
INVX1    g1053(.A(WX1816), .Y(n6644_1));
MX2X1    g1054(.A(n6644_1), .B(n6062), .S0(n5539), .Y(n6645));
MX2X1    g1055(.A(n6643), .B(n6645), .S0(TM1), .Y(n6646));
NOR2X1   g1056(.A(n6646), .B(n5827), .Y(n1894));
INVX1    g1057(.A(CRC_OUT_8_11), .Y(n6648));
XOR2X1   g1058(.A(WX3271), .B(TM0), .Y(n6649_1));
XOR2X1   g1059(.A(n6649_1), .B(WX3335), .Y(n6650));
INVX1    g1060(.A(WX3399), .Y(n6651));
XOR2X1   g1061(.A(WX3463), .B(n6651), .Y(n6652));
XOR2X1   g1062(.A(n6652), .B(n6650), .Y(n6653));
MX2X1    g1063(.A(n6648), .B(n6653), .S0(n5539), .Y(n6655));
INVX1    g1064(.A(WX1818), .Y(n6656));
MX2X1    g1065(.A(n6656), .B(n6074), .S0(n5539), .Y(n6657));
MX2X1    g1066(.A(n6655), .B(n6657), .S0(TM1), .Y(n6658));
NOR2X1   g1067(.A(n6658), .B(n5827), .Y(n1899));
INVX1    g1068(.A(CRC_OUT_8_10), .Y(n6660));
XOR2X1   g1069(.A(WX3273), .B(TM0), .Y(n6661));
XOR2X1   g1070(.A(n6661), .B(WX3337), .Y(n6662));
INVX1    g1071(.A(WX3401), .Y(n6663));
XOR2X1   g1072(.A(WX3465), .B(n6663), .Y(n6664_1));
XOR2X1   g1073(.A(n6664_1), .B(n6662), .Y(n6665));
MX2X1    g1074(.A(n6660), .B(n6665), .S0(n5539), .Y(n6667));
INVX1    g1075(.A(WX1820), .Y(n6668));
MX2X1    g1076(.A(n6668), .B(n6086_1), .S0(n5539), .Y(n6669_1));
MX2X1    g1077(.A(n6667), .B(n6669_1), .S0(TM1), .Y(n6670));
NOR2X1   g1078(.A(n6670), .B(n5827), .Y(n1904));
INVX1    g1079(.A(CRC_OUT_8_9), .Y(n6672));
XOR2X1   g1080(.A(WX3275), .B(TM0), .Y(n6673));
XOR2X1   g1081(.A(n6673), .B(WX3339), .Y(n6674_1));
INVX1    g1082(.A(WX3403), .Y(n6675));
XOR2X1   g1083(.A(WX3467), .B(n6675), .Y(n6676));
XOR2X1   g1084(.A(n6676), .B(n6674_1), .Y(n6677));
MX2X1    g1085(.A(n6672), .B(n6677), .S0(n5539), .Y(n6679_1));
INVX1    g1086(.A(WX1822), .Y(n6680));
MX2X1    g1087(.A(n6680), .B(n6098), .S0(n5539), .Y(n6681));
MX2X1    g1088(.A(n6679_1), .B(n6681), .S0(TM1), .Y(n6682));
NOR2X1   g1089(.A(n6682), .B(n5827), .Y(n1909));
INVX1    g1090(.A(CRC_OUT_8_8), .Y(n6684_1));
XOR2X1   g1091(.A(WX3277), .B(TM0), .Y(n6685));
XOR2X1   g1092(.A(n6685), .B(WX3341), .Y(n6686));
INVX1    g1093(.A(WX3405), .Y(n6687));
XOR2X1   g1094(.A(WX3469), .B(n6687), .Y(n6688));
XOR2X1   g1095(.A(n6688), .B(n6686), .Y(n6689_1));
MX2X1    g1096(.A(n6684_1), .B(n6689_1), .S0(n5539), .Y(n6691));
INVX1    g1097(.A(WX1824), .Y(n6692));
MX2X1    g1098(.A(n6692), .B(n6110), .S0(n5539), .Y(n6693));
MX2X1    g1099(.A(n6691), .B(n6693), .S0(TM1), .Y(n6694_1));
NOR2X1   g1100(.A(n6694_1), .B(n5827), .Y(n1914));
INVX1    g1101(.A(CRC_OUT_8_7), .Y(n6696));
XOR2X1   g1102(.A(WX3279), .B(TM0), .Y(n6697));
XOR2X1   g1103(.A(n6697), .B(WX3343), .Y(n6698));
INVX1    g1104(.A(WX3407), .Y(n6699_1));
XOR2X1   g1105(.A(WX3471), .B(n6699_1), .Y(n6700));
XOR2X1   g1106(.A(n6700), .B(n6698), .Y(n6701));
MX2X1    g1107(.A(n6696), .B(n6701), .S0(n5539), .Y(n6703));
INVX1    g1108(.A(WX1826), .Y(n6704_1));
MX2X1    g1109(.A(n6704_1), .B(n6122), .S0(n5539), .Y(n6705));
MX2X1    g1110(.A(n6703), .B(n6705), .S0(TM1), .Y(n6706));
NOR2X1   g1111(.A(n6706), .B(n5827), .Y(n1919));
INVX1    g1112(.A(CRC_OUT_8_6), .Y(n6708));
XOR2X1   g1113(.A(WX3281), .B(TM0), .Y(n6709_1));
XOR2X1   g1114(.A(n6709_1), .B(WX3345), .Y(n6710));
INVX1    g1115(.A(WX3409), .Y(n6711));
XOR2X1   g1116(.A(WX3473), .B(n6711), .Y(n6712));
XOR2X1   g1117(.A(n6712), .B(n6710), .Y(n6713));
MX2X1    g1118(.A(n6708), .B(n6713), .S0(n5539), .Y(n6715));
INVX1    g1119(.A(WX1828), .Y(n6716));
MX2X1    g1120(.A(n6716), .B(n6134), .S0(n5539), .Y(n6717));
MX2X1    g1121(.A(n6715), .B(n6717), .S0(TM1), .Y(n6718));
NOR2X1   g1122(.A(n6718), .B(n5827), .Y(n1924));
INVX1    g1123(.A(CRC_OUT_8_5), .Y(n6720));
XOR2X1   g1124(.A(WX3283), .B(TM0), .Y(n6721));
XOR2X1   g1125(.A(n6721), .B(WX3347), .Y(n6722));
INVX1    g1126(.A(WX3411), .Y(n6723));
XOR2X1   g1127(.A(WX3475), .B(n6723), .Y(n6724_1));
XOR2X1   g1128(.A(n6724_1), .B(n6722), .Y(n6725));
MX2X1    g1129(.A(n6720), .B(n6725), .S0(n5539), .Y(n6727));
INVX1    g1130(.A(WX1830), .Y(n6728));
MX2X1    g1131(.A(n6728), .B(n6146_1), .S0(n5539), .Y(n6729_1));
MX2X1    g1132(.A(n6727), .B(n6729_1), .S0(TM1), .Y(n6730));
NOR2X1   g1133(.A(n6730), .B(n5827), .Y(n1929));
INVX1    g1134(.A(CRC_OUT_8_4), .Y(n6732));
XOR2X1   g1135(.A(WX3285), .B(TM0), .Y(n6733));
XOR2X1   g1136(.A(n6733), .B(WX3349), .Y(n6734_1));
INVX1    g1137(.A(WX3413), .Y(n6735));
XOR2X1   g1138(.A(WX3477), .B(n6735), .Y(n6736));
XOR2X1   g1139(.A(n6736), .B(n6734_1), .Y(n6737));
MX2X1    g1140(.A(n6732), .B(n6737), .S0(n5539), .Y(n6739_1));
INVX1    g1141(.A(WX1832), .Y(n6740));
MX2X1    g1142(.A(n6740), .B(n6158), .S0(n5539), .Y(n6741));
MX2X1    g1143(.A(n6739_1), .B(n6741), .S0(TM1), .Y(n6742));
NOR2X1   g1144(.A(n6742), .B(n5827), .Y(n1934));
INVX1    g1145(.A(CRC_OUT_8_3), .Y(n6744_1));
XOR2X1   g1146(.A(WX3287), .B(TM0), .Y(n6745));
XOR2X1   g1147(.A(n6745), .B(WX3351), .Y(n6746));
INVX1    g1148(.A(WX3415), .Y(n6747));
XOR2X1   g1149(.A(WX3479), .B(n6747), .Y(n6748));
XOR2X1   g1150(.A(n6748), .B(n6746), .Y(n6749_1));
MX2X1    g1151(.A(n6744_1), .B(n6749_1), .S0(n5539), .Y(n6751));
INVX1    g1152(.A(WX1834), .Y(n6752));
MX2X1    g1153(.A(n6752), .B(n6170), .S0(n5539), .Y(n6753));
MX2X1    g1154(.A(n6751), .B(n6753), .S0(TM1), .Y(n6754_1));
NOR2X1   g1155(.A(n6754_1), .B(n5827), .Y(n1939));
INVX1    g1156(.A(CRC_OUT_8_2), .Y(n6756));
XOR2X1   g1157(.A(WX3289), .B(TM0), .Y(n6757));
XOR2X1   g1158(.A(n6757), .B(WX3353), .Y(n6758));
INVX1    g1159(.A(WX3417), .Y(n6759_1));
XOR2X1   g1160(.A(WX3481), .B(n6759_1), .Y(n6760));
XOR2X1   g1161(.A(n6760), .B(n6758), .Y(n6761));
MX2X1    g1162(.A(n6756), .B(n6761), .S0(n5539), .Y(n6763));
INVX1    g1163(.A(WX1836), .Y(n6764_1));
MX2X1    g1164(.A(n6764_1), .B(n6182), .S0(n5539), .Y(n6765));
MX2X1    g1165(.A(n6763), .B(n6765), .S0(TM1), .Y(n6766));
NOR2X1   g1166(.A(n6766), .B(n5827), .Y(n1944));
INVX1    g1167(.A(CRC_OUT_8_1), .Y(n6768));
XOR2X1   g1168(.A(WX3291), .B(TM0), .Y(n6769_1));
XOR2X1   g1169(.A(n6769_1), .B(WX3355), .Y(n6770));
INVX1    g1170(.A(WX3419), .Y(n6771));
XOR2X1   g1171(.A(WX3483), .B(n6771), .Y(n6772));
XOR2X1   g1172(.A(n6772), .B(n6770), .Y(n6773));
MX2X1    g1173(.A(n6768), .B(n6773), .S0(n5539), .Y(n6775));
INVX1    g1174(.A(WX1838), .Y(n6776));
MX2X1    g1175(.A(n6776), .B(n6194), .S0(n5539), .Y(n6777));
MX2X1    g1176(.A(n6775), .B(n6777), .S0(TM1), .Y(n6778));
NOR2X1   g1177(.A(n6778), .B(n5827), .Y(n1949));
INVX1    g1178(.A(CRC_OUT_8_0), .Y(n6780));
XOR2X1   g1179(.A(WX3293), .B(TM0), .Y(n6781));
XOR2X1   g1180(.A(n6781), .B(WX3357), .Y(n6782));
INVX1    g1181(.A(WX3421), .Y(n6783));
XOR2X1   g1182(.A(WX3485), .B(n6783), .Y(n6784_1));
XOR2X1   g1183(.A(n6784_1), .B(n6782), .Y(n6785));
MX2X1    g1184(.A(n6780), .B(n6785), .S0(n5539), .Y(n6787));
INVX1    g1185(.A(WX1840), .Y(n6788));
MX2X1    g1186(.A(n6788), .B(n6206), .S0(n5539), .Y(n6789_1));
MX2X1    g1187(.A(n6787), .B(n6789_1), .S0(TM1), .Y(n6790));
NOR2X1   g1188(.A(n6790), .B(n5827), .Y(n1954));
AND2X1   g1189(.A(WX1938), .B(RESET), .Y(n1959));
AND2X1   g1190(.A(WX1940), .B(RESET), .Y(n1964));
AND2X1   g1191(.A(WX1942), .B(RESET), .Y(n1969));
AND2X1   g1192(.A(WX1944), .B(RESET), .Y(n1974));
AND2X1   g1193(.A(WX1946), .B(RESET), .Y(n1979));
AND2X1   g1194(.A(WX1948), .B(RESET), .Y(n1984));
AND2X1   g1195(.A(WX1950), .B(RESET), .Y(n1989));
AND2X1   g1196(.A(WX1952), .B(RESET), .Y(n1994));
AND2X1   g1197(.A(WX1954), .B(RESET), .Y(n1999));
AND2X1   g1198(.A(WX1956), .B(RESET), .Y(n2004));
AND2X1   g1199(.A(WX1958), .B(RESET), .Y(n2009));
AND2X1   g1200(.A(WX1960), .B(RESET), .Y(n2014));
AND2X1   g1201(.A(WX1962), .B(RESET), .Y(n2019));
AND2X1   g1202(.A(WX1964), .B(RESET), .Y(n2024));
AND2X1   g1203(.A(WX1966), .B(RESET), .Y(n2029));
AND2X1   g1204(.A(WX1968), .B(RESET), .Y(n2034));
AND2X1   g1205(.A(WX1970), .B(RESET), .Y(n2039));
AND2X1   g1206(.A(WX1972), .B(RESET), .Y(n2044));
AND2X1   g1207(.A(WX1974), .B(RESET), .Y(n2049));
AND2X1   g1208(.A(WX1976), .B(RESET), .Y(n2054));
AND2X1   g1209(.A(WX1978), .B(RESET), .Y(n2059));
AND2X1   g1210(.A(WX1980), .B(RESET), .Y(n2064));
AND2X1   g1211(.A(WX1982), .B(RESET), .Y(n2069));
AND2X1   g1212(.A(WX1984), .B(RESET), .Y(n2074));
AND2X1   g1213(.A(WX1986), .B(RESET), .Y(n2079));
AND2X1   g1214(.A(WX1988), .B(RESET), .Y(n2084));
AND2X1   g1215(.A(WX1990), .B(RESET), .Y(n2089));
AND2X1   g1216(.A(WX1992), .B(RESET), .Y(n2094));
AND2X1   g1217(.A(WX1994), .B(RESET), .Y(n2099));
AND2X1   g1218(.A(WX1996), .B(RESET), .Y(n2104));
AND2X1   g1219(.A(WX1998), .B(RESET), .Y(n2109));
AND2X1   g1220(.A(WX2000), .B(RESET), .Y(n2114));
AND2X1   g1221(.A(WX2002), .B(RESET), .Y(n2119));
AND2X1   g1222(.A(WX2004), .B(RESET), .Y(n2124));
AND2X1   g1223(.A(WX2006), .B(RESET), .Y(n2129));
AND2X1   g1224(.A(WX2008), .B(RESET), .Y(n2134));
AND2X1   g1225(.A(WX2010), .B(RESET), .Y(n2139));
AND2X1   g1226(.A(WX2012), .B(RESET), .Y(n2144));
AND2X1   g1227(.A(WX2014), .B(RESET), .Y(n2149));
AND2X1   g1228(.A(WX2016), .B(RESET), .Y(n2154));
AND2X1   g1229(.A(WX2018), .B(RESET), .Y(n2159));
AND2X1   g1230(.A(WX2020), .B(RESET), .Y(n2164));
AND2X1   g1231(.A(WX2022), .B(RESET), .Y(n2169));
AND2X1   g1232(.A(WX2024), .B(RESET), .Y(n2174));
AND2X1   g1233(.A(WX2026), .B(RESET), .Y(n2179));
AND2X1   g1234(.A(WX2028), .B(RESET), .Y(n2184));
AND2X1   g1235(.A(WX2030), .B(RESET), .Y(n2189));
AND2X1   g1236(.A(WX2032), .B(RESET), .Y(n2194));
AND2X1   g1237(.A(WX2034), .B(RESET), .Y(n2199));
AND2X1   g1238(.A(WX2036), .B(RESET), .Y(n2204));
AND2X1   g1239(.A(WX2038), .B(RESET), .Y(n2209));
AND2X1   g1240(.A(WX2040), .B(RESET), .Y(n2214));
AND2X1   g1241(.A(WX2042), .B(RESET), .Y(n2219));
AND2X1   g1242(.A(WX2044), .B(RESET), .Y(n2224));
AND2X1   g1243(.A(WX2046), .B(RESET), .Y(n2229));
AND2X1   g1244(.A(WX2048), .B(RESET), .Y(n2234));
AND2X1   g1245(.A(WX2050), .B(RESET), .Y(n2239));
AND2X1   g1246(.A(WX2052), .B(RESET), .Y(n2244));
AND2X1   g1247(.A(WX2054), .B(RESET), .Y(n2249));
AND2X1   g1248(.A(WX2056), .B(RESET), .Y(n2254));
AND2X1   g1249(.A(WX2058), .B(RESET), .Y(n2259));
AND2X1   g1250(.A(WX2060), .B(RESET), .Y(n2264));
AND2X1   g1251(.A(WX2062), .B(RESET), .Y(n2269));
AND2X1   g1252(.A(WX2064), .B(RESET), .Y(n2274));
AND2X1   g1253(.A(WX2066), .B(RESET), .Y(n2279));
AND2X1   g1254(.A(WX2068), .B(RESET), .Y(n2284));
AND2X1   g1255(.A(WX2070), .B(RESET), .Y(n2289));
AND2X1   g1256(.A(WX2072), .B(RESET), .Y(n2294));
AND2X1   g1257(.A(WX2074), .B(RESET), .Y(n2299));
AND2X1   g1258(.A(WX2076), .B(RESET), .Y(n2304));
AND2X1   g1259(.A(WX2078), .B(RESET), .Y(n2309));
AND2X1   g1260(.A(WX2080), .B(RESET), .Y(n2314));
AND2X1   g1261(.A(WX2082), .B(RESET), .Y(n2319));
AND2X1   g1262(.A(WX2084), .B(RESET), .Y(n2324));
AND2X1   g1263(.A(WX2086), .B(RESET), .Y(n2329));
AND2X1   g1264(.A(WX2088), .B(RESET), .Y(n2334));
AND2X1   g1265(.A(WX2090), .B(RESET), .Y(n2339));
AND2X1   g1266(.A(WX2092), .B(RESET), .Y(n2344));
AND2X1   g1267(.A(WX2094), .B(RESET), .Y(n2349));
AND2X1   g1268(.A(WX2096), .B(RESET), .Y(n2354));
AND2X1   g1269(.A(WX2098), .B(RESET), .Y(n2359));
AND2X1   g1270(.A(WX2100), .B(RESET), .Y(n2364));
AND2X1   g1271(.A(WX2102), .B(RESET), .Y(n2369));
AND2X1   g1272(.A(WX2104), .B(RESET), .Y(n2374));
AND2X1   g1273(.A(WX2106), .B(RESET), .Y(n2379));
AND2X1   g1274(.A(WX2108), .B(RESET), .Y(n2384));
AND2X1   g1275(.A(WX2110), .B(RESET), .Y(n2389));
AND2X1   g1276(.A(WX2112), .B(RESET), .Y(n2394));
AND2X1   g1277(.A(WX2114), .B(RESET), .Y(n2399));
AND2X1   g1278(.A(WX2116), .B(RESET), .Y(n2404));
AND2X1   g1279(.A(WX2118), .B(RESET), .Y(n2409));
AND2X1   g1280(.A(WX2120), .B(RESET), .Y(n2414));
AND2X1   g1281(.A(WX2122), .B(RESET), .Y(n2419));
AND2X1   g1282(.A(WX2124), .B(RESET), .Y(n2424));
AND2X1   g1283(.A(WX2126), .B(RESET), .Y(n2429));
AND2X1   g1284(.A(WX2128), .B(RESET), .Y(n2434));
XOR2X1   g1285(.A(CRC_OUT_8_31), .B(WX2192), .Y(n6888));
NOR2X1   g1286(.A(n6888), .B(n5827), .Y(CRC_OUT_8_0));
XOR2X1   g1287(.A(CRC_OUT_8_0), .B(WX2190), .Y(n6890));
NOR2X1   g1288(.A(n6890), .B(n5827), .Y(CRC_OUT_8_1));
XOR2X1   g1289(.A(CRC_OUT_8_1), .B(WX2188), .Y(n6892));
NOR2X1   g1290(.A(n6892), .B(n5827), .Y(CRC_OUT_8_2));
XOR2X1   g1291(.A(CRC_OUT_8_2), .B(WX2186), .Y(n6894_1));
NOR2X1   g1292(.A(n6894_1), .B(n5827), .Y(CRC_OUT_8_3));
XOR2X1   g1293(.A(CRC_OUT_8_31), .B(WX2184), .Y(n6896));
XOR2X1   g1294(.A(n6896), .B(CRC_OUT_8_3), .Y(n6897));
NOR2X1   g1295(.A(n6897), .B(n5827), .Y(CRC_OUT_8_4));
XOR2X1   g1296(.A(CRC_OUT_8_4), .B(WX2182), .Y(n6899_1));
NOR2X1   g1297(.A(n6899_1), .B(n5827), .Y(CRC_OUT_8_5));
XOR2X1   g1298(.A(CRC_OUT_8_5), .B(WX2180), .Y(n6901));
NOR2X1   g1299(.A(n6901), .B(n5827), .Y(CRC_OUT_8_6));
XOR2X1   g1300(.A(CRC_OUT_8_6), .B(WX2178), .Y(n6903));
NOR2X1   g1301(.A(n6903), .B(n5827), .Y(CRC_OUT_8_7));
XOR2X1   g1302(.A(CRC_OUT_8_7), .B(WX2176), .Y(n6905));
NOR2X1   g1303(.A(n6905), .B(n5827), .Y(CRC_OUT_8_8));
XOR2X1   g1304(.A(CRC_OUT_8_8), .B(WX2174), .Y(n6907));
NOR2X1   g1305(.A(n6907), .B(n5827), .Y(CRC_OUT_8_9));
XOR2X1   g1306(.A(CRC_OUT_8_9), .B(WX2172), .Y(n6909_1));
NOR2X1   g1307(.A(n6909_1), .B(n5827), .Y(CRC_OUT_8_10));
XOR2X1   g1308(.A(CRC_OUT_8_31), .B(WX2170), .Y(n6911));
XOR2X1   g1309(.A(n6911), .B(CRC_OUT_8_10), .Y(n6912));
NOR2X1   g1310(.A(n6912), .B(n5827), .Y(CRC_OUT_8_11));
XOR2X1   g1311(.A(CRC_OUT_8_11), .B(WX2168), .Y(n6914_1));
NOR2X1   g1312(.A(n6914_1), .B(n5827), .Y(CRC_OUT_8_12));
XOR2X1   g1313(.A(CRC_OUT_8_12), .B(WX2166), .Y(n6916));
NOR2X1   g1314(.A(n6916), .B(n5827), .Y(CRC_OUT_8_13));
XOR2X1   g1315(.A(CRC_OUT_8_13), .B(WX2164), .Y(n6918));
NOR2X1   g1316(.A(n6918), .B(n5827), .Y(CRC_OUT_8_14));
XOR2X1   g1317(.A(CRC_OUT_8_14), .B(WX2162), .Y(n6920));
NOR2X1   g1318(.A(n6920), .B(n5827), .Y(CRC_OUT_8_15));
XOR2X1   g1319(.A(CRC_OUT_8_31), .B(WX2160), .Y(n6922));
XOR2X1   g1320(.A(n6922), .B(CRC_OUT_8_15), .Y(n6923));
NOR2X1   g1321(.A(n6923), .B(n5827), .Y(CRC_OUT_8_16));
XOR2X1   g1322(.A(CRC_OUT_8_16), .B(WX2158), .Y(n6925));
NOR2X1   g1323(.A(n6925), .B(n5827), .Y(CRC_OUT_8_17));
XOR2X1   g1324(.A(CRC_OUT_8_17), .B(WX2156), .Y(n6927));
NOR2X1   g1325(.A(n6927), .B(n5827), .Y(CRC_OUT_8_18));
XOR2X1   g1326(.A(CRC_OUT_8_18), .B(WX2154), .Y(n6929_1));
NOR2X1   g1327(.A(n6929_1), .B(n5827), .Y(CRC_OUT_8_19));
XOR2X1   g1328(.A(CRC_OUT_8_19), .B(WX2152), .Y(n6931));
NOR2X1   g1329(.A(n6931), .B(n5827), .Y(CRC_OUT_8_20));
XOR2X1   g1330(.A(CRC_OUT_8_20), .B(WX2150), .Y(n6933));
NOR2X1   g1331(.A(n6933), .B(n5827), .Y(CRC_OUT_8_21));
XOR2X1   g1332(.A(CRC_OUT_8_21), .B(WX2148), .Y(n6935));
NOR2X1   g1333(.A(n6935), .B(n5827), .Y(CRC_OUT_8_22));
XOR2X1   g1334(.A(CRC_OUT_8_22), .B(WX2146), .Y(n6937));
NOR2X1   g1335(.A(n6937), .B(n5827), .Y(CRC_OUT_8_23));
XOR2X1   g1336(.A(CRC_OUT_8_23), .B(WX2144), .Y(n6939_1));
NOR2X1   g1337(.A(n6939_1), .B(n5827), .Y(CRC_OUT_8_24));
XOR2X1   g1338(.A(CRC_OUT_8_24), .B(WX2142), .Y(n6941));
NOR2X1   g1339(.A(n6941), .B(n5827), .Y(CRC_OUT_8_25));
XOR2X1   g1340(.A(CRC_OUT_8_25), .B(WX2140), .Y(n6943));
NOR2X1   g1341(.A(n6943), .B(n5827), .Y(CRC_OUT_8_26));
XOR2X1   g1342(.A(CRC_OUT_8_26), .B(WX2138), .Y(n6945));
NOR2X1   g1343(.A(n6945), .B(n5827), .Y(CRC_OUT_8_27));
XOR2X1   g1344(.A(CRC_OUT_8_27), .B(WX2136), .Y(n6947));
NOR2X1   g1345(.A(n6947), .B(n5827), .Y(CRC_OUT_8_28));
XOR2X1   g1346(.A(CRC_OUT_8_28), .B(WX2134), .Y(n6949_1));
NOR2X1   g1347(.A(n6949_1), .B(n5827), .Y(CRC_OUT_8_29));
XOR2X1   g1348(.A(CRC_OUT_8_29), .B(WX2132), .Y(n6951));
NOR2X1   g1349(.A(n6951), .B(n5827), .Y(CRC_OUT_8_30));
XOR2X1   g1350(.A(CRC_OUT_8_30), .B(WX2130), .Y(n6953));
NOR2X1   g1351(.A(n6953), .B(n5827), .Y(CRC_OUT_8_31));
AND2X1   g1352(.A(WX3073), .B(RESET), .Y(n2567));
AND2X1   g1353(.A(WX3075), .B(RESET), .Y(n2572));
AND2X1   g1354(.A(WX3077), .B(RESET), .Y(n2577));
AND2X1   g1355(.A(WX3079), .B(RESET), .Y(n2582));
AND2X1   g1356(.A(WX3081), .B(RESET), .Y(n2587));
AND2X1   g1357(.A(WX3083), .B(RESET), .Y(n2592));
AND2X1   g1358(.A(WX3085), .B(RESET), .Y(n2597));
AND2X1   g1359(.A(WX3087), .B(RESET), .Y(n2602));
AND2X1   g1360(.A(WX3089), .B(RESET), .Y(n2607));
AND2X1   g1361(.A(WX3091), .B(RESET), .Y(n2612));
AND2X1   g1362(.A(WX3093), .B(RESET), .Y(n2617));
AND2X1   g1363(.A(WX3095), .B(RESET), .Y(n2622));
AND2X1   g1364(.A(WX3097), .B(RESET), .Y(n2627));
AND2X1   g1365(.A(WX3099), .B(RESET), .Y(n2632));
AND2X1   g1366(.A(WX3101), .B(RESET), .Y(n2637));
AND2X1   g1367(.A(WX3103), .B(RESET), .Y(n2642));
AND2X1   g1368(.A(WX3105), .B(RESET), .Y(n2647));
AND2X1   g1369(.A(WX3107), .B(RESET), .Y(n2652));
AND2X1   g1370(.A(WX3109), .B(RESET), .Y(n2657));
AND2X1   g1371(.A(WX3111), .B(RESET), .Y(n2662));
AND2X1   g1372(.A(WX3113), .B(RESET), .Y(n2667));
AND2X1   g1373(.A(WX3115), .B(RESET), .Y(n2672));
AND2X1   g1374(.A(WX3117), .B(RESET), .Y(n2677));
AND2X1   g1375(.A(WX3119), .B(RESET), .Y(n2682));
AND2X1   g1376(.A(WX3121), .B(RESET), .Y(n2687));
AND2X1   g1377(.A(WX3123), .B(RESET), .Y(n2692));
AND2X1   g1378(.A(WX3125), .B(RESET), .Y(n2697));
AND2X1   g1379(.A(WX3127), .B(RESET), .Y(n2702));
AND2X1   g1380(.A(WX3129), .B(RESET), .Y(n2707));
AND2X1   g1381(.A(WX3131), .B(RESET), .Y(n2712));
AND2X1   g1382(.A(WX3133), .B(RESET), .Y(n2717));
NOR2X1   g1383(.A(WX3071), .B(n5827), .Y(n2722));
INVX1    g1384(.A(CRC_OUT_7_31), .Y(n6987));
XOR2X1   g1385(.A(WX4524), .B(TM1), .Y(n6988));
XOR2X1   g1386(.A(n6988), .B(WX4588), .Y(n6989_1));
INVX1    g1387(.A(WX4652), .Y(n6990));
XOR2X1   g1388(.A(WX4716), .B(n6990), .Y(n6991));
XOR2X1   g1389(.A(n6991), .B(n6989_1), .Y(n6992));
MX2X1    g1390(.A(n6987), .B(n6992), .S0(n5539), .Y(n6994_1));
INVX1    g1391(.A(WX3071), .Y(n6995));
MX2X1    g1392(.A(n6995), .B(n6413), .S0(n5539), .Y(n6996));
MX2X1    g1393(.A(n6994_1), .B(n6996), .S0(TM1), .Y(n6997));
NOR2X1   g1394(.A(n6997), .B(n5827), .Y(n2727));
INVX1    g1395(.A(CRC_OUT_7_30), .Y(n6999_1));
XOR2X1   g1396(.A(WX4526), .B(TM1), .Y(n7000));
XOR2X1   g1397(.A(n7000), .B(WX4590), .Y(n7001));
INVX1    g1398(.A(WX4654), .Y(n7002));
XOR2X1   g1399(.A(WX4718), .B(n7002), .Y(n7003));
XOR2X1   g1400(.A(n7003), .B(n7001), .Y(n7004_1));
MX2X1    g1401(.A(n6999_1), .B(n7004_1), .S0(n5539), .Y(n7006));
INVX1    g1402(.A(WX3073), .Y(n7007));
MX2X1    g1403(.A(n7007), .B(n6425), .S0(n5539), .Y(n7008));
MX2X1    g1404(.A(n7006), .B(n7008), .S0(TM1), .Y(n7009_1));
NOR2X1   g1405(.A(n7009_1), .B(n5827), .Y(n2732));
INVX1    g1406(.A(CRC_OUT_7_29), .Y(n7011));
XOR2X1   g1407(.A(WX4528), .B(TM1), .Y(n7012));
XOR2X1   g1408(.A(n7012), .B(WX4592), .Y(n7013));
INVX1    g1409(.A(WX4656), .Y(n7014_1));
XOR2X1   g1410(.A(WX4720), .B(n7014_1), .Y(n7015));
XOR2X1   g1411(.A(n7015), .B(n7013), .Y(n7016));
MX2X1    g1412(.A(n7011), .B(n7016), .S0(n5539), .Y(n7018));
INVX1    g1413(.A(WX3075), .Y(n7019_1));
MX2X1    g1414(.A(n7019_1), .B(n6437), .S0(n5539), .Y(n7020));
MX2X1    g1415(.A(n7018), .B(n7020), .S0(TM1), .Y(n7021));
NOR2X1   g1416(.A(n7021), .B(n5827), .Y(n2737));
INVX1    g1417(.A(CRC_OUT_7_28), .Y(n7023));
XOR2X1   g1418(.A(WX4530), .B(TM1), .Y(n7024_1));
XOR2X1   g1419(.A(n7024_1), .B(WX4594), .Y(n7025));
INVX1    g1420(.A(WX4658), .Y(n7026));
XOR2X1   g1421(.A(WX4722), .B(n7026), .Y(n7027));
XOR2X1   g1422(.A(n7027), .B(n7025), .Y(n7028));
MX2X1    g1423(.A(n7023), .B(n7028), .S0(n5539), .Y(n7030));
INVX1    g1424(.A(WX3077), .Y(n7031));
MX2X1    g1425(.A(n7031), .B(n6449_1), .S0(n5539), .Y(n7032));
MX2X1    g1426(.A(n7030), .B(n7032), .S0(TM1), .Y(n7033));
NOR2X1   g1427(.A(n7033), .B(n5827), .Y(n2742));
INVX1    g1428(.A(CRC_OUT_7_27), .Y(n7035));
XOR2X1   g1429(.A(WX4532), .B(TM1), .Y(n7036));
XOR2X1   g1430(.A(n7036), .B(WX4596), .Y(n7037));
INVX1    g1431(.A(WX4660), .Y(n7038));
XOR2X1   g1432(.A(WX4724), .B(n7038), .Y(n7039_1));
XOR2X1   g1433(.A(n7039_1), .B(n7037), .Y(n7040));
MX2X1    g1434(.A(n7035), .B(n7040), .S0(n5539), .Y(n7042));
INVX1    g1435(.A(WX3079), .Y(n7043));
MX2X1    g1436(.A(n7043), .B(n6461), .S0(n5539), .Y(n7044_1));
MX2X1    g1437(.A(n7042), .B(n7044_1), .S0(TM1), .Y(n7045));
NOR2X1   g1438(.A(n7045), .B(n5827), .Y(n2747));
INVX1    g1439(.A(CRC_OUT_7_26), .Y(n7047));
XOR2X1   g1440(.A(WX4534), .B(TM1), .Y(n7048));
XOR2X1   g1441(.A(n7048), .B(WX4598), .Y(n7049_1));
INVX1    g1442(.A(WX4662), .Y(n7050));
XOR2X1   g1443(.A(WX4726), .B(n7050), .Y(n7051));
XOR2X1   g1444(.A(n7051), .B(n7049_1), .Y(n7052));
MX2X1    g1445(.A(n7047), .B(n7052), .S0(n5539), .Y(n7054_1));
INVX1    g1446(.A(WX3081), .Y(n7055));
MX2X1    g1447(.A(n7055), .B(n6473), .S0(n5539), .Y(n7056));
MX2X1    g1448(.A(n7054_1), .B(n7056), .S0(TM1), .Y(n7057));
NOR2X1   g1449(.A(n7057), .B(n5827), .Y(n2752));
INVX1    g1450(.A(CRC_OUT_7_25), .Y(n7059_1));
XOR2X1   g1451(.A(WX4536), .B(TM1), .Y(n7060));
XOR2X1   g1452(.A(n7060), .B(WX4600), .Y(n7061));
INVX1    g1453(.A(WX4664), .Y(n7062));
XOR2X1   g1454(.A(WX4728), .B(n7062), .Y(n7063));
XOR2X1   g1455(.A(n7063), .B(n7061), .Y(n7064_1));
MX2X1    g1456(.A(n7059_1), .B(n7064_1), .S0(n5539), .Y(n7066));
INVX1    g1457(.A(WX3083), .Y(n7067));
MX2X1    g1458(.A(n7067), .B(n6485), .S0(n5539), .Y(n7068));
MX2X1    g1459(.A(n7066), .B(n7068), .S0(TM1), .Y(n7069_1));
NOR2X1   g1460(.A(n7069_1), .B(n5827), .Y(n2757));
INVX1    g1461(.A(CRC_OUT_7_24), .Y(n7071));
XOR2X1   g1462(.A(WX4538), .B(TM1), .Y(n7072));
XOR2X1   g1463(.A(n7072), .B(WX4602), .Y(n7073));
INVX1    g1464(.A(WX4666), .Y(n7074_1));
XOR2X1   g1465(.A(WX4730), .B(n7074_1), .Y(n7075));
XOR2X1   g1466(.A(n7075), .B(n7073), .Y(n7076));
MX2X1    g1467(.A(n7071), .B(n7076), .S0(n5539), .Y(n7078));
INVX1    g1468(.A(WX3085), .Y(n7079_1));
MX2X1    g1469(.A(n7079_1), .B(n6497), .S0(n5539), .Y(n7080));
MX2X1    g1470(.A(n7078), .B(n7080), .S0(TM1), .Y(n7081));
NOR2X1   g1471(.A(n7081), .B(n5827), .Y(n2762));
INVX1    g1472(.A(CRC_OUT_7_23), .Y(n7083_1));
XOR2X1   g1473(.A(WX4540), .B(TM1), .Y(n7084));
XOR2X1   g1474(.A(n7084), .B(WX4604), .Y(n7085));
INVX1    g1475(.A(WX4668), .Y(n7086));
XOR2X1   g1476(.A(WX4732), .B(n7086), .Y(n7087_1));
XOR2X1   g1477(.A(n7087_1), .B(n7085), .Y(n7088));
MX2X1    g1478(.A(n7083_1), .B(n7088), .S0(n5539), .Y(n7090));
INVX1    g1479(.A(WX3087), .Y(n7091_1));
MX2X1    g1480(.A(n7091_1), .B(n6509_1), .S0(n5539), .Y(n7092));
MX2X1    g1481(.A(n7090), .B(n7092), .S0(TM1), .Y(n7093));
NOR2X1   g1482(.A(n7093), .B(n5827), .Y(n2767));
INVX1    g1483(.A(CRC_OUT_7_22), .Y(n7095_1));
XOR2X1   g1484(.A(WX4542), .B(TM1), .Y(n7096));
XOR2X1   g1485(.A(n7096), .B(WX4606), .Y(n7097));
INVX1    g1486(.A(WX4670), .Y(n7098));
XOR2X1   g1487(.A(WX4734), .B(n7098), .Y(n7099_1));
XOR2X1   g1488(.A(n7099_1), .B(n7097), .Y(n7100));
MX2X1    g1489(.A(n7095_1), .B(n7100), .S0(n5539), .Y(n7102));
INVX1    g1490(.A(WX3089), .Y(n7103_1));
MX2X1    g1491(.A(n7103_1), .B(n6521), .S0(n5539), .Y(n7104));
MX2X1    g1492(.A(n7102), .B(n7104), .S0(TM1), .Y(n7105));
NOR2X1   g1493(.A(n7105), .B(n5827), .Y(n2772));
INVX1    g1494(.A(CRC_OUT_7_21), .Y(n7107_1));
XOR2X1   g1495(.A(WX4544), .B(TM1), .Y(n7108));
XOR2X1   g1496(.A(n7108), .B(WX4608), .Y(n7109));
INVX1    g1497(.A(WX4672), .Y(n7110));
XOR2X1   g1498(.A(WX4736), .B(n7110), .Y(n7111_1));
XOR2X1   g1499(.A(n7111_1), .B(n7109), .Y(n7112));
MX2X1    g1500(.A(n7107_1), .B(n7112), .S0(n5539), .Y(n7114));
INVX1    g1501(.A(WX3091), .Y(n7115_1));
MX2X1    g1502(.A(n7115_1), .B(n6533), .S0(n5539), .Y(n7116));
MX2X1    g1503(.A(n7114), .B(n7116), .S0(TM1), .Y(n7117));
NOR2X1   g1504(.A(n7117), .B(n5827), .Y(n2777));
INVX1    g1505(.A(CRC_OUT_7_20), .Y(n7119_1));
XOR2X1   g1506(.A(WX4546), .B(TM1), .Y(n7120));
XOR2X1   g1507(.A(n7120), .B(WX4610), .Y(n7121));
INVX1    g1508(.A(WX4674), .Y(n7122));
XOR2X1   g1509(.A(WX4738), .B(n7122), .Y(n7123_1));
XOR2X1   g1510(.A(n7123_1), .B(n7121), .Y(n7124));
MX2X1    g1511(.A(n7119_1), .B(n7124), .S0(n5539), .Y(n7126));
INVX1    g1512(.A(WX3093), .Y(n7127_1));
MX2X1    g1513(.A(n7127_1), .B(n6545), .S0(n5539), .Y(n7128));
MX2X1    g1514(.A(n7126), .B(n7128), .S0(TM1), .Y(n7129));
NOR2X1   g1515(.A(n7129), .B(n5827), .Y(n2782));
INVX1    g1516(.A(CRC_OUT_7_19), .Y(n7131_1));
XOR2X1   g1517(.A(WX4548), .B(TM1), .Y(n7132));
XOR2X1   g1518(.A(n7132), .B(WX4612), .Y(n7133));
INVX1    g1519(.A(WX4676), .Y(n7134));
XOR2X1   g1520(.A(WX4740), .B(n7134), .Y(n7135_1));
XOR2X1   g1521(.A(n7135_1), .B(n7133), .Y(n7136));
MX2X1    g1522(.A(n7131_1), .B(n7136), .S0(n5539), .Y(n7138));
INVX1    g1523(.A(WX3095), .Y(n7139_1));
MX2X1    g1524(.A(n7139_1), .B(n6557), .S0(n5539), .Y(n7140));
MX2X1    g1525(.A(n7138), .B(n7140), .S0(TM1), .Y(n7141));
NOR2X1   g1526(.A(n7141), .B(n5827), .Y(n2787));
INVX1    g1527(.A(CRC_OUT_7_18), .Y(n7143_1));
XOR2X1   g1528(.A(WX4550), .B(TM1), .Y(n7144));
XOR2X1   g1529(.A(n7144), .B(WX4614), .Y(n7145));
INVX1    g1530(.A(WX4678), .Y(n7146));
XOR2X1   g1531(.A(WX4742), .B(n7146), .Y(n7147_1));
XOR2X1   g1532(.A(n7147_1), .B(n7145), .Y(n7148));
MX2X1    g1533(.A(n7143_1), .B(n7148), .S0(n5539), .Y(n7150));
INVX1    g1534(.A(WX3097), .Y(n7151_1));
MX2X1    g1535(.A(n7151_1), .B(n6569_1), .S0(n5539), .Y(n7152));
MX2X1    g1536(.A(n7150), .B(n7152), .S0(TM1), .Y(n7153));
NOR2X1   g1537(.A(n7153), .B(n5827), .Y(n2792));
INVX1    g1538(.A(CRC_OUT_7_17), .Y(n7155_1));
XOR2X1   g1539(.A(WX4552), .B(TM1), .Y(n7156));
XOR2X1   g1540(.A(n7156), .B(WX4616), .Y(n7157));
INVX1    g1541(.A(WX4680), .Y(n7158));
XOR2X1   g1542(.A(WX4744), .B(n7158), .Y(n7159_1));
XOR2X1   g1543(.A(n7159_1), .B(n7157), .Y(n7160));
MX2X1    g1544(.A(n7155_1), .B(n7160), .S0(n5539), .Y(n7162));
INVX1    g1545(.A(WX3099), .Y(n7163_1));
MX2X1    g1546(.A(n7163_1), .B(n6581), .S0(n5539), .Y(n7164));
MX2X1    g1547(.A(n7162), .B(n7164), .S0(TM1), .Y(n7165));
NOR2X1   g1548(.A(n7165), .B(n5827), .Y(n2797));
INVX1    g1549(.A(CRC_OUT_7_16), .Y(n7167_1));
XOR2X1   g1550(.A(WX4554), .B(TM1), .Y(n7168));
XOR2X1   g1551(.A(n7168), .B(WX4618), .Y(n7169));
INVX1    g1552(.A(WX4682), .Y(n7170));
XOR2X1   g1553(.A(WX4746), .B(n7170), .Y(n7171_1));
XOR2X1   g1554(.A(n7171_1), .B(n7169), .Y(n7172));
MX2X1    g1555(.A(n7167_1), .B(n7172), .S0(n5539), .Y(n7174));
INVX1    g1556(.A(WX3101), .Y(n7175_1));
MX2X1    g1557(.A(n7175_1), .B(n6593), .S0(n5539), .Y(n7176));
MX2X1    g1558(.A(n7174), .B(n7176), .S0(TM1), .Y(n7177));
NOR2X1   g1559(.A(n7177), .B(n5827), .Y(n2802));
INVX1    g1560(.A(CRC_OUT_7_15), .Y(n7179_1));
XOR2X1   g1561(.A(WX4556), .B(TM0), .Y(n7180));
XOR2X1   g1562(.A(n7180), .B(WX4620), .Y(n7181));
INVX1    g1563(.A(WX4684), .Y(n7182));
XOR2X1   g1564(.A(WX4748), .B(n7182), .Y(n7183_1));
XOR2X1   g1565(.A(n7183_1), .B(n7181), .Y(n7184));
MX2X1    g1566(.A(n7179_1), .B(n7184), .S0(n5539), .Y(n7186));
INVX1    g1567(.A(WX3103), .Y(n7187_1));
MX2X1    g1568(.A(n7187_1), .B(n6605), .S0(n5539), .Y(n7188));
MX2X1    g1569(.A(n7186), .B(n7188), .S0(TM1), .Y(n7189));
NOR2X1   g1570(.A(n7189), .B(n5827), .Y(n2807));
INVX1    g1571(.A(CRC_OUT_7_14), .Y(n7191_1));
XOR2X1   g1572(.A(WX4558), .B(TM0), .Y(n7192));
XOR2X1   g1573(.A(n7192), .B(WX4622), .Y(n7193));
INVX1    g1574(.A(WX4686), .Y(n7194));
XOR2X1   g1575(.A(WX4750), .B(n7194), .Y(n7195_1));
XOR2X1   g1576(.A(n7195_1), .B(n7193), .Y(n7196));
MX2X1    g1577(.A(n7191_1), .B(n7196), .S0(n5539), .Y(n7198));
INVX1    g1578(.A(WX3105), .Y(n7199_1));
MX2X1    g1579(.A(n7199_1), .B(n6617), .S0(n5539), .Y(n7200));
MX2X1    g1580(.A(n7198), .B(n7200), .S0(TM1), .Y(n7201));
NOR2X1   g1581(.A(n7201), .B(n5827), .Y(n2812));
INVX1    g1582(.A(CRC_OUT_7_13), .Y(n7203_1));
XOR2X1   g1583(.A(WX4560), .B(TM0), .Y(n7204));
XOR2X1   g1584(.A(n7204), .B(WX4624), .Y(n7205));
INVX1    g1585(.A(WX4688), .Y(n7206));
XOR2X1   g1586(.A(WX4752), .B(n7206), .Y(n7207_1));
XOR2X1   g1587(.A(n7207_1), .B(n7205), .Y(n7208));
MX2X1    g1588(.A(n7203_1), .B(n7208), .S0(n5539), .Y(n7210));
INVX1    g1589(.A(WX3107), .Y(n7211));
MX2X1    g1590(.A(n7211), .B(n6629_1), .S0(n5539), .Y(n7212_1));
MX2X1    g1591(.A(n7210), .B(n7212_1), .S0(TM1), .Y(n7213));
NOR2X1   g1592(.A(n7213), .B(n5827), .Y(n2817));
INVX1    g1593(.A(CRC_OUT_7_12), .Y(n7215));
XOR2X1   g1594(.A(WX4562), .B(TM0), .Y(n7216));
XOR2X1   g1595(.A(n7216), .B(WX4626), .Y(n7217_1));
INVX1    g1596(.A(WX4690), .Y(n7218));
XOR2X1   g1597(.A(WX4754), .B(n7218), .Y(n7219));
XOR2X1   g1598(.A(n7219), .B(n7217_1), .Y(n7220));
MX2X1    g1599(.A(n7215), .B(n7220), .S0(n5539), .Y(n7222_1));
INVX1    g1600(.A(WX3109), .Y(n7223));
MX2X1    g1601(.A(n7223), .B(n6641), .S0(n5539), .Y(n7224));
MX2X1    g1602(.A(n7222_1), .B(n7224), .S0(TM1), .Y(n7225));
NOR2X1   g1603(.A(n7225), .B(n5827), .Y(n2822));
INVX1    g1604(.A(CRC_OUT_7_11), .Y(n7227_1));
XOR2X1   g1605(.A(WX4564), .B(TM0), .Y(n7228));
XOR2X1   g1606(.A(n7228), .B(WX4628), .Y(n7229));
INVX1    g1607(.A(WX4692), .Y(n7230));
XOR2X1   g1608(.A(WX4756), .B(n7230), .Y(n7231));
XOR2X1   g1609(.A(n7231), .B(n7229), .Y(n7232_1));
MX2X1    g1610(.A(n7227_1), .B(n7232_1), .S0(n5539), .Y(n7234));
INVX1    g1611(.A(WX3111), .Y(n7235));
MX2X1    g1612(.A(n7235), .B(n6653), .S0(n5539), .Y(n7236));
MX2X1    g1613(.A(n7234), .B(n7236), .S0(TM1), .Y(n7237_1));
NOR2X1   g1614(.A(n7237_1), .B(n5827), .Y(n2827));
INVX1    g1615(.A(CRC_OUT_7_10), .Y(n7239));
XOR2X1   g1616(.A(WX4566), .B(TM0), .Y(n7240));
XOR2X1   g1617(.A(n7240), .B(WX4630), .Y(n7241));
INVX1    g1618(.A(WX4694), .Y(n7242_1));
XOR2X1   g1619(.A(WX4758), .B(n7242_1), .Y(n7243));
XOR2X1   g1620(.A(n7243), .B(n7241), .Y(n7244));
MX2X1    g1621(.A(n7239), .B(n7244), .S0(n5539), .Y(n7246));
INVX1    g1622(.A(WX3113), .Y(n7247_1));
MX2X1    g1623(.A(n7247_1), .B(n6665), .S0(n5539), .Y(n7248));
MX2X1    g1624(.A(n7246), .B(n7248), .S0(TM1), .Y(n7249));
NOR2X1   g1625(.A(n7249), .B(n5827), .Y(n2832));
INVX1    g1626(.A(CRC_OUT_7_9), .Y(n7251));
XOR2X1   g1627(.A(WX4568), .B(TM0), .Y(n7252_1));
XOR2X1   g1628(.A(n7252_1), .B(WX4632), .Y(n7253));
INVX1    g1629(.A(WX4696), .Y(n7254));
XOR2X1   g1630(.A(WX4760), .B(n7254), .Y(n7255));
XOR2X1   g1631(.A(n7255), .B(n7253), .Y(n7256));
MX2X1    g1632(.A(n7251), .B(n7256), .S0(n5539), .Y(n7258));
INVX1    g1633(.A(WX3115), .Y(n7259));
MX2X1    g1634(.A(n7259), .B(n6677), .S0(n5539), .Y(n7260));
MX2X1    g1635(.A(n7258), .B(n7260), .S0(TM1), .Y(n7261));
NOR2X1   g1636(.A(n7261), .B(n5827), .Y(n2837));
INVX1    g1637(.A(CRC_OUT_7_8), .Y(n7263));
XOR2X1   g1638(.A(WX4570), .B(TM0), .Y(n7264));
XOR2X1   g1639(.A(n7264), .B(WX4634), .Y(n7265));
INVX1    g1640(.A(WX4698), .Y(n7266));
XOR2X1   g1641(.A(WX4762), .B(n7266), .Y(n7267_1));
XOR2X1   g1642(.A(n7267_1), .B(n7265), .Y(n7268));
MX2X1    g1643(.A(n7263), .B(n7268), .S0(n5539), .Y(n7270));
INVX1    g1644(.A(WX3117), .Y(n7271));
MX2X1    g1645(.A(n7271), .B(n6689_1), .S0(n5539), .Y(n7272_1));
MX2X1    g1646(.A(n7270), .B(n7272_1), .S0(TM1), .Y(n7273));
NOR2X1   g1647(.A(n7273), .B(n5827), .Y(n2842));
INVX1    g1648(.A(CRC_OUT_7_7), .Y(n7275));
XOR2X1   g1649(.A(WX4572), .B(TM0), .Y(n7276));
XOR2X1   g1650(.A(n7276), .B(WX4636), .Y(n7277_1));
INVX1    g1651(.A(WX4700), .Y(n7278));
XOR2X1   g1652(.A(WX4764), .B(n7278), .Y(n7279));
XOR2X1   g1653(.A(n7279), .B(n7277_1), .Y(n7280));
MX2X1    g1654(.A(n7275), .B(n7280), .S0(n5539), .Y(n7282_1));
INVX1    g1655(.A(WX3119), .Y(n7283));
MX2X1    g1656(.A(n7283), .B(n6701), .S0(n5539), .Y(n7284));
MX2X1    g1657(.A(n7282_1), .B(n7284), .S0(TM1), .Y(n7285));
NOR2X1   g1658(.A(n7285), .B(n5827), .Y(n2847));
INVX1    g1659(.A(CRC_OUT_7_6), .Y(n7287_1));
XOR2X1   g1660(.A(WX4574), .B(TM0), .Y(n7288));
XOR2X1   g1661(.A(n7288), .B(WX4638), .Y(n7289));
INVX1    g1662(.A(WX4702), .Y(n7290));
XOR2X1   g1663(.A(WX4766), .B(n7290), .Y(n7291));
XOR2X1   g1664(.A(n7291), .B(n7289), .Y(n7292_1));
MX2X1    g1665(.A(n7287_1), .B(n7292_1), .S0(n5539), .Y(n7294));
INVX1    g1666(.A(WX3121), .Y(n7295));
MX2X1    g1667(.A(n7295), .B(n6713), .S0(n5539), .Y(n7296));
MX2X1    g1668(.A(n7294), .B(n7296), .S0(TM1), .Y(n7297_1));
NOR2X1   g1669(.A(n7297_1), .B(n5827), .Y(n2852));
INVX1    g1670(.A(CRC_OUT_7_5), .Y(n7299));
XOR2X1   g1671(.A(WX4576), .B(TM0), .Y(n7300));
XOR2X1   g1672(.A(n7300), .B(WX4640), .Y(n7301));
INVX1    g1673(.A(WX4704), .Y(n7302_1));
XOR2X1   g1674(.A(WX4768), .B(n7302_1), .Y(n7303));
XOR2X1   g1675(.A(n7303), .B(n7301), .Y(n7304));
MX2X1    g1676(.A(n7299), .B(n7304), .S0(n5539), .Y(n7306));
INVX1    g1677(.A(WX3123), .Y(n7307_1));
MX2X1    g1678(.A(n7307_1), .B(n6725), .S0(n5539), .Y(n7308));
MX2X1    g1679(.A(n7306), .B(n7308), .S0(TM1), .Y(n7309));
NOR2X1   g1680(.A(n7309), .B(n5827), .Y(n2857));
INVX1    g1681(.A(CRC_OUT_7_4), .Y(n7311));
XOR2X1   g1682(.A(WX4578), .B(TM0), .Y(n7312_1));
XOR2X1   g1683(.A(n7312_1), .B(WX4642), .Y(n7313));
INVX1    g1684(.A(WX4706), .Y(n7314));
XOR2X1   g1685(.A(WX4770), .B(n7314), .Y(n7315));
XOR2X1   g1686(.A(n7315), .B(n7313), .Y(n7316));
MX2X1    g1687(.A(n7311), .B(n7316), .S0(n5539), .Y(n7318));
INVX1    g1688(.A(WX3125), .Y(n7319));
MX2X1    g1689(.A(n7319), .B(n6737), .S0(n5539), .Y(n7320));
MX2X1    g1690(.A(n7318), .B(n7320), .S0(TM1), .Y(n7321));
NOR2X1   g1691(.A(n7321), .B(n5827), .Y(n2862));
INVX1    g1692(.A(CRC_OUT_7_3), .Y(n7323));
XOR2X1   g1693(.A(WX4580), .B(TM0), .Y(n7324));
XOR2X1   g1694(.A(n7324), .B(WX4644), .Y(n7325));
INVX1    g1695(.A(WX4708), .Y(n7326));
XOR2X1   g1696(.A(WX4772), .B(n7326), .Y(n7327_1));
XOR2X1   g1697(.A(n7327_1), .B(n7325), .Y(n7328));
MX2X1    g1698(.A(n7323), .B(n7328), .S0(n5539), .Y(n7330));
INVX1    g1699(.A(WX3127), .Y(n7331));
MX2X1    g1700(.A(n7331), .B(n6749_1), .S0(n5539), .Y(n7332_1));
MX2X1    g1701(.A(n7330), .B(n7332_1), .S0(TM1), .Y(n7333));
NOR2X1   g1702(.A(n7333), .B(n5827), .Y(n2867));
INVX1    g1703(.A(CRC_OUT_7_2), .Y(n7335));
XOR2X1   g1704(.A(WX4582), .B(TM0), .Y(n7336));
XOR2X1   g1705(.A(n7336), .B(WX4646), .Y(n7337_1));
INVX1    g1706(.A(WX4710), .Y(n7338));
XOR2X1   g1707(.A(WX4774), .B(n7338), .Y(n7339));
XOR2X1   g1708(.A(n7339), .B(n7337_1), .Y(n7340));
MX2X1    g1709(.A(n7335), .B(n7340), .S0(n5539), .Y(n7342_1));
INVX1    g1710(.A(WX3129), .Y(n7343));
MX2X1    g1711(.A(n7343), .B(n6761), .S0(n5539), .Y(n7344));
MX2X1    g1712(.A(n7342_1), .B(n7344), .S0(TM1), .Y(n7345));
NOR2X1   g1713(.A(n7345), .B(n5827), .Y(n2872));
INVX1    g1714(.A(CRC_OUT_7_1), .Y(n7347_1));
XOR2X1   g1715(.A(WX4584), .B(TM0), .Y(n7348));
XOR2X1   g1716(.A(n7348), .B(WX4648), .Y(n7349));
INVX1    g1717(.A(WX4712), .Y(n7350));
XOR2X1   g1718(.A(WX4776), .B(n7350), .Y(n7351));
XOR2X1   g1719(.A(n7351), .B(n7349), .Y(n7352_1));
MX2X1    g1720(.A(n7347_1), .B(n7352_1), .S0(n5539), .Y(n7354));
INVX1    g1721(.A(WX3131), .Y(n7355));
MX2X1    g1722(.A(n7355), .B(n6773), .S0(n5539), .Y(n7356));
MX2X1    g1723(.A(n7354), .B(n7356), .S0(TM1), .Y(n7357_1));
NOR2X1   g1724(.A(n7357_1), .B(n5827), .Y(n2877));
INVX1    g1725(.A(CRC_OUT_7_0), .Y(n7359));
XOR2X1   g1726(.A(WX4586), .B(TM0), .Y(n7360));
XOR2X1   g1727(.A(n7360), .B(WX4650), .Y(n7361));
INVX1    g1728(.A(WX4714), .Y(n7362_1));
XOR2X1   g1729(.A(WX4778), .B(n7362_1), .Y(n7363));
XOR2X1   g1730(.A(n7363), .B(n7361), .Y(n7364));
MX2X1    g1731(.A(n7359), .B(n7364), .S0(n5539), .Y(n7366));
INVX1    g1732(.A(WX3133), .Y(n7367_1));
MX2X1    g1733(.A(n7367_1), .B(n6785), .S0(n5539), .Y(n7368));
MX2X1    g1734(.A(n7366), .B(n7368), .S0(TM1), .Y(n7369));
NOR2X1   g1735(.A(n7369), .B(n5827), .Y(n2882));
AND2X1   g1736(.A(WX3231), .B(RESET), .Y(n2887));
AND2X1   g1737(.A(WX3233), .B(RESET), .Y(n2892));
AND2X1   g1738(.A(WX3235), .B(RESET), .Y(n2897));
AND2X1   g1739(.A(WX3237), .B(RESET), .Y(n2902));
AND2X1   g1740(.A(WX3239), .B(RESET), .Y(n2907));
AND2X1   g1741(.A(WX3241), .B(RESET), .Y(n2912));
AND2X1   g1742(.A(WX3243), .B(RESET), .Y(n2917));
AND2X1   g1743(.A(WX3245), .B(RESET), .Y(n2922));
AND2X1   g1744(.A(WX3247), .B(RESET), .Y(n2927));
AND2X1   g1745(.A(WX3249), .B(RESET), .Y(n2932));
AND2X1   g1746(.A(WX3251), .B(RESET), .Y(n2937));
AND2X1   g1747(.A(WX3253), .B(RESET), .Y(n2942));
AND2X1   g1748(.A(WX3255), .B(RESET), .Y(n2947));
AND2X1   g1749(.A(WX3257), .B(RESET), .Y(n2952));
AND2X1   g1750(.A(WX3259), .B(RESET), .Y(n2957));
AND2X1   g1751(.A(WX3261), .B(RESET), .Y(n2962));
AND2X1   g1752(.A(WX3263), .B(RESET), .Y(n2967));
AND2X1   g1753(.A(WX3265), .B(RESET), .Y(n2972));
AND2X1   g1754(.A(WX3267), .B(RESET), .Y(n2977));
AND2X1   g1755(.A(WX3269), .B(RESET), .Y(n2982));
AND2X1   g1756(.A(WX3271), .B(RESET), .Y(n2987));
AND2X1   g1757(.A(WX3273), .B(RESET), .Y(n2992));
AND2X1   g1758(.A(WX3275), .B(RESET), .Y(n2997));
AND2X1   g1759(.A(WX3277), .B(RESET), .Y(n3002));
AND2X1   g1760(.A(WX3279), .B(RESET), .Y(n3007));
AND2X1   g1761(.A(WX3281), .B(RESET), .Y(n3012));
AND2X1   g1762(.A(WX3283), .B(RESET), .Y(n3017));
AND2X1   g1763(.A(WX3285), .B(RESET), .Y(n3022));
AND2X1   g1764(.A(WX3287), .B(RESET), .Y(n3027));
AND2X1   g1765(.A(WX3289), .B(RESET), .Y(n3032));
AND2X1   g1766(.A(WX3291), .B(RESET), .Y(n3037));
AND2X1   g1767(.A(WX3293), .B(RESET), .Y(n3042));
AND2X1   g1768(.A(WX3295), .B(RESET), .Y(n3047));
AND2X1   g1769(.A(WX3297), .B(RESET), .Y(n3052));
AND2X1   g1770(.A(WX3299), .B(RESET), .Y(n3057));
AND2X1   g1771(.A(WX3301), .B(RESET), .Y(n3062));
AND2X1   g1772(.A(WX3303), .B(RESET), .Y(n3067));
AND2X1   g1773(.A(WX3305), .B(RESET), .Y(n3072));
AND2X1   g1774(.A(WX3307), .B(RESET), .Y(n3077));
AND2X1   g1775(.A(WX3309), .B(RESET), .Y(n3082));
AND2X1   g1776(.A(WX3311), .B(RESET), .Y(n3087));
AND2X1   g1777(.A(WX3313), .B(RESET), .Y(n3092));
AND2X1   g1778(.A(WX3315), .B(RESET), .Y(n3097));
AND2X1   g1779(.A(WX3317), .B(RESET), .Y(n3102));
AND2X1   g1780(.A(WX3319), .B(RESET), .Y(n3107));
AND2X1   g1781(.A(WX3321), .B(RESET), .Y(n3112));
AND2X1   g1782(.A(WX3323), .B(RESET), .Y(n3117));
AND2X1   g1783(.A(WX3325), .B(RESET), .Y(n3122));
AND2X1   g1784(.A(WX3327), .B(RESET), .Y(n3127));
AND2X1   g1785(.A(WX3329), .B(RESET), .Y(n3132));
AND2X1   g1786(.A(WX3331), .B(RESET), .Y(n3137));
AND2X1   g1787(.A(WX3333), .B(RESET), .Y(n3142));
AND2X1   g1788(.A(WX3335), .B(RESET), .Y(n3147));
AND2X1   g1789(.A(WX3337), .B(RESET), .Y(n3152));
AND2X1   g1790(.A(WX3339), .B(RESET), .Y(n3157));
AND2X1   g1791(.A(WX3341), .B(RESET), .Y(n3162));
AND2X1   g1792(.A(WX3343), .B(RESET), .Y(n3167));
AND2X1   g1793(.A(WX3345), .B(RESET), .Y(n3172));
AND2X1   g1794(.A(WX3347), .B(RESET), .Y(n3177));
AND2X1   g1795(.A(WX3349), .B(RESET), .Y(n3182));
AND2X1   g1796(.A(WX3351), .B(RESET), .Y(n3187));
AND2X1   g1797(.A(WX3353), .B(RESET), .Y(n3192));
AND2X1   g1798(.A(WX3355), .B(RESET), .Y(n3197));
AND2X1   g1799(.A(WX3357), .B(RESET), .Y(n3202));
AND2X1   g1800(.A(WX3359), .B(RESET), .Y(n3207));
AND2X1   g1801(.A(WX3361), .B(RESET), .Y(n3212));
AND2X1   g1802(.A(WX3363), .B(RESET), .Y(n3217));
AND2X1   g1803(.A(WX3365), .B(RESET), .Y(n3222));
AND2X1   g1804(.A(WX3367), .B(RESET), .Y(n3227));
AND2X1   g1805(.A(WX3369), .B(RESET), .Y(n3232));
AND2X1   g1806(.A(WX3371), .B(RESET), .Y(n3237));
AND2X1   g1807(.A(WX3373), .B(RESET), .Y(n3242));
AND2X1   g1808(.A(WX3375), .B(RESET), .Y(n3247));
AND2X1   g1809(.A(WX3377), .B(RESET), .Y(n3252));
AND2X1   g1810(.A(WX3379), .B(RESET), .Y(n3257));
AND2X1   g1811(.A(WX3381), .B(RESET), .Y(n3262));
AND2X1   g1812(.A(WX3383), .B(RESET), .Y(n3267));
AND2X1   g1813(.A(WX3385), .B(RESET), .Y(n3272));
AND2X1   g1814(.A(WX3387), .B(RESET), .Y(n3277));
AND2X1   g1815(.A(WX3389), .B(RESET), .Y(n3282));
AND2X1   g1816(.A(WX3391), .B(RESET), .Y(n3287));
AND2X1   g1817(.A(WX3393), .B(RESET), .Y(n3292));
AND2X1   g1818(.A(WX3395), .B(RESET), .Y(n3297));
AND2X1   g1819(.A(WX3397), .B(RESET), .Y(n3302));
AND2X1   g1820(.A(WX3399), .B(RESET), .Y(n3307));
AND2X1   g1821(.A(WX3401), .B(RESET), .Y(n3312));
AND2X1   g1822(.A(WX3403), .B(RESET), .Y(n3317));
AND2X1   g1823(.A(WX3405), .B(RESET), .Y(n3322));
AND2X1   g1824(.A(WX3407), .B(RESET), .Y(n3327));
AND2X1   g1825(.A(WX3409), .B(RESET), .Y(n3332));
AND2X1   g1826(.A(WX3411), .B(RESET), .Y(n3337));
AND2X1   g1827(.A(WX3413), .B(RESET), .Y(n3342));
AND2X1   g1828(.A(WX3415), .B(RESET), .Y(n3347));
AND2X1   g1829(.A(WX3417), .B(RESET), .Y(n3352));
AND2X1   g1830(.A(WX3419), .B(RESET), .Y(n3357));
AND2X1   g1831(.A(WX3421), .B(RESET), .Y(n3362));
XOR2X1   g1832(.A(CRC_OUT_7_31), .B(WX3485), .Y(n7467_1));
NOR2X1   g1833(.A(n7467_1), .B(n5827), .Y(CRC_OUT_7_0));
XOR2X1   g1834(.A(CRC_OUT_7_0), .B(WX3483), .Y(n7469));
NOR2X1   g1835(.A(n7469), .B(n5827), .Y(CRC_OUT_7_1));
XOR2X1   g1836(.A(CRC_OUT_7_1), .B(WX3481), .Y(n7471));
NOR2X1   g1837(.A(n7471), .B(n5827), .Y(CRC_OUT_7_2));
XOR2X1   g1838(.A(CRC_OUT_7_2), .B(WX3479), .Y(n7473));
NOR2X1   g1839(.A(n7473), .B(n5827), .Y(CRC_OUT_7_3));
XOR2X1   g1840(.A(CRC_OUT_7_31), .B(WX3477), .Y(n7475));
XOR2X1   g1841(.A(n7475), .B(CRC_OUT_7_3), .Y(n7476));
NOR2X1   g1842(.A(n7476), .B(n5827), .Y(CRC_OUT_7_4));
XOR2X1   g1843(.A(CRC_OUT_7_4), .B(WX3475), .Y(n7478));
NOR2X1   g1844(.A(n7478), .B(n5827), .Y(CRC_OUT_7_5));
XOR2X1   g1845(.A(CRC_OUT_7_5), .B(WX3473), .Y(n7480));
NOR2X1   g1846(.A(n7480), .B(n5827), .Y(CRC_OUT_7_6));
XOR2X1   g1847(.A(CRC_OUT_7_6), .B(WX3471), .Y(n7482_1));
NOR2X1   g1848(.A(n7482_1), .B(n5827), .Y(CRC_OUT_7_7));
XOR2X1   g1849(.A(CRC_OUT_7_7), .B(WX3469), .Y(n7484));
NOR2X1   g1850(.A(n7484), .B(n5827), .Y(CRC_OUT_7_8));
XOR2X1   g1851(.A(CRC_OUT_7_8), .B(WX3467), .Y(n7486));
NOR2X1   g1852(.A(n7486), .B(n5827), .Y(CRC_OUT_7_9));
XOR2X1   g1853(.A(CRC_OUT_7_9), .B(WX3465), .Y(n7488));
NOR2X1   g1854(.A(n7488), .B(n5827), .Y(CRC_OUT_7_10));
XOR2X1   g1855(.A(CRC_OUT_7_31), .B(WX3463), .Y(n7490));
XOR2X1   g1856(.A(n7490), .B(CRC_OUT_7_10), .Y(n7491));
NOR2X1   g1857(.A(n7491), .B(n5827), .Y(CRC_OUT_7_11));
XOR2X1   g1858(.A(CRC_OUT_7_11), .B(WX3461), .Y(n7493));
NOR2X1   g1859(.A(n7493), .B(n5827), .Y(CRC_OUT_7_12));
XOR2X1   g1860(.A(CRC_OUT_7_12), .B(WX3459), .Y(n7495));
NOR2X1   g1861(.A(n7495), .B(n5827), .Y(CRC_OUT_7_13));
XOR2X1   g1862(.A(CRC_OUT_7_13), .B(WX3457), .Y(n7497_1));
NOR2X1   g1863(.A(n7497_1), .B(n5827), .Y(CRC_OUT_7_14));
XOR2X1   g1864(.A(CRC_OUT_7_14), .B(WX3455), .Y(n7499));
NOR2X1   g1865(.A(n7499), .B(n5827), .Y(CRC_OUT_7_15));
XOR2X1   g1866(.A(CRC_OUT_7_31), .B(WX3453), .Y(n7501));
XOR2X1   g1867(.A(n7501), .B(CRC_OUT_7_15), .Y(n7502_1));
NOR2X1   g1868(.A(n7502_1), .B(n5827), .Y(CRC_OUT_7_16));
XOR2X1   g1869(.A(CRC_OUT_7_16), .B(WX3451), .Y(n7504));
NOR2X1   g1870(.A(n7504), .B(n5827), .Y(CRC_OUT_7_17));
XOR2X1   g1871(.A(CRC_OUT_7_17), .B(WX3449), .Y(n7506));
NOR2X1   g1872(.A(n7506), .B(n5827), .Y(CRC_OUT_7_18));
XOR2X1   g1873(.A(CRC_OUT_7_18), .B(WX3447), .Y(n7508));
NOR2X1   g1874(.A(n7508), .B(n5827), .Y(CRC_OUT_7_19));
XOR2X1   g1875(.A(CRC_OUT_7_19), .B(WX3445), .Y(n7510));
NOR2X1   g1876(.A(n7510), .B(n5827), .Y(CRC_OUT_7_20));
XOR2X1   g1877(.A(CRC_OUT_7_20), .B(WX3443), .Y(n7512_1));
NOR2X1   g1878(.A(n7512_1), .B(n5827), .Y(CRC_OUT_7_21));
XOR2X1   g1879(.A(CRC_OUT_7_21), .B(WX3441), .Y(n7514));
NOR2X1   g1880(.A(n7514), .B(n5827), .Y(CRC_OUT_7_22));
XOR2X1   g1881(.A(CRC_OUT_7_22), .B(WX3439), .Y(n7516));
NOR2X1   g1882(.A(n7516), .B(n5827), .Y(CRC_OUT_7_23));
XOR2X1   g1883(.A(CRC_OUT_7_23), .B(WX3437), .Y(n7518));
NOR2X1   g1884(.A(n7518), .B(n5827), .Y(CRC_OUT_7_24));
XOR2X1   g1885(.A(CRC_OUT_7_24), .B(WX3435), .Y(n7520));
NOR2X1   g1886(.A(n7520), .B(n5827), .Y(CRC_OUT_7_25));
XOR2X1   g1887(.A(CRC_OUT_7_25), .B(WX3433), .Y(n7522_1));
NOR2X1   g1888(.A(n7522_1), .B(n5827), .Y(CRC_OUT_7_26));
XOR2X1   g1889(.A(CRC_OUT_7_26), .B(WX3431), .Y(n7524));
NOR2X1   g1890(.A(n7524), .B(n5827), .Y(CRC_OUT_7_27));
XOR2X1   g1891(.A(CRC_OUT_7_27), .B(WX3429), .Y(n7526));
NOR2X1   g1892(.A(n7526), .B(n5827), .Y(CRC_OUT_7_28));
XOR2X1   g1893(.A(CRC_OUT_7_28), .B(WX3427), .Y(n7528));
NOR2X1   g1894(.A(n7528), .B(n5827), .Y(CRC_OUT_7_29));
XOR2X1   g1895(.A(CRC_OUT_7_29), .B(WX3425), .Y(n7530));
NOR2X1   g1896(.A(n7530), .B(n5827), .Y(CRC_OUT_7_30));
XOR2X1   g1897(.A(CRC_OUT_7_30), .B(WX3423), .Y(n7532_1));
NOR2X1   g1898(.A(n7532_1), .B(n5827), .Y(CRC_OUT_7_31));
AND2X1   g1899(.A(WX4366), .B(RESET), .Y(n3495));
AND2X1   g1900(.A(WX4368), .B(RESET), .Y(n3500));
AND2X1   g1901(.A(WX4370), .B(RESET), .Y(n3505));
AND2X1   g1902(.A(WX4372), .B(RESET), .Y(n3510));
AND2X1   g1903(.A(WX4374), .B(RESET), .Y(n3515));
AND2X1   g1904(.A(WX4376), .B(RESET), .Y(n3520));
AND2X1   g1905(.A(WX4378), .B(RESET), .Y(n3525));
AND2X1   g1906(.A(WX4380), .B(RESET), .Y(n3530));
AND2X1   g1907(.A(WX4382), .B(RESET), .Y(n3535));
AND2X1   g1908(.A(WX4384), .B(RESET), .Y(n3540));
AND2X1   g1909(.A(WX4386), .B(RESET), .Y(n3545));
AND2X1   g1910(.A(WX4388), .B(RESET), .Y(n3550));
AND2X1   g1911(.A(WX4390), .B(RESET), .Y(n3555));
AND2X1   g1912(.A(WX4392), .B(RESET), .Y(n3560));
AND2X1   g1913(.A(WX4394), .B(RESET), .Y(n3565));
AND2X1   g1914(.A(WX4396), .B(RESET), .Y(n3570));
AND2X1   g1915(.A(WX4398), .B(RESET), .Y(n3575));
AND2X1   g1916(.A(WX4400), .B(RESET), .Y(n3580));
AND2X1   g1917(.A(WX4402), .B(RESET), .Y(n3585));
AND2X1   g1918(.A(WX4404), .B(RESET), .Y(n3590));
AND2X1   g1919(.A(WX4406), .B(RESET), .Y(n3595));
AND2X1   g1920(.A(WX4408), .B(RESET), .Y(n3600));
AND2X1   g1921(.A(WX4410), .B(RESET), .Y(n3605));
AND2X1   g1922(.A(WX4412), .B(RESET), .Y(n3610));
AND2X1   g1923(.A(WX4414), .B(RESET), .Y(n3615));
AND2X1   g1924(.A(WX4416), .B(RESET), .Y(n3620));
AND2X1   g1925(.A(WX4418), .B(RESET), .Y(n3625));
AND2X1   g1926(.A(WX4420), .B(RESET), .Y(n3630));
AND2X1   g1927(.A(WX4422), .B(RESET), .Y(n3635));
AND2X1   g1928(.A(WX4424), .B(RESET), .Y(n3640));
AND2X1   g1929(.A(WX4426), .B(RESET), .Y(n3645));
NOR2X1   g1930(.A(WX4364), .B(n5827), .Y(n3650));
INVX1    g1931(.A(CRC_OUT_6_31), .Y(n7566));
XOR2X1   g1932(.A(WX5817), .B(TM1), .Y(n7567_1));
XOR2X1   g1933(.A(n7567_1), .B(WX5881), .Y(n7568));
INVX1    g1934(.A(WX5945), .Y(n7569));
XOR2X1   g1935(.A(WX6009), .B(n7569), .Y(n7570));
XOR2X1   g1936(.A(n7570), .B(n7568), .Y(n7571));
MX2X1    g1937(.A(n7566), .B(n7571), .S0(n5539), .Y(n7573));
INVX1    g1938(.A(WX4364), .Y(n7574));
MX2X1    g1939(.A(n7574), .B(n6992), .S0(n5539), .Y(n7575));
MX2X1    g1940(.A(n7573), .B(n7575), .S0(TM1), .Y(n7576));
NOR2X1   g1941(.A(n7576), .B(n5827), .Y(n3655));
INVX1    g1942(.A(CRC_OUT_6_30), .Y(n7578));
XOR2X1   g1943(.A(WX5819), .B(TM1), .Y(n7579));
XOR2X1   g1944(.A(n7579), .B(WX5883), .Y(n7580));
INVX1    g1945(.A(WX5947), .Y(n7581));
XOR2X1   g1946(.A(WX6011), .B(n7581), .Y(n7582_1));
XOR2X1   g1947(.A(n7582_1), .B(n7580), .Y(n7583));
MX2X1    g1948(.A(n7578), .B(n7583), .S0(n5539), .Y(n7585));
INVX1    g1949(.A(WX4366), .Y(n7586));
MX2X1    g1950(.A(n7586), .B(n7004_1), .S0(n5539), .Y(n7587_1));
MX2X1    g1951(.A(n7585), .B(n7587_1), .S0(TM1), .Y(n7588));
NOR2X1   g1952(.A(n7588), .B(n5827), .Y(n3660));
INVX1    g1953(.A(CRC_OUT_6_29), .Y(n7590));
XOR2X1   g1954(.A(WX5821), .B(TM1), .Y(n7591));
XOR2X1   g1955(.A(n7591), .B(WX5885), .Y(n7592_1));
INVX1    g1956(.A(WX5949), .Y(n7593));
XOR2X1   g1957(.A(WX6013), .B(n7593), .Y(n7594));
XOR2X1   g1958(.A(n7594), .B(n7592_1), .Y(n7595));
MX2X1    g1959(.A(n7590), .B(n7595), .S0(n5539), .Y(n7597_1));
INVX1    g1960(.A(WX4368), .Y(n7598));
MX2X1    g1961(.A(n7598), .B(n7016), .S0(n5539), .Y(n7599));
MX2X1    g1962(.A(n7597_1), .B(n7599), .S0(TM1), .Y(n7600));
NOR2X1   g1963(.A(n7600), .B(n5827), .Y(n3665));
INVX1    g1964(.A(CRC_OUT_6_28), .Y(n7602_1));
XOR2X1   g1965(.A(WX5823), .B(TM1), .Y(n7603));
XOR2X1   g1966(.A(n7603), .B(WX5887), .Y(n7604));
INVX1    g1967(.A(WX5951), .Y(n7605));
XOR2X1   g1968(.A(WX6015), .B(n7605), .Y(n7606));
XOR2X1   g1969(.A(n7606), .B(n7604), .Y(n7607_1));
MX2X1    g1970(.A(n7602_1), .B(n7607_1), .S0(n5539), .Y(n7609));
INVX1    g1971(.A(WX4370), .Y(n7610));
MX2X1    g1972(.A(n7610), .B(n7028), .S0(n5539), .Y(n7611));
MX2X1    g1973(.A(n7609), .B(n7611), .S0(TM1), .Y(n7612_1));
NOR2X1   g1974(.A(n7612_1), .B(n5827), .Y(n3670));
INVX1    g1975(.A(CRC_OUT_6_27), .Y(n7614));
XOR2X1   g1976(.A(WX5825), .B(TM1), .Y(n7615));
XOR2X1   g1977(.A(n7615), .B(WX5889), .Y(n7616));
INVX1    g1978(.A(WX5953), .Y(n7617_1));
XOR2X1   g1979(.A(WX6017), .B(n7617_1), .Y(n7618));
XOR2X1   g1980(.A(n7618), .B(n7616), .Y(n7619));
MX2X1    g1981(.A(n7614), .B(n7619), .S0(n5539), .Y(n7621));
INVX1    g1982(.A(WX4372), .Y(n7622_1));
MX2X1    g1983(.A(n7622_1), .B(n7040), .S0(n5539), .Y(n7623));
MX2X1    g1984(.A(n7621), .B(n7623), .S0(TM1), .Y(n7624));
NOR2X1   g1985(.A(n7624), .B(n5827), .Y(n3675));
INVX1    g1986(.A(CRC_OUT_6_26), .Y(n7626));
XOR2X1   g1987(.A(WX5827), .B(TM1), .Y(n7627_1));
XOR2X1   g1988(.A(n7627_1), .B(WX5891), .Y(n7628));
INVX1    g1989(.A(WX5955), .Y(n7629));
XOR2X1   g1990(.A(WX6019), .B(n7629), .Y(n7630));
XOR2X1   g1991(.A(n7630), .B(n7628), .Y(n7631));
MX2X1    g1992(.A(n7626), .B(n7631), .S0(n5539), .Y(n7633));
INVX1    g1993(.A(WX4374), .Y(n7634));
MX2X1    g1994(.A(n7634), .B(n7052), .S0(n5539), .Y(n7635));
MX2X1    g1995(.A(n7633), .B(n7635), .S0(TM1), .Y(n7636));
NOR2X1   g1996(.A(n7636), .B(n5827), .Y(n3680));
INVX1    g1997(.A(CRC_OUT_6_25), .Y(n7638));
XOR2X1   g1998(.A(WX5829), .B(TM1), .Y(n7639));
XOR2X1   g1999(.A(n7639), .B(WX5893), .Y(n7640));
INVX1    g2000(.A(WX5957), .Y(n7641));
XOR2X1   g2001(.A(WX6021), .B(n7641), .Y(n7642_1));
XOR2X1   g2002(.A(n7642_1), .B(n7640), .Y(n7643));
MX2X1    g2003(.A(n7638), .B(n7643), .S0(n5539), .Y(n7645));
INVX1    g2004(.A(WX4376), .Y(n7646));
MX2X1    g2005(.A(n7646), .B(n7064_1), .S0(n5539), .Y(n7647_1));
MX2X1    g2006(.A(n7645), .B(n7647_1), .S0(TM1), .Y(n7648));
NOR2X1   g2007(.A(n7648), .B(n5827), .Y(n3685));
INVX1    g2008(.A(CRC_OUT_6_24), .Y(n7650));
XOR2X1   g2009(.A(WX5831), .B(TM1), .Y(n7651));
XOR2X1   g2010(.A(n7651), .B(WX5895), .Y(n7652_1));
INVX1    g2011(.A(WX5959), .Y(n7653));
XOR2X1   g2012(.A(WX6023), .B(n7653), .Y(n7654));
XOR2X1   g2013(.A(n7654), .B(n7652_1), .Y(n7655));
MX2X1    g2014(.A(n7650), .B(n7655), .S0(n5539), .Y(n7657_1));
INVX1    g2015(.A(WX4378), .Y(n7658));
MX2X1    g2016(.A(n7658), .B(n7076), .S0(n5539), .Y(n7659));
MX2X1    g2017(.A(n7657_1), .B(n7659), .S0(TM1), .Y(n7660));
NOR2X1   g2018(.A(n7660), .B(n5827), .Y(n3690));
INVX1    g2019(.A(CRC_OUT_6_23), .Y(n7662_1));
XOR2X1   g2020(.A(WX5833), .B(TM1), .Y(n7663));
XOR2X1   g2021(.A(n7663), .B(WX5897), .Y(n7664));
INVX1    g2022(.A(WX5961), .Y(n7665));
XOR2X1   g2023(.A(WX6025), .B(n7665), .Y(n7666));
XOR2X1   g2024(.A(n7666), .B(n7664), .Y(n7667_1));
MX2X1    g2025(.A(n7662_1), .B(n7667_1), .S0(n5539), .Y(n7669));
INVX1    g2026(.A(WX4380), .Y(n7670));
MX2X1    g2027(.A(n7670), .B(n7088), .S0(n5539), .Y(n7671));
MX2X1    g2028(.A(n7669), .B(n7671), .S0(TM1), .Y(n7672_1));
NOR2X1   g2029(.A(n7672_1), .B(n5827), .Y(n3695));
INVX1    g2030(.A(CRC_OUT_6_22), .Y(n7674));
XOR2X1   g2031(.A(WX5835), .B(TM1), .Y(n7675));
XOR2X1   g2032(.A(n7675), .B(WX5899), .Y(n7676));
INVX1    g2033(.A(WX5963), .Y(n7677_1));
XOR2X1   g2034(.A(WX6027), .B(n7677_1), .Y(n7678));
XOR2X1   g2035(.A(n7678), .B(n7676), .Y(n7679));
MX2X1    g2036(.A(n7674), .B(n7679), .S0(n5539), .Y(n7681));
INVX1    g2037(.A(WX4382), .Y(n7682_1));
MX2X1    g2038(.A(n7682_1), .B(n7100), .S0(n5539), .Y(n7683));
MX2X1    g2039(.A(n7681), .B(n7683), .S0(TM1), .Y(n7684));
NOR2X1   g2040(.A(n7684), .B(n5827), .Y(n3700));
INVX1    g2041(.A(CRC_OUT_6_21), .Y(n7686));
XOR2X1   g2042(.A(WX5837), .B(TM1), .Y(n7687_1));
XOR2X1   g2043(.A(n7687_1), .B(WX5901), .Y(n7688));
INVX1    g2044(.A(WX5965), .Y(n7689));
XOR2X1   g2045(.A(WX6029), .B(n7689), .Y(n7690));
XOR2X1   g2046(.A(n7690), .B(n7688), .Y(n7691));
MX2X1    g2047(.A(n7686), .B(n7691), .S0(n5539), .Y(n7693));
INVX1    g2048(.A(WX4384), .Y(n7694));
MX2X1    g2049(.A(n7694), .B(n7112), .S0(n5539), .Y(n7695));
MX2X1    g2050(.A(n7693), .B(n7695), .S0(TM1), .Y(n7696));
NOR2X1   g2051(.A(n7696), .B(n5827), .Y(n3705));
INVX1    g2052(.A(CRC_OUT_6_20), .Y(n7698));
XOR2X1   g2053(.A(WX5839), .B(TM1), .Y(n7699));
XOR2X1   g2054(.A(n7699), .B(WX5903), .Y(n7700));
INVX1    g2055(.A(WX5967), .Y(n7701));
XOR2X1   g2056(.A(WX6031), .B(n7701), .Y(n7702_1));
XOR2X1   g2057(.A(n7702_1), .B(n7700), .Y(n7703));
MX2X1    g2058(.A(n7698), .B(n7703), .S0(n5539), .Y(n7705));
INVX1    g2059(.A(WX4386), .Y(n7706));
MX2X1    g2060(.A(n7706), .B(n7124), .S0(n5539), .Y(n7707_1));
MX2X1    g2061(.A(n7705), .B(n7707_1), .S0(TM1), .Y(n7708));
NOR2X1   g2062(.A(n7708), .B(n5827), .Y(n3710));
INVX1    g2063(.A(CRC_OUT_6_19), .Y(n7710));
XOR2X1   g2064(.A(WX5841), .B(TM1), .Y(n7711));
XOR2X1   g2065(.A(n7711), .B(WX5905), .Y(n7712_1));
INVX1    g2066(.A(WX5969), .Y(n7713));
XOR2X1   g2067(.A(WX6033), .B(n7713), .Y(n7714));
XOR2X1   g2068(.A(n7714), .B(n7712_1), .Y(n7715));
MX2X1    g2069(.A(n7710), .B(n7715), .S0(n5539), .Y(n7717_1));
INVX1    g2070(.A(WX4388), .Y(n7718));
MX2X1    g2071(.A(n7718), .B(n7136), .S0(n5539), .Y(n7719));
MX2X1    g2072(.A(n7717_1), .B(n7719), .S0(TM1), .Y(n7720));
NOR2X1   g2073(.A(n7720), .B(n5827), .Y(n3715));
INVX1    g2074(.A(CRC_OUT_6_18), .Y(n7722_1));
XOR2X1   g2075(.A(WX5843), .B(TM1), .Y(n7723));
XOR2X1   g2076(.A(n7723), .B(WX5907), .Y(n7724));
INVX1    g2077(.A(WX5971), .Y(n7725));
XOR2X1   g2078(.A(WX6035), .B(n7725), .Y(n7726));
XOR2X1   g2079(.A(n7726), .B(n7724), .Y(n7727_1));
MX2X1    g2080(.A(n7722_1), .B(n7727_1), .S0(n5539), .Y(n7729));
INVX1    g2081(.A(WX4390), .Y(n7730));
MX2X1    g2082(.A(n7730), .B(n7148), .S0(n5539), .Y(n7731));
MX2X1    g2083(.A(n7729), .B(n7731), .S0(TM1), .Y(n7732_1));
NOR2X1   g2084(.A(n7732_1), .B(n5827), .Y(n3720));
INVX1    g2085(.A(CRC_OUT_6_17), .Y(n7734));
XOR2X1   g2086(.A(WX5845), .B(TM1), .Y(n7735));
XOR2X1   g2087(.A(n7735), .B(WX5909), .Y(n7736));
INVX1    g2088(.A(WX5973), .Y(n7737_1));
XOR2X1   g2089(.A(WX6037), .B(n7737_1), .Y(n7738));
XOR2X1   g2090(.A(n7738), .B(n7736), .Y(n7739));
MX2X1    g2091(.A(n7734), .B(n7739), .S0(n5539), .Y(n7741));
INVX1    g2092(.A(WX4392), .Y(n7742_1));
MX2X1    g2093(.A(n7742_1), .B(n7160), .S0(n5539), .Y(n7743));
MX2X1    g2094(.A(n7741), .B(n7743), .S0(TM1), .Y(n7744));
NOR2X1   g2095(.A(n7744), .B(n5827), .Y(n3725));
INVX1    g2096(.A(CRC_OUT_6_16), .Y(n7746));
XOR2X1   g2097(.A(WX5847), .B(TM1), .Y(n7747_1));
XOR2X1   g2098(.A(n7747_1), .B(WX5911), .Y(n7748));
INVX1    g2099(.A(WX5975), .Y(n7749));
XOR2X1   g2100(.A(WX6039), .B(n7749), .Y(n7750));
XOR2X1   g2101(.A(n7750), .B(n7748), .Y(n7751));
MX2X1    g2102(.A(n7746), .B(n7751), .S0(n5539), .Y(n7753));
INVX1    g2103(.A(WX4394), .Y(n7754));
MX2X1    g2104(.A(n7754), .B(n7172), .S0(n5539), .Y(n7755));
MX2X1    g2105(.A(n7753), .B(n7755), .S0(TM1), .Y(n7756));
NOR2X1   g2106(.A(n7756), .B(n5827), .Y(n3730));
INVX1    g2107(.A(CRC_OUT_6_15), .Y(n7758));
XOR2X1   g2108(.A(WX5849), .B(TM0), .Y(n7759));
XOR2X1   g2109(.A(n7759), .B(WX5913), .Y(n7760));
INVX1    g2110(.A(WX5977), .Y(n7761));
XOR2X1   g2111(.A(WX6041), .B(n7761), .Y(n7762_1));
XOR2X1   g2112(.A(n7762_1), .B(n7760), .Y(n7763));
MX2X1    g2113(.A(n7758), .B(n7763), .S0(n5539), .Y(n7765));
INVX1    g2114(.A(WX4396), .Y(n7766));
MX2X1    g2115(.A(n7766), .B(n7184), .S0(n5539), .Y(n7767_1));
MX2X1    g2116(.A(n7765), .B(n7767_1), .S0(TM1), .Y(n7768));
NOR2X1   g2117(.A(n7768), .B(n5827), .Y(n3735));
INVX1    g2118(.A(CRC_OUT_6_14), .Y(n7770));
XOR2X1   g2119(.A(WX5851), .B(TM0), .Y(n7771));
XOR2X1   g2120(.A(n7771), .B(WX5915), .Y(n7772_1));
INVX1    g2121(.A(WX5979), .Y(n7773));
XOR2X1   g2122(.A(WX6043), .B(n7773), .Y(n7774));
XOR2X1   g2123(.A(n7774), .B(n7772_1), .Y(n7775));
MX2X1    g2124(.A(n7770), .B(n7775), .S0(n5539), .Y(n7777_1));
INVX1    g2125(.A(WX4398), .Y(n7778));
MX2X1    g2126(.A(n7778), .B(n7196), .S0(n5539), .Y(n7779));
MX2X1    g2127(.A(n7777_1), .B(n7779), .S0(TM1), .Y(n7780));
NOR2X1   g2128(.A(n7780), .B(n5827), .Y(n3740));
INVX1    g2129(.A(CRC_OUT_6_13), .Y(n7782_1));
XOR2X1   g2130(.A(WX5853), .B(TM0), .Y(n7783));
XOR2X1   g2131(.A(n7783), .B(WX5917), .Y(n7784));
INVX1    g2132(.A(WX5981), .Y(n7785));
XOR2X1   g2133(.A(WX6045), .B(n7785), .Y(n7786));
XOR2X1   g2134(.A(n7786), .B(n7784), .Y(n7787_1));
MX2X1    g2135(.A(n7782_1), .B(n7787_1), .S0(n5539), .Y(n7789));
INVX1    g2136(.A(WX4400), .Y(n7790));
MX2X1    g2137(.A(n7790), .B(n7208), .S0(n5539), .Y(n7791));
MX2X1    g2138(.A(n7789), .B(n7791), .S0(TM1), .Y(n7792_1));
NOR2X1   g2139(.A(n7792_1), .B(n5827), .Y(n3745));
INVX1    g2140(.A(CRC_OUT_6_12), .Y(n7794));
XOR2X1   g2141(.A(WX5855), .B(TM0), .Y(n7795));
XOR2X1   g2142(.A(n7795), .B(WX5919), .Y(n7796));
INVX1    g2143(.A(WX5983), .Y(n7797_1));
XOR2X1   g2144(.A(WX6047), .B(n7797_1), .Y(n7798));
XOR2X1   g2145(.A(n7798), .B(n7796), .Y(n7799));
MX2X1    g2146(.A(n7794), .B(n7799), .S0(n5539), .Y(n7801));
INVX1    g2147(.A(WX4402), .Y(n7802_1));
MX2X1    g2148(.A(n7802_1), .B(n7220), .S0(n5539), .Y(n7803));
MX2X1    g2149(.A(n7801), .B(n7803), .S0(TM1), .Y(n7804));
NOR2X1   g2150(.A(n7804), .B(n5827), .Y(n3750));
INVX1    g2151(.A(CRC_OUT_6_11), .Y(n7806));
XOR2X1   g2152(.A(WX5857), .B(TM0), .Y(n7807_1));
XOR2X1   g2153(.A(n7807_1), .B(WX5921), .Y(n7808));
INVX1    g2154(.A(WX5985), .Y(n7809));
XOR2X1   g2155(.A(WX6049), .B(n7809), .Y(n7810));
XOR2X1   g2156(.A(n7810), .B(n7808), .Y(n7811));
MX2X1    g2157(.A(n7806), .B(n7811), .S0(n5539), .Y(n7813));
INVX1    g2158(.A(WX4404), .Y(n7814));
MX2X1    g2159(.A(n7814), .B(n7232_1), .S0(n5539), .Y(n7815));
MX2X1    g2160(.A(n7813), .B(n7815), .S0(TM1), .Y(n7816));
NOR2X1   g2161(.A(n7816), .B(n5827), .Y(n3755));
INVX1    g2162(.A(CRC_OUT_6_10), .Y(n7818));
XOR2X1   g2163(.A(WX5859), .B(TM0), .Y(n7819));
XOR2X1   g2164(.A(n7819), .B(WX5923), .Y(n7820));
INVX1    g2165(.A(WX5987), .Y(n7821));
XOR2X1   g2166(.A(WX6051), .B(n7821), .Y(n7822_1));
XOR2X1   g2167(.A(n7822_1), .B(n7820), .Y(n7823));
MX2X1    g2168(.A(n7818), .B(n7823), .S0(n5539), .Y(n7825));
INVX1    g2169(.A(WX4406), .Y(n7826));
MX2X1    g2170(.A(n7826), .B(n7244), .S0(n5539), .Y(n7827_1));
MX2X1    g2171(.A(n7825), .B(n7827_1), .S0(TM1), .Y(n7828));
NOR2X1   g2172(.A(n7828), .B(n5827), .Y(n3760));
INVX1    g2173(.A(CRC_OUT_6_9), .Y(n7830));
XOR2X1   g2174(.A(WX5861), .B(TM0), .Y(n7831));
XOR2X1   g2175(.A(n7831), .B(WX5925), .Y(n7832_1));
INVX1    g2176(.A(WX5989), .Y(n7833));
XOR2X1   g2177(.A(WX6053), .B(n7833), .Y(n7834));
XOR2X1   g2178(.A(n7834), .B(n7832_1), .Y(n7835));
MX2X1    g2179(.A(n7830), .B(n7835), .S0(n5539), .Y(n7837_1));
INVX1    g2180(.A(WX4408), .Y(n7838));
MX2X1    g2181(.A(n7838), .B(n7256), .S0(n5539), .Y(n7839));
MX2X1    g2182(.A(n7837_1), .B(n7839), .S0(TM1), .Y(n7840));
NOR2X1   g2183(.A(n7840), .B(n5827), .Y(n3765));
INVX1    g2184(.A(CRC_OUT_6_8), .Y(n7842_1));
XOR2X1   g2185(.A(WX5863), .B(TM0), .Y(n7843));
XOR2X1   g2186(.A(n7843), .B(WX5927), .Y(n7844));
INVX1    g2187(.A(WX5991), .Y(n7845));
XOR2X1   g2188(.A(WX6055), .B(n7845), .Y(n7846));
XOR2X1   g2189(.A(n7846), .B(n7844), .Y(n7847_1));
MX2X1    g2190(.A(n7842_1), .B(n7847_1), .S0(n5539), .Y(n7849));
INVX1    g2191(.A(WX4410), .Y(n7850));
MX2X1    g2192(.A(n7850), .B(n7268), .S0(n5539), .Y(n7851));
MX2X1    g2193(.A(n7849), .B(n7851), .S0(TM1), .Y(n7852_1));
NOR2X1   g2194(.A(n7852_1), .B(n5827), .Y(n3770));
INVX1    g2195(.A(CRC_OUT_6_7), .Y(n7854));
XOR2X1   g2196(.A(WX5865), .B(TM0), .Y(n7855));
XOR2X1   g2197(.A(n7855), .B(WX5929), .Y(n7856));
INVX1    g2198(.A(WX5993), .Y(n7857_1));
XOR2X1   g2199(.A(WX6057), .B(n7857_1), .Y(n7858));
XOR2X1   g2200(.A(n7858), .B(n7856), .Y(n7859));
MX2X1    g2201(.A(n7854), .B(n7859), .S0(n5539), .Y(n7861));
INVX1    g2202(.A(WX4412), .Y(n7862_1));
MX2X1    g2203(.A(n7862_1), .B(n7280), .S0(n5539), .Y(n7863));
MX2X1    g2204(.A(n7861), .B(n7863), .S0(TM1), .Y(n7864));
NOR2X1   g2205(.A(n7864), .B(n5827), .Y(n3775));
INVX1    g2206(.A(CRC_OUT_6_6), .Y(n7866));
XOR2X1   g2207(.A(WX5867), .B(TM0), .Y(n7867_1));
XOR2X1   g2208(.A(n7867_1), .B(WX5931), .Y(n7868));
INVX1    g2209(.A(WX5995), .Y(n7869));
XOR2X1   g2210(.A(WX6059), .B(n7869), .Y(n7870));
XOR2X1   g2211(.A(n7870), .B(n7868), .Y(n7871));
MX2X1    g2212(.A(n7866), .B(n7871), .S0(n5539), .Y(n7873));
INVX1    g2213(.A(WX4414), .Y(n7874));
MX2X1    g2214(.A(n7874), .B(n7292_1), .S0(n5539), .Y(n7875));
MX2X1    g2215(.A(n7873), .B(n7875), .S0(TM1), .Y(n7876));
NOR2X1   g2216(.A(n7876), .B(n5827), .Y(n3780));
INVX1    g2217(.A(CRC_OUT_6_5), .Y(n7878));
XOR2X1   g2218(.A(WX5869), .B(TM0), .Y(n7879));
XOR2X1   g2219(.A(n7879), .B(WX5933), .Y(n7880));
INVX1    g2220(.A(WX5997), .Y(n7881));
XOR2X1   g2221(.A(WX6061), .B(n7881), .Y(n7882_1));
XOR2X1   g2222(.A(n7882_1), .B(n7880), .Y(n7883));
MX2X1    g2223(.A(n7878), .B(n7883), .S0(n5539), .Y(n7885));
INVX1    g2224(.A(WX4416), .Y(n7886));
MX2X1    g2225(.A(n7886), .B(n7304), .S0(n5539), .Y(n7887_1));
MX2X1    g2226(.A(n7885), .B(n7887_1), .S0(TM1), .Y(n7888));
NOR2X1   g2227(.A(n7888), .B(n5827), .Y(n3785));
INVX1    g2228(.A(CRC_OUT_6_4), .Y(n7890));
XOR2X1   g2229(.A(WX5871), .B(TM0), .Y(n7891));
XOR2X1   g2230(.A(n7891), .B(WX5935), .Y(n7892_1));
INVX1    g2231(.A(WX5999), .Y(n7893));
XOR2X1   g2232(.A(WX6063), .B(n7893), .Y(n7894));
XOR2X1   g2233(.A(n7894), .B(n7892_1), .Y(n7895));
MX2X1    g2234(.A(n7890), .B(n7895), .S0(n5539), .Y(n7897_1));
INVX1    g2235(.A(WX4418), .Y(n7898));
MX2X1    g2236(.A(n7898), .B(n7316), .S0(n5539), .Y(n7899));
MX2X1    g2237(.A(n7897_1), .B(n7899), .S0(TM1), .Y(n7900));
NOR2X1   g2238(.A(n7900), .B(n5827), .Y(n3790));
INVX1    g2239(.A(CRC_OUT_6_3), .Y(n7902_1));
XOR2X1   g2240(.A(WX5873), .B(TM0), .Y(n7903));
XOR2X1   g2241(.A(n7903), .B(WX5937), .Y(n7904));
INVX1    g2242(.A(WX6001), .Y(n7905));
XOR2X1   g2243(.A(WX6065), .B(n7905), .Y(n7906));
XOR2X1   g2244(.A(n7906), .B(n7904), .Y(n7907_1));
MX2X1    g2245(.A(n7902_1), .B(n7907_1), .S0(n5539), .Y(n7909));
INVX1    g2246(.A(WX4420), .Y(n7910));
MX2X1    g2247(.A(n7910), .B(n7328), .S0(n5539), .Y(n7911));
MX2X1    g2248(.A(n7909), .B(n7911), .S0(TM1), .Y(n7912_1));
NOR2X1   g2249(.A(n7912_1), .B(n5827), .Y(n3795));
INVX1    g2250(.A(CRC_OUT_6_2), .Y(n7914));
XOR2X1   g2251(.A(WX5875), .B(TM0), .Y(n7915));
XOR2X1   g2252(.A(n7915), .B(WX5939), .Y(n7916));
INVX1    g2253(.A(WX6003), .Y(n7917_1));
XOR2X1   g2254(.A(WX6067), .B(n7917_1), .Y(n7918));
XOR2X1   g2255(.A(n7918), .B(n7916), .Y(n7919));
MX2X1    g2256(.A(n7914), .B(n7919), .S0(n5539), .Y(n7921));
INVX1    g2257(.A(WX4422), .Y(n7922_1));
MX2X1    g2258(.A(n7922_1), .B(n7340), .S0(n5539), .Y(n7923));
MX2X1    g2259(.A(n7921), .B(n7923), .S0(TM1), .Y(n7924));
NOR2X1   g2260(.A(n7924), .B(n5827), .Y(n3800));
INVX1    g2261(.A(CRC_OUT_6_1), .Y(n7926));
XOR2X1   g2262(.A(WX5877), .B(TM0), .Y(n7927_1));
XOR2X1   g2263(.A(n7927_1), .B(WX5941), .Y(n7928));
INVX1    g2264(.A(WX6005), .Y(n7929));
XOR2X1   g2265(.A(WX6069), .B(n7929), .Y(n7930));
XOR2X1   g2266(.A(n7930), .B(n7928), .Y(n7931));
MX2X1    g2267(.A(n7926), .B(n7931), .S0(n5539), .Y(n7933));
INVX1    g2268(.A(WX4424), .Y(n7934));
MX2X1    g2269(.A(n7934), .B(n7352_1), .S0(n5539), .Y(n7935));
MX2X1    g2270(.A(n7933), .B(n7935), .S0(TM1), .Y(n7936));
NOR2X1   g2271(.A(n7936), .B(n5827), .Y(n3805));
INVX1    g2272(.A(CRC_OUT_6_0), .Y(n7938));
XOR2X1   g2273(.A(WX5879), .B(TM0), .Y(n7939));
XOR2X1   g2274(.A(n7939), .B(WX5943), .Y(n7940));
INVX1    g2275(.A(WX6007), .Y(n7941));
XOR2X1   g2276(.A(WX6071), .B(n7941), .Y(n7942_1));
XOR2X1   g2277(.A(n7942_1), .B(n7940), .Y(n7943));
MX2X1    g2278(.A(n7938), .B(n7943), .S0(n5539), .Y(n7945));
INVX1    g2279(.A(WX4426), .Y(n7946));
MX2X1    g2280(.A(n7946), .B(n7364), .S0(n5539), .Y(n7947_1));
MX2X1    g2281(.A(n7945), .B(n7947_1), .S0(TM1), .Y(n7948));
NOR2X1   g2282(.A(n7948), .B(n5827), .Y(n3810));
AND2X1   g2283(.A(WX4524), .B(RESET), .Y(n3815));
AND2X1   g2284(.A(WX4526), .B(RESET), .Y(n3820));
AND2X1   g2285(.A(WX4528), .B(RESET), .Y(n3825));
AND2X1   g2286(.A(WX4530), .B(RESET), .Y(n3830));
AND2X1   g2287(.A(WX4532), .B(RESET), .Y(n3835));
AND2X1   g2288(.A(WX4534), .B(RESET), .Y(n3840));
AND2X1   g2289(.A(WX4536), .B(RESET), .Y(n3845));
AND2X1   g2290(.A(WX4538), .B(RESET), .Y(n3850));
AND2X1   g2291(.A(WX4540), .B(RESET), .Y(n3855));
AND2X1   g2292(.A(WX4542), .B(RESET), .Y(n3860));
AND2X1   g2293(.A(WX4544), .B(RESET), .Y(n3865));
AND2X1   g2294(.A(WX4546), .B(RESET), .Y(n3870));
AND2X1   g2295(.A(WX4548), .B(RESET), .Y(n3875));
AND2X1   g2296(.A(WX4550), .B(RESET), .Y(n3880));
AND2X1   g2297(.A(WX4552), .B(RESET), .Y(n3885));
AND2X1   g2298(.A(WX4554), .B(RESET), .Y(n3890));
AND2X1   g2299(.A(WX4556), .B(RESET), .Y(n3895));
AND2X1   g2300(.A(WX4558), .B(RESET), .Y(n3900));
AND2X1   g2301(.A(WX4560), .B(RESET), .Y(n3905));
AND2X1   g2302(.A(WX4562), .B(RESET), .Y(n3910));
AND2X1   g2303(.A(WX4564), .B(RESET), .Y(n3915));
AND2X1   g2304(.A(WX4566), .B(RESET), .Y(n3920));
AND2X1   g2305(.A(WX4568), .B(RESET), .Y(n3925));
AND2X1   g2306(.A(WX4570), .B(RESET), .Y(n3930));
AND2X1   g2307(.A(WX4572), .B(RESET), .Y(n3935));
AND2X1   g2308(.A(WX4574), .B(RESET), .Y(n3940));
AND2X1   g2309(.A(WX4576), .B(RESET), .Y(n3945));
AND2X1   g2310(.A(WX4578), .B(RESET), .Y(n3950));
AND2X1   g2311(.A(WX4580), .B(RESET), .Y(n3955));
AND2X1   g2312(.A(WX4582), .B(RESET), .Y(n3960));
AND2X1   g2313(.A(WX4584), .B(RESET), .Y(n3965));
AND2X1   g2314(.A(WX4586), .B(RESET), .Y(n3970));
AND2X1   g2315(.A(WX4588), .B(RESET), .Y(n3975));
AND2X1   g2316(.A(WX4590), .B(RESET), .Y(n3980));
AND2X1   g2317(.A(WX4592), .B(RESET), .Y(n3985));
AND2X1   g2318(.A(WX4594), .B(RESET), .Y(n3990));
AND2X1   g2319(.A(WX4596), .B(RESET), .Y(n3995));
AND2X1   g2320(.A(WX4598), .B(RESET), .Y(n4000));
AND2X1   g2321(.A(WX4600), .B(RESET), .Y(n4005));
AND2X1   g2322(.A(WX4602), .B(RESET), .Y(n4010));
AND2X1   g2323(.A(WX4604), .B(RESET), .Y(n4015));
AND2X1   g2324(.A(WX4606), .B(RESET), .Y(n4020));
AND2X1   g2325(.A(WX4608), .B(RESET), .Y(n4025));
AND2X1   g2326(.A(WX4610), .B(RESET), .Y(n4030));
AND2X1   g2327(.A(WX4612), .B(RESET), .Y(n4035));
AND2X1   g2328(.A(WX4614), .B(RESET), .Y(n4040));
AND2X1   g2329(.A(WX4616), .B(RESET), .Y(n4045));
AND2X1   g2330(.A(WX4618), .B(RESET), .Y(n4050));
AND2X1   g2331(.A(WX4620), .B(RESET), .Y(n4055));
AND2X1   g2332(.A(WX4622), .B(RESET), .Y(n4060));
AND2X1   g2333(.A(WX4624), .B(RESET), .Y(n4065));
AND2X1   g2334(.A(WX4626), .B(RESET), .Y(n4070));
AND2X1   g2335(.A(WX4628), .B(RESET), .Y(n4075));
AND2X1   g2336(.A(WX4630), .B(RESET), .Y(n4080));
AND2X1   g2337(.A(WX4632), .B(RESET), .Y(n4085));
AND2X1   g2338(.A(WX4634), .B(RESET), .Y(n4090));
AND2X1   g2339(.A(WX4636), .B(RESET), .Y(n4095));
AND2X1   g2340(.A(WX4638), .B(RESET), .Y(n4100));
AND2X1   g2341(.A(WX4640), .B(RESET), .Y(n4105));
AND2X1   g2342(.A(WX4642), .B(RESET), .Y(n4110));
AND2X1   g2343(.A(WX4644), .B(RESET), .Y(n4115));
AND2X1   g2344(.A(WX4646), .B(RESET), .Y(n4120));
AND2X1   g2345(.A(WX4648), .B(RESET), .Y(n4125));
AND2X1   g2346(.A(WX4650), .B(RESET), .Y(n4130));
AND2X1   g2347(.A(WX4652), .B(RESET), .Y(n4135));
AND2X1   g2348(.A(WX4654), .B(RESET), .Y(n4140));
AND2X1   g2349(.A(WX4656), .B(RESET), .Y(n4145));
AND2X1   g2350(.A(WX4658), .B(RESET), .Y(n4150));
AND2X1   g2351(.A(WX4660), .B(RESET), .Y(n4155));
AND2X1   g2352(.A(WX4662), .B(RESET), .Y(n4160));
AND2X1   g2353(.A(WX4664), .B(RESET), .Y(n4165));
AND2X1   g2354(.A(WX4666), .B(RESET), .Y(n4170));
AND2X1   g2355(.A(WX4668), .B(RESET), .Y(n4175));
AND2X1   g2356(.A(WX4670), .B(RESET), .Y(n4180));
AND2X1   g2357(.A(WX4672), .B(RESET), .Y(n4185));
AND2X1   g2358(.A(WX4674), .B(RESET), .Y(n4190));
AND2X1   g2359(.A(WX4676), .B(RESET), .Y(n4195));
AND2X1   g2360(.A(WX4678), .B(RESET), .Y(n4200));
AND2X1   g2361(.A(WX4680), .B(RESET), .Y(n4205));
AND2X1   g2362(.A(WX4682), .B(RESET), .Y(n4210));
AND2X1   g2363(.A(WX4684), .B(RESET), .Y(n4215));
AND2X1   g2364(.A(WX4686), .B(RESET), .Y(n4220));
AND2X1   g2365(.A(WX4688), .B(RESET), .Y(n4225));
AND2X1   g2366(.A(WX4690), .B(RESET), .Y(n4230));
AND2X1   g2367(.A(WX4692), .B(RESET), .Y(n4235));
AND2X1   g2368(.A(WX4694), .B(RESET), .Y(n4240));
AND2X1   g2369(.A(WX4696), .B(RESET), .Y(n4245));
AND2X1   g2370(.A(WX4698), .B(RESET), .Y(n4250));
AND2X1   g2371(.A(WX4700), .B(RESET), .Y(n4255));
AND2X1   g2372(.A(WX4702), .B(RESET), .Y(n4260));
AND2X1   g2373(.A(WX4704), .B(RESET), .Y(n4265));
AND2X1   g2374(.A(WX4706), .B(RESET), .Y(n4270));
AND2X1   g2375(.A(WX4708), .B(RESET), .Y(n4275));
AND2X1   g2376(.A(WX4710), .B(RESET), .Y(n4280));
AND2X1   g2377(.A(WX4712), .B(RESET), .Y(n4285));
AND2X1   g2378(.A(WX4714), .B(RESET), .Y(n4290));
XOR2X1   g2379(.A(CRC_OUT_6_31), .B(WX4778), .Y(n8046));
NOR2X1   g2380(.A(n8046), .B(n5827), .Y(CRC_OUT_6_0));
XOR2X1   g2381(.A(CRC_OUT_6_0), .B(WX4776), .Y(n8048));
NOR2X1   g2382(.A(n8048), .B(n5827), .Y(CRC_OUT_6_1));
XOR2X1   g2383(.A(CRC_OUT_6_1), .B(WX4774), .Y(n8050));
NOR2X1   g2384(.A(n8050), .B(n5827), .Y(CRC_OUT_6_2));
XOR2X1   g2385(.A(CRC_OUT_6_2), .B(WX4772), .Y(n8052));
NOR2X1   g2386(.A(n8052), .B(n5827), .Y(CRC_OUT_6_3));
XOR2X1   g2387(.A(CRC_OUT_6_31), .B(WX4770), .Y(n8054));
XOR2X1   g2388(.A(n8054), .B(CRC_OUT_6_3), .Y(n8055_1));
NOR2X1   g2389(.A(n8055_1), .B(n5827), .Y(CRC_OUT_6_4));
XOR2X1   g2390(.A(CRC_OUT_6_4), .B(WX4768), .Y(n8057));
NOR2X1   g2391(.A(n8057), .B(n5827), .Y(CRC_OUT_6_5));
XOR2X1   g2392(.A(CRC_OUT_6_5), .B(WX4766), .Y(n8059_1));
NOR2X1   g2393(.A(n8059_1), .B(n5827), .Y(CRC_OUT_6_6));
XOR2X1   g2394(.A(CRC_OUT_6_6), .B(WX4764), .Y(n8061));
NOR2X1   g2395(.A(n8061), .B(n5827), .Y(CRC_OUT_6_7));
XOR2X1   g2396(.A(CRC_OUT_6_7), .B(WX4762), .Y(n8063_1));
NOR2X1   g2397(.A(n8063_1), .B(n5827), .Y(CRC_OUT_6_8));
XOR2X1   g2398(.A(CRC_OUT_6_8), .B(WX4760), .Y(n8065));
NOR2X1   g2399(.A(n8065), .B(n5827), .Y(CRC_OUT_6_9));
XOR2X1   g2400(.A(CRC_OUT_6_9), .B(WX4758), .Y(n8067_1));
NOR2X1   g2401(.A(n8067_1), .B(n5827), .Y(CRC_OUT_6_10));
XOR2X1   g2402(.A(CRC_OUT_6_31), .B(WX4756), .Y(n8069));
XOR2X1   g2403(.A(n8069), .B(CRC_OUT_6_10), .Y(n8070));
NOR2X1   g2404(.A(n8070), .B(n5827), .Y(CRC_OUT_6_11));
XOR2X1   g2405(.A(CRC_OUT_6_11), .B(WX4754), .Y(n8072));
NOR2X1   g2406(.A(n8072), .B(n5827), .Y(CRC_OUT_6_12));
XOR2X1   g2407(.A(CRC_OUT_6_12), .B(WX4752), .Y(n8074));
NOR2X1   g2408(.A(n8074), .B(n5827), .Y(CRC_OUT_6_13));
XOR2X1   g2409(.A(CRC_OUT_6_13), .B(WX4750), .Y(n8076));
NOR2X1   g2410(.A(n8076), .B(n5827), .Y(CRC_OUT_6_14));
XOR2X1   g2411(.A(CRC_OUT_6_14), .B(WX4748), .Y(n8078));
NOR2X1   g2412(.A(n8078), .B(n5827), .Y(CRC_OUT_6_15));
XOR2X1   g2413(.A(CRC_OUT_6_31), .B(WX4746), .Y(n8080));
XOR2X1   g2414(.A(n8080), .B(CRC_OUT_6_15), .Y(n8081));
NOR2X1   g2415(.A(n8081), .B(n5827), .Y(CRC_OUT_6_16));
XOR2X1   g2416(.A(CRC_OUT_6_16), .B(WX4744), .Y(n8083_1));
NOR2X1   g2417(.A(n8083_1), .B(n5827), .Y(CRC_OUT_6_17));
XOR2X1   g2418(.A(CRC_OUT_6_17), .B(WX4742), .Y(n8085));
NOR2X1   g2419(.A(n8085), .B(n5827), .Y(CRC_OUT_6_18));
XOR2X1   g2420(.A(CRC_OUT_6_18), .B(WX4740), .Y(n8087_1));
NOR2X1   g2421(.A(n8087_1), .B(n5827), .Y(CRC_OUT_6_19));
XOR2X1   g2422(.A(CRC_OUT_6_19), .B(WX4738), .Y(n8089));
NOR2X1   g2423(.A(n8089), .B(n5827), .Y(CRC_OUT_6_20));
XOR2X1   g2424(.A(CRC_OUT_6_20), .B(WX4736), .Y(n8091_1));
NOR2X1   g2425(.A(n8091_1), .B(n5827), .Y(CRC_OUT_6_21));
XOR2X1   g2426(.A(CRC_OUT_6_21), .B(WX4734), .Y(n8093));
NOR2X1   g2427(.A(n8093), .B(n5827), .Y(CRC_OUT_6_22));
XOR2X1   g2428(.A(CRC_OUT_6_22), .B(WX4732), .Y(n8095_1));
NOR2X1   g2429(.A(n8095_1), .B(n5827), .Y(CRC_OUT_6_23));
XOR2X1   g2430(.A(CRC_OUT_6_23), .B(WX4730), .Y(n8097));
NOR2X1   g2431(.A(n8097), .B(n5827), .Y(CRC_OUT_6_24));
XOR2X1   g2432(.A(CRC_OUT_6_24), .B(WX4728), .Y(n8099_1));
NOR2X1   g2433(.A(n8099_1), .B(n5827), .Y(CRC_OUT_6_25));
XOR2X1   g2434(.A(CRC_OUT_6_25), .B(WX4726), .Y(n8101));
NOR2X1   g2435(.A(n8101), .B(n5827), .Y(CRC_OUT_6_26));
XOR2X1   g2436(.A(CRC_OUT_6_26), .B(WX4724), .Y(n8103_1));
NOR2X1   g2437(.A(n8103_1), .B(n5827), .Y(CRC_OUT_6_27));
XOR2X1   g2438(.A(CRC_OUT_6_27), .B(WX4722), .Y(n8105));
NOR2X1   g2439(.A(n8105), .B(n5827), .Y(CRC_OUT_6_28));
XOR2X1   g2440(.A(CRC_OUT_6_28), .B(WX4720), .Y(n8107_1));
NOR2X1   g2441(.A(n8107_1), .B(n5827), .Y(CRC_OUT_6_29));
XOR2X1   g2442(.A(CRC_OUT_6_29), .B(WX4718), .Y(n8109));
NOR2X1   g2443(.A(n8109), .B(n5827), .Y(CRC_OUT_6_30));
XOR2X1   g2444(.A(CRC_OUT_6_30), .B(WX4716), .Y(n8111_1));
NOR2X1   g2445(.A(n8111_1), .B(n5827), .Y(CRC_OUT_6_31));
AND2X1   g2446(.A(WX5659), .B(RESET), .Y(n4423));
AND2X1   g2447(.A(WX5661), .B(RESET), .Y(n4428));
AND2X1   g2448(.A(WX5663), .B(RESET), .Y(n4433));
AND2X1   g2449(.A(WX5665), .B(RESET), .Y(n4438));
AND2X1   g2450(.A(WX5667), .B(RESET), .Y(n4443));
AND2X1   g2451(.A(WX5669), .B(RESET), .Y(n4448));
AND2X1   g2452(.A(WX5671), .B(RESET), .Y(n4453));
AND2X1   g2453(.A(WX5673), .B(RESET), .Y(n4458));
AND2X1   g2454(.A(WX5675), .B(RESET), .Y(n4463));
AND2X1   g2455(.A(WX5677), .B(RESET), .Y(n4468));
AND2X1   g2456(.A(WX5679), .B(RESET), .Y(n4473));
AND2X1   g2457(.A(WX5681), .B(RESET), .Y(n4478));
AND2X1   g2458(.A(WX5683), .B(RESET), .Y(n4483));
AND2X1   g2459(.A(WX5685), .B(RESET), .Y(n4488));
AND2X1   g2460(.A(WX5687), .B(RESET), .Y(n4493));
AND2X1   g2461(.A(WX5689), .B(RESET), .Y(n4498));
AND2X1   g2462(.A(WX5691), .B(RESET), .Y(n4503));
AND2X1   g2463(.A(WX5693), .B(RESET), .Y(n4508));
AND2X1   g2464(.A(WX5695), .B(RESET), .Y(n4513));
AND2X1   g2465(.A(WX5697), .B(RESET), .Y(n4518));
AND2X1   g2466(.A(WX5699), .B(RESET), .Y(n4523));
AND2X1   g2467(.A(WX5701), .B(RESET), .Y(n4528));
AND2X1   g2468(.A(WX5703), .B(RESET), .Y(n4533));
AND2X1   g2469(.A(WX5705), .B(RESET), .Y(n4538));
AND2X1   g2470(.A(WX5707), .B(RESET), .Y(n4543));
AND2X1   g2471(.A(WX5709), .B(RESET), .Y(n4548));
AND2X1   g2472(.A(WX5711), .B(RESET), .Y(n4553));
AND2X1   g2473(.A(WX5713), .B(RESET), .Y(n4558));
AND2X1   g2474(.A(WX5715), .B(RESET), .Y(n4563));
AND2X1   g2475(.A(WX5717), .B(RESET), .Y(n4568));
AND2X1   g2476(.A(WX5719), .B(RESET), .Y(n4573));
NOR2X1   g2477(.A(WX5657), .B(n5827), .Y(n4578));
INVX1    g2478(.A(CRC_OUT_5_31), .Y(n8145_1));
XOR2X1   g2479(.A(WX7110), .B(TM1), .Y(n8146));
XOR2X1   g2480(.A(n8146), .B(WX7174), .Y(n8147));
INVX1    g2481(.A(WX7238), .Y(n8148));
XOR2X1   g2482(.A(WX7302), .B(n8148), .Y(n8149));
XOR2X1   g2483(.A(n8149), .B(n8147), .Y(n8150_1));
MX2X1    g2484(.A(n8145_1), .B(n8150_1), .S0(n5539), .Y(n8152));
INVX1    g2485(.A(WX5657), .Y(n8153));
MX2X1    g2486(.A(n8153), .B(n7571), .S0(n5539), .Y(n8154));
MX2X1    g2487(.A(n8152), .B(n8154), .S0(TM1), .Y(n8155_1));
NOR2X1   g2488(.A(n8155_1), .B(n5827), .Y(n4583));
INVX1    g2489(.A(CRC_OUT_5_30), .Y(n8157));
XOR2X1   g2490(.A(WX7112), .B(TM1), .Y(n8158));
XOR2X1   g2491(.A(n8158), .B(WX7176), .Y(n8159));
INVX1    g2492(.A(WX7240), .Y(n8160_1));
XOR2X1   g2493(.A(WX7304), .B(n8160_1), .Y(n8161));
XOR2X1   g2494(.A(n8161), .B(n8159), .Y(n8162));
MX2X1    g2495(.A(n8157), .B(n8162), .S0(n5539), .Y(n8164));
INVX1    g2496(.A(WX5659), .Y(n8165_1));
MX2X1    g2497(.A(n8165_1), .B(n7583), .S0(n5539), .Y(n8166));
MX2X1    g2498(.A(n8164), .B(n8166), .S0(TM1), .Y(n8167));
NOR2X1   g2499(.A(n8167), .B(n5827), .Y(n4588));
INVX1    g2500(.A(CRC_OUT_5_29), .Y(n8169));
XOR2X1   g2501(.A(WX7114), .B(TM1), .Y(n8170_1));
XOR2X1   g2502(.A(n8170_1), .B(WX7178), .Y(n8171));
INVX1    g2503(.A(WX7242), .Y(n8172));
XOR2X1   g2504(.A(WX7306), .B(n8172), .Y(n8173));
XOR2X1   g2505(.A(n8173), .B(n8171), .Y(n8174));
MX2X1    g2506(.A(n8169), .B(n8174), .S0(n5539), .Y(n8176));
INVX1    g2507(.A(WX5661), .Y(n8177));
MX2X1    g2508(.A(n8177), .B(n7595), .S0(n5539), .Y(n8178));
MX2X1    g2509(.A(n8176), .B(n8178), .S0(TM1), .Y(n8179));
NOR2X1   g2510(.A(n8179), .B(n5827), .Y(n4593));
INVX1    g2511(.A(CRC_OUT_5_28), .Y(n8181));
XOR2X1   g2512(.A(WX7116), .B(TM1), .Y(n8182));
XOR2X1   g2513(.A(n8182), .B(WX7180), .Y(n8183));
INVX1    g2514(.A(WX7244), .Y(n8184));
XOR2X1   g2515(.A(WX7308), .B(n8184), .Y(n8185_1));
XOR2X1   g2516(.A(n8185_1), .B(n8183), .Y(n8186));
MX2X1    g2517(.A(n8181), .B(n8186), .S0(n5539), .Y(n8188));
INVX1    g2518(.A(WX5663), .Y(n8189));
MX2X1    g2519(.A(n8189), .B(n7607_1), .S0(n5539), .Y(n8190_1));
MX2X1    g2520(.A(n8188), .B(n8190_1), .S0(TM1), .Y(n8191));
NOR2X1   g2521(.A(n8191), .B(n5827), .Y(n4598));
INVX1    g2522(.A(CRC_OUT_5_27), .Y(n8193));
XOR2X1   g2523(.A(WX7118), .B(TM1), .Y(n8194));
XOR2X1   g2524(.A(n8194), .B(WX7182), .Y(n8195_1));
INVX1    g2525(.A(WX7246), .Y(n8196));
XOR2X1   g2526(.A(WX7310), .B(n8196), .Y(n8197));
XOR2X1   g2527(.A(n8197), .B(n8195_1), .Y(n8198));
MX2X1    g2528(.A(n8193), .B(n8198), .S0(n5539), .Y(n8200_1));
INVX1    g2529(.A(WX5665), .Y(n8201));
MX2X1    g2530(.A(n8201), .B(n7619), .S0(n5539), .Y(n8202));
MX2X1    g2531(.A(n8200_1), .B(n8202), .S0(TM1), .Y(n8203));
NOR2X1   g2532(.A(n8203), .B(n5827), .Y(n4603));
INVX1    g2533(.A(CRC_OUT_5_26), .Y(n8205_1));
XOR2X1   g2534(.A(WX7120), .B(TM1), .Y(n8206));
XOR2X1   g2535(.A(n8206), .B(WX7184), .Y(n8207));
INVX1    g2536(.A(WX7248), .Y(n8208));
XOR2X1   g2537(.A(WX7312), .B(n8208), .Y(n8209));
XOR2X1   g2538(.A(n8209), .B(n8207), .Y(n8210_1));
MX2X1    g2539(.A(n8205_1), .B(n8210_1), .S0(n5539), .Y(n8212));
INVX1    g2540(.A(WX5667), .Y(n8213));
MX2X1    g2541(.A(n8213), .B(n7631), .S0(n5539), .Y(n8214));
MX2X1    g2542(.A(n8212), .B(n8214), .S0(TM1), .Y(n8215_1));
NOR2X1   g2543(.A(n8215_1), .B(n5827), .Y(n4608));
INVX1    g2544(.A(CRC_OUT_5_25), .Y(n8217));
XOR2X1   g2545(.A(WX7122), .B(TM1), .Y(n8218));
XOR2X1   g2546(.A(n8218), .B(WX7186), .Y(n8219));
INVX1    g2547(.A(WX7250), .Y(n8220_1));
XOR2X1   g2548(.A(WX7314), .B(n8220_1), .Y(n8221));
XOR2X1   g2549(.A(n8221), .B(n8219), .Y(n8222));
MX2X1    g2550(.A(n8217), .B(n8222), .S0(n5539), .Y(n8224));
INVX1    g2551(.A(WX5669), .Y(n8225_1));
MX2X1    g2552(.A(n8225_1), .B(n7643), .S0(n5539), .Y(n8226));
MX2X1    g2553(.A(n8224), .B(n8226), .S0(TM1), .Y(n8227));
NOR2X1   g2554(.A(n8227), .B(n5827), .Y(n4613));
INVX1    g2555(.A(CRC_OUT_5_24), .Y(n8229));
XOR2X1   g2556(.A(WX7124), .B(TM1), .Y(n8230_1));
XOR2X1   g2557(.A(n8230_1), .B(WX7188), .Y(n8231));
INVX1    g2558(.A(WX7252), .Y(n8232));
XOR2X1   g2559(.A(WX7316), .B(n8232), .Y(n8233));
XOR2X1   g2560(.A(n8233), .B(n8231), .Y(n8234));
MX2X1    g2561(.A(n8229), .B(n8234), .S0(n5539), .Y(n8236));
INVX1    g2562(.A(WX5671), .Y(n8237));
MX2X1    g2563(.A(n8237), .B(n7655), .S0(n5539), .Y(n8238));
MX2X1    g2564(.A(n8236), .B(n8238), .S0(TM1), .Y(n8239));
NOR2X1   g2565(.A(n8239), .B(n5827), .Y(n4618));
INVX1    g2566(.A(CRC_OUT_5_23), .Y(n8241));
XOR2X1   g2567(.A(WX7126), .B(TM1), .Y(n8242));
XOR2X1   g2568(.A(n8242), .B(WX7190), .Y(n8243));
INVX1    g2569(.A(WX7254), .Y(n8244));
XOR2X1   g2570(.A(WX7318), .B(n8244), .Y(n8245_1));
XOR2X1   g2571(.A(n8245_1), .B(n8243), .Y(n8246));
MX2X1    g2572(.A(n8241), .B(n8246), .S0(n5539), .Y(n8248));
INVX1    g2573(.A(WX5673), .Y(n8249));
MX2X1    g2574(.A(n8249), .B(n7667_1), .S0(n5539), .Y(n8250_1));
MX2X1    g2575(.A(n8248), .B(n8250_1), .S0(TM1), .Y(n8251));
NOR2X1   g2576(.A(n8251), .B(n5827), .Y(n4623));
INVX1    g2577(.A(CRC_OUT_5_22), .Y(n8253));
XOR2X1   g2578(.A(WX7128), .B(TM1), .Y(n8254));
XOR2X1   g2579(.A(n8254), .B(WX7192), .Y(n8255_1));
INVX1    g2580(.A(WX7256), .Y(n8256));
XOR2X1   g2581(.A(WX7320), .B(n8256), .Y(n8257));
XOR2X1   g2582(.A(n8257), .B(n8255_1), .Y(n8258));
MX2X1    g2583(.A(n8253), .B(n8258), .S0(n5539), .Y(n8260_1));
INVX1    g2584(.A(WX5675), .Y(n8261));
MX2X1    g2585(.A(n8261), .B(n7679), .S0(n5539), .Y(n8262));
MX2X1    g2586(.A(n8260_1), .B(n8262), .S0(TM1), .Y(n8263));
NOR2X1   g2587(.A(n8263), .B(n5827), .Y(n4628));
INVX1    g2588(.A(CRC_OUT_5_21), .Y(n8265_1));
XOR2X1   g2589(.A(WX7130), .B(TM1), .Y(n8266));
XOR2X1   g2590(.A(n8266), .B(WX7194), .Y(n8267));
INVX1    g2591(.A(WX7258), .Y(n8268));
XOR2X1   g2592(.A(WX7322), .B(n8268), .Y(n8269));
XOR2X1   g2593(.A(n8269), .B(n8267), .Y(n8270_1));
MX2X1    g2594(.A(n8265_1), .B(n8270_1), .S0(n5539), .Y(n8272));
INVX1    g2595(.A(WX5677), .Y(n8273));
MX2X1    g2596(.A(n8273), .B(n7691), .S0(n5539), .Y(n8274));
MX2X1    g2597(.A(n8272), .B(n8274), .S0(TM1), .Y(n8275_1));
NOR2X1   g2598(.A(n8275_1), .B(n5827), .Y(n4633));
INVX1    g2599(.A(CRC_OUT_5_20), .Y(n8277));
XOR2X1   g2600(.A(WX7132), .B(TM1), .Y(n8278));
XOR2X1   g2601(.A(n8278), .B(WX7196), .Y(n8279));
INVX1    g2602(.A(WX7260), .Y(n8280_1));
XOR2X1   g2603(.A(WX7324), .B(n8280_1), .Y(n8281));
XOR2X1   g2604(.A(n8281), .B(n8279), .Y(n8282));
MX2X1    g2605(.A(n8277), .B(n8282), .S0(n5539), .Y(n8284));
INVX1    g2606(.A(WX5679), .Y(n8285_1));
MX2X1    g2607(.A(n8285_1), .B(n7703), .S0(n5539), .Y(n8286));
MX2X1    g2608(.A(n8284), .B(n8286), .S0(TM1), .Y(n8287));
NOR2X1   g2609(.A(n8287), .B(n5827), .Y(n4638));
INVX1    g2610(.A(CRC_OUT_5_19), .Y(n8289));
XOR2X1   g2611(.A(WX7134), .B(TM1), .Y(n8290_1));
XOR2X1   g2612(.A(n8290_1), .B(WX7198), .Y(n8291));
INVX1    g2613(.A(WX7262), .Y(n8292));
XOR2X1   g2614(.A(WX7326), .B(n8292), .Y(n8293));
XOR2X1   g2615(.A(n8293), .B(n8291), .Y(n8294));
MX2X1    g2616(.A(n8289), .B(n8294), .S0(n5539), .Y(n8296));
INVX1    g2617(.A(WX5681), .Y(n8297));
MX2X1    g2618(.A(n8297), .B(n7715), .S0(n5539), .Y(n8298));
MX2X1    g2619(.A(n8296), .B(n8298), .S0(TM1), .Y(n8299));
NOR2X1   g2620(.A(n8299), .B(n5827), .Y(n4643));
INVX1    g2621(.A(CRC_OUT_5_18), .Y(n8301));
XOR2X1   g2622(.A(WX7136), .B(TM1), .Y(n8302));
XOR2X1   g2623(.A(n8302), .B(WX7200), .Y(n8303));
INVX1    g2624(.A(WX7264), .Y(n8304));
XOR2X1   g2625(.A(WX7328), .B(n8304), .Y(n8305_1));
XOR2X1   g2626(.A(n8305_1), .B(n8303), .Y(n8306));
MX2X1    g2627(.A(n8301), .B(n8306), .S0(n5539), .Y(n8308));
INVX1    g2628(.A(WX5683), .Y(n8309));
MX2X1    g2629(.A(n8309), .B(n7727_1), .S0(n5539), .Y(n8310_1));
MX2X1    g2630(.A(n8308), .B(n8310_1), .S0(TM1), .Y(n8311));
NOR2X1   g2631(.A(n8311), .B(n5827), .Y(n4648));
INVX1    g2632(.A(CRC_OUT_5_17), .Y(n8313));
XOR2X1   g2633(.A(WX7138), .B(TM1), .Y(n8314));
XOR2X1   g2634(.A(n8314), .B(WX7202), .Y(n8315_1));
INVX1    g2635(.A(WX7266), .Y(n8316));
XOR2X1   g2636(.A(WX7330), .B(n8316), .Y(n8317));
XOR2X1   g2637(.A(n8317), .B(n8315_1), .Y(n8318));
MX2X1    g2638(.A(n8313), .B(n8318), .S0(n5539), .Y(n8320_1));
INVX1    g2639(.A(WX5685), .Y(n8321));
MX2X1    g2640(.A(n8321), .B(n7739), .S0(n5539), .Y(n8322));
MX2X1    g2641(.A(n8320_1), .B(n8322), .S0(TM1), .Y(n8323));
NOR2X1   g2642(.A(n8323), .B(n5827), .Y(n4653));
INVX1    g2643(.A(CRC_OUT_5_16), .Y(n8325_1));
XOR2X1   g2644(.A(WX7140), .B(TM1), .Y(n8326));
XOR2X1   g2645(.A(n8326), .B(WX7204), .Y(n8327));
INVX1    g2646(.A(WX7268), .Y(n8328));
XOR2X1   g2647(.A(WX7332), .B(n8328), .Y(n8329));
XOR2X1   g2648(.A(n8329), .B(n8327), .Y(n8330_1));
MX2X1    g2649(.A(n8325_1), .B(n8330_1), .S0(n5539), .Y(n8332));
INVX1    g2650(.A(WX5687), .Y(n8333));
MX2X1    g2651(.A(n8333), .B(n7751), .S0(n5539), .Y(n8334));
MX2X1    g2652(.A(n8332), .B(n8334), .S0(TM1), .Y(n8335_1));
NOR2X1   g2653(.A(n8335_1), .B(n5827), .Y(n4658));
INVX1    g2654(.A(CRC_OUT_5_15), .Y(n8337));
XOR2X1   g2655(.A(WX7142), .B(TM0), .Y(n8338));
XOR2X1   g2656(.A(n8338), .B(WX7206), .Y(n8339));
INVX1    g2657(.A(WX7270), .Y(n8340_1));
XOR2X1   g2658(.A(WX7334), .B(n8340_1), .Y(n8341));
XOR2X1   g2659(.A(n8341), .B(n8339), .Y(n8342));
MX2X1    g2660(.A(n8337), .B(n8342), .S0(n5539), .Y(n8344));
INVX1    g2661(.A(WX5689), .Y(n8345_1));
MX2X1    g2662(.A(n8345_1), .B(n7763), .S0(n5539), .Y(n8346));
MX2X1    g2663(.A(n8344), .B(n8346), .S0(TM1), .Y(n8347));
NOR2X1   g2664(.A(n8347), .B(n5827), .Y(n4663));
INVX1    g2665(.A(CRC_OUT_5_14), .Y(n8349));
XOR2X1   g2666(.A(WX7144), .B(TM0), .Y(n8350_1));
XOR2X1   g2667(.A(n8350_1), .B(WX7208), .Y(n8351));
INVX1    g2668(.A(WX7272), .Y(n8352));
XOR2X1   g2669(.A(WX7336), .B(n8352), .Y(n8353));
XOR2X1   g2670(.A(n8353), .B(n8351), .Y(n8354));
MX2X1    g2671(.A(n8349), .B(n8354), .S0(n5539), .Y(n8356));
INVX1    g2672(.A(WX5691), .Y(n8357));
MX2X1    g2673(.A(n8357), .B(n7775), .S0(n5539), .Y(n8358));
MX2X1    g2674(.A(n8356), .B(n8358), .S0(TM1), .Y(n8359));
NOR2X1   g2675(.A(n8359), .B(n5827), .Y(n4668));
INVX1    g2676(.A(CRC_OUT_5_13), .Y(n8361));
XOR2X1   g2677(.A(WX7146), .B(TM0), .Y(n8362));
XOR2X1   g2678(.A(n8362), .B(WX7210), .Y(n8363));
INVX1    g2679(.A(WX7274), .Y(n8364));
XOR2X1   g2680(.A(WX7338), .B(n8364), .Y(n8365_1));
XOR2X1   g2681(.A(n8365_1), .B(n8363), .Y(n8366));
MX2X1    g2682(.A(n8361), .B(n8366), .S0(n5539), .Y(n8368));
INVX1    g2683(.A(WX5693), .Y(n8369));
MX2X1    g2684(.A(n8369), .B(n7787_1), .S0(n5539), .Y(n8370_1));
MX2X1    g2685(.A(n8368), .B(n8370_1), .S0(TM1), .Y(n8371));
NOR2X1   g2686(.A(n8371), .B(n5827), .Y(n4673));
INVX1    g2687(.A(CRC_OUT_5_12), .Y(n8373));
XOR2X1   g2688(.A(WX7148), .B(TM0), .Y(n8374));
XOR2X1   g2689(.A(n8374), .B(WX7212), .Y(n8375_1));
INVX1    g2690(.A(WX7276), .Y(n8376));
XOR2X1   g2691(.A(WX7340), .B(n8376), .Y(n8377));
XOR2X1   g2692(.A(n8377), .B(n8375_1), .Y(n8378));
MX2X1    g2693(.A(n8373), .B(n8378), .S0(n5539), .Y(n8380_1));
INVX1    g2694(.A(WX5695), .Y(n8381));
MX2X1    g2695(.A(n8381), .B(n7799), .S0(n5539), .Y(n8382));
MX2X1    g2696(.A(n8380_1), .B(n8382), .S0(TM1), .Y(n8383));
NOR2X1   g2697(.A(n8383), .B(n5827), .Y(n4678));
INVX1    g2698(.A(CRC_OUT_5_11), .Y(n8385_1));
XOR2X1   g2699(.A(WX7150), .B(TM0), .Y(n8386));
XOR2X1   g2700(.A(n8386), .B(WX7214), .Y(n8387));
INVX1    g2701(.A(WX7278), .Y(n8388));
XOR2X1   g2702(.A(WX7342), .B(n8388), .Y(n8389));
XOR2X1   g2703(.A(n8389), .B(n8387), .Y(n8390_1));
MX2X1    g2704(.A(n8385_1), .B(n8390_1), .S0(n5539), .Y(n8392));
INVX1    g2705(.A(WX5697), .Y(n8393));
MX2X1    g2706(.A(n8393), .B(n7811), .S0(n5539), .Y(n8394));
MX2X1    g2707(.A(n8392), .B(n8394), .S0(TM1), .Y(n8395_1));
NOR2X1   g2708(.A(n8395_1), .B(n5827), .Y(n4683));
INVX1    g2709(.A(CRC_OUT_5_10), .Y(n8397));
XOR2X1   g2710(.A(WX7152), .B(TM0), .Y(n8398));
XOR2X1   g2711(.A(n8398), .B(WX7216), .Y(n8399));
INVX1    g2712(.A(WX7280), .Y(n8400_1));
XOR2X1   g2713(.A(WX7344), .B(n8400_1), .Y(n8401));
XOR2X1   g2714(.A(n8401), .B(n8399), .Y(n8402));
MX2X1    g2715(.A(n8397), .B(n8402), .S0(n5539), .Y(n8404));
INVX1    g2716(.A(WX5699), .Y(n8405_1));
MX2X1    g2717(.A(n8405_1), .B(n7823), .S0(n5539), .Y(n8406));
MX2X1    g2718(.A(n8404), .B(n8406), .S0(TM1), .Y(n8407));
NOR2X1   g2719(.A(n8407), .B(n5827), .Y(n4688));
INVX1    g2720(.A(CRC_OUT_5_9), .Y(n8409));
XOR2X1   g2721(.A(WX7154), .B(TM0), .Y(n8410_1));
XOR2X1   g2722(.A(n8410_1), .B(WX7218), .Y(n8411));
INVX1    g2723(.A(WX7282), .Y(n8412));
XOR2X1   g2724(.A(WX7346), .B(n8412), .Y(n8413));
XOR2X1   g2725(.A(n8413), .B(n8411), .Y(n8414));
MX2X1    g2726(.A(n8409), .B(n8414), .S0(n5539), .Y(n8416));
INVX1    g2727(.A(WX5701), .Y(n8417));
MX2X1    g2728(.A(n8417), .B(n7835), .S0(n5539), .Y(n8418));
MX2X1    g2729(.A(n8416), .B(n8418), .S0(TM1), .Y(n8419));
NOR2X1   g2730(.A(n8419), .B(n5827), .Y(n4693));
INVX1    g2731(.A(CRC_OUT_5_8), .Y(n8421));
XOR2X1   g2732(.A(WX7156), .B(TM0), .Y(n8422));
XOR2X1   g2733(.A(n8422), .B(WX7220), .Y(n8423));
INVX1    g2734(.A(WX7284), .Y(n8424));
XOR2X1   g2735(.A(WX7348), .B(n8424), .Y(n8425_1));
XOR2X1   g2736(.A(n8425_1), .B(n8423), .Y(n8426));
MX2X1    g2737(.A(n8421), .B(n8426), .S0(n5539), .Y(n8428));
INVX1    g2738(.A(WX5703), .Y(n8429));
MX2X1    g2739(.A(n8429), .B(n7847_1), .S0(n5539), .Y(n8430_1));
MX2X1    g2740(.A(n8428), .B(n8430_1), .S0(TM1), .Y(n8431));
NOR2X1   g2741(.A(n8431), .B(n5827), .Y(n4698));
INVX1    g2742(.A(CRC_OUT_5_7), .Y(n8433));
XOR2X1   g2743(.A(WX7158), .B(TM0), .Y(n8434));
XOR2X1   g2744(.A(n8434), .B(WX7222), .Y(n8435_1));
INVX1    g2745(.A(WX7286), .Y(n8436));
XOR2X1   g2746(.A(WX7350), .B(n8436), .Y(n8437));
XOR2X1   g2747(.A(n8437), .B(n8435_1), .Y(n8438));
MX2X1    g2748(.A(n8433), .B(n8438), .S0(n5539), .Y(n8440_1));
INVX1    g2749(.A(WX5705), .Y(n8441));
MX2X1    g2750(.A(n8441), .B(n7859), .S0(n5539), .Y(n8442));
MX2X1    g2751(.A(n8440_1), .B(n8442), .S0(TM1), .Y(n8443));
NOR2X1   g2752(.A(n8443), .B(n5827), .Y(n4703));
INVX1    g2753(.A(CRC_OUT_5_6), .Y(n8445_1));
XOR2X1   g2754(.A(WX7160), .B(TM0), .Y(n8446));
XOR2X1   g2755(.A(n8446), .B(WX7224), .Y(n8447));
INVX1    g2756(.A(WX7288), .Y(n8448));
XOR2X1   g2757(.A(WX7352), .B(n8448), .Y(n8449));
XOR2X1   g2758(.A(n8449), .B(n8447), .Y(n8450_1));
MX2X1    g2759(.A(n8445_1), .B(n8450_1), .S0(n5539), .Y(n8452));
INVX1    g2760(.A(WX5707), .Y(n8453));
MX2X1    g2761(.A(n8453), .B(n7871), .S0(n5539), .Y(n8454));
MX2X1    g2762(.A(n8452), .B(n8454), .S0(TM1), .Y(n8455_1));
NOR2X1   g2763(.A(n8455_1), .B(n5827), .Y(n4708));
INVX1    g2764(.A(CRC_OUT_5_5), .Y(n8457));
XOR2X1   g2765(.A(WX7162), .B(TM0), .Y(n8458));
XOR2X1   g2766(.A(n8458), .B(WX7226), .Y(n8459));
INVX1    g2767(.A(WX7290), .Y(n8460_1));
XOR2X1   g2768(.A(WX7354), .B(n8460_1), .Y(n8461));
XOR2X1   g2769(.A(n8461), .B(n8459), .Y(n8462));
MX2X1    g2770(.A(n8457), .B(n8462), .S0(n5539), .Y(n8464));
INVX1    g2771(.A(WX5709), .Y(n8465_1));
MX2X1    g2772(.A(n8465_1), .B(n7883), .S0(n5539), .Y(n8466));
MX2X1    g2773(.A(n8464), .B(n8466), .S0(TM1), .Y(n8467));
NOR2X1   g2774(.A(n8467), .B(n5827), .Y(n4713));
INVX1    g2775(.A(CRC_OUT_5_4), .Y(n8469));
XOR2X1   g2776(.A(WX7164), .B(TM0), .Y(n8470_1));
XOR2X1   g2777(.A(n8470_1), .B(WX7228), .Y(n8471));
INVX1    g2778(.A(WX7292), .Y(n8472));
XOR2X1   g2779(.A(WX7356), .B(n8472), .Y(n8473));
XOR2X1   g2780(.A(n8473), .B(n8471), .Y(n8474));
MX2X1    g2781(.A(n8469), .B(n8474), .S0(n5539), .Y(n8476));
INVX1    g2782(.A(WX5711), .Y(n8477));
MX2X1    g2783(.A(n8477), .B(n7895), .S0(n5539), .Y(n8478));
MX2X1    g2784(.A(n8476), .B(n8478), .S0(TM1), .Y(n8479));
NOR2X1   g2785(.A(n8479), .B(n5827), .Y(n4718));
INVX1    g2786(.A(CRC_OUT_5_3), .Y(n8481));
XOR2X1   g2787(.A(WX7166), .B(TM0), .Y(n8482));
XOR2X1   g2788(.A(n8482), .B(WX7230), .Y(n8483));
INVX1    g2789(.A(WX7294), .Y(n8484));
XOR2X1   g2790(.A(WX7358), .B(n8484), .Y(n8485_1));
XOR2X1   g2791(.A(n8485_1), .B(n8483), .Y(n8486));
MX2X1    g2792(.A(n8481), .B(n8486), .S0(n5539), .Y(n8488));
INVX1    g2793(.A(WX5713), .Y(n8489));
MX2X1    g2794(.A(n8489), .B(n7907_1), .S0(n5539), .Y(n8490_1));
MX2X1    g2795(.A(n8488), .B(n8490_1), .S0(TM1), .Y(n8491));
NOR2X1   g2796(.A(n8491), .B(n5827), .Y(n4723));
INVX1    g2797(.A(CRC_OUT_5_2), .Y(n8493));
XOR2X1   g2798(.A(WX7168), .B(TM0), .Y(n8494));
XOR2X1   g2799(.A(n8494), .B(WX7232), .Y(n8495_1));
INVX1    g2800(.A(WX7296), .Y(n8496));
XOR2X1   g2801(.A(WX7360), .B(n8496), .Y(n8497));
XOR2X1   g2802(.A(n8497), .B(n8495_1), .Y(n8498));
MX2X1    g2803(.A(n8493), .B(n8498), .S0(n5539), .Y(n8500_1));
INVX1    g2804(.A(WX5715), .Y(n8501));
MX2X1    g2805(.A(n8501), .B(n7919), .S0(n5539), .Y(n8502));
MX2X1    g2806(.A(n8500_1), .B(n8502), .S0(TM1), .Y(n8503));
NOR2X1   g2807(.A(n8503), .B(n5827), .Y(n4728));
INVX1    g2808(.A(CRC_OUT_5_1), .Y(n8505_1));
XOR2X1   g2809(.A(WX7170), .B(TM0), .Y(n8506));
XOR2X1   g2810(.A(n8506), .B(WX7234), .Y(n8507));
INVX1    g2811(.A(WX7298), .Y(n8508));
XOR2X1   g2812(.A(WX7362), .B(n8508), .Y(n8509));
XOR2X1   g2813(.A(n8509), .B(n8507), .Y(n8510_1));
MX2X1    g2814(.A(n8505_1), .B(n8510_1), .S0(n5539), .Y(n8512));
INVX1    g2815(.A(WX5717), .Y(n8513));
MX2X1    g2816(.A(n8513), .B(n7931), .S0(n5539), .Y(n8514));
MX2X1    g2817(.A(n8512), .B(n8514), .S0(TM1), .Y(n8515_1));
NOR2X1   g2818(.A(n8515_1), .B(n5827), .Y(n4733));
INVX1    g2819(.A(CRC_OUT_5_0), .Y(n8517));
XOR2X1   g2820(.A(WX7172), .B(TM0), .Y(n8518));
XOR2X1   g2821(.A(n8518), .B(WX7236), .Y(n8519));
INVX1    g2822(.A(WX7300), .Y(n8520_1));
XOR2X1   g2823(.A(WX7364), .B(n8520_1), .Y(n8521));
XOR2X1   g2824(.A(n8521), .B(n8519), .Y(n8522));
MX2X1    g2825(.A(n8517), .B(n8522), .S0(n5539), .Y(n8524));
INVX1    g2826(.A(WX5719), .Y(n8525_1));
MX2X1    g2827(.A(n8525_1), .B(n7943), .S0(n5539), .Y(n8526));
MX2X1    g2828(.A(n8524), .B(n8526), .S0(TM1), .Y(n8527));
NOR2X1   g2829(.A(n8527), .B(n5827), .Y(n4738));
AND2X1   g2830(.A(WX5817), .B(RESET), .Y(n4743));
AND2X1   g2831(.A(WX5819), .B(RESET), .Y(n4748));
AND2X1   g2832(.A(WX5821), .B(RESET), .Y(n4753));
AND2X1   g2833(.A(WX5823), .B(RESET), .Y(n4758));
AND2X1   g2834(.A(WX5825), .B(RESET), .Y(n4763));
AND2X1   g2835(.A(WX5827), .B(RESET), .Y(n4768));
AND2X1   g2836(.A(WX5829), .B(RESET), .Y(n4773));
AND2X1   g2837(.A(WX5831), .B(RESET), .Y(n4778));
AND2X1   g2838(.A(WX5833), .B(RESET), .Y(n4783));
AND2X1   g2839(.A(WX5835), .B(RESET), .Y(n4788));
AND2X1   g2840(.A(WX5837), .B(RESET), .Y(n4793));
AND2X1   g2841(.A(WX5839), .B(RESET), .Y(n4798));
AND2X1   g2842(.A(WX5841), .B(RESET), .Y(n4803));
AND2X1   g2843(.A(WX5843), .B(RESET), .Y(n4808));
AND2X1   g2844(.A(WX5845), .B(RESET), .Y(n4813));
AND2X1   g2845(.A(WX5847), .B(RESET), .Y(n4818));
AND2X1   g2846(.A(WX5849), .B(RESET), .Y(n4823));
AND2X1   g2847(.A(WX5851), .B(RESET), .Y(n4828));
AND2X1   g2848(.A(WX5853), .B(RESET), .Y(n4833));
AND2X1   g2849(.A(WX5855), .B(RESET), .Y(n4838));
AND2X1   g2850(.A(WX5857), .B(RESET), .Y(n4843));
AND2X1   g2851(.A(WX5859), .B(RESET), .Y(n4848));
AND2X1   g2852(.A(WX5861), .B(RESET), .Y(n4853));
AND2X1   g2853(.A(WX5863), .B(RESET), .Y(n4858));
AND2X1   g2854(.A(WX5865), .B(RESET), .Y(n4863));
AND2X1   g2855(.A(WX5867), .B(RESET), .Y(n4868));
AND2X1   g2856(.A(WX5869), .B(RESET), .Y(n4873));
AND2X1   g2857(.A(WX5871), .B(RESET), .Y(n4878));
AND2X1   g2858(.A(WX5873), .B(RESET), .Y(n4883));
AND2X1   g2859(.A(WX5875), .B(RESET), .Y(n4888));
AND2X1   g2860(.A(WX5877), .B(RESET), .Y(n4893));
AND2X1   g2861(.A(WX5879), .B(RESET), .Y(n4898));
AND2X1   g2862(.A(WX5881), .B(RESET), .Y(n4903));
AND2X1   g2863(.A(WX5883), .B(RESET), .Y(n4908));
AND2X1   g2864(.A(WX5885), .B(RESET), .Y(n4913));
AND2X1   g2865(.A(WX5887), .B(RESET), .Y(n4918));
AND2X1   g2866(.A(WX5889), .B(RESET), .Y(n4923));
AND2X1   g2867(.A(WX5891), .B(RESET), .Y(n4928));
AND2X1   g2868(.A(WX5893), .B(RESET), .Y(n4933));
AND2X1   g2869(.A(WX5895), .B(RESET), .Y(n4938));
AND2X1   g2870(.A(WX5897), .B(RESET), .Y(n4943));
AND2X1   g2871(.A(WX5899), .B(RESET), .Y(n4948));
AND2X1   g2872(.A(WX5901), .B(RESET), .Y(n4953));
AND2X1   g2873(.A(WX5903), .B(RESET), .Y(n4958));
AND2X1   g2874(.A(WX5905), .B(RESET), .Y(n4963));
AND2X1   g2875(.A(WX5907), .B(RESET), .Y(n4968));
AND2X1   g2876(.A(WX5909), .B(RESET), .Y(n4973));
AND2X1   g2877(.A(WX5911), .B(RESET), .Y(n4978));
AND2X1   g2878(.A(WX5913), .B(RESET), .Y(n4983));
AND2X1   g2879(.A(WX5915), .B(RESET), .Y(n4988));
AND2X1   g2880(.A(WX5917), .B(RESET), .Y(n4993));
AND2X1   g2881(.A(WX5919), .B(RESET), .Y(n4998));
AND2X1   g2882(.A(WX5921), .B(RESET), .Y(n5003));
AND2X1   g2883(.A(WX5923), .B(RESET), .Y(n5008));
AND2X1   g2884(.A(WX5925), .B(RESET), .Y(n5013));
AND2X1   g2885(.A(WX5927), .B(RESET), .Y(n5018));
AND2X1   g2886(.A(WX5929), .B(RESET), .Y(n5023));
AND2X1   g2887(.A(WX5931), .B(RESET), .Y(n5028));
AND2X1   g2888(.A(WX5933), .B(RESET), .Y(n5033));
AND2X1   g2889(.A(WX5935), .B(RESET), .Y(n5038));
AND2X1   g2890(.A(WX5937), .B(RESET), .Y(n5043));
AND2X1   g2891(.A(WX5939), .B(RESET), .Y(n5048));
AND2X1   g2892(.A(WX5941), .B(RESET), .Y(n5053));
AND2X1   g2893(.A(WX5943), .B(RESET), .Y(n5058));
AND2X1   g2894(.A(WX5945), .B(RESET), .Y(n5063));
AND2X1   g2895(.A(WX5947), .B(RESET), .Y(n5068));
AND2X1   g2896(.A(WX5949), .B(RESET), .Y(n5073));
AND2X1   g2897(.A(WX5951), .B(RESET), .Y(n5078));
AND2X1   g2898(.A(WX5953), .B(RESET), .Y(n5083));
AND2X1   g2899(.A(WX5955), .B(RESET), .Y(n5088));
AND2X1   g2900(.A(WX5957), .B(RESET), .Y(n5093));
AND2X1   g2901(.A(WX5959), .B(RESET), .Y(n5098));
AND2X1   g2902(.A(WX5961), .B(RESET), .Y(n5103));
AND2X1   g2903(.A(WX5963), .B(RESET), .Y(n5108));
AND2X1   g2904(.A(WX5965), .B(RESET), .Y(n5113));
AND2X1   g2905(.A(WX5967), .B(RESET), .Y(n5118));
AND2X1   g2906(.A(WX5969), .B(RESET), .Y(n5123));
AND2X1   g2907(.A(WX5971), .B(RESET), .Y(n5128));
AND2X1   g2908(.A(WX5973), .B(RESET), .Y(n5133));
AND2X1   g2909(.A(WX5975), .B(RESET), .Y(n5138));
AND2X1   g2910(.A(WX5977), .B(RESET), .Y(n5143));
AND2X1   g2911(.A(WX5979), .B(RESET), .Y(n5148));
AND2X1   g2912(.A(WX5981), .B(RESET), .Y(n5153));
AND2X1   g2913(.A(WX5983), .B(RESET), .Y(n5158));
AND2X1   g2914(.A(WX5985), .B(RESET), .Y(n5163));
AND2X1   g2915(.A(WX5987), .B(RESET), .Y(n5168));
AND2X1   g2916(.A(WX5989), .B(RESET), .Y(n5173));
AND2X1   g2917(.A(WX5991), .B(RESET), .Y(n5178));
AND2X1   g2918(.A(WX5993), .B(RESET), .Y(n5183));
AND2X1   g2919(.A(WX5995), .B(RESET), .Y(n5188));
AND2X1   g2920(.A(WX5997), .B(RESET), .Y(n5193));
AND2X1   g2921(.A(WX5999), .B(RESET), .Y(n5198));
AND2X1   g2922(.A(WX6001), .B(RESET), .Y(n5203));
AND2X1   g2923(.A(WX6003), .B(RESET), .Y(n5208));
AND2X1   g2924(.A(WX6005), .B(RESET), .Y(n5213));
AND2X1   g2925(.A(WX6007), .B(RESET), .Y(n5218));
XOR2X1   g2926(.A(CRC_OUT_5_31), .B(WX6071), .Y(n8625_1));
NOR2X1   g2927(.A(n8625_1), .B(n5827), .Y(CRC_OUT_5_0));
XOR2X1   g2928(.A(CRC_OUT_5_0), .B(WX6069), .Y(n8627));
NOR2X1   g2929(.A(n8627), .B(n5827), .Y(CRC_OUT_5_1));
XOR2X1   g2930(.A(CRC_OUT_5_1), .B(WX6067), .Y(n8629));
NOR2X1   g2931(.A(n8629), .B(n5827), .Y(CRC_OUT_5_2));
XOR2X1   g2932(.A(CRC_OUT_5_2), .B(WX6065), .Y(n8631));
NOR2X1   g2933(.A(n8631), .B(n5827), .Y(CRC_OUT_5_3));
XOR2X1   g2934(.A(CRC_OUT_5_31), .B(WX6063), .Y(n8633));
XOR2X1   g2935(.A(n8633), .B(CRC_OUT_5_3), .Y(n8634));
NOR2X1   g2936(.A(n8634), .B(n5827), .Y(CRC_OUT_5_4));
XOR2X1   g2937(.A(CRC_OUT_5_4), .B(WX6061), .Y(n8636));
NOR2X1   g2938(.A(n8636), .B(n5827), .Y(CRC_OUT_5_5));
XOR2X1   g2939(.A(CRC_OUT_5_5), .B(WX6059), .Y(n8638));
NOR2X1   g2940(.A(n8638), .B(n5827), .Y(CRC_OUT_5_6));
XOR2X1   g2941(.A(CRC_OUT_5_6), .B(WX6057), .Y(n8640_1));
NOR2X1   g2942(.A(n8640_1), .B(n5827), .Y(CRC_OUT_5_7));
XOR2X1   g2943(.A(CRC_OUT_5_7), .B(WX6055), .Y(n8642));
NOR2X1   g2944(.A(n8642), .B(n5827), .Y(CRC_OUT_5_8));
XOR2X1   g2945(.A(CRC_OUT_5_8), .B(WX6053), .Y(n8644));
NOR2X1   g2946(.A(n8644), .B(n5827), .Y(CRC_OUT_5_9));
XOR2X1   g2947(.A(CRC_OUT_5_9), .B(WX6051), .Y(n8646));
NOR2X1   g2948(.A(n8646), .B(n5827), .Y(CRC_OUT_5_10));
XOR2X1   g2949(.A(CRC_OUT_5_31), .B(WX6049), .Y(n8648));
XOR2X1   g2950(.A(n8648), .B(CRC_OUT_5_10), .Y(n8649));
NOR2X1   g2951(.A(n8649), .B(n5827), .Y(CRC_OUT_5_11));
XOR2X1   g2952(.A(CRC_OUT_5_11), .B(WX6047), .Y(n8651));
NOR2X1   g2953(.A(n8651), .B(n5827), .Y(CRC_OUT_5_12));
XOR2X1   g2954(.A(CRC_OUT_5_12), .B(WX6045), .Y(n8653));
NOR2X1   g2955(.A(n8653), .B(n5827), .Y(CRC_OUT_5_13));
XOR2X1   g2956(.A(CRC_OUT_5_13), .B(WX6043), .Y(n8655_1));
NOR2X1   g2957(.A(n8655_1), .B(n5827), .Y(CRC_OUT_5_14));
XOR2X1   g2958(.A(CRC_OUT_5_14), .B(WX6041), .Y(n8657));
NOR2X1   g2959(.A(n8657), .B(n5827), .Y(CRC_OUT_5_15));
XOR2X1   g2960(.A(CRC_OUT_5_31), .B(WX6039), .Y(n8659));
XOR2X1   g2961(.A(n8659), .B(CRC_OUT_5_15), .Y(n8660_1));
NOR2X1   g2962(.A(n8660_1), .B(n5827), .Y(CRC_OUT_5_16));
XOR2X1   g2963(.A(CRC_OUT_5_16), .B(WX6037), .Y(n8662));
NOR2X1   g2964(.A(n8662), .B(n5827), .Y(CRC_OUT_5_17));
XOR2X1   g2965(.A(CRC_OUT_5_17), .B(WX6035), .Y(n8664));
NOR2X1   g2966(.A(n8664), .B(n5827), .Y(CRC_OUT_5_18));
XOR2X1   g2967(.A(CRC_OUT_5_18), .B(WX6033), .Y(n8666));
NOR2X1   g2968(.A(n8666), .B(n5827), .Y(CRC_OUT_5_19));
XOR2X1   g2969(.A(CRC_OUT_5_19), .B(WX6031), .Y(n8668));
NOR2X1   g2970(.A(n8668), .B(n5827), .Y(CRC_OUT_5_20));
XOR2X1   g2971(.A(CRC_OUT_5_20), .B(WX6029), .Y(n8670_1));
NOR2X1   g2972(.A(n8670_1), .B(n5827), .Y(CRC_OUT_5_21));
XOR2X1   g2973(.A(CRC_OUT_5_21), .B(WX6027), .Y(n8672));
NOR2X1   g2974(.A(n8672), .B(n5827), .Y(CRC_OUT_5_22));
XOR2X1   g2975(.A(CRC_OUT_5_22), .B(WX6025), .Y(n8674));
NOR2X1   g2976(.A(n8674), .B(n5827), .Y(CRC_OUT_5_23));
XOR2X1   g2977(.A(CRC_OUT_5_23), .B(WX6023), .Y(n8676));
NOR2X1   g2978(.A(n8676), .B(n5827), .Y(CRC_OUT_5_24));
XOR2X1   g2979(.A(CRC_OUT_5_24), .B(WX6021), .Y(n8678));
NOR2X1   g2980(.A(n8678), .B(n5827), .Y(CRC_OUT_5_25));
XOR2X1   g2981(.A(CRC_OUT_5_25), .B(WX6019), .Y(n8680_1));
NOR2X1   g2982(.A(n8680_1), .B(n5827), .Y(CRC_OUT_5_26));
XOR2X1   g2983(.A(CRC_OUT_5_26), .B(WX6017), .Y(n8682));
NOR2X1   g2984(.A(n8682), .B(n5827), .Y(CRC_OUT_5_27));
XOR2X1   g2985(.A(CRC_OUT_5_27), .B(WX6015), .Y(n8684));
NOR2X1   g2986(.A(n8684), .B(n5827), .Y(CRC_OUT_5_28));
XOR2X1   g2987(.A(CRC_OUT_5_28), .B(WX6013), .Y(n8686));
NOR2X1   g2988(.A(n8686), .B(n5827), .Y(CRC_OUT_5_29));
XOR2X1   g2989(.A(CRC_OUT_5_29), .B(WX6011), .Y(n8688));
NOR2X1   g2990(.A(n8688), .B(n5827), .Y(CRC_OUT_5_30));
XOR2X1   g2991(.A(CRC_OUT_5_30), .B(WX6009), .Y(n8690_1));
NOR2X1   g2992(.A(n8690_1), .B(n5827), .Y(CRC_OUT_5_31));
AND2X1   g2993(.A(WX6952), .B(RESET), .Y(n5351));
AND2X1   g2994(.A(WX6954), .B(RESET), .Y(n5356));
AND2X1   g2995(.A(WX6956), .B(RESET), .Y(n5361));
AND2X1   g2996(.A(WX6958), .B(RESET), .Y(n5366));
AND2X1   g2997(.A(WX6960), .B(RESET), .Y(n5371));
AND2X1   g2998(.A(WX6962), .B(RESET), .Y(n5376));
AND2X1   g2999(.A(WX6964), .B(RESET), .Y(n5381));
AND2X1   g3000(.A(WX6966), .B(RESET), .Y(n5386));
AND2X1   g3001(.A(WX6968), .B(RESET), .Y(n5391));
AND2X1   g3002(.A(WX6970), .B(RESET), .Y(n5396));
AND2X1   g3003(.A(WX6972), .B(RESET), .Y(n5401));
AND2X1   g3004(.A(WX6974), .B(RESET), .Y(n5406));
AND2X1   g3005(.A(WX6976), .B(RESET), .Y(n5411));
AND2X1   g3006(.A(WX6978), .B(RESET), .Y(n5416));
AND2X1   g3007(.A(WX6980), .B(RESET), .Y(n5421));
AND2X1   g3008(.A(WX6982), .B(RESET), .Y(n5426));
AND2X1   g3009(.A(WX6984), .B(RESET), .Y(n5431));
AND2X1   g3010(.A(WX6986), .B(RESET), .Y(n5436));
AND2X1   g3011(.A(WX6988), .B(RESET), .Y(n5441));
AND2X1   g3012(.A(WX6990), .B(RESET), .Y(n5446));
AND2X1   g3013(.A(WX6992), .B(RESET), .Y(n5451));
AND2X1   g3014(.A(WX6994), .B(RESET), .Y(n5456));
AND2X1   g3015(.A(WX6996), .B(RESET), .Y(n5461));
AND2X1   g3016(.A(WX6998), .B(RESET), .Y(n5466));
AND2X1   g3017(.A(WX7000), .B(RESET), .Y(n5471));
AND2X1   g3018(.A(WX7002), .B(RESET), .Y(n5476));
AND2X1   g3019(.A(WX7004), .B(RESET), .Y(n5481));
AND2X1   g3020(.A(WX7006), .B(RESET), .Y(n5486));
AND2X1   g3021(.A(WX7008), .B(RESET), .Y(n5491));
AND2X1   g3022(.A(WX7010), .B(RESET), .Y(n5496));
AND2X1   g3023(.A(WX7012), .B(RESET), .Y(n5501));
NOR2X1   g3024(.A(WX6950), .B(n5827), .Y(n5506));
INVX1    g3025(.A(CRC_OUT_4_31), .Y(n8724));
XOR2X1   g3026(.A(WX8403), .B(TM1), .Y(n8725_1));
XOR2X1   g3027(.A(n8725_1), .B(WX8467), .Y(n8726));
INVX1    g3028(.A(WX8531), .Y(n8727));
XOR2X1   g3029(.A(WX8595), .B(n8727), .Y(n8728));
XOR2X1   g3030(.A(n8728), .B(n8726), .Y(n8729));
MX2X1    g3031(.A(n8724), .B(n8729), .S0(n5539), .Y(n8731));
INVX1    g3032(.A(WX6950), .Y(n8732));
MX2X1    g3033(.A(n8732), .B(n8150_1), .S0(n5539), .Y(n8733));
MX2X1    g3034(.A(n8731), .B(n8733), .S0(TM1), .Y(n8734));
NOR2X1   g3035(.A(n8734), .B(n5827), .Y(n5511));
INVX1    g3036(.A(CRC_OUT_4_30), .Y(n8736));
XOR2X1   g3037(.A(WX8405), .B(TM1), .Y(n8737));
XOR2X1   g3038(.A(n8737), .B(WX8469), .Y(n8738));
INVX1    g3039(.A(WX8533), .Y(n8739));
XOR2X1   g3040(.A(WX8597), .B(n8739), .Y(n8740_1));
XOR2X1   g3041(.A(n8740_1), .B(n8738), .Y(n8741));
MX2X1    g3042(.A(n8736), .B(n8741), .S0(n5539), .Y(n8743));
INVX1    g3043(.A(WX6952), .Y(n8744));
MX2X1    g3044(.A(n8744), .B(n8162), .S0(n5539), .Y(n8745_1));
MX2X1    g3045(.A(n8743), .B(n8745_1), .S0(TM1), .Y(n8746));
NOR2X1   g3046(.A(n8746), .B(n5827), .Y(n5516));
INVX1    g3047(.A(CRC_OUT_4_29), .Y(n8748));
XOR2X1   g3048(.A(WX8407), .B(TM1), .Y(n8749));
XOR2X1   g3049(.A(n8749), .B(WX8471), .Y(n8750_1));
INVX1    g3050(.A(WX8535), .Y(n8751));
XOR2X1   g3051(.A(WX8599), .B(n8751), .Y(n8752));
XOR2X1   g3052(.A(n8752), .B(n8750_1), .Y(n8753));
MX2X1    g3053(.A(n8748), .B(n8753), .S0(n5539), .Y(n8755_1));
INVX1    g3054(.A(WX6954), .Y(n8756));
MX2X1    g3055(.A(n8756), .B(n8174), .S0(n5539), .Y(n8757));
MX2X1    g3056(.A(n8755_1), .B(n8757), .S0(TM1), .Y(n8758));
NOR2X1   g3057(.A(n8758), .B(n5827), .Y(n5521));
INVX1    g3058(.A(CRC_OUT_4_28), .Y(n8760_1));
XOR2X1   g3059(.A(WX8409), .B(TM1), .Y(n8761));
XOR2X1   g3060(.A(n8761), .B(WX8473), .Y(n8762));
INVX1    g3061(.A(WX8537), .Y(n8763));
XOR2X1   g3062(.A(WX8601), .B(n8763), .Y(n8764));
XOR2X1   g3063(.A(n8764), .B(n8762), .Y(n8765_1));
MX2X1    g3064(.A(n8760_1), .B(n8765_1), .S0(n5539), .Y(n8767));
INVX1    g3065(.A(WX6956), .Y(n8768));
MX2X1    g3066(.A(n8768), .B(n8186), .S0(n5539), .Y(n8769));
MX2X1    g3067(.A(n8767), .B(n8769), .S0(TM1), .Y(n8770_1));
NOR2X1   g3068(.A(n8770_1), .B(n5827), .Y(n5526));
INVX1    g3069(.A(CRC_OUT_4_27), .Y(n8772));
XOR2X1   g3070(.A(WX8411), .B(TM1), .Y(n8773));
XOR2X1   g3071(.A(n8773), .B(WX8475), .Y(n8774));
INVX1    g3072(.A(WX8539), .Y(n8775_1));
XOR2X1   g3073(.A(WX8603), .B(n8775_1), .Y(n8776));
XOR2X1   g3074(.A(n8776), .B(n8774), .Y(n8777));
MX2X1    g3075(.A(n8772), .B(n8777), .S0(n5539), .Y(n8779));
INVX1    g3076(.A(WX6958), .Y(n8780_1));
MX2X1    g3077(.A(n8780_1), .B(n8198), .S0(n5539), .Y(n8781));
MX2X1    g3078(.A(n8779), .B(n8781), .S0(TM1), .Y(n8782));
NOR2X1   g3079(.A(n8782), .B(n5827), .Y(n5531));
INVX1    g3080(.A(CRC_OUT_4_26), .Y(n8784));
XOR2X1   g3081(.A(WX8413), .B(TM1), .Y(n8785_1));
XOR2X1   g3082(.A(n8785_1), .B(WX8477), .Y(n8786));
INVX1    g3083(.A(WX8541), .Y(n8787));
XOR2X1   g3084(.A(WX8605), .B(n8787), .Y(n8788));
XOR2X1   g3085(.A(n8788), .B(n8786), .Y(n8789));
MX2X1    g3086(.A(n8784), .B(n8789), .S0(n5539), .Y(n8791));
INVX1    g3087(.A(WX6960), .Y(n8792));
MX2X1    g3088(.A(n8792), .B(n8210_1), .S0(n5539), .Y(n8793));
MX2X1    g3089(.A(n8791), .B(n8793), .S0(TM1), .Y(n8794));
NOR2X1   g3090(.A(n8794), .B(n5827), .Y(n5536));
INVX1    g3091(.A(CRC_OUT_4_25), .Y(n8796));
XOR2X1   g3092(.A(WX8415), .B(TM1), .Y(n8797));
XOR2X1   g3093(.A(n8797), .B(WX8479), .Y(n8798));
INVX1    g3094(.A(WX8543), .Y(n8799));
XOR2X1   g3095(.A(WX8607), .B(n8799), .Y(n8800_1));
XOR2X1   g3096(.A(n8800_1), .B(n8798), .Y(n8801));
MX2X1    g3097(.A(n8796), .B(n8801), .S0(n5539), .Y(n8803));
INVX1    g3098(.A(WX6962), .Y(n8804));
MX2X1    g3099(.A(n8804), .B(n8222), .S0(n5539), .Y(n8805_1));
MX2X1    g3100(.A(n8803), .B(n8805_1), .S0(TM1), .Y(n8806));
NOR2X1   g3101(.A(n8806), .B(n5827), .Y(n5541));
INVX1    g3102(.A(CRC_OUT_4_24), .Y(n8808));
XOR2X1   g3103(.A(WX8417), .B(TM1), .Y(n8809));
XOR2X1   g3104(.A(n8809), .B(WX8481), .Y(n8810_1));
INVX1    g3105(.A(WX8545), .Y(n8811));
XOR2X1   g3106(.A(WX8609), .B(n8811), .Y(n8812));
XOR2X1   g3107(.A(n8812), .B(n8810_1), .Y(n8813));
MX2X1    g3108(.A(n8808), .B(n8813), .S0(n5539), .Y(n8815_1));
INVX1    g3109(.A(WX6964), .Y(n8816));
MX2X1    g3110(.A(n8816), .B(n8234), .S0(n5539), .Y(n8817));
MX2X1    g3111(.A(n8815_1), .B(n8817), .S0(TM1), .Y(n8818));
NOR2X1   g3112(.A(n8818), .B(n5827), .Y(n5546));
INVX1    g3113(.A(CRC_OUT_4_23), .Y(n8820_1));
XOR2X1   g3114(.A(WX8419), .B(TM1), .Y(n8821));
XOR2X1   g3115(.A(n8821), .B(WX8483), .Y(n8822));
INVX1    g3116(.A(WX8547), .Y(n8823));
XOR2X1   g3117(.A(WX8611), .B(n8823), .Y(n8824));
XOR2X1   g3118(.A(n8824), .B(n8822), .Y(n8825_1));
MX2X1    g3119(.A(n8820_1), .B(n8825_1), .S0(n5539), .Y(n8827));
INVX1    g3120(.A(WX6966), .Y(n8828));
MX2X1    g3121(.A(n8828), .B(n8246), .S0(n5539), .Y(n8829));
MX2X1    g3122(.A(n8827), .B(n8829), .S0(TM1), .Y(n8830_1));
NOR2X1   g3123(.A(n8830_1), .B(n5827), .Y(n5551));
INVX1    g3124(.A(CRC_OUT_4_22), .Y(n8832));
XOR2X1   g3125(.A(WX8421), .B(TM1), .Y(n8833));
XOR2X1   g3126(.A(n8833), .B(WX8485), .Y(n8834));
INVX1    g3127(.A(WX8549), .Y(n8835_1));
XOR2X1   g3128(.A(WX8613), .B(n8835_1), .Y(n8836));
XOR2X1   g3129(.A(n8836), .B(n8834), .Y(n8837));
MX2X1    g3130(.A(n8832), .B(n8837), .S0(n5539), .Y(n8839));
INVX1    g3131(.A(WX6968), .Y(n8840_1));
MX2X1    g3132(.A(n8840_1), .B(n8258), .S0(n5539), .Y(n8841));
MX2X1    g3133(.A(n8839), .B(n8841), .S0(TM1), .Y(n8842));
NOR2X1   g3134(.A(n8842), .B(n5827), .Y(n5556));
INVX1    g3135(.A(CRC_OUT_4_21), .Y(n8844));
XOR2X1   g3136(.A(WX8423), .B(TM1), .Y(n8845_1));
XOR2X1   g3137(.A(n8845_1), .B(WX8487), .Y(n8846));
INVX1    g3138(.A(WX8551), .Y(n8847));
XOR2X1   g3139(.A(WX8615), .B(n8847), .Y(n8848));
XOR2X1   g3140(.A(n8848), .B(n8846), .Y(n8849));
MX2X1    g3141(.A(n8844), .B(n8849), .S0(n5539), .Y(n8851));
INVX1    g3142(.A(WX6970), .Y(n8852));
MX2X1    g3143(.A(n8852), .B(n8270_1), .S0(n5539), .Y(n8853));
MX2X1    g3144(.A(n8851), .B(n8853), .S0(TM1), .Y(n8854));
NOR2X1   g3145(.A(n8854), .B(n5827), .Y(n5561));
INVX1    g3146(.A(CRC_OUT_4_20), .Y(n8856));
XOR2X1   g3147(.A(WX8425), .B(TM1), .Y(n8857));
XOR2X1   g3148(.A(n8857), .B(WX8489), .Y(n8858));
INVX1    g3149(.A(WX8553), .Y(n8859));
XOR2X1   g3150(.A(WX8617), .B(n8859), .Y(n8860_1));
XOR2X1   g3151(.A(n8860_1), .B(n8858), .Y(n8861));
MX2X1    g3152(.A(n8856), .B(n8861), .S0(n5539), .Y(n8863));
INVX1    g3153(.A(WX6972), .Y(n8864));
MX2X1    g3154(.A(n8864), .B(n8282), .S0(n5539), .Y(n8865_1));
MX2X1    g3155(.A(n8863), .B(n8865_1), .S0(TM1), .Y(n8866));
NOR2X1   g3156(.A(n8866), .B(n5827), .Y(n5566));
INVX1    g3157(.A(CRC_OUT_4_19), .Y(n8868));
XOR2X1   g3158(.A(WX8427), .B(TM1), .Y(n8869));
XOR2X1   g3159(.A(n8869), .B(WX8491), .Y(n8870_1));
INVX1    g3160(.A(WX8555), .Y(n8871));
XOR2X1   g3161(.A(WX8619), .B(n8871), .Y(n8872));
XOR2X1   g3162(.A(n8872), .B(n8870_1), .Y(n8873));
MX2X1    g3163(.A(n8868), .B(n8873), .S0(n5539), .Y(n8875_1));
INVX1    g3164(.A(WX6974), .Y(n8876));
MX2X1    g3165(.A(n8876), .B(n8294), .S0(n5539), .Y(n8877));
MX2X1    g3166(.A(n8875_1), .B(n8877), .S0(TM1), .Y(n8878));
NOR2X1   g3167(.A(n8878), .B(n5827), .Y(n5571));
INVX1    g3168(.A(CRC_OUT_4_18), .Y(n8880_1));
XOR2X1   g3169(.A(WX8429), .B(TM1), .Y(n8881));
XOR2X1   g3170(.A(n8881), .B(WX8493), .Y(n8882));
INVX1    g3171(.A(WX8557), .Y(n8883));
XOR2X1   g3172(.A(WX8621), .B(n8883), .Y(n8884));
XOR2X1   g3173(.A(n8884), .B(n8882), .Y(n8885_1));
MX2X1    g3174(.A(n8880_1), .B(n8885_1), .S0(n5539), .Y(n8887));
INVX1    g3175(.A(WX6976), .Y(n8888));
MX2X1    g3176(.A(n8888), .B(n8306), .S0(n5539), .Y(n8889));
MX2X1    g3177(.A(n8887), .B(n8889), .S0(TM1), .Y(n8890_1));
NOR2X1   g3178(.A(n8890_1), .B(n5827), .Y(n5576));
INVX1    g3179(.A(CRC_OUT_4_17), .Y(n8892));
XOR2X1   g3180(.A(WX8431), .B(TM1), .Y(n8893));
XOR2X1   g3181(.A(n8893), .B(WX8495), .Y(n8894));
INVX1    g3182(.A(WX8559), .Y(n8895_1));
XOR2X1   g3183(.A(WX8623), .B(n8895_1), .Y(n8896));
XOR2X1   g3184(.A(n8896), .B(n8894), .Y(n8897));
MX2X1    g3185(.A(n8892), .B(n8897), .S0(n5539), .Y(n8899));
INVX1    g3186(.A(WX6978), .Y(n8900_1));
MX2X1    g3187(.A(n8900_1), .B(n8318), .S0(n5539), .Y(n8901));
MX2X1    g3188(.A(n8899), .B(n8901), .S0(TM1), .Y(n8902));
NOR2X1   g3189(.A(n8902), .B(n5827), .Y(n5581));
INVX1    g3190(.A(CRC_OUT_4_16), .Y(n8904));
XOR2X1   g3191(.A(WX8433), .B(TM1), .Y(n8905_1));
XOR2X1   g3192(.A(n8905_1), .B(WX8497), .Y(n8906));
INVX1    g3193(.A(WX8561), .Y(n8907));
XOR2X1   g3194(.A(WX8625), .B(n8907), .Y(n8908));
XOR2X1   g3195(.A(n8908), .B(n8906), .Y(n8909));
MX2X1    g3196(.A(n8904), .B(n8909), .S0(n5539), .Y(n8911));
INVX1    g3197(.A(WX6980), .Y(n8912));
MX2X1    g3198(.A(n8912), .B(n8330_1), .S0(n5539), .Y(n8913));
MX2X1    g3199(.A(n8911), .B(n8913), .S0(TM1), .Y(n8914));
NOR2X1   g3200(.A(n8914), .B(n5827), .Y(n5586));
INVX1    g3201(.A(CRC_OUT_4_15), .Y(n8916));
XOR2X1   g3202(.A(WX8435), .B(TM0), .Y(n8917));
XOR2X1   g3203(.A(n8917), .B(WX8499), .Y(n8918));
INVX1    g3204(.A(WX8563), .Y(n8919));
XOR2X1   g3205(.A(WX8627), .B(n8919), .Y(n8920_1));
XOR2X1   g3206(.A(n8920_1), .B(n8918), .Y(n8921));
MX2X1    g3207(.A(n8916), .B(n8921), .S0(n5539), .Y(n8923));
INVX1    g3208(.A(WX6982), .Y(n8924));
MX2X1    g3209(.A(n8924), .B(n8342), .S0(n5539), .Y(n8925_1));
MX2X1    g3210(.A(n8923), .B(n8925_1), .S0(TM1), .Y(n8926));
NOR2X1   g3211(.A(n8926), .B(n5827), .Y(n5591));
INVX1    g3212(.A(CRC_OUT_4_14), .Y(n8928));
XOR2X1   g3213(.A(WX8437), .B(TM0), .Y(n8929));
XOR2X1   g3214(.A(n8929), .B(WX8501), .Y(n8930_1));
INVX1    g3215(.A(WX8565), .Y(n8931));
XOR2X1   g3216(.A(WX8629), .B(n8931), .Y(n8932));
XOR2X1   g3217(.A(n8932), .B(n8930_1), .Y(n8933));
MX2X1    g3218(.A(n8928), .B(n8933), .S0(n5539), .Y(n8935_1));
INVX1    g3219(.A(WX6984), .Y(n8936));
MX2X1    g3220(.A(n8936), .B(n8354), .S0(n5539), .Y(n8937));
MX2X1    g3221(.A(n8935_1), .B(n8937), .S0(TM1), .Y(n8938));
NOR2X1   g3222(.A(n8938), .B(n5827), .Y(n5596));
INVX1    g3223(.A(CRC_OUT_4_13), .Y(n8940));
XOR2X1   g3224(.A(WX8439), .B(TM0), .Y(n8941));
XOR2X1   g3225(.A(n8941), .B(WX8503), .Y(n8942));
INVX1    g3226(.A(WX8567), .Y(n8943_1));
XOR2X1   g3227(.A(WX8631), .B(n8943_1), .Y(n8944));
XOR2X1   g3228(.A(n8944), .B(n8942), .Y(n8945));
MX2X1    g3229(.A(n8940), .B(n8945), .S0(n5539), .Y(n8947_1));
INVX1    g3230(.A(WX6986), .Y(n8948));
MX2X1    g3231(.A(n8948), .B(n8366), .S0(n5539), .Y(n8949));
MX2X1    g3232(.A(n8947_1), .B(n8949), .S0(TM1), .Y(n8950));
NOR2X1   g3233(.A(n8950), .B(n5827), .Y(n5601));
INVX1    g3234(.A(CRC_OUT_4_12), .Y(n8952));
XOR2X1   g3235(.A(WX8441), .B(TM0), .Y(n8953));
XOR2X1   g3236(.A(n8953), .B(WX8505), .Y(n8954));
INVX1    g3237(.A(WX8569), .Y(n8955_1));
XOR2X1   g3238(.A(WX8633), .B(n8955_1), .Y(n8956));
XOR2X1   g3239(.A(n8956), .B(n8954), .Y(n8957));
MX2X1    g3240(.A(n8952), .B(n8957), .S0(n5539), .Y(n8959_1));
INVX1    g3241(.A(WX6988), .Y(n8960));
MX2X1    g3242(.A(n8960), .B(n8378), .S0(n5539), .Y(n8961));
MX2X1    g3243(.A(n8959_1), .B(n8961), .S0(TM1), .Y(n8962));
NOR2X1   g3244(.A(n8962), .B(n5827), .Y(n5606));
INVX1    g3245(.A(CRC_OUT_4_11), .Y(n8964));
XOR2X1   g3246(.A(WX8443), .B(TM0), .Y(n8965));
XOR2X1   g3247(.A(n8965), .B(WX8507), .Y(n8966));
INVX1    g3248(.A(WX8571), .Y(n8967_1));
XOR2X1   g3249(.A(WX8635), .B(n8967_1), .Y(n8968));
XOR2X1   g3250(.A(n8968), .B(n8966), .Y(n8969));
MX2X1    g3251(.A(n8964), .B(n8969), .S0(n5539), .Y(n8971_1));
INVX1    g3252(.A(WX6990), .Y(n8972));
MX2X1    g3253(.A(n8972), .B(n8390_1), .S0(n5539), .Y(n8973));
MX2X1    g3254(.A(n8971_1), .B(n8973), .S0(TM1), .Y(n8974));
NOR2X1   g3255(.A(n8974), .B(n5827), .Y(n5611));
INVX1    g3256(.A(CRC_OUT_4_10), .Y(n8976));
XOR2X1   g3257(.A(WX8445), .B(TM0), .Y(n8977));
XOR2X1   g3258(.A(n8977), .B(WX8509), .Y(n8978));
INVX1    g3259(.A(WX8573), .Y(n8979_1));
XOR2X1   g3260(.A(WX8637), .B(n8979_1), .Y(n8980));
XOR2X1   g3261(.A(n8980), .B(n8978), .Y(n8981));
MX2X1    g3262(.A(n8976), .B(n8981), .S0(n5539), .Y(n8983_1));
INVX1    g3263(.A(WX6992), .Y(n8984));
MX2X1    g3264(.A(n8984), .B(n8402), .S0(n5539), .Y(n8985));
MX2X1    g3265(.A(n8983_1), .B(n8985), .S0(TM1), .Y(n8986));
NOR2X1   g3266(.A(n8986), .B(n5827), .Y(n5616));
INVX1    g3267(.A(CRC_OUT_4_9), .Y(n8988));
XOR2X1   g3268(.A(WX8447), .B(TM0), .Y(n8989));
XOR2X1   g3269(.A(n8989), .B(WX8511), .Y(n8990));
INVX1    g3270(.A(WX8575), .Y(n8991_1));
XOR2X1   g3271(.A(WX8639), .B(n8991_1), .Y(n8992));
XOR2X1   g3272(.A(n8992), .B(n8990), .Y(n8993));
MX2X1    g3273(.A(n8988), .B(n8993), .S0(n5539), .Y(n8995_1));
INVX1    g3274(.A(WX6994), .Y(n8996));
MX2X1    g3275(.A(n8996), .B(n8414), .S0(n5539), .Y(n8997));
MX2X1    g3276(.A(n8995_1), .B(n8997), .S0(TM1), .Y(n8998));
NOR2X1   g3277(.A(n8998), .B(n5827), .Y(n5621));
INVX1    g3278(.A(CRC_OUT_4_8), .Y(n9000));
XOR2X1   g3279(.A(WX8449), .B(TM0), .Y(n9001));
XOR2X1   g3280(.A(n9001), .B(WX8513), .Y(n9002));
INVX1    g3281(.A(WX8577), .Y(n9003_1));
XOR2X1   g3282(.A(WX8641), .B(n9003_1), .Y(n9004));
XOR2X1   g3283(.A(n9004), .B(n9002), .Y(n9005));
MX2X1    g3284(.A(n9000), .B(n9005), .S0(n5539), .Y(n9007_1));
INVX1    g3285(.A(WX6996), .Y(n9008));
MX2X1    g3286(.A(n9008), .B(n8426), .S0(n5539), .Y(n9009));
MX2X1    g3287(.A(n9007_1), .B(n9009), .S0(TM1), .Y(n9010));
NOR2X1   g3288(.A(n9010), .B(n5827), .Y(n5626));
INVX1    g3289(.A(CRC_OUT_4_7), .Y(n9012));
XOR2X1   g3290(.A(WX8451), .B(TM0), .Y(n9013));
XOR2X1   g3291(.A(n9013), .B(WX8515), .Y(n9014));
INVX1    g3292(.A(WX8579), .Y(n9015_1));
XOR2X1   g3293(.A(WX8643), .B(n9015_1), .Y(n9016));
XOR2X1   g3294(.A(n9016), .B(n9014), .Y(n9017));
MX2X1    g3295(.A(n9012), .B(n9017), .S0(n5539), .Y(n9019_1));
INVX1    g3296(.A(WX6998), .Y(n9020));
MX2X1    g3297(.A(n9020), .B(n8438), .S0(n5539), .Y(n9021));
MX2X1    g3298(.A(n9019_1), .B(n9021), .S0(TM1), .Y(n9022));
NOR2X1   g3299(.A(n9022), .B(n5827), .Y(n5631));
INVX1    g3300(.A(CRC_OUT_4_6), .Y(n9024));
XOR2X1   g3301(.A(WX8453), .B(TM0), .Y(n9025));
XOR2X1   g3302(.A(n9025), .B(WX8517), .Y(n9026));
INVX1    g3303(.A(WX8581), .Y(n9027_1));
XOR2X1   g3304(.A(WX8645), .B(n9027_1), .Y(n9028));
XOR2X1   g3305(.A(n9028), .B(n9026), .Y(n9029));
MX2X1    g3306(.A(n9024), .B(n9029), .S0(n5539), .Y(n9031_1));
INVX1    g3307(.A(WX7000), .Y(n9032));
MX2X1    g3308(.A(n9032), .B(n8450_1), .S0(n5539), .Y(n9033));
MX2X1    g3309(.A(n9031_1), .B(n9033), .S0(TM1), .Y(n9034));
NOR2X1   g3310(.A(n9034), .B(n5827), .Y(n5636));
INVX1    g3311(.A(CRC_OUT_4_5), .Y(n9036));
XOR2X1   g3312(.A(WX8455), .B(TM0), .Y(n9037));
XOR2X1   g3313(.A(n9037), .B(WX8519), .Y(n9038));
INVX1    g3314(.A(WX8583), .Y(n9039_1));
XOR2X1   g3315(.A(WX8647), .B(n9039_1), .Y(n9040));
XOR2X1   g3316(.A(n9040), .B(n9038), .Y(n9041));
MX2X1    g3317(.A(n9036), .B(n9041), .S0(n5539), .Y(n9043_1));
INVX1    g3318(.A(WX7002), .Y(n9044));
MX2X1    g3319(.A(n9044), .B(n8462), .S0(n5539), .Y(n9045));
MX2X1    g3320(.A(n9043_1), .B(n9045), .S0(TM1), .Y(n9046));
NOR2X1   g3321(.A(n9046), .B(n5827), .Y(n5641));
INVX1    g3322(.A(CRC_OUT_4_4), .Y(n9048));
XOR2X1   g3323(.A(WX8457), .B(TM0), .Y(n9049));
XOR2X1   g3324(.A(n9049), .B(WX8521), .Y(n9050));
INVX1    g3325(.A(WX8585), .Y(n9051_1));
XOR2X1   g3326(.A(WX8649), .B(n9051_1), .Y(n9052));
XOR2X1   g3327(.A(n9052), .B(n9050), .Y(n9053));
MX2X1    g3328(.A(n9048), .B(n9053), .S0(n5539), .Y(n9055_1));
INVX1    g3329(.A(WX7004), .Y(n9056));
MX2X1    g3330(.A(n9056), .B(n8474), .S0(n5539), .Y(n9057));
MX2X1    g3331(.A(n9055_1), .B(n9057), .S0(TM1), .Y(n9058));
NOR2X1   g3332(.A(n9058), .B(n5827), .Y(n5646));
INVX1    g3333(.A(CRC_OUT_4_3), .Y(n9060));
XOR2X1   g3334(.A(WX8459), .B(TM0), .Y(n9061));
XOR2X1   g3335(.A(n9061), .B(WX8523), .Y(n9062));
INVX1    g3336(.A(WX8587), .Y(n9063));
XOR2X1   g3337(.A(WX8651), .B(n9063), .Y(n9064));
XOR2X1   g3338(.A(n9064), .B(n9062), .Y(n9065));
MX2X1    g3339(.A(n9060), .B(n9065), .S0(n5539), .Y(n9067));
INVX1    g3340(.A(WX7006), .Y(n9068));
MX2X1    g3341(.A(n9068), .B(n8486), .S0(n5539), .Y(n9069));
MX2X1    g3342(.A(n9067), .B(n9069), .S0(TM1), .Y(n9070));
NOR2X1   g3343(.A(n9070), .B(n5827), .Y(n5651));
INVX1    g3344(.A(CRC_OUT_4_2), .Y(n9072));
XOR2X1   g3345(.A(WX8461), .B(TM0), .Y(n9073));
XOR2X1   g3346(.A(n9073), .B(WX8525), .Y(n9074));
INVX1    g3347(.A(WX8589), .Y(n9075));
XOR2X1   g3348(.A(WX8653), .B(n9075), .Y(n9076));
XOR2X1   g3349(.A(n9076), .B(n9074), .Y(n9077));
MX2X1    g3350(.A(n9072), .B(n9077), .S0(n5539), .Y(n9079));
INVX1    g3351(.A(WX7008), .Y(n9080));
MX2X1    g3352(.A(n9080), .B(n8498), .S0(n5539), .Y(n9081));
MX2X1    g3353(.A(n9079), .B(n9081), .S0(TM1), .Y(n9082));
NOR2X1   g3354(.A(n9082), .B(n5827), .Y(n5656));
INVX1    g3355(.A(CRC_OUT_4_1), .Y(n9084));
XOR2X1   g3356(.A(WX8463), .B(TM0), .Y(n9085));
XOR2X1   g3357(.A(n9085), .B(WX8527), .Y(n9086));
INVX1    g3358(.A(WX8591), .Y(n9087));
XOR2X1   g3359(.A(WX8655), .B(n9087), .Y(n9088));
XOR2X1   g3360(.A(n9088), .B(n9086), .Y(n9089));
MX2X1    g3361(.A(n9084), .B(n9089), .S0(n5539), .Y(n9091));
INVX1    g3362(.A(WX7010), .Y(n9092));
MX2X1    g3363(.A(n9092), .B(n8510_1), .S0(n5539), .Y(n9093));
MX2X1    g3364(.A(n9091), .B(n9093), .S0(TM1), .Y(n9094));
NOR2X1   g3365(.A(n9094), .B(n5827), .Y(n5661));
INVX1    g3366(.A(CRC_OUT_4_0), .Y(n9096));
XOR2X1   g3367(.A(WX8465), .B(TM0), .Y(n9097));
XOR2X1   g3368(.A(n9097), .B(WX8529), .Y(n9098));
INVX1    g3369(.A(WX8593), .Y(n9099));
XOR2X1   g3370(.A(WX8657), .B(n9099), .Y(n9100));
XOR2X1   g3371(.A(n9100), .B(n9098), .Y(n9101));
MX2X1    g3372(.A(n9096), .B(n9101), .S0(n5539), .Y(n9103));
INVX1    g3373(.A(WX7012), .Y(n9104));
MX2X1    g3374(.A(n9104), .B(n8522), .S0(n5539), .Y(n9105));
MX2X1    g3375(.A(n9103), .B(n9105), .S0(TM1), .Y(n9106));
NOR2X1   g3376(.A(n9106), .B(n5827), .Y(n5666));
AND2X1   g3377(.A(WX7110), .B(RESET), .Y(n5671));
AND2X1   g3378(.A(WX7112), .B(RESET), .Y(n5676));
AND2X1   g3379(.A(WX7114), .B(RESET), .Y(n5681));
AND2X1   g3380(.A(WX7116), .B(RESET), .Y(n5686));
AND2X1   g3381(.A(WX7118), .B(RESET), .Y(n5691));
AND2X1   g3382(.A(WX7120), .B(RESET), .Y(n5696));
AND2X1   g3383(.A(WX7122), .B(RESET), .Y(n5701));
AND2X1   g3384(.A(WX7124), .B(RESET), .Y(n5706));
AND2X1   g3385(.A(WX7126), .B(RESET), .Y(n5711));
AND2X1   g3386(.A(WX7128), .B(RESET), .Y(n5716));
AND2X1   g3387(.A(WX7130), .B(RESET), .Y(n5721));
AND2X1   g3388(.A(WX7132), .B(RESET), .Y(n5726));
AND2X1   g3389(.A(WX7134), .B(RESET), .Y(n5731));
AND2X1   g3390(.A(WX7136), .B(RESET), .Y(n5736));
AND2X1   g3391(.A(WX7138), .B(RESET), .Y(n5741));
AND2X1   g3392(.A(WX7140), .B(RESET), .Y(n5746));
AND2X1   g3393(.A(WX7142), .B(RESET), .Y(n5751));
AND2X1   g3394(.A(WX7144), .B(RESET), .Y(n5756));
AND2X1   g3395(.A(WX7146), .B(RESET), .Y(n5761));
AND2X1   g3396(.A(WX7148), .B(RESET), .Y(n5766));
AND2X1   g3397(.A(WX7150), .B(RESET), .Y(n5771));
AND2X1   g3398(.A(WX7152), .B(RESET), .Y(n5776));
AND2X1   g3399(.A(WX7154), .B(RESET), .Y(n5781));
AND2X1   g3400(.A(WX7156), .B(RESET), .Y(n5786));
AND2X1   g3401(.A(WX7158), .B(RESET), .Y(n5791));
AND2X1   g3402(.A(WX7160), .B(RESET), .Y(n5796));
AND2X1   g3403(.A(WX7162), .B(RESET), .Y(n5801));
AND2X1   g3404(.A(WX7164), .B(RESET), .Y(n5806));
AND2X1   g3405(.A(WX7166), .B(RESET), .Y(n5811));
AND2X1   g3406(.A(WX7168), .B(RESET), .Y(n5816));
AND2X1   g3407(.A(WX7170), .B(RESET), .Y(n5821));
AND2X1   g3408(.A(WX7172), .B(RESET), .Y(n5826));
AND2X1   g3409(.A(WX7174), .B(RESET), .Y(n5831));
AND2X1   g3410(.A(WX7176), .B(RESET), .Y(n5836));
AND2X1   g3411(.A(WX7178), .B(RESET), .Y(n5841));
AND2X1   g3412(.A(WX7180), .B(RESET), .Y(n5846));
AND2X1   g3413(.A(WX7182), .B(RESET), .Y(n5851));
AND2X1   g3414(.A(WX7184), .B(RESET), .Y(n5856));
AND2X1   g3415(.A(WX7186), .B(RESET), .Y(n5861));
AND2X1   g3416(.A(WX7188), .B(RESET), .Y(n5866));
AND2X1   g3417(.A(WX7190), .B(RESET), .Y(n5871));
AND2X1   g3418(.A(WX7192), .B(RESET), .Y(n5876));
AND2X1   g3419(.A(WX7194), .B(RESET), .Y(n5881));
AND2X1   g3420(.A(WX7196), .B(RESET), .Y(n5886));
AND2X1   g3421(.A(WX7198), .B(RESET), .Y(n5891));
AND2X1   g3422(.A(WX7200), .B(RESET), .Y(n5896));
AND2X1   g3423(.A(WX7202), .B(RESET), .Y(n5901));
AND2X1   g3424(.A(WX7204), .B(RESET), .Y(n5906));
AND2X1   g3425(.A(WX7206), .B(RESET), .Y(n5911));
AND2X1   g3426(.A(WX7208), .B(RESET), .Y(n5916));
AND2X1   g3427(.A(WX7210), .B(RESET), .Y(n5921));
AND2X1   g3428(.A(WX7212), .B(RESET), .Y(n5926));
AND2X1   g3429(.A(WX7214), .B(RESET), .Y(n5931));
AND2X1   g3430(.A(WX7216), .B(RESET), .Y(n5936));
AND2X1   g3431(.A(WX7218), .B(RESET), .Y(n5941));
AND2X1   g3432(.A(WX7220), .B(RESET), .Y(n5946));
AND2X1   g3433(.A(WX7222), .B(RESET), .Y(n5951));
AND2X1   g3434(.A(WX7224), .B(RESET), .Y(n5956));
AND2X1   g3435(.A(WX7226), .B(RESET), .Y(n5961));
AND2X1   g3436(.A(WX7228), .B(RESET), .Y(n5966));
AND2X1   g3437(.A(WX7230), .B(RESET), .Y(n5971));
AND2X1   g3438(.A(WX7232), .B(RESET), .Y(n5976));
AND2X1   g3439(.A(WX7234), .B(RESET), .Y(n5981));
AND2X1   g3440(.A(WX7236), .B(RESET), .Y(n5986));
AND2X1   g3441(.A(WX7238), .B(RESET), .Y(n5991));
AND2X1   g3442(.A(WX7240), .B(RESET), .Y(n5996));
AND2X1   g3443(.A(WX7242), .B(RESET), .Y(n6001));
AND2X1   g3444(.A(WX7244), .B(RESET), .Y(n6006));
AND2X1   g3445(.A(WX7246), .B(RESET), .Y(n6011));
AND2X1   g3446(.A(WX7248), .B(RESET), .Y(n6016));
AND2X1   g3447(.A(WX7250), .B(RESET), .Y(n6021));
AND2X1   g3448(.A(WX7252), .B(RESET), .Y(n6026));
AND2X1   g3449(.A(WX7254), .B(RESET), .Y(n6031));
AND2X1   g3450(.A(WX7256), .B(RESET), .Y(n6036));
AND2X1   g3451(.A(WX7258), .B(RESET), .Y(n6041));
AND2X1   g3452(.A(WX7260), .B(RESET), .Y(n6046));
AND2X1   g3453(.A(WX7262), .B(RESET), .Y(n6051));
AND2X1   g3454(.A(WX7264), .B(RESET), .Y(n6056));
AND2X1   g3455(.A(WX7266), .B(RESET), .Y(n6061));
AND2X1   g3456(.A(WX7268), .B(RESET), .Y(n6066));
AND2X1   g3457(.A(WX7270), .B(RESET), .Y(n6071));
AND2X1   g3458(.A(WX7272), .B(RESET), .Y(n6076));
AND2X1   g3459(.A(WX7274), .B(RESET), .Y(n6081));
AND2X1   g3460(.A(WX7276), .B(RESET), .Y(n6086));
AND2X1   g3461(.A(WX7278), .B(RESET), .Y(n6091));
AND2X1   g3462(.A(WX7280), .B(RESET), .Y(n6096));
AND2X1   g3463(.A(WX7282), .B(RESET), .Y(n6101));
AND2X1   g3464(.A(WX7284), .B(RESET), .Y(n6106));
AND2X1   g3465(.A(WX7286), .B(RESET), .Y(n6111));
AND2X1   g3466(.A(WX7288), .B(RESET), .Y(n6116));
AND2X1   g3467(.A(WX7290), .B(RESET), .Y(n6121));
AND2X1   g3468(.A(WX7292), .B(RESET), .Y(n6126));
AND2X1   g3469(.A(WX7294), .B(RESET), .Y(n6131));
AND2X1   g3470(.A(WX7296), .B(RESET), .Y(n6136));
AND2X1   g3471(.A(WX7298), .B(RESET), .Y(n6141));
AND2X1   g3472(.A(WX7300), .B(RESET), .Y(n6146));
XOR2X1   g3473(.A(CRC_OUT_4_31), .B(WX7364), .Y(n9204));
NOR2X1   g3474(.A(n9204), .B(n5827), .Y(CRC_OUT_4_0));
XOR2X1   g3475(.A(CRC_OUT_4_0), .B(WX7362), .Y(n9206));
NOR2X1   g3476(.A(n9206), .B(n5827), .Y(CRC_OUT_4_1));
XOR2X1   g3477(.A(CRC_OUT_4_1), .B(WX7360), .Y(n9208));
NOR2X1   g3478(.A(n9208), .B(n5827), .Y(CRC_OUT_4_2));
XOR2X1   g3479(.A(CRC_OUT_4_2), .B(WX7358), .Y(n9210));
NOR2X1   g3480(.A(n9210), .B(n5827), .Y(CRC_OUT_4_3));
XOR2X1   g3481(.A(CRC_OUT_4_31), .B(WX7356), .Y(n9212));
XOR2X1   g3482(.A(n9212), .B(CRC_OUT_4_3), .Y(n9213));
NOR2X1   g3483(.A(n9213), .B(n5827), .Y(CRC_OUT_4_4));
XOR2X1   g3484(.A(CRC_OUT_4_4), .B(WX7354), .Y(n9215));
NOR2X1   g3485(.A(n9215), .B(n5827), .Y(CRC_OUT_4_5));
XOR2X1   g3486(.A(CRC_OUT_4_5), .B(WX7352), .Y(n9217));
NOR2X1   g3487(.A(n9217), .B(n5827), .Y(CRC_OUT_4_6));
XOR2X1   g3488(.A(CRC_OUT_4_6), .B(WX7350), .Y(n9219));
NOR2X1   g3489(.A(n9219), .B(n5827), .Y(CRC_OUT_4_7));
XOR2X1   g3490(.A(CRC_OUT_4_7), .B(WX7348), .Y(n9221));
NOR2X1   g3491(.A(n9221), .B(n5827), .Y(CRC_OUT_4_8));
XOR2X1   g3492(.A(CRC_OUT_4_8), .B(WX7346), .Y(n9223));
NOR2X1   g3493(.A(n9223), .B(n5827), .Y(CRC_OUT_4_9));
XOR2X1   g3494(.A(CRC_OUT_4_9), .B(WX7344), .Y(n9225));
NOR2X1   g3495(.A(n9225), .B(n5827), .Y(CRC_OUT_4_10));
XOR2X1   g3496(.A(CRC_OUT_4_31), .B(WX7342), .Y(n9227));
XOR2X1   g3497(.A(n9227), .B(CRC_OUT_4_10), .Y(n9228));
NOR2X1   g3498(.A(n9228), .B(n5827), .Y(CRC_OUT_4_11));
XOR2X1   g3499(.A(CRC_OUT_4_11), .B(WX7340), .Y(n9230));
NOR2X1   g3500(.A(n9230), .B(n5827), .Y(CRC_OUT_4_12));
XOR2X1   g3501(.A(CRC_OUT_4_12), .B(WX7338), .Y(n9232));
NOR2X1   g3502(.A(n9232), .B(n5827), .Y(CRC_OUT_4_13));
XOR2X1   g3503(.A(CRC_OUT_4_13), .B(WX7336), .Y(n9234));
NOR2X1   g3504(.A(n9234), .B(n5827), .Y(CRC_OUT_4_14));
XOR2X1   g3505(.A(CRC_OUT_4_14), .B(WX7334), .Y(n9236));
NOR2X1   g3506(.A(n9236), .B(n5827), .Y(CRC_OUT_4_15));
XOR2X1   g3507(.A(CRC_OUT_4_31), .B(WX7332), .Y(n9238));
XOR2X1   g3508(.A(n9238), .B(CRC_OUT_4_15), .Y(n9239));
NOR2X1   g3509(.A(n9239), .B(n5827), .Y(CRC_OUT_4_16));
XOR2X1   g3510(.A(CRC_OUT_4_16), .B(WX7330), .Y(n9241));
NOR2X1   g3511(.A(n9241), .B(n5827), .Y(CRC_OUT_4_17));
XOR2X1   g3512(.A(CRC_OUT_4_17), .B(WX7328), .Y(n9243));
NOR2X1   g3513(.A(n9243), .B(n5827), .Y(CRC_OUT_4_18));
XOR2X1   g3514(.A(CRC_OUT_4_18), .B(WX7326), .Y(n9245));
NOR2X1   g3515(.A(n9245), .B(n5827), .Y(CRC_OUT_4_19));
XOR2X1   g3516(.A(CRC_OUT_4_19), .B(WX7324), .Y(n9247));
NOR2X1   g3517(.A(n9247), .B(n5827), .Y(CRC_OUT_4_20));
XOR2X1   g3518(.A(CRC_OUT_4_20), .B(WX7322), .Y(n9249));
NOR2X1   g3519(.A(n9249), .B(n5827), .Y(CRC_OUT_4_21));
XOR2X1   g3520(.A(CRC_OUT_4_21), .B(WX7320), .Y(n9251));
NOR2X1   g3521(.A(n9251), .B(n5827), .Y(CRC_OUT_4_22));
XOR2X1   g3522(.A(CRC_OUT_4_22), .B(WX7318), .Y(n9253));
NOR2X1   g3523(.A(n9253), .B(n5827), .Y(CRC_OUT_4_23));
XOR2X1   g3524(.A(CRC_OUT_4_23), .B(WX7316), .Y(n9255));
NOR2X1   g3525(.A(n9255), .B(n5827), .Y(CRC_OUT_4_24));
XOR2X1   g3526(.A(CRC_OUT_4_24), .B(WX7314), .Y(n9257));
NOR2X1   g3527(.A(n9257), .B(n5827), .Y(CRC_OUT_4_25));
XOR2X1   g3528(.A(CRC_OUT_4_25), .B(WX7312), .Y(n9259));
NOR2X1   g3529(.A(n9259), .B(n5827), .Y(CRC_OUT_4_26));
XOR2X1   g3530(.A(CRC_OUT_4_26), .B(WX7310), .Y(n9261));
NOR2X1   g3531(.A(n9261), .B(n5827), .Y(CRC_OUT_4_27));
XOR2X1   g3532(.A(CRC_OUT_4_27), .B(WX7308), .Y(n9263));
NOR2X1   g3533(.A(n9263), .B(n5827), .Y(CRC_OUT_4_28));
XOR2X1   g3534(.A(CRC_OUT_4_28), .B(WX7306), .Y(n9265));
NOR2X1   g3535(.A(n9265), .B(n5827), .Y(CRC_OUT_4_29));
XOR2X1   g3536(.A(CRC_OUT_4_29), .B(WX7304), .Y(n9267));
NOR2X1   g3537(.A(n9267), .B(n5827), .Y(CRC_OUT_4_30));
XOR2X1   g3538(.A(CRC_OUT_4_30), .B(WX7302), .Y(n9269));
NOR2X1   g3539(.A(n9269), .B(n5827), .Y(CRC_OUT_4_31));
AND2X1   g3540(.A(WX8245), .B(RESET), .Y(n6279));
AND2X1   g3541(.A(WX8247), .B(RESET), .Y(n6284));
AND2X1   g3542(.A(WX8249), .B(RESET), .Y(n6289));
AND2X1   g3543(.A(WX8251), .B(RESET), .Y(n6294));
AND2X1   g3544(.A(WX8253), .B(RESET), .Y(n6299));
AND2X1   g3545(.A(WX8255), .B(RESET), .Y(n6304));
AND2X1   g3546(.A(WX8257), .B(RESET), .Y(n6309));
AND2X1   g3547(.A(WX8259), .B(RESET), .Y(n6314));
AND2X1   g3548(.A(WX8261), .B(RESET), .Y(n6319));
AND2X1   g3549(.A(WX8263), .B(RESET), .Y(n6324));
AND2X1   g3550(.A(WX8265), .B(RESET), .Y(n6329));
AND2X1   g3551(.A(WX8267), .B(RESET), .Y(n6334));
AND2X1   g3552(.A(WX8269), .B(RESET), .Y(n6339));
AND2X1   g3553(.A(WX8271), .B(RESET), .Y(n6344));
AND2X1   g3554(.A(WX8273), .B(RESET), .Y(n6349));
AND2X1   g3555(.A(WX8275), .B(RESET), .Y(n6354));
AND2X1   g3556(.A(WX8277), .B(RESET), .Y(n6359));
AND2X1   g3557(.A(WX8279), .B(RESET), .Y(n6364));
AND2X1   g3558(.A(WX8281), .B(RESET), .Y(n6369));
AND2X1   g3559(.A(WX8283), .B(RESET), .Y(n6374));
AND2X1   g3560(.A(WX8285), .B(RESET), .Y(n6379));
AND2X1   g3561(.A(WX8287), .B(RESET), .Y(n6384));
AND2X1   g3562(.A(WX8289), .B(RESET), .Y(n6389));
AND2X1   g3563(.A(WX8291), .B(RESET), .Y(n6394));
AND2X1   g3564(.A(WX8293), .B(RESET), .Y(n6399));
AND2X1   g3565(.A(WX8295), .B(RESET), .Y(n6404));
AND2X1   g3566(.A(WX8297), .B(RESET), .Y(n6409));
AND2X1   g3567(.A(WX8299), .B(RESET), .Y(n6414));
AND2X1   g3568(.A(WX8301), .B(RESET), .Y(n6419));
AND2X1   g3569(.A(WX8303), .B(RESET), .Y(n6424));
AND2X1   g3570(.A(WX8305), .B(RESET), .Y(n6429));
NOR2X1   g3571(.A(WX8243), .B(n5827), .Y(n6434));
INVX1    g3572(.A(CRC_OUT_3_31), .Y(n9303));
XOR2X1   g3573(.A(WX9696), .B(TM1), .Y(n9304));
XOR2X1   g3574(.A(n9304), .B(WX9760), .Y(n9305));
INVX1    g3575(.A(WX9824), .Y(n9306));
XOR2X1   g3576(.A(WX9888), .B(n9306), .Y(n9307));
XOR2X1   g3577(.A(n9307), .B(n9305), .Y(n9308));
MX2X1    g3578(.A(n9303), .B(n9308), .S0(n5539), .Y(n9310));
INVX1    g3579(.A(WX8243), .Y(n9311));
MX2X1    g3580(.A(n9311), .B(n8729), .S0(n5539), .Y(n9312));
MX2X1    g3581(.A(n9310), .B(n9312), .S0(TM1), .Y(n9313));
NOR2X1   g3582(.A(n9313), .B(n5827), .Y(n6439));
INVX1    g3583(.A(CRC_OUT_3_30), .Y(n9315));
XOR2X1   g3584(.A(WX9698), .B(TM1), .Y(n9316));
XOR2X1   g3585(.A(n9316), .B(WX9762), .Y(n9317));
INVX1    g3586(.A(WX9826), .Y(n9318));
XOR2X1   g3587(.A(WX9890), .B(n9318), .Y(n9319));
XOR2X1   g3588(.A(n9319), .B(n9317), .Y(n9320));
MX2X1    g3589(.A(n9315), .B(n9320), .S0(n5539), .Y(n9322));
INVX1    g3590(.A(WX8245), .Y(n9323));
MX2X1    g3591(.A(n9323), .B(n8741), .S0(n5539), .Y(n9324));
MX2X1    g3592(.A(n9322), .B(n9324), .S0(TM1), .Y(n9325));
NOR2X1   g3593(.A(n9325), .B(n5827), .Y(n6444));
INVX1    g3594(.A(CRC_OUT_3_29), .Y(n9327));
XOR2X1   g3595(.A(WX9700), .B(TM1), .Y(n9328));
XOR2X1   g3596(.A(n9328), .B(WX9764), .Y(n9329));
INVX1    g3597(.A(WX9828), .Y(n9330));
XOR2X1   g3598(.A(WX9892), .B(n9330), .Y(n9331));
XOR2X1   g3599(.A(n9331), .B(n9329), .Y(n9332));
MX2X1    g3600(.A(n9327), .B(n9332), .S0(n5539), .Y(n9334));
INVX1    g3601(.A(WX8247), .Y(n9335));
MX2X1    g3602(.A(n9335), .B(n8753), .S0(n5539), .Y(n9336));
MX2X1    g3603(.A(n9334), .B(n9336), .S0(TM1), .Y(n9337));
NOR2X1   g3604(.A(n9337), .B(n5827), .Y(n6449));
INVX1    g3605(.A(CRC_OUT_3_28), .Y(n9339));
XOR2X1   g3606(.A(WX9702), .B(TM1), .Y(n9340));
XOR2X1   g3607(.A(n9340), .B(WX9766), .Y(n9341));
INVX1    g3608(.A(WX9830), .Y(n9342));
XOR2X1   g3609(.A(WX9894), .B(n9342), .Y(n9343));
XOR2X1   g3610(.A(n9343), .B(n9341), .Y(n9344));
MX2X1    g3611(.A(n9339), .B(n9344), .S0(n5539), .Y(n9346));
INVX1    g3612(.A(WX8249), .Y(n9347));
MX2X1    g3613(.A(n9347), .B(n8765_1), .S0(n5539), .Y(n9348));
MX2X1    g3614(.A(n9346), .B(n9348), .S0(TM1), .Y(n9349));
NOR2X1   g3615(.A(n9349), .B(n5827), .Y(n6454));
INVX1    g3616(.A(CRC_OUT_3_27), .Y(n9351));
XOR2X1   g3617(.A(WX9704), .B(TM1), .Y(n9352));
XOR2X1   g3618(.A(n9352), .B(WX9768), .Y(n9353));
INVX1    g3619(.A(WX9832), .Y(n9354));
XOR2X1   g3620(.A(WX9896), .B(n9354), .Y(n9355));
XOR2X1   g3621(.A(n9355), .B(n9353), .Y(n9356));
MX2X1    g3622(.A(n9351), .B(n9356), .S0(n5539), .Y(n9358));
INVX1    g3623(.A(WX8251), .Y(n9359));
MX2X1    g3624(.A(n9359), .B(n8777), .S0(n5539), .Y(n9360));
MX2X1    g3625(.A(n9358), .B(n9360), .S0(TM1), .Y(n9361));
NOR2X1   g3626(.A(n9361), .B(n5827), .Y(n6459));
INVX1    g3627(.A(CRC_OUT_3_26), .Y(n9363));
XOR2X1   g3628(.A(WX9706), .B(TM1), .Y(n9364));
XOR2X1   g3629(.A(n9364), .B(WX9770), .Y(n9365));
INVX1    g3630(.A(WX9834), .Y(n9366));
XOR2X1   g3631(.A(WX9898), .B(n9366), .Y(n9367));
XOR2X1   g3632(.A(n9367), .B(n9365), .Y(n9368));
MX2X1    g3633(.A(n9363), .B(n9368), .S0(n5539), .Y(n9370));
INVX1    g3634(.A(WX8253), .Y(n9371));
MX2X1    g3635(.A(n9371), .B(n8789), .S0(n5539), .Y(n9372));
MX2X1    g3636(.A(n9370), .B(n9372), .S0(TM1), .Y(n9373));
NOR2X1   g3637(.A(n9373), .B(n5827), .Y(n6464));
INVX1    g3638(.A(CRC_OUT_3_25), .Y(n9375));
XOR2X1   g3639(.A(WX9708), .B(TM1), .Y(n9376));
XOR2X1   g3640(.A(n9376), .B(WX9772), .Y(n9377));
INVX1    g3641(.A(WX9836), .Y(n9378));
XOR2X1   g3642(.A(WX9900), .B(n9378), .Y(n9379));
XOR2X1   g3643(.A(n9379), .B(n9377), .Y(n9380));
MX2X1    g3644(.A(n9375), .B(n9380), .S0(n5539), .Y(n9382));
INVX1    g3645(.A(WX8255), .Y(n9383));
MX2X1    g3646(.A(n9383), .B(n8801), .S0(n5539), .Y(n9384));
MX2X1    g3647(.A(n9382), .B(n9384), .S0(TM1), .Y(n9385));
NOR2X1   g3648(.A(n9385), .B(n5827), .Y(n6469));
INVX1    g3649(.A(CRC_OUT_3_24), .Y(n9387));
XOR2X1   g3650(.A(WX9710), .B(TM1), .Y(n9388));
XOR2X1   g3651(.A(n9388), .B(WX9774), .Y(n9389));
INVX1    g3652(.A(WX9838), .Y(n9390));
XOR2X1   g3653(.A(WX9902), .B(n9390), .Y(n9391));
XOR2X1   g3654(.A(n9391), .B(n9389), .Y(n9392));
MX2X1    g3655(.A(n9387), .B(n9392), .S0(n5539), .Y(n9394));
INVX1    g3656(.A(WX8257), .Y(n9395));
MX2X1    g3657(.A(n9395), .B(n8813), .S0(n5539), .Y(n9396));
MX2X1    g3658(.A(n9394), .B(n9396), .S0(TM1), .Y(n9397));
NOR2X1   g3659(.A(n9397), .B(n5827), .Y(n6474));
INVX1    g3660(.A(CRC_OUT_3_23), .Y(n9399));
XOR2X1   g3661(.A(WX9712), .B(TM1), .Y(n9400));
XOR2X1   g3662(.A(n9400), .B(WX9776), .Y(n9401));
INVX1    g3663(.A(WX9840), .Y(n9402));
XOR2X1   g3664(.A(WX9904), .B(n9402), .Y(n9403));
XOR2X1   g3665(.A(n9403), .B(n9401), .Y(n9404));
MX2X1    g3666(.A(n9399), .B(n9404), .S0(n5539), .Y(n9406));
INVX1    g3667(.A(WX8259), .Y(n9407));
MX2X1    g3668(.A(n9407), .B(n8825_1), .S0(n5539), .Y(n9408));
MX2X1    g3669(.A(n9406), .B(n9408), .S0(TM1), .Y(n9409));
NOR2X1   g3670(.A(n9409), .B(n5827), .Y(n6479));
INVX1    g3671(.A(CRC_OUT_3_22), .Y(n9411));
XOR2X1   g3672(.A(WX9714), .B(TM1), .Y(n9412));
XOR2X1   g3673(.A(n9412), .B(WX9778), .Y(n9413));
INVX1    g3674(.A(WX9842), .Y(n9414));
XOR2X1   g3675(.A(WX9906), .B(n9414), .Y(n9415));
XOR2X1   g3676(.A(n9415), .B(n9413), .Y(n9416));
MX2X1    g3677(.A(n9411), .B(n9416), .S0(n5539), .Y(n9418));
INVX1    g3678(.A(WX8261), .Y(n9419));
MX2X1    g3679(.A(n9419), .B(n8837), .S0(n5539), .Y(n9420));
MX2X1    g3680(.A(n9418), .B(n9420), .S0(TM1), .Y(n9421));
NOR2X1   g3681(.A(n9421), .B(n5827), .Y(n6484));
INVX1    g3682(.A(CRC_OUT_3_21), .Y(n9423));
XOR2X1   g3683(.A(WX9716), .B(TM1), .Y(n9424));
XOR2X1   g3684(.A(n9424), .B(WX9780), .Y(n9425));
INVX1    g3685(.A(WX9844), .Y(n9426));
XOR2X1   g3686(.A(WX9908), .B(n9426), .Y(n9427));
XOR2X1   g3687(.A(n9427), .B(n9425), .Y(n9428));
MX2X1    g3688(.A(n9423), .B(n9428), .S0(n5539), .Y(n9430));
INVX1    g3689(.A(WX8263), .Y(n9431));
MX2X1    g3690(.A(n9431), .B(n8849), .S0(n5539), .Y(n9432));
MX2X1    g3691(.A(n9430), .B(n9432), .S0(TM1), .Y(n9433));
NOR2X1   g3692(.A(n9433), .B(n5827), .Y(n6489));
INVX1    g3693(.A(CRC_OUT_3_20), .Y(n9435));
XOR2X1   g3694(.A(WX9718), .B(TM1), .Y(n9436));
XOR2X1   g3695(.A(n9436), .B(WX9782), .Y(n9437));
INVX1    g3696(.A(WX9846), .Y(n9438));
XOR2X1   g3697(.A(WX9910), .B(n9438), .Y(n9439));
XOR2X1   g3698(.A(n9439), .B(n9437), .Y(n9440));
MX2X1    g3699(.A(n9435), .B(n9440), .S0(n5539), .Y(n9442));
INVX1    g3700(.A(WX8265), .Y(n9443));
MX2X1    g3701(.A(n9443), .B(n8861), .S0(n5539), .Y(n9444));
MX2X1    g3702(.A(n9442), .B(n9444), .S0(TM1), .Y(n9445));
NOR2X1   g3703(.A(n9445), .B(n5827), .Y(n6494));
INVX1    g3704(.A(CRC_OUT_3_19), .Y(n9447));
XOR2X1   g3705(.A(WX9720), .B(TM1), .Y(n9448));
XOR2X1   g3706(.A(n9448), .B(WX9784), .Y(n9449));
INVX1    g3707(.A(WX9848), .Y(n9450));
XOR2X1   g3708(.A(WX9912), .B(n9450), .Y(n9451));
XOR2X1   g3709(.A(n9451), .B(n9449), .Y(n9452));
MX2X1    g3710(.A(n9447), .B(n9452), .S0(n5539), .Y(n9454));
INVX1    g3711(.A(WX8267), .Y(n9455));
MX2X1    g3712(.A(n9455), .B(n8873), .S0(n5539), .Y(n9456));
MX2X1    g3713(.A(n9454), .B(n9456), .S0(TM1), .Y(n9457));
NOR2X1   g3714(.A(n9457), .B(n5827), .Y(n6499));
INVX1    g3715(.A(CRC_OUT_3_18), .Y(n9459));
XOR2X1   g3716(.A(WX9722), .B(TM1), .Y(n9460));
XOR2X1   g3717(.A(n9460), .B(WX9786), .Y(n9461));
INVX1    g3718(.A(WX9850), .Y(n9462));
XOR2X1   g3719(.A(WX9914), .B(n9462), .Y(n9463));
XOR2X1   g3720(.A(n9463), .B(n9461), .Y(n9464));
MX2X1    g3721(.A(n9459), .B(n9464), .S0(n5539), .Y(n9466));
INVX1    g3722(.A(WX8269), .Y(n9467));
MX2X1    g3723(.A(n9467), .B(n8885_1), .S0(n5539), .Y(n9468));
MX2X1    g3724(.A(n9466), .B(n9468), .S0(TM1), .Y(n9469));
NOR2X1   g3725(.A(n9469), .B(n5827), .Y(n6504));
INVX1    g3726(.A(CRC_OUT_3_17), .Y(n9471));
XOR2X1   g3727(.A(WX9724), .B(TM1), .Y(n9472));
XOR2X1   g3728(.A(n9472), .B(WX9788), .Y(n9473));
INVX1    g3729(.A(WX9852), .Y(n9474));
XOR2X1   g3730(.A(WX9916), .B(n9474), .Y(n9475));
XOR2X1   g3731(.A(n9475), .B(n9473), .Y(n9476));
MX2X1    g3732(.A(n9471), .B(n9476), .S0(n5539), .Y(n9478));
INVX1    g3733(.A(WX8271), .Y(n9479));
MX2X1    g3734(.A(n9479), .B(n8897), .S0(n5539), .Y(n9480));
MX2X1    g3735(.A(n9478), .B(n9480), .S0(TM1), .Y(n9481));
NOR2X1   g3736(.A(n9481), .B(n5827), .Y(n6509));
INVX1    g3737(.A(CRC_OUT_3_16), .Y(n9483));
XOR2X1   g3738(.A(WX9726), .B(TM1), .Y(n9484));
XOR2X1   g3739(.A(n9484), .B(WX9790), .Y(n9485));
INVX1    g3740(.A(WX9854), .Y(n9486));
XOR2X1   g3741(.A(WX9918), .B(n9486), .Y(n9487));
XOR2X1   g3742(.A(n9487), .B(n9485), .Y(n9488));
MX2X1    g3743(.A(n9483), .B(n9488), .S0(n5539), .Y(n9490));
INVX1    g3744(.A(WX8273), .Y(n9491));
MX2X1    g3745(.A(n9491), .B(n8909), .S0(n5539), .Y(n9492));
MX2X1    g3746(.A(n9490), .B(n9492), .S0(TM1), .Y(n9493));
NOR2X1   g3747(.A(n9493), .B(n5827), .Y(n6514));
INVX1    g3748(.A(CRC_OUT_3_15), .Y(n9495));
XOR2X1   g3749(.A(WX9728), .B(TM0), .Y(n9496));
XOR2X1   g3750(.A(n9496), .B(WX9792), .Y(n9497));
INVX1    g3751(.A(WX9856), .Y(n9498));
XOR2X1   g3752(.A(WX9920), .B(n9498), .Y(n9499));
XOR2X1   g3753(.A(n9499), .B(n9497), .Y(n9500));
MX2X1    g3754(.A(n9495), .B(n9500), .S0(n5539), .Y(n9502));
INVX1    g3755(.A(WX8275), .Y(n9503));
MX2X1    g3756(.A(n9503), .B(n8921), .S0(n5539), .Y(n9504));
MX2X1    g3757(.A(n9502), .B(n9504), .S0(TM1), .Y(n9505));
NOR2X1   g3758(.A(n9505), .B(n5827), .Y(n6519));
INVX1    g3759(.A(CRC_OUT_3_14), .Y(n9507));
XOR2X1   g3760(.A(WX9730), .B(TM0), .Y(n9508));
XOR2X1   g3761(.A(n9508), .B(WX9794), .Y(n9509));
INVX1    g3762(.A(WX9858), .Y(n9510));
XOR2X1   g3763(.A(WX9922), .B(n9510), .Y(n9511));
XOR2X1   g3764(.A(n9511), .B(n9509), .Y(n9512));
MX2X1    g3765(.A(n9507), .B(n9512), .S0(n5539), .Y(n9514));
INVX1    g3766(.A(WX8277), .Y(n9515));
MX2X1    g3767(.A(n9515), .B(n8933), .S0(n5539), .Y(n9516));
MX2X1    g3768(.A(n9514), .B(n9516), .S0(TM1), .Y(n9517));
NOR2X1   g3769(.A(n9517), .B(n5827), .Y(n6524));
INVX1    g3770(.A(CRC_OUT_3_13), .Y(n9519));
XOR2X1   g3771(.A(WX9732), .B(TM0), .Y(n9520));
XOR2X1   g3772(.A(n9520), .B(WX9796), .Y(n9521));
INVX1    g3773(.A(WX9860), .Y(n9522));
XOR2X1   g3774(.A(WX9924), .B(n9522), .Y(n9523));
XOR2X1   g3775(.A(n9523), .B(n9521), .Y(n9524));
MX2X1    g3776(.A(n9519), .B(n9524), .S0(n5539), .Y(n9526));
INVX1    g3777(.A(WX8279), .Y(n9527));
MX2X1    g3778(.A(n9527), .B(n8945), .S0(n5539), .Y(n9528));
MX2X1    g3779(.A(n9526), .B(n9528), .S0(TM1), .Y(n9529));
NOR2X1   g3780(.A(n9529), .B(n5827), .Y(n6529));
INVX1    g3781(.A(CRC_OUT_3_12), .Y(n9531));
XOR2X1   g3782(.A(WX9734), .B(TM0), .Y(n9532));
XOR2X1   g3783(.A(n9532), .B(WX9798), .Y(n9533));
INVX1    g3784(.A(WX9862), .Y(n9534));
XOR2X1   g3785(.A(WX9926), .B(n9534), .Y(n9535));
XOR2X1   g3786(.A(n9535), .B(n9533), .Y(n9536));
MX2X1    g3787(.A(n9531), .B(n9536), .S0(n5539), .Y(n9538));
INVX1    g3788(.A(WX8281), .Y(n9539));
MX2X1    g3789(.A(n9539), .B(n8957), .S0(n5539), .Y(n9540));
MX2X1    g3790(.A(n9538), .B(n9540), .S0(TM1), .Y(n9541));
NOR2X1   g3791(.A(n9541), .B(n5827), .Y(n6534));
INVX1    g3792(.A(CRC_OUT_3_11), .Y(n9543));
XOR2X1   g3793(.A(WX9736), .B(TM0), .Y(n9544));
XOR2X1   g3794(.A(n9544), .B(WX9800), .Y(n9545));
INVX1    g3795(.A(WX9864), .Y(n9546));
XOR2X1   g3796(.A(WX9928), .B(n9546), .Y(n9547));
XOR2X1   g3797(.A(n9547), .B(n9545), .Y(n9548));
MX2X1    g3798(.A(n9543), .B(n9548), .S0(n5539), .Y(n9550));
INVX1    g3799(.A(WX8283), .Y(n9551));
MX2X1    g3800(.A(n9551), .B(n8969), .S0(n5539), .Y(n9552));
MX2X1    g3801(.A(n9550), .B(n9552), .S0(TM1), .Y(n9553));
NOR2X1   g3802(.A(n9553), .B(n5827), .Y(n6539));
INVX1    g3803(.A(CRC_OUT_3_10), .Y(n9555));
XOR2X1   g3804(.A(WX9738), .B(TM0), .Y(n9556));
XOR2X1   g3805(.A(n9556), .B(WX9802), .Y(n9557));
INVX1    g3806(.A(WX9866), .Y(n9558));
XOR2X1   g3807(.A(WX9930), .B(n9558), .Y(n9559));
XOR2X1   g3808(.A(n9559), .B(n9557), .Y(n9560));
MX2X1    g3809(.A(n9555), .B(n9560), .S0(n5539), .Y(n9562));
INVX1    g3810(.A(WX8285), .Y(n9563));
MX2X1    g3811(.A(n9563), .B(n8981), .S0(n5539), .Y(n9564));
MX2X1    g3812(.A(n9562), .B(n9564), .S0(TM1), .Y(n9565));
NOR2X1   g3813(.A(n9565), .B(n5827), .Y(n6544));
INVX1    g3814(.A(CRC_OUT_3_9), .Y(n9567));
XOR2X1   g3815(.A(WX9740), .B(TM0), .Y(n9568));
XOR2X1   g3816(.A(n9568), .B(WX9804), .Y(n9569));
INVX1    g3817(.A(WX9868), .Y(n9570));
XOR2X1   g3818(.A(WX9932), .B(n9570), .Y(n9571));
XOR2X1   g3819(.A(n9571), .B(n9569), .Y(n9572));
MX2X1    g3820(.A(n9567), .B(n9572), .S0(n5539), .Y(n9574));
INVX1    g3821(.A(WX8287), .Y(n9575));
MX2X1    g3822(.A(n9575), .B(n8993), .S0(n5539), .Y(n9576));
MX2X1    g3823(.A(n9574), .B(n9576), .S0(TM1), .Y(n9577));
NOR2X1   g3824(.A(n9577), .B(n5827), .Y(n6549));
INVX1    g3825(.A(CRC_OUT_3_8), .Y(n9579));
XOR2X1   g3826(.A(WX9742), .B(TM0), .Y(n9580));
XOR2X1   g3827(.A(n9580), .B(WX9806), .Y(n9581));
INVX1    g3828(.A(WX9870), .Y(n9582));
XOR2X1   g3829(.A(WX9934), .B(n9582), .Y(n9583));
XOR2X1   g3830(.A(n9583), .B(n9581), .Y(n9584));
MX2X1    g3831(.A(n9579), .B(n9584), .S0(n5539), .Y(n9586));
INVX1    g3832(.A(WX8289), .Y(n9587));
MX2X1    g3833(.A(n9587), .B(n9005), .S0(n5539), .Y(n9588));
MX2X1    g3834(.A(n9586), .B(n9588), .S0(TM1), .Y(n9589));
NOR2X1   g3835(.A(n9589), .B(n5827), .Y(n6554));
INVX1    g3836(.A(CRC_OUT_3_7), .Y(n9591));
XOR2X1   g3837(.A(WX9744), .B(TM0), .Y(n9592));
XOR2X1   g3838(.A(n9592), .B(WX9808), .Y(n9593));
INVX1    g3839(.A(WX9872), .Y(n9594));
XOR2X1   g3840(.A(WX9936), .B(n9594), .Y(n9595));
XOR2X1   g3841(.A(n9595), .B(n9593), .Y(n9596));
MX2X1    g3842(.A(n9591), .B(n9596), .S0(n5539), .Y(n9598));
INVX1    g3843(.A(WX8291), .Y(n9599));
MX2X1    g3844(.A(n9599), .B(n9017), .S0(n5539), .Y(n9600));
MX2X1    g3845(.A(n9598), .B(n9600), .S0(TM1), .Y(n9601));
NOR2X1   g3846(.A(n9601), .B(n5827), .Y(n6559));
INVX1    g3847(.A(CRC_OUT_3_6), .Y(n9603));
XOR2X1   g3848(.A(WX9746), .B(TM0), .Y(n9604));
XOR2X1   g3849(.A(n9604), .B(WX9810), .Y(n9605));
INVX1    g3850(.A(WX9874), .Y(n9606));
XOR2X1   g3851(.A(WX9938), .B(n9606), .Y(n9607));
XOR2X1   g3852(.A(n9607), .B(n9605), .Y(n9608));
MX2X1    g3853(.A(n9603), .B(n9608), .S0(n5539), .Y(n9610));
INVX1    g3854(.A(WX8293), .Y(n9611));
MX2X1    g3855(.A(n9611), .B(n9029), .S0(n5539), .Y(n9612));
MX2X1    g3856(.A(n9610), .B(n9612), .S0(TM1), .Y(n9613));
NOR2X1   g3857(.A(n9613), .B(n5827), .Y(n6564));
INVX1    g3858(.A(CRC_OUT_3_5), .Y(n9615));
XOR2X1   g3859(.A(WX9748), .B(TM0), .Y(n9616));
XOR2X1   g3860(.A(n9616), .B(WX9812), .Y(n9617));
INVX1    g3861(.A(WX9876), .Y(n9618));
XOR2X1   g3862(.A(WX9940), .B(n9618), .Y(n9619));
XOR2X1   g3863(.A(n9619), .B(n9617), .Y(n9620));
MX2X1    g3864(.A(n9615), .B(n9620), .S0(n5539), .Y(n9622));
INVX1    g3865(.A(WX8295), .Y(n9623));
MX2X1    g3866(.A(n9623), .B(n9041), .S0(n5539), .Y(n9624));
MX2X1    g3867(.A(n9622), .B(n9624), .S0(TM1), .Y(n9625));
NOR2X1   g3868(.A(n9625), .B(n5827), .Y(n6569));
INVX1    g3869(.A(CRC_OUT_3_4), .Y(n9627));
XOR2X1   g3870(.A(WX9750), .B(TM0), .Y(n9628));
XOR2X1   g3871(.A(n9628), .B(WX9814), .Y(n9629));
INVX1    g3872(.A(WX9878), .Y(n9630));
XOR2X1   g3873(.A(WX9942), .B(n9630), .Y(n9631));
XOR2X1   g3874(.A(n9631), .B(n9629), .Y(n9632));
MX2X1    g3875(.A(n9627), .B(n9632), .S0(n5539), .Y(n9634));
INVX1    g3876(.A(WX8297), .Y(n9635));
MX2X1    g3877(.A(n9635), .B(n9053), .S0(n5539), .Y(n9636));
MX2X1    g3878(.A(n9634), .B(n9636), .S0(TM1), .Y(n9637));
NOR2X1   g3879(.A(n9637), .B(n5827), .Y(n6574));
INVX1    g3880(.A(CRC_OUT_3_3), .Y(n9639));
XOR2X1   g3881(.A(WX9752), .B(TM0), .Y(n9640));
XOR2X1   g3882(.A(n9640), .B(WX9816), .Y(n9641));
INVX1    g3883(.A(WX9880), .Y(n9642));
XOR2X1   g3884(.A(WX9944), .B(n9642), .Y(n9643));
XOR2X1   g3885(.A(n9643), .B(n9641), .Y(n9644));
MX2X1    g3886(.A(n9639), .B(n9644), .S0(n5539), .Y(n9646));
INVX1    g3887(.A(WX8299), .Y(n9647));
MX2X1    g3888(.A(n9647), .B(n9065), .S0(n5539), .Y(n9648));
MX2X1    g3889(.A(n9646), .B(n9648), .S0(TM1), .Y(n9649));
NOR2X1   g3890(.A(n9649), .B(n5827), .Y(n6579));
INVX1    g3891(.A(CRC_OUT_3_2), .Y(n9651));
XOR2X1   g3892(.A(WX9754), .B(TM0), .Y(n9652));
XOR2X1   g3893(.A(n9652), .B(WX9818), .Y(n9653));
INVX1    g3894(.A(WX9882), .Y(n9654));
XOR2X1   g3895(.A(WX9946), .B(n9654), .Y(n9655));
XOR2X1   g3896(.A(n9655), .B(n9653), .Y(n9656));
MX2X1    g3897(.A(n9651), .B(n9656), .S0(n5539), .Y(n9658));
INVX1    g3898(.A(WX8301), .Y(n9659));
MX2X1    g3899(.A(n9659), .B(n9077), .S0(n5539), .Y(n9660));
MX2X1    g3900(.A(n9658), .B(n9660), .S0(TM1), .Y(n9661));
NOR2X1   g3901(.A(n9661), .B(n5827), .Y(n6584));
INVX1    g3902(.A(CRC_OUT_3_1), .Y(n9663));
XOR2X1   g3903(.A(WX9756), .B(TM0), .Y(n9664));
XOR2X1   g3904(.A(n9664), .B(WX9820), .Y(n9665));
INVX1    g3905(.A(WX9884), .Y(n9666));
XOR2X1   g3906(.A(WX9948), .B(n9666), .Y(n9667));
XOR2X1   g3907(.A(n9667), .B(n9665), .Y(n9668));
MX2X1    g3908(.A(n9663), .B(n9668), .S0(n5539), .Y(n9670));
INVX1    g3909(.A(WX8303), .Y(n9671));
MX2X1    g3910(.A(n9671), .B(n9089), .S0(n5539), .Y(n9672));
MX2X1    g3911(.A(n9670), .B(n9672), .S0(TM1), .Y(n9673));
NOR2X1   g3912(.A(n9673), .B(n5827), .Y(n6589));
INVX1    g3913(.A(CRC_OUT_3_0), .Y(n9675));
XOR2X1   g3914(.A(WX9758), .B(TM0), .Y(n9676));
XOR2X1   g3915(.A(n9676), .B(WX9822), .Y(n9677));
INVX1    g3916(.A(WX9886), .Y(n9678));
XOR2X1   g3917(.A(WX9950), .B(n9678), .Y(n9679));
XOR2X1   g3918(.A(n9679), .B(n9677), .Y(n9680));
MX2X1    g3919(.A(n9675), .B(n9680), .S0(n5539), .Y(n9682));
INVX1    g3920(.A(WX8305), .Y(n9683));
MX2X1    g3921(.A(n9683), .B(n9101), .S0(n5539), .Y(n9684));
MX2X1    g3922(.A(n9682), .B(n9684), .S0(TM1), .Y(n9685));
NOR2X1   g3923(.A(n9685), .B(n5827), .Y(n6594));
AND2X1   g3924(.A(WX8403), .B(RESET), .Y(n6599));
AND2X1   g3925(.A(WX8405), .B(RESET), .Y(n6604));
AND2X1   g3926(.A(WX8407), .B(RESET), .Y(n6609));
AND2X1   g3927(.A(WX8409), .B(RESET), .Y(n6614));
AND2X1   g3928(.A(WX8411), .B(RESET), .Y(n6619));
AND2X1   g3929(.A(WX8413), .B(RESET), .Y(n6624));
AND2X1   g3930(.A(WX8415), .B(RESET), .Y(n6629));
AND2X1   g3931(.A(WX8417), .B(RESET), .Y(n6634));
AND2X1   g3932(.A(WX8419), .B(RESET), .Y(n6639));
AND2X1   g3933(.A(WX8421), .B(RESET), .Y(n6644));
AND2X1   g3934(.A(WX8423), .B(RESET), .Y(n6649));
AND2X1   g3935(.A(WX8425), .B(RESET), .Y(n6654));
AND2X1   g3936(.A(WX8427), .B(RESET), .Y(n6659));
AND2X1   g3937(.A(WX8429), .B(RESET), .Y(n6664));
AND2X1   g3938(.A(WX8431), .B(RESET), .Y(n6669));
AND2X1   g3939(.A(WX8433), .B(RESET), .Y(n6674));
AND2X1   g3940(.A(WX8435), .B(RESET), .Y(n6679));
AND2X1   g3941(.A(WX8437), .B(RESET), .Y(n6684));
AND2X1   g3942(.A(WX8439), .B(RESET), .Y(n6689));
AND2X1   g3943(.A(WX8441), .B(RESET), .Y(n6694));
AND2X1   g3944(.A(WX8443), .B(RESET), .Y(n6699));
AND2X1   g3945(.A(WX8445), .B(RESET), .Y(n6704));
AND2X1   g3946(.A(WX8447), .B(RESET), .Y(n6709));
AND2X1   g3947(.A(WX8449), .B(RESET), .Y(n6714));
AND2X1   g3948(.A(WX8451), .B(RESET), .Y(n6719));
AND2X1   g3949(.A(WX8453), .B(RESET), .Y(n6724));
AND2X1   g3950(.A(WX8455), .B(RESET), .Y(n6729));
AND2X1   g3951(.A(WX8457), .B(RESET), .Y(n6734));
AND2X1   g3952(.A(WX8459), .B(RESET), .Y(n6739));
AND2X1   g3953(.A(WX8461), .B(RESET), .Y(n6744));
AND2X1   g3954(.A(WX8463), .B(RESET), .Y(n6749));
AND2X1   g3955(.A(WX8465), .B(RESET), .Y(n6754));
AND2X1   g3956(.A(WX8467), .B(RESET), .Y(n6759));
AND2X1   g3957(.A(WX8469), .B(RESET), .Y(n6764));
AND2X1   g3958(.A(WX8471), .B(RESET), .Y(n6769));
AND2X1   g3959(.A(WX8473), .B(RESET), .Y(n6774));
AND2X1   g3960(.A(WX8475), .B(RESET), .Y(n6779));
AND2X1   g3961(.A(WX8477), .B(RESET), .Y(n6784));
AND2X1   g3962(.A(WX8479), .B(RESET), .Y(n6789));
AND2X1   g3963(.A(WX8481), .B(RESET), .Y(n6794));
AND2X1   g3964(.A(WX8483), .B(RESET), .Y(n6799));
AND2X1   g3965(.A(WX8485), .B(RESET), .Y(n6804));
AND2X1   g3966(.A(WX8487), .B(RESET), .Y(n6809));
AND2X1   g3967(.A(WX8489), .B(RESET), .Y(n6814));
AND2X1   g3968(.A(WX8491), .B(RESET), .Y(n6819));
AND2X1   g3969(.A(WX8493), .B(RESET), .Y(n6824));
AND2X1   g3970(.A(WX8495), .B(RESET), .Y(n6829));
AND2X1   g3971(.A(WX8497), .B(RESET), .Y(n6834));
AND2X1   g3972(.A(WX8499), .B(RESET), .Y(n6839));
AND2X1   g3973(.A(WX8501), .B(RESET), .Y(n6844));
AND2X1   g3974(.A(WX8503), .B(RESET), .Y(n6849));
AND2X1   g3975(.A(WX8505), .B(RESET), .Y(n6854));
AND2X1   g3976(.A(WX8507), .B(RESET), .Y(n6859));
AND2X1   g3977(.A(WX8509), .B(RESET), .Y(n6864));
AND2X1   g3978(.A(WX8511), .B(RESET), .Y(n6869));
AND2X1   g3979(.A(WX8513), .B(RESET), .Y(n6874));
AND2X1   g3980(.A(WX8515), .B(RESET), .Y(n6879));
AND2X1   g3981(.A(WX8517), .B(RESET), .Y(n6884));
AND2X1   g3982(.A(WX8519), .B(RESET), .Y(n6889));
AND2X1   g3983(.A(WX8521), .B(RESET), .Y(n6894));
AND2X1   g3984(.A(WX8523), .B(RESET), .Y(n6899));
AND2X1   g3985(.A(WX8525), .B(RESET), .Y(n6904));
AND2X1   g3986(.A(WX8527), .B(RESET), .Y(n6909));
AND2X1   g3987(.A(WX8529), .B(RESET), .Y(n6914));
AND2X1   g3988(.A(WX8531), .B(RESET), .Y(n6919));
AND2X1   g3989(.A(WX8533), .B(RESET), .Y(n6924));
AND2X1   g3990(.A(WX8535), .B(RESET), .Y(n6929));
AND2X1   g3991(.A(WX8537), .B(RESET), .Y(n6934));
AND2X1   g3992(.A(WX8539), .B(RESET), .Y(n6939));
AND2X1   g3993(.A(WX8541), .B(RESET), .Y(n6944));
AND2X1   g3994(.A(WX8543), .B(RESET), .Y(n6949));
AND2X1   g3995(.A(WX8545), .B(RESET), .Y(n6954));
AND2X1   g3996(.A(WX8547), .B(RESET), .Y(n6959));
AND2X1   g3997(.A(WX8549), .B(RESET), .Y(n6964));
AND2X1   g3998(.A(WX8551), .B(RESET), .Y(n6969));
AND2X1   g3999(.A(WX8553), .B(RESET), .Y(n6974));
AND2X1   g4000(.A(WX8555), .B(RESET), .Y(n6979));
AND2X1   g4001(.A(WX8557), .B(RESET), .Y(n6984));
AND2X1   g4002(.A(WX8559), .B(RESET), .Y(n6989));
AND2X1   g4003(.A(WX8561), .B(RESET), .Y(n6994));
AND2X1   g4004(.A(WX8563), .B(RESET), .Y(n6999));
AND2X1   g4005(.A(WX8565), .B(RESET), .Y(n7004));
AND2X1   g4006(.A(WX8567), .B(RESET), .Y(n7009));
AND2X1   g4007(.A(WX8569), .B(RESET), .Y(n7014));
AND2X1   g4008(.A(WX8571), .B(RESET), .Y(n7019));
AND2X1   g4009(.A(WX8573), .B(RESET), .Y(n7024));
AND2X1   g4010(.A(WX8575), .B(RESET), .Y(n7029));
AND2X1   g4011(.A(WX8577), .B(RESET), .Y(n7034));
AND2X1   g4012(.A(WX8579), .B(RESET), .Y(n7039));
AND2X1   g4013(.A(WX8581), .B(RESET), .Y(n7044));
AND2X1   g4014(.A(WX8583), .B(RESET), .Y(n7049));
AND2X1   g4015(.A(WX8585), .B(RESET), .Y(n7054));
AND2X1   g4016(.A(WX8587), .B(RESET), .Y(n7059));
AND2X1   g4017(.A(WX8589), .B(RESET), .Y(n7064));
AND2X1   g4018(.A(WX8591), .B(RESET), .Y(n7069));
AND2X1   g4019(.A(WX8593), .B(RESET), .Y(n7074));
XOR2X1   g4020(.A(CRC_OUT_3_31), .B(WX8657), .Y(n9783));
NOR2X1   g4021(.A(n9783), .B(n5827), .Y(CRC_OUT_3_0));
XOR2X1   g4022(.A(CRC_OUT_3_0), .B(WX8655), .Y(n9785));
NOR2X1   g4023(.A(n9785), .B(n5827), .Y(CRC_OUT_3_1));
XOR2X1   g4024(.A(CRC_OUT_3_1), .B(WX8653), .Y(n9787));
NOR2X1   g4025(.A(n9787), .B(n5827), .Y(CRC_OUT_3_2));
XOR2X1   g4026(.A(CRC_OUT_3_2), .B(WX8651), .Y(n9789));
NOR2X1   g4027(.A(n9789), .B(n5827), .Y(CRC_OUT_3_3));
XOR2X1   g4028(.A(CRC_OUT_3_31), .B(WX8649), .Y(n9791));
XOR2X1   g4029(.A(n9791), .B(CRC_OUT_3_3), .Y(n9792));
NOR2X1   g4030(.A(n9792), .B(n5827), .Y(CRC_OUT_3_4));
XOR2X1   g4031(.A(CRC_OUT_3_4), .B(WX8647), .Y(n9794));
NOR2X1   g4032(.A(n9794), .B(n5827), .Y(CRC_OUT_3_5));
XOR2X1   g4033(.A(CRC_OUT_3_5), .B(WX8645), .Y(n9796));
NOR2X1   g4034(.A(n9796), .B(n5827), .Y(CRC_OUT_3_6));
XOR2X1   g4035(.A(CRC_OUT_3_6), .B(WX8643), .Y(n9798));
NOR2X1   g4036(.A(n9798), .B(n5827), .Y(CRC_OUT_3_7));
XOR2X1   g4037(.A(CRC_OUT_3_7), .B(WX8641), .Y(n9800));
NOR2X1   g4038(.A(n9800), .B(n5827), .Y(CRC_OUT_3_8));
XOR2X1   g4039(.A(CRC_OUT_3_8), .B(WX8639), .Y(n9802));
NOR2X1   g4040(.A(n9802), .B(n5827), .Y(CRC_OUT_3_9));
XOR2X1   g4041(.A(CRC_OUT_3_9), .B(WX8637), .Y(n9804));
NOR2X1   g4042(.A(n9804), .B(n5827), .Y(CRC_OUT_3_10));
XOR2X1   g4043(.A(CRC_OUT_3_31), .B(WX8635), .Y(n9806));
XOR2X1   g4044(.A(n9806), .B(CRC_OUT_3_10), .Y(n9807));
NOR2X1   g4045(.A(n9807), .B(n5827), .Y(CRC_OUT_3_11));
XOR2X1   g4046(.A(CRC_OUT_3_11), .B(WX8633), .Y(n9809));
NOR2X1   g4047(.A(n9809), .B(n5827), .Y(CRC_OUT_3_12));
XOR2X1   g4048(.A(CRC_OUT_3_12), .B(WX8631), .Y(n9811));
NOR2X1   g4049(.A(n9811), .B(n5827), .Y(CRC_OUT_3_13));
XOR2X1   g4050(.A(CRC_OUT_3_13), .B(WX8629), .Y(n9813));
NOR2X1   g4051(.A(n9813), .B(n5827), .Y(CRC_OUT_3_14));
XOR2X1   g4052(.A(CRC_OUT_3_14), .B(WX8627), .Y(n9815));
NOR2X1   g4053(.A(n9815), .B(n5827), .Y(CRC_OUT_3_15));
XOR2X1   g4054(.A(CRC_OUT_3_31), .B(WX8625), .Y(n9817));
XOR2X1   g4055(.A(n9817), .B(CRC_OUT_3_15), .Y(n9818));
NOR2X1   g4056(.A(n9818), .B(n5827), .Y(CRC_OUT_3_16));
XOR2X1   g4057(.A(CRC_OUT_3_16), .B(WX8623), .Y(n9820));
NOR2X1   g4058(.A(n9820), .B(n5827), .Y(CRC_OUT_3_17));
XOR2X1   g4059(.A(CRC_OUT_3_17), .B(WX8621), .Y(n9822));
NOR2X1   g4060(.A(n9822), .B(n5827), .Y(CRC_OUT_3_18));
XOR2X1   g4061(.A(CRC_OUT_3_18), .B(WX8619), .Y(n9824));
NOR2X1   g4062(.A(n9824), .B(n5827), .Y(CRC_OUT_3_19));
XOR2X1   g4063(.A(CRC_OUT_3_19), .B(WX8617), .Y(n9826));
NOR2X1   g4064(.A(n9826), .B(n5827), .Y(CRC_OUT_3_20));
XOR2X1   g4065(.A(CRC_OUT_3_20), .B(WX8615), .Y(n9828));
NOR2X1   g4066(.A(n9828), .B(n5827), .Y(CRC_OUT_3_21));
XOR2X1   g4067(.A(CRC_OUT_3_21), .B(WX8613), .Y(n9830));
NOR2X1   g4068(.A(n9830), .B(n5827), .Y(CRC_OUT_3_22));
XOR2X1   g4069(.A(CRC_OUT_3_22), .B(WX8611), .Y(n9832));
NOR2X1   g4070(.A(n9832), .B(n5827), .Y(CRC_OUT_3_23));
XOR2X1   g4071(.A(CRC_OUT_3_23), .B(WX8609), .Y(n9834));
NOR2X1   g4072(.A(n9834), .B(n5827), .Y(CRC_OUT_3_24));
XOR2X1   g4073(.A(CRC_OUT_3_24), .B(WX8607), .Y(n9836));
NOR2X1   g4074(.A(n9836), .B(n5827), .Y(CRC_OUT_3_25));
XOR2X1   g4075(.A(CRC_OUT_3_25), .B(WX8605), .Y(n9838));
NOR2X1   g4076(.A(n9838), .B(n5827), .Y(CRC_OUT_3_26));
XOR2X1   g4077(.A(CRC_OUT_3_26), .B(WX8603), .Y(n9840));
NOR2X1   g4078(.A(n9840), .B(n5827), .Y(CRC_OUT_3_27));
XOR2X1   g4079(.A(CRC_OUT_3_27), .B(WX8601), .Y(n9842));
NOR2X1   g4080(.A(n9842), .B(n5827), .Y(CRC_OUT_3_28));
XOR2X1   g4081(.A(CRC_OUT_3_28), .B(WX8599), .Y(n9844));
NOR2X1   g4082(.A(n9844), .B(n5827), .Y(CRC_OUT_3_29));
XOR2X1   g4083(.A(CRC_OUT_3_29), .B(WX8597), .Y(n9846));
NOR2X1   g4084(.A(n9846), .B(n5827), .Y(CRC_OUT_3_30));
XOR2X1   g4085(.A(CRC_OUT_3_30), .B(WX8595), .Y(n9848));
NOR2X1   g4086(.A(n9848), .B(n5827), .Y(CRC_OUT_3_31));
AND2X1   g4087(.A(WX9538), .B(RESET), .Y(n7207));
AND2X1   g4088(.A(WX9540), .B(RESET), .Y(n7212));
AND2X1   g4089(.A(WX9542), .B(RESET), .Y(n7217));
AND2X1   g4090(.A(WX9544), .B(RESET), .Y(n7222));
AND2X1   g4091(.A(WX9546), .B(RESET), .Y(n7227));
AND2X1   g4092(.A(WX9548), .B(RESET), .Y(n7232));
AND2X1   g4093(.A(WX9550), .B(RESET), .Y(n7237));
AND2X1   g4094(.A(WX9552), .B(RESET), .Y(n7242));
AND2X1   g4095(.A(WX9554), .B(RESET), .Y(n7247));
AND2X1   g4096(.A(WX9556), .B(RESET), .Y(n7252));
AND2X1   g4097(.A(WX9558), .B(RESET), .Y(n7257));
AND2X1   g4098(.A(WX9560), .B(RESET), .Y(n7262));
AND2X1   g4099(.A(WX9562), .B(RESET), .Y(n7267));
AND2X1   g4100(.A(WX9564), .B(RESET), .Y(n7272));
AND2X1   g4101(.A(WX9566), .B(RESET), .Y(n7277));
AND2X1   g4102(.A(WX9568), .B(RESET), .Y(n7282));
AND2X1   g4103(.A(WX9570), .B(RESET), .Y(n7287));
AND2X1   g4104(.A(WX9572), .B(RESET), .Y(n7292));
AND2X1   g4105(.A(WX9574), .B(RESET), .Y(n7297));
AND2X1   g4106(.A(WX9576), .B(RESET), .Y(n7302));
AND2X1   g4107(.A(WX9578), .B(RESET), .Y(n7307));
AND2X1   g4108(.A(WX9580), .B(RESET), .Y(n7312));
AND2X1   g4109(.A(WX9582), .B(RESET), .Y(n7317));
AND2X1   g4110(.A(WX9584), .B(RESET), .Y(n7322));
AND2X1   g4111(.A(WX9586), .B(RESET), .Y(n7327));
AND2X1   g4112(.A(WX9588), .B(RESET), .Y(n7332));
AND2X1   g4113(.A(WX9590), .B(RESET), .Y(n7337));
AND2X1   g4114(.A(WX9592), .B(RESET), .Y(n7342));
AND2X1   g4115(.A(WX9594), .B(RESET), .Y(n7347));
AND2X1   g4116(.A(WX9596), .B(RESET), .Y(n7352));
AND2X1   g4117(.A(WX9598), .B(RESET), .Y(n7357));
NOR2X1   g4118(.A(WX9536), .B(n5827), .Y(n7362));
INVX1    g4119(.A(CRC_OUT_2_31), .Y(n9882));
XOR2X1   g4120(.A(WX10989), .B(TM1), .Y(n9883));
XOR2X1   g4121(.A(n9883), .B(WX11053), .Y(n9884));
INVX1    g4122(.A(WX11117), .Y(n9885));
XOR2X1   g4123(.A(WX11181), .B(n9885), .Y(n9886));
XOR2X1   g4124(.A(n9886), .B(n9884), .Y(n9887));
MX2X1    g4125(.A(n9882), .B(n9887), .S0(n5539), .Y(n9889));
INVX1    g4126(.A(WX9536), .Y(n9890));
MX2X1    g4127(.A(n9890), .B(n9308), .S0(n5539), .Y(n9891));
MX2X1    g4128(.A(n9889), .B(n9891), .S0(TM1), .Y(n9892));
NOR2X1   g4129(.A(n9892), .B(n5827), .Y(n7367));
INVX1    g4130(.A(CRC_OUT_2_30), .Y(n9894));
XOR2X1   g4131(.A(WX10991), .B(TM1), .Y(n9895));
XOR2X1   g4132(.A(n9895), .B(WX11055), .Y(n9896));
INVX1    g4133(.A(WX11119), .Y(n9897));
XOR2X1   g4134(.A(WX11183), .B(n9897), .Y(n9898));
XOR2X1   g4135(.A(n9898), .B(n9896), .Y(n9899));
MX2X1    g4136(.A(n9894), .B(n9899), .S0(n5539), .Y(n9901));
INVX1    g4137(.A(WX9538), .Y(n9902));
MX2X1    g4138(.A(n9902), .B(n9320), .S0(n5539), .Y(n9903));
MX2X1    g4139(.A(n9901), .B(n9903), .S0(TM1), .Y(n9904));
NOR2X1   g4140(.A(n9904), .B(n5827), .Y(n7372));
INVX1    g4141(.A(CRC_OUT_2_29), .Y(n9906));
XOR2X1   g4142(.A(WX10993), .B(TM1), .Y(n9907));
XOR2X1   g4143(.A(n9907), .B(WX11057), .Y(n9908));
INVX1    g4144(.A(WX11121), .Y(n9909));
XOR2X1   g4145(.A(WX11185), .B(n9909), .Y(n9910));
XOR2X1   g4146(.A(n9910), .B(n9908), .Y(n9911));
MX2X1    g4147(.A(n9906), .B(n9911), .S0(n5539), .Y(n9913));
INVX1    g4148(.A(WX9540), .Y(n9914));
MX2X1    g4149(.A(n9914), .B(n9332), .S0(n5539), .Y(n9915));
MX2X1    g4150(.A(n9913), .B(n9915), .S0(TM1), .Y(n9916));
NOR2X1   g4151(.A(n9916), .B(n5827), .Y(n7377));
INVX1    g4152(.A(CRC_OUT_2_28), .Y(n9918));
XOR2X1   g4153(.A(WX10995), .B(TM1), .Y(n9919));
XOR2X1   g4154(.A(n9919), .B(WX11059), .Y(n9920));
INVX1    g4155(.A(WX11123), .Y(n9921));
XOR2X1   g4156(.A(WX11187), .B(n9921), .Y(n9922));
XOR2X1   g4157(.A(n9922), .B(n9920), .Y(n9923));
MX2X1    g4158(.A(n9918), .B(n9923), .S0(n5539), .Y(n9925));
INVX1    g4159(.A(WX9542), .Y(n9926));
MX2X1    g4160(.A(n9926), .B(n9344), .S0(n5539), .Y(n9927));
MX2X1    g4161(.A(n9925), .B(n9927), .S0(TM1), .Y(n9928));
NOR2X1   g4162(.A(n9928), .B(n5827), .Y(n7382));
INVX1    g4163(.A(CRC_OUT_2_27), .Y(n9930));
XOR2X1   g4164(.A(WX10997), .B(TM1), .Y(n9931));
XOR2X1   g4165(.A(n9931), .B(WX11061), .Y(n9932));
INVX1    g4166(.A(WX11125), .Y(n9933));
XOR2X1   g4167(.A(WX11189), .B(n9933), .Y(n9934));
XOR2X1   g4168(.A(n9934), .B(n9932), .Y(n9935));
MX2X1    g4169(.A(n9930), .B(n9935), .S0(n5539), .Y(n9937));
INVX1    g4170(.A(WX9544), .Y(n9938));
MX2X1    g4171(.A(n9938), .B(n9356), .S0(n5539), .Y(n9939));
MX2X1    g4172(.A(n9937), .B(n9939), .S0(TM1), .Y(n9940));
NOR2X1   g4173(.A(n9940), .B(n5827), .Y(n7387));
INVX1    g4174(.A(CRC_OUT_2_26), .Y(n9942));
XOR2X1   g4175(.A(WX10999), .B(TM1), .Y(n9943));
XOR2X1   g4176(.A(n9943), .B(WX11063), .Y(n9944));
INVX1    g4177(.A(WX11127), .Y(n9945));
XOR2X1   g4178(.A(WX11191), .B(n9945), .Y(n9946));
XOR2X1   g4179(.A(n9946), .B(n9944), .Y(n9947));
MX2X1    g4180(.A(n9942), .B(n9947), .S0(n5539), .Y(n9949));
INVX1    g4181(.A(WX9546), .Y(n9950));
MX2X1    g4182(.A(n9950), .B(n9368), .S0(n5539), .Y(n9951));
MX2X1    g4183(.A(n9949), .B(n9951), .S0(TM1), .Y(n9952));
NOR2X1   g4184(.A(n9952), .B(n5827), .Y(n7392));
INVX1    g4185(.A(CRC_OUT_2_25), .Y(n9954));
XOR2X1   g4186(.A(WX11001), .B(TM1), .Y(n9955));
XOR2X1   g4187(.A(n9955), .B(WX11065), .Y(n9956));
INVX1    g4188(.A(WX11129), .Y(n9957));
XOR2X1   g4189(.A(WX11193), .B(n9957), .Y(n9958));
XOR2X1   g4190(.A(n9958), .B(n9956), .Y(n9959));
MX2X1    g4191(.A(n9954), .B(n9959), .S0(n5539), .Y(n9961));
INVX1    g4192(.A(WX9548), .Y(n9962));
MX2X1    g4193(.A(n9962), .B(n9380), .S0(n5539), .Y(n9963));
MX2X1    g4194(.A(n9961), .B(n9963), .S0(TM1), .Y(n9964));
NOR2X1   g4195(.A(n9964), .B(n5827), .Y(n7397));
INVX1    g4196(.A(CRC_OUT_2_24), .Y(n9966));
XOR2X1   g4197(.A(WX11003), .B(TM1), .Y(n9967));
XOR2X1   g4198(.A(n9967), .B(WX11067), .Y(n9968));
INVX1    g4199(.A(WX11131), .Y(n9969));
XOR2X1   g4200(.A(WX11195), .B(n9969), .Y(n9970));
XOR2X1   g4201(.A(n9970), .B(n9968), .Y(n9971));
MX2X1    g4202(.A(n9966), .B(n9971), .S0(n5539), .Y(n9973));
INVX1    g4203(.A(WX9550), .Y(n9974));
MX2X1    g4204(.A(n9974), .B(n9392), .S0(n5539), .Y(n9975));
MX2X1    g4205(.A(n9973), .B(n9975), .S0(TM1), .Y(n9976));
NOR2X1   g4206(.A(n9976), .B(n5827), .Y(n7402));
INVX1    g4207(.A(CRC_OUT_2_23), .Y(n9978));
XOR2X1   g4208(.A(WX11005), .B(TM1), .Y(n9979));
XOR2X1   g4209(.A(n9979), .B(WX11069), .Y(n9980));
INVX1    g4210(.A(WX11133), .Y(n9981));
XOR2X1   g4211(.A(WX11197), .B(n9981), .Y(n9982));
XOR2X1   g4212(.A(n9982), .B(n9980), .Y(n9983));
MX2X1    g4213(.A(n9978), .B(n9983), .S0(n5539), .Y(n9985));
INVX1    g4214(.A(WX9552), .Y(n9986));
MX2X1    g4215(.A(n9986), .B(n9404), .S0(n5539), .Y(n9987));
MX2X1    g4216(.A(n9985), .B(n9987), .S0(TM1), .Y(n9988));
NOR2X1   g4217(.A(n9988), .B(n5827), .Y(n7407));
INVX1    g4218(.A(CRC_OUT_2_22), .Y(n9990));
XOR2X1   g4219(.A(WX11007), .B(TM1), .Y(n9991));
XOR2X1   g4220(.A(n9991), .B(WX11071), .Y(n9992));
INVX1    g4221(.A(WX11135), .Y(n9993));
XOR2X1   g4222(.A(WX11199), .B(n9993), .Y(n9994));
XOR2X1   g4223(.A(n9994), .B(n9992), .Y(n9995));
MX2X1    g4224(.A(n9990), .B(n9995), .S0(n5539), .Y(n9997));
INVX1    g4225(.A(WX9554), .Y(n9998));
MX2X1    g4226(.A(n9998), .B(n9416), .S0(n5539), .Y(n9999));
MX2X1    g4227(.A(n9997), .B(n9999), .S0(TM1), .Y(n10000));
NOR2X1   g4228(.A(n10000), .B(n5827), .Y(n7412));
INVX1    g4229(.A(CRC_OUT_2_21), .Y(n10002));
XOR2X1   g4230(.A(WX11009), .B(TM1), .Y(n10003));
XOR2X1   g4231(.A(n10003), .B(WX11073), .Y(n10004));
INVX1    g4232(.A(WX11137), .Y(n10005));
XOR2X1   g4233(.A(WX11201), .B(n10005), .Y(n10006));
XOR2X1   g4234(.A(n10006), .B(n10004), .Y(n10007));
MX2X1    g4235(.A(n10002), .B(n10007), .S0(n5539), .Y(n10009));
INVX1    g4236(.A(WX9556), .Y(n10010));
MX2X1    g4237(.A(n10010), .B(n9428), .S0(n5539), .Y(n10011));
MX2X1    g4238(.A(n10009), .B(n10011), .S0(TM1), .Y(n10012));
NOR2X1   g4239(.A(n10012), .B(n5827), .Y(n7417));
INVX1    g4240(.A(CRC_OUT_2_20), .Y(n10014));
XOR2X1   g4241(.A(WX11011), .B(TM1), .Y(n10015));
XOR2X1   g4242(.A(n10015), .B(WX11075), .Y(n10016));
INVX1    g4243(.A(WX11139), .Y(n10017));
XOR2X1   g4244(.A(WX11203), .B(n10017), .Y(n10018));
XOR2X1   g4245(.A(n10018), .B(n10016), .Y(n10019));
MX2X1    g4246(.A(n10014), .B(n10019), .S0(n5539), .Y(n10021));
INVX1    g4247(.A(WX9558), .Y(n10022));
MX2X1    g4248(.A(n10022), .B(n9440), .S0(n5539), .Y(n10023));
MX2X1    g4249(.A(n10021), .B(n10023), .S0(TM1), .Y(n10024));
NOR2X1   g4250(.A(n10024), .B(n5827), .Y(n7422));
INVX1    g4251(.A(CRC_OUT_2_19), .Y(n10026));
XOR2X1   g4252(.A(WX11013), .B(TM1), .Y(n10027));
XOR2X1   g4253(.A(n10027), .B(WX11077), .Y(n10028));
INVX1    g4254(.A(WX11141), .Y(n10029));
XOR2X1   g4255(.A(WX11205), .B(n10029), .Y(n10030));
XOR2X1   g4256(.A(n10030), .B(n10028), .Y(n10031));
MX2X1    g4257(.A(n10026), .B(n10031), .S0(n5539), .Y(n10033));
INVX1    g4258(.A(WX9560), .Y(n10034));
MX2X1    g4259(.A(n10034), .B(n9452), .S0(n5539), .Y(n10035));
MX2X1    g4260(.A(n10033), .B(n10035), .S0(TM1), .Y(n10036));
NOR2X1   g4261(.A(n10036), .B(n5827), .Y(n7427));
INVX1    g4262(.A(CRC_OUT_2_18), .Y(n10038));
XOR2X1   g4263(.A(WX11015), .B(TM1), .Y(n10039));
XOR2X1   g4264(.A(n10039), .B(WX11079), .Y(n10040));
INVX1    g4265(.A(WX11143), .Y(n10041));
XOR2X1   g4266(.A(WX11207), .B(n10041), .Y(n10042));
XOR2X1   g4267(.A(n10042), .B(n10040), .Y(n10043));
MX2X1    g4268(.A(n10038), .B(n10043), .S0(n5539), .Y(n10045));
INVX1    g4269(.A(WX9562), .Y(n10046));
MX2X1    g4270(.A(n10046), .B(n9464), .S0(n5539), .Y(n10047));
MX2X1    g4271(.A(n10045), .B(n10047), .S0(TM1), .Y(n10048));
NOR2X1   g4272(.A(n10048), .B(n5827), .Y(n7432));
INVX1    g4273(.A(CRC_OUT_2_17), .Y(n10050));
XOR2X1   g4274(.A(WX11017), .B(TM1), .Y(n10051));
XOR2X1   g4275(.A(n10051), .B(WX11081), .Y(n10052));
INVX1    g4276(.A(WX11145), .Y(n10053));
XOR2X1   g4277(.A(WX11209), .B(n10053), .Y(n10054));
XOR2X1   g4278(.A(n10054), .B(n10052), .Y(n10055));
MX2X1    g4279(.A(n10050), .B(n10055), .S0(n5539), .Y(n10057));
INVX1    g4280(.A(WX9564), .Y(n10058));
MX2X1    g4281(.A(n10058), .B(n9476), .S0(n5539), .Y(n10059));
MX2X1    g4282(.A(n10057), .B(n10059), .S0(TM1), .Y(n10060));
NOR2X1   g4283(.A(n10060), .B(n5827), .Y(n7437));
INVX1    g4284(.A(CRC_OUT_2_16), .Y(n10062));
XOR2X1   g4285(.A(WX11019), .B(TM1), .Y(n10063));
XOR2X1   g4286(.A(n10063), .B(WX11083), .Y(n10064));
INVX1    g4287(.A(WX11147), .Y(n10065));
XOR2X1   g4288(.A(WX11211), .B(n10065), .Y(n10066));
XOR2X1   g4289(.A(n10066), .B(n10064), .Y(n10067));
MX2X1    g4290(.A(n10062), .B(n10067), .S0(n5539), .Y(n10069));
INVX1    g4291(.A(WX9566), .Y(n10070));
MX2X1    g4292(.A(n10070), .B(n9488), .S0(n5539), .Y(n10071));
MX2X1    g4293(.A(n10069), .B(n10071), .S0(TM1), .Y(n10072));
NOR2X1   g4294(.A(n10072), .B(n5827), .Y(n7442));
INVX1    g4295(.A(CRC_OUT_2_15), .Y(n10074));
XOR2X1   g4296(.A(WX11021), .B(TM0), .Y(n10075));
XOR2X1   g4297(.A(n10075), .B(WX11085), .Y(n10076));
INVX1    g4298(.A(WX11149), .Y(n10077));
XOR2X1   g4299(.A(WX11213), .B(n10077), .Y(n10078));
XOR2X1   g4300(.A(n10078), .B(n10076), .Y(n10079));
MX2X1    g4301(.A(n10074), .B(n10079), .S0(n5539), .Y(n10081));
INVX1    g4302(.A(WX9568), .Y(n10082));
MX2X1    g4303(.A(n10082), .B(n9500), .S0(n5539), .Y(n10083));
MX2X1    g4304(.A(n10081), .B(n10083), .S0(TM1), .Y(n10084));
NOR2X1   g4305(.A(n10084), .B(n5827), .Y(n7447));
INVX1    g4306(.A(CRC_OUT_2_14), .Y(n10086));
XOR2X1   g4307(.A(WX11023), .B(TM0), .Y(n10087));
XOR2X1   g4308(.A(n10087), .B(WX11087), .Y(n10088));
INVX1    g4309(.A(WX11151), .Y(n10089));
XOR2X1   g4310(.A(WX11215), .B(n10089), .Y(n10090));
XOR2X1   g4311(.A(n10090), .B(n10088), .Y(n10091));
MX2X1    g4312(.A(n10086), .B(n10091), .S0(n5539), .Y(n10093));
INVX1    g4313(.A(WX9570), .Y(n10094));
MX2X1    g4314(.A(n10094), .B(n9512), .S0(n5539), .Y(n10095));
MX2X1    g4315(.A(n10093), .B(n10095), .S0(TM1), .Y(n10096));
NOR2X1   g4316(.A(n10096), .B(n5827), .Y(n7452));
INVX1    g4317(.A(CRC_OUT_2_13), .Y(n10098));
XOR2X1   g4318(.A(WX11025), .B(TM0), .Y(n10099));
XOR2X1   g4319(.A(n10099), .B(WX11089), .Y(n10100));
INVX1    g4320(.A(WX11153), .Y(n10101));
XOR2X1   g4321(.A(WX11217), .B(n10101), .Y(n10102));
XOR2X1   g4322(.A(n10102), .B(n10100), .Y(n10103));
MX2X1    g4323(.A(n10098), .B(n10103), .S0(n5539), .Y(n10105));
INVX1    g4324(.A(WX9572), .Y(n10106));
MX2X1    g4325(.A(n10106), .B(n9524), .S0(n5539), .Y(n10107));
MX2X1    g4326(.A(n10105), .B(n10107), .S0(TM1), .Y(n10108));
NOR2X1   g4327(.A(n10108), .B(n5827), .Y(n7457));
INVX1    g4328(.A(CRC_OUT_2_12), .Y(n10110));
XOR2X1   g4329(.A(WX11027), .B(TM0), .Y(n10111));
XOR2X1   g4330(.A(n10111), .B(WX11091), .Y(n10112));
INVX1    g4331(.A(WX11155), .Y(n10113));
XOR2X1   g4332(.A(WX11219), .B(n10113), .Y(n10114));
XOR2X1   g4333(.A(n10114), .B(n10112), .Y(n10115));
MX2X1    g4334(.A(n10110), .B(n10115), .S0(n5539), .Y(n10117));
INVX1    g4335(.A(WX9574), .Y(n10118));
MX2X1    g4336(.A(n10118), .B(n9536), .S0(n5539), .Y(n10119));
MX2X1    g4337(.A(n10117), .B(n10119), .S0(TM1), .Y(n10120));
NOR2X1   g4338(.A(n10120), .B(n5827), .Y(n7462));
INVX1    g4339(.A(CRC_OUT_2_11), .Y(n10122));
XOR2X1   g4340(.A(WX11029), .B(TM0), .Y(n10123));
XOR2X1   g4341(.A(n10123), .B(WX11093), .Y(n10124));
INVX1    g4342(.A(WX11157), .Y(n10125));
XOR2X1   g4343(.A(WX11221), .B(n10125), .Y(n10126));
XOR2X1   g4344(.A(n10126), .B(n10124), .Y(n10127));
MX2X1    g4345(.A(n10122), .B(n10127), .S0(n5539), .Y(n10129));
INVX1    g4346(.A(WX9576), .Y(n10130));
MX2X1    g4347(.A(n10130), .B(n9548), .S0(n5539), .Y(n10131));
MX2X1    g4348(.A(n10129), .B(n10131), .S0(TM1), .Y(n10132));
NOR2X1   g4349(.A(n10132), .B(n5827), .Y(n7467));
INVX1    g4350(.A(CRC_OUT_2_10), .Y(n10134));
XOR2X1   g4351(.A(WX11031), .B(TM0), .Y(n10135));
XOR2X1   g4352(.A(n10135), .B(WX11095), .Y(n10136));
INVX1    g4353(.A(WX11159), .Y(n10137));
XOR2X1   g4354(.A(WX11223), .B(n10137), .Y(n10138));
XOR2X1   g4355(.A(n10138), .B(n10136), .Y(n10139));
MX2X1    g4356(.A(n10134), .B(n10139), .S0(n5539), .Y(n10141));
INVX1    g4357(.A(WX9578), .Y(n10142));
MX2X1    g4358(.A(n10142), .B(n9560), .S0(n5539), .Y(n10143));
MX2X1    g4359(.A(n10141), .B(n10143), .S0(TM1), .Y(n10144));
NOR2X1   g4360(.A(n10144), .B(n5827), .Y(n7472));
INVX1    g4361(.A(CRC_OUT_2_9), .Y(n10146));
XOR2X1   g4362(.A(WX11033), .B(TM0), .Y(n10147));
XOR2X1   g4363(.A(n10147), .B(WX11097), .Y(n10148));
INVX1    g4364(.A(WX11161), .Y(n10149));
XOR2X1   g4365(.A(WX11225), .B(n10149), .Y(n10150));
XOR2X1   g4366(.A(n10150), .B(n10148), .Y(n10151));
MX2X1    g4367(.A(n10146), .B(n10151), .S0(n5539), .Y(n10153));
INVX1    g4368(.A(WX9580), .Y(n10154));
MX2X1    g4369(.A(n10154), .B(n9572), .S0(n5539), .Y(n10155));
MX2X1    g4370(.A(n10153), .B(n10155), .S0(TM1), .Y(n10156));
NOR2X1   g4371(.A(n10156), .B(n5827), .Y(n7477));
INVX1    g4372(.A(CRC_OUT_2_8), .Y(n10158));
XOR2X1   g4373(.A(WX11035), .B(TM0), .Y(n10159));
XOR2X1   g4374(.A(n10159), .B(WX11099), .Y(n10160));
INVX1    g4375(.A(WX11163), .Y(n10161));
XOR2X1   g4376(.A(WX11227), .B(n10161), .Y(n10162));
XOR2X1   g4377(.A(n10162), .B(n10160), .Y(n10163));
MX2X1    g4378(.A(n10158), .B(n10163), .S0(n5539), .Y(n10165));
INVX1    g4379(.A(WX9582), .Y(n10166));
MX2X1    g4380(.A(n10166), .B(n9584), .S0(n5539), .Y(n10167));
MX2X1    g4381(.A(n10165), .B(n10167), .S0(TM1), .Y(n10168));
NOR2X1   g4382(.A(n10168), .B(n5827), .Y(n7482));
INVX1    g4383(.A(CRC_OUT_2_7), .Y(n10170));
XOR2X1   g4384(.A(WX11037), .B(TM0), .Y(n10171));
XOR2X1   g4385(.A(n10171), .B(WX11101), .Y(n10172));
INVX1    g4386(.A(WX11165), .Y(n10173));
XOR2X1   g4387(.A(WX11229), .B(n10173), .Y(n10174));
XOR2X1   g4388(.A(n10174), .B(n10172), .Y(n10175));
MX2X1    g4389(.A(n10170), .B(n10175), .S0(n5539), .Y(n10177));
INVX1    g4390(.A(WX9584), .Y(n10178));
MX2X1    g4391(.A(n10178), .B(n9596), .S0(n5539), .Y(n10179));
MX2X1    g4392(.A(n10177), .B(n10179), .S0(TM1), .Y(n10180));
NOR2X1   g4393(.A(n10180), .B(n5827), .Y(n7487));
INVX1    g4394(.A(CRC_OUT_2_6), .Y(n10182));
XOR2X1   g4395(.A(WX11039), .B(TM0), .Y(n10183));
XOR2X1   g4396(.A(n10183), .B(WX11103), .Y(n10184));
INVX1    g4397(.A(WX11167), .Y(n10185));
XOR2X1   g4398(.A(WX11231), .B(n10185), .Y(n10186));
XOR2X1   g4399(.A(n10186), .B(n10184), .Y(n10187));
MX2X1    g4400(.A(n10182), .B(n10187), .S0(n5539), .Y(n10189));
INVX1    g4401(.A(WX9586), .Y(n10190));
MX2X1    g4402(.A(n10190), .B(n9608), .S0(n5539), .Y(n10191));
MX2X1    g4403(.A(n10189), .B(n10191), .S0(TM1), .Y(n10192));
NOR2X1   g4404(.A(n10192), .B(n5827), .Y(n7492));
INVX1    g4405(.A(CRC_OUT_2_5), .Y(n10194));
XOR2X1   g4406(.A(WX11041), .B(TM0), .Y(n10195));
XOR2X1   g4407(.A(n10195), .B(WX11105), .Y(n10196));
INVX1    g4408(.A(WX11169), .Y(n10197));
XOR2X1   g4409(.A(WX11233), .B(n10197), .Y(n10198));
XOR2X1   g4410(.A(n10198), .B(n10196), .Y(n10199));
MX2X1    g4411(.A(n10194), .B(n10199), .S0(n5539), .Y(n10201));
INVX1    g4412(.A(WX9588), .Y(n10202));
MX2X1    g4413(.A(n10202), .B(n9620), .S0(n5539), .Y(n10203));
MX2X1    g4414(.A(n10201), .B(n10203), .S0(TM1), .Y(n10204));
NOR2X1   g4415(.A(n10204), .B(n5827), .Y(n7497));
INVX1    g4416(.A(CRC_OUT_2_4), .Y(n10206));
XOR2X1   g4417(.A(WX11043), .B(TM0), .Y(n10207));
XOR2X1   g4418(.A(n10207), .B(WX11107), .Y(n10208));
INVX1    g4419(.A(WX11171), .Y(n10209));
XOR2X1   g4420(.A(WX11235), .B(n10209), .Y(n10210));
XOR2X1   g4421(.A(n10210), .B(n10208), .Y(n10211));
MX2X1    g4422(.A(n10206), .B(n10211), .S0(n5539), .Y(n10213));
INVX1    g4423(.A(WX9590), .Y(n10214));
MX2X1    g4424(.A(n10214), .B(n9632), .S0(n5539), .Y(n10215));
MX2X1    g4425(.A(n10213), .B(n10215), .S0(TM1), .Y(n10216));
NOR2X1   g4426(.A(n10216), .B(n5827), .Y(n7502));
INVX1    g4427(.A(CRC_OUT_2_3), .Y(n10218));
XOR2X1   g4428(.A(WX11045), .B(TM0), .Y(n10219));
XOR2X1   g4429(.A(n10219), .B(WX11109), .Y(n10220));
INVX1    g4430(.A(WX11173), .Y(n10221));
XOR2X1   g4431(.A(WX11237), .B(n10221), .Y(n10222));
XOR2X1   g4432(.A(n10222), .B(n10220), .Y(n10223));
MX2X1    g4433(.A(n10218), .B(n10223), .S0(n5539), .Y(n10225));
INVX1    g4434(.A(WX9592), .Y(n10226));
MX2X1    g4435(.A(n10226), .B(n9644), .S0(n5539), .Y(n10227));
MX2X1    g4436(.A(n10225), .B(n10227), .S0(TM1), .Y(n10228));
NOR2X1   g4437(.A(n10228), .B(n5827), .Y(n7507));
INVX1    g4438(.A(CRC_OUT_2_2), .Y(n10230));
XOR2X1   g4439(.A(WX11047), .B(TM0), .Y(n10231));
XOR2X1   g4440(.A(n10231), .B(WX11111), .Y(n10232));
INVX1    g4441(.A(WX11175), .Y(n10233));
XOR2X1   g4442(.A(WX11239), .B(n10233), .Y(n10234));
XOR2X1   g4443(.A(n10234), .B(n10232), .Y(n10235));
MX2X1    g4444(.A(n10230), .B(n10235), .S0(n5539), .Y(n10237));
INVX1    g4445(.A(WX9594), .Y(n10238));
MX2X1    g4446(.A(n10238), .B(n9656), .S0(n5539), .Y(n10239));
MX2X1    g4447(.A(n10237), .B(n10239), .S0(TM1), .Y(n10240));
NOR2X1   g4448(.A(n10240), .B(n5827), .Y(n7512));
INVX1    g4449(.A(CRC_OUT_2_1), .Y(n10242));
XOR2X1   g4450(.A(WX11049), .B(TM0), .Y(n10243));
XOR2X1   g4451(.A(n10243), .B(WX11113), .Y(n10244));
INVX1    g4452(.A(WX11177), .Y(n10245));
XOR2X1   g4453(.A(WX11241), .B(n10245), .Y(n10246));
XOR2X1   g4454(.A(n10246), .B(n10244), .Y(n10247));
MX2X1    g4455(.A(n10242), .B(n10247), .S0(n5539), .Y(n10249));
INVX1    g4456(.A(WX9596), .Y(n10250));
MX2X1    g4457(.A(n10250), .B(n9668), .S0(n5539), .Y(n10251));
MX2X1    g4458(.A(n10249), .B(n10251), .S0(TM1), .Y(n10252));
NOR2X1   g4459(.A(n10252), .B(n5827), .Y(n7517));
INVX1    g4460(.A(CRC_OUT_2_0), .Y(n10254));
XOR2X1   g4461(.A(WX11051), .B(TM0), .Y(n10255));
XOR2X1   g4462(.A(n10255), .B(WX11115), .Y(n10256));
INVX1    g4463(.A(WX11179), .Y(n10257));
XOR2X1   g4464(.A(WX11243), .B(n10257), .Y(n10258));
XOR2X1   g4465(.A(n10258), .B(n10256), .Y(n10259));
MX2X1    g4466(.A(n10254), .B(n10259), .S0(n5539), .Y(n10261));
INVX1    g4467(.A(WX9598), .Y(n10262));
MX2X1    g4468(.A(n10262), .B(n9680), .S0(n5539), .Y(n10263));
MX2X1    g4469(.A(n10261), .B(n10263), .S0(TM1), .Y(n10264));
NOR2X1   g4470(.A(n10264), .B(n5827), .Y(n7522));
AND2X1   g4471(.A(WX9696), .B(RESET), .Y(n7527));
AND2X1   g4472(.A(WX9698), .B(RESET), .Y(n7532));
AND2X1   g4473(.A(WX9700), .B(RESET), .Y(n7537));
AND2X1   g4474(.A(WX9702), .B(RESET), .Y(n7542));
AND2X1   g4475(.A(WX9704), .B(RESET), .Y(n7547));
AND2X1   g4476(.A(WX9706), .B(RESET), .Y(n7552));
AND2X1   g4477(.A(WX9708), .B(RESET), .Y(n7557));
AND2X1   g4478(.A(WX9710), .B(RESET), .Y(n7562));
AND2X1   g4479(.A(WX9712), .B(RESET), .Y(n7567));
AND2X1   g4480(.A(WX9714), .B(RESET), .Y(n7572));
AND2X1   g4481(.A(WX9716), .B(RESET), .Y(n7577));
AND2X1   g4482(.A(WX9718), .B(RESET), .Y(n7582));
AND2X1   g4483(.A(WX9720), .B(RESET), .Y(n7587));
AND2X1   g4484(.A(WX9722), .B(RESET), .Y(n7592));
AND2X1   g4485(.A(WX9724), .B(RESET), .Y(n7597));
AND2X1   g4486(.A(WX9726), .B(RESET), .Y(n7602));
AND2X1   g4487(.A(WX9728), .B(RESET), .Y(n7607));
AND2X1   g4488(.A(WX9730), .B(RESET), .Y(n7612));
AND2X1   g4489(.A(WX9732), .B(RESET), .Y(n7617));
AND2X1   g4490(.A(WX9734), .B(RESET), .Y(n7622));
AND2X1   g4491(.A(WX9736), .B(RESET), .Y(n7627));
AND2X1   g4492(.A(WX9738), .B(RESET), .Y(n7632));
AND2X1   g4493(.A(WX9740), .B(RESET), .Y(n7637));
AND2X1   g4494(.A(WX9742), .B(RESET), .Y(n7642));
AND2X1   g4495(.A(WX9744), .B(RESET), .Y(n7647));
AND2X1   g4496(.A(WX9746), .B(RESET), .Y(n7652));
AND2X1   g4497(.A(WX9748), .B(RESET), .Y(n7657));
AND2X1   g4498(.A(WX9750), .B(RESET), .Y(n7662));
AND2X1   g4499(.A(WX9752), .B(RESET), .Y(n7667));
AND2X1   g4500(.A(WX9754), .B(RESET), .Y(n7672));
AND2X1   g4501(.A(WX9756), .B(RESET), .Y(n7677));
AND2X1   g4502(.A(WX9758), .B(RESET), .Y(n7682));
AND2X1   g4503(.A(WX9760), .B(RESET), .Y(n7687));
AND2X1   g4504(.A(WX9762), .B(RESET), .Y(n7692));
AND2X1   g4505(.A(WX9764), .B(RESET), .Y(n7697));
AND2X1   g4506(.A(WX9766), .B(RESET), .Y(n7702));
AND2X1   g4507(.A(WX9768), .B(RESET), .Y(n7707));
AND2X1   g4508(.A(WX9770), .B(RESET), .Y(n7712));
AND2X1   g4509(.A(WX9772), .B(RESET), .Y(n7717));
AND2X1   g4510(.A(WX9774), .B(RESET), .Y(n7722));
AND2X1   g4511(.A(WX9776), .B(RESET), .Y(n7727));
AND2X1   g4512(.A(WX9778), .B(RESET), .Y(n7732));
AND2X1   g4513(.A(WX9780), .B(RESET), .Y(n7737));
AND2X1   g4514(.A(WX9782), .B(RESET), .Y(n7742));
AND2X1   g4515(.A(WX9784), .B(RESET), .Y(n7747));
AND2X1   g4516(.A(WX9786), .B(RESET), .Y(n7752));
AND2X1   g4517(.A(WX9788), .B(RESET), .Y(n7757));
AND2X1   g4518(.A(WX9790), .B(RESET), .Y(n7762));
AND2X1   g4519(.A(WX9792), .B(RESET), .Y(n7767));
AND2X1   g4520(.A(WX9794), .B(RESET), .Y(n7772));
AND2X1   g4521(.A(WX9796), .B(RESET), .Y(n7777));
AND2X1   g4522(.A(WX9798), .B(RESET), .Y(n7782));
AND2X1   g4523(.A(WX9800), .B(RESET), .Y(n7787));
AND2X1   g4524(.A(WX9802), .B(RESET), .Y(n7792));
AND2X1   g4525(.A(WX9804), .B(RESET), .Y(n7797));
AND2X1   g4526(.A(WX9806), .B(RESET), .Y(n7802));
AND2X1   g4527(.A(WX9808), .B(RESET), .Y(n7807));
AND2X1   g4528(.A(WX9810), .B(RESET), .Y(n7812));
AND2X1   g4529(.A(WX9812), .B(RESET), .Y(n7817));
AND2X1   g4530(.A(WX9814), .B(RESET), .Y(n7822));
AND2X1   g4531(.A(WX9816), .B(RESET), .Y(n7827));
AND2X1   g4532(.A(WX9818), .B(RESET), .Y(n7832));
AND2X1   g4533(.A(WX9820), .B(RESET), .Y(n7837));
AND2X1   g4534(.A(WX9822), .B(RESET), .Y(n7842));
AND2X1   g4535(.A(WX9824), .B(RESET), .Y(n7847));
AND2X1   g4536(.A(WX9826), .B(RESET), .Y(n7852));
AND2X1   g4537(.A(WX9828), .B(RESET), .Y(n7857));
AND2X1   g4538(.A(WX9830), .B(RESET), .Y(n7862));
AND2X1   g4539(.A(WX9832), .B(RESET), .Y(n7867));
AND2X1   g4540(.A(WX9834), .B(RESET), .Y(n7872));
AND2X1   g4541(.A(WX9836), .B(RESET), .Y(n7877));
AND2X1   g4542(.A(WX9838), .B(RESET), .Y(n7882));
AND2X1   g4543(.A(WX9840), .B(RESET), .Y(n7887));
AND2X1   g4544(.A(WX9842), .B(RESET), .Y(n7892));
AND2X1   g4545(.A(WX9844), .B(RESET), .Y(n7897));
AND2X1   g4546(.A(WX9846), .B(RESET), .Y(n7902));
AND2X1   g4547(.A(WX9848), .B(RESET), .Y(n7907));
AND2X1   g4548(.A(WX9850), .B(RESET), .Y(n7912));
AND2X1   g4549(.A(WX9852), .B(RESET), .Y(n7917));
AND2X1   g4550(.A(WX9854), .B(RESET), .Y(n7922));
AND2X1   g4551(.A(WX9856), .B(RESET), .Y(n7927));
AND2X1   g4552(.A(WX9858), .B(RESET), .Y(n7932));
AND2X1   g4553(.A(WX9860), .B(RESET), .Y(n7937));
AND2X1   g4554(.A(WX9862), .B(RESET), .Y(n7942));
AND2X1   g4555(.A(WX9864), .B(RESET), .Y(n7947));
AND2X1   g4556(.A(WX9866), .B(RESET), .Y(n7952));
AND2X1   g4557(.A(WX9868), .B(RESET), .Y(n7957));
AND2X1   g4558(.A(WX9870), .B(RESET), .Y(n7962));
AND2X1   g4559(.A(WX9872), .B(RESET), .Y(n7967));
AND2X1   g4560(.A(WX9874), .B(RESET), .Y(n7972));
AND2X1   g4561(.A(WX9876), .B(RESET), .Y(n7977));
AND2X1   g4562(.A(WX9878), .B(RESET), .Y(n7982));
AND2X1   g4563(.A(WX9880), .B(RESET), .Y(n7987));
AND2X1   g4564(.A(WX9882), .B(RESET), .Y(n7992));
AND2X1   g4565(.A(WX9884), .B(RESET), .Y(n7997));
AND2X1   g4566(.A(WX9886), .B(RESET), .Y(n8002));
XOR2X1   g4567(.A(CRC_OUT_2_31), .B(WX9950), .Y(n10362));
NOR2X1   g4568(.A(n10362), .B(n5827), .Y(CRC_OUT_2_0));
XOR2X1   g4569(.A(CRC_OUT_2_0), .B(WX9948), .Y(n10364));
NOR2X1   g4570(.A(n10364), .B(n5827), .Y(CRC_OUT_2_1));
XOR2X1   g4571(.A(CRC_OUT_2_1), .B(WX9946), .Y(n10366));
NOR2X1   g4572(.A(n10366), .B(n5827), .Y(CRC_OUT_2_2));
XOR2X1   g4573(.A(CRC_OUT_2_2), .B(WX9944), .Y(n10368));
NOR2X1   g4574(.A(n10368), .B(n5827), .Y(CRC_OUT_2_3));
XOR2X1   g4575(.A(CRC_OUT_2_31), .B(WX9942), .Y(n10370));
XOR2X1   g4576(.A(n10370), .B(CRC_OUT_2_3), .Y(n10371));
NOR2X1   g4577(.A(n10371), .B(n5827), .Y(CRC_OUT_2_4));
XOR2X1   g4578(.A(CRC_OUT_2_4), .B(WX9940), .Y(n10373));
NOR2X1   g4579(.A(n10373), .B(n5827), .Y(CRC_OUT_2_5));
XOR2X1   g4580(.A(CRC_OUT_2_5), .B(WX9938), .Y(n10375));
NOR2X1   g4581(.A(n10375), .B(n5827), .Y(CRC_OUT_2_6));
XOR2X1   g4582(.A(CRC_OUT_2_6), .B(WX9936), .Y(n10377));
NOR2X1   g4583(.A(n10377), .B(n5827), .Y(CRC_OUT_2_7));
XOR2X1   g4584(.A(CRC_OUT_2_7), .B(WX9934), .Y(n10379));
NOR2X1   g4585(.A(n10379), .B(n5827), .Y(CRC_OUT_2_8));
XOR2X1   g4586(.A(CRC_OUT_2_8), .B(WX9932), .Y(n10381));
NOR2X1   g4587(.A(n10381), .B(n5827), .Y(CRC_OUT_2_9));
XOR2X1   g4588(.A(CRC_OUT_2_9), .B(WX9930), .Y(n10383));
NOR2X1   g4589(.A(n10383), .B(n5827), .Y(CRC_OUT_2_10));
XOR2X1   g4590(.A(CRC_OUT_2_31), .B(WX9928), .Y(n10385));
XOR2X1   g4591(.A(n10385), .B(CRC_OUT_2_10), .Y(n10386));
NOR2X1   g4592(.A(n10386), .B(n5827), .Y(CRC_OUT_2_11));
XOR2X1   g4593(.A(CRC_OUT_2_11), .B(WX9926), .Y(n10388));
NOR2X1   g4594(.A(n10388), .B(n5827), .Y(CRC_OUT_2_12));
XOR2X1   g4595(.A(CRC_OUT_2_12), .B(WX9924), .Y(n10390));
NOR2X1   g4596(.A(n10390), .B(n5827), .Y(CRC_OUT_2_13));
XOR2X1   g4597(.A(CRC_OUT_2_13), .B(WX9922), .Y(n10392));
NOR2X1   g4598(.A(n10392), .B(n5827), .Y(CRC_OUT_2_14));
XOR2X1   g4599(.A(CRC_OUT_2_14), .B(WX9920), .Y(n10394));
NOR2X1   g4600(.A(n10394), .B(n5827), .Y(CRC_OUT_2_15));
XOR2X1   g4601(.A(CRC_OUT_2_31), .B(WX9918), .Y(n10396));
XOR2X1   g4602(.A(n10396), .B(CRC_OUT_2_15), .Y(n10397));
NOR2X1   g4603(.A(n10397), .B(n5827), .Y(CRC_OUT_2_16));
XOR2X1   g4604(.A(CRC_OUT_2_16), .B(WX9916), .Y(n10399));
NOR2X1   g4605(.A(n10399), .B(n5827), .Y(CRC_OUT_2_17));
XOR2X1   g4606(.A(CRC_OUT_2_17), .B(WX9914), .Y(n10401));
NOR2X1   g4607(.A(n10401), .B(n5827), .Y(CRC_OUT_2_18));
XOR2X1   g4608(.A(CRC_OUT_2_18), .B(WX9912), .Y(n10403));
NOR2X1   g4609(.A(n10403), .B(n5827), .Y(CRC_OUT_2_19));
XOR2X1   g4610(.A(CRC_OUT_2_19), .B(WX9910), .Y(n10405));
NOR2X1   g4611(.A(n10405), .B(n5827), .Y(CRC_OUT_2_20));
XOR2X1   g4612(.A(CRC_OUT_2_20), .B(WX9908), .Y(n10407));
NOR2X1   g4613(.A(n10407), .B(n5827), .Y(CRC_OUT_2_21));
XOR2X1   g4614(.A(CRC_OUT_2_21), .B(WX9906), .Y(n10409));
NOR2X1   g4615(.A(n10409), .B(n5827), .Y(CRC_OUT_2_22));
XOR2X1   g4616(.A(CRC_OUT_2_22), .B(WX9904), .Y(n10411));
NOR2X1   g4617(.A(n10411), .B(n5827), .Y(CRC_OUT_2_23));
XOR2X1   g4618(.A(CRC_OUT_2_23), .B(WX9902), .Y(n10413));
NOR2X1   g4619(.A(n10413), .B(n5827), .Y(CRC_OUT_2_24));
XOR2X1   g4620(.A(CRC_OUT_2_24), .B(WX9900), .Y(n10415));
NOR2X1   g4621(.A(n10415), .B(n5827), .Y(CRC_OUT_2_25));
XOR2X1   g4622(.A(CRC_OUT_2_25), .B(WX9898), .Y(n10417));
NOR2X1   g4623(.A(n10417), .B(n5827), .Y(CRC_OUT_2_26));
XOR2X1   g4624(.A(CRC_OUT_2_26), .B(WX9896), .Y(n10419));
NOR2X1   g4625(.A(n10419), .B(n5827), .Y(CRC_OUT_2_27));
XOR2X1   g4626(.A(CRC_OUT_2_27), .B(WX9894), .Y(n10421));
NOR2X1   g4627(.A(n10421), .B(n5827), .Y(CRC_OUT_2_28));
XOR2X1   g4628(.A(CRC_OUT_2_28), .B(WX9892), .Y(n10423));
NOR2X1   g4629(.A(n10423), .B(n5827), .Y(CRC_OUT_2_29));
XOR2X1   g4630(.A(CRC_OUT_2_29), .B(WX9890), .Y(n10425));
NOR2X1   g4631(.A(n10425), .B(n5827), .Y(CRC_OUT_2_30));
XOR2X1   g4632(.A(CRC_OUT_2_30), .B(WX9888), .Y(n10427));
NOR2X1   g4633(.A(n10427), .B(n5827), .Y(CRC_OUT_2_31));
AND2X1   g4634(.A(WX10831), .B(RESET), .Y(n8135));
AND2X1   g4635(.A(WX10833), .B(RESET), .Y(n8140));
AND2X1   g4636(.A(WX10835), .B(RESET), .Y(n8145));
AND2X1   g4637(.A(WX10837), .B(RESET), .Y(n8150));
AND2X1   g4638(.A(WX10839), .B(RESET), .Y(n8155));
AND2X1   g4639(.A(WX10841), .B(RESET), .Y(n8160));
AND2X1   g4640(.A(WX10843), .B(RESET), .Y(n8165));
AND2X1   g4641(.A(WX10845), .B(RESET), .Y(n8170));
AND2X1   g4642(.A(WX10847), .B(RESET), .Y(n8175));
AND2X1   g4643(.A(WX10849), .B(RESET), .Y(n8180));
AND2X1   g4644(.A(WX10851), .B(RESET), .Y(n8185));
AND2X1   g4645(.A(WX10853), .B(RESET), .Y(n8190));
AND2X1   g4646(.A(WX10855), .B(RESET), .Y(n8195));
AND2X1   g4647(.A(WX10857), .B(RESET), .Y(n8200));
AND2X1   g4648(.A(WX10859), .B(RESET), .Y(n8205));
AND2X1   g4649(.A(WX10861), .B(RESET), .Y(n8210));
AND2X1   g4650(.A(WX10863), .B(RESET), .Y(n8215));
AND2X1   g4651(.A(WX10865), .B(RESET), .Y(n8220));
AND2X1   g4652(.A(WX10867), .B(RESET), .Y(n8225));
AND2X1   g4653(.A(WX10869), .B(RESET), .Y(n8230));
AND2X1   g4654(.A(WX10871), .B(RESET), .Y(n8235));
AND2X1   g4655(.A(WX10873), .B(RESET), .Y(n8240));
AND2X1   g4656(.A(WX10875), .B(RESET), .Y(n8245));
AND2X1   g4657(.A(WX10877), .B(RESET), .Y(n8250));
AND2X1   g4658(.A(WX10879), .B(RESET), .Y(n8255));
AND2X1   g4659(.A(WX10881), .B(RESET), .Y(n8260));
AND2X1   g4660(.A(WX10883), .B(RESET), .Y(n8265));
AND2X1   g4661(.A(WX10885), .B(RESET), .Y(n8270));
AND2X1   g4662(.A(WX10887), .B(RESET), .Y(n8275));
AND2X1   g4663(.A(WX10889), .B(RESET), .Y(n8280));
AND2X1   g4664(.A(WX10891), .B(RESET), .Y(n8285));
NOR2X1   g4665(.A(WX10829), .B(n5827), .Y(n8290));
AND2X1   g4666(.A(CRC_OUT_1_31), .B(TM0), .Y(n10461));
AOI21X1  g4667(.A0(n5539), .A1(DATA_0_31), .B0(n10461), .Y(n10462));
INVX1    g4668(.A(WX10829), .Y(n10463));
MX2X1    g4669(.A(n10463), .B(n9887), .S0(n5539), .Y(n10464));
MX2X1    g4670(.A(n10462), .B(n10464), .S0(TM1), .Y(n10465));
NOR2X1   g4671(.A(n10465), .B(n5827), .Y(n8295));
AND2X1   g4672(.A(CRC_OUT_1_30), .B(TM0), .Y(n10467));
AOI21X1  g4673(.A0(n5539), .A1(DATA_0_30), .B0(n10467), .Y(n10468));
INVX1    g4674(.A(WX10831), .Y(n10469));
MX2X1    g4675(.A(n10469), .B(n9899), .S0(n5539), .Y(n10470));
MX2X1    g4676(.A(n10468), .B(n10470), .S0(TM1), .Y(n10471));
NOR2X1   g4677(.A(n10471), .B(n5827), .Y(n8300));
AND2X1   g4678(.A(CRC_OUT_1_29), .B(TM0), .Y(n10473));
AOI21X1  g4679(.A0(n5539), .A1(DATA_0_29), .B0(n10473), .Y(n10474));
INVX1    g4680(.A(WX10833), .Y(n10475));
MX2X1    g4681(.A(n10475), .B(n9911), .S0(n5539), .Y(n10476));
MX2X1    g4682(.A(n10474), .B(n10476), .S0(TM1), .Y(n10477));
NOR2X1   g4683(.A(n10477), .B(n5827), .Y(n8305));
AND2X1   g4684(.A(CRC_OUT_1_28), .B(TM0), .Y(n10479));
AOI21X1  g4685(.A0(n5539), .A1(DATA_0_28), .B0(n10479), .Y(n10480));
INVX1    g4686(.A(WX10835), .Y(n10481));
MX2X1    g4687(.A(n10481), .B(n9923), .S0(n5539), .Y(n10482));
MX2X1    g4688(.A(n10480), .B(n10482), .S0(TM1), .Y(n10483));
NOR2X1   g4689(.A(n10483), .B(n5827), .Y(n8310));
AND2X1   g4690(.A(CRC_OUT_1_27), .B(TM0), .Y(n10485));
AOI21X1  g4691(.A0(n5539), .A1(DATA_0_27), .B0(n10485), .Y(n10486));
INVX1    g4692(.A(WX10837), .Y(n10487));
MX2X1    g4693(.A(n10487), .B(n9935), .S0(n5539), .Y(n10488));
MX2X1    g4694(.A(n10486), .B(n10488), .S0(TM1), .Y(n10489));
NOR2X1   g4695(.A(n10489), .B(n5827), .Y(n8315));
AND2X1   g4696(.A(CRC_OUT_1_26), .B(TM0), .Y(n10491));
AOI21X1  g4697(.A0(n5539), .A1(DATA_0_26), .B0(n10491), .Y(n10492));
INVX1    g4698(.A(WX10839), .Y(n10493));
MX2X1    g4699(.A(n10493), .B(n9947), .S0(n5539), .Y(n10494));
MX2X1    g4700(.A(n10492), .B(n10494), .S0(TM1), .Y(n10495));
NOR2X1   g4701(.A(n10495), .B(n5827), .Y(n8320));
AND2X1   g4702(.A(CRC_OUT_1_25), .B(TM0), .Y(n10497));
AOI21X1  g4703(.A0(n5539), .A1(DATA_0_25), .B0(n10497), .Y(n10498));
INVX1    g4704(.A(WX10841), .Y(n10499));
MX2X1    g4705(.A(n10499), .B(n9959), .S0(n5539), .Y(n10500));
MX2X1    g4706(.A(n10498), .B(n10500), .S0(TM1), .Y(n10501));
NOR2X1   g4707(.A(n10501), .B(n5827), .Y(n8325));
AND2X1   g4708(.A(CRC_OUT_1_24), .B(TM0), .Y(n10503));
AOI21X1  g4709(.A0(n5539), .A1(DATA_0_24), .B0(n10503), .Y(n10504));
INVX1    g4710(.A(WX10843), .Y(n10505));
MX2X1    g4711(.A(n10505), .B(n9971), .S0(n5539), .Y(n10506));
MX2X1    g4712(.A(n10504), .B(n10506), .S0(TM1), .Y(n10507));
NOR2X1   g4713(.A(n10507), .B(n5827), .Y(n8330));
AND2X1   g4714(.A(CRC_OUT_1_23), .B(TM0), .Y(n10509));
AOI21X1  g4715(.A0(n5539), .A1(DATA_0_23), .B0(n10509), .Y(n10510));
INVX1    g4716(.A(WX10845), .Y(n10511));
MX2X1    g4717(.A(n10511), .B(n9983), .S0(n5539), .Y(n10512));
MX2X1    g4718(.A(n10510), .B(n10512), .S0(TM1), .Y(n10513));
NOR2X1   g4719(.A(n10513), .B(n5827), .Y(n8335));
AND2X1   g4720(.A(CRC_OUT_1_22), .B(TM0), .Y(n10515));
AOI21X1  g4721(.A0(n5539), .A1(DATA_0_22), .B0(n10515), .Y(n10516));
INVX1    g4722(.A(WX10847), .Y(n10517));
MX2X1    g4723(.A(n10517), .B(n9995), .S0(n5539), .Y(n10518));
MX2X1    g4724(.A(n10516), .B(n10518), .S0(TM1), .Y(n10519));
NOR2X1   g4725(.A(n10519), .B(n5827), .Y(n8340));
AND2X1   g4726(.A(CRC_OUT_1_21), .B(TM0), .Y(n10521));
AOI21X1  g4727(.A0(n5539), .A1(DATA_0_21), .B0(n10521), .Y(n10522));
INVX1    g4728(.A(WX10849), .Y(n10523));
MX2X1    g4729(.A(n10523), .B(n10007), .S0(n5539), .Y(n10524));
MX2X1    g4730(.A(n10522), .B(n10524), .S0(TM1), .Y(n10525));
NOR2X1   g4731(.A(n10525), .B(n5827), .Y(n8345));
AND2X1   g4732(.A(CRC_OUT_1_20), .B(TM0), .Y(n10527));
AOI21X1  g4733(.A0(n5539), .A1(DATA_0_20), .B0(n10527), .Y(n10528));
INVX1    g4734(.A(WX10851), .Y(n10529));
MX2X1    g4735(.A(n10529), .B(n10019), .S0(n5539), .Y(n10530));
MX2X1    g4736(.A(n10528), .B(n10530), .S0(TM1), .Y(n10531));
NOR2X1   g4737(.A(n10531), .B(n5827), .Y(n8350));
AND2X1   g4738(.A(CRC_OUT_1_19), .B(TM0), .Y(n10533));
AOI21X1  g4739(.A0(n5539), .A1(DATA_0_19), .B0(n10533), .Y(n10534));
INVX1    g4740(.A(WX10853), .Y(n10535));
MX2X1    g4741(.A(n10535), .B(n10031), .S0(n5539), .Y(n10536));
MX2X1    g4742(.A(n10534), .B(n10536), .S0(TM1), .Y(n10537));
NOR2X1   g4743(.A(n10537), .B(n5827), .Y(n8355));
AND2X1   g4744(.A(CRC_OUT_1_18), .B(TM0), .Y(n10539));
AOI21X1  g4745(.A0(n5539), .A1(DATA_0_18), .B0(n10539), .Y(n10540));
INVX1    g4746(.A(WX10855), .Y(n10541));
MX2X1    g4747(.A(n10541), .B(n10043), .S0(n5539), .Y(n10542));
MX2X1    g4748(.A(n10540), .B(n10542), .S0(TM1), .Y(n10543));
NOR2X1   g4749(.A(n10543), .B(n5827), .Y(n8360));
AND2X1   g4750(.A(CRC_OUT_1_17), .B(TM0), .Y(n10545));
AOI21X1  g4751(.A0(n5539), .A1(DATA_0_17), .B0(n10545), .Y(n10546));
INVX1    g4752(.A(WX10857), .Y(n10547));
MX2X1    g4753(.A(n10547), .B(n10055), .S0(n5539), .Y(n10548));
MX2X1    g4754(.A(n10546), .B(n10548), .S0(TM1), .Y(n10549));
NOR2X1   g4755(.A(n10549), .B(n5827), .Y(n8365));
AND2X1   g4756(.A(CRC_OUT_1_16), .B(TM0), .Y(n10551));
AOI21X1  g4757(.A0(n5539), .A1(DATA_0_16), .B0(n10551), .Y(n10552));
INVX1    g4758(.A(WX10859), .Y(n10553));
MX2X1    g4759(.A(n10553), .B(n10067), .S0(n5539), .Y(n10554));
MX2X1    g4760(.A(n10552), .B(n10554), .S0(TM1), .Y(n10555));
NOR2X1   g4761(.A(n10555), .B(n5827), .Y(n8370));
AND2X1   g4762(.A(CRC_OUT_1_15), .B(TM0), .Y(n10557));
AOI21X1  g4763(.A0(n5539), .A1(DATA_0_15), .B0(n10557), .Y(n10558));
INVX1    g4764(.A(WX10861), .Y(n10559));
MX2X1    g4765(.A(n10559), .B(n10079), .S0(n5539), .Y(n10560));
MX2X1    g4766(.A(n10558), .B(n10560), .S0(TM1), .Y(n10561));
NOR2X1   g4767(.A(n10561), .B(n5827), .Y(n8375));
AND2X1   g4768(.A(CRC_OUT_1_14), .B(TM0), .Y(n10563));
AOI21X1  g4769(.A0(n5539), .A1(DATA_0_14), .B0(n10563), .Y(n10564));
INVX1    g4770(.A(WX10863), .Y(n10565));
MX2X1    g4771(.A(n10565), .B(n10091), .S0(n5539), .Y(n10566));
MX2X1    g4772(.A(n10564), .B(n10566), .S0(TM1), .Y(n10567));
NOR2X1   g4773(.A(n10567), .B(n5827), .Y(n8380));
AND2X1   g4774(.A(CRC_OUT_1_13), .B(TM0), .Y(n10569));
AOI21X1  g4775(.A0(n5539), .A1(DATA_0_13), .B0(n10569), .Y(n10570));
INVX1    g4776(.A(WX10865), .Y(n10571));
MX2X1    g4777(.A(n10571), .B(n10103), .S0(n5539), .Y(n10572));
MX2X1    g4778(.A(n10570), .B(n10572), .S0(TM1), .Y(n10573));
NOR2X1   g4779(.A(n10573), .B(n5827), .Y(n8385));
AND2X1   g4780(.A(CRC_OUT_1_12), .B(TM0), .Y(n10575));
AOI21X1  g4781(.A0(n5539), .A1(DATA_0_12), .B0(n10575), .Y(n10576));
INVX1    g4782(.A(WX10867), .Y(n10577));
MX2X1    g4783(.A(n10577), .B(n10115), .S0(n5539), .Y(n10578));
MX2X1    g4784(.A(n10576), .B(n10578), .S0(TM1), .Y(n10579));
NOR2X1   g4785(.A(n10579), .B(n5827), .Y(n8390));
AND2X1   g4786(.A(CRC_OUT_1_11), .B(TM0), .Y(n10581));
AOI21X1  g4787(.A0(n5539), .A1(DATA_0_11), .B0(n10581), .Y(n10582));
INVX1    g4788(.A(WX10869), .Y(n10583));
MX2X1    g4789(.A(n10583), .B(n10127), .S0(n5539), .Y(n10584));
MX2X1    g4790(.A(n10582), .B(n10584), .S0(TM1), .Y(n10585));
NOR2X1   g4791(.A(n10585), .B(n5827), .Y(n8395));
AND2X1   g4792(.A(CRC_OUT_1_10), .B(TM0), .Y(n10587));
AOI21X1  g4793(.A0(n5539), .A1(DATA_0_10), .B0(n10587), .Y(n10588));
INVX1    g4794(.A(WX10871), .Y(n10589));
MX2X1    g4795(.A(n10589), .B(n10139), .S0(n5539), .Y(n10590));
MX2X1    g4796(.A(n10588), .B(n10590), .S0(TM1), .Y(n10591));
NOR2X1   g4797(.A(n10591), .B(n5827), .Y(n8400));
AND2X1   g4798(.A(CRC_OUT_1_9), .B(TM0), .Y(n10593));
AOI21X1  g4799(.A0(n5539), .A1(DATA_0_9), .B0(n10593), .Y(n10594));
INVX1    g4800(.A(WX10873), .Y(n10595));
MX2X1    g4801(.A(n10595), .B(n10151), .S0(n5539), .Y(n10596));
MX2X1    g4802(.A(n10594), .B(n10596), .S0(TM1), .Y(n10597));
NOR2X1   g4803(.A(n10597), .B(n5827), .Y(n8405));
AND2X1   g4804(.A(CRC_OUT_1_8), .B(TM0), .Y(n10599));
AOI21X1  g4805(.A0(n5539), .A1(DATA_0_8), .B0(n10599), .Y(n10600));
INVX1    g4806(.A(WX10875), .Y(n10601));
MX2X1    g4807(.A(n10601), .B(n10163), .S0(n5539), .Y(n10602));
MX2X1    g4808(.A(n10600), .B(n10602), .S0(TM1), .Y(n10603));
NOR2X1   g4809(.A(n10603), .B(n5827), .Y(n8410));
AND2X1   g4810(.A(CRC_OUT_1_7), .B(TM0), .Y(n10605));
AOI21X1  g4811(.A0(n5539), .A1(DATA_0_7), .B0(n10605), .Y(n10606));
INVX1    g4812(.A(WX10877), .Y(n10607));
MX2X1    g4813(.A(n10607), .B(n10175), .S0(n5539), .Y(n10608));
MX2X1    g4814(.A(n10606), .B(n10608), .S0(TM1), .Y(n10609));
NOR2X1   g4815(.A(n10609), .B(n5827), .Y(n8415));
AND2X1   g4816(.A(CRC_OUT_1_6), .B(TM0), .Y(n10611));
AOI21X1  g4817(.A0(n5539), .A1(DATA_0_6), .B0(n10611), .Y(n10612));
INVX1    g4818(.A(WX10879), .Y(n10613));
MX2X1    g4819(.A(n10613), .B(n10187), .S0(n5539), .Y(n10614));
MX2X1    g4820(.A(n10612), .B(n10614), .S0(TM1), .Y(n10615));
NOR2X1   g4821(.A(n10615), .B(n5827), .Y(n8420));
AND2X1   g4822(.A(CRC_OUT_1_5), .B(TM0), .Y(n10617));
AOI21X1  g4823(.A0(n5539), .A1(DATA_0_5), .B0(n10617), .Y(n10618));
INVX1    g4824(.A(WX10881), .Y(n10619));
MX2X1    g4825(.A(n10619), .B(n10199), .S0(n5539), .Y(n10620));
MX2X1    g4826(.A(n10618), .B(n10620), .S0(TM1), .Y(n10621));
NOR2X1   g4827(.A(n10621), .B(n5827), .Y(n8425));
AND2X1   g4828(.A(CRC_OUT_1_4), .B(TM0), .Y(n10623));
AOI21X1  g4829(.A0(n5539), .A1(DATA_0_4), .B0(n10623), .Y(n10624));
INVX1    g4830(.A(WX10883), .Y(n10625));
MX2X1    g4831(.A(n10625), .B(n10211), .S0(n5539), .Y(n10626));
MX2X1    g4832(.A(n10624), .B(n10626), .S0(TM1), .Y(n10627));
NOR2X1   g4833(.A(n10627), .B(n5827), .Y(n8430));
AND2X1   g4834(.A(CRC_OUT_1_3), .B(TM0), .Y(n10629));
AOI21X1  g4835(.A0(n5539), .A1(DATA_0_3), .B0(n10629), .Y(n10630));
INVX1    g4836(.A(WX10885), .Y(n10631));
MX2X1    g4837(.A(n10631), .B(n10223), .S0(n5539), .Y(n10632));
MX2X1    g4838(.A(n10630), .B(n10632), .S0(TM1), .Y(n10633));
NOR2X1   g4839(.A(n10633), .B(n5827), .Y(n8435));
AND2X1   g4840(.A(CRC_OUT_1_2), .B(TM0), .Y(n10635));
AOI21X1  g4841(.A0(n5539), .A1(DATA_0_2), .B0(n10635), .Y(n10636));
INVX1    g4842(.A(WX10887), .Y(n10637));
MX2X1    g4843(.A(n10637), .B(n10235), .S0(n5539), .Y(n10638));
MX2X1    g4844(.A(n10636), .B(n10638), .S0(TM1), .Y(n10639));
NOR2X1   g4845(.A(n10639), .B(n5827), .Y(n8440));
AND2X1   g4846(.A(CRC_OUT_1_1), .B(TM0), .Y(n10641));
AOI21X1  g4847(.A0(n5539), .A1(DATA_0_1), .B0(n10641), .Y(n10642));
INVX1    g4848(.A(WX10889), .Y(n10643));
MX2X1    g4849(.A(n10643), .B(n10247), .S0(n5539), .Y(n10644));
MX2X1    g4850(.A(n10642), .B(n10644), .S0(TM1), .Y(n10645));
NOR2X1   g4851(.A(n10645), .B(n5827), .Y(n8445));
AND2X1   g4852(.A(CRC_OUT_1_0), .B(TM0), .Y(n10647));
AOI21X1  g4853(.A0(n5539), .A1(DATA_0_0), .B0(n10647), .Y(n10648));
INVX1    g4854(.A(WX10891), .Y(n10649));
MX2X1    g4855(.A(n10649), .B(n10259), .S0(n5539), .Y(n10650));
MX2X1    g4856(.A(n10648), .B(n10650), .S0(TM1), .Y(n10651));
NOR2X1   g4857(.A(n10651), .B(n5827), .Y(n8450));
AND2X1   g4858(.A(WX10989), .B(RESET), .Y(n8455));
AND2X1   g4859(.A(WX10991), .B(RESET), .Y(n8460));
AND2X1   g4860(.A(WX10993), .B(RESET), .Y(n8465));
AND2X1   g4861(.A(WX10995), .B(RESET), .Y(n8470));
AND2X1   g4862(.A(WX10997), .B(RESET), .Y(n8475));
AND2X1   g4863(.A(WX10999), .B(RESET), .Y(n8480));
AND2X1   g4864(.A(WX11001), .B(RESET), .Y(n8485));
AND2X1   g4865(.A(WX11003), .B(RESET), .Y(n8490));
AND2X1   g4866(.A(WX11005), .B(RESET), .Y(n8495));
AND2X1   g4867(.A(WX11007), .B(RESET), .Y(n8500));
AND2X1   g4868(.A(WX11009), .B(RESET), .Y(n8505));
AND2X1   g4869(.A(WX11011), .B(RESET), .Y(n8510));
AND2X1   g4870(.A(WX11013), .B(RESET), .Y(n8515));
AND2X1   g4871(.A(WX11015), .B(RESET), .Y(n8520));
AND2X1   g4872(.A(WX11017), .B(RESET), .Y(n8525));
AND2X1   g4873(.A(WX11019), .B(RESET), .Y(n8530));
AND2X1   g4874(.A(WX11021), .B(RESET), .Y(n8535));
AND2X1   g4875(.A(WX11023), .B(RESET), .Y(n8540));
AND2X1   g4876(.A(WX11025), .B(RESET), .Y(n8545));
AND2X1   g4877(.A(WX11027), .B(RESET), .Y(n8550));
AND2X1   g4878(.A(WX11029), .B(RESET), .Y(n8555));
AND2X1   g4879(.A(WX11031), .B(RESET), .Y(n8560));
AND2X1   g4880(.A(WX11033), .B(RESET), .Y(n8565));
AND2X1   g4881(.A(WX11035), .B(RESET), .Y(n8570));
AND2X1   g4882(.A(WX11037), .B(RESET), .Y(n8575));
AND2X1   g4883(.A(WX11039), .B(RESET), .Y(n8580));
AND2X1   g4884(.A(WX11041), .B(RESET), .Y(n8585));
AND2X1   g4885(.A(WX11043), .B(RESET), .Y(n8590));
AND2X1   g4886(.A(WX11045), .B(RESET), .Y(n8595));
AND2X1   g4887(.A(WX11047), .B(RESET), .Y(n8600));
AND2X1   g4888(.A(WX11049), .B(RESET), .Y(n8605));
AND2X1   g4889(.A(WX11051), .B(RESET), .Y(n8610));
AND2X1   g4890(.A(WX11053), .B(RESET), .Y(n8615));
AND2X1   g4891(.A(WX11055), .B(RESET), .Y(n8620));
AND2X1   g4892(.A(WX11057), .B(RESET), .Y(n8625));
AND2X1   g4893(.A(WX11059), .B(RESET), .Y(n8630));
AND2X1   g4894(.A(WX11061), .B(RESET), .Y(n8635));
AND2X1   g4895(.A(WX11063), .B(RESET), .Y(n8640));
AND2X1   g4896(.A(WX11065), .B(RESET), .Y(n8645));
AND2X1   g4897(.A(WX11067), .B(RESET), .Y(n8650));
AND2X1   g4898(.A(WX11069), .B(RESET), .Y(n8655));
AND2X1   g4899(.A(WX11071), .B(RESET), .Y(n8660));
AND2X1   g4900(.A(WX11073), .B(RESET), .Y(n8665));
AND2X1   g4901(.A(WX11075), .B(RESET), .Y(n8670));
AND2X1   g4902(.A(WX11077), .B(RESET), .Y(n8675));
AND2X1   g4903(.A(WX11079), .B(RESET), .Y(n8680));
AND2X1   g4904(.A(WX11081), .B(RESET), .Y(n8685));
AND2X1   g4905(.A(WX11083), .B(RESET), .Y(n8690));
AND2X1   g4906(.A(WX11085), .B(RESET), .Y(n8695));
AND2X1   g4907(.A(WX11087), .B(RESET), .Y(n8700));
AND2X1   g4908(.A(WX11089), .B(RESET), .Y(n8705));
AND2X1   g4909(.A(WX11091), .B(RESET), .Y(n8710));
AND2X1   g4910(.A(WX11093), .B(RESET), .Y(n8715));
AND2X1   g4911(.A(WX11095), .B(RESET), .Y(n8720));
AND2X1   g4912(.A(WX11097), .B(RESET), .Y(n8725));
AND2X1   g4913(.A(WX11099), .B(RESET), .Y(n8730));
AND2X1   g4914(.A(WX11101), .B(RESET), .Y(n8735));
AND2X1   g4915(.A(WX11103), .B(RESET), .Y(n8740));
AND2X1   g4916(.A(WX11105), .B(RESET), .Y(n8745));
AND2X1   g4917(.A(WX11107), .B(RESET), .Y(n8750));
AND2X1   g4918(.A(WX11109), .B(RESET), .Y(n8755));
AND2X1   g4919(.A(WX11111), .B(RESET), .Y(n8760));
AND2X1   g4920(.A(WX11113), .B(RESET), .Y(n8765));
AND2X1   g4921(.A(WX11115), .B(RESET), .Y(n8770));
AND2X1   g4922(.A(WX11117), .B(RESET), .Y(n8775));
AND2X1   g4923(.A(WX11119), .B(RESET), .Y(n8780));
AND2X1   g4924(.A(WX11121), .B(RESET), .Y(n8785));
AND2X1   g4925(.A(WX11123), .B(RESET), .Y(n8790));
AND2X1   g4926(.A(WX11125), .B(RESET), .Y(n8795));
AND2X1   g4927(.A(WX11127), .B(RESET), .Y(n8800));
AND2X1   g4928(.A(WX11129), .B(RESET), .Y(n8805));
AND2X1   g4929(.A(WX11131), .B(RESET), .Y(n8810));
AND2X1   g4930(.A(WX11133), .B(RESET), .Y(n8815));
AND2X1   g4931(.A(WX11135), .B(RESET), .Y(n8820));
AND2X1   g4932(.A(WX11137), .B(RESET), .Y(n8825));
AND2X1   g4933(.A(WX11139), .B(RESET), .Y(n8830));
AND2X1   g4934(.A(WX11141), .B(RESET), .Y(n8835));
AND2X1   g4935(.A(WX11143), .B(RESET), .Y(n8840));
AND2X1   g4936(.A(WX11145), .B(RESET), .Y(n8845));
AND2X1   g4937(.A(WX11147), .B(RESET), .Y(n8850));
AND2X1   g4938(.A(WX11149), .B(RESET), .Y(n8855));
AND2X1   g4939(.A(WX11151), .B(RESET), .Y(n8860));
AND2X1   g4940(.A(WX11153), .B(RESET), .Y(n8865));
AND2X1   g4941(.A(WX11155), .B(RESET), .Y(n8870));
AND2X1   g4942(.A(WX11157), .B(RESET), .Y(n8875));
AND2X1   g4943(.A(WX11159), .B(RESET), .Y(n8880));
AND2X1   g4944(.A(WX11161), .B(RESET), .Y(n8885));
AND2X1   g4945(.A(WX11163), .B(RESET), .Y(n8890));
AND2X1   g4946(.A(WX11165), .B(RESET), .Y(n8895));
AND2X1   g4947(.A(WX11167), .B(RESET), .Y(n8900));
AND2X1   g4948(.A(WX11169), .B(RESET), .Y(n8905));
AND2X1   g4949(.A(WX11171), .B(RESET), .Y(n8910));
AND2X1   g4950(.A(WX11173), .B(RESET), .Y(n8915));
AND2X1   g4951(.A(WX11175), .B(RESET), .Y(n8920));
AND2X1   g4952(.A(WX11177), .B(RESET), .Y(n8925));
AND2X1   g4953(.A(WX11179), .B(RESET), .Y(n8930));
XOR2X1   g4954(.A(CRC_OUT_1_31), .B(WX11243), .Y(n10749));
NOR2X1   g4955(.A(n10749), .B(n5827), .Y(CRC_OUT_1_0));
XOR2X1   g4956(.A(CRC_OUT_1_0), .B(WX11241), .Y(n10751));
NOR2X1   g4957(.A(n10751), .B(n5827), .Y(CRC_OUT_1_1));
XOR2X1   g4958(.A(CRC_OUT_1_1), .B(WX11239), .Y(n10753));
NOR2X1   g4959(.A(n10753), .B(n5827), .Y(CRC_OUT_1_2));
XOR2X1   g4960(.A(CRC_OUT_1_2), .B(WX11237), .Y(n10755));
NOR2X1   g4961(.A(n10755), .B(n5827), .Y(CRC_OUT_1_3));
XOR2X1   g4962(.A(CRC_OUT_1_31), .B(WX11235), .Y(n10757));
XOR2X1   g4963(.A(n10757), .B(CRC_OUT_1_3), .Y(n10758));
NOR2X1   g4964(.A(n10758), .B(n5827), .Y(CRC_OUT_1_4));
XOR2X1   g4965(.A(CRC_OUT_1_4), .B(WX11233), .Y(n10760));
NOR2X1   g4966(.A(n10760), .B(n5827), .Y(CRC_OUT_1_5));
XOR2X1   g4967(.A(CRC_OUT_1_5), .B(WX11231), .Y(n10762));
NOR2X1   g4968(.A(n10762), .B(n5827), .Y(CRC_OUT_1_6));
XOR2X1   g4969(.A(CRC_OUT_1_6), .B(WX11229), .Y(n10764));
NOR2X1   g4970(.A(n10764), .B(n5827), .Y(CRC_OUT_1_7));
XOR2X1   g4971(.A(CRC_OUT_1_7), .B(WX11227), .Y(n10766));
NOR2X1   g4972(.A(n10766), .B(n5827), .Y(CRC_OUT_1_8));
XOR2X1   g4973(.A(CRC_OUT_1_8), .B(WX11225), .Y(n10768));
NOR2X1   g4974(.A(n10768), .B(n5827), .Y(CRC_OUT_1_9));
XOR2X1   g4975(.A(CRC_OUT_1_9), .B(WX11223), .Y(n10770));
NOR2X1   g4976(.A(n10770), .B(n5827), .Y(CRC_OUT_1_10));
XOR2X1   g4977(.A(CRC_OUT_1_31), .B(WX11221), .Y(n10772));
XOR2X1   g4978(.A(n10772), .B(CRC_OUT_1_10), .Y(n10773));
NOR2X1   g4979(.A(n10773), .B(n5827), .Y(CRC_OUT_1_11));
XOR2X1   g4980(.A(CRC_OUT_1_11), .B(WX11219), .Y(n10775));
NOR2X1   g4981(.A(n10775), .B(n5827), .Y(CRC_OUT_1_12));
XOR2X1   g4982(.A(CRC_OUT_1_12), .B(WX11217), .Y(n10777));
NOR2X1   g4983(.A(n10777), .B(n5827), .Y(CRC_OUT_1_13));
XOR2X1   g4984(.A(CRC_OUT_1_13), .B(WX11215), .Y(n10779));
NOR2X1   g4985(.A(n10779), .B(n5827), .Y(CRC_OUT_1_14));
XOR2X1   g4986(.A(CRC_OUT_1_14), .B(WX11213), .Y(n10781));
NOR2X1   g4987(.A(n10781), .B(n5827), .Y(CRC_OUT_1_15));
XOR2X1   g4988(.A(CRC_OUT_1_31), .B(WX11211), .Y(n10783));
XOR2X1   g4989(.A(n10783), .B(CRC_OUT_1_15), .Y(n10784));
NOR2X1   g4990(.A(n10784), .B(n5827), .Y(CRC_OUT_1_16));
XOR2X1   g4991(.A(CRC_OUT_1_16), .B(WX11209), .Y(n10786));
NOR2X1   g4992(.A(n10786), .B(n5827), .Y(CRC_OUT_1_17));
XOR2X1   g4993(.A(CRC_OUT_1_17), .B(WX11207), .Y(n10788));
NOR2X1   g4994(.A(n10788), .B(n5827), .Y(CRC_OUT_1_18));
XOR2X1   g4995(.A(CRC_OUT_1_18), .B(WX11205), .Y(n10790));
NOR2X1   g4996(.A(n10790), .B(n5827), .Y(CRC_OUT_1_19));
XOR2X1   g4997(.A(CRC_OUT_1_19), .B(WX11203), .Y(n10792));
NOR2X1   g4998(.A(n10792), .B(n5827), .Y(CRC_OUT_1_20));
XOR2X1   g4999(.A(CRC_OUT_1_20), .B(WX11201), .Y(n10794));
NOR2X1   g5000(.A(n10794), .B(n5827), .Y(CRC_OUT_1_21));
XOR2X1   g5001(.A(CRC_OUT_1_21), .B(WX11199), .Y(n10796));
NOR2X1   g5002(.A(n10796), .B(n5827), .Y(CRC_OUT_1_22));
XOR2X1   g5003(.A(CRC_OUT_1_22), .B(WX11197), .Y(n10798));
NOR2X1   g5004(.A(n10798), .B(n5827), .Y(CRC_OUT_1_23));
XOR2X1   g5005(.A(CRC_OUT_1_23), .B(WX11195), .Y(n10800));
NOR2X1   g5006(.A(n10800), .B(n5827), .Y(CRC_OUT_1_24));
XOR2X1   g5007(.A(CRC_OUT_1_24), .B(WX11193), .Y(n10802));
NOR2X1   g5008(.A(n10802), .B(n5827), .Y(CRC_OUT_1_25));
XOR2X1   g5009(.A(CRC_OUT_1_25), .B(WX11191), .Y(n10804));
NOR2X1   g5010(.A(n10804), .B(n5827), .Y(CRC_OUT_1_26));
XOR2X1   g5011(.A(CRC_OUT_1_26), .B(WX11189), .Y(n10806));
NOR2X1   g5012(.A(n10806), .B(n5827), .Y(CRC_OUT_1_27));
XOR2X1   g5013(.A(CRC_OUT_1_27), .B(WX11187), .Y(n10808));
NOR2X1   g5014(.A(n10808), .B(n5827), .Y(CRC_OUT_1_28));
XOR2X1   g5015(.A(CRC_OUT_1_28), .B(WX11185), .Y(n10810));
NOR2X1   g5016(.A(n10810), .B(n5827), .Y(CRC_OUT_1_29));
XOR2X1   g5017(.A(CRC_OUT_1_29), .B(WX11183), .Y(n10812));
NOR2X1   g5018(.A(n10812), .B(n5827), .Y(CRC_OUT_1_30));
XOR2X1   g5019(.A(CRC_OUT_1_30), .B(WX11181), .Y(n10814));
NOR2X1   g5020(.A(n10814), .B(n5827), .Y(CRC_OUT_1_31));
endmodule
